library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs: in std_logic_vector(1023 downto 0);
        outputs: out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs: std_logic_vector(7679 downto 0);
    signal layer1_outputs: std_logic_vector(7679 downto 0);
    signal layer2_outputs: std_logic_vector(7679 downto 0);

begin
    layer0_outputs(0) <= a and not b;
    layer0_outputs(1) <= not a;
    layer0_outputs(2) <= a or b;
    layer0_outputs(3) <= a or b;
    layer0_outputs(4) <= not (a or b);
    layer0_outputs(5) <= a or b;
    layer0_outputs(6) <= a and b;
    layer0_outputs(7) <= a or b;
    layer0_outputs(8) <= not b;
    layer0_outputs(9) <= not (a or b);
    layer0_outputs(10) <= a and not b;
    layer0_outputs(11) <= not (a or b);
    layer0_outputs(12) <= a xor b;
    layer0_outputs(13) <= a and not b;
    layer0_outputs(14) <= a;
    layer0_outputs(15) <= a xor b;
    layer0_outputs(16) <= a or b;
    layer0_outputs(17) <= a;
    layer0_outputs(18) <= not (a xor b);
    layer0_outputs(19) <= not a;
    layer0_outputs(20) <= not (a or b);
    layer0_outputs(21) <= not b;
    layer0_outputs(22) <= a;
    layer0_outputs(23) <= a or b;
    layer0_outputs(24) <= not b or a;
    layer0_outputs(25) <= not (a xor b);
    layer0_outputs(26) <= b and not a;
    layer0_outputs(27) <= not b;
    layer0_outputs(28) <= not (a or b);
    layer0_outputs(29) <= b;
    layer0_outputs(30) <= a;
    layer0_outputs(31) <= 1'b0;
    layer0_outputs(32) <= not (a or b);
    layer0_outputs(33) <= a or b;
    layer0_outputs(34) <= not b;
    layer0_outputs(35) <= not (a and b);
    layer0_outputs(36) <= not (a xor b);
    layer0_outputs(37) <= a and not b;
    layer0_outputs(38) <= not a or b;
    layer0_outputs(39) <= a or b;
    layer0_outputs(40) <= a xor b;
    layer0_outputs(41) <= not (a or b);
    layer0_outputs(42) <= not b;
    layer0_outputs(43) <= not a;
    layer0_outputs(44) <= not a;
    layer0_outputs(45) <= b and not a;
    layer0_outputs(46) <= a or b;
    layer0_outputs(47) <= not b or a;
    layer0_outputs(48) <= not (a or b);
    layer0_outputs(49) <= b and not a;
    layer0_outputs(50) <= not (a xor b);
    layer0_outputs(51) <= not b or a;
    layer0_outputs(52) <= 1'b0;
    layer0_outputs(53) <= a or b;
    layer0_outputs(54) <= a and not b;
    layer0_outputs(55) <= a xor b;
    layer0_outputs(56) <= a or b;
    layer0_outputs(57) <= not (a and b);
    layer0_outputs(58) <= a and b;
    layer0_outputs(59) <= b;
    layer0_outputs(60) <= 1'b1;
    layer0_outputs(61) <= 1'b1;
    layer0_outputs(62) <= b and not a;
    layer0_outputs(63) <= not (a or b);
    layer0_outputs(64) <= not (a xor b);
    layer0_outputs(65) <= b;
    layer0_outputs(66) <= not a or b;
    layer0_outputs(67) <= not (a xor b);
    layer0_outputs(68) <= a xor b;
    layer0_outputs(69) <= b;
    layer0_outputs(70) <= not b or a;
    layer0_outputs(71) <= not (a xor b);
    layer0_outputs(72) <= a or b;
    layer0_outputs(73) <= a and not b;
    layer0_outputs(74) <= 1'b1;
    layer0_outputs(75) <= not (a or b);
    layer0_outputs(76) <= not (a or b);
    layer0_outputs(77) <= a and not b;
    layer0_outputs(78) <= not (a xor b);
    layer0_outputs(79) <= not a or b;
    layer0_outputs(80) <= b;
    layer0_outputs(81) <= not (a or b);
    layer0_outputs(82) <= a or b;
    layer0_outputs(83) <= a xor b;
    layer0_outputs(84) <= a;
    layer0_outputs(85) <= not b;
    layer0_outputs(86) <= not b;
    layer0_outputs(87) <= not b;
    layer0_outputs(88) <= a;
    layer0_outputs(89) <= not (a and b);
    layer0_outputs(90) <= not (a xor b);
    layer0_outputs(91) <= a and b;
    layer0_outputs(92) <= b;
    layer0_outputs(93) <= b;
    layer0_outputs(94) <= a or b;
    layer0_outputs(95) <= a;
    layer0_outputs(96) <= not (a xor b);
    layer0_outputs(97) <= not (a or b);
    layer0_outputs(98) <= b and not a;
    layer0_outputs(99) <= a xor b;
    layer0_outputs(100) <= 1'b0;
    layer0_outputs(101) <= a xor b;
    layer0_outputs(102) <= not (a or b);
    layer0_outputs(103) <= a or b;
    layer0_outputs(104) <= a and not b;
    layer0_outputs(105) <= not a or b;
    layer0_outputs(106) <= b;
    layer0_outputs(107) <= a and not b;
    layer0_outputs(108) <= a and not b;
    layer0_outputs(109) <= not b or a;
    layer0_outputs(110) <= not a or b;
    layer0_outputs(111) <= not (a or b);
    layer0_outputs(112) <= not (a or b);
    layer0_outputs(113) <= a and not b;
    layer0_outputs(114) <= 1'b1;
    layer0_outputs(115) <= not a;
    layer0_outputs(116) <= not b;
    layer0_outputs(117) <= not (a xor b);
    layer0_outputs(118) <= a;
    layer0_outputs(119) <= a and not b;
    layer0_outputs(120) <= not a or b;
    layer0_outputs(121) <= not a;
    layer0_outputs(122) <= b and not a;
    layer0_outputs(123) <= a xor b;
    layer0_outputs(124) <= 1'b0;
    layer0_outputs(125) <= not (a xor b);
    layer0_outputs(126) <= not (a and b);
    layer0_outputs(127) <= not (a or b);
    layer0_outputs(128) <= a or b;
    layer0_outputs(129) <= not (a or b);
    layer0_outputs(130) <= not a;
    layer0_outputs(131) <= a or b;
    layer0_outputs(132) <= a or b;
    layer0_outputs(133) <= a;
    layer0_outputs(134) <= a and not b;
    layer0_outputs(135) <= not a;
    layer0_outputs(136) <= not b;
    layer0_outputs(137) <= a and not b;
    layer0_outputs(138) <= not b or a;
    layer0_outputs(139) <= not (a or b);
    layer0_outputs(140) <= b and not a;
    layer0_outputs(141) <= a and not b;
    layer0_outputs(142) <= not a;
    layer0_outputs(143) <= not b or a;
    layer0_outputs(144) <= a and b;
    layer0_outputs(145) <= a and b;
    layer0_outputs(146) <= a and not b;
    layer0_outputs(147) <= not b;
    layer0_outputs(148) <= b and not a;
    layer0_outputs(149) <= not (a xor b);
    layer0_outputs(150) <= not (a or b);
    layer0_outputs(151) <= not a;
    layer0_outputs(152) <= a and b;
    layer0_outputs(153) <= a and b;
    layer0_outputs(154) <= not b or a;
    layer0_outputs(155) <= not (a or b);
    layer0_outputs(156) <= not (a xor b);
    layer0_outputs(157) <= a or b;
    layer0_outputs(158) <= a or b;
    layer0_outputs(159) <= not b or a;
    layer0_outputs(160) <= not (a and b);
    layer0_outputs(161) <= a;
    layer0_outputs(162) <= b;
    layer0_outputs(163) <= b and not a;
    layer0_outputs(164) <= a;
    layer0_outputs(165) <= not b;
    layer0_outputs(166) <= b;
    layer0_outputs(167) <= a xor b;
    layer0_outputs(168) <= not a or b;
    layer0_outputs(169) <= not (a xor b);
    layer0_outputs(170) <= a or b;
    layer0_outputs(171) <= b and not a;
    layer0_outputs(172) <= not b;
    layer0_outputs(173) <= a or b;
    layer0_outputs(174) <= b and not a;
    layer0_outputs(175) <= not (a or b);
    layer0_outputs(176) <= not (a xor b);
    layer0_outputs(177) <= a or b;
    layer0_outputs(178) <= not b or a;
    layer0_outputs(179) <= 1'b1;
    layer0_outputs(180) <= not a;
    layer0_outputs(181) <= b and not a;
    layer0_outputs(182) <= not b;
    layer0_outputs(183) <= not a;
    layer0_outputs(184) <= a and not b;
    layer0_outputs(185) <= b and not a;
    layer0_outputs(186) <= not b;
    layer0_outputs(187) <= a and not b;
    layer0_outputs(188) <= not a or b;
    layer0_outputs(189) <= b;
    layer0_outputs(190) <= not b or a;
    layer0_outputs(191) <= not (a or b);
    layer0_outputs(192) <= not b or a;
    layer0_outputs(193) <= a;
    layer0_outputs(194) <= not (a or b);
    layer0_outputs(195) <= 1'b1;
    layer0_outputs(196) <= not b;
    layer0_outputs(197) <= a and not b;
    layer0_outputs(198) <= not b or a;
    layer0_outputs(199) <= a or b;
    layer0_outputs(200) <= not (a xor b);
    layer0_outputs(201) <= a xor b;
    layer0_outputs(202) <= 1'b1;
    layer0_outputs(203) <= not a;
    layer0_outputs(204) <= a xor b;
    layer0_outputs(205) <= not (a xor b);
    layer0_outputs(206) <= not a;
    layer0_outputs(207) <= a xor b;
    layer0_outputs(208) <= a and not b;
    layer0_outputs(209) <= b;
    layer0_outputs(210) <= a;
    layer0_outputs(211) <= 1'b1;
    layer0_outputs(212) <= 1'b1;
    layer0_outputs(213) <= not (a and b);
    layer0_outputs(214) <= not b;
    layer0_outputs(215) <= a and not b;
    layer0_outputs(216) <= b and not a;
    layer0_outputs(217) <= not b or a;
    layer0_outputs(218) <= not a or b;
    layer0_outputs(219) <= a;
    layer0_outputs(220) <= a;
    layer0_outputs(221) <= not a or b;
    layer0_outputs(222) <= not a or b;
    layer0_outputs(223) <= a and not b;
    layer0_outputs(224) <= a and b;
    layer0_outputs(225) <= not b;
    layer0_outputs(226) <= 1'b0;
    layer0_outputs(227) <= not b;
    layer0_outputs(228) <= a and not b;
    layer0_outputs(229) <= not (a or b);
    layer0_outputs(230) <= a and not b;
    layer0_outputs(231) <= not a;
    layer0_outputs(232) <= not a;
    layer0_outputs(233) <= not (a xor b);
    layer0_outputs(234) <= b and not a;
    layer0_outputs(235) <= b;
    layer0_outputs(236) <= a xor b;
    layer0_outputs(237) <= not b;
    layer0_outputs(238) <= not (a or b);
    layer0_outputs(239) <= not b;
    layer0_outputs(240) <= not b;
    layer0_outputs(241) <= a or b;
    layer0_outputs(242) <= b;
    layer0_outputs(243) <= not b;
    layer0_outputs(244) <= a xor b;
    layer0_outputs(245) <= a or b;
    layer0_outputs(246) <= not a;
    layer0_outputs(247) <= a or b;
    layer0_outputs(248) <= 1'b0;
    layer0_outputs(249) <= a;
    layer0_outputs(250) <= not (a or b);
    layer0_outputs(251) <= a or b;
    layer0_outputs(252) <= not (a or b);
    layer0_outputs(253) <= not (a xor b);
    layer0_outputs(254) <= a or b;
    layer0_outputs(255) <= a and not b;
    layer0_outputs(256) <= a and b;
    layer0_outputs(257) <= b and not a;
    layer0_outputs(258) <= b and not a;
    layer0_outputs(259) <= b;
    layer0_outputs(260) <= a xor b;
    layer0_outputs(261) <= not b;
    layer0_outputs(262) <= not a or b;
    layer0_outputs(263) <= a and not b;
    layer0_outputs(264) <= a and b;
    layer0_outputs(265) <= not (a or b);
    layer0_outputs(266) <= a and not b;
    layer0_outputs(267) <= a and b;
    layer0_outputs(268) <= b and not a;
    layer0_outputs(269) <= b;
    layer0_outputs(270) <= b and not a;
    layer0_outputs(271) <= not b;
    layer0_outputs(272) <= not b or a;
    layer0_outputs(273) <= not a or b;
    layer0_outputs(274) <= not a or b;
    layer0_outputs(275) <= a or b;
    layer0_outputs(276) <= not b;
    layer0_outputs(277) <= b;
    layer0_outputs(278) <= not b;
    layer0_outputs(279) <= not a;
    layer0_outputs(280) <= b;
    layer0_outputs(281) <= not (a or b);
    layer0_outputs(282) <= not b or a;
    layer0_outputs(283) <= a xor b;
    layer0_outputs(284) <= a and not b;
    layer0_outputs(285) <= a or b;
    layer0_outputs(286) <= not (a xor b);
    layer0_outputs(287) <= not a;
    layer0_outputs(288) <= a;
    layer0_outputs(289) <= not (a or b);
    layer0_outputs(290) <= a and not b;
    layer0_outputs(291) <= not b;
    layer0_outputs(292) <= not (a and b);
    layer0_outputs(293) <= b;
    layer0_outputs(294) <= not a;
    layer0_outputs(295) <= a xor b;
    layer0_outputs(296) <= not b or a;
    layer0_outputs(297) <= a;
    layer0_outputs(298) <= a;
    layer0_outputs(299) <= a or b;
    layer0_outputs(300) <= a xor b;
    layer0_outputs(301) <= a;
    layer0_outputs(302) <= 1'b0;
    layer0_outputs(303) <= b;
    layer0_outputs(304) <= not (a or b);
    layer0_outputs(305) <= b and not a;
    layer0_outputs(306) <= a or b;
    layer0_outputs(307) <= a and not b;
    layer0_outputs(308) <= not (a or b);
    layer0_outputs(309) <= a xor b;
    layer0_outputs(310) <= a;
    layer0_outputs(311) <= not a;
    layer0_outputs(312) <= not a or b;
    layer0_outputs(313) <= a or b;
    layer0_outputs(314) <= b;
    layer0_outputs(315) <= a;
    layer0_outputs(316) <= not a;
    layer0_outputs(317) <= not (a or b);
    layer0_outputs(318) <= 1'b0;
    layer0_outputs(319) <= not (a xor b);
    layer0_outputs(320) <= not (a and b);
    layer0_outputs(321) <= a and not b;
    layer0_outputs(322) <= not (a xor b);
    layer0_outputs(323) <= a and b;
    layer0_outputs(324) <= a or b;
    layer0_outputs(325) <= a or b;
    layer0_outputs(326) <= not a or b;
    layer0_outputs(327) <= not (a xor b);
    layer0_outputs(328) <= a and not b;
    layer0_outputs(329) <= not b;
    layer0_outputs(330) <= a;
    layer0_outputs(331) <= not (a and b);
    layer0_outputs(332) <= not (a xor b);
    layer0_outputs(333) <= a or b;
    layer0_outputs(334) <= a xor b;
    layer0_outputs(335) <= a or b;
    layer0_outputs(336) <= a;
    layer0_outputs(337) <= a;
    layer0_outputs(338) <= a;
    layer0_outputs(339) <= b;
    layer0_outputs(340) <= not (a or b);
    layer0_outputs(341) <= 1'b0;
    layer0_outputs(342) <= not a;
    layer0_outputs(343) <= a xor b;
    layer0_outputs(344) <= a or b;
    layer0_outputs(345) <= b and not a;
    layer0_outputs(346) <= not a;
    layer0_outputs(347) <= not b;
    layer0_outputs(348) <= not b or a;
    layer0_outputs(349) <= not b;
    layer0_outputs(350) <= b;
    layer0_outputs(351) <= not (a xor b);
    layer0_outputs(352) <= not b;
    layer0_outputs(353) <= not (a or b);
    layer0_outputs(354) <= not (a xor b);
    layer0_outputs(355) <= not (a or b);
    layer0_outputs(356) <= b and not a;
    layer0_outputs(357) <= b and not a;
    layer0_outputs(358) <= a and not b;
    layer0_outputs(359) <= a xor b;
    layer0_outputs(360) <= not a;
    layer0_outputs(361) <= a or b;
    layer0_outputs(362) <= not (a or b);
    layer0_outputs(363) <= not (a or b);
    layer0_outputs(364) <= a;
    layer0_outputs(365) <= b and not a;
    layer0_outputs(366) <= not (a and b);
    layer0_outputs(367) <= b and not a;
    layer0_outputs(368) <= not b or a;
    layer0_outputs(369) <= not (a xor b);
    layer0_outputs(370) <= not (a and b);
    layer0_outputs(371) <= a xor b;
    layer0_outputs(372) <= 1'b0;
    layer0_outputs(373) <= not a;
    layer0_outputs(374) <= not b;
    layer0_outputs(375) <= not b or a;
    layer0_outputs(376) <= not a;
    layer0_outputs(377) <= not (a xor b);
    layer0_outputs(378) <= not a or b;
    layer0_outputs(379) <= a or b;
    layer0_outputs(380) <= not (a or b);
    layer0_outputs(381) <= not b or a;
    layer0_outputs(382) <= 1'b1;
    layer0_outputs(383) <= not b or a;
    layer0_outputs(384) <= a xor b;
    layer0_outputs(385) <= not (a or b);
    layer0_outputs(386) <= b and not a;
    layer0_outputs(387) <= 1'b0;
    layer0_outputs(388) <= b;
    layer0_outputs(389) <= a;
    layer0_outputs(390) <= b and not a;
    layer0_outputs(391) <= a and not b;
    layer0_outputs(392) <= a xor b;
    layer0_outputs(393) <= not a or b;
    layer0_outputs(394) <= not (a or b);
    layer0_outputs(395) <= not (a or b);
    layer0_outputs(396) <= a or b;
    layer0_outputs(397) <= not a;
    layer0_outputs(398) <= b and not a;
    layer0_outputs(399) <= not (a or b);
    layer0_outputs(400) <= b and not a;
    layer0_outputs(401) <= not b or a;
    layer0_outputs(402) <= a xor b;
    layer0_outputs(403) <= b;
    layer0_outputs(404) <= b and not a;
    layer0_outputs(405) <= not a or b;
    layer0_outputs(406) <= not b;
    layer0_outputs(407) <= not (a xor b);
    layer0_outputs(408) <= not a;
    layer0_outputs(409) <= not b or a;
    layer0_outputs(410) <= not b or a;
    layer0_outputs(411) <= a;
    layer0_outputs(412) <= a and b;
    layer0_outputs(413) <= a and b;
    layer0_outputs(414) <= 1'b1;
    layer0_outputs(415) <= not (a or b);
    layer0_outputs(416) <= not b or a;
    layer0_outputs(417) <= a or b;
    layer0_outputs(418) <= a and not b;
    layer0_outputs(419) <= a or b;
    layer0_outputs(420) <= b;
    layer0_outputs(421) <= not (a xor b);
    layer0_outputs(422) <= a or b;
    layer0_outputs(423) <= a;
    layer0_outputs(424) <= a xor b;
    layer0_outputs(425) <= a and b;
    layer0_outputs(426) <= not b;
    layer0_outputs(427) <= not a;
    layer0_outputs(428) <= a or b;
    layer0_outputs(429) <= not (a or b);
    layer0_outputs(430) <= not a or b;
    layer0_outputs(431) <= a and not b;
    layer0_outputs(432) <= not (a and b);
    layer0_outputs(433) <= not (a or b);
    layer0_outputs(434) <= not b;
    layer0_outputs(435) <= not b;
    layer0_outputs(436) <= b;
    layer0_outputs(437) <= not (a or b);
    layer0_outputs(438) <= b and not a;
    layer0_outputs(439) <= b;
    layer0_outputs(440) <= b;
    layer0_outputs(441) <= b and not a;
    layer0_outputs(442) <= a;
    layer0_outputs(443) <= b and not a;
    layer0_outputs(444) <= a;
    layer0_outputs(445) <= a xor b;
    layer0_outputs(446) <= a xor b;
    layer0_outputs(447) <= not (a or b);
    layer0_outputs(448) <= not (a xor b);
    layer0_outputs(449) <= b and not a;
    layer0_outputs(450) <= not (a or b);
    layer0_outputs(451) <= not (a or b);
    layer0_outputs(452) <= a or b;
    layer0_outputs(453) <= not (a or b);
    layer0_outputs(454) <= a or b;
    layer0_outputs(455) <= not a;
    layer0_outputs(456) <= b;
    layer0_outputs(457) <= not a or b;
    layer0_outputs(458) <= not a;
    layer0_outputs(459) <= a or b;
    layer0_outputs(460) <= not (a xor b);
    layer0_outputs(461) <= b and not a;
    layer0_outputs(462) <= not a;
    layer0_outputs(463) <= not a;
    layer0_outputs(464) <= a or b;
    layer0_outputs(465) <= a and not b;
    layer0_outputs(466) <= not a or b;
    layer0_outputs(467) <= a and not b;
    layer0_outputs(468) <= not b;
    layer0_outputs(469) <= a;
    layer0_outputs(470) <= not (a and b);
    layer0_outputs(471) <= a and not b;
    layer0_outputs(472) <= a or b;
    layer0_outputs(473) <= a and not b;
    layer0_outputs(474) <= 1'b1;
    layer0_outputs(475) <= not (a and b);
    layer0_outputs(476) <= not (a or b);
    layer0_outputs(477) <= not b;
    layer0_outputs(478) <= not a or b;
    layer0_outputs(479) <= 1'b0;
    layer0_outputs(480) <= 1'b0;
    layer0_outputs(481) <= a;
    layer0_outputs(482) <= not (a xor b);
    layer0_outputs(483) <= not b;
    layer0_outputs(484) <= not a or b;
    layer0_outputs(485) <= not a or b;
    layer0_outputs(486) <= b and not a;
    layer0_outputs(487) <= not b or a;
    layer0_outputs(488) <= not (a or b);
    layer0_outputs(489) <= not a or b;
    layer0_outputs(490) <= a;
    layer0_outputs(491) <= a and not b;
    layer0_outputs(492) <= b and not a;
    layer0_outputs(493) <= not b or a;
    layer0_outputs(494) <= a or b;
    layer0_outputs(495) <= a and not b;
    layer0_outputs(496) <= not (a and b);
    layer0_outputs(497) <= a and not b;
    layer0_outputs(498) <= b and not a;
    layer0_outputs(499) <= not a;
    layer0_outputs(500) <= not (a or b);
    layer0_outputs(501) <= a or b;
    layer0_outputs(502) <= a or b;
    layer0_outputs(503) <= not (a or b);
    layer0_outputs(504) <= not (a or b);
    layer0_outputs(505) <= a and not b;
    layer0_outputs(506) <= a;
    layer0_outputs(507) <= a or b;
    layer0_outputs(508) <= not a or b;
    layer0_outputs(509) <= a xor b;
    layer0_outputs(510) <= a xor b;
    layer0_outputs(511) <= not (a or b);
    layer0_outputs(512) <= not (a or b);
    layer0_outputs(513) <= b and not a;
    layer0_outputs(514) <= not b or a;
    layer0_outputs(515) <= a xor b;
    layer0_outputs(516) <= not b or a;
    layer0_outputs(517) <= a and b;
    layer0_outputs(518) <= a xor b;
    layer0_outputs(519) <= a and not b;
    layer0_outputs(520) <= not a or b;
    layer0_outputs(521) <= not (a or b);
    layer0_outputs(522) <= not (a xor b);
    layer0_outputs(523) <= a xor b;
    layer0_outputs(524) <= not b;
    layer0_outputs(525) <= a or b;
    layer0_outputs(526) <= not a;
    layer0_outputs(527) <= b;
    layer0_outputs(528) <= not b or a;
    layer0_outputs(529) <= a;
    layer0_outputs(530) <= not (a and b);
    layer0_outputs(531) <= not b;
    layer0_outputs(532) <= b;
    layer0_outputs(533) <= a xor b;
    layer0_outputs(534) <= b and not a;
    layer0_outputs(535) <= not a;
    layer0_outputs(536) <= a and not b;
    layer0_outputs(537) <= b;
    layer0_outputs(538) <= not b or a;
    layer0_outputs(539) <= a or b;
    layer0_outputs(540) <= not (a xor b);
    layer0_outputs(541) <= a xor b;
    layer0_outputs(542) <= b;
    layer0_outputs(543) <= not b or a;
    layer0_outputs(544) <= a xor b;
    layer0_outputs(545) <= not a or b;
    layer0_outputs(546) <= b;
    layer0_outputs(547) <= 1'b0;
    layer0_outputs(548) <= a;
    layer0_outputs(549) <= not b or a;
    layer0_outputs(550) <= not (a or b);
    layer0_outputs(551) <= not (a xor b);
    layer0_outputs(552) <= a and not b;
    layer0_outputs(553) <= a or b;
    layer0_outputs(554) <= not (a or b);
    layer0_outputs(555) <= a;
    layer0_outputs(556) <= not (a xor b);
    layer0_outputs(557) <= not a;
    layer0_outputs(558) <= a;
    layer0_outputs(559) <= b;
    layer0_outputs(560) <= b and not a;
    layer0_outputs(561) <= not (a or b);
    layer0_outputs(562) <= a and b;
    layer0_outputs(563) <= 1'b0;
    layer0_outputs(564) <= a and not b;
    layer0_outputs(565) <= not (a or b);
    layer0_outputs(566) <= a and b;
    layer0_outputs(567) <= 1'b0;
    layer0_outputs(568) <= not (a and b);
    layer0_outputs(569) <= not b or a;
    layer0_outputs(570) <= not (a or b);
    layer0_outputs(571) <= a or b;
    layer0_outputs(572) <= a;
    layer0_outputs(573) <= not (a or b);
    layer0_outputs(574) <= not (a or b);
    layer0_outputs(575) <= not (a xor b);
    layer0_outputs(576) <= not b;
    layer0_outputs(577) <= not b;
    layer0_outputs(578) <= b and not a;
    layer0_outputs(579) <= a xor b;
    layer0_outputs(580) <= not a or b;
    layer0_outputs(581) <= not a;
    layer0_outputs(582) <= not (a and b);
    layer0_outputs(583) <= not (a and b);
    layer0_outputs(584) <= not a or b;
    layer0_outputs(585) <= b and not a;
    layer0_outputs(586) <= a or b;
    layer0_outputs(587) <= a xor b;
    layer0_outputs(588) <= a xor b;
    layer0_outputs(589) <= a or b;
    layer0_outputs(590) <= not a or b;
    layer0_outputs(591) <= not (a and b);
    layer0_outputs(592) <= not b;
    layer0_outputs(593) <= b and not a;
    layer0_outputs(594) <= a xor b;
    layer0_outputs(595) <= not (a or b);
    layer0_outputs(596) <= a;
    layer0_outputs(597) <= not b;
    layer0_outputs(598) <= b and not a;
    layer0_outputs(599) <= b;
    layer0_outputs(600) <= not b or a;
    layer0_outputs(601) <= not a or b;
    layer0_outputs(602) <= a and b;
    layer0_outputs(603) <= not (a or b);
    layer0_outputs(604) <= 1'b0;
    layer0_outputs(605) <= not (a and b);
    layer0_outputs(606) <= not a;
    layer0_outputs(607) <= not a or b;
    layer0_outputs(608) <= 1'b1;
    layer0_outputs(609) <= a or b;
    layer0_outputs(610) <= not b;
    layer0_outputs(611) <= not a;
    layer0_outputs(612) <= 1'b1;
    layer0_outputs(613) <= b;
    layer0_outputs(614) <= a and not b;
    layer0_outputs(615) <= not (a and b);
    layer0_outputs(616) <= not (a xor b);
    layer0_outputs(617) <= a and b;
    layer0_outputs(618) <= a or b;
    layer0_outputs(619) <= a and b;
    layer0_outputs(620) <= not (a xor b);
    layer0_outputs(621) <= not b or a;
    layer0_outputs(622) <= not a;
    layer0_outputs(623) <= not b or a;
    layer0_outputs(624) <= not (a or b);
    layer0_outputs(625) <= not b;
    layer0_outputs(626) <= not (a or b);
    layer0_outputs(627) <= b;
    layer0_outputs(628) <= a xor b;
    layer0_outputs(629) <= not (a or b);
    layer0_outputs(630) <= not a;
    layer0_outputs(631) <= not (a or b);
    layer0_outputs(632) <= not (a or b);
    layer0_outputs(633) <= a or b;
    layer0_outputs(634) <= not a;
    layer0_outputs(635) <= not b;
    layer0_outputs(636) <= not (a or b);
    layer0_outputs(637) <= not a;
    layer0_outputs(638) <= not b;
    layer0_outputs(639) <= b;
    layer0_outputs(640) <= 1'b0;
    layer0_outputs(641) <= b;
    layer0_outputs(642) <= a and b;
    layer0_outputs(643) <= not (a xor b);
    layer0_outputs(644) <= a xor b;
    layer0_outputs(645) <= not a or b;
    layer0_outputs(646) <= not a;
    layer0_outputs(647) <= not b;
    layer0_outputs(648) <= not b or a;
    layer0_outputs(649) <= not b;
    layer0_outputs(650) <= a or b;
    layer0_outputs(651) <= a and not b;
    layer0_outputs(652) <= a or b;
    layer0_outputs(653) <= not a or b;
    layer0_outputs(654) <= not b;
    layer0_outputs(655) <= not b or a;
    layer0_outputs(656) <= a or b;
    layer0_outputs(657) <= a or b;
    layer0_outputs(658) <= b and not a;
    layer0_outputs(659) <= a;
    layer0_outputs(660) <= b and not a;
    layer0_outputs(661) <= b and not a;
    layer0_outputs(662) <= a;
    layer0_outputs(663) <= a or b;
    layer0_outputs(664) <= not a or b;
    layer0_outputs(665) <= not (a and b);
    layer0_outputs(666) <= not b;
    layer0_outputs(667) <= not (a xor b);
    layer0_outputs(668) <= not b or a;
    layer0_outputs(669) <= not (a xor b);
    layer0_outputs(670) <= a or b;
    layer0_outputs(671) <= not (a or b);
    layer0_outputs(672) <= a;
    layer0_outputs(673) <= a;
    layer0_outputs(674) <= a or b;
    layer0_outputs(675) <= not b or a;
    layer0_outputs(676) <= a and not b;
    layer0_outputs(677) <= not (a or b);
    layer0_outputs(678) <= not b;
    layer0_outputs(679) <= not (a and b);
    layer0_outputs(680) <= not a or b;
    layer0_outputs(681) <= a and not b;
    layer0_outputs(682) <= not (a or b);
    layer0_outputs(683) <= b and not a;
    layer0_outputs(684) <= a and b;
    layer0_outputs(685) <= not b;
    layer0_outputs(686) <= a xor b;
    layer0_outputs(687) <= not a or b;
    layer0_outputs(688) <= not b or a;
    layer0_outputs(689) <= b;
    layer0_outputs(690) <= not (a or b);
    layer0_outputs(691) <= a or b;
    layer0_outputs(692) <= a;
    layer0_outputs(693) <= 1'b0;
    layer0_outputs(694) <= a or b;
    layer0_outputs(695) <= not b;
    layer0_outputs(696) <= b and not a;
    layer0_outputs(697) <= not b or a;
    layer0_outputs(698) <= a xor b;
    layer0_outputs(699) <= not (a xor b);
    layer0_outputs(700) <= not b or a;
    layer0_outputs(701) <= not (a or b);
    layer0_outputs(702) <= b and not a;
    layer0_outputs(703) <= 1'b0;
    layer0_outputs(704) <= not (a or b);
    layer0_outputs(705) <= a or b;
    layer0_outputs(706) <= not a;
    layer0_outputs(707) <= not (a or b);
    layer0_outputs(708) <= not (a xor b);
    layer0_outputs(709) <= not b;
    layer0_outputs(710) <= a and not b;
    layer0_outputs(711) <= a or b;
    layer0_outputs(712) <= not a;
    layer0_outputs(713) <= a xor b;
    layer0_outputs(714) <= not (a xor b);
    layer0_outputs(715) <= a and not b;
    layer0_outputs(716) <= not (a or b);
    layer0_outputs(717) <= 1'b0;
    layer0_outputs(718) <= not a;
    layer0_outputs(719) <= not (a xor b);
    layer0_outputs(720) <= b and not a;
    layer0_outputs(721) <= a xor b;
    layer0_outputs(722) <= not (a or b);
    layer0_outputs(723) <= a;
    layer0_outputs(724) <= not b;
    layer0_outputs(725) <= b and not a;
    layer0_outputs(726) <= not (a or b);
    layer0_outputs(727) <= a xor b;
    layer0_outputs(728) <= a or b;
    layer0_outputs(729) <= not a;
    layer0_outputs(730) <= not (a or b);
    layer0_outputs(731) <= not (a or b);
    layer0_outputs(732) <= not b or a;
    layer0_outputs(733) <= a xor b;
    layer0_outputs(734) <= a xor b;
    layer0_outputs(735) <= a or b;
    layer0_outputs(736) <= not (a or b);
    layer0_outputs(737) <= b;
    layer0_outputs(738) <= not a;
    layer0_outputs(739) <= not a or b;
    layer0_outputs(740) <= a or b;
    layer0_outputs(741) <= a;
    layer0_outputs(742) <= not a;
    layer0_outputs(743) <= a;
    layer0_outputs(744) <= not (a or b);
    layer0_outputs(745) <= a or b;
    layer0_outputs(746) <= not (a xor b);
    layer0_outputs(747) <= a or b;
    layer0_outputs(748) <= a and not b;
    layer0_outputs(749) <= b and not a;
    layer0_outputs(750) <= a;
    layer0_outputs(751) <= not b or a;
    layer0_outputs(752) <= not a;
    layer0_outputs(753) <= b and not a;
    layer0_outputs(754) <= not a or b;
    layer0_outputs(755) <= not (a or b);
    layer0_outputs(756) <= not a;
    layer0_outputs(757) <= not (a xor b);
    layer0_outputs(758) <= 1'b0;
    layer0_outputs(759) <= not a;
    layer0_outputs(760) <= a or b;
    layer0_outputs(761) <= a xor b;
    layer0_outputs(762) <= b;
    layer0_outputs(763) <= not (a xor b);
    layer0_outputs(764) <= not b;
    layer0_outputs(765) <= not (a xor b);
    layer0_outputs(766) <= a xor b;
    layer0_outputs(767) <= not (a or b);
    layer0_outputs(768) <= not b;
    layer0_outputs(769) <= not (a or b);
    layer0_outputs(770) <= b and not a;
    layer0_outputs(771) <= not a;
    layer0_outputs(772) <= not b or a;
    layer0_outputs(773) <= not b;
    layer0_outputs(774) <= 1'b0;
    layer0_outputs(775) <= a and not b;
    layer0_outputs(776) <= 1'b0;
    layer0_outputs(777) <= not b or a;
    layer0_outputs(778) <= b;
    layer0_outputs(779) <= not (a or b);
    layer0_outputs(780) <= a xor b;
    layer0_outputs(781) <= a;
    layer0_outputs(782) <= b and not a;
    layer0_outputs(783) <= a or b;
    layer0_outputs(784) <= not (a xor b);
    layer0_outputs(785) <= not b;
    layer0_outputs(786) <= a;
    layer0_outputs(787) <= a or b;
    layer0_outputs(788) <= not (a or b);
    layer0_outputs(789) <= a and not b;
    layer0_outputs(790) <= a;
    layer0_outputs(791) <= 1'b0;
    layer0_outputs(792) <= a and not b;
    layer0_outputs(793) <= not b;
    layer0_outputs(794) <= b;
    layer0_outputs(795) <= not b or a;
    layer0_outputs(796) <= b and not a;
    layer0_outputs(797) <= not (a or b);
    layer0_outputs(798) <= b;
    layer0_outputs(799) <= not a or b;
    layer0_outputs(800) <= 1'b1;
    layer0_outputs(801) <= a and not b;
    layer0_outputs(802) <= not (a or b);
    layer0_outputs(803) <= not a;
    layer0_outputs(804) <= a and not b;
    layer0_outputs(805) <= b;
    layer0_outputs(806) <= a;
    layer0_outputs(807) <= a xor b;
    layer0_outputs(808) <= not (a xor b);
    layer0_outputs(809) <= not a;
    layer0_outputs(810) <= a xor b;
    layer0_outputs(811) <= not (a and b);
    layer0_outputs(812) <= not (a xor b);
    layer0_outputs(813) <= a and b;
    layer0_outputs(814) <= b;
    layer0_outputs(815) <= not a;
    layer0_outputs(816) <= not a;
    layer0_outputs(817) <= not (a or b);
    layer0_outputs(818) <= not b;
    layer0_outputs(819) <= a;
    layer0_outputs(820) <= not (a or b);
    layer0_outputs(821) <= not (a or b);
    layer0_outputs(822) <= a xor b;
    layer0_outputs(823) <= a or b;
    layer0_outputs(824) <= not b;
    layer0_outputs(825) <= b;
    layer0_outputs(826) <= a and not b;
    layer0_outputs(827) <= b and not a;
    layer0_outputs(828) <= b and not a;
    layer0_outputs(829) <= not (a or b);
    layer0_outputs(830) <= a and not b;
    layer0_outputs(831) <= not (a xor b);
    layer0_outputs(832) <= not (a or b);
    layer0_outputs(833) <= a or b;
    layer0_outputs(834) <= a or b;
    layer0_outputs(835) <= not (a or b);
    layer0_outputs(836) <= b;
    layer0_outputs(837) <= a xor b;
    layer0_outputs(838) <= a and not b;
    layer0_outputs(839) <= a;
    layer0_outputs(840) <= not b;
    layer0_outputs(841) <= not b;
    layer0_outputs(842) <= not b;
    layer0_outputs(843) <= not a;
    layer0_outputs(844) <= not a or b;
    layer0_outputs(845) <= not (a or b);
    layer0_outputs(846) <= not (a or b);
    layer0_outputs(847) <= not (a or b);
    layer0_outputs(848) <= 1'b0;
    layer0_outputs(849) <= a or b;
    layer0_outputs(850) <= not b;
    layer0_outputs(851) <= a and b;
    layer0_outputs(852) <= a xor b;
    layer0_outputs(853) <= 1'b1;
    layer0_outputs(854) <= not a or b;
    layer0_outputs(855) <= not b;
    layer0_outputs(856) <= not b or a;
    layer0_outputs(857) <= not b;
    layer0_outputs(858) <= not (a or b);
    layer0_outputs(859) <= b and not a;
    layer0_outputs(860) <= not (a or b);
    layer0_outputs(861) <= not (a or b);
    layer0_outputs(862) <= not (a and b);
    layer0_outputs(863) <= a;
    layer0_outputs(864) <= not a or b;
    layer0_outputs(865) <= not (a xor b);
    layer0_outputs(866) <= not (a or b);
    layer0_outputs(867) <= not (a xor b);
    layer0_outputs(868) <= not b or a;
    layer0_outputs(869) <= a;
    layer0_outputs(870) <= a or b;
    layer0_outputs(871) <= not (a xor b);
    layer0_outputs(872) <= a and not b;
    layer0_outputs(873) <= not (a or b);
    layer0_outputs(874) <= a xor b;
    layer0_outputs(875) <= not (a xor b);
    layer0_outputs(876) <= b;
    layer0_outputs(877) <= a or b;
    layer0_outputs(878) <= a or b;
    layer0_outputs(879) <= not (a or b);
    layer0_outputs(880) <= not (a or b);
    layer0_outputs(881) <= a;
    layer0_outputs(882) <= a or b;
    layer0_outputs(883) <= b and not a;
    layer0_outputs(884) <= a xor b;
    layer0_outputs(885) <= b and not a;
    layer0_outputs(886) <= not (a xor b);
    layer0_outputs(887) <= a;
    layer0_outputs(888) <= a or b;
    layer0_outputs(889) <= not (a xor b);
    layer0_outputs(890) <= not a or b;
    layer0_outputs(891) <= a xor b;
    layer0_outputs(892) <= a xor b;
    layer0_outputs(893) <= a and not b;
    layer0_outputs(894) <= b;
    layer0_outputs(895) <= a and b;
    layer0_outputs(896) <= not b;
    layer0_outputs(897) <= not (a or b);
    layer0_outputs(898) <= b and not a;
    layer0_outputs(899) <= not a or b;
    layer0_outputs(900) <= 1'b1;
    layer0_outputs(901) <= not (a or b);
    layer0_outputs(902) <= not (a xor b);
    layer0_outputs(903) <= not a or b;
    layer0_outputs(904) <= not a or b;
    layer0_outputs(905) <= b;
    layer0_outputs(906) <= not b or a;
    layer0_outputs(907) <= not a;
    layer0_outputs(908) <= not b or a;
    layer0_outputs(909) <= 1'b0;
    layer0_outputs(910) <= b and not a;
    layer0_outputs(911) <= not a or b;
    layer0_outputs(912) <= a or b;
    layer0_outputs(913) <= a;
    layer0_outputs(914) <= a xor b;
    layer0_outputs(915) <= 1'b0;
    layer0_outputs(916) <= a xor b;
    layer0_outputs(917) <= a or b;
    layer0_outputs(918) <= b and not a;
    layer0_outputs(919) <= a;
    layer0_outputs(920) <= b and not a;
    layer0_outputs(921) <= not a or b;
    layer0_outputs(922) <= b and not a;
    layer0_outputs(923) <= not (a xor b);
    layer0_outputs(924) <= not b or a;
    layer0_outputs(925) <= b;
    layer0_outputs(926) <= not a or b;
    layer0_outputs(927) <= not a;
    layer0_outputs(928) <= a or b;
    layer0_outputs(929) <= a;
    layer0_outputs(930) <= not (a or b);
    layer0_outputs(931) <= a and not b;
    layer0_outputs(932) <= not a;
    layer0_outputs(933) <= not (a or b);
    layer0_outputs(934) <= not a;
    layer0_outputs(935) <= not b or a;
    layer0_outputs(936) <= 1'b0;
    layer0_outputs(937) <= not a or b;
    layer0_outputs(938) <= not a;
    layer0_outputs(939) <= a xor b;
    layer0_outputs(940) <= a xor b;
    layer0_outputs(941) <= not a;
    layer0_outputs(942) <= not (a xor b);
    layer0_outputs(943) <= b and not a;
    layer0_outputs(944) <= a xor b;
    layer0_outputs(945) <= a or b;
    layer0_outputs(946) <= b and not a;
    layer0_outputs(947) <= a xor b;
    layer0_outputs(948) <= a xor b;
    layer0_outputs(949) <= a;
    layer0_outputs(950) <= b and not a;
    layer0_outputs(951) <= not (a or b);
    layer0_outputs(952) <= b;
    layer0_outputs(953) <= a or b;
    layer0_outputs(954) <= not (a or b);
    layer0_outputs(955) <= a;
    layer0_outputs(956) <= not a;
    layer0_outputs(957) <= a or b;
    layer0_outputs(958) <= not b or a;
    layer0_outputs(959) <= a or b;
    layer0_outputs(960) <= not a or b;
    layer0_outputs(961) <= a or b;
    layer0_outputs(962) <= b;
    layer0_outputs(963) <= not (a xor b);
    layer0_outputs(964) <= not (a xor b);
    layer0_outputs(965) <= a xor b;
    layer0_outputs(966) <= a or b;
    layer0_outputs(967) <= a and not b;
    layer0_outputs(968) <= a or b;
    layer0_outputs(969) <= not b;
    layer0_outputs(970) <= not b;
    layer0_outputs(971) <= a or b;
    layer0_outputs(972) <= not (a xor b);
    layer0_outputs(973) <= a and not b;
    layer0_outputs(974) <= not b;
    layer0_outputs(975) <= not (a xor b);
    layer0_outputs(976) <= a and not b;
    layer0_outputs(977) <= not a or b;
    layer0_outputs(978) <= not (a or b);
    layer0_outputs(979) <= not b or a;
    layer0_outputs(980) <= not a;
    layer0_outputs(981) <= not a;
    layer0_outputs(982) <= b and not a;
    layer0_outputs(983) <= not a;
    layer0_outputs(984) <= 1'b0;
    layer0_outputs(985) <= not a or b;
    layer0_outputs(986) <= not b or a;
    layer0_outputs(987) <= not (a xor b);
    layer0_outputs(988) <= not a or b;
    layer0_outputs(989) <= a or b;
    layer0_outputs(990) <= a xor b;
    layer0_outputs(991) <= b;
    layer0_outputs(992) <= not (a or b);
    layer0_outputs(993) <= a and b;
    layer0_outputs(994) <= a and not b;
    layer0_outputs(995) <= not a or b;
    layer0_outputs(996) <= a and not b;
    layer0_outputs(997) <= not b or a;
    layer0_outputs(998) <= a and b;
    layer0_outputs(999) <= not b;
    layer0_outputs(1000) <= a;
    layer0_outputs(1001) <= not b;
    layer0_outputs(1002) <= a or b;
    layer0_outputs(1003) <= not (a xor b);
    layer0_outputs(1004) <= not b or a;
    layer0_outputs(1005) <= not a;
    layer0_outputs(1006) <= not b;
    layer0_outputs(1007) <= b and not a;
    layer0_outputs(1008) <= not (a or b);
    layer0_outputs(1009) <= not b or a;
    layer0_outputs(1010) <= not b;
    layer0_outputs(1011) <= not (a and b);
    layer0_outputs(1012) <= b and not a;
    layer0_outputs(1013) <= not a or b;
    layer0_outputs(1014) <= a or b;
    layer0_outputs(1015) <= a or b;
    layer0_outputs(1016) <= b;
    layer0_outputs(1017) <= a or b;
    layer0_outputs(1018) <= a;
    layer0_outputs(1019) <= not (a or b);
    layer0_outputs(1020) <= a and not b;
    layer0_outputs(1021) <= b;
    layer0_outputs(1022) <= not (a or b);
    layer0_outputs(1023) <= not (a xor b);
    layer0_outputs(1024) <= not b;
    layer0_outputs(1025) <= not (a or b);
    layer0_outputs(1026) <= a;
    layer0_outputs(1027) <= 1'b1;
    layer0_outputs(1028) <= not (a or b);
    layer0_outputs(1029) <= a or b;
    layer0_outputs(1030) <= not (a xor b);
    layer0_outputs(1031) <= a xor b;
    layer0_outputs(1032) <= a or b;
    layer0_outputs(1033) <= not (a or b);
    layer0_outputs(1034) <= not (a or b);
    layer0_outputs(1035) <= not a or b;
    layer0_outputs(1036) <= not a;
    layer0_outputs(1037) <= a or b;
    layer0_outputs(1038) <= not (a xor b);
    layer0_outputs(1039) <= not a;
    layer0_outputs(1040) <= a or b;
    layer0_outputs(1041) <= not b;
    layer0_outputs(1042) <= a and b;
    layer0_outputs(1043) <= not (a or b);
    layer0_outputs(1044) <= a and b;
    layer0_outputs(1045) <= 1'b0;
    layer0_outputs(1046) <= a or b;
    layer0_outputs(1047) <= not (a or b);
    layer0_outputs(1048) <= a or b;
    layer0_outputs(1049) <= not (a or b);
    layer0_outputs(1050) <= not b or a;
    layer0_outputs(1051) <= not a;
    layer0_outputs(1052) <= a;
    layer0_outputs(1053) <= not (a or b);
    layer0_outputs(1054) <= b;
    layer0_outputs(1055) <= not (a xor b);
    layer0_outputs(1056) <= not b or a;
    layer0_outputs(1057) <= not (a or b);
    layer0_outputs(1058) <= a xor b;
    layer0_outputs(1059) <= not b;
    layer0_outputs(1060) <= not a or b;
    layer0_outputs(1061) <= a or b;
    layer0_outputs(1062) <= not b;
    layer0_outputs(1063) <= not a or b;
    layer0_outputs(1064) <= not (a xor b);
    layer0_outputs(1065) <= a and not b;
    layer0_outputs(1066) <= b;
    layer0_outputs(1067) <= a xor b;
    layer0_outputs(1068) <= not (a or b);
    layer0_outputs(1069) <= not (a xor b);
    layer0_outputs(1070) <= a and not b;
    layer0_outputs(1071) <= 1'b1;
    layer0_outputs(1072) <= a and not b;
    layer0_outputs(1073) <= a xor b;
    layer0_outputs(1074) <= not a;
    layer0_outputs(1075) <= 1'b1;
    layer0_outputs(1076) <= b;
    layer0_outputs(1077) <= not (a xor b);
    layer0_outputs(1078) <= b;
    layer0_outputs(1079) <= a;
    layer0_outputs(1080) <= not (a or b);
    layer0_outputs(1081) <= not (a and b);
    layer0_outputs(1082) <= not a or b;
    layer0_outputs(1083) <= b;
    layer0_outputs(1084) <= a and not b;
    layer0_outputs(1085) <= not (a or b);
    layer0_outputs(1086) <= a xor b;
    layer0_outputs(1087) <= not b;
    layer0_outputs(1088) <= not b or a;
    layer0_outputs(1089) <= not a or b;
    layer0_outputs(1090) <= not a;
    layer0_outputs(1091) <= a and b;
    layer0_outputs(1092) <= b and not a;
    layer0_outputs(1093) <= not a;
    layer0_outputs(1094) <= not a or b;
    layer0_outputs(1095) <= b;
    layer0_outputs(1096) <= not a;
    layer0_outputs(1097) <= a xor b;
    layer0_outputs(1098) <= a;
    layer0_outputs(1099) <= not (a xor b);
    layer0_outputs(1100) <= not b;
    layer0_outputs(1101) <= a;
    layer0_outputs(1102) <= a or b;
    layer0_outputs(1103) <= b;
    layer0_outputs(1104) <= b;
    layer0_outputs(1105) <= a xor b;
    layer0_outputs(1106) <= a;
    layer0_outputs(1107) <= a xor b;
    layer0_outputs(1108) <= not (a and b);
    layer0_outputs(1109) <= b and not a;
    layer0_outputs(1110) <= not a;
    layer0_outputs(1111) <= not a or b;
    layer0_outputs(1112) <= a xor b;
    layer0_outputs(1113) <= a xor b;
    layer0_outputs(1114) <= a or b;
    layer0_outputs(1115) <= not (a xor b);
    layer0_outputs(1116) <= not (a xor b);
    layer0_outputs(1117) <= a or b;
    layer0_outputs(1118) <= a and not b;
    layer0_outputs(1119) <= not (a or b);
    layer0_outputs(1120) <= b;
    layer0_outputs(1121) <= not (a or b);
    layer0_outputs(1122) <= a or b;
    layer0_outputs(1123) <= a xor b;
    layer0_outputs(1124) <= not (a or b);
    layer0_outputs(1125) <= not b or a;
    layer0_outputs(1126) <= a and b;
    layer0_outputs(1127) <= not b or a;
    layer0_outputs(1128) <= not b;
    layer0_outputs(1129) <= not (a xor b);
    layer0_outputs(1130) <= not a or b;
    layer0_outputs(1131) <= a or b;
    layer0_outputs(1132) <= a or b;
    layer0_outputs(1133) <= a or b;
    layer0_outputs(1134) <= not (a or b);
    layer0_outputs(1135) <= a or b;
    layer0_outputs(1136) <= not (a xor b);
    layer0_outputs(1137) <= a xor b;
    layer0_outputs(1138) <= not (a and b);
    layer0_outputs(1139) <= b;
    layer0_outputs(1140) <= not a or b;
    layer0_outputs(1141) <= a or b;
    layer0_outputs(1142) <= 1'b0;
    layer0_outputs(1143) <= a;
    layer0_outputs(1144) <= not b;
    layer0_outputs(1145) <= 1'b0;
    layer0_outputs(1146) <= not (a or b);
    layer0_outputs(1147) <= not (a xor b);
    layer0_outputs(1148) <= not (a xor b);
    layer0_outputs(1149) <= not b;
    layer0_outputs(1150) <= not b;
    layer0_outputs(1151) <= not (a or b);
    layer0_outputs(1152) <= a;
    layer0_outputs(1153) <= b;
    layer0_outputs(1154) <= not (a and b);
    layer0_outputs(1155) <= not (a or b);
    layer0_outputs(1156) <= not (a xor b);
    layer0_outputs(1157) <= b and not a;
    layer0_outputs(1158) <= a xor b;
    layer0_outputs(1159) <= b;
    layer0_outputs(1160) <= a or b;
    layer0_outputs(1161) <= b and not a;
    layer0_outputs(1162) <= a or b;
    layer0_outputs(1163) <= a;
    layer0_outputs(1164) <= not b or a;
    layer0_outputs(1165) <= not a or b;
    layer0_outputs(1166) <= not (a or b);
    layer0_outputs(1167) <= not b or a;
    layer0_outputs(1168) <= not (a and b);
    layer0_outputs(1169) <= a or b;
    layer0_outputs(1170) <= not b;
    layer0_outputs(1171) <= a xor b;
    layer0_outputs(1172) <= 1'b1;
    layer0_outputs(1173) <= not a or b;
    layer0_outputs(1174) <= b and not a;
    layer0_outputs(1175) <= a;
    layer0_outputs(1176) <= b;
    layer0_outputs(1177) <= a;
    layer0_outputs(1178) <= not (a or b);
    layer0_outputs(1179) <= b;
    layer0_outputs(1180) <= a or b;
    layer0_outputs(1181) <= not a or b;
    layer0_outputs(1182) <= b;
    layer0_outputs(1183) <= not (a xor b);
    layer0_outputs(1184) <= a;
    layer0_outputs(1185) <= not a or b;
    layer0_outputs(1186) <= 1'b1;
    layer0_outputs(1187) <= not (a or b);
    layer0_outputs(1188) <= a and not b;
    layer0_outputs(1189) <= b;
    layer0_outputs(1190) <= not (a and b);
    layer0_outputs(1191) <= not b;
    layer0_outputs(1192) <= not b or a;
    layer0_outputs(1193) <= not b or a;
    layer0_outputs(1194) <= b;
    layer0_outputs(1195) <= not a;
    layer0_outputs(1196) <= a and not b;
    layer0_outputs(1197) <= 1'b0;
    layer0_outputs(1198) <= a or b;
    layer0_outputs(1199) <= a or b;
    layer0_outputs(1200) <= not b;
    layer0_outputs(1201) <= not (a xor b);
    layer0_outputs(1202) <= not (a or b);
    layer0_outputs(1203) <= a or b;
    layer0_outputs(1204) <= not b;
    layer0_outputs(1205) <= not (a or b);
    layer0_outputs(1206) <= not b;
    layer0_outputs(1207) <= not a;
    layer0_outputs(1208) <= a or b;
    layer0_outputs(1209) <= not b;
    layer0_outputs(1210) <= a or b;
    layer0_outputs(1211) <= not a or b;
    layer0_outputs(1212) <= b;
    layer0_outputs(1213) <= b and not a;
    layer0_outputs(1214) <= not a or b;
    layer0_outputs(1215) <= 1'b1;
    layer0_outputs(1216) <= not (a or b);
    layer0_outputs(1217) <= a or b;
    layer0_outputs(1218) <= not b;
    layer0_outputs(1219) <= a;
    layer0_outputs(1220) <= not (a and b);
    layer0_outputs(1221) <= not (a and b);
    layer0_outputs(1222) <= not (a and b);
    layer0_outputs(1223) <= not a;
    layer0_outputs(1224) <= not (a xor b);
    layer0_outputs(1225) <= not b;
    layer0_outputs(1226) <= b;
    layer0_outputs(1227) <= not b;
    layer0_outputs(1228) <= a;
    layer0_outputs(1229) <= not (a and b);
    layer0_outputs(1230) <= b;
    layer0_outputs(1231) <= not b;
    layer0_outputs(1232) <= not a;
    layer0_outputs(1233) <= a or b;
    layer0_outputs(1234) <= b;
    layer0_outputs(1235) <= not (a or b);
    layer0_outputs(1236) <= b;
    layer0_outputs(1237) <= not a;
    layer0_outputs(1238) <= not b or a;
    layer0_outputs(1239) <= not a;
    layer0_outputs(1240) <= not b;
    layer0_outputs(1241) <= not b;
    layer0_outputs(1242) <= not (a or b);
    layer0_outputs(1243) <= not (a or b);
    layer0_outputs(1244) <= not b;
    layer0_outputs(1245) <= not (a xor b);
    layer0_outputs(1246) <= not a or b;
    layer0_outputs(1247) <= not (a or b);
    layer0_outputs(1248) <= not a;
    layer0_outputs(1249) <= not a or b;
    layer0_outputs(1250) <= not b;
    layer0_outputs(1251) <= not (a xor b);
    layer0_outputs(1252) <= not b or a;
    layer0_outputs(1253) <= b;
    layer0_outputs(1254) <= not b;
    layer0_outputs(1255) <= not a;
    layer0_outputs(1256) <= not b;
    layer0_outputs(1257) <= a;
    layer0_outputs(1258) <= not b;
    layer0_outputs(1259) <= a or b;
    layer0_outputs(1260) <= not (a xor b);
    layer0_outputs(1261) <= a and not b;
    layer0_outputs(1262) <= a or b;
    layer0_outputs(1263) <= not b;
    layer0_outputs(1264) <= not b;
    layer0_outputs(1265) <= not b;
    layer0_outputs(1266) <= a and b;
    layer0_outputs(1267) <= not (a xor b);
    layer0_outputs(1268) <= a xor b;
    layer0_outputs(1269) <= a or b;
    layer0_outputs(1270) <= a;
    layer0_outputs(1271) <= b and not a;
    layer0_outputs(1272) <= not a;
    layer0_outputs(1273) <= b and not a;
    layer0_outputs(1274) <= not (a or b);
    layer0_outputs(1275) <= b and not a;
    layer0_outputs(1276) <= a;
    layer0_outputs(1277) <= not (a xor b);
    layer0_outputs(1278) <= not b or a;
    layer0_outputs(1279) <= not a;
    layer0_outputs(1280) <= not a;
    layer0_outputs(1281) <= a;
    layer0_outputs(1282) <= a or b;
    layer0_outputs(1283) <= not (a or b);
    layer0_outputs(1284) <= not b;
    layer0_outputs(1285) <= not b or a;
    layer0_outputs(1286) <= a xor b;
    layer0_outputs(1287) <= not (a or b);
    layer0_outputs(1288) <= a and not b;
    layer0_outputs(1289) <= b;
    layer0_outputs(1290) <= not (a xor b);
    layer0_outputs(1291) <= 1'b1;
    layer0_outputs(1292) <= not (a xor b);
    layer0_outputs(1293) <= not a or b;
    layer0_outputs(1294) <= a or b;
    layer0_outputs(1295) <= not (a xor b);
    layer0_outputs(1296) <= a xor b;
    layer0_outputs(1297) <= not a or b;
    layer0_outputs(1298) <= not (a or b);
    layer0_outputs(1299) <= a and not b;
    layer0_outputs(1300) <= not a;
    layer0_outputs(1301) <= not a;
    layer0_outputs(1302) <= a xor b;
    layer0_outputs(1303) <= a or b;
    layer0_outputs(1304) <= a or b;
    layer0_outputs(1305) <= not a;
    layer0_outputs(1306) <= a or b;
    layer0_outputs(1307) <= not b;
    layer0_outputs(1308) <= a xor b;
    layer0_outputs(1309) <= not a or b;
    layer0_outputs(1310) <= b and not a;
    layer0_outputs(1311) <= a and b;
    layer0_outputs(1312) <= b and not a;
    layer0_outputs(1313) <= not b;
    layer0_outputs(1314) <= not (a or b);
    layer0_outputs(1315) <= not a;
    layer0_outputs(1316) <= not a or b;
    layer0_outputs(1317) <= b;
    layer0_outputs(1318) <= 1'b1;
    layer0_outputs(1319) <= b;
    layer0_outputs(1320) <= not b or a;
    layer0_outputs(1321) <= a xor b;
    layer0_outputs(1322) <= not (a and b);
    layer0_outputs(1323) <= not a or b;
    layer0_outputs(1324) <= not (a or b);
    layer0_outputs(1325) <= a;
    layer0_outputs(1326) <= b and not a;
    layer0_outputs(1327) <= not b or a;
    layer0_outputs(1328) <= b and not a;
    layer0_outputs(1329) <= not a or b;
    layer0_outputs(1330) <= b and not a;
    layer0_outputs(1331) <= a or b;
    layer0_outputs(1332) <= a xor b;
    layer0_outputs(1333) <= not a;
    layer0_outputs(1334) <= a xor b;
    layer0_outputs(1335) <= a and not b;
    layer0_outputs(1336) <= b and not a;
    layer0_outputs(1337) <= a;
    layer0_outputs(1338) <= a xor b;
    layer0_outputs(1339) <= not (a and b);
    layer0_outputs(1340) <= a xor b;
    layer0_outputs(1341) <= not (a xor b);
    layer0_outputs(1342) <= a;
    layer0_outputs(1343) <= not (a xor b);
    layer0_outputs(1344) <= not b;
    layer0_outputs(1345) <= not a or b;
    layer0_outputs(1346) <= not (a xor b);
    layer0_outputs(1347) <= 1'b0;
    layer0_outputs(1348) <= not b;
    layer0_outputs(1349) <= not a;
    layer0_outputs(1350) <= a xor b;
    layer0_outputs(1351) <= a;
    layer0_outputs(1352) <= b;
    layer0_outputs(1353) <= a and not b;
    layer0_outputs(1354) <= b and not a;
    layer0_outputs(1355) <= not a;
    layer0_outputs(1356) <= a and not b;
    layer0_outputs(1357) <= b and not a;
    layer0_outputs(1358) <= a or b;
    layer0_outputs(1359) <= not a or b;
    layer0_outputs(1360) <= b and not a;
    layer0_outputs(1361) <= not b;
    layer0_outputs(1362) <= a xor b;
    layer0_outputs(1363) <= a and not b;
    layer0_outputs(1364) <= not a or b;
    layer0_outputs(1365) <= a;
    layer0_outputs(1366) <= not (a or b);
    layer0_outputs(1367) <= a or b;
    layer0_outputs(1368) <= a;
    layer0_outputs(1369) <= not a;
    layer0_outputs(1370) <= a or b;
    layer0_outputs(1371) <= not (a xor b);
    layer0_outputs(1372) <= a;
    layer0_outputs(1373) <= not a;
    layer0_outputs(1374) <= not (a or b);
    layer0_outputs(1375) <= not b;
    layer0_outputs(1376) <= b;
    layer0_outputs(1377) <= a and not b;
    layer0_outputs(1378) <= 1'b1;
    layer0_outputs(1379) <= 1'b1;
    layer0_outputs(1380) <= not (a or b);
    layer0_outputs(1381) <= not (a or b);
    layer0_outputs(1382) <= a and b;
    layer0_outputs(1383) <= a;
    layer0_outputs(1384) <= a and not b;
    layer0_outputs(1385) <= a and not b;
    layer0_outputs(1386) <= a or b;
    layer0_outputs(1387) <= b and not a;
    layer0_outputs(1388) <= not b;
    layer0_outputs(1389) <= 1'b0;
    layer0_outputs(1390) <= 1'b0;
    layer0_outputs(1391) <= a or b;
    layer0_outputs(1392) <= a or b;
    layer0_outputs(1393) <= not (a or b);
    layer0_outputs(1394) <= b and not a;
    layer0_outputs(1395) <= b;
    layer0_outputs(1396) <= a xor b;
    layer0_outputs(1397) <= not (a or b);
    layer0_outputs(1398) <= not b or a;
    layer0_outputs(1399) <= not (a xor b);
    layer0_outputs(1400) <= b;
    layer0_outputs(1401) <= a or b;
    layer0_outputs(1402) <= not b;
    layer0_outputs(1403) <= b and not a;
    layer0_outputs(1404) <= not (a or b);
    layer0_outputs(1405) <= a or b;
    layer0_outputs(1406) <= not b;
    layer0_outputs(1407) <= not (a and b);
    layer0_outputs(1408) <= 1'b0;
    layer0_outputs(1409) <= a or b;
    layer0_outputs(1410) <= b;
    layer0_outputs(1411) <= b and not a;
    layer0_outputs(1412) <= not (a xor b);
    layer0_outputs(1413) <= not a or b;
    layer0_outputs(1414) <= a;
    layer0_outputs(1415) <= not b or a;
    layer0_outputs(1416) <= not a or b;
    layer0_outputs(1417) <= a;
    layer0_outputs(1418) <= b;
    layer0_outputs(1419) <= 1'b0;
    layer0_outputs(1420) <= not b or a;
    layer0_outputs(1421) <= a;
    layer0_outputs(1422) <= not b or a;
    layer0_outputs(1423) <= a or b;
    layer0_outputs(1424) <= a;
    layer0_outputs(1425) <= 1'b0;
    layer0_outputs(1426) <= not b or a;
    layer0_outputs(1427) <= not (a xor b);
    layer0_outputs(1428) <= a or b;
    layer0_outputs(1429) <= a xor b;
    layer0_outputs(1430) <= not (a xor b);
    layer0_outputs(1431) <= not b;
    layer0_outputs(1432) <= b;
    layer0_outputs(1433) <= not (a or b);
    layer0_outputs(1434) <= not b or a;
    layer0_outputs(1435) <= a;
    layer0_outputs(1436) <= not (a or b);
    layer0_outputs(1437) <= b and not a;
    layer0_outputs(1438) <= 1'b0;
    layer0_outputs(1439) <= b and not a;
    layer0_outputs(1440) <= a or b;
    layer0_outputs(1441) <= not b;
    layer0_outputs(1442) <= not (a or b);
    layer0_outputs(1443) <= a;
    layer0_outputs(1444) <= a or b;
    layer0_outputs(1445) <= not (a or b);
    layer0_outputs(1446) <= not b or a;
    layer0_outputs(1447) <= not b;
    layer0_outputs(1448) <= a or b;
    layer0_outputs(1449) <= a or b;
    layer0_outputs(1450) <= not (a or b);
    layer0_outputs(1451) <= a xor b;
    layer0_outputs(1452) <= not b;
    layer0_outputs(1453) <= not a;
    layer0_outputs(1454) <= not b;
    layer0_outputs(1455) <= a xor b;
    layer0_outputs(1456) <= not a;
    layer0_outputs(1457) <= a;
    layer0_outputs(1458) <= not b or a;
    layer0_outputs(1459) <= a;
    layer0_outputs(1460) <= not (a or b);
    layer0_outputs(1461) <= a or b;
    layer0_outputs(1462) <= b and not a;
    layer0_outputs(1463) <= not (a or b);
    layer0_outputs(1464) <= a;
    layer0_outputs(1465) <= not b;
    layer0_outputs(1466) <= not a;
    layer0_outputs(1467) <= a or b;
    layer0_outputs(1468) <= not (a xor b);
    layer0_outputs(1469) <= not (a or b);
    layer0_outputs(1470) <= not a;
    layer0_outputs(1471) <= a;
    layer0_outputs(1472) <= a xor b;
    layer0_outputs(1473) <= b and not a;
    layer0_outputs(1474) <= not (a or b);
    layer0_outputs(1475) <= not (a or b);
    layer0_outputs(1476) <= not (a xor b);
    layer0_outputs(1477) <= not b;
    layer0_outputs(1478) <= not b or a;
    layer0_outputs(1479) <= a xor b;
    layer0_outputs(1480) <= not b or a;
    layer0_outputs(1481) <= not a;
    layer0_outputs(1482) <= a;
    layer0_outputs(1483) <= not (a and b);
    layer0_outputs(1484) <= not (a xor b);
    layer0_outputs(1485) <= a and not b;
    layer0_outputs(1486) <= not a;
    layer0_outputs(1487) <= not (a xor b);
    layer0_outputs(1488) <= a xor b;
    layer0_outputs(1489) <= not a;
    layer0_outputs(1490) <= a and not b;
    layer0_outputs(1491) <= a;
    layer0_outputs(1492) <= a xor b;
    layer0_outputs(1493) <= not b or a;
    layer0_outputs(1494) <= b;
    layer0_outputs(1495) <= not b;
    layer0_outputs(1496) <= not a;
    layer0_outputs(1497) <= not a or b;
    layer0_outputs(1498) <= not a or b;
    layer0_outputs(1499) <= not b;
    layer0_outputs(1500) <= not a;
    layer0_outputs(1501) <= not a;
    layer0_outputs(1502) <= a or b;
    layer0_outputs(1503) <= not a;
    layer0_outputs(1504) <= a and not b;
    layer0_outputs(1505) <= a or b;
    layer0_outputs(1506) <= not (a and b);
    layer0_outputs(1507) <= not b or a;
    layer0_outputs(1508) <= not b;
    layer0_outputs(1509) <= not (a xor b);
    layer0_outputs(1510) <= not (a or b);
    layer0_outputs(1511) <= not (a xor b);
    layer0_outputs(1512) <= a and not b;
    layer0_outputs(1513) <= a or b;
    layer0_outputs(1514) <= a or b;
    layer0_outputs(1515) <= a xor b;
    layer0_outputs(1516) <= a and b;
    layer0_outputs(1517) <= a and not b;
    layer0_outputs(1518) <= not (a or b);
    layer0_outputs(1519) <= not a;
    layer0_outputs(1520) <= a;
    layer0_outputs(1521) <= not (a or b);
    layer0_outputs(1522) <= not (a or b);
    layer0_outputs(1523) <= not (a xor b);
    layer0_outputs(1524) <= a xor b;
    layer0_outputs(1525) <= a;
    layer0_outputs(1526) <= not a or b;
    layer0_outputs(1527) <= not b or a;
    layer0_outputs(1528) <= not (a xor b);
    layer0_outputs(1529) <= not a or b;
    layer0_outputs(1530) <= a or b;
    layer0_outputs(1531) <= not (a and b);
    layer0_outputs(1532) <= a or b;
    layer0_outputs(1533) <= a xor b;
    layer0_outputs(1534) <= not a;
    layer0_outputs(1535) <= b and not a;
    layer0_outputs(1536) <= not a or b;
    layer0_outputs(1537) <= a xor b;
    layer0_outputs(1538) <= b and not a;
    layer0_outputs(1539) <= a and not b;
    layer0_outputs(1540) <= not b;
    layer0_outputs(1541) <= not b;
    layer0_outputs(1542) <= not a;
    layer0_outputs(1543) <= 1'b0;
    layer0_outputs(1544) <= b and not a;
    layer0_outputs(1545) <= not (a or b);
    layer0_outputs(1546) <= not (a or b);
    layer0_outputs(1547) <= not (a and b);
    layer0_outputs(1548) <= not (a xor b);
    layer0_outputs(1549) <= a xor b;
    layer0_outputs(1550) <= not b or a;
    layer0_outputs(1551) <= a and not b;
    layer0_outputs(1552) <= a or b;
    layer0_outputs(1553) <= a and not b;
    layer0_outputs(1554) <= 1'b0;
    layer0_outputs(1555) <= b;
    layer0_outputs(1556) <= not a or b;
    layer0_outputs(1557) <= not b;
    layer0_outputs(1558) <= not a or b;
    layer0_outputs(1559) <= a or b;
    layer0_outputs(1560) <= not (a and b);
    layer0_outputs(1561) <= a xor b;
    layer0_outputs(1562) <= not b;
    layer0_outputs(1563) <= not b;
    layer0_outputs(1564) <= b;
    layer0_outputs(1565) <= a xor b;
    layer0_outputs(1566) <= b and not a;
    layer0_outputs(1567) <= not a or b;
    layer0_outputs(1568) <= a or b;
    layer0_outputs(1569) <= not (a or b);
    layer0_outputs(1570) <= a or b;
    layer0_outputs(1571) <= not (a xor b);
    layer0_outputs(1572) <= a or b;
    layer0_outputs(1573) <= not (a xor b);
    layer0_outputs(1574) <= a;
    layer0_outputs(1575) <= not (a or b);
    layer0_outputs(1576) <= a or b;
    layer0_outputs(1577) <= a or b;
    layer0_outputs(1578) <= a and not b;
    layer0_outputs(1579) <= b;
    layer0_outputs(1580) <= b;
    layer0_outputs(1581) <= 1'b0;
    layer0_outputs(1582) <= a;
    layer0_outputs(1583) <= b and not a;
    layer0_outputs(1584) <= not a;
    layer0_outputs(1585) <= 1'b1;
    layer0_outputs(1586) <= a and b;
    layer0_outputs(1587) <= a and b;
    layer0_outputs(1588) <= a and not b;
    layer0_outputs(1589) <= not b or a;
    layer0_outputs(1590) <= a xor b;
    layer0_outputs(1591) <= a or b;
    layer0_outputs(1592) <= not (a or b);
    layer0_outputs(1593) <= 1'b0;
    layer0_outputs(1594) <= b;
    layer0_outputs(1595) <= a or b;
    layer0_outputs(1596) <= a or b;
    layer0_outputs(1597) <= not (a or b);
    layer0_outputs(1598) <= b and not a;
    layer0_outputs(1599) <= 1'b0;
    layer0_outputs(1600) <= a and b;
    layer0_outputs(1601) <= not a or b;
    layer0_outputs(1602) <= not (a or b);
    layer0_outputs(1603) <= a and b;
    layer0_outputs(1604) <= not a;
    layer0_outputs(1605) <= a and b;
    layer0_outputs(1606) <= not (a and b);
    layer0_outputs(1607) <= not b or a;
    layer0_outputs(1608) <= not (a xor b);
    layer0_outputs(1609) <= not a or b;
    layer0_outputs(1610) <= not a;
    layer0_outputs(1611) <= b and not a;
    layer0_outputs(1612) <= not (a xor b);
    layer0_outputs(1613) <= 1'b1;
    layer0_outputs(1614) <= not (a and b);
    layer0_outputs(1615) <= not (a or b);
    layer0_outputs(1616) <= b;
    layer0_outputs(1617) <= not a or b;
    layer0_outputs(1618) <= not b or a;
    layer0_outputs(1619) <= a and not b;
    layer0_outputs(1620) <= not b or a;
    layer0_outputs(1621) <= not (a or b);
    layer0_outputs(1622) <= a xor b;
    layer0_outputs(1623) <= not (a xor b);
    layer0_outputs(1624) <= a xor b;
    layer0_outputs(1625) <= a and b;
    layer0_outputs(1626) <= not a;
    layer0_outputs(1627) <= not a or b;
    layer0_outputs(1628) <= b and not a;
    layer0_outputs(1629) <= a xor b;
    layer0_outputs(1630) <= not a;
    layer0_outputs(1631) <= not (a xor b);
    layer0_outputs(1632) <= not b;
    layer0_outputs(1633) <= not (a xor b);
    layer0_outputs(1634) <= b;
    layer0_outputs(1635) <= not (a or b);
    layer0_outputs(1636) <= not a or b;
    layer0_outputs(1637) <= b and not a;
    layer0_outputs(1638) <= not (a xor b);
    layer0_outputs(1639) <= 1'b0;
    layer0_outputs(1640) <= not b;
    layer0_outputs(1641) <= a;
    layer0_outputs(1642) <= not b;
    layer0_outputs(1643) <= not b or a;
    layer0_outputs(1644) <= not (a or b);
    layer0_outputs(1645) <= not b;
    layer0_outputs(1646) <= not (a or b);
    layer0_outputs(1647) <= a or b;
    layer0_outputs(1648) <= not (a or b);
    layer0_outputs(1649) <= not (a or b);
    layer0_outputs(1650) <= not a or b;
    layer0_outputs(1651) <= a xor b;
    layer0_outputs(1652) <= a xor b;
    layer0_outputs(1653) <= a;
    layer0_outputs(1654) <= not b;
    layer0_outputs(1655) <= a or b;
    layer0_outputs(1656) <= not b or a;
    layer0_outputs(1657) <= not (a xor b);
    layer0_outputs(1658) <= not (a or b);
    layer0_outputs(1659) <= not a or b;
    layer0_outputs(1660) <= b and not a;
    layer0_outputs(1661) <= not a;
    layer0_outputs(1662) <= not (a or b);
    layer0_outputs(1663) <= not (a xor b);
    layer0_outputs(1664) <= not a;
    layer0_outputs(1665) <= not (a xor b);
    layer0_outputs(1666) <= not (a and b);
    layer0_outputs(1667) <= a and b;
    layer0_outputs(1668) <= a xor b;
    layer0_outputs(1669) <= b;
    layer0_outputs(1670) <= not (a xor b);
    layer0_outputs(1671) <= b;
    layer0_outputs(1672) <= not a or b;
    layer0_outputs(1673) <= not a;
    layer0_outputs(1674) <= not (a or b);
    layer0_outputs(1675) <= a or b;
    layer0_outputs(1676) <= not (a xor b);
    layer0_outputs(1677) <= not (a xor b);
    layer0_outputs(1678) <= not a or b;
    layer0_outputs(1679) <= not b;
    layer0_outputs(1680) <= not (a xor b);
    layer0_outputs(1681) <= b and not a;
    layer0_outputs(1682) <= a xor b;
    layer0_outputs(1683) <= not (a or b);
    layer0_outputs(1684) <= not (a and b);
    layer0_outputs(1685) <= a xor b;
    layer0_outputs(1686) <= not (a xor b);
    layer0_outputs(1687) <= not a;
    layer0_outputs(1688) <= not (a or b);
    layer0_outputs(1689) <= not (a and b);
    layer0_outputs(1690) <= not a;
    layer0_outputs(1691) <= a;
    layer0_outputs(1692) <= a and not b;
    layer0_outputs(1693) <= not a or b;
    layer0_outputs(1694) <= not b;
    layer0_outputs(1695) <= a and b;
    layer0_outputs(1696) <= not b or a;
    layer0_outputs(1697) <= a and not b;
    layer0_outputs(1698) <= not (a and b);
    layer0_outputs(1699) <= b and not a;
    layer0_outputs(1700) <= not b or a;
    layer0_outputs(1701) <= not (a or b);
    layer0_outputs(1702) <= not b;
    layer0_outputs(1703) <= b;
    layer0_outputs(1704) <= not b;
    layer0_outputs(1705) <= b;
    layer0_outputs(1706) <= a;
    layer0_outputs(1707) <= not (a or b);
    layer0_outputs(1708) <= a xor b;
    layer0_outputs(1709) <= a or b;
    layer0_outputs(1710) <= not b or a;
    layer0_outputs(1711) <= not (a and b);
    layer0_outputs(1712) <= not a;
    layer0_outputs(1713) <= not (a xor b);
    layer0_outputs(1714) <= not b;
    layer0_outputs(1715) <= a;
    layer0_outputs(1716) <= b;
    layer0_outputs(1717) <= b and not a;
    layer0_outputs(1718) <= not b or a;
    layer0_outputs(1719) <= not a;
    layer0_outputs(1720) <= b;
    layer0_outputs(1721) <= not (a and b);
    layer0_outputs(1722) <= not (a and b);
    layer0_outputs(1723) <= not (a or b);
    layer0_outputs(1724) <= a or b;
    layer0_outputs(1725) <= not b or a;
    layer0_outputs(1726) <= not a or b;
    layer0_outputs(1727) <= not (a or b);
    layer0_outputs(1728) <= b;
    layer0_outputs(1729) <= not a or b;
    layer0_outputs(1730) <= b;
    layer0_outputs(1731) <= a or b;
    layer0_outputs(1732) <= 1'b1;
    layer0_outputs(1733) <= b;
    layer0_outputs(1734) <= not a or b;
    layer0_outputs(1735) <= not a;
    layer0_outputs(1736) <= a;
    layer0_outputs(1737) <= b and not a;
    layer0_outputs(1738) <= 1'b1;
    layer0_outputs(1739) <= not b;
    layer0_outputs(1740) <= not (a xor b);
    layer0_outputs(1741) <= not a;
    layer0_outputs(1742) <= b;
    layer0_outputs(1743) <= not a or b;
    layer0_outputs(1744) <= not (a xor b);
    layer0_outputs(1745) <= a xor b;
    layer0_outputs(1746) <= not (a and b);
    layer0_outputs(1747) <= not (a xor b);
    layer0_outputs(1748) <= a or b;
    layer0_outputs(1749) <= b and not a;
    layer0_outputs(1750) <= not b;
    layer0_outputs(1751) <= not a or b;
    layer0_outputs(1752) <= not a or b;
    layer0_outputs(1753) <= a;
    layer0_outputs(1754) <= a xor b;
    layer0_outputs(1755) <= b;
    layer0_outputs(1756) <= not a or b;
    layer0_outputs(1757) <= not (a or b);
    layer0_outputs(1758) <= not a;
    layer0_outputs(1759) <= a or b;
    layer0_outputs(1760) <= a and not b;
    layer0_outputs(1761) <= not b;
    layer0_outputs(1762) <= not a;
    layer0_outputs(1763) <= b;
    layer0_outputs(1764) <= a;
    layer0_outputs(1765) <= a xor b;
    layer0_outputs(1766) <= a or b;
    layer0_outputs(1767) <= not (a xor b);
    layer0_outputs(1768) <= a and b;
    layer0_outputs(1769) <= 1'b1;
    layer0_outputs(1770) <= not b;
    layer0_outputs(1771) <= a and b;
    layer0_outputs(1772) <= not a or b;
    layer0_outputs(1773) <= not (a or b);
    layer0_outputs(1774) <= not b or a;
    layer0_outputs(1775) <= not (a or b);
    layer0_outputs(1776) <= not (a or b);
    layer0_outputs(1777) <= b;
    layer0_outputs(1778) <= not a;
    layer0_outputs(1779) <= not b;
    layer0_outputs(1780) <= a;
    layer0_outputs(1781) <= not a;
    layer0_outputs(1782) <= a and b;
    layer0_outputs(1783) <= a;
    layer0_outputs(1784) <= a and not b;
    layer0_outputs(1785) <= not (a and b);
    layer0_outputs(1786) <= not b;
    layer0_outputs(1787) <= not a;
    layer0_outputs(1788) <= b and not a;
    layer0_outputs(1789) <= not (a xor b);
    layer0_outputs(1790) <= a xor b;
    layer0_outputs(1791) <= not b;
    layer0_outputs(1792) <= a xor b;
    layer0_outputs(1793) <= not a or b;
    layer0_outputs(1794) <= a or b;
    layer0_outputs(1795) <= not b or a;
    layer0_outputs(1796) <= not (a and b);
    layer0_outputs(1797) <= 1'b0;
    layer0_outputs(1798) <= a or b;
    layer0_outputs(1799) <= not (a or b);
    layer0_outputs(1800) <= a xor b;
    layer0_outputs(1801) <= a;
    layer0_outputs(1802) <= not b;
    layer0_outputs(1803) <= not a or b;
    layer0_outputs(1804) <= not (a or b);
    layer0_outputs(1805) <= a or b;
    layer0_outputs(1806) <= not b or a;
    layer0_outputs(1807) <= a xor b;
    layer0_outputs(1808) <= a xor b;
    layer0_outputs(1809) <= a and not b;
    layer0_outputs(1810) <= not (a xor b);
    layer0_outputs(1811) <= a and not b;
    layer0_outputs(1812) <= not a or b;
    layer0_outputs(1813) <= a or b;
    layer0_outputs(1814) <= not (a or b);
    layer0_outputs(1815) <= b;
    layer0_outputs(1816) <= a and not b;
    layer0_outputs(1817) <= a or b;
    layer0_outputs(1818) <= not (a xor b);
    layer0_outputs(1819) <= a or b;
    layer0_outputs(1820) <= b;
    layer0_outputs(1821) <= a or b;
    layer0_outputs(1822) <= a xor b;
    layer0_outputs(1823) <= not (a and b);
    layer0_outputs(1824) <= b and not a;
    layer0_outputs(1825) <= a or b;
    layer0_outputs(1826) <= a or b;
    layer0_outputs(1827) <= not (a or b);
    layer0_outputs(1828) <= not a;
    layer0_outputs(1829) <= not (a xor b);
    layer0_outputs(1830) <= a;
    layer0_outputs(1831) <= not (a xor b);
    layer0_outputs(1832) <= not a;
    layer0_outputs(1833) <= a or b;
    layer0_outputs(1834) <= not a or b;
    layer0_outputs(1835) <= not b;
    layer0_outputs(1836) <= a;
    layer0_outputs(1837) <= not b or a;
    layer0_outputs(1838) <= a and not b;
    layer0_outputs(1839) <= not (a or b);
    layer0_outputs(1840) <= a and b;
    layer0_outputs(1841) <= not (a or b);
    layer0_outputs(1842) <= not (a xor b);
    layer0_outputs(1843) <= not (a xor b);
    layer0_outputs(1844) <= not b or a;
    layer0_outputs(1845) <= not b or a;
    layer0_outputs(1846) <= b and not a;
    layer0_outputs(1847) <= b;
    layer0_outputs(1848) <= a;
    layer0_outputs(1849) <= a;
    layer0_outputs(1850) <= a xor b;
    layer0_outputs(1851) <= 1'b0;
    layer0_outputs(1852) <= not (a or b);
    layer0_outputs(1853) <= a or b;
    layer0_outputs(1854) <= b;
    layer0_outputs(1855) <= b;
    layer0_outputs(1856) <= not b;
    layer0_outputs(1857) <= a xor b;
    layer0_outputs(1858) <= not a or b;
    layer0_outputs(1859) <= a or b;
    layer0_outputs(1860) <= not (a xor b);
    layer0_outputs(1861) <= 1'b0;
    layer0_outputs(1862) <= b;
    layer0_outputs(1863) <= not a;
    layer0_outputs(1864) <= a xor b;
    layer0_outputs(1865) <= not (a or b);
    layer0_outputs(1866) <= not a or b;
    layer0_outputs(1867) <= not (a or b);
    layer0_outputs(1868) <= not (a or b);
    layer0_outputs(1869) <= not a or b;
    layer0_outputs(1870) <= not (a xor b);
    layer0_outputs(1871) <= not (a or b);
    layer0_outputs(1872) <= not (a or b);
    layer0_outputs(1873) <= b and not a;
    layer0_outputs(1874) <= not (a or b);
    layer0_outputs(1875) <= a or b;
    layer0_outputs(1876) <= not a or b;
    layer0_outputs(1877) <= a and not b;
    layer0_outputs(1878) <= a xor b;
    layer0_outputs(1879) <= not a;
    layer0_outputs(1880) <= b and not a;
    layer0_outputs(1881) <= b and not a;
    layer0_outputs(1882) <= not (a or b);
    layer0_outputs(1883) <= b;
    layer0_outputs(1884) <= a and not b;
    layer0_outputs(1885) <= not a;
    layer0_outputs(1886) <= not b;
    layer0_outputs(1887) <= not (a xor b);
    layer0_outputs(1888) <= not a;
    layer0_outputs(1889) <= a xor b;
    layer0_outputs(1890) <= not a or b;
    layer0_outputs(1891) <= a and b;
    layer0_outputs(1892) <= not (a xor b);
    layer0_outputs(1893) <= a;
    layer0_outputs(1894) <= not b;
    layer0_outputs(1895) <= not b or a;
    layer0_outputs(1896) <= not a;
    layer0_outputs(1897) <= b and not a;
    layer0_outputs(1898) <= not a or b;
    layer0_outputs(1899) <= not (a and b);
    layer0_outputs(1900) <= b and not a;
    layer0_outputs(1901) <= a or b;
    layer0_outputs(1902) <= b and not a;
    layer0_outputs(1903) <= a xor b;
    layer0_outputs(1904) <= a;
    layer0_outputs(1905) <= 1'b0;
    layer0_outputs(1906) <= b and not a;
    layer0_outputs(1907) <= a xor b;
    layer0_outputs(1908) <= a;
    layer0_outputs(1909) <= not (a xor b);
    layer0_outputs(1910) <= a or b;
    layer0_outputs(1911) <= not (a or b);
    layer0_outputs(1912) <= not (a xor b);
    layer0_outputs(1913) <= a xor b;
    layer0_outputs(1914) <= not b;
    layer0_outputs(1915) <= not (a xor b);
    layer0_outputs(1916) <= b;
    layer0_outputs(1917) <= a or b;
    layer0_outputs(1918) <= not (a or b);
    layer0_outputs(1919) <= b;
    layer0_outputs(1920) <= a xor b;
    layer0_outputs(1921) <= not (a or b);
    layer0_outputs(1922) <= not b;
    layer0_outputs(1923) <= not (a xor b);
    layer0_outputs(1924) <= not b;
    layer0_outputs(1925) <= b;
    layer0_outputs(1926) <= not (a or b);
    layer0_outputs(1927) <= not a or b;
    layer0_outputs(1928) <= b;
    layer0_outputs(1929) <= a or b;
    layer0_outputs(1930) <= not a;
    layer0_outputs(1931) <= not (a or b);
    layer0_outputs(1932) <= a or b;
    layer0_outputs(1933) <= not a;
    layer0_outputs(1934) <= not (a and b);
    layer0_outputs(1935) <= not (a or b);
    layer0_outputs(1936) <= not (a and b);
    layer0_outputs(1937) <= not (a xor b);
    layer0_outputs(1938) <= not b;
    layer0_outputs(1939) <= a or b;
    layer0_outputs(1940) <= a or b;
    layer0_outputs(1941) <= not b or a;
    layer0_outputs(1942) <= a and not b;
    layer0_outputs(1943) <= b and not a;
    layer0_outputs(1944) <= a and b;
    layer0_outputs(1945) <= a and not b;
    layer0_outputs(1946) <= not (a or b);
    layer0_outputs(1947) <= not a;
    layer0_outputs(1948) <= 1'b1;
    layer0_outputs(1949) <= not a;
    layer0_outputs(1950) <= a xor b;
    layer0_outputs(1951) <= not b;
    layer0_outputs(1952) <= a xor b;
    layer0_outputs(1953) <= a or b;
    layer0_outputs(1954) <= a or b;
    layer0_outputs(1955) <= 1'b1;
    layer0_outputs(1956) <= a and b;
    layer0_outputs(1957) <= a and b;
    layer0_outputs(1958) <= not (a and b);
    layer0_outputs(1959) <= not b;
    layer0_outputs(1960) <= a;
    layer0_outputs(1961) <= b;
    layer0_outputs(1962) <= not (a or b);
    layer0_outputs(1963) <= a or b;
    layer0_outputs(1964) <= not a;
    layer0_outputs(1965) <= not a;
    layer0_outputs(1966) <= a;
    layer0_outputs(1967) <= 1'b1;
    layer0_outputs(1968) <= a and b;
    layer0_outputs(1969) <= not a or b;
    layer0_outputs(1970) <= not a;
    layer0_outputs(1971) <= a xor b;
    layer0_outputs(1972) <= b;
    layer0_outputs(1973) <= 1'b0;
    layer0_outputs(1974) <= not a;
    layer0_outputs(1975) <= not b or a;
    layer0_outputs(1976) <= a and b;
    layer0_outputs(1977) <= a or b;
    layer0_outputs(1978) <= a or b;
    layer0_outputs(1979) <= not a or b;
    layer0_outputs(1980) <= 1'b1;
    layer0_outputs(1981) <= not a or b;
    layer0_outputs(1982) <= not b;
    layer0_outputs(1983) <= not (a or b);
    layer0_outputs(1984) <= not b or a;
    layer0_outputs(1985) <= a or b;
    layer0_outputs(1986) <= not b;
    layer0_outputs(1987) <= b;
    layer0_outputs(1988) <= not (a xor b);
    layer0_outputs(1989) <= not a;
    layer0_outputs(1990) <= a and not b;
    layer0_outputs(1991) <= not a or b;
    layer0_outputs(1992) <= a or b;
    layer0_outputs(1993) <= b and not a;
    layer0_outputs(1994) <= not b;
    layer0_outputs(1995) <= a;
    layer0_outputs(1996) <= not b or a;
    layer0_outputs(1997) <= not a;
    layer0_outputs(1998) <= not a;
    layer0_outputs(1999) <= not b or a;
    layer0_outputs(2000) <= 1'b1;
    layer0_outputs(2001) <= a and not b;
    layer0_outputs(2002) <= not a or b;
    layer0_outputs(2003) <= not b or a;
    layer0_outputs(2004) <= not a or b;
    layer0_outputs(2005) <= not a;
    layer0_outputs(2006) <= not a;
    layer0_outputs(2007) <= not (a or b);
    layer0_outputs(2008) <= not b or a;
    layer0_outputs(2009) <= not (a xor b);
    layer0_outputs(2010) <= not b or a;
    layer0_outputs(2011) <= b;
    layer0_outputs(2012) <= not b or a;
    layer0_outputs(2013) <= not (a xor b);
    layer0_outputs(2014) <= a or b;
    layer0_outputs(2015) <= a and not b;
    layer0_outputs(2016) <= not b;
    layer0_outputs(2017) <= not (a xor b);
    layer0_outputs(2018) <= not b;
    layer0_outputs(2019) <= not (a xor b);
    layer0_outputs(2020) <= a and not b;
    layer0_outputs(2021) <= not (a or b);
    layer0_outputs(2022) <= a xor b;
    layer0_outputs(2023) <= not a;
    layer0_outputs(2024) <= a and not b;
    layer0_outputs(2025) <= 1'b1;
    layer0_outputs(2026) <= a and b;
    layer0_outputs(2027) <= not (a xor b);
    layer0_outputs(2028) <= a or b;
    layer0_outputs(2029) <= not (a or b);
    layer0_outputs(2030) <= a and not b;
    layer0_outputs(2031) <= not (a and b);
    layer0_outputs(2032) <= a;
    layer0_outputs(2033) <= a;
    layer0_outputs(2034) <= a or b;
    layer0_outputs(2035) <= a;
    layer0_outputs(2036) <= not (a or b);
    layer0_outputs(2037) <= b and not a;
    layer0_outputs(2038) <= not (a or b);
    layer0_outputs(2039) <= a;
    layer0_outputs(2040) <= 1'b0;
    layer0_outputs(2041) <= not a;
    layer0_outputs(2042) <= not (a or b);
    layer0_outputs(2043) <= not b;
    layer0_outputs(2044) <= not (a or b);
    layer0_outputs(2045) <= not (a or b);
    layer0_outputs(2046) <= a or b;
    layer0_outputs(2047) <= not (a or b);
    layer0_outputs(2048) <= 1'b1;
    layer0_outputs(2049) <= not a or b;
    layer0_outputs(2050) <= not (a or b);
    layer0_outputs(2051) <= not (a or b);
    layer0_outputs(2052) <= a xor b;
    layer0_outputs(2053) <= not (a or b);
    layer0_outputs(2054) <= a xor b;
    layer0_outputs(2055) <= not b or a;
    layer0_outputs(2056) <= not (a and b);
    layer0_outputs(2057) <= 1'b0;
    layer0_outputs(2058) <= not b or a;
    layer0_outputs(2059) <= a xor b;
    layer0_outputs(2060) <= a;
    layer0_outputs(2061) <= a xor b;
    layer0_outputs(2062) <= b;
    layer0_outputs(2063) <= a xor b;
    layer0_outputs(2064) <= a;
    layer0_outputs(2065) <= not (a or b);
    layer0_outputs(2066) <= not a;
    layer0_outputs(2067) <= a;
    layer0_outputs(2068) <= a;
    layer0_outputs(2069) <= a;
    layer0_outputs(2070) <= not b or a;
    layer0_outputs(2071) <= not b;
    layer0_outputs(2072) <= not b;
    layer0_outputs(2073) <= not (a and b);
    layer0_outputs(2074) <= not a;
    layer0_outputs(2075) <= b;
    layer0_outputs(2076) <= not (a or b);
    layer0_outputs(2077) <= b and not a;
    layer0_outputs(2078) <= b;
    layer0_outputs(2079) <= not b;
    layer0_outputs(2080) <= a xor b;
    layer0_outputs(2081) <= not b or a;
    layer0_outputs(2082) <= not a or b;
    layer0_outputs(2083) <= a or b;
    layer0_outputs(2084) <= a or b;
    layer0_outputs(2085) <= not a;
    layer0_outputs(2086) <= not a or b;
    layer0_outputs(2087) <= not (a or b);
    layer0_outputs(2088) <= a and not b;
    layer0_outputs(2089) <= not (a or b);
    layer0_outputs(2090) <= not (a and b);
    layer0_outputs(2091) <= not a;
    layer0_outputs(2092) <= not (a and b);
    layer0_outputs(2093) <= a or b;
    layer0_outputs(2094) <= a;
    layer0_outputs(2095) <= not (a or b);
    layer0_outputs(2096) <= not a;
    layer0_outputs(2097) <= not b;
    layer0_outputs(2098) <= not (a or b);
    layer0_outputs(2099) <= a and not b;
    layer0_outputs(2100) <= not (a xor b);
    layer0_outputs(2101) <= a and b;
    layer0_outputs(2102) <= a or b;
    layer0_outputs(2103) <= not b;
    layer0_outputs(2104) <= 1'b1;
    layer0_outputs(2105) <= a and not b;
    layer0_outputs(2106) <= b and not a;
    layer0_outputs(2107) <= a or b;
    layer0_outputs(2108) <= a and not b;
    layer0_outputs(2109) <= not b or a;
    layer0_outputs(2110) <= b and not a;
    layer0_outputs(2111) <= a or b;
    layer0_outputs(2112) <= not a;
    layer0_outputs(2113) <= not (a or b);
    layer0_outputs(2114) <= 1'b1;
    layer0_outputs(2115) <= not (a xor b);
    layer0_outputs(2116) <= a or b;
    layer0_outputs(2117) <= b;
    layer0_outputs(2118) <= a xor b;
    layer0_outputs(2119) <= not a;
    layer0_outputs(2120) <= 1'b1;
    layer0_outputs(2121) <= not (a or b);
    layer0_outputs(2122) <= b;
    layer0_outputs(2123) <= not b or a;
    layer0_outputs(2124) <= not a;
    layer0_outputs(2125) <= not b or a;
    layer0_outputs(2126) <= not a or b;
    layer0_outputs(2127) <= b;
    layer0_outputs(2128) <= a and not b;
    layer0_outputs(2129) <= not b;
    layer0_outputs(2130) <= not (a xor b);
    layer0_outputs(2131) <= a xor b;
    layer0_outputs(2132) <= a or b;
    layer0_outputs(2133) <= 1'b1;
    layer0_outputs(2134) <= not a;
    layer0_outputs(2135) <= not b or a;
    layer0_outputs(2136) <= b and not a;
    layer0_outputs(2137) <= not (a xor b);
    layer0_outputs(2138) <= not a;
    layer0_outputs(2139) <= a;
    layer0_outputs(2140) <= b and not a;
    layer0_outputs(2141) <= not (a or b);
    layer0_outputs(2142) <= a or b;
    layer0_outputs(2143) <= not b;
    layer0_outputs(2144) <= a and not b;
    layer0_outputs(2145) <= not (a or b);
    layer0_outputs(2146) <= a xor b;
    layer0_outputs(2147) <= not (a or b);
    layer0_outputs(2148) <= not (a or b);
    layer0_outputs(2149) <= b;
    layer0_outputs(2150) <= not b or a;
    layer0_outputs(2151) <= a or b;
    layer0_outputs(2152) <= a and not b;
    layer0_outputs(2153) <= a;
    layer0_outputs(2154) <= not a or b;
    layer0_outputs(2155) <= not (a or b);
    layer0_outputs(2156) <= 1'b1;
    layer0_outputs(2157) <= 1'b0;
    layer0_outputs(2158) <= b;
    layer0_outputs(2159) <= b and not a;
    layer0_outputs(2160) <= not a;
    layer0_outputs(2161) <= not b;
    layer0_outputs(2162) <= not (a xor b);
    layer0_outputs(2163) <= a or b;
    layer0_outputs(2164) <= not a;
    layer0_outputs(2165) <= not b or a;
    layer0_outputs(2166) <= not b;
    layer0_outputs(2167) <= not (a or b);
    layer0_outputs(2168) <= not b;
    layer0_outputs(2169) <= b;
    layer0_outputs(2170) <= b and not a;
    layer0_outputs(2171) <= not (a or b);
    layer0_outputs(2172) <= not a;
    layer0_outputs(2173) <= 1'b1;
    layer0_outputs(2174) <= a;
    layer0_outputs(2175) <= not b;
    layer0_outputs(2176) <= a and not b;
    layer0_outputs(2177) <= not (a or b);
    layer0_outputs(2178) <= 1'b0;
    layer0_outputs(2179) <= not b;
    layer0_outputs(2180) <= not a;
    layer0_outputs(2181) <= not a or b;
    layer0_outputs(2182) <= not a or b;
    layer0_outputs(2183) <= not (a or b);
    layer0_outputs(2184) <= not b;
    layer0_outputs(2185) <= a;
    layer0_outputs(2186) <= a xor b;
    layer0_outputs(2187) <= b;
    layer0_outputs(2188) <= b and not a;
    layer0_outputs(2189) <= not a;
    layer0_outputs(2190) <= b;
    layer0_outputs(2191) <= a;
    layer0_outputs(2192) <= 1'b0;
    layer0_outputs(2193) <= a;
    layer0_outputs(2194) <= b;
    layer0_outputs(2195) <= not (a xor b);
    layer0_outputs(2196) <= b and not a;
    layer0_outputs(2197) <= not a or b;
    layer0_outputs(2198) <= a xor b;
    layer0_outputs(2199) <= a and not b;
    layer0_outputs(2200) <= not b or a;
    layer0_outputs(2201) <= a xor b;
    layer0_outputs(2202) <= a xor b;
    layer0_outputs(2203) <= a xor b;
    layer0_outputs(2204) <= b and not a;
    layer0_outputs(2205) <= b;
    layer0_outputs(2206) <= b and not a;
    layer0_outputs(2207) <= not a;
    layer0_outputs(2208) <= not a or b;
    layer0_outputs(2209) <= b and not a;
    layer0_outputs(2210) <= not (a or b);
    layer0_outputs(2211) <= b and not a;
    layer0_outputs(2212) <= not (a xor b);
    layer0_outputs(2213) <= a;
    layer0_outputs(2214) <= not b;
    layer0_outputs(2215) <= b;
    layer0_outputs(2216) <= b;
    layer0_outputs(2217) <= not (a xor b);
    layer0_outputs(2218) <= a and not b;
    layer0_outputs(2219) <= a xor b;
    layer0_outputs(2220) <= not a;
    layer0_outputs(2221) <= not a;
    layer0_outputs(2222) <= a or b;
    layer0_outputs(2223) <= not b;
    layer0_outputs(2224) <= a xor b;
    layer0_outputs(2225) <= a or b;
    layer0_outputs(2226) <= b and not a;
    layer0_outputs(2227) <= not b;
    layer0_outputs(2228) <= not b;
    layer0_outputs(2229) <= not a or b;
    layer0_outputs(2230) <= not (a and b);
    layer0_outputs(2231) <= a and not b;
    layer0_outputs(2232) <= a or b;
    layer0_outputs(2233) <= b and not a;
    layer0_outputs(2234) <= a xor b;
    layer0_outputs(2235) <= not b or a;
    layer0_outputs(2236) <= 1'b1;
    layer0_outputs(2237) <= not a or b;
    layer0_outputs(2238) <= not (a or b);
    layer0_outputs(2239) <= not a;
    layer0_outputs(2240) <= not (a and b);
    layer0_outputs(2241) <= a or b;
    layer0_outputs(2242) <= a xor b;
    layer0_outputs(2243) <= a;
    layer0_outputs(2244) <= not b or a;
    layer0_outputs(2245) <= a or b;
    layer0_outputs(2246) <= not b;
    layer0_outputs(2247) <= not (a and b);
    layer0_outputs(2248) <= not (a or b);
    layer0_outputs(2249) <= a xor b;
    layer0_outputs(2250) <= not (a or b);
    layer0_outputs(2251) <= not b or a;
    layer0_outputs(2252) <= not (a and b);
    layer0_outputs(2253) <= a or b;
    layer0_outputs(2254) <= not (a xor b);
    layer0_outputs(2255) <= not (a or b);
    layer0_outputs(2256) <= a xor b;
    layer0_outputs(2257) <= not (a or b);
    layer0_outputs(2258) <= a xor b;
    layer0_outputs(2259) <= not (a and b);
    layer0_outputs(2260) <= a xor b;
    layer0_outputs(2261) <= not (a or b);
    layer0_outputs(2262) <= not a;
    layer0_outputs(2263) <= not b or a;
    layer0_outputs(2264) <= b and not a;
    layer0_outputs(2265) <= not a or b;
    layer0_outputs(2266) <= b and not a;
    layer0_outputs(2267) <= not (a or b);
    layer0_outputs(2268) <= a xor b;
    layer0_outputs(2269) <= not a;
    layer0_outputs(2270) <= a or b;
    layer0_outputs(2271) <= a;
    layer0_outputs(2272) <= not b or a;
    layer0_outputs(2273) <= b and not a;
    layer0_outputs(2274) <= not b;
    layer0_outputs(2275) <= b and not a;
    layer0_outputs(2276) <= a or b;
    layer0_outputs(2277) <= a and not b;
    layer0_outputs(2278) <= a or b;
    layer0_outputs(2279) <= 1'b1;
    layer0_outputs(2280) <= a and not b;
    layer0_outputs(2281) <= a xor b;
    layer0_outputs(2282) <= a;
    layer0_outputs(2283) <= not a;
    layer0_outputs(2284) <= a and not b;
    layer0_outputs(2285) <= a xor b;
    layer0_outputs(2286) <= not b;
    layer0_outputs(2287) <= not b or a;
    layer0_outputs(2288) <= not a or b;
    layer0_outputs(2289) <= b and not a;
    layer0_outputs(2290) <= 1'b0;
    layer0_outputs(2291) <= a or b;
    layer0_outputs(2292) <= not (a or b);
    layer0_outputs(2293) <= a and b;
    layer0_outputs(2294) <= not (a or b);
    layer0_outputs(2295) <= b and not a;
    layer0_outputs(2296) <= not b or a;
    layer0_outputs(2297) <= a xor b;
    layer0_outputs(2298) <= 1'b1;
    layer0_outputs(2299) <= not b or a;
    layer0_outputs(2300) <= b and not a;
    layer0_outputs(2301) <= not b;
    layer0_outputs(2302) <= a and not b;
    layer0_outputs(2303) <= a or b;
    layer0_outputs(2304) <= not b;
    layer0_outputs(2305) <= not a;
    layer0_outputs(2306) <= not (a or b);
    layer0_outputs(2307) <= a and not b;
    layer0_outputs(2308) <= a or b;
    layer0_outputs(2309) <= not a or b;
    layer0_outputs(2310) <= a and b;
    layer0_outputs(2311) <= a xor b;
    layer0_outputs(2312) <= a or b;
    layer0_outputs(2313) <= not a or b;
    layer0_outputs(2314) <= a and not b;
    layer0_outputs(2315) <= not (a xor b);
    layer0_outputs(2316) <= not b;
    layer0_outputs(2317) <= a;
    layer0_outputs(2318) <= 1'b0;
    layer0_outputs(2319) <= not (a or b);
    layer0_outputs(2320) <= a or b;
    layer0_outputs(2321) <= not b or a;
    layer0_outputs(2322) <= a and not b;
    layer0_outputs(2323) <= not (a xor b);
    layer0_outputs(2324) <= a and not b;
    layer0_outputs(2325) <= not a;
    layer0_outputs(2326) <= not a;
    layer0_outputs(2327) <= a and b;
    layer0_outputs(2328) <= a;
    layer0_outputs(2329) <= not b or a;
    layer0_outputs(2330) <= not (a xor b);
    layer0_outputs(2331) <= not b or a;
    layer0_outputs(2332) <= not b;
    layer0_outputs(2333) <= b and not a;
    layer0_outputs(2334) <= a or b;
    layer0_outputs(2335) <= a;
    layer0_outputs(2336) <= a or b;
    layer0_outputs(2337) <= not (a xor b);
    layer0_outputs(2338) <= a xor b;
    layer0_outputs(2339) <= not a;
    layer0_outputs(2340) <= not a;
    layer0_outputs(2341) <= b and not a;
    layer0_outputs(2342) <= not (a or b);
    layer0_outputs(2343) <= a xor b;
    layer0_outputs(2344) <= b and not a;
    layer0_outputs(2345) <= not (a or b);
    layer0_outputs(2346) <= not (a or b);
    layer0_outputs(2347) <= not (a and b);
    layer0_outputs(2348) <= not b;
    layer0_outputs(2349) <= not (a xor b);
    layer0_outputs(2350) <= b;
    layer0_outputs(2351) <= 1'b0;
    layer0_outputs(2352) <= not a or b;
    layer0_outputs(2353) <= b;
    layer0_outputs(2354) <= b;
    layer0_outputs(2355) <= not b or a;
    layer0_outputs(2356) <= a xor b;
    layer0_outputs(2357) <= a and b;
    layer0_outputs(2358) <= not a;
    layer0_outputs(2359) <= not (a or b);
    layer0_outputs(2360) <= a or b;
    layer0_outputs(2361) <= a xor b;
    layer0_outputs(2362) <= a or b;
    layer0_outputs(2363) <= a or b;
    layer0_outputs(2364) <= not a;
    layer0_outputs(2365) <= a;
    layer0_outputs(2366) <= not b;
    layer0_outputs(2367) <= a or b;
    layer0_outputs(2368) <= a and b;
    layer0_outputs(2369) <= a xor b;
    layer0_outputs(2370) <= a or b;
    layer0_outputs(2371) <= a or b;
    layer0_outputs(2372) <= a and not b;
    layer0_outputs(2373) <= not (a or b);
    layer0_outputs(2374) <= not b;
    layer0_outputs(2375) <= a and not b;
    layer0_outputs(2376) <= not (a or b);
    layer0_outputs(2377) <= not b or a;
    layer0_outputs(2378) <= not b or a;
    layer0_outputs(2379) <= a and not b;
    layer0_outputs(2380) <= not (a and b);
    layer0_outputs(2381) <= not (a or b);
    layer0_outputs(2382) <= a and b;
    layer0_outputs(2383) <= a or b;
    layer0_outputs(2384) <= a;
    layer0_outputs(2385) <= 1'b1;
    layer0_outputs(2386) <= not (a xor b);
    layer0_outputs(2387) <= not b or a;
    layer0_outputs(2388) <= not (a xor b);
    layer0_outputs(2389) <= 1'b0;
    layer0_outputs(2390) <= not a or b;
    layer0_outputs(2391) <= not a;
    layer0_outputs(2392) <= a or b;
    layer0_outputs(2393) <= a xor b;
    layer0_outputs(2394) <= a and not b;
    layer0_outputs(2395) <= a;
    layer0_outputs(2396) <= a;
    layer0_outputs(2397) <= not (a or b);
    layer0_outputs(2398) <= a and b;
    layer0_outputs(2399) <= a and not b;
    layer0_outputs(2400) <= b and not a;
    layer0_outputs(2401) <= not b or a;
    layer0_outputs(2402) <= not (a or b);
    layer0_outputs(2403) <= a and not b;
    layer0_outputs(2404) <= not (a or b);
    layer0_outputs(2405) <= not a or b;
    layer0_outputs(2406) <= not (a xor b);
    layer0_outputs(2407) <= not (a or b);
    layer0_outputs(2408) <= a or b;
    layer0_outputs(2409) <= not a;
    layer0_outputs(2410) <= not b or a;
    layer0_outputs(2411) <= a or b;
    layer0_outputs(2412) <= a and not b;
    layer0_outputs(2413) <= not a;
    layer0_outputs(2414) <= not (a and b);
    layer0_outputs(2415) <= b;
    layer0_outputs(2416) <= a and not b;
    layer0_outputs(2417) <= not a or b;
    layer0_outputs(2418) <= a;
    layer0_outputs(2419) <= not (a or b);
    layer0_outputs(2420) <= a;
    layer0_outputs(2421) <= not (a or b);
    layer0_outputs(2422) <= a and not b;
    layer0_outputs(2423) <= not a or b;
    layer0_outputs(2424) <= a xor b;
    layer0_outputs(2425) <= b and not a;
    layer0_outputs(2426) <= not (a or b);
    layer0_outputs(2427) <= not a;
    layer0_outputs(2428) <= not (a or b);
    layer0_outputs(2429) <= not (a xor b);
    layer0_outputs(2430) <= 1'b0;
    layer0_outputs(2431) <= not (a xor b);
    layer0_outputs(2432) <= not (a or b);
    layer0_outputs(2433) <= a and not b;
    layer0_outputs(2434) <= not (a xor b);
    layer0_outputs(2435) <= not (a xor b);
    layer0_outputs(2436) <= a or b;
    layer0_outputs(2437) <= not a or b;
    layer0_outputs(2438) <= a xor b;
    layer0_outputs(2439) <= a;
    layer0_outputs(2440) <= a or b;
    layer0_outputs(2441) <= a xor b;
    layer0_outputs(2442) <= not (a or b);
    layer0_outputs(2443) <= a or b;
    layer0_outputs(2444) <= not b or a;
    layer0_outputs(2445) <= a xor b;
    layer0_outputs(2446) <= not b or a;
    layer0_outputs(2447) <= 1'b0;
    layer0_outputs(2448) <= not (a xor b);
    layer0_outputs(2449) <= a and not b;
    layer0_outputs(2450) <= not a;
    layer0_outputs(2451) <= not (a or b);
    layer0_outputs(2452) <= not b;
    layer0_outputs(2453) <= not b;
    layer0_outputs(2454) <= not a;
    layer0_outputs(2455) <= b and not a;
    layer0_outputs(2456) <= not (a and b);
    layer0_outputs(2457) <= a xor b;
    layer0_outputs(2458) <= not (a or b);
    layer0_outputs(2459) <= not (a or b);
    layer0_outputs(2460) <= a and b;
    layer0_outputs(2461) <= not b or a;
    layer0_outputs(2462) <= a xor b;
    layer0_outputs(2463) <= a and b;
    layer0_outputs(2464) <= 1'b1;
    layer0_outputs(2465) <= a xor b;
    layer0_outputs(2466) <= a or b;
    layer0_outputs(2467) <= a xor b;
    layer0_outputs(2468) <= not (a and b);
    layer0_outputs(2469) <= b;
    layer0_outputs(2470) <= not a or b;
    layer0_outputs(2471) <= b;
    layer0_outputs(2472) <= b;
    layer0_outputs(2473) <= not (a or b);
    layer0_outputs(2474) <= 1'b0;
    layer0_outputs(2475) <= not (a or b);
    layer0_outputs(2476) <= not a;
    layer0_outputs(2477) <= a or b;
    layer0_outputs(2478) <= b and not a;
    layer0_outputs(2479) <= a and not b;
    layer0_outputs(2480) <= not a or b;
    layer0_outputs(2481) <= not a or b;
    layer0_outputs(2482) <= not b;
    layer0_outputs(2483) <= b;
    layer0_outputs(2484) <= not (a xor b);
    layer0_outputs(2485) <= not a or b;
    layer0_outputs(2486) <= a xor b;
    layer0_outputs(2487) <= b and not a;
    layer0_outputs(2488) <= not a;
    layer0_outputs(2489) <= not (a or b);
    layer0_outputs(2490) <= a;
    layer0_outputs(2491) <= a and not b;
    layer0_outputs(2492) <= not (a and b);
    layer0_outputs(2493) <= not (a or b);
    layer0_outputs(2494) <= not a or b;
    layer0_outputs(2495) <= not (a or b);
    layer0_outputs(2496) <= a and b;
    layer0_outputs(2497) <= a xor b;
    layer0_outputs(2498) <= a xor b;
    layer0_outputs(2499) <= not b;
    layer0_outputs(2500) <= a;
    layer0_outputs(2501) <= a xor b;
    layer0_outputs(2502) <= b and not a;
    layer0_outputs(2503) <= not b;
    layer0_outputs(2504) <= b;
    layer0_outputs(2505) <= 1'b0;
    layer0_outputs(2506) <= not a or b;
    layer0_outputs(2507) <= a xor b;
    layer0_outputs(2508) <= not (a or b);
    layer0_outputs(2509) <= b and not a;
    layer0_outputs(2510) <= b;
    layer0_outputs(2511) <= b;
    layer0_outputs(2512) <= not b or a;
    layer0_outputs(2513) <= a;
    layer0_outputs(2514) <= a or b;
    layer0_outputs(2515) <= not a;
    layer0_outputs(2516) <= a or b;
    layer0_outputs(2517) <= not b;
    layer0_outputs(2518) <= a and not b;
    layer0_outputs(2519) <= a xor b;
    layer0_outputs(2520) <= not (a xor b);
    layer0_outputs(2521) <= not (a xor b);
    layer0_outputs(2522) <= not (a or b);
    layer0_outputs(2523) <= not a or b;
    layer0_outputs(2524) <= not (a or b);
    layer0_outputs(2525) <= not b;
    layer0_outputs(2526) <= not (a xor b);
    layer0_outputs(2527) <= a;
    layer0_outputs(2528) <= b;
    layer0_outputs(2529) <= a and not b;
    layer0_outputs(2530) <= a and not b;
    layer0_outputs(2531) <= b;
    layer0_outputs(2532) <= not b;
    layer0_outputs(2533) <= a or b;
    layer0_outputs(2534) <= 1'b0;
    layer0_outputs(2535) <= a xor b;
    layer0_outputs(2536) <= a;
    layer0_outputs(2537) <= b and not a;
    layer0_outputs(2538) <= a and not b;
    layer0_outputs(2539) <= a xor b;
    layer0_outputs(2540) <= not b or a;
    layer0_outputs(2541) <= not a or b;
    layer0_outputs(2542) <= b;
    layer0_outputs(2543) <= not a or b;
    layer0_outputs(2544) <= b;
    layer0_outputs(2545) <= not a or b;
    layer0_outputs(2546) <= a xor b;
    layer0_outputs(2547) <= 1'b1;
    layer0_outputs(2548) <= not (a or b);
    layer0_outputs(2549) <= a;
    layer0_outputs(2550) <= a xor b;
    layer0_outputs(2551) <= not (a or b);
    layer0_outputs(2552) <= not (a or b);
    layer0_outputs(2553) <= a or b;
    layer0_outputs(2554) <= not (a and b);
    layer0_outputs(2555) <= a;
    layer0_outputs(2556) <= a or b;
    layer0_outputs(2557) <= not b or a;
    layer0_outputs(2558) <= not (a xor b);
    layer0_outputs(2559) <= b;
    layer0_outputs(2560) <= not a or b;
    layer0_outputs(2561) <= a or b;
    layer0_outputs(2562) <= not a;
    layer0_outputs(2563) <= not a;
    layer0_outputs(2564) <= not a;
    layer0_outputs(2565) <= not (a or b);
    layer0_outputs(2566) <= not a or b;
    layer0_outputs(2567) <= b;
    layer0_outputs(2568) <= b;
    layer0_outputs(2569) <= b;
    layer0_outputs(2570) <= a or b;
    layer0_outputs(2571) <= a and not b;
    layer0_outputs(2572) <= 1'b0;
    layer0_outputs(2573) <= a;
    layer0_outputs(2574) <= not b;
    layer0_outputs(2575) <= not (a or b);
    layer0_outputs(2576) <= b;
    layer0_outputs(2577) <= not (a or b);
    layer0_outputs(2578) <= b and not a;
    layer0_outputs(2579) <= a or b;
    layer0_outputs(2580) <= a or b;
    layer0_outputs(2581) <= not (a xor b);
    layer0_outputs(2582) <= a or b;
    layer0_outputs(2583) <= not a or b;
    layer0_outputs(2584) <= b;
    layer0_outputs(2585) <= a and not b;
    layer0_outputs(2586) <= a;
    layer0_outputs(2587) <= a or b;
    layer0_outputs(2588) <= a and b;
    layer0_outputs(2589) <= not b or a;
    layer0_outputs(2590) <= a xor b;
    layer0_outputs(2591) <= not (a xor b);
    layer0_outputs(2592) <= not (a xor b);
    layer0_outputs(2593) <= b;
    layer0_outputs(2594) <= not (a xor b);
    layer0_outputs(2595) <= not a;
    layer0_outputs(2596) <= not b or a;
    layer0_outputs(2597) <= not b;
    layer0_outputs(2598) <= a;
    layer0_outputs(2599) <= 1'b0;
    layer0_outputs(2600) <= a or b;
    layer0_outputs(2601) <= not b;
    layer0_outputs(2602) <= a or b;
    layer0_outputs(2603) <= not b or a;
    layer0_outputs(2604) <= b;
    layer0_outputs(2605) <= a xor b;
    layer0_outputs(2606) <= b;
    layer0_outputs(2607) <= a or b;
    layer0_outputs(2608) <= 1'b0;
    layer0_outputs(2609) <= a;
    layer0_outputs(2610) <= 1'b1;
    layer0_outputs(2611) <= not (a or b);
    layer0_outputs(2612) <= not a or b;
    layer0_outputs(2613) <= a and not b;
    layer0_outputs(2614) <= not (a and b);
    layer0_outputs(2615) <= a xor b;
    layer0_outputs(2616) <= a and not b;
    layer0_outputs(2617) <= a;
    layer0_outputs(2618) <= a or b;
    layer0_outputs(2619) <= b and not a;
    layer0_outputs(2620) <= a xor b;
    layer0_outputs(2621) <= a xor b;
    layer0_outputs(2622) <= not a;
    layer0_outputs(2623) <= not a or b;
    layer0_outputs(2624) <= a or b;
    layer0_outputs(2625) <= not b;
    layer0_outputs(2626) <= b and not a;
    layer0_outputs(2627) <= b;
    layer0_outputs(2628) <= a xor b;
    layer0_outputs(2629) <= b and not a;
    layer0_outputs(2630) <= not a or b;
    layer0_outputs(2631) <= a and b;
    layer0_outputs(2632) <= not b or a;
    layer0_outputs(2633) <= not (a or b);
    layer0_outputs(2634) <= not b;
    layer0_outputs(2635) <= not (a or b);
    layer0_outputs(2636) <= a or b;
    layer0_outputs(2637) <= not a;
    layer0_outputs(2638) <= not a;
    layer0_outputs(2639) <= a;
    layer0_outputs(2640) <= a xor b;
    layer0_outputs(2641) <= a and b;
    layer0_outputs(2642) <= not b;
    layer0_outputs(2643) <= not a or b;
    layer0_outputs(2644) <= not a or b;
    layer0_outputs(2645) <= a;
    layer0_outputs(2646) <= a and b;
    layer0_outputs(2647) <= a or b;
    layer0_outputs(2648) <= not b or a;
    layer0_outputs(2649) <= b and not a;
    layer0_outputs(2650) <= b and not a;
    layer0_outputs(2651) <= a;
    layer0_outputs(2652) <= b;
    layer0_outputs(2653) <= a and b;
    layer0_outputs(2654) <= not b;
    layer0_outputs(2655) <= a xor b;
    layer0_outputs(2656) <= not b;
    layer0_outputs(2657) <= a;
    layer0_outputs(2658) <= not (a and b);
    layer0_outputs(2659) <= not (a or b);
    layer0_outputs(2660) <= a and not b;
    layer0_outputs(2661) <= not (a xor b);
    layer0_outputs(2662) <= not (a xor b);
    layer0_outputs(2663) <= not (a or b);
    layer0_outputs(2664) <= a and not b;
    layer0_outputs(2665) <= a and not b;
    layer0_outputs(2666) <= not a;
    layer0_outputs(2667) <= not (a xor b);
    layer0_outputs(2668) <= not b or a;
    layer0_outputs(2669) <= a or b;
    layer0_outputs(2670) <= a and b;
    layer0_outputs(2671) <= not a;
    layer0_outputs(2672) <= not b;
    layer0_outputs(2673) <= not a;
    layer0_outputs(2674) <= 1'b1;
    layer0_outputs(2675) <= a and not b;
    layer0_outputs(2676) <= a xor b;
    layer0_outputs(2677) <= not (a or b);
    layer0_outputs(2678) <= b;
    layer0_outputs(2679) <= a and b;
    layer0_outputs(2680) <= b;
    layer0_outputs(2681) <= a or b;
    layer0_outputs(2682) <= a xor b;
    layer0_outputs(2683) <= not a;
    layer0_outputs(2684) <= a xor b;
    layer0_outputs(2685) <= b;
    layer0_outputs(2686) <= not a or b;
    layer0_outputs(2687) <= not b or a;
    layer0_outputs(2688) <= not (a or b);
    layer0_outputs(2689) <= a;
    layer0_outputs(2690) <= not a or b;
    layer0_outputs(2691) <= not (a or b);
    layer0_outputs(2692) <= b and not a;
    layer0_outputs(2693) <= not b;
    layer0_outputs(2694) <= a or b;
    layer0_outputs(2695) <= not b or a;
    layer0_outputs(2696) <= not (a xor b);
    layer0_outputs(2697) <= a or b;
    layer0_outputs(2698) <= not (a xor b);
    layer0_outputs(2699) <= not b;
    layer0_outputs(2700) <= not (a and b);
    layer0_outputs(2701) <= a xor b;
    layer0_outputs(2702) <= not (a or b);
    layer0_outputs(2703) <= a or b;
    layer0_outputs(2704) <= not (a or b);
    layer0_outputs(2705) <= not (a xor b);
    layer0_outputs(2706) <= not b or a;
    layer0_outputs(2707) <= not b or a;
    layer0_outputs(2708) <= not (a and b);
    layer0_outputs(2709) <= not a;
    layer0_outputs(2710) <= a;
    layer0_outputs(2711) <= a;
    layer0_outputs(2712) <= a or b;
    layer0_outputs(2713) <= a or b;
    layer0_outputs(2714) <= not a;
    layer0_outputs(2715) <= a;
    layer0_outputs(2716) <= not b;
    layer0_outputs(2717) <= a;
    layer0_outputs(2718) <= not (a xor b);
    layer0_outputs(2719) <= not b;
    layer0_outputs(2720) <= a;
    layer0_outputs(2721) <= a xor b;
    layer0_outputs(2722) <= b;
    layer0_outputs(2723) <= not a or b;
    layer0_outputs(2724) <= not b;
    layer0_outputs(2725) <= not b;
    layer0_outputs(2726) <= a or b;
    layer0_outputs(2727) <= b;
    layer0_outputs(2728) <= not (a xor b);
    layer0_outputs(2729) <= a;
    layer0_outputs(2730) <= a and not b;
    layer0_outputs(2731) <= not b or a;
    layer0_outputs(2732) <= a or b;
    layer0_outputs(2733) <= a or b;
    layer0_outputs(2734) <= not b;
    layer0_outputs(2735) <= not a;
    layer0_outputs(2736) <= not (a or b);
    layer0_outputs(2737) <= not (a or b);
    layer0_outputs(2738) <= not (a xor b);
    layer0_outputs(2739) <= b and not a;
    layer0_outputs(2740) <= a or b;
    layer0_outputs(2741) <= a xor b;
    layer0_outputs(2742) <= a;
    layer0_outputs(2743) <= a or b;
    layer0_outputs(2744) <= not a;
    layer0_outputs(2745) <= not (a xor b);
    layer0_outputs(2746) <= 1'b1;
    layer0_outputs(2747) <= not (a or b);
    layer0_outputs(2748) <= not b;
    layer0_outputs(2749) <= not a;
    layer0_outputs(2750) <= not (a or b);
    layer0_outputs(2751) <= a and not b;
    layer0_outputs(2752) <= not b or a;
    layer0_outputs(2753) <= not (a or b);
    layer0_outputs(2754) <= not a or b;
    layer0_outputs(2755) <= 1'b0;
    layer0_outputs(2756) <= a and b;
    layer0_outputs(2757) <= a or b;
    layer0_outputs(2758) <= a or b;
    layer0_outputs(2759) <= not a;
    layer0_outputs(2760) <= b;
    layer0_outputs(2761) <= not (a xor b);
    layer0_outputs(2762) <= a or b;
    layer0_outputs(2763) <= not a or b;
    layer0_outputs(2764) <= a or b;
    layer0_outputs(2765) <= a xor b;
    layer0_outputs(2766) <= 1'b0;
    layer0_outputs(2767) <= 1'b0;
    layer0_outputs(2768) <= not (a xor b);
    layer0_outputs(2769) <= not (a xor b);
    layer0_outputs(2770) <= a and b;
    layer0_outputs(2771) <= not b;
    layer0_outputs(2772) <= not (a or b);
    layer0_outputs(2773) <= not (a and b);
    layer0_outputs(2774) <= not a or b;
    layer0_outputs(2775) <= a and not b;
    layer0_outputs(2776) <= b;
    layer0_outputs(2777) <= not (a and b);
    layer0_outputs(2778) <= b;
    layer0_outputs(2779) <= a or b;
    layer0_outputs(2780) <= not (a or b);
    layer0_outputs(2781) <= not b;
    layer0_outputs(2782) <= not (a or b);
    layer0_outputs(2783) <= b;
    layer0_outputs(2784) <= b and not a;
    layer0_outputs(2785) <= not (a or b);
    layer0_outputs(2786) <= not (a or b);
    layer0_outputs(2787) <= not b;
    layer0_outputs(2788) <= b and not a;
    layer0_outputs(2789) <= not b;
    layer0_outputs(2790) <= not (a or b);
    layer0_outputs(2791) <= not b or a;
    layer0_outputs(2792) <= b and not a;
    layer0_outputs(2793) <= a;
    layer0_outputs(2794) <= b;
    layer0_outputs(2795) <= not a or b;
    layer0_outputs(2796) <= a;
    layer0_outputs(2797) <= not b;
    layer0_outputs(2798) <= a or b;
    layer0_outputs(2799) <= 1'b0;
    layer0_outputs(2800) <= not a;
    layer0_outputs(2801) <= not (a xor b);
    layer0_outputs(2802) <= a and not b;
    layer0_outputs(2803) <= a or b;
    layer0_outputs(2804) <= not (a or b);
    layer0_outputs(2805) <= not (a or b);
    layer0_outputs(2806) <= b;
    layer0_outputs(2807) <= a xor b;
    layer0_outputs(2808) <= a or b;
    layer0_outputs(2809) <= not b or a;
    layer0_outputs(2810) <= not a or b;
    layer0_outputs(2811) <= not b or a;
    layer0_outputs(2812) <= a xor b;
    layer0_outputs(2813) <= a;
    layer0_outputs(2814) <= not a;
    layer0_outputs(2815) <= b and not a;
    layer0_outputs(2816) <= not b;
    layer0_outputs(2817) <= a and not b;
    layer0_outputs(2818) <= not (a and b);
    layer0_outputs(2819) <= a xor b;
    layer0_outputs(2820) <= a and not b;
    layer0_outputs(2821) <= not b;
    layer0_outputs(2822) <= a and not b;
    layer0_outputs(2823) <= b and not a;
    layer0_outputs(2824) <= not (a xor b);
    layer0_outputs(2825) <= not b;
    layer0_outputs(2826) <= not (a or b);
    layer0_outputs(2827) <= not (a or b);
    layer0_outputs(2828) <= b and not a;
    layer0_outputs(2829) <= a xor b;
    layer0_outputs(2830) <= a and not b;
    layer0_outputs(2831) <= a or b;
    layer0_outputs(2832) <= a xor b;
    layer0_outputs(2833) <= a or b;
    layer0_outputs(2834) <= a or b;
    layer0_outputs(2835) <= a xor b;
    layer0_outputs(2836) <= a or b;
    layer0_outputs(2837) <= not (a or b);
    layer0_outputs(2838) <= b and not a;
    layer0_outputs(2839) <= not b;
    layer0_outputs(2840) <= not a;
    layer0_outputs(2841) <= not b;
    layer0_outputs(2842) <= not a;
    layer0_outputs(2843) <= a xor b;
    layer0_outputs(2844) <= 1'b0;
    layer0_outputs(2845) <= not (a and b);
    layer0_outputs(2846) <= b;
    layer0_outputs(2847) <= not (a or b);
    layer0_outputs(2848) <= not a or b;
    layer0_outputs(2849) <= a or b;
    layer0_outputs(2850) <= not b;
    layer0_outputs(2851) <= a and b;
    layer0_outputs(2852) <= not b;
    layer0_outputs(2853) <= not b or a;
    layer0_outputs(2854) <= not b;
    layer0_outputs(2855) <= 1'b1;
    layer0_outputs(2856) <= not (a xor b);
    layer0_outputs(2857) <= not a;
    layer0_outputs(2858) <= b;
    layer0_outputs(2859) <= not b;
    layer0_outputs(2860) <= not (a or b);
    layer0_outputs(2861) <= b;
    layer0_outputs(2862) <= not (a or b);
    layer0_outputs(2863) <= not b;
    layer0_outputs(2864) <= a and not b;
    layer0_outputs(2865) <= a xor b;
    layer0_outputs(2866) <= not a;
    layer0_outputs(2867) <= b;
    layer0_outputs(2868) <= a or b;
    layer0_outputs(2869) <= a;
    layer0_outputs(2870) <= a and b;
    layer0_outputs(2871) <= a xor b;
    layer0_outputs(2872) <= a or b;
    layer0_outputs(2873) <= a and not b;
    layer0_outputs(2874) <= not a or b;
    layer0_outputs(2875) <= not b or a;
    layer0_outputs(2876) <= a xor b;
    layer0_outputs(2877) <= 1'b1;
    layer0_outputs(2878) <= not (a or b);
    layer0_outputs(2879) <= not b or a;
    layer0_outputs(2880) <= not (a or b);
    layer0_outputs(2881) <= a;
    layer0_outputs(2882) <= not a or b;
    layer0_outputs(2883) <= a and b;
    layer0_outputs(2884) <= a;
    layer0_outputs(2885) <= a or b;
    layer0_outputs(2886) <= not b;
    layer0_outputs(2887) <= a xor b;
    layer0_outputs(2888) <= not b;
    layer0_outputs(2889) <= b;
    layer0_outputs(2890) <= a and not b;
    layer0_outputs(2891) <= not (a or b);
    layer0_outputs(2892) <= not (a or b);
    layer0_outputs(2893) <= a;
    layer0_outputs(2894) <= b and not a;
    layer0_outputs(2895) <= not (a xor b);
    layer0_outputs(2896) <= not a or b;
    layer0_outputs(2897) <= b and not a;
    layer0_outputs(2898) <= b and not a;
    layer0_outputs(2899) <= not a or b;
    layer0_outputs(2900) <= not a;
    layer0_outputs(2901) <= not (a or b);
    layer0_outputs(2902) <= not b;
    layer0_outputs(2903) <= not (a xor b);
    layer0_outputs(2904) <= a or b;
    layer0_outputs(2905) <= not (a xor b);
    layer0_outputs(2906) <= not a;
    layer0_outputs(2907) <= 1'b0;
    layer0_outputs(2908) <= not a or b;
    layer0_outputs(2909) <= not b;
    layer0_outputs(2910) <= a and not b;
    layer0_outputs(2911) <= a;
    layer0_outputs(2912) <= a xor b;
    layer0_outputs(2913) <= b;
    layer0_outputs(2914) <= b and not a;
    layer0_outputs(2915) <= b;
    layer0_outputs(2916) <= not (a or b);
    layer0_outputs(2917) <= a or b;
    layer0_outputs(2918) <= a or b;
    layer0_outputs(2919) <= not a or b;
    layer0_outputs(2920) <= a or b;
    layer0_outputs(2921) <= not a or b;
    layer0_outputs(2922) <= not a or b;
    layer0_outputs(2923) <= a or b;
    layer0_outputs(2924) <= a;
    layer0_outputs(2925) <= not (a or b);
    layer0_outputs(2926) <= a or b;
    layer0_outputs(2927) <= a and not b;
    layer0_outputs(2928) <= a and not b;
    layer0_outputs(2929) <= 1'b0;
    layer0_outputs(2930) <= a and b;
    layer0_outputs(2931) <= not (a xor b);
    layer0_outputs(2932) <= not b;
    layer0_outputs(2933) <= a and not b;
    layer0_outputs(2934) <= not (a or b);
    layer0_outputs(2935) <= not a;
    layer0_outputs(2936) <= not b or a;
    layer0_outputs(2937) <= not b;
    layer0_outputs(2938) <= not (a and b);
    layer0_outputs(2939) <= b and not a;
    layer0_outputs(2940) <= b and not a;
    layer0_outputs(2941) <= a and b;
    layer0_outputs(2942) <= not (a or b);
    layer0_outputs(2943) <= not b or a;
    layer0_outputs(2944) <= not a or b;
    layer0_outputs(2945) <= a and not b;
    layer0_outputs(2946) <= a or b;
    layer0_outputs(2947) <= b and not a;
    layer0_outputs(2948) <= b;
    layer0_outputs(2949) <= not (a and b);
    layer0_outputs(2950) <= not (a and b);
    layer0_outputs(2951) <= b;
    layer0_outputs(2952) <= not (a or b);
    layer0_outputs(2953) <= a and not b;
    layer0_outputs(2954) <= b and not a;
    layer0_outputs(2955) <= not (a or b);
    layer0_outputs(2956) <= not (a xor b);
    layer0_outputs(2957) <= not b or a;
    layer0_outputs(2958) <= b and not a;
    layer0_outputs(2959) <= a and not b;
    layer0_outputs(2960) <= b;
    layer0_outputs(2961) <= not b or a;
    layer0_outputs(2962) <= not b;
    layer0_outputs(2963) <= b;
    layer0_outputs(2964) <= a and not b;
    layer0_outputs(2965) <= not (a xor b);
    layer0_outputs(2966) <= a and not b;
    layer0_outputs(2967) <= a;
    layer0_outputs(2968) <= not (a and b);
    layer0_outputs(2969) <= not (a xor b);
    layer0_outputs(2970) <= a xor b;
    layer0_outputs(2971) <= 1'b0;
    layer0_outputs(2972) <= a xor b;
    layer0_outputs(2973) <= not (a or b);
    layer0_outputs(2974) <= not b;
    layer0_outputs(2975) <= not a;
    layer0_outputs(2976) <= not a;
    layer0_outputs(2977) <= not a or b;
    layer0_outputs(2978) <= not a;
    layer0_outputs(2979) <= a or b;
    layer0_outputs(2980) <= not (a and b);
    layer0_outputs(2981) <= a or b;
    layer0_outputs(2982) <= not (a and b);
    layer0_outputs(2983) <= not a or b;
    layer0_outputs(2984) <= a;
    layer0_outputs(2985) <= not (a or b);
    layer0_outputs(2986) <= 1'b0;
    layer0_outputs(2987) <= not (a or b);
    layer0_outputs(2988) <= not (a or b);
    layer0_outputs(2989) <= a xor b;
    layer0_outputs(2990) <= not (a xor b);
    layer0_outputs(2991) <= not a;
    layer0_outputs(2992) <= not a;
    layer0_outputs(2993) <= 1'b0;
    layer0_outputs(2994) <= not a;
    layer0_outputs(2995) <= a xor b;
    layer0_outputs(2996) <= b and not a;
    layer0_outputs(2997) <= 1'b1;
    layer0_outputs(2998) <= not b;
    layer0_outputs(2999) <= a or b;
    layer0_outputs(3000) <= not a or b;
    layer0_outputs(3001) <= a xor b;
    layer0_outputs(3002) <= a or b;
    layer0_outputs(3003) <= not b;
    layer0_outputs(3004) <= b and not a;
    layer0_outputs(3005) <= 1'b0;
    layer0_outputs(3006) <= b and not a;
    layer0_outputs(3007) <= a;
    layer0_outputs(3008) <= not (a and b);
    layer0_outputs(3009) <= not (a xor b);
    layer0_outputs(3010) <= not b or a;
    layer0_outputs(3011) <= 1'b1;
    layer0_outputs(3012) <= a or b;
    layer0_outputs(3013) <= a or b;
    layer0_outputs(3014) <= a or b;
    layer0_outputs(3015) <= a xor b;
    layer0_outputs(3016) <= a and b;
    layer0_outputs(3017) <= a;
    layer0_outputs(3018) <= a or b;
    layer0_outputs(3019) <= a or b;
    layer0_outputs(3020) <= a or b;
    layer0_outputs(3021) <= a or b;
    layer0_outputs(3022) <= a xor b;
    layer0_outputs(3023) <= not a;
    layer0_outputs(3024) <= not b;
    layer0_outputs(3025) <= b and not a;
    layer0_outputs(3026) <= not a;
    layer0_outputs(3027) <= not b or a;
    layer0_outputs(3028) <= a;
    layer0_outputs(3029) <= not (a and b);
    layer0_outputs(3030) <= b;
    layer0_outputs(3031) <= not (a and b);
    layer0_outputs(3032) <= not (a or b);
    layer0_outputs(3033) <= b and not a;
    layer0_outputs(3034) <= not (a xor b);
    layer0_outputs(3035) <= a;
    layer0_outputs(3036) <= not b;
    layer0_outputs(3037) <= a or b;
    layer0_outputs(3038) <= not (a and b);
    layer0_outputs(3039) <= a and b;
    layer0_outputs(3040) <= not (a xor b);
    layer0_outputs(3041) <= a and not b;
    layer0_outputs(3042) <= a xor b;
    layer0_outputs(3043) <= not (a xor b);
    layer0_outputs(3044) <= not b;
    layer0_outputs(3045) <= 1'b1;
    layer0_outputs(3046) <= a or b;
    layer0_outputs(3047) <= not b;
    layer0_outputs(3048) <= a xor b;
    layer0_outputs(3049) <= not (a xor b);
    layer0_outputs(3050) <= 1'b1;
    layer0_outputs(3051) <= 1'b1;
    layer0_outputs(3052) <= a xor b;
    layer0_outputs(3053) <= a and not b;
    layer0_outputs(3054) <= a or b;
    layer0_outputs(3055) <= not b;
    layer0_outputs(3056) <= b and not a;
    layer0_outputs(3057) <= 1'b0;
    layer0_outputs(3058) <= not (a or b);
    layer0_outputs(3059) <= a xor b;
    layer0_outputs(3060) <= a or b;
    layer0_outputs(3061) <= a;
    layer0_outputs(3062) <= b and not a;
    layer0_outputs(3063) <= b;
    layer0_outputs(3064) <= not b;
    layer0_outputs(3065) <= not a;
    layer0_outputs(3066) <= a;
    layer0_outputs(3067) <= not b or a;
    layer0_outputs(3068) <= b;
    layer0_outputs(3069) <= not a or b;
    layer0_outputs(3070) <= not (a and b);
    layer0_outputs(3071) <= 1'b0;
    layer0_outputs(3072) <= a xor b;
    layer0_outputs(3073) <= a or b;
    layer0_outputs(3074) <= not b;
    layer0_outputs(3075) <= b and not a;
    layer0_outputs(3076) <= a;
    layer0_outputs(3077) <= a and not b;
    layer0_outputs(3078) <= b;
    layer0_outputs(3079) <= not (a xor b);
    layer0_outputs(3080) <= not (a or b);
    layer0_outputs(3081) <= a and not b;
    layer0_outputs(3082) <= not (a and b);
    layer0_outputs(3083) <= a or b;
    layer0_outputs(3084) <= not a or b;
    layer0_outputs(3085) <= a and not b;
    layer0_outputs(3086) <= a and not b;
    layer0_outputs(3087) <= a or b;
    layer0_outputs(3088) <= a and b;
    layer0_outputs(3089) <= not a;
    layer0_outputs(3090) <= a or b;
    layer0_outputs(3091) <= a or b;
    layer0_outputs(3092) <= a and not b;
    layer0_outputs(3093) <= a;
    layer0_outputs(3094) <= not a;
    layer0_outputs(3095) <= a;
    layer0_outputs(3096) <= b;
    layer0_outputs(3097) <= not (a or b);
    layer0_outputs(3098) <= a or b;
    layer0_outputs(3099) <= not (a or b);
    layer0_outputs(3100) <= a xor b;
    layer0_outputs(3101) <= not a;
    layer0_outputs(3102) <= not (a or b);
    layer0_outputs(3103) <= not b or a;
    layer0_outputs(3104) <= not (a xor b);
    layer0_outputs(3105) <= a xor b;
    layer0_outputs(3106) <= 1'b1;
    layer0_outputs(3107) <= a or b;
    layer0_outputs(3108) <= not (a or b);
    layer0_outputs(3109) <= a and not b;
    layer0_outputs(3110) <= not b;
    layer0_outputs(3111) <= b;
    layer0_outputs(3112) <= b;
    layer0_outputs(3113) <= b and not a;
    layer0_outputs(3114) <= a and not b;
    layer0_outputs(3115) <= not (a xor b);
    layer0_outputs(3116) <= a and not b;
    layer0_outputs(3117) <= a xor b;
    layer0_outputs(3118) <= a and not b;
    layer0_outputs(3119) <= a or b;
    layer0_outputs(3120) <= a and not b;
    layer0_outputs(3121) <= not (a or b);
    layer0_outputs(3122) <= not b;
    layer0_outputs(3123) <= not (a or b);
    layer0_outputs(3124) <= 1'b0;
    layer0_outputs(3125) <= a and not b;
    layer0_outputs(3126) <= b and not a;
    layer0_outputs(3127) <= a and not b;
    layer0_outputs(3128) <= not b or a;
    layer0_outputs(3129) <= a;
    layer0_outputs(3130) <= a and not b;
    layer0_outputs(3131) <= not b or a;
    layer0_outputs(3132) <= a xor b;
    layer0_outputs(3133) <= not (a or b);
    layer0_outputs(3134) <= a xor b;
    layer0_outputs(3135) <= b and not a;
    layer0_outputs(3136) <= 1'b0;
    layer0_outputs(3137) <= 1'b0;
    layer0_outputs(3138) <= a or b;
    layer0_outputs(3139) <= not a or b;
    layer0_outputs(3140) <= not (a or b);
    layer0_outputs(3141) <= not (a or b);
    layer0_outputs(3142) <= a or b;
    layer0_outputs(3143) <= a and b;
    layer0_outputs(3144) <= b;
    layer0_outputs(3145) <= not (a or b);
    layer0_outputs(3146) <= not b or a;
    layer0_outputs(3147) <= b;
    layer0_outputs(3148) <= a and not b;
    layer0_outputs(3149) <= a;
    layer0_outputs(3150) <= not b;
    layer0_outputs(3151) <= not b;
    layer0_outputs(3152) <= b and not a;
    layer0_outputs(3153) <= a and b;
    layer0_outputs(3154) <= a or b;
    layer0_outputs(3155) <= not a;
    layer0_outputs(3156) <= b;
    layer0_outputs(3157) <= not (a or b);
    layer0_outputs(3158) <= b and not a;
    layer0_outputs(3159) <= a or b;
    layer0_outputs(3160) <= a or b;
    layer0_outputs(3161) <= b;
    layer0_outputs(3162) <= a or b;
    layer0_outputs(3163) <= not a or b;
    layer0_outputs(3164) <= not b;
    layer0_outputs(3165) <= b and not a;
    layer0_outputs(3166) <= not (a or b);
    layer0_outputs(3167) <= b and not a;
    layer0_outputs(3168) <= not b;
    layer0_outputs(3169) <= not a;
    layer0_outputs(3170) <= not a;
    layer0_outputs(3171) <= b and not a;
    layer0_outputs(3172) <= a xor b;
    layer0_outputs(3173) <= a and not b;
    layer0_outputs(3174) <= a;
    layer0_outputs(3175) <= not a;
    layer0_outputs(3176) <= not (a and b);
    layer0_outputs(3177) <= a and not b;
    layer0_outputs(3178) <= not a or b;
    layer0_outputs(3179) <= a or b;
    layer0_outputs(3180) <= not b;
    layer0_outputs(3181) <= a and not b;
    layer0_outputs(3182) <= not (a or b);
    layer0_outputs(3183) <= a or b;
    layer0_outputs(3184) <= not (a xor b);
    layer0_outputs(3185) <= not a;
    layer0_outputs(3186) <= not (a or b);
    layer0_outputs(3187) <= a or b;
    layer0_outputs(3188) <= not (a or b);
    layer0_outputs(3189) <= a or b;
    layer0_outputs(3190) <= a xor b;
    layer0_outputs(3191) <= not b or a;
    layer0_outputs(3192) <= not (a or b);
    layer0_outputs(3193) <= a xor b;
    layer0_outputs(3194) <= not b;
    layer0_outputs(3195) <= a and not b;
    layer0_outputs(3196) <= a or b;
    layer0_outputs(3197) <= not (a or b);
    layer0_outputs(3198) <= not (a or b);
    layer0_outputs(3199) <= a or b;
    layer0_outputs(3200) <= not b;
    layer0_outputs(3201) <= not a or b;
    layer0_outputs(3202) <= not b;
    layer0_outputs(3203) <= not (a or b);
    layer0_outputs(3204) <= 1'b0;
    layer0_outputs(3205) <= not (a xor b);
    layer0_outputs(3206) <= a or b;
    layer0_outputs(3207) <= a or b;
    layer0_outputs(3208) <= a or b;
    layer0_outputs(3209) <= not b or a;
    layer0_outputs(3210) <= not a or b;
    layer0_outputs(3211) <= not b;
    layer0_outputs(3212) <= not b or a;
    layer0_outputs(3213) <= not (a or b);
    layer0_outputs(3214) <= a and not b;
    layer0_outputs(3215) <= a and not b;
    layer0_outputs(3216) <= not a or b;
    layer0_outputs(3217) <= not (a or b);
    layer0_outputs(3218) <= not a or b;
    layer0_outputs(3219) <= b;
    layer0_outputs(3220) <= a or b;
    layer0_outputs(3221) <= not b;
    layer0_outputs(3222) <= not (a or b);
    layer0_outputs(3223) <= b;
    layer0_outputs(3224) <= not (a or b);
    layer0_outputs(3225) <= a xor b;
    layer0_outputs(3226) <= a or b;
    layer0_outputs(3227) <= a or b;
    layer0_outputs(3228) <= a or b;
    layer0_outputs(3229) <= a and not b;
    layer0_outputs(3230) <= 1'b1;
    layer0_outputs(3231) <= not (a xor b);
    layer0_outputs(3232) <= a xor b;
    layer0_outputs(3233) <= a or b;
    layer0_outputs(3234) <= not b;
    layer0_outputs(3235) <= b;
    layer0_outputs(3236) <= not (a or b);
    layer0_outputs(3237) <= b and not a;
    layer0_outputs(3238) <= not a or b;
    layer0_outputs(3239) <= not (a and b);
    layer0_outputs(3240) <= a xor b;
    layer0_outputs(3241) <= a;
    layer0_outputs(3242) <= not a;
    layer0_outputs(3243) <= a or b;
    layer0_outputs(3244) <= not b;
    layer0_outputs(3245) <= a or b;
    layer0_outputs(3246) <= 1'b0;
    layer0_outputs(3247) <= not b or a;
    layer0_outputs(3248) <= b;
    layer0_outputs(3249) <= a;
    layer0_outputs(3250) <= b;
    layer0_outputs(3251) <= 1'b1;
    layer0_outputs(3252) <= not (a xor b);
    layer0_outputs(3253) <= not (a or b);
    layer0_outputs(3254) <= not (a or b);
    layer0_outputs(3255) <= a or b;
    layer0_outputs(3256) <= not a;
    layer0_outputs(3257) <= a and not b;
    layer0_outputs(3258) <= 1'b1;
    layer0_outputs(3259) <= 1'b1;
    layer0_outputs(3260) <= not a or b;
    layer0_outputs(3261) <= not a or b;
    layer0_outputs(3262) <= not (a and b);
    layer0_outputs(3263) <= a;
    layer0_outputs(3264) <= not b or a;
    layer0_outputs(3265) <= not (a xor b);
    layer0_outputs(3266) <= not (a or b);
    layer0_outputs(3267) <= a and not b;
    layer0_outputs(3268) <= a;
    layer0_outputs(3269) <= a xor b;
    layer0_outputs(3270) <= a or b;
    layer0_outputs(3271) <= a or b;
    layer0_outputs(3272) <= not (a or b);
    layer0_outputs(3273) <= a and not b;
    layer0_outputs(3274) <= 1'b1;
    layer0_outputs(3275) <= not (a or b);
    layer0_outputs(3276) <= not a;
    layer0_outputs(3277) <= not a;
    layer0_outputs(3278) <= not b;
    layer0_outputs(3279) <= not a or b;
    layer0_outputs(3280) <= not (a xor b);
    layer0_outputs(3281) <= b;
    layer0_outputs(3282) <= b;
    layer0_outputs(3283) <= a and not b;
    layer0_outputs(3284) <= a xor b;
    layer0_outputs(3285) <= not (a and b);
    layer0_outputs(3286) <= a and not b;
    layer0_outputs(3287) <= not b;
    layer0_outputs(3288) <= a or b;
    layer0_outputs(3289) <= 1'b0;
    layer0_outputs(3290) <= b and not a;
    layer0_outputs(3291) <= not (a or b);
    layer0_outputs(3292) <= b and not a;
    layer0_outputs(3293) <= not (a or b);
    layer0_outputs(3294) <= b and not a;
    layer0_outputs(3295) <= not (a xor b);
    layer0_outputs(3296) <= a and b;
    layer0_outputs(3297) <= not (a or b);
    layer0_outputs(3298) <= not a;
    layer0_outputs(3299) <= not b or a;
    layer0_outputs(3300) <= b;
    layer0_outputs(3301) <= a or b;
    layer0_outputs(3302) <= b;
    layer0_outputs(3303) <= not b or a;
    layer0_outputs(3304) <= not a or b;
    layer0_outputs(3305) <= a or b;
    layer0_outputs(3306) <= not (a or b);
    layer0_outputs(3307) <= b;
    layer0_outputs(3308) <= 1'b1;
    layer0_outputs(3309) <= not a;
    layer0_outputs(3310) <= not a or b;
    layer0_outputs(3311) <= not (a and b);
    layer0_outputs(3312) <= 1'b1;
    layer0_outputs(3313) <= not (a or b);
    layer0_outputs(3314) <= not b or a;
    layer0_outputs(3315) <= b;
    layer0_outputs(3316) <= not a;
    layer0_outputs(3317) <= not a;
    layer0_outputs(3318) <= not (a xor b);
    layer0_outputs(3319) <= not (a xor b);
    layer0_outputs(3320) <= a or b;
    layer0_outputs(3321) <= not (a or b);
    layer0_outputs(3322) <= not a or b;
    layer0_outputs(3323) <= not a;
    layer0_outputs(3324) <= b;
    layer0_outputs(3325) <= b;
    layer0_outputs(3326) <= a;
    layer0_outputs(3327) <= not a;
    layer0_outputs(3328) <= a;
    layer0_outputs(3329) <= not (a xor b);
    layer0_outputs(3330) <= a;
    layer0_outputs(3331) <= b and not a;
    layer0_outputs(3332) <= b and not a;
    layer0_outputs(3333) <= not (a xor b);
    layer0_outputs(3334) <= a;
    layer0_outputs(3335) <= not (a and b);
    layer0_outputs(3336) <= not a;
    layer0_outputs(3337) <= a and not b;
    layer0_outputs(3338) <= not (a or b);
    layer0_outputs(3339) <= not (a and b);
    layer0_outputs(3340) <= a or b;
    layer0_outputs(3341) <= not (a and b);
    layer0_outputs(3342) <= b and not a;
    layer0_outputs(3343) <= a or b;
    layer0_outputs(3344) <= not b or a;
    layer0_outputs(3345) <= not a;
    layer0_outputs(3346) <= a and not b;
    layer0_outputs(3347) <= not a or b;
    layer0_outputs(3348) <= a and not b;
    layer0_outputs(3349) <= a;
    layer0_outputs(3350) <= not a;
    layer0_outputs(3351) <= b;
    layer0_outputs(3352) <= a;
    layer0_outputs(3353) <= not (a or b);
    layer0_outputs(3354) <= 1'b0;
    layer0_outputs(3355) <= not (a and b);
    layer0_outputs(3356) <= a or b;
    layer0_outputs(3357) <= not (a or b);
    layer0_outputs(3358) <= not b or a;
    layer0_outputs(3359) <= not b;
    layer0_outputs(3360) <= not a or b;
    layer0_outputs(3361) <= not (a xor b);
    layer0_outputs(3362) <= a;
    layer0_outputs(3363) <= a and not b;
    layer0_outputs(3364) <= a or b;
    layer0_outputs(3365) <= b and not a;
    layer0_outputs(3366) <= 1'b1;
    layer0_outputs(3367) <= b and not a;
    layer0_outputs(3368) <= a and not b;
    layer0_outputs(3369) <= not a or b;
    layer0_outputs(3370) <= not (a or b);
    layer0_outputs(3371) <= 1'b1;
    layer0_outputs(3372) <= not b;
    layer0_outputs(3373) <= not (a or b);
    layer0_outputs(3374) <= not a or b;
    layer0_outputs(3375) <= not (a xor b);
    layer0_outputs(3376) <= b and not a;
    layer0_outputs(3377) <= a;
    layer0_outputs(3378) <= not (a or b);
    layer0_outputs(3379) <= not (a xor b);
    layer0_outputs(3380) <= not b;
    layer0_outputs(3381) <= a and b;
    layer0_outputs(3382) <= not a or b;
    layer0_outputs(3383) <= a or b;
    layer0_outputs(3384) <= a and not b;
    layer0_outputs(3385) <= a and b;
    layer0_outputs(3386) <= not b or a;
    layer0_outputs(3387) <= b and not a;
    layer0_outputs(3388) <= not (a or b);
    layer0_outputs(3389) <= not a or b;
    layer0_outputs(3390) <= not a;
    layer0_outputs(3391) <= b;
    layer0_outputs(3392) <= not (a or b);
    layer0_outputs(3393) <= not (a or b);
    layer0_outputs(3394) <= not (a xor b);
    layer0_outputs(3395) <= b and not a;
    layer0_outputs(3396) <= b;
    layer0_outputs(3397) <= not a or b;
    layer0_outputs(3398) <= not b;
    layer0_outputs(3399) <= not (a xor b);
    layer0_outputs(3400) <= not (a or b);
    layer0_outputs(3401) <= 1'b0;
    layer0_outputs(3402) <= b;
    layer0_outputs(3403) <= a;
    layer0_outputs(3404) <= a or b;
    layer0_outputs(3405) <= not (a or b);
    layer0_outputs(3406) <= a;
    layer0_outputs(3407) <= b;
    layer0_outputs(3408) <= not (a and b);
    layer0_outputs(3409) <= 1'b1;
    layer0_outputs(3410) <= not (a xor b);
    layer0_outputs(3411) <= not (a or b);
    layer0_outputs(3412) <= a or b;
    layer0_outputs(3413) <= not (a or b);
    layer0_outputs(3414) <= a xor b;
    layer0_outputs(3415) <= b and not a;
    layer0_outputs(3416) <= a;
    layer0_outputs(3417) <= a xor b;
    layer0_outputs(3418) <= b;
    layer0_outputs(3419) <= not b;
    layer0_outputs(3420) <= not (a xor b);
    layer0_outputs(3421) <= not b;
    layer0_outputs(3422) <= b;
    layer0_outputs(3423) <= not (a or b);
    layer0_outputs(3424) <= a or b;
    layer0_outputs(3425) <= a;
    layer0_outputs(3426) <= not a;
    layer0_outputs(3427) <= b;
    layer0_outputs(3428) <= not (a xor b);
    layer0_outputs(3429) <= 1'b0;
    layer0_outputs(3430) <= a or b;
    layer0_outputs(3431) <= 1'b0;
    layer0_outputs(3432) <= 1'b0;
    layer0_outputs(3433) <= b and not a;
    layer0_outputs(3434) <= not b;
    layer0_outputs(3435) <= a or b;
    layer0_outputs(3436) <= not b;
    layer0_outputs(3437) <= not a;
    layer0_outputs(3438) <= not (a or b);
    layer0_outputs(3439) <= not a or b;
    layer0_outputs(3440) <= not (a xor b);
    layer0_outputs(3441) <= a or b;
    layer0_outputs(3442) <= not (a or b);
    layer0_outputs(3443) <= not b or a;
    layer0_outputs(3444) <= not b;
    layer0_outputs(3445) <= not (a xor b);
    layer0_outputs(3446) <= not b;
    layer0_outputs(3447) <= not b or a;
    layer0_outputs(3448) <= a and not b;
    layer0_outputs(3449) <= a or b;
    layer0_outputs(3450) <= not (a xor b);
    layer0_outputs(3451) <= not b or a;
    layer0_outputs(3452) <= a xor b;
    layer0_outputs(3453) <= 1'b0;
    layer0_outputs(3454) <= a;
    layer0_outputs(3455) <= not a or b;
    layer0_outputs(3456) <= b;
    layer0_outputs(3457) <= a or b;
    layer0_outputs(3458) <= not b or a;
    layer0_outputs(3459) <= b;
    layer0_outputs(3460) <= a;
    layer0_outputs(3461) <= not (a or b);
    layer0_outputs(3462) <= a;
    layer0_outputs(3463) <= not a;
    layer0_outputs(3464) <= not (a and b);
    layer0_outputs(3465) <= not a;
    layer0_outputs(3466) <= a and not b;
    layer0_outputs(3467) <= not (a xor b);
    layer0_outputs(3468) <= not (a xor b);
    layer0_outputs(3469) <= a and not b;
    layer0_outputs(3470) <= not b;
    layer0_outputs(3471) <= a xor b;
    layer0_outputs(3472) <= a and not b;
    layer0_outputs(3473) <= a and not b;
    layer0_outputs(3474) <= a or b;
    layer0_outputs(3475) <= a or b;
    layer0_outputs(3476) <= b;
    layer0_outputs(3477) <= b and not a;
    layer0_outputs(3478) <= not (a xor b);
    layer0_outputs(3479) <= b;
    layer0_outputs(3480) <= not b;
    layer0_outputs(3481) <= 1'b1;
    layer0_outputs(3482) <= not a;
    layer0_outputs(3483) <= a and b;
    layer0_outputs(3484) <= b and not a;
    layer0_outputs(3485) <= not a;
    layer0_outputs(3486) <= a xor b;
    layer0_outputs(3487) <= a xor b;
    layer0_outputs(3488) <= not (a and b);
    layer0_outputs(3489) <= not b;
    layer0_outputs(3490) <= not b;
    layer0_outputs(3491) <= not a or b;
    layer0_outputs(3492) <= a and not b;
    layer0_outputs(3493) <= a or b;
    layer0_outputs(3494) <= a;
    layer0_outputs(3495) <= b;
    layer0_outputs(3496) <= not a or b;
    layer0_outputs(3497) <= b and not a;
    layer0_outputs(3498) <= a or b;
    layer0_outputs(3499) <= a or b;
    layer0_outputs(3500) <= a or b;
    layer0_outputs(3501) <= not (a xor b);
    layer0_outputs(3502) <= b;
    layer0_outputs(3503) <= not b;
    layer0_outputs(3504) <= a;
    layer0_outputs(3505) <= not b;
    layer0_outputs(3506) <= a or b;
    layer0_outputs(3507) <= not a;
    layer0_outputs(3508) <= b;
    layer0_outputs(3509) <= a and b;
    layer0_outputs(3510) <= a or b;
    layer0_outputs(3511) <= not (a or b);
    layer0_outputs(3512) <= not (a or b);
    layer0_outputs(3513) <= a;
    layer0_outputs(3514) <= not (a or b);
    layer0_outputs(3515) <= not (a or b);
    layer0_outputs(3516) <= 1'b0;
    layer0_outputs(3517) <= not (a or b);
    layer0_outputs(3518) <= not (a xor b);
    layer0_outputs(3519) <= b and not a;
    layer0_outputs(3520) <= b and not a;
    layer0_outputs(3521) <= not b;
    layer0_outputs(3522) <= b and not a;
    layer0_outputs(3523) <= a xor b;
    layer0_outputs(3524) <= b;
    layer0_outputs(3525) <= not (a or b);
    layer0_outputs(3526) <= a or b;
    layer0_outputs(3527) <= not a or b;
    layer0_outputs(3528) <= not (a or b);
    layer0_outputs(3529) <= not b;
    layer0_outputs(3530) <= a xor b;
    layer0_outputs(3531) <= not b or a;
    layer0_outputs(3532) <= not (a or b);
    layer0_outputs(3533) <= b and not a;
    layer0_outputs(3534) <= not (a or b);
    layer0_outputs(3535) <= b;
    layer0_outputs(3536) <= not (a or b);
    layer0_outputs(3537) <= not a;
    layer0_outputs(3538) <= b;
    layer0_outputs(3539) <= not (a xor b);
    layer0_outputs(3540) <= a xor b;
    layer0_outputs(3541) <= not (a xor b);
    layer0_outputs(3542) <= a and not b;
    layer0_outputs(3543) <= not a;
    layer0_outputs(3544) <= not (a or b);
    layer0_outputs(3545) <= not (a or b);
    layer0_outputs(3546) <= not b or a;
    layer0_outputs(3547) <= a xor b;
    layer0_outputs(3548) <= not (a xor b);
    layer0_outputs(3549) <= 1'b0;
    layer0_outputs(3550) <= not (a and b);
    layer0_outputs(3551) <= not b or a;
    layer0_outputs(3552) <= not (a xor b);
    layer0_outputs(3553) <= b and not a;
    layer0_outputs(3554) <= a or b;
    layer0_outputs(3555) <= a;
    layer0_outputs(3556) <= b and not a;
    layer0_outputs(3557) <= a and not b;
    layer0_outputs(3558) <= 1'b1;
    layer0_outputs(3559) <= b;
    layer0_outputs(3560) <= a or b;
    layer0_outputs(3561) <= not a;
    layer0_outputs(3562) <= not (a xor b);
    layer0_outputs(3563) <= not (a or b);
    layer0_outputs(3564) <= not a;
    layer0_outputs(3565) <= a and b;
    layer0_outputs(3566) <= not (a or b);
    layer0_outputs(3567) <= b and not a;
    layer0_outputs(3568) <= not (a xor b);
    layer0_outputs(3569) <= a;
    layer0_outputs(3570) <= not (a xor b);
    layer0_outputs(3571) <= not (a xor b);
    layer0_outputs(3572) <= not a or b;
    layer0_outputs(3573) <= not a or b;
    layer0_outputs(3574) <= 1'b1;
    layer0_outputs(3575) <= not (a or b);
    layer0_outputs(3576) <= b and not a;
    layer0_outputs(3577) <= a xor b;
    layer0_outputs(3578) <= not a or b;
    layer0_outputs(3579) <= a and not b;
    layer0_outputs(3580) <= 1'b1;
    layer0_outputs(3581) <= a;
    layer0_outputs(3582) <= a xor b;
    layer0_outputs(3583) <= b;
    layer0_outputs(3584) <= b and not a;
    layer0_outputs(3585) <= a or b;
    layer0_outputs(3586) <= not (a or b);
    layer0_outputs(3587) <= a and not b;
    layer0_outputs(3588) <= a;
    layer0_outputs(3589) <= not b;
    layer0_outputs(3590) <= a or b;
    layer0_outputs(3591) <= not b;
    layer0_outputs(3592) <= not (a xor b);
    layer0_outputs(3593) <= b and not a;
    layer0_outputs(3594) <= not a or b;
    layer0_outputs(3595) <= not (a or b);
    layer0_outputs(3596) <= not (a or b);
    layer0_outputs(3597) <= not (a or b);
    layer0_outputs(3598) <= a or b;
    layer0_outputs(3599) <= not b;
    layer0_outputs(3600) <= b and not a;
    layer0_outputs(3601) <= not (a xor b);
    layer0_outputs(3602) <= not (a xor b);
    layer0_outputs(3603) <= 1'b1;
    layer0_outputs(3604) <= not (a xor b);
    layer0_outputs(3605) <= a and not b;
    layer0_outputs(3606) <= not a or b;
    layer0_outputs(3607) <= not a or b;
    layer0_outputs(3608) <= b;
    layer0_outputs(3609) <= a xor b;
    layer0_outputs(3610) <= a or b;
    layer0_outputs(3611) <= a and not b;
    layer0_outputs(3612) <= b;
    layer0_outputs(3613) <= not b;
    layer0_outputs(3614) <= a or b;
    layer0_outputs(3615) <= a xor b;
    layer0_outputs(3616) <= not (a or b);
    layer0_outputs(3617) <= a;
    layer0_outputs(3618) <= a and not b;
    layer0_outputs(3619) <= a and not b;
    layer0_outputs(3620) <= 1'b1;
    layer0_outputs(3621) <= not (a and b);
    layer0_outputs(3622) <= b;
    layer0_outputs(3623) <= a;
    layer0_outputs(3624) <= not (a or b);
    layer0_outputs(3625) <= a;
    layer0_outputs(3626) <= b and not a;
    layer0_outputs(3627) <= a xor b;
    layer0_outputs(3628) <= a and not b;
    layer0_outputs(3629) <= a and b;
    layer0_outputs(3630) <= a;
    layer0_outputs(3631) <= not (a xor b);
    layer0_outputs(3632) <= a or b;
    layer0_outputs(3633) <= a;
    layer0_outputs(3634) <= not (a xor b);
    layer0_outputs(3635) <= not b;
    layer0_outputs(3636) <= not (a or b);
    layer0_outputs(3637) <= b;
    layer0_outputs(3638) <= b;
    layer0_outputs(3639) <= a and not b;
    layer0_outputs(3640) <= a xor b;
    layer0_outputs(3641) <= a and b;
    layer0_outputs(3642) <= a xor b;
    layer0_outputs(3643) <= a xor b;
    layer0_outputs(3644) <= not (a or b);
    layer0_outputs(3645) <= a xor b;
    layer0_outputs(3646) <= not b or a;
    layer0_outputs(3647) <= a or b;
    layer0_outputs(3648) <= not b or a;
    layer0_outputs(3649) <= not a;
    layer0_outputs(3650) <= a or b;
    layer0_outputs(3651) <= not (a xor b);
    layer0_outputs(3652) <= not b or a;
    layer0_outputs(3653) <= a or b;
    layer0_outputs(3654) <= not a or b;
    layer0_outputs(3655) <= a;
    layer0_outputs(3656) <= b;
    layer0_outputs(3657) <= b;
    layer0_outputs(3658) <= not (a or b);
    layer0_outputs(3659) <= not b or a;
    layer0_outputs(3660) <= b and not a;
    layer0_outputs(3661) <= not (a xor b);
    layer0_outputs(3662) <= a;
    layer0_outputs(3663) <= a and not b;
    layer0_outputs(3664) <= not a;
    layer0_outputs(3665) <= not (a or b);
    layer0_outputs(3666) <= a or b;
    layer0_outputs(3667) <= not b or a;
    layer0_outputs(3668) <= a or b;
    layer0_outputs(3669) <= not a or b;
    layer0_outputs(3670) <= not a or b;
    layer0_outputs(3671) <= a or b;
    layer0_outputs(3672) <= a xor b;
    layer0_outputs(3673) <= a xor b;
    layer0_outputs(3674) <= not (a or b);
    layer0_outputs(3675) <= not b or a;
    layer0_outputs(3676) <= b and not a;
    layer0_outputs(3677) <= a;
    layer0_outputs(3678) <= not (a xor b);
    layer0_outputs(3679) <= 1'b1;
    layer0_outputs(3680) <= not a;
    layer0_outputs(3681) <= not b;
    layer0_outputs(3682) <= a and not b;
    layer0_outputs(3683) <= not b;
    layer0_outputs(3684) <= b;
    layer0_outputs(3685) <= a and not b;
    layer0_outputs(3686) <= not (a xor b);
    layer0_outputs(3687) <= not a;
    layer0_outputs(3688) <= not a or b;
    layer0_outputs(3689) <= a or b;
    layer0_outputs(3690) <= not b or a;
    layer0_outputs(3691) <= a and not b;
    layer0_outputs(3692) <= not (a or b);
    layer0_outputs(3693) <= b;
    layer0_outputs(3694) <= not (a and b);
    layer0_outputs(3695) <= b;
    layer0_outputs(3696) <= not (a xor b);
    layer0_outputs(3697) <= not b or a;
    layer0_outputs(3698) <= a xor b;
    layer0_outputs(3699) <= not (a or b);
    layer0_outputs(3700) <= a or b;
    layer0_outputs(3701) <= not b or a;
    layer0_outputs(3702) <= not (a or b);
    layer0_outputs(3703) <= a and not b;
    layer0_outputs(3704) <= a or b;
    layer0_outputs(3705) <= not a;
    layer0_outputs(3706) <= a or b;
    layer0_outputs(3707) <= a and not b;
    layer0_outputs(3708) <= a and b;
    layer0_outputs(3709) <= not (a or b);
    layer0_outputs(3710) <= not (a or b);
    layer0_outputs(3711) <= b and not a;
    layer0_outputs(3712) <= a and not b;
    layer0_outputs(3713) <= not (a xor b);
    layer0_outputs(3714) <= not (a or b);
    layer0_outputs(3715) <= not (a xor b);
    layer0_outputs(3716) <= not a;
    layer0_outputs(3717) <= b and not a;
    layer0_outputs(3718) <= a;
    layer0_outputs(3719) <= a;
    layer0_outputs(3720) <= a or b;
    layer0_outputs(3721) <= not a;
    layer0_outputs(3722) <= a xor b;
    layer0_outputs(3723) <= a;
    layer0_outputs(3724) <= a and not b;
    layer0_outputs(3725) <= a or b;
    layer0_outputs(3726) <= b;
    layer0_outputs(3727) <= 1'b0;
    layer0_outputs(3728) <= a and b;
    layer0_outputs(3729) <= not (a or b);
    layer0_outputs(3730) <= b and not a;
    layer0_outputs(3731) <= b;
    layer0_outputs(3732) <= not a;
    layer0_outputs(3733) <= not (a xor b);
    layer0_outputs(3734) <= a;
    layer0_outputs(3735) <= not (a or b);
    layer0_outputs(3736) <= not (a or b);
    layer0_outputs(3737) <= not (a and b);
    layer0_outputs(3738) <= not a;
    layer0_outputs(3739) <= not b or a;
    layer0_outputs(3740) <= not (a or b);
    layer0_outputs(3741) <= not (a or b);
    layer0_outputs(3742) <= 1'b1;
    layer0_outputs(3743) <= not (a or b);
    layer0_outputs(3744) <= not b;
    layer0_outputs(3745) <= not a or b;
    layer0_outputs(3746) <= a or b;
    layer0_outputs(3747) <= not (a xor b);
    layer0_outputs(3748) <= a or b;
    layer0_outputs(3749) <= a or b;
    layer0_outputs(3750) <= not a or b;
    layer0_outputs(3751) <= a or b;
    layer0_outputs(3752) <= a or b;
    layer0_outputs(3753) <= not b or a;
    layer0_outputs(3754) <= not (a or b);
    layer0_outputs(3755) <= not (a or b);
    layer0_outputs(3756) <= not (a xor b);
    layer0_outputs(3757) <= not a;
    layer0_outputs(3758) <= 1'b1;
    layer0_outputs(3759) <= not b;
    layer0_outputs(3760) <= not (a xor b);
    layer0_outputs(3761) <= not a;
    layer0_outputs(3762) <= a and b;
    layer0_outputs(3763) <= a xor b;
    layer0_outputs(3764) <= not a or b;
    layer0_outputs(3765) <= a and not b;
    layer0_outputs(3766) <= a xor b;
    layer0_outputs(3767) <= a or b;
    layer0_outputs(3768) <= b;
    layer0_outputs(3769) <= not b;
    layer0_outputs(3770) <= not a;
    layer0_outputs(3771) <= a or b;
    layer0_outputs(3772) <= 1'b0;
    layer0_outputs(3773) <= a and not b;
    layer0_outputs(3774) <= not (a xor b);
    layer0_outputs(3775) <= not a;
    layer0_outputs(3776) <= not b;
    layer0_outputs(3777) <= not (a or b);
    layer0_outputs(3778) <= not a;
    layer0_outputs(3779) <= a or b;
    layer0_outputs(3780) <= a or b;
    layer0_outputs(3781) <= a;
    layer0_outputs(3782) <= not a;
    layer0_outputs(3783) <= b and not a;
    layer0_outputs(3784) <= not a or b;
    layer0_outputs(3785) <= not b;
    layer0_outputs(3786) <= b and not a;
    layer0_outputs(3787) <= a;
    layer0_outputs(3788) <= b and not a;
    layer0_outputs(3789) <= not a;
    layer0_outputs(3790) <= not (a xor b);
    layer0_outputs(3791) <= a or b;
    layer0_outputs(3792) <= a;
    layer0_outputs(3793) <= b and not a;
    layer0_outputs(3794) <= not b or a;
    layer0_outputs(3795) <= a or b;
    layer0_outputs(3796) <= not b;
    layer0_outputs(3797) <= b and not a;
    layer0_outputs(3798) <= not b;
    layer0_outputs(3799) <= a xor b;
    layer0_outputs(3800) <= not (a xor b);
    layer0_outputs(3801) <= a or b;
    layer0_outputs(3802) <= a or b;
    layer0_outputs(3803) <= a and b;
    layer0_outputs(3804) <= not a;
    layer0_outputs(3805) <= not a;
    layer0_outputs(3806) <= 1'b1;
    layer0_outputs(3807) <= not (a xor b);
    layer0_outputs(3808) <= not b or a;
    layer0_outputs(3809) <= a or b;
    layer0_outputs(3810) <= not b;
    layer0_outputs(3811) <= a and b;
    layer0_outputs(3812) <= not b;
    layer0_outputs(3813) <= a;
    layer0_outputs(3814) <= a;
    layer0_outputs(3815) <= 1'b0;
    layer0_outputs(3816) <= not b;
    layer0_outputs(3817) <= a or b;
    layer0_outputs(3818) <= b and not a;
    layer0_outputs(3819) <= not (a or b);
    layer0_outputs(3820) <= b;
    layer0_outputs(3821) <= a and not b;
    layer0_outputs(3822) <= not b;
    layer0_outputs(3823) <= b and not a;
    layer0_outputs(3824) <= not b or a;
    layer0_outputs(3825) <= not b;
    layer0_outputs(3826) <= not (a or b);
    layer0_outputs(3827) <= a or b;
    layer0_outputs(3828) <= not a or b;
    layer0_outputs(3829) <= a xor b;
    layer0_outputs(3830) <= not (a or b);
    layer0_outputs(3831) <= a;
    layer0_outputs(3832) <= a xor b;
    layer0_outputs(3833) <= not b or a;
    layer0_outputs(3834) <= not b or a;
    layer0_outputs(3835) <= not a;
    layer0_outputs(3836) <= a;
    layer0_outputs(3837) <= a or b;
    layer0_outputs(3838) <= a or b;
    layer0_outputs(3839) <= a;
    layer0_outputs(3840) <= a or b;
    layer0_outputs(3841) <= a and not b;
    layer0_outputs(3842) <= not (a or b);
    layer0_outputs(3843) <= not a;
    layer0_outputs(3844) <= b and not a;
    layer0_outputs(3845) <= not a;
    layer0_outputs(3846) <= not (a and b);
    layer0_outputs(3847) <= not b;
    layer0_outputs(3848) <= not b;
    layer0_outputs(3849) <= not a;
    layer0_outputs(3850) <= not (a or b);
    layer0_outputs(3851) <= not (a xor b);
    layer0_outputs(3852) <= a and b;
    layer0_outputs(3853) <= a;
    layer0_outputs(3854) <= not (a xor b);
    layer0_outputs(3855) <= a or b;
    layer0_outputs(3856) <= not b;
    layer0_outputs(3857) <= b and not a;
    layer0_outputs(3858) <= 1'b0;
    layer0_outputs(3859) <= 1'b1;
    layer0_outputs(3860) <= a;
    layer0_outputs(3861) <= not (a xor b);
    layer0_outputs(3862) <= not a or b;
    layer0_outputs(3863) <= not b or a;
    layer0_outputs(3864) <= a xor b;
    layer0_outputs(3865) <= a;
    layer0_outputs(3866) <= not b or a;
    layer0_outputs(3867) <= a or b;
    layer0_outputs(3868) <= not b;
    layer0_outputs(3869) <= b;
    layer0_outputs(3870) <= a;
    layer0_outputs(3871) <= not a or b;
    layer0_outputs(3872) <= b and not a;
    layer0_outputs(3873) <= not a or b;
    layer0_outputs(3874) <= not (a or b);
    layer0_outputs(3875) <= 1'b0;
    layer0_outputs(3876) <= not (a xor b);
    layer0_outputs(3877) <= a;
    layer0_outputs(3878) <= a or b;
    layer0_outputs(3879) <= not a or b;
    layer0_outputs(3880) <= a or b;
    layer0_outputs(3881) <= a and not b;
    layer0_outputs(3882) <= not (a and b);
    layer0_outputs(3883) <= a or b;
    layer0_outputs(3884) <= a or b;
    layer0_outputs(3885) <= 1'b1;
    layer0_outputs(3886) <= a xor b;
    layer0_outputs(3887) <= not (a xor b);
    layer0_outputs(3888) <= b;
    layer0_outputs(3889) <= not (a and b);
    layer0_outputs(3890) <= b;
    layer0_outputs(3891) <= 1'b1;
    layer0_outputs(3892) <= not a or b;
    layer0_outputs(3893) <= a xor b;
    layer0_outputs(3894) <= not (a and b);
    layer0_outputs(3895) <= not a or b;
    layer0_outputs(3896) <= not (a xor b);
    layer0_outputs(3897) <= a;
    layer0_outputs(3898) <= not a or b;
    layer0_outputs(3899) <= not (a xor b);
    layer0_outputs(3900) <= not (a and b);
    layer0_outputs(3901) <= a;
    layer0_outputs(3902) <= b and not a;
    layer0_outputs(3903) <= not a;
    layer0_outputs(3904) <= not (a or b);
    layer0_outputs(3905) <= not (a or b);
    layer0_outputs(3906) <= a and not b;
    layer0_outputs(3907) <= a or b;
    layer0_outputs(3908) <= not (a and b);
    layer0_outputs(3909) <= a and not b;
    layer0_outputs(3910) <= a xor b;
    layer0_outputs(3911) <= b;
    layer0_outputs(3912) <= not (a xor b);
    layer0_outputs(3913) <= a xor b;
    layer0_outputs(3914) <= not (a xor b);
    layer0_outputs(3915) <= a or b;
    layer0_outputs(3916) <= a;
    layer0_outputs(3917) <= not a or b;
    layer0_outputs(3918) <= not b;
    layer0_outputs(3919) <= not b or a;
    layer0_outputs(3920) <= not b or a;
    layer0_outputs(3921) <= not (a or b);
    layer0_outputs(3922) <= not b;
    layer0_outputs(3923) <= a;
    layer0_outputs(3924) <= not (a xor b);
    layer0_outputs(3925) <= a or b;
    layer0_outputs(3926) <= a or b;
    layer0_outputs(3927) <= a or b;
    layer0_outputs(3928) <= 1'b1;
    layer0_outputs(3929) <= a xor b;
    layer0_outputs(3930) <= not b or a;
    layer0_outputs(3931) <= not a or b;
    layer0_outputs(3932) <= not b;
    layer0_outputs(3933) <= not a;
    layer0_outputs(3934) <= not (a xor b);
    layer0_outputs(3935) <= a;
    layer0_outputs(3936) <= not (a and b);
    layer0_outputs(3937) <= not b or a;
    layer0_outputs(3938) <= a or b;
    layer0_outputs(3939) <= b and not a;
    layer0_outputs(3940) <= b;
    layer0_outputs(3941) <= not b;
    layer0_outputs(3942) <= not (a or b);
    layer0_outputs(3943) <= a and not b;
    layer0_outputs(3944) <= not (a and b);
    layer0_outputs(3945) <= b;
    layer0_outputs(3946) <= 1'b0;
    layer0_outputs(3947) <= a xor b;
    layer0_outputs(3948) <= not (a or b);
    layer0_outputs(3949) <= a and not b;
    layer0_outputs(3950) <= a and not b;
    layer0_outputs(3951) <= a or b;
    layer0_outputs(3952) <= a xor b;
    layer0_outputs(3953) <= a xor b;
    layer0_outputs(3954) <= not b;
    layer0_outputs(3955) <= a and not b;
    layer0_outputs(3956) <= not (a xor b);
    layer0_outputs(3957) <= not a;
    layer0_outputs(3958) <= not (a or b);
    layer0_outputs(3959) <= not b;
    layer0_outputs(3960) <= a xor b;
    layer0_outputs(3961) <= a xor b;
    layer0_outputs(3962) <= a;
    layer0_outputs(3963) <= a;
    layer0_outputs(3964) <= a or b;
    layer0_outputs(3965) <= 1'b0;
    layer0_outputs(3966) <= b;
    layer0_outputs(3967) <= a;
    layer0_outputs(3968) <= not (a or b);
    layer0_outputs(3969) <= not (a or b);
    layer0_outputs(3970) <= a or b;
    layer0_outputs(3971) <= not a;
    layer0_outputs(3972) <= not a;
    layer0_outputs(3973) <= a and not b;
    layer0_outputs(3974) <= not a;
    layer0_outputs(3975) <= not (a or b);
    layer0_outputs(3976) <= not (a or b);
    layer0_outputs(3977) <= not b;
    layer0_outputs(3978) <= b and not a;
    layer0_outputs(3979) <= b;
    layer0_outputs(3980) <= not a or b;
    layer0_outputs(3981) <= a or b;
    layer0_outputs(3982) <= b and not a;
    layer0_outputs(3983) <= a;
    layer0_outputs(3984) <= a;
    layer0_outputs(3985) <= not b or a;
    layer0_outputs(3986) <= not (a xor b);
    layer0_outputs(3987) <= not (a or b);
    layer0_outputs(3988) <= a and not b;
    layer0_outputs(3989) <= a or b;
    layer0_outputs(3990) <= not a or b;
    layer0_outputs(3991) <= a and not b;
    layer0_outputs(3992) <= not (a and b);
    layer0_outputs(3993) <= a xor b;
    layer0_outputs(3994) <= not a or b;
    layer0_outputs(3995) <= a or b;
    layer0_outputs(3996) <= not b or a;
    layer0_outputs(3997) <= a xor b;
    layer0_outputs(3998) <= not b;
    layer0_outputs(3999) <= b and not a;
    layer0_outputs(4000) <= a and b;
    layer0_outputs(4001) <= not (a xor b);
    layer0_outputs(4002) <= not b or a;
    layer0_outputs(4003) <= not b or a;
    layer0_outputs(4004) <= not (a or b);
    layer0_outputs(4005) <= b and not a;
    layer0_outputs(4006) <= b and not a;
    layer0_outputs(4007) <= not (a xor b);
    layer0_outputs(4008) <= a or b;
    layer0_outputs(4009) <= not (a or b);
    layer0_outputs(4010) <= a and b;
    layer0_outputs(4011) <= 1'b0;
    layer0_outputs(4012) <= not a;
    layer0_outputs(4013) <= not a or b;
    layer0_outputs(4014) <= b;
    layer0_outputs(4015) <= not (a or b);
    layer0_outputs(4016) <= a xor b;
    layer0_outputs(4017) <= a and not b;
    layer0_outputs(4018) <= not a or b;
    layer0_outputs(4019) <= b and not a;
    layer0_outputs(4020) <= not a or b;
    layer0_outputs(4021) <= a;
    layer0_outputs(4022) <= not (a xor b);
    layer0_outputs(4023) <= a or b;
    layer0_outputs(4024) <= not (a or b);
    layer0_outputs(4025) <= a and not b;
    layer0_outputs(4026) <= not (a xor b);
    layer0_outputs(4027) <= a xor b;
    layer0_outputs(4028) <= b and not a;
    layer0_outputs(4029) <= a xor b;
    layer0_outputs(4030) <= not b or a;
    layer0_outputs(4031) <= not a;
    layer0_outputs(4032) <= b and not a;
    layer0_outputs(4033) <= not a or b;
    layer0_outputs(4034) <= not a or b;
    layer0_outputs(4035) <= not b or a;
    layer0_outputs(4036) <= not (a xor b);
    layer0_outputs(4037) <= a xor b;
    layer0_outputs(4038) <= not (a or b);
    layer0_outputs(4039) <= 1'b0;
    layer0_outputs(4040) <= not (a or b);
    layer0_outputs(4041) <= not (a or b);
    layer0_outputs(4042) <= a or b;
    layer0_outputs(4043) <= a and b;
    layer0_outputs(4044) <= not b;
    layer0_outputs(4045) <= not (a xor b);
    layer0_outputs(4046) <= not a;
    layer0_outputs(4047) <= not (a and b);
    layer0_outputs(4048) <= a;
    layer0_outputs(4049) <= a or b;
    layer0_outputs(4050) <= not (a and b);
    layer0_outputs(4051) <= not (a and b);
    layer0_outputs(4052) <= b;
    layer0_outputs(4053) <= a or b;
    layer0_outputs(4054) <= 1'b0;
    layer0_outputs(4055) <= a xor b;
    layer0_outputs(4056) <= not b or a;
    layer0_outputs(4057) <= not a;
    layer0_outputs(4058) <= a xor b;
    layer0_outputs(4059) <= not b or a;
    layer0_outputs(4060) <= not b or a;
    layer0_outputs(4061) <= not (a or b);
    layer0_outputs(4062) <= not (a or b);
    layer0_outputs(4063) <= b and not a;
    layer0_outputs(4064) <= a or b;
    layer0_outputs(4065) <= not (a xor b);
    layer0_outputs(4066) <= not b;
    layer0_outputs(4067) <= 1'b1;
    layer0_outputs(4068) <= 1'b1;
    layer0_outputs(4069) <= b and not a;
    layer0_outputs(4070) <= a or b;
    layer0_outputs(4071) <= b and not a;
    layer0_outputs(4072) <= not b or a;
    layer0_outputs(4073) <= not (a or b);
    layer0_outputs(4074) <= not a;
    layer0_outputs(4075) <= a xor b;
    layer0_outputs(4076) <= not (a or b);
    layer0_outputs(4077) <= not b;
    layer0_outputs(4078) <= not (a or b);
    layer0_outputs(4079) <= not a;
    layer0_outputs(4080) <= not (a or b);
    layer0_outputs(4081) <= b;
    layer0_outputs(4082) <= not (a or b);
    layer0_outputs(4083) <= a and not b;
    layer0_outputs(4084) <= b and not a;
    layer0_outputs(4085) <= a or b;
    layer0_outputs(4086) <= a and b;
    layer0_outputs(4087) <= not (a or b);
    layer0_outputs(4088) <= 1'b1;
    layer0_outputs(4089) <= a and not b;
    layer0_outputs(4090) <= a;
    layer0_outputs(4091) <= not b or a;
    layer0_outputs(4092) <= not b;
    layer0_outputs(4093) <= not (a xor b);
    layer0_outputs(4094) <= not a;
    layer0_outputs(4095) <= not (a or b);
    layer0_outputs(4096) <= b;
    layer0_outputs(4097) <= b;
    layer0_outputs(4098) <= not b or a;
    layer0_outputs(4099) <= b and not a;
    layer0_outputs(4100) <= a or b;
    layer0_outputs(4101) <= a and not b;
    layer0_outputs(4102) <= b and not a;
    layer0_outputs(4103) <= not (a xor b);
    layer0_outputs(4104) <= not a;
    layer0_outputs(4105) <= a xor b;
    layer0_outputs(4106) <= a or b;
    layer0_outputs(4107) <= b;
    layer0_outputs(4108) <= not (a xor b);
    layer0_outputs(4109) <= a;
    layer0_outputs(4110) <= not b;
    layer0_outputs(4111) <= not a or b;
    layer0_outputs(4112) <= not (a xor b);
    layer0_outputs(4113) <= b and not a;
    layer0_outputs(4114) <= not (a or b);
    layer0_outputs(4115) <= a or b;
    layer0_outputs(4116) <= not a;
    layer0_outputs(4117) <= not a;
    layer0_outputs(4118) <= not (a or b);
    layer0_outputs(4119) <= 1'b1;
    layer0_outputs(4120) <= a or b;
    layer0_outputs(4121) <= 1'b0;
    layer0_outputs(4122) <= 1'b0;
    layer0_outputs(4123) <= not a;
    layer0_outputs(4124) <= a;
    layer0_outputs(4125) <= 1'b0;
    layer0_outputs(4126) <= a xor b;
    layer0_outputs(4127) <= a xor b;
    layer0_outputs(4128) <= not (a or b);
    layer0_outputs(4129) <= not a or b;
    layer0_outputs(4130) <= 1'b1;
    layer0_outputs(4131) <= a or b;
    layer0_outputs(4132) <= a;
    layer0_outputs(4133) <= not (a or b);
    layer0_outputs(4134) <= not (a and b);
    layer0_outputs(4135) <= a;
    layer0_outputs(4136) <= not a;
    layer0_outputs(4137) <= a;
    layer0_outputs(4138) <= not a or b;
    layer0_outputs(4139) <= not b or a;
    layer0_outputs(4140) <= not (a and b);
    layer0_outputs(4141) <= a and not b;
    layer0_outputs(4142) <= not b or a;
    layer0_outputs(4143) <= a;
    layer0_outputs(4144) <= a;
    layer0_outputs(4145) <= not (a or b);
    layer0_outputs(4146) <= not (a xor b);
    layer0_outputs(4147) <= not b;
    layer0_outputs(4148) <= a or b;
    layer0_outputs(4149) <= 1'b1;
    layer0_outputs(4150) <= b and not a;
    layer0_outputs(4151) <= a xor b;
    layer0_outputs(4152) <= a;
    layer0_outputs(4153) <= a or b;
    layer0_outputs(4154) <= a or b;
    layer0_outputs(4155) <= not b;
    layer0_outputs(4156) <= b;
    layer0_outputs(4157) <= b;
    layer0_outputs(4158) <= a xor b;
    layer0_outputs(4159) <= not b;
    layer0_outputs(4160) <= 1'b1;
    layer0_outputs(4161) <= not b;
    layer0_outputs(4162) <= not b or a;
    layer0_outputs(4163) <= a and not b;
    layer0_outputs(4164) <= not (a or b);
    layer0_outputs(4165) <= not (a or b);
    layer0_outputs(4166) <= b;
    layer0_outputs(4167) <= not (a xor b);
    layer0_outputs(4168) <= not b;
    layer0_outputs(4169) <= not (a or b);
    layer0_outputs(4170) <= not (a xor b);
    layer0_outputs(4171) <= a and not b;
    layer0_outputs(4172) <= a xor b;
    layer0_outputs(4173) <= 1'b1;
    layer0_outputs(4174) <= a xor b;
    layer0_outputs(4175) <= not (a or b);
    layer0_outputs(4176) <= b and not a;
    layer0_outputs(4177) <= a;
    layer0_outputs(4178) <= a or b;
    layer0_outputs(4179) <= a or b;
    layer0_outputs(4180) <= not a or b;
    layer0_outputs(4181) <= not a or b;
    layer0_outputs(4182) <= b;
    layer0_outputs(4183) <= a and b;
    layer0_outputs(4184) <= not a;
    layer0_outputs(4185) <= not a or b;
    layer0_outputs(4186) <= not (a or b);
    layer0_outputs(4187) <= not (a or b);
    layer0_outputs(4188) <= 1'b0;
    layer0_outputs(4189) <= not (a or b);
    layer0_outputs(4190) <= a or b;
    layer0_outputs(4191) <= a or b;
    layer0_outputs(4192) <= 1'b1;
    layer0_outputs(4193) <= a or b;
    layer0_outputs(4194) <= not (a or b);
    layer0_outputs(4195) <= not (a or b);
    layer0_outputs(4196) <= a or b;
    layer0_outputs(4197) <= a or b;
    layer0_outputs(4198) <= not (a xor b);
    layer0_outputs(4199) <= a;
    layer0_outputs(4200) <= not b or a;
    layer0_outputs(4201) <= not a or b;
    layer0_outputs(4202) <= not b;
    layer0_outputs(4203) <= b;
    layer0_outputs(4204) <= a and not b;
    layer0_outputs(4205) <= 1'b0;
    layer0_outputs(4206) <= a and b;
    layer0_outputs(4207) <= 1'b1;
    layer0_outputs(4208) <= b and not a;
    layer0_outputs(4209) <= b and not a;
    layer0_outputs(4210) <= not b;
    layer0_outputs(4211) <= not a or b;
    layer0_outputs(4212) <= b;
    layer0_outputs(4213) <= a or b;
    layer0_outputs(4214) <= a xor b;
    layer0_outputs(4215) <= b and not a;
    layer0_outputs(4216) <= a and not b;
    layer0_outputs(4217) <= not a or b;
    layer0_outputs(4218) <= not a or b;
    layer0_outputs(4219) <= a and not b;
    layer0_outputs(4220) <= not (a xor b);
    layer0_outputs(4221) <= a;
    layer0_outputs(4222) <= not a or b;
    layer0_outputs(4223) <= a xor b;
    layer0_outputs(4224) <= not a or b;
    layer0_outputs(4225) <= a;
    layer0_outputs(4226) <= b;
    layer0_outputs(4227) <= not (a xor b);
    layer0_outputs(4228) <= not (a xor b);
    layer0_outputs(4229) <= a and b;
    layer0_outputs(4230) <= not a or b;
    layer0_outputs(4231) <= a and not b;
    layer0_outputs(4232) <= b;
    layer0_outputs(4233) <= b;
    layer0_outputs(4234) <= not (a xor b);
    layer0_outputs(4235) <= not a or b;
    layer0_outputs(4236) <= not a;
    layer0_outputs(4237) <= b and not a;
    layer0_outputs(4238) <= b and not a;
    layer0_outputs(4239) <= a and b;
    layer0_outputs(4240) <= not a or b;
    layer0_outputs(4241) <= a and not b;
    layer0_outputs(4242) <= not (a or b);
    layer0_outputs(4243) <= not b or a;
    layer0_outputs(4244) <= not (a or b);
    layer0_outputs(4245) <= a xor b;
    layer0_outputs(4246) <= b;
    layer0_outputs(4247) <= b;
    layer0_outputs(4248) <= a and not b;
    layer0_outputs(4249) <= a;
    layer0_outputs(4250) <= a or b;
    layer0_outputs(4251) <= not (a or b);
    layer0_outputs(4252) <= a and b;
    layer0_outputs(4253) <= 1'b1;
    layer0_outputs(4254) <= a xor b;
    layer0_outputs(4255) <= b and not a;
    layer0_outputs(4256) <= not a or b;
    layer0_outputs(4257) <= a xor b;
    layer0_outputs(4258) <= 1'b1;
    layer0_outputs(4259) <= not (a or b);
    layer0_outputs(4260) <= not (a or b);
    layer0_outputs(4261) <= not (a or b);
    layer0_outputs(4262) <= not b;
    layer0_outputs(4263) <= a or b;
    layer0_outputs(4264) <= not (a or b);
    layer0_outputs(4265) <= 1'b0;
    layer0_outputs(4266) <= not a;
    layer0_outputs(4267) <= a or b;
    layer0_outputs(4268) <= b and not a;
    layer0_outputs(4269) <= a;
    layer0_outputs(4270) <= not a;
    layer0_outputs(4271) <= 1'b0;
    layer0_outputs(4272) <= not a or b;
    layer0_outputs(4273) <= a or b;
    layer0_outputs(4274) <= not (a xor b);
    layer0_outputs(4275) <= not a;
    layer0_outputs(4276) <= not (a xor b);
    layer0_outputs(4277) <= b and not a;
    layer0_outputs(4278) <= a xor b;
    layer0_outputs(4279) <= not a or b;
    layer0_outputs(4280) <= not (a or b);
    layer0_outputs(4281) <= not a or b;
    layer0_outputs(4282) <= not b or a;
    layer0_outputs(4283) <= not b;
    layer0_outputs(4284) <= a;
    layer0_outputs(4285) <= not (a or b);
    layer0_outputs(4286) <= a or b;
    layer0_outputs(4287) <= 1'b0;
    layer0_outputs(4288) <= not b;
    layer0_outputs(4289) <= not a;
    layer0_outputs(4290) <= b;
    layer0_outputs(4291) <= a or b;
    layer0_outputs(4292) <= not a or b;
    layer0_outputs(4293) <= b;
    layer0_outputs(4294) <= not (a and b);
    layer0_outputs(4295) <= a and b;
    layer0_outputs(4296) <= a or b;
    layer0_outputs(4297) <= b and not a;
    layer0_outputs(4298) <= a and not b;
    layer0_outputs(4299) <= a or b;
    layer0_outputs(4300) <= a or b;
    layer0_outputs(4301) <= not (a or b);
    layer0_outputs(4302) <= a or b;
    layer0_outputs(4303) <= not (a or b);
    layer0_outputs(4304) <= a;
    layer0_outputs(4305) <= b and not a;
    layer0_outputs(4306) <= not a;
    layer0_outputs(4307) <= not (a or b);
    layer0_outputs(4308) <= not a;
    layer0_outputs(4309) <= not a;
    layer0_outputs(4310) <= not b;
    layer0_outputs(4311) <= b and not a;
    layer0_outputs(4312) <= not b or a;
    layer0_outputs(4313) <= a;
    layer0_outputs(4314) <= a and not b;
    layer0_outputs(4315) <= a xor b;
    layer0_outputs(4316) <= not a;
    layer0_outputs(4317) <= not a or b;
    layer0_outputs(4318) <= not (a or b);
    layer0_outputs(4319) <= b;
    layer0_outputs(4320) <= a;
    layer0_outputs(4321) <= a;
    layer0_outputs(4322) <= not b or a;
    layer0_outputs(4323) <= 1'b1;
    layer0_outputs(4324) <= a or b;
    layer0_outputs(4325) <= not (a or b);
    layer0_outputs(4326) <= b and not a;
    layer0_outputs(4327) <= not b or a;
    layer0_outputs(4328) <= not (a xor b);
    layer0_outputs(4329) <= not a;
    layer0_outputs(4330) <= not a;
    layer0_outputs(4331) <= b and not a;
    layer0_outputs(4332) <= not (a or b);
    layer0_outputs(4333) <= a or b;
    layer0_outputs(4334) <= not b or a;
    layer0_outputs(4335) <= a;
    layer0_outputs(4336) <= not b or a;
    layer0_outputs(4337) <= a and not b;
    layer0_outputs(4338) <= b and not a;
    layer0_outputs(4339) <= not b;
    layer0_outputs(4340) <= a or b;
    layer0_outputs(4341) <= not (a or b);
    layer0_outputs(4342) <= not a or b;
    layer0_outputs(4343) <= not (a or b);
    layer0_outputs(4344) <= not b;
    layer0_outputs(4345) <= a xor b;
    layer0_outputs(4346) <= not (a xor b);
    layer0_outputs(4347) <= not b;
    layer0_outputs(4348) <= b;
    layer0_outputs(4349) <= not a or b;
    layer0_outputs(4350) <= not b;
    layer0_outputs(4351) <= a xor b;
    layer0_outputs(4352) <= not a or b;
    layer0_outputs(4353) <= not a;
    layer0_outputs(4354) <= b;
    layer0_outputs(4355) <= not a;
    layer0_outputs(4356) <= b;
    layer0_outputs(4357) <= a;
    layer0_outputs(4358) <= b and not a;
    layer0_outputs(4359) <= a and b;
    layer0_outputs(4360) <= 1'b0;
    layer0_outputs(4361) <= b;
    layer0_outputs(4362) <= not a or b;
    layer0_outputs(4363) <= a and not b;
    layer0_outputs(4364) <= not b;
    layer0_outputs(4365) <= not a or b;
    layer0_outputs(4366) <= not (a xor b);
    layer0_outputs(4367) <= not (a or b);
    layer0_outputs(4368) <= not b;
    layer0_outputs(4369) <= not a or b;
    layer0_outputs(4370) <= a;
    layer0_outputs(4371) <= a xor b;
    layer0_outputs(4372) <= not b;
    layer0_outputs(4373) <= a or b;
    layer0_outputs(4374) <= not b or a;
    layer0_outputs(4375) <= not (a or b);
    layer0_outputs(4376) <= not (a and b);
    layer0_outputs(4377) <= a and not b;
    layer0_outputs(4378) <= a and not b;
    layer0_outputs(4379) <= not (a and b);
    layer0_outputs(4380) <= 1'b1;
    layer0_outputs(4381) <= not a or b;
    layer0_outputs(4382) <= b;
    layer0_outputs(4383) <= not (a and b);
    layer0_outputs(4384) <= b and not a;
    layer0_outputs(4385) <= a or b;
    layer0_outputs(4386) <= not b;
    layer0_outputs(4387) <= a xor b;
    layer0_outputs(4388) <= a or b;
    layer0_outputs(4389) <= b;
    layer0_outputs(4390) <= not b;
    layer0_outputs(4391) <= a or b;
    layer0_outputs(4392) <= not (a or b);
    layer0_outputs(4393) <= b;
    layer0_outputs(4394) <= not a or b;
    layer0_outputs(4395) <= not (a or b);
    layer0_outputs(4396) <= a and b;
    layer0_outputs(4397) <= a and b;
    layer0_outputs(4398) <= not (a xor b);
    layer0_outputs(4399) <= a and not b;
    layer0_outputs(4400) <= not b or a;
    layer0_outputs(4401) <= not a or b;
    layer0_outputs(4402) <= not b or a;
    layer0_outputs(4403) <= not (a or b);
    layer0_outputs(4404) <= not b or a;
    layer0_outputs(4405) <= a or b;
    layer0_outputs(4406) <= not a or b;
    layer0_outputs(4407) <= a and not b;
    layer0_outputs(4408) <= not (a and b);
    layer0_outputs(4409) <= not (a xor b);
    layer0_outputs(4410) <= a xor b;
    layer0_outputs(4411) <= not (a or b);
    layer0_outputs(4412) <= not (a or b);
    layer0_outputs(4413) <= b and not a;
    layer0_outputs(4414) <= not (a or b);
    layer0_outputs(4415) <= not a;
    layer0_outputs(4416) <= a or b;
    layer0_outputs(4417) <= not a or b;
    layer0_outputs(4418) <= a and b;
    layer0_outputs(4419) <= 1'b0;
    layer0_outputs(4420) <= not b or a;
    layer0_outputs(4421) <= a or b;
    layer0_outputs(4422) <= a;
    layer0_outputs(4423) <= a xor b;
    layer0_outputs(4424) <= a or b;
    layer0_outputs(4425) <= b and not a;
    layer0_outputs(4426) <= not a;
    layer0_outputs(4427) <= a or b;
    layer0_outputs(4428) <= not (a or b);
    layer0_outputs(4429) <= not a or b;
    layer0_outputs(4430) <= not (a and b);
    layer0_outputs(4431) <= not a;
    layer0_outputs(4432) <= a;
    layer0_outputs(4433) <= not b or a;
    layer0_outputs(4434) <= 1'b0;
    layer0_outputs(4435) <= a and not b;
    layer0_outputs(4436) <= not a;
    layer0_outputs(4437) <= b;
    layer0_outputs(4438) <= not b;
    layer0_outputs(4439) <= not (a xor b);
    layer0_outputs(4440) <= not a or b;
    layer0_outputs(4441) <= not b;
    layer0_outputs(4442) <= not (a or b);
    layer0_outputs(4443) <= a or b;
    layer0_outputs(4444) <= not a or b;
    layer0_outputs(4445) <= a and not b;
    layer0_outputs(4446) <= not (a xor b);
    layer0_outputs(4447) <= not (a xor b);
    layer0_outputs(4448) <= a or b;
    layer0_outputs(4449) <= not (a or b);
    layer0_outputs(4450) <= not (a and b);
    layer0_outputs(4451) <= not (a or b);
    layer0_outputs(4452) <= a or b;
    layer0_outputs(4453) <= b;
    layer0_outputs(4454) <= not (a or b);
    layer0_outputs(4455) <= not b;
    layer0_outputs(4456) <= a;
    layer0_outputs(4457) <= not b;
    layer0_outputs(4458) <= b and not a;
    layer0_outputs(4459) <= not (a or b);
    layer0_outputs(4460) <= not a;
    layer0_outputs(4461) <= not b;
    layer0_outputs(4462) <= b and not a;
    layer0_outputs(4463) <= 1'b1;
    layer0_outputs(4464) <= not (a xor b);
    layer0_outputs(4465) <= a xor b;
    layer0_outputs(4466) <= 1'b1;
    layer0_outputs(4467) <= not (a and b);
    layer0_outputs(4468) <= b and not a;
    layer0_outputs(4469) <= a xor b;
    layer0_outputs(4470) <= a or b;
    layer0_outputs(4471) <= b and not a;
    layer0_outputs(4472) <= not (a xor b);
    layer0_outputs(4473) <= b and not a;
    layer0_outputs(4474) <= not b;
    layer0_outputs(4475) <= not (a xor b);
    layer0_outputs(4476) <= not a or b;
    layer0_outputs(4477) <= not b;
    layer0_outputs(4478) <= 1'b0;
    layer0_outputs(4479) <= a or b;
    layer0_outputs(4480) <= not b;
    layer0_outputs(4481) <= a or b;
    layer0_outputs(4482) <= not (a or b);
    layer0_outputs(4483) <= not (a or b);
    layer0_outputs(4484) <= not a;
    layer0_outputs(4485) <= not (a or b);
    layer0_outputs(4486) <= not a or b;
    layer0_outputs(4487) <= not (a and b);
    layer0_outputs(4488) <= not b or a;
    layer0_outputs(4489) <= a or b;
    layer0_outputs(4490) <= 1'b0;
    layer0_outputs(4491) <= b and not a;
    layer0_outputs(4492) <= not a or b;
    layer0_outputs(4493) <= a;
    layer0_outputs(4494) <= a or b;
    layer0_outputs(4495) <= a or b;
    layer0_outputs(4496) <= a or b;
    layer0_outputs(4497) <= not a;
    layer0_outputs(4498) <= 1'b1;
    layer0_outputs(4499) <= not (a or b);
    layer0_outputs(4500) <= b and not a;
    layer0_outputs(4501) <= not (a or b);
    layer0_outputs(4502) <= a xor b;
    layer0_outputs(4503) <= b;
    layer0_outputs(4504) <= b;
    layer0_outputs(4505) <= 1'b0;
    layer0_outputs(4506) <= not a;
    layer0_outputs(4507) <= not (a or b);
    layer0_outputs(4508) <= a and not b;
    layer0_outputs(4509) <= a or b;
    layer0_outputs(4510) <= b and not a;
    layer0_outputs(4511) <= a or b;
    layer0_outputs(4512) <= not b;
    layer0_outputs(4513) <= a xor b;
    layer0_outputs(4514) <= not (a or b);
    layer0_outputs(4515) <= not (a or b);
    layer0_outputs(4516) <= not (a or b);
    layer0_outputs(4517) <= a;
    layer0_outputs(4518) <= not b;
    layer0_outputs(4519) <= a and not b;
    layer0_outputs(4520) <= not a;
    layer0_outputs(4521) <= a and not b;
    layer0_outputs(4522) <= a or b;
    layer0_outputs(4523) <= a or b;
    layer0_outputs(4524) <= not a;
    layer0_outputs(4525) <= 1'b1;
    layer0_outputs(4526) <= 1'b1;
    layer0_outputs(4527) <= 1'b1;
    layer0_outputs(4528) <= a xor b;
    layer0_outputs(4529) <= b;
    layer0_outputs(4530) <= a and b;
    layer0_outputs(4531) <= a xor b;
    layer0_outputs(4532) <= not (a or b);
    layer0_outputs(4533) <= not a;
    layer0_outputs(4534) <= a;
    layer0_outputs(4535) <= a;
    layer0_outputs(4536) <= not (a xor b);
    layer0_outputs(4537) <= b;
    layer0_outputs(4538) <= not a or b;
    layer0_outputs(4539) <= a or b;
    layer0_outputs(4540) <= not a;
    layer0_outputs(4541) <= a xor b;
    layer0_outputs(4542) <= not b;
    layer0_outputs(4543) <= 1'b1;
    layer0_outputs(4544) <= 1'b0;
    layer0_outputs(4545) <= not a or b;
    layer0_outputs(4546) <= not (a xor b);
    layer0_outputs(4547) <= a and not b;
    layer0_outputs(4548) <= not a;
    layer0_outputs(4549) <= not a or b;
    layer0_outputs(4550) <= a or b;
    layer0_outputs(4551) <= not (a or b);
    layer0_outputs(4552) <= b;
    layer0_outputs(4553) <= b;
    layer0_outputs(4554) <= not b;
    layer0_outputs(4555) <= a;
    layer0_outputs(4556) <= b;
    layer0_outputs(4557) <= a or b;
    layer0_outputs(4558) <= a or b;
    layer0_outputs(4559) <= a and b;
    layer0_outputs(4560) <= a or b;
    layer0_outputs(4561) <= a;
    layer0_outputs(4562) <= not a;
    layer0_outputs(4563) <= not b;
    layer0_outputs(4564) <= not (a or b);
    layer0_outputs(4565) <= b;
    layer0_outputs(4566) <= not (a and b);
    layer0_outputs(4567) <= not b;
    layer0_outputs(4568) <= a and not b;
    layer0_outputs(4569) <= not a or b;
    layer0_outputs(4570) <= a and not b;
    layer0_outputs(4571) <= not (a xor b);
    layer0_outputs(4572) <= a or b;
    layer0_outputs(4573) <= not a;
    layer0_outputs(4574) <= b and not a;
    layer0_outputs(4575) <= not b;
    layer0_outputs(4576) <= not a;
    layer0_outputs(4577) <= not b;
    layer0_outputs(4578) <= a or b;
    layer0_outputs(4579) <= not (a xor b);
    layer0_outputs(4580) <= b;
    layer0_outputs(4581) <= a and not b;
    layer0_outputs(4582) <= not (a xor b);
    layer0_outputs(4583) <= not a or b;
    layer0_outputs(4584) <= a or b;
    layer0_outputs(4585) <= b;
    layer0_outputs(4586) <= not b or a;
    layer0_outputs(4587) <= a and not b;
    layer0_outputs(4588) <= not b or a;
    layer0_outputs(4589) <= not b;
    layer0_outputs(4590) <= b and not a;
    layer0_outputs(4591) <= not b or a;
    layer0_outputs(4592) <= a and not b;
    layer0_outputs(4593) <= b;
    layer0_outputs(4594) <= not (a or b);
    layer0_outputs(4595) <= not a;
    layer0_outputs(4596) <= not (a or b);
    layer0_outputs(4597) <= b and not a;
    layer0_outputs(4598) <= not b;
    layer0_outputs(4599) <= not (a xor b);
    layer0_outputs(4600) <= a or b;
    layer0_outputs(4601) <= a and not b;
    layer0_outputs(4602) <= b;
    layer0_outputs(4603) <= 1'b0;
    layer0_outputs(4604) <= a;
    layer0_outputs(4605) <= b;
    layer0_outputs(4606) <= not b;
    layer0_outputs(4607) <= b and not a;
    layer0_outputs(4608) <= a xor b;
    layer0_outputs(4609) <= b;
    layer0_outputs(4610) <= not (a or b);
    layer0_outputs(4611) <= a xor b;
    layer0_outputs(4612) <= 1'b0;
    layer0_outputs(4613) <= a;
    layer0_outputs(4614) <= not (a xor b);
    layer0_outputs(4615) <= a xor b;
    layer0_outputs(4616) <= a;
    layer0_outputs(4617) <= not a;
    layer0_outputs(4618) <= not b;
    layer0_outputs(4619) <= not b or a;
    layer0_outputs(4620) <= not (a xor b);
    layer0_outputs(4621) <= a or b;
    layer0_outputs(4622) <= a and not b;
    layer0_outputs(4623) <= a xor b;
    layer0_outputs(4624) <= a;
    layer0_outputs(4625) <= not a;
    layer0_outputs(4626) <= not b;
    layer0_outputs(4627) <= not a;
    layer0_outputs(4628) <= a;
    layer0_outputs(4629) <= not (a xor b);
    layer0_outputs(4630) <= not b or a;
    layer0_outputs(4631) <= b;
    layer0_outputs(4632) <= a and b;
    layer0_outputs(4633) <= not (a or b);
    layer0_outputs(4634) <= a or b;
    layer0_outputs(4635) <= b;
    layer0_outputs(4636) <= b and not a;
    layer0_outputs(4637) <= not b or a;
    layer0_outputs(4638) <= a or b;
    layer0_outputs(4639) <= not b;
    layer0_outputs(4640) <= not (a or b);
    layer0_outputs(4641) <= not b;
    layer0_outputs(4642) <= a;
    layer0_outputs(4643) <= b;
    layer0_outputs(4644) <= b and not a;
    layer0_outputs(4645) <= a or b;
    layer0_outputs(4646) <= a or b;
    layer0_outputs(4647) <= a or b;
    layer0_outputs(4648) <= b and not a;
    layer0_outputs(4649) <= a;
    layer0_outputs(4650) <= not b or a;
    layer0_outputs(4651) <= b;
    layer0_outputs(4652) <= a or b;
    layer0_outputs(4653) <= not b or a;
    layer0_outputs(4654) <= a xor b;
    layer0_outputs(4655) <= not (a xor b);
    layer0_outputs(4656) <= not (a xor b);
    layer0_outputs(4657) <= a;
    layer0_outputs(4658) <= not a or b;
    layer0_outputs(4659) <= a xor b;
    layer0_outputs(4660) <= a and not b;
    layer0_outputs(4661) <= a or b;
    layer0_outputs(4662) <= 1'b1;
    layer0_outputs(4663) <= not a;
    layer0_outputs(4664) <= b;
    layer0_outputs(4665) <= b;
    layer0_outputs(4666) <= not b;
    layer0_outputs(4667) <= b and not a;
    layer0_outputs(4668) <= not b or a;
    layer0_outputs(4669) <= 1'b1;
    layer0_outputs(4670) <= not a or b;
    layer0_outputs(4671) <= 1'b0;
    layer0_outputs(4672) <= b;
    layer0_outputs(4673) <= not b or a;
    layer0_outputs(4674) <= not a or b;
    layer0_outputs(4675) <= not b or a;
    layer0_outputs(4676) <= not (a xor b);
    layer0_outputs(4677) <= not (a xor b);
    layer0_outputs(4678) <= not (a or b);
    layer0_outputs(4679) <= a and not b;
    layer0_outputs(4680) <= b;
    layer0_outputs(4681) <= a or b;
    layer0_outputs(4682) <= not b or a;
    layer0_outputs(4683) <= not b or a;
    layer0_outputs(4684) <= not a;
    layer0_outputs(4685) <= b and not a;
    layer0_outputs(4686) <= b and not a;
    layer0_outputs(4687) <= not (a or b);
    layer0_outputs(4688) <= b and not a;
    layer0_outputs(4689) <= not (a or b);
    layer0_outputs(4690) <= not (a or b);
    layer0_outputs(4691) <= not a or b;
    layer0_outputs(4692) <= a xor b;
    layer0_outputs(4693) <= not (a or b);
    layer0_outputs(4694) <= not a;
    layer0_outputs(4695) <= b and not a;
    layer0_outputs(4696) <= not b;
    layer0_outputs(4697) <= not (a and b);
    layer0_outputs(4698) <= a xor b;
    layer0_outputs(4699) <= b;
    layer0_outputs(4700) <= a and not b;
    layer0_outputs(4701) <= a or b;
    layer0_outputs(4702) <= not a or b;
    layer0_outputs(4703) <= b;
    layer0_outputs(4704) <= not a;
    layer0_outputs(4705) <= a or b;
    layer0_outputs(4706) <= a or b;
    layer0_outputs(4707) <= not b;
    layer0_outputs(4708) <= a or b;
    layer0_outputs(4709) <= not (a and b);
    layer0_outputs(4710) <= a and not b;
    layer0_outputs(4711) <= a xor b;
    layer0_outputs(4712) <= not (a or b);
    layer0_outputs(4713) <= not (a and b);
    layer0_outputs(4714) <= 1'b1;
    layer0_outputs(4715) <= not a or b;
    layer0_outputs(4716) <= not (a or b);
    layer0_outputs(4717) <= not a;
    layer0_outputs(4718) <= a or b;
    layer0_outputs(4719) <= not b;
    layer0_outputs(4720) <= a;
    layer0_outputs(4721) <= not (a xor b);
    layer0_outputs(4722) <= a xor b;
    layer0_outputs(4723) <= a or b;
    layer0_outputs(4724) <= b;
    layer0_outputs(4725) <= not a or b;
    layer0_outputs(4726) <= a xor b;
    layer0_outputs(4727) <= a or b;
    layer0_outputs(4728) <= a and not b;
    layer0_outputs(4729) <= not a;
    layer0_outputs(4730) <= not (a and b);
    layer0_outputs(4731) <= a and not b;
    layer0_outputs(4732) <= not b or a;
    layer0_outputs(4733) <= a;
    layer0_outputs(4734) <= b;
    layer0_outputs(4735) <= not (a and b);
    layer0_outputs(4736) <= not b;
    layer0_outputs(4737) <= a and not b;
    layer0_outputs(4738) <= a and not b;
    layer0_outputs(4739) <= not (a xor b);
    layer0_outputs(4740) <= a xor b;
    layer0_outputs(4741) <= not b or a;
    layer0_outputs(4742) <= a or b;
    layer0_outputs(4743) <= b;
    layer0_outputs(4744) <= a or b;
    layer0_outputs(4745) <= not b or a;
    layer0_outputs(4746) <= not a;
    layer0_outputs(4747) <= a xor b;
    layer0_outputs(4748) <= a or b;
    layer0_outputs(4749) <= not (a xor b);
    layer0_outputs(4750) <= b and not a;
    layer0_outputs(4751) <= a;
    layer0_outputs(4752) <= b;
    layer0_outputs(4753) <= not (a xor b);
    layer0_outputs(4754) <= a xor b;
    layer0_outputs(4755) <= not (a and b);
    layer0_outputs(4756) <= not b;
    layer0_outputs(4757) <= not (a or b);
    layer0_outputs(4758) <= a or b;
    layer0_outputs(4759) <= b;
    layer0_outputs(4760) <= a and b;
    layer0_outputs(4761) <= not (a or b);
    layer0_outputs(4762) <= not b or a;
    layer0_outputs(4763) <= a xor b;
    layer0_outputs(4764) <= a or b;
    layer0_outputs(4765) <= a and not b;
    layer0_outputs(4766) <= a and not b;
    layer0_outputs(4767) <= not a;
    layer0_outputs(4768) <= a xor b;
    layer0_outputs(4769) <= not a;
    layer0_outputs(4770) <= a;
    layer0_outputs(4771) <= not (a xor b);
    layer0_outputs(4772) <= not (a or b);
    layer0_outputs(4773) <= not (a xor b);
    layer0_outputs(4774) <= a xor b;
    layer0_outputs(4775) <= a;
    layer0_outputs(4776) <= a and not b;
    layer0_outputs(4777) <= 1'b0;
    layer0_outputs(4778) <= b and not a;
    layer0_outputs(4779) <= a;
    layer0_outputs(4780) <= a xor b;
    layer0_outputs(4781) <= a or b;
    layer0_outputs(4782) <= not b or a;
    layer0_outputs(4783) <= a;
    layer0_outputs(4784) <= not (a or b);
    layer0_outputs(4785) <= not a;
    layer0_outputs(4786) <= a and not b;
    layer0_outputs(4787) <= not a;
    layer0_outputs(4788) <= a xor b;
    layer0_outputs(4789) <= 1'b1;
    layer0_outputs(4790) <= b;
    layer0_outputs(4791) <= a and not b;
    layer0_outputs(4792) <= not b;
    layer0_outputs(4793) <= b and not a;
    layer0_outputs(4794) <= not a;
    layer0_outputs(4795) <= a and b;
    layer0_outputs(4796) <= a and b;
    layer0_outputs(4797) <= not (a or b);
    layer0_outputs(4798) <= not b or a;
    layer0_outputs(4799) <= a xor b;
    layer0_outputs(4800) <= not b or a;
    layer0_outputs(4801) <= a and b;
    layer0_outputs(4802) <= not (a xor b);
    layer0_outputs(4803) <= a or b;
    layer0_outputs(4804) <= a xor b;
    layer0_outputs(4805) <= a or b;
    layer0_outputs(4806) <= b and not a;
    layer0_outputs(4807) <= not (a xor b);
    layer0_outputs(4808) <= not (a or b);
    layer0_outputs(4809) <= a or b;
    layer0_outputs(4810) <= b;
    layer0_outputs(4811) <= not b or a;
    layer0_outputs(4812) <= 1'b0;
    layer0_outputs(4813) <= not (a or b);
    layer0_outputs(4814) <= a xor b;
    layer0_outputs(4815) <= a xor b;
    layer0_outputs(4816) <= b;
    layer0_outputs(4817) <= not b;
    layer0_outputs(4818) <= 1'b1;
    layer0_outputs(4819) <= a;
    layer0_outputs(4820) <= not a;
    layer0_outputs(4821) <= not a;
    layer0_outputs(4822) <= a;
    layer0_outputs(4823) <= a;
    layer0_outputs(4824) <= not (a or b);
    layer0_outputs(4825) <= a or b;
    layer0_outputs(4826) <= a or b;
    layer0_outputs(4827) <= not b or a;
    layer0_outputs(4828) <= b;
    layer0_outputs(4829) <= b and not a;
    layer0_outputs(4830) <= a xor b;
    layer0_outputs(4831) <= not b or a;
    layer0_outputs(4832) <= not b;
    layer0_outputs(4833) <= a or b;
    layer0_outputs(4834) <= a or b;
    layer0_outputs(4835) <= a or b;
    layer0_outputs(4836) <= not (a or b);
    layer0_outputs(4837) <= not b;
    layer0_outputs(4838) <= not b or a;
    layer0_outputs(4839) <= a and not b;
    layer0_outputs(4840) <= not (a or b);
    layer0_outputs(4841) <= not a or b;
    layer0_outputs(4842) <= a or b;
    layer0_outputs(4843) <= not (a or b);
    layer0_outputs(4844) <= not (a or b);
    layer0_outputs(4845) <= not b or a;
    layer0_outputs(4846) <= not b;
    layer0_outputs(4847) <= not (a or b);
    layer0_outputs(4848) <= b;
    layer0_outputs(4849) <= b;
    layer0_outputs(4850) <= not a;
    layer0_outputs(4851) <= a and not b;
    layer0_outputs(4852) <= a and not b;
    layer0_outputs(4853) <= a or b;
    layer0_outputs(4854) <= not a;
    layer0_outputs(4855) <= a and not b;
    layer0_outputs(4856) <= not (a xor b);
    layer0_outputs(4857) <= a or b;
    layer0_outputs(4858) <= not b or a;
    layer0_outputs(4859) <= not b;
    layer0_outputs(4860) <= not b;
    layer0_outputs(4861) <= a or b;
    layer0_outputs(4862) <= a and not b;
    layer0_outputs(4863) <= a xor b;
    layer0_outputs(4864) <= not (a or b);
    layer0_outputs(4865) <= not a or b;
    layer0_outputs(4866) <= a and not b;
    layer0_outputs(4867) <= not b;
    layer0_outputs(4868) <= 1'b1;
    layer0_outputs(4869) <= not (a and b);
    layer0_outputs(4870) <= not (a or b);
    layer0_outputs(4871) <= a;
    layer0_outputs(4872) <= not b or a;
    layer0_outputs(4873) <= 1'b1;
    layer0_outputs(4874) <= not (a xor b);
    layer0_outputs(4875) <= b and not a;
    layer0_outputs(4876) <= a;
    layer0_outputs(4877) <= not b;
    layer0_outputs(4878) <= a and not b;
    layer0_outputs(4879) <= b and not a;
    layer0_outputs(4880) <= not a;
    layer0_outputs(4881) <= a;
    layer0_outputs(4882) <= a or b;
    layer0_outputs(4883) <= not b or a;
    layer0_outputs(4884) <= a xor b;
    layer0_outputs(4885) <= a xor b;
    layer0_outputs(4886) <= 1'b1;
    layer0_outputs(4887) <= not a;
    layer0_outputs(4888) <= a and b;
    layer0_outputs(4889) <= not (a or b);
    layer0_outputs(4890) <= a or b;
    layer0_outputs(4891) <= not b or a;
    layer0_outputs(4892) <= a xor b;
    layer0_outputs(4893) <= a and b;
    layer0_outputs(4894) <= a and not b;
    layer0_outputs(4895) <= 1'b1;
    layer0_outputs(4896) <= 1'b1;
    layer0_outputs(4897) <= b;
    layer0_outputs(4898) <= not b or a;
    layer0_outputs(4899) <= not a;
    layer0_outputs(4900) <= 1'b0;
    layer0_outputs(4901) <= not a or b;
    layer0_outputs(4902) <= a xor b;
    layer0_outputs(4903) <= a and b;
    layer0_outputs(4904) <= not (a xor b);
    layer0_outputs(4905) <= a and not b;
    layer0_outputs(4906) <= 1'b0;
    layer0_outputs(4907) <= not (a or b);
    layer0_outputs(4908) <= 1'b1;
    layer0_outputs(4909) <= not a or b;
    layer0_outputs(4910) <= a xor b;
    layer0_outputs(4911) <= a;
    layer0_outputs(4912) <= a or b;
    layer0_outputs(4913) <= b;
    layer0_outputs(4914) <= not b or a;
    layer0_outputs(4915) <= b;
    layer0_outputs(4916) <= b;
    layer0_outputs(4917) <= a or b;
    layer0_outputs(4918) <= a or b;
    layer0_outputs(4919) <= a or b;
    layer0_outputs(4920) <= not b;
    layer0_outputs(4921) <= a;
    layer0_outputs(4922) <= a or b;
    layer0_outputs(4923) <= a xor b;
    layer0_outputs(4924) <= not b;
    layer0_outputs(4925) <= 1'b1;
    layer0_outputs(4926) <= 1'b0;
    layer0_outputs(4927) <= not b or a;
    layer0_outputs(4928) <= 1'b0;
    layer0_outputs(4929) <= not (a or b);
    layer0_outputs(4930) <= a or b;
    layer0_outputs(4931) <= a;
    layer0_outputs(4932) <= not a;
    layer0_outputs(4933) <= b;
    layer0_outputs(4934) <= not (a or b);
    layer0_outputs(4935) <= a or b;
    layer0_outputs(4936) <= a or b;
    layer0_outputs(4937) <= a xor b;
    layer0_outputs(4938) <= 1'b1;
    layer0_outputs(4939) <= a and b;
    layer0_outputs(4940) <= a or b;
    layer0_outputs(4941) <= a or b;
    layer0_outputs(4942) <= a and not b;
    layer0_outputs(4943) <= not (a and b);
    layer0_outputs(4944) <= not (a or b);
    layer0_outputs(4945) <= not a;
    layer0_outputs(4946) <= not (a or b);
    layer0_outputs(4947) <= not b;
    layer0_outputs(4948) <= not a;
    layer0_outputs(4949) <= b and not a;
    layer0_outputs(4950) <= not (a xor b);
    layer0_outputs(4951) <= a xor b;
    layer0_outputs(4952) <= not b or a;
    layer0_outputs(4953) <= a or b;
    layer0_outputs(4954) <= a;
    layer0_outputs(4955) <= a and not b;
    layer0_outputs(4956) <= a xor b;
    layer0_outputs(4957) <= not (a or b);
    layer0_outputs(4958) <= a;
    layer0_outputs(4959) <= a and not b;
    layer0_outputs(4960) <= not a;
    layer0_outputs(4961) <= a and not b;
    layer0_outputs(4962) <= not (a xor b);
    layer0_outputs(4963) <= not b;
    layer0_outputs(4964) <= not (a or b);
    layer0_outputs(4965) <= not (a or b);
    layer0_outputs(4966) <= not (a or b);
    layer0_outputs(4967) <= a or b;
    layer0_outputs(4968) <= not (a xor b);
    layer0_outputs(4969) <= not (a or b);
    layer0_outputs(4970) <= not a;
    layer0_outputs(4971) <= not (a or b);
    layer0_outputs(4972) <= a or b;
    layer0_outputs(4973) <= not (a and b);
    layer0_outputs(4974) <= not b;
    layer0_outputs(4975) <= not (a or b);
    layer0_outputs(4976) <= a;
    layer0_outputs(4977) <= not b;
    layer0_outputs(4978) <= b;
    layer0_outputs(4979) <= not (a or b);
    layer0_outputs(4980) <= not (a xor b);
    layer0_outputs(4981) <= not a or b;
    layer0_outputs(4982) <= a and not b;
    layer0_outputs(4983) <= b and not a;
    layer0_outputs(4984) <= a and not b;
    layer0_outputs(4985) <= a or b;
    layer0_outputs(4986) <= not a or b;
    layer0_outputs(4987) <= a xor b;
    layer0_outputs(4988) <= a;
    layer0_outputs(4989) <= not a or b;
    layer0_outputs(4990) <= b;
    layer0_outputs(4991) <= not b or a;
    layer0_outputs(4992) <= not (a and b);
    layer0_outputs(4993) <= b and not a;
    layer0_outputs(4994) <= a xor b;
    layer0_outputs(4995) <= a and b;
    layer0_outputs(4996) <= not b;
    layer0_outputs(4997) <= not a or b;
    layer0_outputs(4998) <= a or b;
    layer0_outputs(4999) <= a and not b;
    layer0_outputs(5000) <= a or b;
    layer0_outputs(5001) <= a or b;
    layer0_outputs(5002) <= not a;
    layer0_outputs(5003) <= a or b;
    layer0_outputs(5004) <= not (a xor b);
    layer0_outputs(5005) <= b and not a;
    layer0_outputs(5006) <= a xor b;
    layer0_outputs(5007) <= not (a and b);
    layer0_outputs(5008) <= a;
    layer0_outputs(5009) <= not b or a;
    layer0_outputs(5010) <= not b or a;
    layer0_outputs(5011) <= not b;
    layer0_outputs(5012) <= a;
    layer0_outputs(5013) <= not (a or b);
    layer0_outputs(5014) <= not b or a;
    layer0_outputs(5015) <= not b;
    layer0_outputs(5016) <= b and not a;
    layer0_outputs(5017) <= not a;
    layer0_outputs(5018) <= a or b;
    layer0_outputs(5019) <= a and not b;
    layer0_outputs(5020) <= a or b;
    layer0_outputs(5021) <= 1'b0;
    layer0_outputs(5022) <= not (a and b);
    layer0_outputs(5023) <= not (a and b);
    layer0_outputs(5024) <= a and not b;
    layer0_outputs(5025) <= a or b;
    layer0_outputs(5026) <= 1'b0;
    layer0_outputs(5027) <= not b;
    layer0_outputs(5028) <= 1'b0;
    layer0_outputs(5029) <= a;
    layer0_outputs(5030) <= a xor b;
    layer0_outputs(5031) <= a or b;
    layer0_outputs(5032) <= not (a xor b);
    layer0_outputs(5033) <= a or b;
    layer0_outputs(5034) <= not a or b;
    layer0_outputs(5035) <= not a or b;
    layer0_outputs(5036) <= not a or b;
    layer0_outputs(5037) <= not a or b;
    layer0_outputs(5038) <= b;
    layer0_outputs(5039) <= a xor b;
    layer0_outputs(5040) <= not b or a;
    layer0_outputs(5041) <= b;
    layer0_outputs(5042) <= not (a or b);
    layer0_outputs(5043) <= a and b;
    layer0_outputs(5044) <= not (a or b);
    layer0_outputs(5045) <= a and not b;
    layer0_outputs(5046) <= a and not b;
    layer0_outputs(5047) <= not b or a;
    layer0_outputs(5048) <= not b or a;
    layer0_outputs(5049) <= not (a xor b);
    layer0_outputs(5050) <= a;
    layer0_outputs(5051) <= not (a xor b);
    layer0_outputs(5052) <= b;
    layer0_outputs(5053) <= not a or b;
    layer0_outputs(5054) <= not a or b;
    layer0_outputs(5055) <= 1'b0;
    layer0_outputs(5056) <= not (a or b);
    layer0_outputs(5057) <= a or b;
    layer0_outputs(5058) <= not a;
    layer0_outputs(5059) <= not (a or b);
    layer0_outputs(5060) <= b;
    layer0_outputs(5061) <= not (a or b);
    layer0_outputs(5062) <= not b or a;
    layer0_outputs(5063) <= not (a xor b);
    layer0_outputs(5064) <= not a;
    layer0_outputs(5065) <= not b or a;
    layer0_outputs(5066) <= a or b;
    layer0_outputs(5067) <= not a or b;
    layer0_outputs(5068) <= a;
    layer0_outputs(5069) <= not b;
    layer0_outputs(5070) <= not (a xor b);
    layer0_outputs(5071) <= not a;
    layer0_outputs(5072) <= not a;
    layer0_outputs(5073) <= b and not a;
    layer0_outputs(5074) <= b and not a;
    layer0_outputs(5075) <= not a;
    layer0_outputs(5076) <= not a or b;
    layer0_outputs(5077) <= b;
    layer0_outputs(5078) <= not a;
    layer0_outputs(5079) <= not b;
    layer0_outputs(5080) <= a or b;
    layer0_outputs(5081) <= not a or b;
    layer0_outputs(5082) <= not (a and b);
    layer0_outputs(5083) <= not (a xor b);
    layer0_outputs(5084) <= not (a or b);
    layer0_outputs(5085) <= a and not b;
    layer0_outputs(5086) <= not a;
    layer0_outputs(5087) <= not (a xor b);
    layer0_outputs(5088) <= a;
    layer0_outputs(5089) <= not b;
    layer0_outputs(5090) <= b;
    layer0_outputs(5091) <= b and not a;
    layer0_outputs(5092) <= a;
    layer0_outputs(5093) <= not b or a;
    layer0_outputs(5094) <= not (a xor b);
    layer0_outputs(5095) <= not (a xor b);
    layer0_outputs(5096) <= b and not a;
    layer0_outputs(5097) <= not (a xor b);
    layer0_outputs(5098) <= a and not b;
    layer0_outputs(5099) <= not a or b;
    layer0_outputs(5100) <= not a;
    layer0_outputs(5101) <= not b or a;
    layer0_outputs(5102) <= b and not a;
    layer0_outputs(5103) <= not (a xor b);
    layer0_outputs(5104) <= a and not b;
    layer0_outputs(5105) <= 1'b0;
    layer0_outputs(5106) <= not a or b;
    layer0_outputs(5107) <= b;
    layer0_outputs(5108) <= b;
    layer0_outputs(5109) <= b and not a;
    layer0_outputs(5110) <= not (a or b);
    layer0_outputs(5111) <= not a;
    layer0_outputs(5112) <= not a or b;
    layer0_outputs(5113) <= b;
    layer0_outputs(5114) <= a xor b;
    layer0_outputs(5115) <= a;
    layer0_outputs(5116) <= not b;
    layer0_outputs(5117) <= not a;
    layer0_outputs(5118) <= not (a xor b);
    layer0_outputs(5119) <= not b;
    layer0_outputs(5120) <= a or b;
    layer0_outputs(5121) <= a and not b;
    layer0_outputs(5122) <= b;
    layer0_outputs(5123) <= b;
    layer0_outputs(5124) <= not a;
    layer0_outputs(5125) <= b and not a;
    layer0_outputs(5126) <= a or b;
    layer0_outputs(5127) <= 1'b0;
    layer0_outputs(5128) <= a and not b;
    layer0_outputs(5129) <= a and not b;
    layer0_outputs(5130) <= b;
    layer0_outputs(5131) <= a and not b;
    layer0_outputs(5132) <= a xor b;
    layer0_outputs(5133) <= a or b;
    layer0_outputs(5134) <= not (a and b);
    layer0_outputs(5135) <= a or b;
    layer0_outputs(5136) <= not (a or b);
    layer0_outputs(5137) <= a or b;
    layer0_outputs(5138) <= not a;
    layer0_outputs(5139) <= a xor b;
    layer0_outputs(5140) <= a or b;
    layer0_outputs(5141) <= a or b;
    layer0_outputs(5142) <= not (a xor b);
    layer0_outputs(5143) <= a xor b;
    layer0_outputs(5144) <= not (a or b);
    layer0_outputs(5145) <= not a;
    layer0_outputs(5146) <= not a;
    layer0_outputs(5147) <= not b or a;
    layer0_outputs(5148) <= not a or b;
    layer0_outputs(5149) <= not (a or b);
    layer0_outputs(5150) <= not (a and b);
    layer0_outputs(5151) <= not b or a;
    layer0_outputs(5152) <= not a or b;
    layer0_outputs(5153) <= not (a or b);
    layer0_outputs(5154) <= a;
    layer0_outputs(5155) <= a xor b;
    layer0_outputs(5156) <= not a;
    layer0_outputs(5157) <= a;
    layer0_outputs(5158) <= a or b;
    layer0_outputs(5159) <= a xor b;
    layer0_outputs(5160) <= b and not a;
    layer0_outputs(5161) <= not a or b;
    layer0_outputs(5162) <= not (a xor b);
    layer0_outputs(5163) <= a and not b;
    layer0_outputs(5164) <= b and not a;
    layer0_outputs(5165) <= a xor b;
    layer0_outputs(5166) <= a;
    layer0_outputs(5167) <= a or b;
    layer0_outputs(5168) <= not (a or b);
    layer0_outputs(5169) <= not a or b;
    layer0_outputs(5170) <= not a;
    layer0_outputs(5171) <= not b or a;
    layer0_outputs(5172) <= not a or b;
    layer0_outputs(5173) <= a and not b;
    layer0_outputs(5174) <= not (a or b);
    layer0_outputs(5175) <= not (a xor b);
    layer0_outputs(5176) <= not b;
    layer0_outputs(5177) <= b;
    layer0_outputs(5178) <= a;
    layer0_outputs(5179) <= not a;
    layer0_outputs(5180) <= 1'b1;
    layer0_outputs(5181) <= not a or b;
    layer0_outputs(5182) <= not (a or b);
    layer0_outputs(5183) <= not (a xor b);
    layer0_outputs(5184) <= a or b;
    layer0_outputs(5185) <= a and not b;
    layer0_outputs(5186) <= a xor b;
    layer0_outputs(5187) <= not (a or b);
    layer0_outputs(5188) <= not a;
    layer0_outputs(5189) <= a and not b;
    layer0_outputs(5190) <= a or b;
    layer0_outputs(5191) <= b and not a;
    layer0_outputs(5192) <= a or b;
    layer0_outputs(5193) <= not (a xor b);
    layer0_outputs(5194) <= not (a xor b);
    layer0_outputs(5195) <= not a or b;
    layer0_outputs(5196) <= a;
    layer0_outputs(5197) <= a or b;
    layer0_outputs(5198) <= b and not a;
    layer0_outputs(5199) <= not a;
    layer0_outputs(5200) <= 1'b1;
    layer0_outputs(5201) <= not b or a;
    layer0_outputs(5202) <= a or b;
    layer0_outputs(5203) <= not a;
    layer0_outputs(5204) <= b and not a;
    layer0_outputs(5205) <= not b;
    layer0_outputs(5206) <= not (a and b);
    layer0_outputs(5207) <= b and not a;
    layer0_outputs(5208) <= not (a or b);
    layer0_outputs(5209) <= not b or a;
    layer0_outputs(5210) <= not b;
    layer0_outputs(5211) <= not a or b;
    layer0_outputs(5212) <= not a or b;
    layer0_outputs(5213) <= b;
    layer0_outputs(5214) <= 1'b0;
    layer0_outputs(5215) <= not a;
    layer0_outputs(5216) <= not a;
    layer0_outputs(5217) <= b;
    layer0_outputs(5218) <= a or b;
    layer0_outputs(5219) <= not (a or b);
    layer0_outputs(5220) <= 1'b1;
    layer0_outputs(5221) <= a or b;
    layer0_outputs(5222) <= a xor b;
    layer0_outputs(5223) <= 1'b0;
    layer0_outputs(5224) <= a or b;
    layer0_outputs(5225) <= not (a or b);
    layer0_outputs(5226) <= not a or b;
    layer0_outputs(5227) <= not b;
    layer0_outputs(5228) <= a;
    layer0_outputs(5229) <= b;
    layer0_outputs(5230) <= a or b;
    layer0_outputs(5231) <= not b or a;
    layer0_outputs(5232) <= a xor b;
    layer0_outputs(5233) <= b and not a;
    layer0_outputs(5234) <= a or b;
    layer0_outputs(5235) <= not b;
    layer0_outputs(5236) <= 1'b0;
    layer0_outputs(5237) <= a;
    layer0_outputs(5238) <= b;
    layer0_outputs(5239) <= a or b;
    layer0_outputs(5240) <= a;
    layer0_outputs(5241) <= not a;
    layer0_outputs(5242) <= a;
    layer0_outputs(5243) <= a;
    layer0_outputs(5244) <= not (a and b);
    layer0_outputs(5245) <= a;
    layer0_outputs(5246) <= not b or a;
    layer0_outputs(5247) <= not (a and b);
    layer0_outputs(5248) <= not (a xor b);
    layer0_outputs(5249) <= a xor b;
    layer0_outputs(5250) <= not b or a;
    layer0_outputs(5251) <= not a;
    layer0_outputs(5252) <= not b;
    layer0_outputs(5253) <= not (a or b);
    layer0_outputs(5254) <= b;
    layer0_outputs(5255) <= a xor b;
    layer0_outputs(5256) <= not (a and b);
    layer0_outputs(5257) <= not a;
    layer0_outputs(5258) <= not (a xor b);
    layer0_outputs(5259) <= a or b;
    layer0_outputs(5260) <= not (a and b);
    layer0_outputs(5261) <= b;
    layer0_outputs(5262) <= a;
    layer0_outputs(5263) <= not (a xor b);
    layer0_outputs(5264) <= b;
    layer0_outputs(5265) <= a xor b;
    layer0_outputs(5266) <= a and not b;
    layer0_outputs(5267) <= not b or a;
    layer0_outputs(5268) <= not a or b;
    layer0_outputs(5269) <= a and not b;
    layer0_outputs(5270) <= a and not b;
    layer0_outputs(5271) <= b and not a;
    layer0_outputs(5272) <= not b or a;
    layer0_outputs(5273) <= not (a xor b);
    layer0_outputs(5274) <= a or b;
    layer0_outputs(5275) <= not (a and b);
    layer0_outputs(5276) <= not b or a;
    layer0_outputs(5277) <= b and not a;
    layer0_outputs(5278) <= a or b;
    layer0_outputs(5279) <= b;
    layer0_outputs(5280) <= a and b;
    layer0_outputs(5281) <= a;
    layer0_outputs(5282) <= a;
    layer0_outputs(5283) <= not b;
    layer0_outputs(5284) <= not (a or b);
    layer0_outputs(5285) <= a or b;
    layer0_outputs(5286) <= b;
    layer0_outputs(5287) <= 1'b0;
    layer0_outputs(5288) <= a or b;
    layer0_outputs(5289) <= not b;
    layer0_outputs(5290) <= not b or a;
    layer0_outputs(5291) <= 1'b0;
    layer0_outputs(5292) <= b and not a;
    layer0_outputs(5293) <= not b or a;
    layer0_outputs(5294) <= not (a xor b);
    layer0_outputs(5295) <= 1'b0;
    layer0_outputs(5296) <= not (a or b);
    layer0_outputs(5297) <= not (a xor b);
    layer0_outputs(5298) <= b;
    layer0_outputs(5299) <= not (a xor b);
    layer0_outputs(5300) <= not (a xor b);
    layer0_outputs(5301) <= not b or a;
    layer0_outputs(5302) <= a;
    layer0_outputs(5303) <= b and not a;
    layer0_outputs(5304) <= a or b;
    layer0_outputs(5305) <= not (a or b);
    layer0_outputs(5306) <= a xor b;
    layer0_outputs(5307) <= a or b;
    layer0_outputs(5308) <= not a;
    layer0_outputs(5309) <= not (a or b);
    layer0_outputs(5310) <= 1'b1;
    layer0_outputs(5311) <= not a;
    layer0_outputs(5312) <= a xor b;
    layer0_outputs(5313) <= not (a or b);
    layer0_outputs(5314) <= not (a xor b);
    layer0_outputs(5315) <= a and not b;
    layer0_outputs(5316) <= a xor b;
    layer0_outputs(5317) <= a xor b;
    layer0_outputs(5318) <= not a;
    layer0_outputs(5319) <= not a or b;
    layer0_outputs(5320) <= not b;
    layer0_outputs(5321) <= a or b;
    layer0_outputs(5322) <= not a;
    layer0_outputs(5323) <= a or b;
    layer0_outputs(5324) <= a or b;
    layer0_outputs(5325) <= not a or b;
    layer0_outputs(5326) <= not a or b;
    layer0_outputs(5327) <= not (a xor b);
    layer0_outputs(5328) <= b;
    layer0_outputs(5329) <= not a;
    layer0_outputs(5330) <= b and not a;
    layer0_outputs(5331) <= a;
    layer0_outputs(5332) <= b;
    layer0_outputs(5333) <= a or b;
    layer0_outputs(5334) <= not (a xor b);
    layer0_outputs(5335) <= a;
    layer0_outputs(5336) <= a and not b;
    layer0_outputs(5337) <= a and not b;
    layer0_outputs(5338) <= not a;
    layer0_outputs(5339) <= b;
    layer0_outputs(5340) <= 1'b0;
    layer0_outputs(5341) <= not a or b;
    layer0_outputs(5342) <= not b or a;
    layer0_outputs(5343) <= not a or b;
    layer0_outputs(5344) <= not (a xor b);
    layer0_outputs(5345) <= not (a or b);
    layer0_outputs(5346) <= not (a xor b);
    layer0_outputs(5347) <= not (a or b);
    layer0_outputs(5348) <= not (a or b);
    layer0_outputs(5349) <= b;
    layer0_outputs(5350) <= not b;
    layer0_outputs(5351) <= not (a xor b);
    layer0_outputs(5352) <= not b or a;
    layer0_outputs(5353) <= a xor b;
    layer0_outputs(5354) <= 1'b1;
    layer0_outputs(5355) <= a or b;
    layer0_outputs(5356) <= a xor b;
    layer0_outputs(5357) <= a;
    layer0_outputs(5358) <= b;
    layer0_outputs(5359) <= a;
    layer0_outputs(5360) <= a;
    layer0_outputs(5361) <= 1'b0;
    layer0_outputs(5362) <= a and b;
    layer0_outputs(5363) <= a xor b;
    layer0_outputs(5364) <= a and not b;
    layer0_outputs(5365) <= a or b;
    layer0_outputs(5366) <= a and b;
    layer0_outputs(5367) <= a or b;
    layer0_outputs(5368) <= 1'b1;
    layer0_outputs(5369) <= not a or b;
    layer0_outputs(5370) <= b;
    layer0_outputs(5371) <= 1'b0;
    layer0_outputs(5372) <= a or b;
    layer0_outputs(5373) <= not a;
    layer0_outputs(5374) <= b;
    layer0_outputs(5375) <= not a or b;
    layer0_outputs(5376) <= b;
    layer0_outputs(5377) <= 1'b0;
    layer0_outputs(5378) <= not (a or b);
    layer0_outputs(5379) <= a xor b;
    layer0_outputs(5380) <= b and not a;
    layer0_outputs(5381) <= 1'b0;
    layer0_outputs(5382) <= not (a xor b);
    layer0_outputs(5383) <= not a;
    layer0_outputs(5384) <= b;
    layer0_outputs(5385) <= b and not a;
    layer0_outputs(5386) <= not (a and b);
    layer0_outputs(5387) <= not b;
    layer0_outputs(5388) <= not b;
    layer0_outputs(5389) <= not a;
    layer0_outputs(5390) <= not a or b;
    layer0_outputs(5391) <= b and not a;
    layer0_outputs(5392) <= not (a or b);
    layer0_outputs(5393) <= not (a and b);
    layer0_outputs(5394) <= not b or a;
    layer0_outputs(5395) <= not (a or b);
    layer0_outputs(5396) <= not b or a;
    layer0_outputs(5397) <= not a;
    layer0_outputs(5398) <= not (a or b);
    layer0_outputs(5399) <= not (a xor b);
    layer0_outputs(5400) <= a or b;
    layer0_outputs(5401) <= 1'b1;
    layer0_outputs(5402) <= not b;
    layer0_outputs(5403) <= not (a and b);
    layer0_outputs(5404) <= not b;
    layer0_outputs(5405) <= not b or a;
    layer0_outputs(5406) <= a or b;
    layer0_outputs(5407) <= not a;
    layer0_outputs(5408) <= a or b;
    layer0_outputs(5409) <= b and not a;
    layer0_outputs(5410) <= b;
    layer0_outputs(5411) <= a and b;
    layer0_outputs(5412) <= 1'b1;
    layer0_outputs(5413) <= a xor b;
    layer0_outputs(5414) <= not (a or b);
    layer0_outputs(5415) <= not b or a;
    layer0_outputs(5416) <= not b or a;
    layer0_outputs(5417) <= not a or b;
    layer0_outputs(5418) <= b and not a;
    layer0_outputs(5419) <= not a;
    layer0_outputs(5420) <= not (a xor b);
    layer0_outputs(5421) <= not b or a;
    layer0_outputs(5422) <= a xor b;
    layer0_outputs(5423) <= not b;
    layer0_outputs(5424) <= not a or b;
    layer0_outputs(5425) <= a or b;
    layer0_outputs(5426) <= not a or b;
    layer0_outputs(5427) <= not a;
    layer0_outputs(5428) <= not a;
    layer0_outputs(5429) <= a and not b;
    layer0_outputs(5430) <= not (a or b);
    layer0_outputs(5431) <= a or b;
    layer0_outputs(5432) <= a or b;
    layer0_outputs(5433) <= a xor b;
    layer0_outputs(5434) <= not a or b;
    layer0_outputs(5435) <= b;
    layer0_outputs(5436) <= not a or b;
    layer0_outputs(5437) <= b;
    layer0_outputs(5438) <= a and b;
    layer0_outputs(5439) <= not a or b;
    layer0_outputs(5440) <= a;
    layer0_outputs(5441) <= not (a xor b);
    layer0_outputs(5442) <= not b or a;
    layer0_outputs(5443) <= not (a or b);
    layer0_outputs(5444) <= not (a xor b);
    layer0_outputs(5445) <= not (a xor b);
    layer0_outputs(5446) <= 1'b0;
    layer0_outputs(5447) <= not b or a;
    layer0_outputs(5448) <= not (a and b);
    layer0_outputs(5449) <= 1'b0;
    layer0_outputs(5450) <= 1'b0;
    layer0_outputs(5451) <= not (a or b);
    layer0_outputs(5452) <= 1'b0;
    layer0_outputs(5453) <= a or b;
    layer0_outputs(5454) <= a xor b;
    layer0_outputs(5455) <= not b;
    layer0_outputs(5456) <= not (a or b);
    layer0_outputs(5457) <= not a or b;
    layer0_outputs(5458) <= not (a or b);
    layer0_outputs(5459) <= not (a or b);
    layer0_outputs(5460) <= not a;
    layer0_outputs(5461) <= a;
    layer0_outputs(5462) <= a;
    layer0_outputs(5463) <= not (a and b);
    layer0_outputs(5464) <= not a;
    layer0_outputs(5465) <= not a or b;
    layer0_outputs(5466) <= not (a or b);
    layer0_outputs(5467) <= not (a or b);
    layer0_outputs(5468) <= not (a or b);
    layer0_outputs(5469) <= 1'b1;
    layer0_outputs(5470) <= not (a or b);
    layer0_outputs(5471) <= a or b;
    layer0_outputs(5472) <= a and not b;
    layer0_outputs(5473) <= not (a and b);
    layer0_outputs(5474) <= a and b;
    layer0_outputs(5475) <= b;
    layer0_outputs(5476) <= not a or b;
    layer0_outputs(5477) <= not b;
    layer0_outputs(5478) <= a and not b;
    layer0_outputs(5479) <= not (a xor b);
    layer0_outputs(5480) <= not (a or b);
    layer0_outputs(5481) <= a;
    layer0_outputs(5482) <= not a or b;
    layer0_outputs(5483) <= not (a or b);
    layer0_outputs(5484) <= not b;
    layer0_outputs(5485) <= a;
    layer0_outputs(5486) <= not (a or b);
    layer0_outputs(5487) <= a or b;
    layer0_outputs(5488) <= b and not a;
    layer0_outputs(5489) <= not b or a;
    layer0_outputs(5490) <= not (a xor b);
    layer0_outputs(5491) <= not (a xor b);
    layer0_outputs(5492) <= not a or b;
    layer0_outputs(5493) <= not (a xor b);
    layer0_outputs(5494) <= 1'b0;
    layer0_outputs(5495) <= not a or b;
    layer0_outputs(5496) <= b and not a;
    layer0_outputs(5497) <= a or b;
    layer0_outputs(5498) <= a xor b;
    layer0_outputs(5499) <= b and not a;
    layer0_outputs(5500) <= a and not b;
    layer0_outputs(5501) <= not (a xor b);
    layer0_outputs(5502) <= a or b;
    layer0_outputs(5503) <= not b or a;
    layer0_outputs(5504) <= not a or b;
    layer0_outputs(5505) <= not a or b;
    layer0_outputs(5506) <= a or b;
    layer0_outputs(5507) <= not (a or b);
    layer0_outputs(5508) <= not (a and b);
    layer0_outputs(5509) <= a;
    layer0_outputs(5510) <= not b;
    layer0_outputs(5511) <= a and b;
    layer0_outputs(5512) <= b and not a;
    layer0_outputs(5513) <= 1'b0;
    layer0_outputs(5514) <= 1'b0;
    layer0_outputs(5515) <= a or b;
    layer0_outputs(5516) <= a or b;
    layer0_outputs(5517) <= a xor b;
    layer0_outputs(5518) <= a and not b;
    layer0_outputs(5519) <= not a or b;
    layer0_outputs(5520) <= not (a xor b);
    layer0_outputs(5521) <= a xor b;
    layer0_outputs(5522) <= not b;
    layer0_outputs(5523) <= a or b;
    layer0_outputs(5524) <= not (a xor b);
    layer0_outputs(5525) <= b;
    layer0_outputs(5526) <= a or b;
    layer0_outputs(5527) <= a or b;
    layer0_outputs(5528) <= not a;
    layer0_outputs(5529) <= a and not b;
    layer0_outputs(5530) <= not (a xor b);
    layer0_outputs(5531) <= a or b;
    layer0_outputs(5532) <= not b or a;
    layer0_outputs(5533) <= a or b;
    layer0_outputs(5534) <= not (a or b);
    layer0_outputs(5535) <= not (a or b);
    layer0_outputs(5536) <= b and not a;
    layer0_outputs(5537) <= b;
    layer0_outputs(5538) <= not (a xor b);
    layer0_outputs(5539) <= a and not b;
    layer0_outputs(5540) <= not (a and b);
    layer0_outputs(5541) <= not b or a;
    layer0_outputs(5542) <= not a;
    layer0_outputs(5543) <= a xor b;
    layer0_outputs(5544) <= not b;
    layer0_outputs(5545) <= b and not a;
    layer0_outputs(5546) <= a xor b;
    layer0_outputs(5547) <= b;
    layer0_outputs(5548) <= a and not b;
    layer0_outputs(5549) <= not a;
    layer0_outputs(5550) <= not (a xor b);
    layer0_outputs(5551) <= a xor b;
    layer0_outputs(5552) <= a and not b;
    layer0_outputs(5553) <= b;
    layer0_outputs(5554) <= a;
    layer0_outputs(5555) <= 1'b0;
    layer0_outputs(5556) <= not b or a;
    layer0_outputs(5557) <= a or b;
    layer0_outputs(5558) <= not (a xor b);
    layer0_outputs(5559) <= b and not a;
    layer0_outputs(5560) <= not (a xor b);
    layer0_outputs(5561) <= a and not b;
    layer0_outputs(5562) <= not (a or b);
    layer0_outputs(5563) <= not a;
    layer0_outputs(5564) <= b;
    layer0_outputs(5565) <= a;
    layer0_outputs(5566) <= not a or b;
    layer0_outputs(5567) <= b and not a;
    layer0_outputs(5568) <= 1'b1;
    layer0_outputs(5569) <= not b;
    layer0_outputs(5570) <= not a or b;
    layer0_outputs(5571) <= b;
    layer0_outputs(5572) <= not (a xor b);
    layer0_outputs(5573) <= a and b;
    layer0_outputs(5574) <= b and not a;
    layer0_outputs(5575) <= a xor b;
    layer0_outputs(5576) <= a and not b;
    layer0_outputs(5577) <= not b;
    layer0_outputs(5578) <= a or b;
    layer0_outputs(5579) <= not a;
    layer0_outputs(5580) <= not b or a;
    layer0_outputs(5581) <= a or b;
    layer0_outputs(5582) <= a;
    layer0_outputs(5583) <= a and not b;
    layer0_outputs(5584) <= a xor b;
    layer0_outputs(5585) <= 1'b0;
    layer0_outputs(5586) <= a xor b;
    layer0_outputs(5587) <= not a or b;
    layer0_outputs(5588) <= not a;
    layer0_outputs(5589) <= a or b;
    layer0_outputs(5590) <= not b;
    layer0_outputs(5591) <= not a;
    layer0_outputs(5592) <= b and not a;
    layer0_outputs(5593) <= not a;
    layer0_outputs(5594) <= a;
    layer0_outputs(5595) <= a or b;
    layer0_outputs(5596) <= b and not a;
    layer0_outputs(5597) <= a;
    layer0_outputs(5598) <= a or b;
    layer0_outputs(5599) <= a;
    layer0_outputs(5600) <= a;
    layer0_outputs(5601) <= not a;
    layer0_outputs(5602) <= not a;
    layer0_outputs(5603) <= not a;
    layer0_outputs(5604) <= a and not b;
    layer0_outputs(5605) <= b;
    layer0_outputs(5606) <= 1'b1;
    layer0_outputs(5607) <= a or b;
    layer0_outputs(5608) <= not a;
    layer0_outputs(5609) <= a or b;
    layer0_outputs(5610) <= not (a xor b);
    layer0_outputs(5611) <= not b;
    layer0_outputs(5612) <= a or b;
    layer0_outputs(5613) <= not b;
    layer0_outputs(5614) <= not (a xor b);
    layer0_outputs(5615) <= a and not b;
    layer0_outputs(5616) <= not (a xor b);
    layer0_outputs(5617) <= not a or b;
    layer0_outputs(5618) <= a and not b;
    layer0_outputs(5619) <= not (a or b);
    layer0_outputs(5620) <= not a;
    layer0_outputs(5621) <= a xor b;
    layer0_outputs(5622) <= a or b;
    layer0_outputs(5623) <= not (a xor b);
    layer0_outputs(5624) <= not (a or b);
    layer0_outputs(5625) <= 1'b1;
    layer0_outputs(5626) <= b;
    layer0_outputs(5627) <= b and not a;
    layer0_outputs(5628) <= not b or a;
    layer0_outputs(5629) <= not (a or b);
    layer0_outputs(5630) <= a xor b;
    layer0_outputs(5631) <= not a or b;
    layer0_outputs(5632) <= not a or b;
    layer0_outputs(5633) <= a;
    layer0_outputs(5634) <= not (a and b);
    layer0_outputs(5635) <= a or b;
    layer0_outputs(5636) <= b;
    layer0_outputs(5637) <= not (a xor b);
    layer0_outputs(5638) <= not (a xor b);
    layer0_outputs(5639) <= b and not a;
    layer0_outputs(5640) <= not (a or b);
    layer0_outputs(5641) <= 1'b1;
    layer0_outputs(5642) <= a and not b;
    layer0_outputs(5643) <= a and not b;
    layer0_outputs(5644) <= not (a xor b);
    layer0_outputs(5645) <= a xor b;
    layer0_outputs(5646) <= a xor b;
    layer0_outputs(5647) <= not (a or b);
    layer0_outputs(5648) <= a;
    layer0_outputs(5649) <= not a;
    layer0_outputs(5650) <= not (a or b);
    layer0_outputs(5651) <= not a or b;
    layer0_outputs(5652) <= not b;
    layer0_outputs(5653) <= not (a xor b);
    layer0_outputs(5654) <= a;
    layer0_outputs(5655) <= not b or a;
    layer0_outputs(5656) <= not b or a;
    layer0_outputs(5657) <= not (a xor b);
    layer0_outputs(5658) <= a and b;
    layer0_outputs(5659) <= a xor b;
    layer0_outputs(5660) <= b;
    layer0_outputs(5661) <= not a;
    layer0_outputs(5662) <= not (a xor b);
    layer0_outputs(5663) <= not a;
    layer0_outputs(5664) <= a or b;
    layer0_outputs(5665) <= not a;
    layer0_outputs(5666) <= b and not a;
    layer0_outputs(5667) <= a xor b;
    layer0_outputs(5668) <= not a;
    layer0_outputs(5669) <= 1'b0;
    layer0_outputs(5670) <= not (a xor b);
    layer0_outputs(5671) <= a or b;
    layer0_outputs(5672) <= not b or a;
    layer0_outputs(5673) <= a or b;
    layer0_outputs(5674) <= 1'b0;
    layer0_outputs(5675) <= a or b;
    layer0_outputs(5676) <= not (a xor b);
    layer0_outputs(5677) <= a;
    layer0_outputs(5678) <= not a or b;
    layer0_outputs(5679) <= b;
    layer0_outputs(5680) <= b and not a;
    layer0_outputs(5681) <= a xor b;
    layer0_outputs(5682) <= a xor b;
    layer0_outputs(5683) <= 1'b1;
    layer0_outputs(5684) <= a xor b;
    layer0_outputs(5685) <= a or b;
    layer0_outputs(5686) <= not b or a;
    layer0_outputs(5687) <= a or b;
    layer0_outputs(5688) <= not b or a;
    layer0_outputs(5689) <= not a or b;
    layer0_outputs(5690) <= not a or b;
    layer0_outputs(5691) <= not (a or b);
    layer0_outputs(5692) <= 1'b1;
    layer0_outputs(5693) <= not (a or b);
    layer0_outputs(5694) <= a and not b;
    layer0_outputs(5695) <= not (a or b);
    layer0_outputs(5696) <= a;
    layer0_outputs(5697) <= a or b;
    layer0_outputs(5698) <= b;
    layer0_outputs(5699) <= a xor b;
    layer0_outputs(5700) <= not b or a;
    layer0_outputs(5701) <= b and not a;
    layer0_outputs(5702) <= a or b;
    layer0_outputs(5703) <= not b;
    layer0_outputs(5704) <= not a or b;
    layer0_outputs(5705) <= a;
    layer0_outputs(5706) <= a or b;
    layer0_outputs(5707) <= a or b;
    layer0_outputs(5708) <= not (a xor b);
    layer0_outputs(5709) <= not (a or b);
    layer0_outputs(5710) <= not (a or b);
    layer0_outputs(5711) <= 1'b1;
    layer0_outputs(5712) <= a or b;
    layer0_outputs(5713) <= a xor b;
    layer0_outputs(5714) <= not (a or b);
    layer0_outputs(5715) <= not b or a;
    layer0_outputs(5716) <= a or b;
    layer0_outputs(5717) <= not (a or b);
    layer0_outputs(5718) <= b;
    layer0_outputs(5719) <= not (a or b);
    layer0_outputs(5720) <= a and not b;
    layer0_outputs(5721) <= not b or a;
    layer0_outputs(5722) <= not b;
    layer0_outputs(5723) <= a or b;
    layer0_outputs(5724) <= not b or a;
    layer0_outputs(5725) <= b;
    layer0_outputs(5726) <= not b;
    layer0_outputs(5727) <= not (a or b);
    layer0_outputs(5728) <= not b or a;
    layer0_outputs(5729) <= a;
    layer0_outputs(5730) <= not (a or b);
    layer0_outputs(5731) <= a xor b;
    layer0_outputs(5732) <= not b or a;
    layer0_outputs(5733) <= a or b;
    layer0_outputs(5734) <= 1'b0;
    layer0_outputs(5735) <= not b or a;
    layer0_outputs(5736) <= not (a or b);
    layer0_outputs(5737) <= a or b;
    layer0_outputs(5738) <= a xor b;
    layer0_outputs(5739) <= not (a xor b);
    layer0_outputs(5740) <= b;
    layer0_outputs(5741) <= a or b;
    layer0_outputs(5742) <= b and not a;
    layer0_outputs(5743) <= b;
    layer0_outputs(5744) <= b and not a;
    layer0_outputs(5745) <= a xor b;
    layer0_outputs(5746) <= not (a and b);
    layer0_outputs(5747) <= a or b;
    layer0_outputs(5748) <= a or b;
    layer0_outputs(5749) <= not b or a;
    layer0_outputs(5750) <= not (a or b);
    layer0_outputs(5751) <= b;
    layer0_outputs(5752) <= a and b;
    layer0_outputs(5753) <= b and not a;
    layer0_outputs(5754) <= not (a or b);
    layer0_outputs(5755) <= not (a xor b);
    layer0_outputs(5756) <= not b;
    layer0_outputs(5757) <= not b or a;
    layer0_outputs(5758) <= a or b;
    layer0_outputs(5759) <= b;
    layer0_outputs(5760) <= not a;
    layer0_outputs(5761) <= b and not a;
    layer0_outputs(5762) <= not (a or b);
    layer0_outputs(5763) <= a or b;
    layer0_outputs(5764) <= a and not b;
    layer0_outputs(5765) <= not a;
    layer0_outputs(5766) <= a or b;
    layer0_outputs(5767) <= b and not a;
    layer0_outputs(5768) <= a or b;
    layer0_outputs(5769) <= not b;
    layer0_outputs(5770) <= a or b;
    layer0_outputs(5771) <= a xor b;
    layer0_outputs(5772) <= not (a or b);
    layer0_outputs(5773) <= b;
    layer0_outputs(5774) <= not (a xor b);
    layer0_outputs(5775) <= not b or a;
    layer0_outputs(5776) <= a;
    layer0_outputs(5777) <= a or b;
    layer0_outputs(5778) <= a and b;
    layer0_outputs(5779) <= 1'b1;
    layer0_outputs(5780) <= not a;
    layer0_outputs(5781) <= b;
    layer0_outputs(5782) <= b and not a;
    layer0_outputs(5783) <= not a or b;
    layer0_outputs(5784) <= not (a xor b);
    layer0_outputs(5785) <= not (a or b);
    layer0_outputs(5786) <= a or b;
    layer0_outputs(5787) <= not b;
    layer0_outputs(5788) <= not (a or b);
    layer0_outputs(5789) <= not a;
    layer0_outputs(5790) <= not a;
    layer0_outputs(5791) <= not a;
    layer0_outputs(5792) <= 1'b0;
    layer0_outputs(5793) <= not b or a;
    layer0_outputs(5794) <= b;
    layer0_outputs(5795) <= a and not b;
    layer0_outputs(5796) <= b;
    layer0_outputs(5797) <= not (a and b);
    layer0_outputs(5798) <= a;
    layer0_outputs(5799) <= a or b;
    layer0_outputs(5800) <= a xor b;
    layer0_outputs(5801) <= not (a or b);
    layer0_outputs(5802) <= not a or b;
    layer0_outputs(5803) <= not (a or b);
    layer0_outputs(5804) <= not (a xor b);
    layer0_outputs(5805) <= not b or a;
    layer0_outputs(5806) <= b;
    layer0_outputs(5807) <= not b;
    layer0_outputs(5808) <= not (a and b);
    layer0_outputs(5809) <= not (a or b);
    layer0_outputs(5810) <= 1'b1;
    layer0_outputs(5811) <= not a or b;
    layer0_outputs(5812) <= b;
    layer0_outputs(5813) <= not a;
    layer0_outputs(5814) <= not b;
    layer0_outputs(5815) <= not b;
    layer0_outputs(5816) <= not a or b;
    layer0_outputs(5817) <= not a;
    layer0_outputs(5818) <= b;
    layer0_outputs(5819) <= b and not a;
    layer0_outputs(5820) <= not a;
    layer0_outputs(5821) <= not a;
    layer0_outputs(5822) <= a;
    layer0_outputs(5823) <= not (a xor b);
    layer0_outputs(5824) <= a and not b;
    layer0_outputs(5825) <= not (a or b);
    layer0_outputs(5826) <= 1'b1;
    layer0_outputs(5827) <= not a or b;
    layer0_outputs(5828) <= not a;
    layer0_outputs(5829) <= a and not b;
    layer0_outputs(5830) <= a xor b;
    layer0_outputs(5831) <= a xor b;
    layer0_outputs(5832) <= not a or b;
    layer0_outputs(5833) <= not (a or b);
    layer0_outputs(5834) <= not b;
    layer0_outputs(5835) <= not (a xor b);
    layer0_outputs(5836) <= 1'b1;
    layer0_outputs(5837) <= a or b;
    layer0_outputs(5838) <= 1'b1;
    layer0_outputs(5839) <= not a;
    layer0_outputs(5840) <= a or b;
    layer0_outputs(5841) <= not (a or b);
    layer0_outputs(5842) <= a;
    layer0_outputs(5843) <= not (a xor b);
    layer0_outputs(5844) <= a;
    layer0_outputs(5845) <= a xor b;
    layer0_outputs(5846) <= not b;
    layer0_outputs(5847) <= a and b;
    layer0_outputs(5848) <= a or b;
    layer0_outputs(5849) <= not a or b;
    layer0_outputs(5850) <= not (a xor b);
    layer0_outputs(5851) <= not a or b;
    layer0_outputs(5852) <= b;
    layer0_outputs(5853) <= a or b;
    layer0_outputs(5854) <= b and not a;
    layer0_outputs(5855) <= not (a or b);
    layer0_outputs(5856) <= not b;
    layer0_outputs(5857) <= 1'b1;
    layer0_outputs(5858) <= not (a xor b);
    layer0_outputs(5859) <= not b or a;
    layer0_outputs(5860) <= not a or b;
    layer0_outputs(5861) <= not a or b;
    layer0_outputs(5862) <= b;
    layer0_outputs(5863) <= 1'b1;
    layer0_outputs(5864) <= a;
    layer0_outputs(5865) <= b;
    layer0_outputs(5866) <= not a;
    layer0_outputs(5867) <= a xor b;
    layer0_outputs(5868) <= a and not b;
    layer0_outputs(5869) <= a xor b;
    layer0_outputs(5870) <= not a or b;
    layer0_outputs(5871) <= a xor b;
    layer0_outputs(5872) <= not b;
    layer0_outputs(5873) <= a;
    layer0_outputs(5874) <= not b or a;
    layer0_outputs(5875) <= a or b;
    layer0_outputs(5876) <= not (a or b);
    layer0_outputs(5877) <= a or b;
    layer0_outputs(5878) <= not b or a;
    layer0_outputs(5879) <= not a;
    layer0_outputs(5880) <= not (a xor b);
    layer0_outputs(5881) <= not (a or b);
    layer0_outputs(5882) <= b;
    layer0_outputs(5883) <= 1'b0;
    layer0_outputs(5884) <= not a;
    layer0_outputs(5885) <= 1'b0;
    layer0_outputs(5886) <= not b;
    layer0_outputs(5887) <= b;
    layer0_outputs(5888) <= not a or b;
    layer0_outputs(5889) <= not (a or b);
    layer0_outputs(5890) <= not (a xor b);
    layer0_outputs(5891) <= not b or a;
    layer0_outputs(5892) <= not (a xor b);
    layer0_outputs(5893) <= a and not b;
    layer0_outputs(5894) <= a or b;
    layer0_outputs(5895) <= not b;
    layer0_outputs(5896) <= a xor b;
    layer0_outputs(5897) <= not a or b;
    layer0_outputs(5898) <= a or b;
    layer0_outputs(5899) <= not (a or b);
    layer0_outputs(5900) <= a and not b;
    layer0_outputs(5901) <= not (a xor b);
    layer0_outputs(5902) <= not (a or b);
    layer0_outputs(5903) <= a xor b;
    layer0_outputs(5904) <= not a;
    layer0_outputs(5905) <= b and not a;
    layer0_outputs(5906) <= not a;
    layer0_outputs(5907) <= a xor b;
    layer0_outputs(5908) <= a or b;
    layer0_outputs(5909) <= not b;
    layer0_outputs(5910) <= a and not b;
    layer0_outputs(5911) <= not b;
    layer0_outputs(5912) <= b and not a;
    layer0_outputs(5913) <= not b or a;
    layer0_outputs(5914) <= a;
    layer0_outputs(5915) <= not (a xor b);
    layer0_outputs(5916) <= not a or b;
    layer0_outputs(5917) <= not (a or b);
    layer0_outputs(5918) <= not (a xor b);
    layer0_outputs(5919) <= not (a xor b);
    layer0_outputs(5920) <= 1'b1;
    layer0_outputs(5921) <= not (a or b);
    layer0_outputs(5922) <= not a or b;
    layer0_outputs(5923) <= 1'b1;
    layer0_outputs(5924) <= not (a xor b);
    layer0_outputs(5925) <= not b or a;
    layer0_outputs(5926) <= not a;
    layer0_outputs(5927) <= a;
    layer0_outputs(5928) <= not b or a;
    layer0_outputs(5929) <= b and not a;
    layer0_outputs(5930) <= a and not b;
    layer0_outputs(5931) <= 1'b1;
    layer0_outputs(5932) <= not (a xor b);
    layer0_outputs(5933) <= not b;
    layer0_outputs(5934) <= a or b;
    layer0_outputs(5935) <= b;
    layer0_outputs(5936) <= a and not b;
    layer0_outputs(5937) <= a;
    layer0_outputs(5938) <= not (a or b);
    layer0_outputs(5939) <= not (a or b);
    layer0_outputs(5940) <= not (a xor b);
    layer0_outputs(5941) <= not (a or b);
    layer0_outputs(5942) <= a and b;
    layer0_outputs(5943) <= a or b;
    layer0_outputs(5944) <= a;
    layer0_outputs(5945) <= 1'b0;
    layer0_outputs(5946) <= not (a and b);
    layer0_outputs(5947) <= not (a or b);
    layer0_outputs(5948) <= not a;
    layer0_outputs(5949) <= not a;
    layer0_outputs(5950) <= a or b;
    layer0_outputs(5951) <= a xor b;
    layer0_outputs(5952) <= a and b;
    layer0_outputs(5953) <= a or b;
    layer0_outputs(5954) <= a or b;
    layer0_outputs(5955) <= not (a or b);
    layer0_outputs(5956) <= not (a xor b);
    layer0_outputs(5957) <= not a or b;
    layer0_outputs(5958) <= not b or a;
    layer0_outputs(5959) <= b;
    layer0_outputs(5960) <= a xor b;
    layer0_outputs(5961) <= not a;
    layer0_outputs(5962) <= not (a and b);
    layer0_outputs(5963) <= a and not b;
    layer0_outputs(5964) <= a xor b;
    layer0_outputs(5965) <= a and b;
    layer0_outputs(5966) <= not (a and b);
    layer0_outputs(5967) <= not (a or b);
    layer0_outputs(5968) <= not a or b;
    layer0_outputs(5969) <= 1'b0;
    layer0_outputs(5970) <= a xor b;
    layer0_outputs(5971) <= a or b;
    layer0_outputs(5972) <= a xor b;
    layer0_outputs(5973) <= not b;
    layer0_outputs(5974) <= b;
    layer0_outputs(5975) <= not (a or b);
    layer0_outputs(5976) <= not a;
    layer0_outputs(5977) <= not (a xor b);
    layer0_outputs(5978) <= not a;
    layer0_outputs(5979) <= not b;
    layer0_outputs(5980) <= not a or b;
    layer0_outputs(5981) <= a and not b;
    layer0_outputs(5982) <= b;
    layer0_outputs(5983) <= a and not b;
    layer0_outputs(5984) <= a;
    layer0_outputs(5985) <= not a;
    layer0_outputs(5986) <= a xor b;
    layer0_outputs(5987) <= not a or b;
    layer0_outputs(5988) <= 1'b1;
    layer0_outputs(5989) <= a or b;
    layer0_outputs(5990) <= a and b;
    layer0_outputs(5991) <= not (a and b);
    layer0_outputs(5992) <= not (a or b);
    layer0_outputs(5993) <= not (a or b);
    layer0_outputs(5994) <= a xor b;
    layer0_outputs(5995) <= a;
    layer0_outputs(5996) <= 1'b0;
    layer0_outputs(5997) <= not (a or b);
    layer0_outputs(5998) <= 1'b0;
    layer0_outputs(5999) <= a and not b;
    layer0_outputs(6000) <= b;
    layer0_outputs(6001) <= a or b;
    layer0_outputs(6002) <= not (a and b);
    layer0_outputs(6003) <= not a;
    layer0_outputs(6004) <= not b;
    layer0_outputs(6005) <= not b;
    layer0_outputs(6006) <= not (a and b);
    layer0_outputs(6007) <= not (a or b);
    layer0_outputs(6008) <= a and not b;
    layer0_outputs(6009) <= b;
    layer0_outputs(6010) <= not a;
    layer0_outputs(6011) <= a and not b;
    layer0_outputs(6012) <= not (a or b);
    layer0_outputs(6013) <= a or b;
    layer0_outputs(6014) <= b;
    layer0_outputs(6015) <= a and not b;
    layer0_outputs(6016) <= b and not a;
    layer0_outputs(6017) <= not a or b;
    layer0_outputs(6018) <= not a;
    layer0_outputs(6019) <= a and b;
    layer0_outputs(6020) <= a and b;
    layer0_outputs(6021) <= not (a or b);
    layer0_outputs(6022) <= a xor b;
    layer0_outputs(6023) <= a and not b;
    layer0_outputs(6024) <= a and not b;
    layer0_outputs(6025) <= a or b;
    layer0_outputs(6026) <= not a or b;
    layer0_outputs(6027) <= b;
    layer0_outputs(6028) <= not b or a;
    layer0_outputs(6029) <= not (a or b);
    layer0_outputs(6030) <= a or b;
    layer0_outputs(6031) <= a or b;
    layer0_outputs(6032) <= not b or a;
    layer0_outputs(6033) <= not b;
    layer0_outputs(6034) <= not a or b;
    layer0_outputs(6035) <= not (a xor b);
    layer0_outputs(6036) <= a and not b;
    layer0_outputs(6037) <= not a;
    layer0_outputs(6038) <= not b;
    layer0_outputs(6039) <= not b;
    layer0_outputs(6040) <= a and b;
    layer0_outputs(6041) <= not (a xor b);
    layer0_outputs(6042) <= not b or a;
    layer0_outputs(6043) <= not b or a;
    layer0_outputs(6044) <= not (a or b);
    layer0_outputs(6045) <= 1'b0;
    layer0_outputs(6046) <= a and not b;
    layer0_outputs(6047) <= b;
    layer0_outputs(6048) <= not (a xor b);
    layer0_outputs(6049) <= not b or a;
    layer0_outputs(6050) <= not (a xor b);
    layer0_outputs(6051) <= a xor b;
    layer0_outputs(6052) <= not b;
    layer0_outputs(6053) <= b;
    layer0_outputs(6054) <= a and not b;
    layer0_outputs(6055) <= not (a xor b);
    layer0_outputs(6056) <= b and not a;
    layer0_outputs(6057) <= not a or b;
    layer0_outputs(6058) <= not (a or b);
    layer0_outputs(6059) <= a;
    layer0_outputs(6060) <= not b;
    layer0_outputs(6061) <= b and not a;
    layer0_outputs(6062) <= a xor b;
    layer0_outputs(6063) <= not b or a;
    layer0_outputs(6064) <= a xor b;
    layer0_outputs(6065) <= b;
    layer0_outputs(6066) <= not (a or b);
    layer0_outputs(6067) <= b;
    layer0_outputs(6068) <= a and not b;
    layer0_outputs(6069) <= b;
    layer0_outputs(6070) <= a or b;
    layer0_outputs(6071) <= 1'b1;
    layer0_outputs(6072) <= not (a xor b);
    layer0_outputs(6073) <= not (a xor b);
    layer0_outputs(6074) <= b and not a;
    layer0_outputs(6075) <= a and not b;
    layer0_outputs(6076) <= a or b;
    layer0_outputs(6077) <= a;
    layer0_outputs(6078) <= not (a xor b);
    layer0_outputs(6079) <= a;
    layer0_outputs(6080) <= not b;
    layer0_outputs(6081) <= not (a or b);
    layer0_outputs(6082) <= 1'b1;
    layer0_outputs(6083) <= 1'b1;
    layer0_outputs(6084) <= a xor b;
    layer0_outputs(6085) <= 1'b1;
    layer0_outputs(6086) <= b and not a;
    layer0_outputs(6087) <= not b;
    layer0_outputs(6088) <= not a;
    layer0_outputs(6089) <= b;
    layer0_outputs(6090) <= a and b;
    layer0_outputs(6091) <= a;
    layer0_outputs(6092) <= a xor b;
    layer0_outputs(6093) <= a xor b;
    layer0_outputs(6094) <= not a;
    layer0_outputs(6095) <= a;
    layer0_outputs(6096) <= a or b;
    layer0_outputs(6097) <= not a or b;
    layer0_outputs(6098) <= b and not a;
    layer0_outputs(6099) <= b and not a;
    layer0_outputs(6100) <= 1'b1;
    layer0_outputs(6101) <= 1'b1;
    layer0_outputs(6102) <= b and not a;
    layer0_outputs(6103) <= a xor b;
    layer0_outputs(6104) <= a or b;
    layer0_outputs(6105) <= not a or b;
    layer0_outputs(6106) <= a;
    layer0_outputs(6107) <= not (a and b);
    layer0_outputs(6108) <= a or b;
    layer0_outputs(6109) <= not (a xor b);
    layer0_outputs(6110) <= not (a xor b);
    layer0_outputs(6111) <= a xor b;
    layer0_outputs(6112) <= not b;
    layer0_outputs(6113) <= b;
    layer0_outputs(6114) <= a or b;
    layer0_outputs(6115) <= a or b;
    layer0_outputs(6116) <= not b or a;
    layer0_outputs(6117) <= b;
    layer0_outputs(6118) <= a or b;
    layer0_outputs(6119) <= b;
    layer0_outputs(6120) <= b and not a;
    layer0_outputs(6121) <= not b;
    layer0_outputs(6122) <= not (a or b);
    layer0_outputs(6123) <= a;
    layer0_outputs(6124) <= not (a xor b);
    layer0_outputs(6125) <= a and b;
    layer0_outputs(6126) <= b and not a;
    layer0_outputs(6127) <= b and not a;
    layer0_outputs(6128) <= a xor b;
    layer0_outputs(6129) <= a or b;
    layer0_outputs(6130) <= not (a xor b);
    layer0_outputs(6131) <= a or b;
    layer0_outputs(6132) <= not a;
    layer0_outputs(6133) <= 1'b1;
    layer0_outputs(6134) <= not (a or b);
    layer0_outputs(6135) <= b;
    layer0_outputs(6136) <= not a;
    layer0_outputs(6137) <= a xor b;
    layer0_outputs(6138) <= a or b;
    layer0_outputs(6139) <= not b or a;
    layer0_outputs(6140) <= b;
    layer0_outputs(6141) <= not a;
    layer0_outputs(6142) <= not (a or b);
    layer0_outputs(6143) <= not b;
    layer0_outputs(6144) <= a or b;
    layer0_outputs(6145) <= a;
    layer0_outputs(6146) <= not a;
    layer0_outputs(6147) <= a xor b;
    layer0_outputs(6148) <= a and not b;
    layer0_outputs(6149) <= a;
    layer0_outputs(6150) <= not (a or b);
    layer0_outputs(6151) <= a or b;
    layer0_outputs(6152) <= a;
    layer0_outputs(6153) <= a or b;
    layer0_outputs(6154) <= a;
    layer0_outputs(6155) <= a or b;
    layer0_outputs(6156) <= 1'b0;
    layer0_outputs(6157) <= a or b;
    layer0_outputs(6158) <= not (a xor b);
    layer0_outputs(6159) <= not (a xor b);
    layer0_outputs(6160) <= b;
    layer0_outputs(6161) <= a or b;
    layer0_outputs(6162) <= a or b;
    layer0_outputs(6163) <= not a;
    layer0_outputs(6164) <= not a or b;
    layer0_outputs(6165) <= not (a or b);
    layer0_outputs(6166) <= not (a xor b);
    layer0_outputs(6167) <= not b or a;
    layer0_outputs(6168) <= b and not a;
    layer0_outputs(6169) <= not (a or b);
    layer0_outputs(6170) <= not (a or b);
    layer0_outputs(6171) <= not (a xor b);
    layer0_outputs(6172) <= not (a xor b);
    layer0_outputs(6173) <= a xor b;
    layer0_outputs(6174) <= b;
    layer0_outputs(6175) <= b;
    layer0_outputs(6176) <= not b;
    layer0_outputs(6177) <= not (a and b);
    layer0_outputs(6178) <= not b or a;
    layer0_outputs(6179) <= not b or a;
    layer0_outputs(6180) <= not a or b;
    layer0_outputs(6181) <= a xor b;
    layer0_outputs(6182) <= not a or b;
    layer0_outputs(6183) <= a xor b;
    layer0_outputs(6184) <= a xor b;
    layer0_outputs(6185) <= not (a or b);
    layer0_outputs(6186) <= a or b;
    layer0_outputs(6187) <= not a or b;
    layer0_outputs(6188) <= not (a xor b);
    layer0_outputs(6189) <= not a or b;
    layer0_outputs(6190) <= not b;
    layer0_outputs(6191) <= b and not a;
    layer0_outputs(6192) <= not (a or b);
    layer0_outputs(6193) <= a xor b;
    layer0_outputs(6194) <= not a;
    layer0_outputs(6195) <= not a or b;
    layer0_outputs(6196) <= a xor b;
    layer0_outputs(6197) <= not b or a;
    layer0_outputs(6198) <= a and not b;
    layer0_outputs(6199) <= not (a xor b);
    layer0_outputs(6200) <= 1'b1;
    layer0_outputs(6201) <= a or b;
    layer0_outputs(6202) <= b;
    layer0_outputs(6203) <= not (a xor b);
    layer0_outputs(6204) <= a and not b;
    layer0_outputs(6205) <= not b or a;
    layer0_outputs(6206) <= not (a xor b);
    layer0_outputs(6207) <= not b;
    layer0_outputs(6208) <= a;
    layer0_outputs(6209) <= not a or b;
    layer0_outputs(6210) <= 1'b0;
    layer0_outputs(6211) <= 1'b0;
    layer0_outputs(6212) <= a xor b;
    layer0_outputs(6213) <= not (a or b);
    layer0_outputs(6214) <= a;
    layer0_outputs(6215) <= a xor b;
    layer0_outputs(6216) <= not b;
    layer0_outputs(6217) <= b and not a;
    layer0_outputs(6218) <= a xor b;
    layer0_outputs(6219) <= a and not b;
    layer0_outputs(6220) <= not a;
    layer0_outputs(6221) <= a and b;
    layer0_outputs(6222) <= not a;
    layer0_outputs(6223) <= not b or a;
    layer0_outputs(6224) <= b and not a;
    layer0_outputs(6225) <= a xor b;
    layer0_outputs(6226) <= a or b;
    layer0_outputs(6227) <= not a;
    layer0_outputs(6228) <= not (a or b);
    layer0_outputs(6229) <= not b;
    layer0_outputs(6230) <= not (a or b);
    layer0_outputs(6231) <= a or b;
    layer0_outputs(6232) <= a and not b;
    layer0_outputs(6233) <= a;
    layer0_outputs(6234) <= a or b;
    layer0_outputs(6235) <= not (a or b);
    layer0_outputs(6236) <= not a;
    layer0_outputs(6237) <= not (a or b);
    layer0_outputs(6238) <= a and b;
    layer0_outputs(6239) <= not (a or b);
    layer0_outputs(6240) <= not (a or b);
    layer0_outputs(6241) <= a xor b;
    layer0_outputs(6242) <= not b or a;
    layer0_outputs(6243) <= a and not b;
    layer0_outputs(6244) <= not a;
    layer0_outputs(6245) <= a;
    layer0_outputs(6246) <= not (a or b);
    layer0_outputs(6247) <= not (a xor b);
    layer0_outputs(6248) <= not a or b;
    layer0_outputs(6249) <= a or b;
    layer0_outputs(6250) <= not b or a;
    layer0_outputs(6251) <= not (a xor b);
    layer0_outputs(6252) <= not b;
    layer0_outputs(6253) <= a and not b;
    layer0_outputs(6254) <= not a;
    layer0_outputs(6255) <= a and not b;
    layer0_outputs(6256) <= not a or b;
    layer0_outputs(6257) <= not (a or b);
    layer0_outputs(6258) <= b and not a;
    layer0_outputs(6259) <= not a or b;
    layer0_outputs(6260) <= a and not b;
    layer0_outputs(6261) <= a xor b;
    layer0_outputs(6262) <= b and not a;
    layer0_outputs(6263) <= a xor b;
    layer0_outputs(6264) <= not (a or b);
    layer0_outputs(6265) <= not a;
    layer0_outputs(6266) <= a and not b;
    layer0_outputs(6267) <= b;
    layer0_outputs(6268) <= not b or a;
    layer0_outputs(6269) <= not b or a;
    layer0_outputs(6270) <= not b or a;
    layer0_outputs(6271) <= not (a xor b);
    layer0_outputs(6272) <= not b;
    layer0_outputs(6273) <= a;
    layer0_outputs(6274) <= a;
    layer0_outputs(6275) <= b;
    layer0_outputs(6276) <= a or b;
    layer0_outputs(6277) <= a or b;
    layer0_outputs(6278) <= a xor b;
    layer0_outputs(6279) <= a;
    layer0_outputs(6280) <= a or b;
    layer0_outputs(6281) <= a;
    layer0_outputs(6282) <= a xor b;
    layer0_outputs(6283) <= b;
    layer0_outputs(6284) <= a;
    layer0_outputs(6285) <= not b;
    layer0_outputs(6286) <= b;
    layer0_outputs(6287) <= not (a or b);
    layer0_outputs(6288) <= a xor b;
    layer0_outputs(6289) <= 1'b0;
    layer0_outputs(6290) <= 1'b0;
    layer0_outputs(6291) <= not (a or b);
    layer0_outputs(6292) <= a or b;
    layer0_outputs(6293) <= b and not a;
    layer0_outputs(6294) <= not a or b;
    layer0_outputs(6295) <= not (a xor b);
    layer0_outputs(6296) <= not b or a;
    layer0_outputs(6297) <= not (a or b);
    layer0_outputs(6298) <= a;
    layer0_outputs(6299) <= not b or a;
    layer0_outputs(6300) <= not b;
    layer0_outputs(6301) <= not (a or b);
    layer0_outputs(6302) <= b;
    layer0_outputs(6303) <= not (a and b);
    layer0_outputs(6304) <= a or b;
    layer0_outputs(6305) <= not (a xor b);
    layer0_outputs(6306) <= a;
    layer0_outputs(6307) <= not (a or b);
    layer0_outputs(6308) <= not a;
    layer0_outputs(6309) <= a and b;
    layer0_outputs(6310) <= a or b;
    layer0_outputs(6311) <= a or b;
    layer0_outputs(6312) <= b and not a;
    layer0_outputs(6313) <= 1'b1;
    layer0_outputs(6314) <= b;
    layer0_outputs(6315) <= not (a and b);
    layer0_outputs(6316) <= b;
    layer0_outputs(6317) <= b and not a;
    layer0_outputs(6318) <= not a;
    layer0_outputs(6319) <= a or b;
    layer0_outputs(6320) <= a or b;
    layer0_outputs(6321) <= b;
    layer0_outputs(6322) <= not (a or b);
    layer0_outputs(6323) <= 1'b1;
    layer0_outputs(6324) <= not (a or b);
    layer0_outputs(6325) <= a;
    layer0_outputs(6326) <= not a;
    layer0_outputs(6327) <= not (a xor b);
    layer0_outputs(6328) <= not (a or b);
    layer0_outputs(6329) <= not (a or b);
    layer0_outputs(6330) <= a and not b;
    layer0_outputs(6331) <= not b or a;
    layer0_outputs(6332) <= a or b;
    layer0_outputs(6333) <= a;
    layer0_outputs(6334) <= not b;
    layer0_outputs(6335) <= a xor b;
    layer0_outputs(6336) <= not a;
    layer0_outputs(6337) <= a xor b;
    layer0_outputs(6338) <= not a;
    layer0_outputs(6339) <= not a;
    layer0_outputs(6340) <= not b;
    layer0_outputs(6341) <= not a;
    layer0_outputs(6342) <= b and not a;
    layer0_outputs(6343) <= not (a xor b);
    layer0_outputs(6344) <= a xor b;
    layer0_outputs(6345) <= not a;
    layer0_outputs(6346) <= not (a or b);
    layer0_outputs(6347) <= not a or b;
    layer0_outputs(6348) <= 1'b1;
    layer0_outputs(6349) <= not a;
    layer0_outputs(6350) <= 1'b0;
    layer0_outputs(6351) <= 1'b0;
    layer0_outputs(6352) <= not b or a;
    layer0_outputs(6353) <= b;
    layer0_outputs(6354) <= not (a xor b);
    layer0_outputs(6355) <= a xor b;
    layer0_outputs(6356) <= b and not a;
    layer0_outputs(6357) <= a or b;
    layer0_outputs(6358) <= a or b;
    layer0_outputs(6359) <= a xor b;
    layer0_outputs(6360) <= not b;
    layer0_outputs(6361) <= b;
    layer0_outputs(6362) <= a xor b;
    layer0_outputs(6363) <= b;
    layer0_outputs(6364) <= a or b;
    layer0_outputs(6365) <= not (a xor b);
    layer0_outputs(6366) <= not (a xor b);
    layer0_outputs(6367) <= not a or b;
    layer0_outputs(6368) <= b;
    layer0_outputs(6369) <= not (a or b);
    layer0_outputs(6370) <= not a or b;
    layer0_outputs(6371) <= not b or a;
    layer0_outputs(6372) <= not (a or b);
    layer0_outputs(6373) <= a or b;
    layer0_outputs(6374) <= a or b;
    layer0_outputs(6375) <= b;
    layer0_outputs(6376) <= not b or a;
    layer0_outputs(6377) <= a;
    layer0_outputs(6378) <= b;
    layer0_outputs(6379) <= a or b;
    layer0_outputs(6380) <= a or b;
    layer0_outputs(6381) <= a and b;
    layer0_outputs(6382) <= a and not b;
    layer0_outputs(6383) <= a xor b;
    layer0_outputs(6384) <= not b;
    layer0_outputs(6385) <= a and not b;
    layer0_outputs(6386) <= not (a and b);
    layer0_outputs(6387) <= not b;
    layer0_outputs(6388) <= not (a or b);
    layer0_outputs(6389) <= not a;
    layer0_outputs(6390) <= b;
    layer0_outputs(6391) <= a or b;
    layer0_outputs(6392) <= not (a and b);
    layer0_outputs(6393) <= a xor b;
    layer0_outputs(6394) <= a;
    layer0_outputs(6395) <= not b;
    layer0_outputs(6396) <= a and not b;
    layer0_outputs(6397) <= a or b;
    layer0_outputs(6398) <= not b or a;
    layer0_outputs(6399) <= not b;
    layer0_outputs(6400) <= a;
    layer0_outputs(6401) <= a and b;
    layer0_outputs(6402) <= not a or b;
    layer0_outputs(6403) <= b;
    layer0_outputs(6404) <= b and not a;
    layer0_outputs(6405) <= a or b;
    layer0_outputs(6406) <= a xor b;
    layer0_outputs(6407) <= a and b;
    layer0_outputs(6408) <= not a or b;
    layer0_outputs(6409) <= 1'b0;
    layer0_outputs(6410) <= not b;
    layer0_outputs(6411) <= not b or a;
    layer0_outputs(6412) <= a or b;
    layer0_outputs(6413) <= a;
    layer0_outputs(6414) <= a xor b;
    layer0_outputs(6415) <= not a;
    layer0_outputs(6416) <= not (a or b);
    layer0_outputs(6417) <= a or b;
    layer0_outputs(6418) <= not a or b;
    layer0_outputs(6419) <= not a or b;
    layer0_outputs(6420) <= not b or a;
    layer0_outputs(6421) <= not (a and b);
    layer0_outputs(6422) <= not (a or b);
    layer0_outputs(6423) <= b;
    layer0_outputs(6424) <= b and not a;
    layer0_outputs(6425) <= not (a xor b);
    layer0_outputs(6426) <= not (a xor b);
    layer0_outputs(6427) <= b and not a;
    layer0_outputs(6428) <= 1'b1;
    layer0_outputs(6429) <= not b;
    layer0_outputs(6430) <= a and not b;
    layer0_outputs(6431) <= b and not a;
    layer0_outputs(6432) <= not (a or b);
    layer0_outputs(6433) <= not (a or b);
    layer0_outputs(6434) <= a xor b;
    layer0_outputs(6435) <= not (a or b);
    layer0_outputs(6436) <= 1'b0;
    layer0_outputs(6437) <= a;
    layer0_outputs(6438) <= not (a and b);
    layer0_outputs(6439) <= 1'b1;
    layer0_outputs(6440) <= not b or a;
    layer0_outputs(6441) <= b;
    layer0_outputs(6442) <= a;
    layer0_outputs(6443) <= 1'b0;
    layer0_outputs(6444) <= b and not a;
    layer0_outputs(6445) <= a xor b;
    layer0_outputs(6446) <= not b;
    layer0_outputs(6447) <= b;
    layer0_outputs(6448) <= not a;
    layer0_outputs(6449) <= not b;
    layer0_outputs(6450) <= not b;
    layer0_outputs(6451) <= a;
    layer0_outputs(6452) <= b;
    layer0_outputs(6453) <= 1'b1;
    layer0_outputs(6454) <= a and b;
    layer0_outputs(6455) <= a xor b;
    layer0_outputs(6456) <= not b;
    layer0_outputs(6457) <= not (a and b);
    layer0_outputs(6458) <= a and not b;
    layer0_outputs(6459) <= not (a xor b);
    layer0_outputs(6460) <= not (a and b);
    layer0_outputs(6461) <= not b;
    layer0_outputs(6462) <= a or b;
    layer0_outputs(6463) <= b;
    layer0_outputs(6464) <= a and not b;
    layer0_outputs(6465) <= a xor b;
    layer0_outputs(6466) <= a;
    layer0_outputs(6467) <= not (a or b);
    layer0_outputs(6468) <= not (a xor b);
    layer0_outputs(6469) <= b;
    layer0_outputs(6470) <= a;
    layer0_outputs(6471) <= not b or a;
    layer0_outputs(6472) <= b;
    layer0_outputs(6473) <= a xor b;
    layer0_outputs(6474) <= b;
    layer0_outputs(6475) <= not a or b;
    layer0_outputs(6476) <= a or b;
    layer0_outputs(6477) <= b;
    layer0_outputs(6478) <= a and not b;
    layer0_outputs(6479) <= a;
    layer0_outputs(6480) <= not b;
    layer0_outputs(6481) <= not a or b;
    layer0_outputs(6482) <= a or b;
    layer0_outputs(6483) <= not (a xor b);
    layer0_outputs(6484) <= a;
    layer0_outputs(6485) <= not a;
    layer0_outputs(6486) <= a and not b;
    layer0_outputs(6487) <= not (a or b);
    layer0_outputs(6488) <= not (a xor b);
    layer0_outputs(6489) <= a or b;
    layer0_outputs(6490) <= a;
    layer0_outputs(6491) <= a xor b;
    layer0_outputs(6492) <= a and not b;
    layer0_outputs(6493) <= a;
    layer0_outputs(6494) <= not (a or b);
    layer0_outputs(6495) <= not (a and b);
    layer0_outputs(6496) <= b;
    layer0_outputs(6497) <= a or b;
    layer0_outputs(6498) <= not b;
    layer0_outputs(6499) <= a;
    layer0_outputs(6500) <= not (a and b);
    layer0_outputs(6501) <= a xor b;
    layer0_outputs(6502) <= 1'b1;
    layer0_outputs(6503) <= not (a or b);
    layer0_outputs(6504) <= b;
    layer0_outputs(6505) <= b;
    layer0_outputs(6506) <= not (a or b);
    layer0_outputs(6507) <= a and b;
    layer0_outputs(6508) <= b;
    layer0_outputs(6509) <= not a;
    layer0_outputs(6510) <= not (a or b);
    layer0_outputs(6511) <= not a or b;
    layer0_outputs(6512) <= not a or b;
    layer0_outputs(6513) <= a;
    layer0_outputs(6514) <= b;
    layer0_outputs(6515) <= not (a and b);
    layer0_outputs(6516) <= a xor b;
    layer0_outputs(6517) <= not a;
    layer0_outputs(6518) <= not a or b;
    layer0_outputs(6519) <= a or b;
    layer0_outputs(6520) <= not (a and b);
    layer0_outputs(6521) <= not (a xor b);
    layer0_outputs(6522) <= not b;
    layer0_outputs(6523) <= not b or a;
    layer0_outputs(6524) <= b and not a;
    layer0_outputs(6525) <= a;
    layer0_outputs(6526) <= not a;
    layer0_outputs(6527) <= not (a or b);
    layer0_outputs(6528) <= a and not b;
    layer0_outputs(6529) <= not (a xor b);
    layer0_outputs(6530) <= not (a xor b);
    layer0_outputs(6531) <= 1'b0;
    layer0_outputs(6532) <= not a;
    layer0_outputs(6533) <= 1'b1;
    layer0_outputs(6534) <= a;
    layer0_outputs(6535) <= b;
    layer0_outputs(6536) <= a or b;
    layer0_outputs(6537) <= b and not a;
    layer0_outputs(6538) <= 1'b1;
    layer0_outputs(6539) <= not (a xor b);
    layer0_outputs(6540) <= not b or a;
    layer0_outputs(6541) <= a or b;
    layer0_outputs(6542) <= not a;
    layer0_outputs(6543) <= 1'b1;
    layer0_outputs(6544) <= a xor b;
    layer0_outputs(6545) <= a;
    layer0_outputs(6546) <= b;
    layer0_outputs(6547) <= not (a xor b);
    layer0_outputs(6548) <= a xor b;
    layer0_outputs(6549) <= not (a xor b);
    layer0_outputs(6550) <= not (a or b);
    layer0_outputs(6551) <= a or b;
    layer0_outputs(6552) <= 1'b1;
    layer0_outputs(6553) <= not b;
    layer0_outputs(6554) <= not (a and b);
    layer0_outputs(6555) <= not a;
    layer0_outputs(6556) <= not b or a;
    layer0_outputs(6557) <= 1'b1;
    layer0_outputs(6558) <= not a;
    layer0_outputs(6559) <= not (a or b);
    layer0_outputs(6560) <= not b or a;
    layer0_outputs(6561) <= a or b;
    layer0_outputs(6562) <= not (a xor b);
    layer0_outputs(6563) <= a xor b;
    layer0_outputs(6564) <= a and not b;
    layer0_outputs(6565) <= a xor b;
    layer0_outputs(6566) <= not a or b;
    layer0_outputs(6567) <= not (a or b);
    layer0_outputs(6568) <= a;
    layer0_outputs(6569) <= b and not a;
    layer0_outputs(6570) <= a xor b;
    layer0_outputs(6571) <= a or b;
    layer0_outputs(6572) <= not (a or b);
    layer0_outputs(6573) <= a and not b;
    layer0_outputs(6574) <= not (a xor b);
    layer0_outputs(6575) <= not (a xor b);
    layer0_outputs(6576) <= 1'b0;
    layer0_outputs(6577) <= not (a xor b);
    layer0_outputs(6578) <= b;
    layer0_outputs(6579) <= a and not b;
    layer0_outputs(6580) <= b and not a;
    layer0_outputs(6581) <= a or b;
    layer0_outputs(6582) <= not (a or b);
    layer0_outputs(6583) <= not a;
    layer0_outputs(6584) <= b and not a;
    layer0_outputs(6585) <= not b or a;
    layer0_outputs(6586) <= b;
    layer0_outputs(6587) <= a xor b;
    layer0_outputs(6588) <= not (a xor b);
    layer0_outputs(6589) <= not (a or b);
    layer0_outputs(6590) <= not (a or b);
    layer0_outputs(6591) <= not b or a;
    layer0_outputs(6592) <= a and not b;
    layer0_outputs(6593) <= 1'b1;
    layer0_outputs(6594) <= a or b;
    layer0_outputs(6595) <= not b or a;
    layer0_outputs(6596) <= a xor b;
    layer0_outputs(6597) <= a or b;
    layer0_outputs(6598) <= a and not b;
    layer0_outputs(6599) <= 1'b0;
    layer0_outputs(6600) <= not (a xor b);
    layer0_outputs(6601) <= a and b;
    layer0_outputs(6602) <= a and b;
    layer0_outputs(6603) <= a;
    layer0_outputs(6604) <= not a;
    layer0_outputs(6605) <= a or b;
    layer0_outputs(6606) <= b and not a;
    layer0_outputs(6607) <= a xor b;
    layer0_outputs(6608) <= not b or a;
    layer0_outputs(6609) <= not a or b;
    layer0_outputs(6610) <= not (a and b);
    layer0_outputs(6611) <= not (a xor b);
    layer0_outputs(6612) <= a and b;
    layer0_outputs(6613) <= not b;
    layer0_outputs(6614) <= not b or a;
    layer0_outputs(6615) <= not a or b;
    layer0_outputs(6616) <= a or b;
    layer0_outputs(6617) <= not (a xor b);
    layer0_outputs(6618) <= not b or a;
    layer0_outputs(6619) <= a or b;
    layer0_outputs(6620) <= not (a or b);
    layer0_outputs(6621) <= not (a xor b);
    layer0_outputs(6622) <= not (a or b);
    layer0_outputs(6623) <= not (a or b);
    layer0_outputs(6624) <= not b;
    layer0_outputs(6625) <= b;
    layer0_outputs(6626) <= not b or a;
    layer0_outputs(6627) <= a and not b;
    layer0_outputs(6628) <= not (a or b);
    layer0_outputs(6629) <= a or b;
    layer0_outputs(6630) <= a and not b;
    layer0_outputs(6631) <= not a;
    layer0_outputs(6632) <= not a;
    layer0_outputs(6633) <= 1'b0;
    layer0_outputs(6634) <= not a;
    layer0_outputs(6635) <= not a or b;
    layer0_outputs(6636) <= not (a and b);
    layer0_outputs(6637) <= a;
    layer0_outputs(6638) <= not a or b;
    layer0_outputs(6639) <= a and b;
    layer0_outputs(6640) <= not (a xor b);
    layer0_outputs(6641) <= not (a or b);
    layer0_outputs(6642) <= not a or b;
    layer0_outputs(6643) <= not b or a;
    layer0_outputs(6644) <= 1'b1;
    layer0_outputs(6645) <= not (a or b);
    layer0_outputs(6646) <= a xor b;
    layer0_outputs(6647) <= not b or a;
    layer0_outputs(6648) <= a and not b;
    layer0_outputs(6649) <= not (a and b);
    layer0_outputs(6650) <= a or b;
    layer0_outputs(6651) <= not a or b;
    layer0_outputs(6652) <= not b;
    layer0_outputs(6653) <= not a;
    layer0_outputs(6654) <= a or b;
    layer0_outputs(6655) <= not a or b;
    layer0_outputs(6656) <= b and not a;
    layer0_outputs(6657) <= not (a or b);
    layer0_outputs(6658) <= b and not a;
    layer0_outputs(6659) <= not a or b;
    layer0_outputs(6660) <= b;
    layer0_outputs(6661) <= not (a or b);
    layer0_outputs(6662) <= 1'b1;
    layer0_outputs(6663) <= a or b;
    layer0_outputs(6664) <= a or b;
    layer0_outputs(6665) <= not (a xor b);
    layer0_outputs(6666) <= not a;
    layer0_outputs(6667) <= a or b;
    layer0_outputs(6668) <= b;
    layer0_outputs(6669) <= not b;
    layer0_outputs(6670) <= not b or a;
    layer0_outputs(6671) <= not (a xor b);
    layer0_outputs(6672) <= not a;
    layer0_outputs(6673) <= b and not a;
    layer0_outputs(6674) <= a or b;
    layer0_outputs(6675) <= not (a or b);
    layer0_outputs(6676) <= not a;
    layer0_outputs(6677) <= b;
    layer0_outputs(6678) <= not b;
    layer0_outputs(6679) <= a xor b;
    layer0_outputs(6680) <= not b or a;
    layer0_outputs(6681) <= a or b;
    layer0_outputs(6682) <= not a;
    layer0_outputs(6683) <= not a;
    layer0_outputs(6684) <= not b;
    layer0_outputs(6685) <= not a;
    layer0_outputs(6686) <= not b or a;
    layer0_outputs(6687) <= not a;
    layer0_outputs(6688) <= not (a or b);
    layer0_outputs(6689) <= a and b;
    layer0_outputs(6690) <= b and not a;
    layer0_outputs(6691) <= a xor b;
    layer0_outputs(6692) <= a or b;
    layer0_outputs(6693) <= not a or b;
    layer0_outputs(6694) <= not (a or b);
    layer0_outputs(6695) <= not b;
    layer0_outputs(6696) <= not a or b;
    layer0_outputs(6697) <= a xor b;
    layer0_outputs(6698) <= not b;
    layer0_outputs(6699) <= a or b;
    layer0_outputs(6700) <= not (a and b);
    layer0_outputs(6701) <= a or b;
    layer0_outputs(6702) <= a;
    layer0_outputs(6703) <= not b;
    layer0_outputs(6704) <= a;
    layer0_outputs(6705) <= 1'b1;
    layer0_outputs(6706) <= a and not b;
    layer0_outputs(6707) <= not (a xor b);
    layer0_outputs(6708) <= a xor b;
    layer0_outputs(6709) <= not a;
    layer0_outputs(6710) <= a xor b;
    layer0_outputs(6711) <= not (a xor b);
    layer0_outputs(6712) <= not b or a;
    layer0_outputs(6713) <= not (a or b);
    layer0_outputs(6714) <= not a or b;
    layer0_outputs(6715) <= not a;
    layer0_outputs(6716) <= not (a or b);
    layer0_outputs(6717) <= a and b;
    layer0_outputs(6718) <= not (a or b);
    layer0_outputs(6719) <= not b or a;
    layer0_outputs(6720) <= not b;
    layer0_outputs(6721) <= not b;
    layer0_outputs(6722) <= b and not a;
    layer0_outputs(6723) <= not (a xor b);
    layer0_outputs(6724) <= 1'b1;
    layer0_outputs(6725) <= 1'b1;
    layer0_outputs(6726) <= a or b;
    layer0_outputs(6727) <= a or b;
    layer0_outputs(6728) <= not a;
    layer0_outputs(6729) <= not (a xor b);
    layer0_outputs(6730) <= b;
    layer0_outputs(6731) <= a and b;
    layer0_outputs(6732) <= b;
    layer0_outputs(6733) <= not (a or b);
    layer0_outputs(6734) <= not a;
    layer0_outputs(6735) <= not (a or b);
    layer0_outputs(6736) <= not (a or b);
    layer0_outputs(6737) <= 1'b0;
    layer0_outputs(6738) <= a xor b;
    layer0_outputs(6739) <= b;
    layer0_outputs(6740) <= b;
    layer0_outputs(6741) <= not b or a;
    layer0_outputs(6742) <= b and not a;
    layer0_outputs(6743) <= a and b;
    layer0_outputs(6744) <= not a;
    layer0_outputs(6745) <= not a or b;
    layer0_outputs(6746) <= 1'b1;
    layer0_outputs(6747) <= b;
    layer0_outputs(6748) <= a;
    layer0_outputs(6749) <= b and not a;
    layer0_outputs(6750) <= not a or b;
    layer0_outputs(6751) <= a or b;
    layer0_outputs(6752) <= a or b;
    layer0_outputs(6753) <= not b or a;
    layer0_outputs(6754) <= not a;
    layer0_outputs(6755) <= not (a or b);
    layer0_outputs(6756) <= 1'b1;
    layer0_outputs(6757) <= b and not a;
    layer0_outputs(6758) <= a;
    layer0_outputs(6759) <= not (a xor b);
    layer0_outputs(6760) <= a or b;
    layer0_outputs(6761) <= a and b;
    layer0_outputs(6762) <= b and not a;
    layer0_outputs(6763) <= b;
    layer0_outputs(6764) <= not a or b;
    layer0_outputs(6765) <= not b or a;
    layer0_outputs(6766) <= not b or a;
    layer0_outputs(6767) <= not a;
    layer0_outputs(6768) <= not b or a;
    layer0_outputs(6769) <= not b or a;
    layer0_outputs(6770) <= a and b;
    layer0_outputs(6771) <= not (a xor b);
    layer0_outputs(6772) <= not a;
    layer0_outputs(6773) <= not a or b;
    layer0_outputs(6774) <= not a or b;
    layer0_outputs(6775) <= a or b;
    layer0_outputs(6776) <= 1'b1;
    layer0_outputs(6777) <= b and not a;
    layer0_outputs(6778) <= not a;
    layer0_outputs(6779) <= b and not a;
    layer0_outputs(6780) <= not (a and b);
    layer0_outputs(6781) <= b and not a;
    layer0_outputs(6782) <= b;
    layer0_outputs(6783) <= a or b;
    layer0_outputs(6784) <= not a or b;
    layer0_outputs(6785) <= 1'b0;
    layer0_outputs(6786) <= a xor b;
    layer0_outputs(6787) <= not (a or b);
    layer0_outputs(6788) <= not a;
    layer0_outputs(6789) <= a xor b;
    layer0_outputs(6790) <= a and b;
    layer0_outputs(6791) <= not (a or b);
    layer0_outputs(6792) <= not (a or b);
    layer0_outputs(6793) <= not a or b;
    layer0_outputs(6794) <= not (a or b);
    layer0_outputs(6795) <= b and not a;
    layer0_outputs(6796) <= a;
    layer0_outputs(6797) <= 1'b1;
    layer0_outputs(6798) <= a or b;
    layer0_outputs(6799) <= not b or a;
    layer0_outputs(6800) <= not (a or b);
    layer0_outputs(6801) <= a or b;
    layer0_outputs(6802) <= a or b;
    layer0_outputs(6803) <= a xor b;
    layer0_outputs(6804) <= a;
    layer0_outputs(6805) <= not (a and b);
    layer0_outputs(6806) <= not a or b;
    layer0_outputs(6807) <= a or b;
    layer0_outputs(6808) <= b and not a;
    layer0_outputs(6809) <= not b or a;
    layer0_outputs(6810) <= a or b;
    layer0_outputs(6811) <= a xor b;
    layer0_outputs(6812) <= not a;
    layer0_outputs(6813) <= not (a and b);
    layer0_outputs(6814) <= not a or b;
    layer0_outputs(6815) <= a xor b;
    layer0_outputs(6816) <= not b or a;
    layer0_outputs(6817) <= a or b;
    layer0_outputs(6818) <= a or b;
    layer0_outputs(6819) <= not (a or b);
    layer0_outputs(6820) <= a;
    layer0_outputs(6821) <= not b or a;
    layer0_outputs(6822) <= not b or a;
    layer0_outputs(6823) <= b and not a;
    layer0_outputs(6824) <= b and not a;
    layer0_outputs(6825) <= not b or a;
    layer0_outputs(6826) <= not b or a;
    layer0_outputs(6827) <= b and not a;
    layer0_outputs(6828) <= not a or b;
    layer0_outputs(6829) <= not a;
    layer0_outputs(6830) <= not (a or b);
    layer0_outputs(6831) <= a or b;
    layer0_outputs(6832) <= a or b;
    layer0_outputs(6833) <= a or b;
    layer0_outputs(6834) <= a or b;
    layer0_outputs(6835) <= b and not a;
    layer0_outputs(6836) <= a;
    layer0_outputs(6837) <= not a;
    layer0_outputs(6838) <= b and not a;
    layer0_outputs(6839) <= not a;
    layer0_outputs(6840) <= b;
    layer0_outputs(6841) <= not (a xor b);
    layer0_outputs(6842) <= not (a xor b);
    layer0_outputs(6843) <= not b;
    layer0_outputs(6844) <= a xor b;
    layer0_outputs(6845) <= not b;
    layer0_outputs(6846) <= not (a xor b);
    layer0_outputs(6847) <= not a or b;
    layer0_outputs(6848) <= a or b;
    layer0_outputs(6849) <= not b or a;
    layer0_outputs(6850) <= not b or a;
    layer0_outputs(6851) <= not b;
    layer0_outputs(6852) <= a xor b;
    layer0_outputs(6853) <= not b;
    layer0_outputs(6854) <= not b;
    layer0_outputs(6855) <= a or b;
    layer0_outputs(6856) <= a or b;
    layer0_outputs(6857) <= not a or b;
    layer0_outputs(6858) <= a or b;
    layer0_outputs(6859) <= b and not a;
    layer0_outputs(6860) <= a xor b;
    layer0_outputs(6861) <= not a;
    layer0_outputs(6862) <= not (a or b);
    layer0_outputs(6863) <= not (a or b);
    layer0_outputs(6864) <= not (a or b);
    layer0_outputs(6865) <= not a;
    layer0_outputs(6866) <= not a or b;
    layer0_outputs(6867) <= b;
    layer0_outputs(6868) <= b;
    layer0_outputs(6869) <= not a;
    layer0_outputs(6870) <= b and not a;
    layer0_outputs(6871) <= not (a xor b);
    layer0_outputs(6872) <= not a or b;
    layer0_outputs(6873) <= a and not b;
    layer0_outputs(6874) <= a xor b;
    layer0_outputs(6875) <= a xor b;
    layer0_outputs(6876) <= a xor b;
    layer0_outputs(6877) <= not (a xor b);
    layer0_outputs(6878) <= b and not a;
    layer0_outputs(6879) <= not a;
    layer0_outputs(6880) <= b and not a;
    layer0_outputs(6881) <= not b or a;
    layer0_outputs(6882) <= a and not b;
    layer0_outputs(6883) <= not a;
    layer0_outputs(6884) <= not (a and b);
    layer0_outputs(6885) <= a;
    layer0_outputs(6886) <= not a;
    layer0_outputs(6887) <= a or b;
    layer0_outputs(6888) <= not (a xor b);
    layer0_outputs(6889) <= a or b;
    layer0_outputs(6890) <= b;
    layer0_outputs(6891) <= b;
    layer0_outputs(6892) <= not b or a;
    layer0_outputs(6893) <= a or b;
    layer0_outputs(6894) <= not a or b;
    layer0_outputs(6895) <= not a or b;
    layer0_outputs(6896) <= not (a or b);
    layer0_outputs(6897) <= a or b;
    layer0_outputs(6898) <= not (a xor b);
    layer0_outputs(6899) <= not a or b;
    layer0_outputs(6900) <= not (a or b);
    layer0_outputs(6901) <= not (a or b);
    layer0_outputs(6902) <= not (a and b);
    layer0_outputs(6903) <= b and not a;
    layer0_outputs(6904) <= not a;
    layer0_outputs(6905) <= a and b;
    layer0_outputs(6906) <= not a;
    layer0_outputs(6907) <= b and not a;
    layer0_outputs(6908) <= not (a and b);
    layer0_outputs(6909) <= a or b;
    layer0_outputs(6910) <= b;
    layer0_outputs(6911) <= b;
    layer0_outputs(6912) <= 1'b1;
    layer0_outputs(6913) <= a and b;
    layer0_outputs(6914) <= a or b;
    layer0_outputs(6915) <= a or b;
    layer0_outputs(6916) <= not a;
    layer0_outputs(6917) <= not b;
    layer0_outputs(6918) <= not b or a;
    layer0_outputs(6919) <= b and not a;
    layer0_outputs(6920) <= not b or a;
    layer0_outputs(6921) <= not (a or b);
    layer0_outputs(6922) <= not b;
    layer0_outputs(6923) <= 1'b1;
    layer0_outputs(6924) <= not (a and b);
    layer0_outputs(6925) <= b;
    layer0_outputs(6926) <= not b;
    layer0_outputs(6927) <= not (a or b);
    layer0_outputs(6928) <= not (a or b);
    layer0_outputs(6929) <= not (a and b);
    layer0_outputs(6930) <= not (a or b);
    layer0_outputs(6931) <= not (a xor b);
    layer0_outputs(6932) <= not (a or b);
    layer0_outputs(6933) <= a and not b;
    layer0_outputs(6934) <= not b or a;
    layer0_outputs(6935) <= a and b;
    layer0_outputs(6936) <= 1'b0;
    layer0_outputs(6937) <= a or b;
    layer0_outputs(6938) <= not (a or b);
    layer0_outputs(6939) <= not b or a;
    layer0_outputs(6940) <= not (a or b);
    layer0_outputs(6941) <= not (a xor b);
    layer0_outputs(6942) <= a xor b;
    layer0_outputs(6943) <= not (a and b);
    layer0_outputs(6944) <= b and not a;
    layer0_outputs(6945) <= b and not a;
    layer0_outputs(6946) <= not (a or b);
    layer0_outputs(6947) <= not b or a;
    layer0_outputs(6948) <= a and not b;
    layer0_outputs(6949) <= not (a xor b);
    layer0_outputs(6950) <= a;
    layer0_outputs(6951) <= a xor b;
    layer0_outputs(6952) <= not b or a;
    layer0_outputs(6953) <= b;
    layer0_outputs(6954) <= not (a or b);
    layer0_outputs(6955) <= a or b;
    layer0_outputs(6956) <= not (a xor b);
    layer0_outputs(6957) <= not b or a;
    layer0_outputs(6958) <= not (a xor b);
    layer0_outputs(6959) <= not (a or b);
    layer0_outputs(6960) <= a or b;
    layer0_outputs(6961) <= a or b;
    layer0_outputs(6962) <= a or b;
    layer0_outputs(6963) <= b and not a;
    layer0_outputs(6964) <= not (a or b);
    layer0_outputs(6965) <= a;
    layer0_outputs(6966) <= not a or b;
    layer0_outputs(6967) <= a;
    layer0_outputs(6968) <= not a;
    layer0_outputs(6969) <= b;
    layer0_outputs(6970) <= a and not b;
    layer0_outputs(6971) <= a and not b;
    layer0_outputs(6972) <= not (a or b);
    layer0_outputs(6973) <= not (a xor b);
    layer0_outputs(6974) <= 1'b0;
    layer0_outputs(6975) <= not a or b;
    layer0_outputs(6976) <= not (a or b);
    layer0_outputs(6977) <= not (a xor b);
    layer0_outputs(6978) <= a or b;
    layer0_outputs(6979) <= a xor b;
    layer0_outputs(6980) <= not b or a;
    layer0_outputs(6981) <= a xor b;
    layer0_outputs(6982) <= not (a xor b);
    layer0_outputs(6983) <= not (a or b);
    layer0_outputs(6984) <= a;
    layer0_outputs(6985) <= not a or b;
    layer0_outputs(6986) <= not (a xor b);
    layer0_outputs(6987) <= b;
    layer0_outputs(6988) <= a;
    layer0_outputs(6989) <= 1'b1;
    layer0_outputs(6990) <= not (a xor b);
    layer0_outputs(6991) <= not (a xor b);
    layer0_outputs(6992) <= a or b;
    layer0_outputs(6993) <= not (a xor b);
    layer0_outputs(6994) <= not a or b;
    layer0_outputs(6995) <= not (a xor b);
    layer0_outputs(6996) <= not a or b;
    layer0_outputs(6997) <= a xor b;
    layer0_outputs(6998) <= a xor b;
    layer0_outputs(6999) <= a xor b;
    layer0_outputs(7000) <= a xor b;
    layer0_outputs(7001) <= not a;
    layer0_outputs(7002) <= not (a and b);
    layer0_outputs(7003) <= not (a xor b);
    layer0_outputs(7004) <= a or b;
    layer0_outputs(7005) <= a or b;
    layer0_outputs(7006) <= a;
    layer0_outputs(7007) <= a or b;
    layer0_outputs(7008) <= not b or a;
    layer0_outputs(7009) <= not (a or b);
    layer0_outputs(7010) <= not a;
    layer0_outputs(7011) <= not (a or b);
    layer0_outputs(7012) <= not b;
    layer0_outputs(7013) <= 1'b1;
    layer0_outputs(7014) <= b;
    layer0_outputs(7015) <= not (a xor b);
    layer0_outputs(7016) <= a and b;
    layer0_outputs(7017) <= not a;
    layer0_outputs(7018) <= b;
    layer0_outputs(7019) <= b and not a;
    layer0_outputs(7020) <= b;
    layer0_outputs(7021) <= not b;
    layer0_outputs(7022) <= not a;
    layer0_outputs(7023) <= a;
    layer0_outputs(7024) <= not (a xor b);
    layer0_outputs(7025) <= not (a or b);
    layer0_outputs(7026) <= not (a xor b);
    layer0_outputs(7027) <= not (a xor b);
    layer0_outputs(7028) <= not (a xor b);
    layer0_outputs(7029) <= not a or b;
    layer0_outputs(7030) <= a;
    layer0_outputs(7031) <= not b;
    layer0_outputs(7032) <= 1'b0;
    layer0_outputs(7033) <= b;
    layer0_outputs(7034) <= a and b;
    layer0_outputs(7035) <= 1'b1;
    layer0_outputs(7036) <= not (a or b);
    layer0_outputs(7037) <= a or b;
    layer0_outputs(7038) <= a;
    layer0_outputs(7039) <= not b;
    layer0_outputs(7040) <= not b;
    layer0_outputs(7041) <= a;
    layer0_outputs(7042) <= 1'b1;
    layer0_outputs(7043) <= a xor b;
    layer0_outputs(7044) <= not (a or b);
    layer0_outputs(7045) <= not a;
    layer0_outputs(7046) <= not b or a;
    layer0_outputs(7047) <= a;
    layer0_outputs(7048) <= a xor b;
    layer0_outputs(7049) <= a xor b;
    layer0_outputs(7050) <= not b;
    layer0_outputs(7051) <= b;
    layer0_outputs(7052) <= not (a or b);
    layer0_outputs(7053) <= not (a or b);
    layer0_outputs(7054) <= not b;
    layer0_outputs(7055) <= a and b;
    layer0_outputs(7056) <= not b;
    layer0_outputs(7057) <= not a;
    layer0_outputs(7058) <= not a or b;
    layer0_outputs(7059) <= a xor b;
    layer0_outputs(7060) <= not (a or b);
    layer0_outputs(7061) <= not (a or b);
    layer0_outputs(7062) <= not a;
    layer0_outputs(7063) <= a xor b;
    layer0_outputs(7064) <= not b or a;
    layer0_outputs(7065) <= not a;
    layer0_outputs(7066) <= a or b;
    layer0_outputs(7067) <= b;
    layer0_outputs(7068) <= b and not a;
    layer0_outputs(7069) <= not b;
    layer0_outputs(7070) <= a xor b;
    layer0_outputs(7071) <= a xor b;
    layer0_outputs(7072) <= not (a xor b);
    layer0_outputs(7073) <= not (a or b);
    layer0_outputs(7074) <= not a;
    layer0_outputs(7075) <= not (a or b);
    layer0_outputs(7076) <= not b;
    layer0_outputs(7077) <= 1'b0;
    layer0_outputs(7078) <= b;
    layer0_outputs(7079) <= not b;
    layer0_outputs(7080) <= not (a and b);
    layer0_outputs(7081) <= a and b;
    layer0_outputs(7082) <= not (a xor b);
    layer0_outputs(7083) <= a or b;
    layer0_outputs(7084) <= a and not b;
    layer0_outputs(7085) <= 1'b1;
    layer0_outputs(7086) <= a and not b;
    layer0_outputs(7087) <= not b;
    layer0_outputs(7088) <= not b;
    layer0_outputs(7089) <= a and not b;
    layer0_outputs(7090) <= not b or a;
    layer0_outputs(7091) <= b and not a;
    layer0_outputs(7092) <= a and not b;
    layer0_outputs(7093) <= not (a or b);
    layer0_outputs(7094) <= b and not a;
    layer0_outputs(7095) <= a;
    layer0_outputs(7096) <= a;
    layer0_outputs(7097) <= a or b;
    layer0_outputs(7098) <= b;
    layer0_outputs(7099) <= a and not b;
    layer0_outputs(7100) <= b;
    layer0_outputs(7101) <= not b or a;
    layer0_outputs(7102) <= not b or a;
    layer0_outputs(7103) <= not (a and b);
    layer0_outputs(7104) <= not (a and b);
    layer0_outputs(7105) <= b;
    layer0_outputs(7106) <= not a;
    layer0_outputs(7107) <= not b or a;
    layer0_outputs(7108) <= not a or b;
    layer0_outputs(7109) <= not a or b;
    layer0_outputs(7110) <= a or b;
    layer0_outputs(7111) <= not a;
    layer0_outputs(7112) <= a;
    layer0_outputs(7113) <= not a or b;
    layer0_outputs(7114) <= not b or a;
    layer0_outputs(7115) <= not b;
    layer0_outputs(7116) <= a xor b;
    layer0_outputs(7117) <= b and not a;
    layer0_outputs(7118) <= not (a xor b);
    layer0_outputs(7119) <= b and not a;
    layer0_outputs(7120) <= b;
    layer0_outputs(7121) <= 1'b0;
    layer0_outputs(7122) <= not b;
    layer0_outputs(7123) <= a and b;
    layer0_outputs(7124) <= not a or b;
    layer0_outputs(7125) <= not (a or b);
    layer0_outputs(7126) <= not (a or b);
    layer0_outputs(7127) <= b and not a;
    layer0_outputs(7128) <= a xor b;
    layer0_outputs(7129) <= b and not a;
    layer0_outputs(7130) <= not (a or b);
    layer0_outputs(7131) <= not (a or b);
    layer0_outputs(7132) <= a;
    layer0_outputs(7133) <= a xor b;
    layer0_outputs(7134) <= a or b;
    layer0_outputs(7135) <= a and not b;
    layer0_outputs(7136) <= a or b;
    layer0_outputs(7137) <= a and not b;
    layer0_outputs(7138) <= 1'b0;
    layer0_outputs(7139) <= not b or a;
    layer0_outputs(7140) <= b;
    layer0_outputs(7141) <= not b;
    layer0_outputs(7142) <= not a or b;
    layer0_outputs(7143) <= not (a or b);
    layer0_outputs(7144) <= not a or b;
    layer0_outputs(7145) <= a and not b;
    layer0_outputs(7146) <= not (a xor b);
    layer0_outputs(7147) <= not b or a;
    layer0_outputs(7148) <= 1'b0;
    layer0_outputs(7149) <= not (a or b);
    layer0_outputs(7150) <= a or b;
    layer0_outputs(7151) <= not b;
    layer0_outputs(7152) <= a and not b;
    layer0_outputs(7153) <= not (a or b);
    layer0_outputs(7154) <= 1'b1;
    layer0_outputs(7155) <= not b;
    layer0_outputs(7156) <= b and not a;
    layer0_outputs(7157) <= a or b;
    layer0_outputs(7158) <= b and not a;
    layer0_outputs(7159) <= a and b;
    layer0_outputs(7160) <= a xor b;
    layer0_outputs(7161) <= not (a or b);
    layer0_outputs(7162) <= a;
    layer0_outputs(7163) <= a;
    layer0_outputs(7164) <= a or b;
    layer0_outputs(7165) <= not a;
    layer0_outputs(7166) <= a;
    layer0_outputs(7167) <= not b;
    layer0_outputs(7168) <= not b;
    layer0_outputs(7169) <= not b or a;
    layer0_outputs(7170) <= not a or b;
    layer0_outputs(7171) <= not a;
    layer0_outputs(7172) <= not b or a;
    layer0_outputs(7173) <= not a or b;
    layer0_outputs(7174) <= a xor b;
    layer0_outputs(7175) <= a;
    layer0_outputs(7176) <= not b;
    layer0_outputs(7177) <= a and b;
    layer0_outputs(7178) <= not a;
    layer0_outputs(7179) <= a xor b;
    layer0_outputs(7180) <= b and not a;
    layer0_outputs(7181) <= b;
    layer0_outputs(7182) <= a or b;
    layer0_outputs(7183) <= a or b;
    layer0_outputs(7184) <= not b;
    layer0_outputs(7185) <= a;
    layer0_outputs(7186) <= a or b;
    layer0_outputs(7187) <= not b or a;
    layer0_outputs(7188) <= a;
    layer0_outputs(7189) <= a and not b;
    layer0_outputs(7190) <= a xor b;
    layer0_outputs(7191) <= a and not b;
    layer0_outputs(7192) <= a xor b;
    layer0_outputs(7193) <= not a;
    layer0_outputs(7194) <= not b;
    layer0_outputs(7195) <= not b;
    layer0_outputs(7196) <= a and not b;
    layer0_outputs(7197) <= not a or b;
    layer0_outputs(7198) <= a xor b;
    layer0_outputs(7199) <= not (a xor b);
    layer0_outputs(7200) <= not a or b;
    layer0_outputs(7201) <= a xor b;
    layer0_outputs(7202) <= not (a or b);
    layer0_outputs(7203) <= a;
    layer0_outputs(7204) <= a and not b;
    layer0_outputs(7205) <= a and not b;
    layer0_outputs(7206) <= a and b;
    layer0_outputs(7207) <= a and not b;
    layer0_outputs(7208) <= not a or b;
    layer0_outputs(7209) <= b and not a;
    layer0_outputs(7210) <= not (a xor b);
    layer0_outputs(7211) <= a;
    layer0_outputs(7212) <= not b or a;
    layer0_outputs(7213) <= not b;
    layer0_outputs(7214) <= a xor b;
    layer0_outputs(7215) <= not (a or b);
    layer0_outputs(7216) <= a or b;
    layer0_outputs(7217) <= a;
    layer0_outputs(7218) <= a and b;
    layer0_outputs(7219) <= not (a or b);
    layer0_outputs(7220) <= not (a and b);
    layer0_outputs(7221) <= not (a or b);
    layer0_outputs(7222) <= a or b;
    layer0_outputs(7223) <= a and not b;
    layer0_outputs(7224) <= not (a or b);
    layer0_outputs(7225) <= a and not b;
    layer0_outputs(7226) <= not (a or b);
    layer0_outputs(7227) <= 1'b0;
    layer0_outputs(7228) <= not a;
    layer0_outputs(7229) <= not b;
    layer0_outputs(7230) <= b and not a;
    layer0_outputs(7231) <= a xor b;
    layer0_outputs(7232) <= not b;
    layer0_outputs(7233) <= b and not a;
    layer0_outputs(7234) <= a and b;
    layer0_outputs(7235) <= not a or b;
    layer0_outputs(7236) <= not (a or b);
    layer0_outputs(7237) <= a;
    layer0_outputs(7238) <= a and not b;
    layer0_outputs(7239) <= a or b;
    layer0_outputs(7240) <= b;
    layer0_outputs(7241) <= not b or a;
    layer0_outputs(7242) <= a or b;
    layer0_outputs(7243) <= b;
    layer0_outputs(7244) <= not b;
    layer0_outputs(7245) <= a xor b;
    layer0_outputs(7246) <= a or b;
    layer0_outputs(7247) <= not b or a;
    layer0_outputs(7248) <= not (a or b);
    layer0_outputs(7249) <= a xor b;
    layer0_outputs(7250) <= not (a and b);
    layer0_outputs(7251) <= not b;
    layer0_outputs(7252) <= a or b;
    layer0_outputs(7253) <= 1'b0;
    layer0_outputs(7254) <= not (a or b);
    layer0_outputs(7255) <= a xor b;
    layer0_outputs(7256) <= not (a or b);
    layer0_outputs(7257) <= a or b;
    layer0_outputs(7258) <= a;
    layer0_outputs(7259) <= not b or a;
    layer0_outputs(7260) <= not b or a;
    layer0_outputs(7261) <= not a or b;
    layer0_outputs(7262) <= not a;
    layer0_outputs(7263) <= 1'b1;
    layer0_outputs(7264) <= not (a and b);
    layer0_outputs(7265) <= a xor b;
    layer0_outputs(7266) <= a xor b;
    layer0_outputs(7267) <= not a or b;
    layer0_outputs(7268) <= a or b;
    layer0_outputs(7269) <= not (a xor b);
    layer0_outputs(7270) <= a and not b;
    layer0_outputs(7271) <= b and not a;
    layer0_outputs(7272) <= a or b;
    layer0_outputs(7273) <= not a;
    layer0_outputs(7274) <= b;
    layer0_outputs(7275) <= 1'b0;
    layer0_outputs(7276) <= not b or a;
    layer0_outputs(7277) <= b;
    layer0_outputs(7278) <= not (a or b);
    layer0_outputs(7279) <= not (a or b);
    layer0_outputs(7280) <= not a or b;
    layer0_outputs(7281) <= not a or b;
    layer0_outputs(7282) <= a xor b;
    layer0_outputs(7283) <= a or b;
    layer0_outputs(7284) <= a and not b;
    layer0_outputs(7285) <= a;
    layer0_outputs(7286) <= not (a xor b);
    layer0_outputs(7287) <= b;
    layer0_outputs(7288) <= not (a xor b);
    layer0_outputs(7289) <= not b or a;
    layer0_outputs(7290) <= a and not b;
    layer0_outputs(7291) <= not (a xor b);
    layer0_outputs(7292) <= a xor b;
    layer0_outputs(7293) <= b;
    layer0_outputs(7294) <= a or b;
    layer0_outputs(7295) <= not (a or b);
    layer0_outputs(7296) <= b;
    layer0_outputs(7297) <= not (a xor b);
    layer0_outputs(7298) <= not b;
    layer0_outputs(7299) <= not b;
    layer0_outputs(7300) <= a xor b;
    layer0_outputs(7301) <= 1'b1;
    layer0_outputs(7302) <= not b;
    layer0_outputs(7303) <= not a;
    layer0_outputs(7304) <= a and not b;
    layer0_outputs(7305) <= not (a xor b);
    layer0_outputs(7306) <= a or b;
    layer0_outputs(7307) <= not (a or b);
    layer0_outputs(7308) <= b and not a;
    layer0_outputs(7309) <= not (a or b);
    layer0_outputs(7310) <= not a or b;
    layer0_outputs(7311) <= not (a and b);
    layer0_outputs(7312) <= not (a or b);
    layer0_outputs(7313) <= not a or b;
    layer0_outputs(7314) <= a or b;
    layer0_outputs(7315) <= a;
    layer0_outputs(7316) <= not b or a;
    layer0_outputs(7317) <= a;
    layer0_outputs(7318) <= a xor b;
    layer0_outputs(7319) <= b;
    layer0_outputs(7320) <= not (a or b);
    layer0_outputs(7321) <= b;
    layer0_outputs(7322) <= not (a xor b);
    layer0_outputs(7323) <= not b;
    layer0_outputs(7324) <= not (a or b);
    layer0_outputs(7325) <= not a;
    layer0_outputs(7326) <= not a or b;
    layer0_outputs(7327) <= b and not a;
    layer0_outputs(7328) <= b and not a;
    layer0_outputs(7329) <= not a;
    layer0_outputs(7330) <= not (a or b);
    layer0_outputs(7331) <= not a or b;
    layer0_outputs(7332) <= not b;
    layer0_outputs(7333) <= not a or b;
    layer0_outputs(7334) <= not a;
    layer0_outputs(7335) <= not (a or b);
    layer0_outputs(7336) <= b;
    layer0_outputs(7337) <= b and not a;
    layer0_outputs(7338) <= not a;
    layer0_outputs(7339) <= 1'b0;
    layer0_outputs(7340) <= b;
    layer0_outputs(7341) <= not (a or b);
    layer0_outputs(7342) <= not a or b;
    layer0_outputs(7343) <= a or b;
    layer0_outputs(7344) <= a and not b;
    layer0_outputs(7345) <= not (a xor b);
    layer0_outputs(7346) <= not (a xor b);
    layer0_outputs(7347) <= a xor b;
    layer0_outputs(7348) <= not (a or b);
    layer0_outputs(7349) <= not (a xor b);
    layer0_outputs(7350) <= not (a xor b);
    layer0_outputs(7351) <= not b or a;
    layer0_outputs(7352) <= not (a and b);
    layer0_outputs(7353) <= not (a xor b);
    layer0_outputs(7354) <= b;
    layer0_outputs(7355) <= a xor b;
    layer0_outputs(7356) <= b and not a;
    layer0_outputs(7357) <= a;
    layer0_outputs(7358) <= a and b;
    layer0_outputs(7359) <= not a or b;
    layer0_outputs(7360) <= not (a xor b);
    layer0_outputs(7361) <= not (a or b);
    layer0_outputs(7362) <= not (a xor b);
    layer0_outputs(7363) <= a;
    layer0_outputs(7364) <= not b or a;
    layer0_outputs(7365) <= a and b;
    layer0_outputs(7366) <= a or b;
    layer0_outputs(7367) <= 1'b0;
    layer0_outputs(7368) <= not (a or b);
    layer0_outputs(7369) <= a xor b;
    layer0_outputs(7370) <= not (a or b);
    layer0_outputs(7371) <= not a or b;
    layer0_outputs(7372) <= not (a and b);
    layer0_outputs(7373) <= not (a or b);
    layer0_outputs(7374) <= not (a or b);
    layer0_outputs(7375) <= a and not b;
    layer0_outputs(7376) <= not (a or b);
    layer0_outputs(7377) <= not a;
    layer0_outputs(7378) <= not a;
    layer0_outputs(7379) <= not a;
    layer0_outputs(7380) <= 1'b1;
    layer0_outputs(7381) <= a xor b;
    layer0_outputs(7382) <= b;
    layer0_outputs(7383) <= a or b;
    layer0_outputs(7384) <= a or b;
    layer0_outputs(7385) <= not b;
    layer0_outputs(7386) <= a and b;
    layer0_outputs(7387) <= a or b;
    layer0_outputs(7388) <= not (a and b);
    layer0_outputs(7389) <= not (a or b);
    layer0_outputs(7390) <= not (a or b);
    layer0_outputs(7391) <= a xor b;
    layer0_outputs(7392) <= not a or b;
    layer0_outputs(7393) <= b and not a;
    layer0_outputs(7394) <= not b or a;
    layer0_outputs(7395) <= a;
    layer0_outputs(7396) <= a xor b;
    layer0_outputs(7397) <= not (a or b);
    layer0_outputs(7398) <= not (a or b);
    layer0_outputs(7399) <= not (a or b);
    layer0_outputs(7400) <= a;
    layer0_outputs(7401) <= a or b;
    layer0_outputs(7402) <= not (a and b);
    layer0_outputs(7403) <= not b;
    layer0_outputs(7404) <= a xor b;
    layer0_outputs(7405) <= a xor b;
    layer0_outputs(7406) <= 1'b0;
    layer0_outputs(7407) <= not (a xor b);
    layer0_outputs(7408) <= a and b;
    layer0_outputs(7409) <= not b;
    layer0_outputs(7410) <= 1'b1;
    layer0_outputs(7411) <= not b or a;
    layer0_outputs(7412) <= a;
    layer0_outputs(7413) <= not a or b;
    layer0_outputs(7414) <= 1'b0;
    layer0_outputs(7415) <= not (a or b);
    layer0_outputs(7416) <= not a or b;
    layer0_outputs(7417) <= not (a xor b);
    layer0_outputs(7418) <= not a;
    layer0_outputs(7419) <= b;
    layer0_outputs(7420) <= a or b;
    layer0_outputs(7421) <= not b;
    layer0_outputs(7422) <= a and not b;
    layer0_outputs(7423) <= b;
    layer0_outputs(7424) <= a and not b;
    layer0_outputs(7425) <= a and not b;
    layer0_outputs(7426) <= 1'b0;
    layer0_outputs(7427) <= a;
    layer0_outputs(7428) <= a xor b;
    layer0_outputs(7429) <= b and not a;
    layer0_outputs(7430) <= a or b;
    layer0_outputs(7431) <= not (a and b);
    layer0_outputs(7432) <= b;
    layer0_outputs(7433) <= not a;
    layer0_outputs(7434) <= a;
    layer0_outputs(7435) <= a or b;
    layer0_outputs(7436) <= not b or a;
    layer0_outputs(7437) <= not a;
    layer0_outputs(7438) <= not a or b;
    layer0_outputs(7439) <= not a;
    layer0_outputs(7440) <= not b;
    layer0_outputs(7441) <= not b;
    layer0_outputs(7442) <= not b or a;
    layer0_outputs(7443) <= 1'b1;
    layer0_outputs(7444) <= a or b;
    layer0_outputs(7445) <= a or b;
    layer0_outputs(7446) <= a or b;
    layer0_outputs(7447) <= not (a or b);
    layer0_outputs(7448) <= not (a or b);
    layer0_outputs(7449) <= not a;
    layer0_outputs(7450) <= b;
    layer0_outputs(7451) <= a xor b;
    layer0_outputs(7452) <= a xor b;
    layer0_outputs(7453) <= not (a or b);
    layer0_outputs(7454) <= 1'b0;
    layer0_outputs(7455) <= a xor b;
    layer0_outputs(7456) <= not (a xor b);
    layer0_outputs(7457) <= a xor b;
    layer0_outputs(7458) <= not a;
    layer0_outputs(7459) <= not (a and b);
    layer0_outputs(7460) <= a or b;
    layer0_outputs(7461) <= a or b;
    layer0_outputs(7462) <= a xor b;
    layer0_outputs(7463) <= a;
    layer0_outputs(7464) <= not b;
    layer0_outputs(7465) <= not a;
    layer0_outputs(7466) <= a or b;
    layer0_outputs(7467) <= a and not b;
    layer0_outputs(7468) <= b;
    layer0_outputs(7469) <= b;
    layer0_outputs(7470) <= a or b;
    layer0_outputs(7471) <= not (a or b);
    layer0_outputs(7472) <= b;
    layer0_outputs(7473) <= not (a xor b);
    layer0_outputs(7474) <= not (a xor b);
    layer0_outputs(7475) <= b and not a;
    layer0_outputs(7476) <= not (a or b);
    layer0_outputs(7477) <= a and b;
    layer0_outputs(7478) <= b;
    layer0_outputs(7479) <= not b;
    layer0_outputs(7480) <= a and not b;
    layer0_outputs(7481) <= 1'b0;
    layer0_outputs(7482) <= not (a xor b);
    layer0_outputs(7483) <= a and not b;
    layer0_outputs(7484) <= not b;
    layer0_outputs(7485) <= a or b;
    layer0_outputs(7486) <= not a;
    layer0_outputs(7487) <= not a or b;
    layer0_outputs(7488) <= not a;
    layer0_outputs(7489) <= b and not a;
    layer0_outputs(7490) <= not (a and b);
    layer0_outputs(7491) <= not (a or b);
    layer0_outputs(7492) <= a and b;
    layer0_outputs(7493) <= not b or a;
    layer0_outputs(7494) <= b and not a;
    layer0_outputs(7495) <= a xor b;
    layer0_outputs(7496) <= not b or a;
    layer0_outputs(7497) <= a;
    layer0_outputs(7498) <= not a or b;
    layer0_outputs(7499) <= not b;
    layer0_outputs(7500) <= a and b;
    layer0_outputs(7501) <= not a;
    layer0_outputs(7502) <= a or b;
    layer0_outputs(7503) <= not (a or b);
    layer0_outputs(7504) <= not a;
    layer0_outputs(7505) <= not a;
    layer0_outputs(7506) <= not b;
    layer0_outputs(7507) <= not a;
    layer0_outputs(7508) <= not b or a;
    layer0_outputs(7509) <= b;
    layer0_outputs(7510) <= a xor b;
    layer0_outputs(7511) <= not (a and b);
    layer0_outputs(7512) <= a or b;
    layer0_outputs(7513) <= a;
    layer0_outputs(7514) <= a xor b;
    layer0_outputs(7515) <= not (a or b);
    layer0_outputs(7516) <= not a;
    layer0_outputs(7517) <= not (a xor b);
    layer0_outputs(7518) <= a xor b;
    layer0_outputs(7519) <= 1'b1;
    layer0_outputs(7520) <= not a;
    layer0_outputs(7521) <= a;
    layer0_outputs(7522) <= b;
    layer0_outputs(7523) <= not (a or b);
    layer0_outputs(7524) <= a xor b;
    layer0_outputs(7525) <= a or b;
    layer0_outputs(7526) <= not (a xor b);
    layer0_outputs(7527) <= 1'b1;
    layer0_outputs(7528) <= not b or a;
    layer0_outputs(7529) <= not (a xor b);
    layer0_outputs(7530) <= not (a xor b);
    layer0_outputs(7531) <= not (a xor b);
    layer0_outputs(7532) <= a;
    layer0_outputs(7533) <= not b;
    layer0_outputs(7534) <= b and not a;
    layer0_outputs(7535) <= not a or b;
    layer0_outputs(7536) <= a xor b;
    layer0_outputs(7537) <= a xor b;
    layer0_outputs(7538) <= not (a and b);
    layer0_outputs(7539) <= a xor b;
    layer0_outputs(7540) <= a or b;
    layer0_outputs(7541) <= b and not a;
    layer0_outputs(7542) <= not (a or b);
    layer0_outputs(7543) <= a and not b;
    layer0_outputs(7544) <= b and not a;
    layer0_outputs(7545) <= not a;
    layer0_outputs(7546) <= a and not b;
    layer0_outputs(7547) <= a or b;
    layer0_outputs(7548) <= not b;
    layer0_outputs(7549) <= a xor b;
    layer0_outputs(7550) <= not (a or b);
    layer0_outputs(7551) <= not b or a;
    layer0_outputs(7552) <= not a or b;
    layer0_outputs(7553) <= a xor b;
    layer0_outputs(7554) <= a xor b;
    layer0_outputs(7555) <= a;
    layer0_outputs(7556) <= not b;
    layer0_outputs(7557) <= not (a or b);
    layer0_outputs(7558) <= b and not a;
    layer0_outputs(7559) <= a;
    layer0_outputs(7560) <= a or b;
    layer0_outputs(7561) <= not b or a;
    layer0_outputs(7562) <= a or b;
    layer0_outputs(7563) <= not (a or b);
    layer0_outputs(7564) <= a or b;
    layer0_outputs(7565) <= b;
    layer0_outputs(7566) <= not (a and b);
    layer0_outputs(7567) <= not (a or b);
    layer0_outputs(7568) <= not (a xor b);
    layer0_outputs(7569) <= not (a xor b);
    layer0_outputs(7570) <= b and not a;
    layer0_outputs(7571) <= a and not b;
    layer0_outputs(7572) <= a or b;
    layer0_outputs(7573) <= not (a xor b);
    layer0_outputs(7574) <= not (a or b);
    layer0_outputs(7575) <= b;
    layer0_outputs(7576) <= not (a or b);
    layer0_outputs(7577) <= a xor b;
    layer0_outputs(7578) <= a and not b;
    layer0_outputs(7579) <= not (a xor b);
    layer0_outputs(7580) <= not (a xor b);
    layer0_outputs(7581) <= not a or b;
    layer0_outputs(7582) <= a or b;
    layer0_outputs(7583) <= not (a or b);
    layer0_outputs(7584) <= not (a xor b);
    layer0_outputs(7585) <= a;
    layer0_outputs(7586) <= a and b;
    layer0_outputs(7587) <= not a;
    layer0_outputs(7588) <= b and not a;
    layer0_outputs(7589) <= a and not b;
    layer0_outputs(7590) <= not (a xor b);
    layer0_outputs(7591) <= a;
    layer0_outputs(7592) <= b;
    layer0_outputs(7593) <= a;
    layer0_outputs(7594) <= not (a xor b);
    layer0_outputs(7595) <= 1'b0;
    layer0_outputs(7596) <= not (a or b);
    layer0_outputs(7597) <= a;
    layer0_outputs(7598) <= b and not a;
    layer0_outputs(7599) <= not b or a;
    layer0_outputs(7600) <= a or b;
    layer0_outputs(7601) <= a and b;
    layer0_outputs(7602) <= not a;
    layer0_outputs(7603) <= a or b;
    layer0_outputs(7604) <= a;
    layer0_outputs(7605) <= a;
    layer0_outputs(7606) <= not (a or b);
    layer0_outputs(7607) <= not a;
    layer0_outputs(7608) <= not b or a;
    layer0_outputs(7609) <= not a;
    layer0_outputs(7610) <= not a;
    layer0_outputs(7611) <= a and not b;
    layer0_outputs(7612) <= a or b;
    layer0_outputs(7613) <= a and not b;
    layer0_outputs(7614) <= not (a or b);
    layer0_outputs(7615) <= not b or a;
    layer0_outputs(7616) <= not (a and b);
    layer0_outputs(7617) <= a or b;
    layer0_outputs(7618) <= a;
    layer0_outputs(7619) <= not b or a;
    layer0_outputs(7620) <= not b;
    layer0_outputs(7621) <= a or b;
    layer0_outputs(7622) <= a;
    layer0_outputs(7623) <= not a or b;
    layer0_outputs(7624) <= a and not b;
    layer0_outputs(7625) <= not (a or b);
    layer0_outputs(7626) <= a;
    layer0_outputs(7627) <= not b;
    layer0_outputs(7628) <= a or b;
    layer0_outputs(7629) <= not b;
    layer0_outputs(7630) <= a xor b;
    layer0_outputs(7631) <= b;
    layer0_outputs(7632) <= not a;
    layer0_outputs(7633) <= a and not b;
    layer0_outputs(7634) <= not (a or b);
    layer0_outputs(7635) <= not a;
    layer0_outputs(7636) <= not b or a;
    layer0_outputs(7637) <= 1'b1;
    layer0_outputs(7638) <= not a;
    layer0_outputs(7639) <= a;
    layer0_outputs(7640) <= not (a or b);
    layer0_outputs(7641) <= not (a or b);
    layer0_outputs(7642) <= 1'b0;
    layer0_outputs(7643) <= not (a and b);
    layer0_outputs(7644) <= not a or b;
    layer0_outputs(7645) <= a;
    layer0_outputs(7646) <= not (a or b);
    layer0_outputs(7647) <= b and not a;
    layer0_outputs(7648) <= a;
    layer0_outputs(7649) <= a and not b;
    layer0_outputs(7650) <= not (a or b);
    layer0_outputs(7651) <= a xor b;
    layer0_outputs(7652) <= a and b;
    layer0_outputs(7653) <= not a or b;
    layer0_outputs(7654) <= not (a or b);
    layer0_outputs(7655) <= not b or a;
    layer0_outputs(7656) <= 1'b1;
    layer0_outputs(7657) <= a;
    layer0_outputs(7658) <= a or b;
    layer0_outputs(7659) <= not (a or b);
    layer0_outputs(7660) <= a and b;
    layer0_outputs(7661) <= not (a or b);
    layer0_outputs(7662) <= a and not b;
    layer0_outputs(7663) <= not (a xor b);
    layer0_outputs(7664) <= not a or b;
    layer0_outputs(7665) <= 1'b0;
    layer0_outputs(7666) <= not (a xor b);
    layer0_outputs(7667) <= a and not b;
    layer0_outputs(7668) <= not (a xor b);
    layer0_outputs(7669) <= a and not b;
    layer0_outputs(7670) <= not (a xor b);
    layer0_outputs(7671) <= 1'b1;
    layer0_outputs(7672) <= b and not a;
    layer0_outputs(7673) <= not b or a;
    layer0_outputs(7674) <= b;
    layer0_outputs(7675) <= a xor b;
    layer0_outputs(7676) <= a or b;
    layer0_outputs(7677) <= not b or a;
    layer0_outputs(7678) <= b and not a;
    layer0_outputs(7679) <= 1'b0;
    layer1_outputs(0) <= b and not a;
    layer1_outputs(1) <= a and b;
    layer1_outputs(2) <= not (a xor b);
    layer1_outputs(3) <= not (a and b);
    layer1_outputs(4) <= a or b;
    layer1_outputs(5) <= 1'b0;
    layer1_outputs(6) <= not a;
    layer1_outputs(7) <= not a;
    layer1_outputs(8) <= not b;
    layer1_outputs(9) <= a xor b;
    layer1_outputs(10) <= not a or b;
    layer1_outputs(11) <= not (a and b);
    layer1_outputs(12) <= b and not a;
    layer1_outputs(13) <= not b;
    layer1_outputs(14) <= b;
    layer1_outputs(15) <= not (a and b);
    layer1_outputs(16) <= a or b;
    layer1_outputs(17) <= b and not a;
    layer1_outputs(18) <= a xor b;
    layer1_outputs(19) <= b;
    layer1_outputs(20) <= not (a xor b);
    layer1_outputs(21) <= a and not b;
    layer1_outputs(22) <= a or b;
    layer1_outputs(23) <= a and b;
    layer1_outputs(24) <= a xor b;
    layer1_outputs(25) <= a;
    layer1_outputs(26) <= not b or a;
    layer1_outputs(27) <= a or b;
    layer1_outputs(28) <= a and b;
    layer1_outputs(29) <= not b;
    layer1_outputs(30) <= b;
    layer1_outputs(31) <= not b or a;
    layer1_outputs(32) <= not b or a;
    layer1_outputs(33) <= not (a or b);
    layer1_outputs(34) <= not (a xor b);
    layer1_outputs(35) <= b;
    layer1_outputs(36) <= a;
    layer1_outputs(37) <= a;
    layer1_outputs(38) <= a xor b;
    layer1_outputs(39) <= not b or a;
    layer1_outputs(40) <= a or b;
    layer1_outputs(41) <= a and b;
    layer1_outputs(42) <= b;
    layer1_outputs(43) <= not b;
    layer1_outputs(44) <= a xor b;
    layer1_outputs(45) <= a and not b;
    layer1_outputs(46) <= not b;
    layer1_outputs(47) <= not b;
    layer1_outputs(48) <= a;
    layer1_outputs(49) <= a xor b;
    layer1_outputs(50) <= not a or b;
    layer1_outputs(51) <= not a;
    layer1_outputs(52) <= not (a xor b);
    layer1_outputs(53) <= not a;
    layer1_outputs(54) <= a and not b;
    layer1_outputs(55) <= a and b;
    layer1_outputs(56) <= not a;
    layer1_outputs(57) <= not b or a;
    layer1_outputs(58) <= a or b;
    layer1_outputs(59) <= a and not b;
    layer1_outputs(60) <= not (a xor b);
    layer1_outputs(61) <= a and b;
    layer1_outputs(62) <= not a or b;
    layer1_outputs(63) <= a xor b;
    layer1_outputs(64) <= a and not b;
    layer1_outputs(65) <= not a;
    layer1_outputs(66) <= not b or a;
    layer1_outputs(67) <= a;
    layer1_outputs(68) <= a xor b;
    layer1_outputs(69) <= not (a xor b);
    layer1_outputs(70) <= a and b;
    layer1_outputs(71) <= 1'b0;
    layer1_outputs(72) <= b;
    layer1_outputs(73) <= not a;
    layer1_outputs(74) <= not a or b;
    layer1_outputs(75) <= b;
    layer1_outputs(76) <= not b or a;
    layer1_outputs(77) <= a;
    layer1_outputs(78) <= a xor b;
    layer1_outputs(79) <= b and not a;
    layer1_outputs(80) <= b;
    layer1_outputs(81) <= not b;
    layer1_outputs(82) <= b;
    layer1_outputs(83) <= a and not b;
    layer1_outputs(84) <= not b;
    layer1_outputs(85) <= a;
    layer1_outputs(86) <= b and not a;
    layer1_outputs(87) <= a and not b;
    layer1_outputs(88) <= b and not a;
    layer1_outputs(89) <= not (a and b);
    layer1_outputs(90) <= a and b;
    layer1_outputs(91) <= b and not a;
    layer1_outputs(92) <= a or b;
    layer1_outputs(93) <= a and not b;
    layer1_outputs(94) <= a or b;
    layer1_outputs(95) <= a and not b;
    layer1_outputs(96) <= a xor b;
    layer1_outputs(97) <= a or b;
    layer1_outputs(98) <= b and not a;
    layer1_outputs(99) <= not b;
    layer1_outputs(100) <= not a or b;
    layer1_outputs(101) <= b and not a;
    layer1_outputs(102) <= not b;
    layer1_outputs(103) <= not (a or b);
    layer1_outputs(104) <= not b;
    layer1_outputs(105) <= 1'b1;
    layer1_outputs(106) <= not (a and b);
    layer1_outputs(107) <= not (a xor b);
    layer1_outputs(108) <= a and not b;
    layer1_outputs(109) <= b and not a;
    layer1_outputs(110) <= not a or b;
    layer1_outputs(111) <= not b;
    layer1_outputs(112) <= a xor b;
    layer1_outputs(113) <= not b or a;
    layer1_outputs(114) <= a xor b;
    layer1_outputs(115) <= a;
    layer1_outputs(116) <= a;
    layer1_outputs(117) <= a xor b;
    layer1_outputs(118) <= a;
    layer1_outputs(119) <= a xor b;
    layer1_outputs(120) <= a;
    layer1_outputs(121) <= b and not a;
    layer1_outputs(122) <= not (a xor b);
    layer1_outputs(123) <= b and not a;
    layer1_outputs(124) <= a xor b;
    layer1_outputs(125) <= not a;
    layer1_outputs(126) <= a and not b;
    layer1_outputs(127) <= a or b;
    layer1_outputs(128) <= not (a or b);
    layer1_outputs(129) <= not a;
    layer1_outputs(130) <= not b;
    layer1_outputs(131) <= b;
    layer1_outputs(132) <= a and b;
    layer1_outputs(133) <= b and not a;
    layer1_outputs(134) <= a and not b;
    layer1_outputs(135) <= a;
    layer1_outputs(136) <= not b;
    layer1_outputs(137) <= a and b;
    layer1_outputs(138) <= a and b;
    layer1_outputs(139) <= not b or a;
    layer1_outputs(140) <= a;
    layer1_outputs(141) <= not b;
    layer1_outputs(142) <= a and not b;
    layer1_outputs(143) <= b;
    layer1_outputs(144) <= a or b;
    layer1_outputs(145) <= not b or a;
    layer1_outputs(146) <= a and b;
    layer1_outputs(147) <= a and b;
    layer1_outputs(148) <= b and not a;
    layer1_outputs(149) <= a;
    layer1_outputs(150) <= b and not a;
    layer1_outputs(151) <= not (a or b);
    layer1_outputs(152) <= not b;
    layer1_outputs(153) <= not b or a;
    layer1_outputs(154) <= b and not a;
    layer1_outputs(155) <= not (a or b);
    layer1_outputs(156) <= a and b;
    layer1_outputs(157) <= not a;
    layer1_outputs(158) <= a and not b;
    layer1_outputs(159) <= not b;
    layer1_outputs(160) <= not a;
    layer1_outputs(161) <= 1'b0;
    layer1_outputs(162) <= b;
    layer1_outputs(163) <= not (a xor b);
    layer1_outputs(164) <= not a or b;
    layer1_outputs(165) <= a or b;
    layer1_outputs(166) <= not (a xor b);
    layer1_outputs(167) <= not a or b;
    layer1_outputs(168) <= a xor b;
    layer1_outputs(169) <= not b;
    layer1_outputs(170) <= not a;
    layer1_outputs(171) <= a and b;
    layer1_outputs(172) <= b and not a;
    layer1_outputs(173) <= not (a and b);
    layer1_outputs(174) <= 1'b0;
    layer1_outputs(175) <= a;
    layer1_outputs(176) <= not (a and b);
    layer1_outputs(177) <= a and not b;
    layer1_outputs(178) <= not a;
    layer1_outputs(179) <= not a;
    layer1_outputs(180) <= not (a or b);
    layer1_outputs(181) <= not a;
    layer1_outputs(182) <= not b or a;
    layer1_outputs(183) <= b;
    layer1_outputs(184) <= b and not a;
    layer1_outputs(185) <= not (a and b);
    layer1_outputs(186) <= a and b;
    layer1_outputs(187) <= not a or b;
    layer1_outputs(188) <= not (a or b);
    layer1_outputs(189) <= not b or a;
    layer1_outputs(190) <= a and b;
    layer1_outputs(191) <= not (a or b);
    layer1_outputs(192) <= not a or b;
    layer1_outputs(193) <= a and b;
    layer1_outputs(194) <= not (a or b);
    layer1_outputs(195) <= not b;
    layer1_outputs(196) <= not (a or b);
    layer1_outputs(197) <= 1'b0;
    layer1_outputs(198) <= not a or b;
    layer1_outputs(199) <= not (a xor b);
    layer1_outputs(200) <= not b;
    layer1_outputs(201) <= a and not b;
    layer1_outputs(202) <= not (a and b);
    layer1_outputs(203) <= a or b;
    layer1_outputs(204) <= not (a xor b);
    layer1_outputs(205) <= b and not a;
    layer1_outputs(206) <= a;
    layer1_outputs(207) <= b;
    layer1_outputs(208) <= not (a xor b);
    layer1_outputs(209) <= not a;
    layer1_outputs(210) <= a;
    layer1_outputs(211) <= a and not b;
    layer1_outputs(212) <= a;
    layer1_outputs(213) <= b;
    layer1_outputs(214) <= a and not b;
    layer1_outputs(215) <= a or b;
    layer1_outputs(216) <= a;
    layer1_outputs(217) <= 1'b1;
    layer1_outputs(218) <= b and not a;
    layer1_outputs(219) <= not (a and b);
    layer1_outputs(220) <= not (a xor b);
    layer1_outputs(221) <= b;
    layer1_outputs(222) <= a or b;
    layer1_outputs(223) <= a xor b;
    layer1_outputs(224) <= b and not a;
    layer1_outputs(225) <= not (a xor b);
    layer1_outputs(226) <= b;
    layer1_outputs(227) <= b;
    layer1_outputs(228) <= a and b;
    layer1_outputs(229) <= not a or b;
    layer1_outputs(230) <= 1'b1;
    layer1_outputs(231) <= not a or b;
    layer1_outputs(232) <= b;
    layer1_outputs(233) <= not (a xor b);
    layer1_outputs(234) <= not (a xor b);
    layer1_outputs(235) <= b;
    layer1_outputs(236) <= b;
    layer1_outputs(237) <= a and b;
    layer1_outputs(238) <= a xor b;
    layer1_outputs(239) <= a and b;
    layer1_outputs(240) <= not b;
    layer1_outputs(241) <= not (a or b);
    layer1_outputs(242) <= not (a or b);
    layer1_outputs(243) <= not b or a;
    layer1_outputs(244) <= not (a or b);
    layer1_outputs(245) <= not a or b;
    layer1_outputs(246) <= a xor b;
    layer1_outputs(247) <= b;
    layer1_outputs(248) <= a and b;
    layer1_outputs(249) <= a xor b;
    layer1_outputs(250) <= b and not a;
    layer1_outputs(251) <= a and b;
    layer1_outputs(252) <= a;
    layer1_outputs(253) <= b;
    layer1_outputs(254) <= a and b;
    layer1_outputs(255) <= a;
    layer1_outputs(256) <= not (a xor b);
    layer1_outputs(257) <= b;
    layer1_outputs(258) <= not b or a;
    layer1_outputs(259) <= a xor b;
    layer1_outputs(260) <= b;
    layer1_outputs(261) <= a or b;
    layer1_outputs(262) <= a or b;
    layer1_outputs(263) <= a and not b;
    layer1_outputs(264) <= b and not a;
    layer1_outputs(265) <= not (a or b);
    layer1_outputs(266) <= not (a xor b);
    layer1_outputs(267) <= not (a or b);
    layer1_outputs(268) <= not (a xor b);
    layer1_outputs(269) <= not a;
    layer1_outputs(270) <= not (a or b);
    layer1_outputs(271) <= b and not a;
    layer1_outputs(272) <= not a;
    layer1_outputs(273) <= not b;
    layer1_outputs(274) <= not b;
    layer1_outputs(275) <= a and b;
    layer1_outputs(276) <= not a or b;
    layer1_outputs(277) <= a and not b;
    layer1_outputs(278) <= a and b;
    layer1_outputs(279) <= not (a and b);
    layer1_outputs(280) <= not b;
    layer1_outputs(281) <= b;
    layer1_outputs(282) <= a or b;
    layer1_outputs(283) <= b;
    layer1_outputs(284) <= not (a and b);
    layer1_outputs(285) <= not (a and b);
    layer1_outputs(286) <= b;
    layer1_outputs(287) <= a xor b;
    layer1_outputs(288) <= not a;
    layer1_outputs(289) <= a xor b;
    layer1_outputs(290) <= not (a xor b);
    layer1_outputs(291) <= b;
    layer1_outputs(292) <= b;
    layer1_outputs(293) <= a and not b;
    layer1_outputs(294) <= a and b;
    layer1_outputs(295) <= a and not b;
    layer1_outputs(296) <= a and b;
    layer1_outputs(297) <= a;
    layer1_outputs(298) <= a xor b;
    layer1_outputs(299) <= not (a and b);
    layer1_outputs(300) <= a and not b;
    layer1_outputs(301) <= 1'b0;
    layer1_outputs(302) <= not a or b;
    layer1_outputs(303) <= not (a xor b);
    layer1_outputs(304) <= not a;
    layer1_outputs(305) <= a and b;
    layer1_outputs(306) <= a;
    layer1_outputs(307) <= a and b;
    layer1_outputs(308) <= a or b;
    layer1_outputs(309) <= b and not a;
    layer1_outputs(310) <= a and not b;
    layer1_outputs(311) <= b;
    layer1_outputs(312) <= not (a xor b);
    layer1_outputs(313) <= a and b;
    layer1_outputs(314) <= not (a or b);
    layer1_outputs(315) <= a xor b;
    layer1_outputs(316) <= a or b;
    layer1_outputs(317) <= not (a or b);
    layer1_outputs(318) <= not b;
    layer1_outputs(319) <= not (a and b);
    layer1_outputs(320) <= not (a or b);
    layer1_outputs(321) <= not (a or b);
    layer1_outputs(322) <= not a;
    layer1_outputs(323) <= not (a and b);
    layer1_outputs(324) <= a xor b;
    layer1_outputs(325) <= a xor b;
    layer1_outputs(326) <= not b;
    layer1_outputs(327) <= not b or a;
    layer1_outputs(328) <= not a or b;
    layer1_outputs(329) <= a and b;
    layer1_outputs(330) <= a and b;
    layer1_outputs(331) <= not (a or b);
    layer1_outputs(332) <= b;
    layer1_outputs(333) <= b and not a;
    layer1_outputs(334) <= not b;
    layer1_outputs(335) <= a and not b;
    layer1_outputs(336) <= b;
    layer1_outputs(337) <= not b;
    layer1_outputs(338) <= b;
    layer1_outputs(339) <= a xor b;
    layer1_outputs(340) <= not b or a;
    layer1_outputs(341) <= a xor b;
    layer1_outputs(342) <= not (a xor b);
    layer1_outputs(343) <= not (a or b);
    layer1_outputs(344) <= a;
    layer1_outputs(345) <= not b;
    layer1_outputs(346) <= not (a xor b);
    layer1_outputs(347) <= not (a and b);
    layer1_outputs(348) <= not (a and b);
    layer1_outputs(349) <= a and not b;
    layer1_outputs(350) <= b;
    layer1_outputs(351) <= not (a xor b);
    layer1_outputs(352) <= not b or a;
    layer1_outputs(353) <= not (a xor b);
    layer1_outputs(354) <= not (a xor b);
    layer1_outputs(355) <= not a;
    layer1_outputs(356) <= a;
    layer1_outputs(357) <= not a;
    layer1_outputs(358) <= not a;
    layer1_outputs(359) <= not b or a;
    layer1_outputs(360) <= a xor b;
    layer1_outputs(361) <= a or b;
    layer1_outputs(362) <= a xor b;
    layer1_outputs(363) <= b and not a;
    layer1_outputs(364) <= not b or a;
    layer1_outputs(365) <= not (a and b);
    layer1_outputs(366) <= not (a xor b);
    layer1_outputs(367) <= b and not a;
    layer1_outputs(368) <= not b or a;
    layer1_outputs(369) <= not b;
    layer1_outputs(370) <= not a;
    layer1_outputs(371) <= b and not a;
    layer1_outputs(372) <= 1'b1;
    layer1_outputs(373) <= not a or b;
    layer1_outputs(374) <= a;
    layer1_outputs(375) <= a xor b;
    layer1_outputs(376) <= b;
    layer1_outputs(377) <= a;
    layer1_outputs(378) <= not (a or b);
    layer1_outputs(379) <= 1'b1;
    layer1_outputs(380) <= not (a xor b);
    layer1_outputs(381) <= not (a or b);
    layer1_outputs(382) <= not a;
    layer1_outputs(383) <= b;
    layer1_outputs(384) <= a xor b;
    layer1_outputs(385) <= not b;
    layer1_outputs(386) <= not b;
    layer1_outputs(387) <= not (a or b);
    layer1_outputs(388) <= not (a xor b);
    layer1_outputs(389) <= b;
    layer1_outputs(390) <= not a;
    layer1_outputs(391) <= b and not a;
    layer1_outputs(392) <= a xor b;
    layer1_outputs(393) <= b;
    layer1_outputs(394) <= not a or b;
    layer1_outputs(395) <= a;
    layer1_outputs(396) <= a and b;
    layer1_outputs(397) <= a and not b;
    layer1_outputs(398) <= not a;
    layer1_outputs(399) <= a;
    layer1_outputs(400) <= a xor b;
    layer1_outputs(401) <= a;
    layer1_outputs(402) <= a;
    layer1_outputs(403) <= a and not b;
    layer1_outputs(404) <= a and not b;
    layer1_outputs(405) <= b;
    layer1_outputs(406) <= b;
    layer1_outputs(407) <= a or b;
    layer1_outputs(408) <= a or b;
    layer1_outputs(409) <= not a or b;
    layer1_outputs(410) <= b;
    layer1_outputs(411) <= not (a and b);
    layer1_outputs(412) <= not (a and b);
    layer1_outputs(413) <= not a;
    layer1_outputs(414) <= not b;
    layer1_outputs(415) <= not b or a;
    layer1_outputs(416) <= not a;
    layer1_outputs(417) <= a or b;
    layer1_outputs(418) <= not (a or b);
    layer1_outputs(419) <= not a or b;
    layer1_outputs(420) <= not (a or b);
    layer1_outputs(421) <= not b or a;
    layer1_outputs(422) <= not a;
    layer1_outputs(423) <= a xor b;
    layer1_outputs(424) <= a xor b;
    layer1_outputs(425) <= a xor b;
    layer1_outputs(426) <= not (a and b);
    layer1_outputs(427) <= a xor b;
    layer1_outputs(428) <= not b or a;
    layer1_outputs(429) <= 1'b0;
    layer1_outputs(430) <= not b;
    layer1_outputs(431) <= 1'b0;
    layer1_outputs(432) <= a or b;
    layer1_outputs(433) <= 1'b1;
    layer1_outputs(434) <= not (a and b);
    layer1_outputs(435) <= a and not b;
    layer1_outputs(436) <= a;
    layer1_outputs(437) <= not a or b;
    layer1_outputs(438) <= not (a and b);
    layer1_outputs(439) <= b and not a;
    layer1_outputs(440) <= not (a xor b);
    layer1_outputs(441) <= not (a and b);
    layer1_outputs(442) <= b and not a;
    layer1_outputs(443) <= 1'b1;
    layer1_outputs(444) <= not b or a;
    layer1_outputs(445) <= a and b;
    layer1_outputs(446) <= a;
    layer1_outputs(447) <= a and b;
    layer1_outputs(448) <= a and b;
    layer1_outputs(449) <= a or b;
    layer1_outputs(450) <= a and not b;
    layer1_outputs(451) <= a and b;
    layer1_outputs(452) <= not (a or b);
    layer1_outputs(453) <= not b or a;
    layer1_outputs(454) <= not a or b;
    layer1_outputs(455) <= not (a xor b);
    layer1_outputs(456) <= a or b;
    layer1_outputs(457) <= a and not b;
    layer1_outputs(458) <= not a or b;
    layer1_outputs(459) <= a and b;
    layer1_outputs(460) <= 1'b1;
    layer1_outputs(461) <= a and b;
    layer1_outputs(462) <= not b;
    layer1_outputs(463) <= b and not a;
    layer1_outputs(464) <= a and b;
    layer1_outputs(465) <= not a;
    layer1_outputs(466) <= not (a or b);
    layer1_outputs(467) <= a and b;
    layer1_outputs(468) <= not a;
    layer1_outputs(469) <= not a or b;
    layer1_outputs(470) <= b and not a;
    layer1_outputs(471) <= not (a xor b);
    layer1_outputs(472) <= a and b;
    layer1_outputs(473) <= not b or a;
    layer1_outputs(474) <= a;
    layer1_outputs(475) <= a or b;
    layer1_outputs(476) <= a and b;
    layer1_outputs(477) <= a xor b;
    layer1_outputs(478) <= a;
    layer1_outputs(479) <= a or b;
    layer1_outputs(480) <= b;
    layer1_outputs(481) <= not a or b;
    layer1_outputs(482) <= a and b;
    layer1_outputs(483) <= a or b;
    layer1_outputs(484) <= a and not b;
    layer1_outputs(485) <= not b or a;
    layer1_outputs(486) <= a and b;
    layer1_outputs(487) <= not a;
    layer1_outputs(488) <= not a;
    layer1_outputs(489) <= not a or b;
    layer1_outputs(490) <= a and b;
    layer1_outputs(491) <= not b or a;
    layer1_outputs(492) <= not (a xor b);
    layer1_outputs(493) <= not a;
    layer1_outputs(494) <= b and not a;
    layer1_outputs(495) <= b;
    layer1_outputs(496) <= a;
    layer1_outputs(497) <= not a or b;
    layer1_outputs(498) <= not b or a;
    layer1_outputs(499) <= 1'b0;
    layer1_outputs(500) <= not a;
    layer1_outputs(501) <= not a or b;
    layer1_outputs(502) <= a;
    layer1_outputs(503) <= a xor b;
    layer1_outputs(504) <= not a;
    layer1_outputs(505) <= b and not a;
    layer1_outputs(506) <= not b;
    layer1_outputs(507) <= a and not b;
    layer1_outputs(508) <= a and b;
    layer1_outputs(509) <= a or b;
    layer1_outputs(510) <= not (a xor b);
    layer1_outputs(511) <= a or b;
    layer1_outputs(512) <= b;
    layer1_outputs(513) <= not (a xor b);
    layer1_outputs(514) <= a xor b;
    layer1_outputs(515) <= not b or a;
    layer1_outputs(516) <= not a or b;
    layer1_outputs(517) <= not (a and b);
    layer1_outputs(518) <= b and not a;
    layer1_outputs(519) <= not a or b;
    layer1_outputs(520) <= not (a or b);
    layer1_outputs(521) <= not (a and b);
    layer1_outputs(522) <= b;
    layer1_outputs(523) <= not (a xor b);
    layer1_outputs(524) <= not (a or b);
    layer1_outputs(525) <= a;
    layer1_outputs(526) <= not (a xor b);
    layer1_outputs(527) <= not a;
    layer1_outputs(528) <= not a or b;
    layer1_outputs(529) <= a and not b;
    layer1_outputs(530) <= not (a xor b);
    layer1_outputs(531) <= not a;
    layer1_outputs(532) <= a and b;
    layer1_outputs(533) <= b and not a;
    layer1_outputs(534) <= not b or a;
    layer1_outputs(535) <= b;
    layer1_outputs(536) <= not (a xor b);
    layer1_outputs(537) <= a and not b;
    layer1_outputs(538) <= not b;
    layer1_outputs(539) <= b;
    layer1_outputs(540) <= a xor b;
    layer1_outputs(541) <= b;
    layer1_outputs(542) <= not (a xor b);
    layer1_outputs(543) <= a and b;
    layer1_outputs(544) <= a;
    layer1_outputs(545) <= a;
    layer1_outputs(546) <= a;
    layer1_outputs(547) <= a xor b;
    layer1_outputs(548) <= a;
    layer1_outputs(549) <= a or b;
    layer1_outputs(550) <= not (a and b);
    layer1_outputs(551) <= b and not a;
    layer1_outputs(552) <= not (a xor b);
    layer1_outputs(553) <= a;
    layer1_outputs(554) <= b;
    layer1_outputs(555) <= a xor b;
    layer1_outputs(556) <= b and not a;
    layer1_outputs(557) <= a;
    layer1_outputs(558) <= not b or a;
    layer1_outputs(559) <= not (a or b);
    layer1_outputs(560) <= not (a xor b);
    layer1_outputs(561) <= a and not b;
    layer1_outputs(562) <= not b;
    layer1_outputs(563) <= a xor b;
    layer1_outputs(564) <= not (a and b);
    layer1_outputs(565) <= not b;
    layer1_outputs(566) <= not (a and b);
    layer1_outputs(567) <= not a or b;
    layer1_outputs(568) <= not b or a;
    layer1_outputs(569) <= a;
    layer1_outputs(570) <= not b or a;
    layer1_outputs(571) <= not a;
    layer1_outputs(572) <= a and b;
    layer1_outputs(573) <= not b or a;
    layer1_outputs(574) <= 1'b0;
    layer1_outputs(575) <= not b or a;
    layer1_outputs(576) <= a and b;
    layer1_outputs(577) <= a and b;
    layer1_outputs(578) <= not (a and b);
    layer1_outputs(579) <= a and b;
    layer1_outputs(580) <= a;
    layer1_outputs(581) <= not b;
    layer1_outputs(582) <= a and not b;
    layer1_outputs(583) <= not b;
    layer1_outputs(584) <= b;
    layer1_outputs(585) <= a and not b;
    layer1_outputs(586) <= not (a and b);
    layer1_outputs(587) <= not a;
    layer1_outputs(588) <= b and not a;
    layer1_outputs(589) <= not (a xor b);
    layer1_outputs(590) <= a and b;
    layer1_outputs(591) <= not (a and b);
    layer1_outputs(592) <= a and b;
    layer1_outputs(593) <= not a;
    layer1_outputs(594) <= a or b;
    layer1_outputs(595) <= not b;
    layer1_outputs(596) <= not (a and b);
    layer1_outputs(597) <= b;
    layer1_outputs(598) <= a xor b;
    layer1_outputs(599) <= b and not a;
    layer1_outputs(600) <= not (a or b);
    layer1_outputs(601) <= not (a or b);
    layer1_outputs(602) <= not (a or b);
    layer1_outputs(603) <= a and b;
    layer1_outputs(604) <= b;
    layer1_outputs(605) <= a;
    layer1_outputs(606) <= not (a and b);
    layer1_outputs(607) <= a;
    layer1_outputs(608) <= not b or a;
    layer1_outputs(609) <= not b;
    layer1_outputs(610) <= not (a and b);
    layer1_outputs(611) <= a or b;
    layer1_outputs(612) <= a and b;
    layer1_outputs(613) <= b;
    layer1_outputs(614) <= not b or a;
    layer1_outputs(615) <= a and not b;
    layer1_outputs(616) <= b;
    layer1_outputs(617) <= not (a and b);
    layer1_outputs(618) <= a;
    layer1_outputs(619) <= b;
    layer1_outputs(620) <= a and b;
    layer1_outputs(621) <= not a;
    layer1_outputs(622) <= not (a or b);
    layer1_outputs(623) <= not a or b;
    layer1_outputs(624) <= a xor b;
    layer1_outputs(625) <= a;
    layer1_outputs(626) <= b;
    layer1_outputs(627) <= not (a xor b);
    layer1_outputs(628) <= not (a or b);
    layer1_outputs(629) <= not a or b;
    layer1_outputs(630) <= 1'b1;
    layer1_outputs(631) <= a and b;
    layer1_outputs(632) <= a and not b;
    layer1_outputs(633) <= not b or a;
    layer1_outputs(634) <= b;
    layer1_outputs(635) <= not b or a;
    layer1_outputs(636) <= b;
    layer1_outputs(637) <= not a or b;
    layer1_outputs(638) <= a and not b;
    layer1_outputs(639) <= not (a or b);
    layer1_outputs(640) <= a;
    layer1_outputs(641) <= not b;
    layer1_outputs(642) <= not (a xor b);
    layer1_outputs(643) <= not b or a;
    layer1_outputs(644) <= not b;
    layer1_outputs(645) <= not b;
    layer1_outputs(646) <= not a;
    layer1_outputs(647) <= not (a or b);
    layer1_outputs(648) <= not b;
    layer1_outputs(649) <= not (a xor b);
    layer1_outputs(650) <= a and b;
    layer1_outputs(651) <= not (a or b);
    layer1_outputs(652) <= b;
    layer1_outputs(653) <= not (a xor b);
    layer1_outputs(654) <= not b;
    layer1_outputs(655) <= not a;
    layer1_outputs(656) <= a;
    layer1_outputs(657) <= b;
    layer1_outputs(658) <= a and b;
    layer1_outputs(659) <= not b;
    layer1_outputs(660) <= not b;
    layer1_outputs(661) <= not a;
    layer1_outputs(662) <= a and b;
    layer1_outputs(663) <= not a;
    layer1_outputs(664) <= a and not b;
    layer1_outputs(665) <= b;
    layer1_outputs(666) <= not (a or b);
    layer1_outputs(667) <= a xor b;
    layer1_outputs(668) <= 1'b0;
    layer1_outputs(669) <= not (a or b);
    layer1_outputs(670) <= a;
    layer1_outputs(671) <= not (a xor b);
    layer1_outputs(672) <= b;
    layer1_outputs(673) <= b and not a;
    layer1_outputs(674) <= not b or a;
    layer1_outputs(675) <= a or b;
    layer1_outputs(676) <= a xor b;
    layer1_outputs(677) <= a and b;
    layer1_outputs(678) <= not a;
    layer1_outputs(679) <= a or b;
    layer1_outputs(680) <= a xor b;
    layer1_outputs(681) <= b;
    layer1_outputs(682) <= a;
    layer1_outputs(683) <= not b;
    layer1_outputs(684) <= a and b;
    layer1_outputs(685) <= not b;
    layer1_outputs(686) <= a and not b;
    layer1_outputs(687) <= not (a or b);
    layer1_outputs(688) <= a xor b;
    layer1_outputs(689) <= a xor b;
    layer1_outputs(690) <= not (a xor b);
    layer1_outputs(691) <= not b;
    layer1_outputs(692) <= not a;
    layer1_outputs(693) <= a and b;
    layer1_outputs(694) <= a xor b;
    layer1_outputs(695) <= b and not a;
    layer1_outputs(696) <= not (a or b);
    layer1_outputs(697) <= not (a and b);
    layer1_outputs(698) <= not (a xor b);
    layer1_outputs(699) <= a xor b;
    layer1_outputs(700) <= a xor b;
    layer1_outputs(701) <= a;
    layer1_outputs(702) <= a and b;
    layer1_outputs(703) <= not b;
    layer1_outputs(704) <= a or b;
    layer1_outputs(705) <= a;
    layer1_outputs(706) <= a and not b;
    layer1_outputs(707) <= not (a or b);
    layer1_outputs(708) <= not b or a;
    layer1_outputs(709) <= a;
    layer1_outputs(710) <= not (a or b);
    layer1_outputs(711) <= not a;
    layer1_outputs(712) <= not (a or b);
    layer1_outputs(713) <= not (a or b);
    layer1_outputs(714) <= not (a and b);
    layer1_outputs(715) <= b;
    layer1_outputs(716) <= not a or b;
    layer1_outputs(717) <= b;
    layer1_outputs(718) <= a xor b;
    layer1_outputs(719) <= a;
    layer1_outputs(720) <= b;
    layer1_outputs(721) <= not a or b;
    layer1_outputs(722) <= a;
    layer1_outputs(723) <= b and not a;
    layer1_outputs(724) <= not b or a;
    layer1_outputs(725) <= not (a xor b);
    layer1_outputs(726) <= not b or a;
    layer1_outputs(727) <= not b;
    layer1_outputs(728) <= not (a xor b);
    layer1_outputs(729) <= a and not b;
    layer1_outputs(730) <= not b;
    layer1_outputs(731) <= a and not b;
    layer1_outputs(732) <= a xor b;
    layer1_outputs(733) <= not a;
    layer1_outputs(734) <= not (a and b);
    layer1_outputs(735) <= a or b;
    layer1_outputs(736) <= a;
    layer1_outputs(737) <= not a or b;
    layer1_outputs(738) <= a or b;
    layer1_outputs(739) <= a or b;
    layer1_outputs(740) <= not b;
    layer1_outputs(741) <= a xor b;
    layer1_outputs(742) <= a or b;
    layer1_outputs(743) <= not a or b;
    layer1_outputs(744) <= not a;
    layer1_outputs(745) <= a;
    layer1_outputs(746) <= b;
    layer1_outputs(747) <= not (a or b);
    layer1_outputs(748) <= not b or a;
    layer1_outputs(749) <= not a;
    layer1_outputs(750) <= a;
    layer1_outputs(751) <= not a or b;
    layer1_outputs(752) <= a;
    layer1_outputs(753) <= not b or a;
    layer1_outputs(754) <= b and not a;
    layer1_outputs(755) <= a or b;
    layer1_outputs(756) <= 1'b1;
    layer1_outputs(757) <= a and b;
    layer1_outputs(758) <= not b or a;
    layer1_outputs(759) <= not a or b;
    layer1_outputs(760) <= b;
    layer1_outputs(761) <= not (a or b);
    layer1_outputs(762) <= not (a xor b);
    layer1_outputs(763) <= not b or a;
    layer1_outputs(764) <= not b or a;
    layer1_outputs(765) <= b;
    layer1_outputs(766) <= not a;
    layer1_outputs(767) <= a and b;
    layer1_outputs(768) <= a;
    layer1_outputs(769) <= a and b;
    layer1_outputs(770) <= not (a and b);
    layer1_outputs(771) <= not b;
    layer1_outputs(772) <= not a or b;
    layer1_outputs(773) <= not b;
    layer1_outputs(774) <= a;
    layer1_outputs(775) <= not b;
    layer1_outputs(776) <= b;
    layer1_outputs(777) <= b;
    layer1_outputs(778) <= not b or a;
    layer1_outputs(779) <= not b or a;
    layer1_outputs(780) <= not (a and b);
    layer1_outputs(781) <= not (a or b);
    layer1_outputs(782) <= not a;
    layer1_outputs(783) <= 1'b0;
    layer1_outputs(784) <= not a or b;
    layer1_outputs(785) <= not a or b;
    layer1_outputs(786) <= a and b;
    layer1_outputs(787) <= not a;
    layer1_outputs(788) <= a and b;
    layer1_outputs(789) <= 1'b1;
    layer1_outputs(790) <= a and b;
    layer1_outputs(791) <= not b or a;
    layer1_outputs(792) <= not (a or b);
    layer1_outputs(793) <= not (a xor b);
    layer1_outputs(794) <= not (a or b);
    layer1_outputs(795) <= not b;
    layer1_outputs(796) <= a or b;
    layer1_outputs(797) <= a or b;
    layer1_outputs(798) <= b;
    layer1_outputs(799) <= a xor b;
    layer1_outputs(800) <= not (a xor b);
    layer1_outputs(801) <= a or b;
    layer1_outputs(802) <= a and b;
    layer1_outputs(803) <= a;
    layer1_outputs(804) <= not b or a;
    layer1_outputs(805) <= a and not b;
    layer1_outputs(806) <= a xor b;
    layer1_outputs(807) <= not b;
    layer1_outputs(808) <= not a or b;
    layer1_outputs(809) <= not a;
    layer1_outputs(810) <= not b or a;
    layer1_outputs(811) <= a xor b;
    layer1_outputs(812) <= not a or b;
    layer1_outputs(813) <= not a;
    layer1_outputs(814) <= b;
    layer1_outputs(815) <= b;
    layer1_outputs(816) <= not a or b;
    layer1_outputs(817) <= not a or b;
    layer1_outputs(818) <= b;
    layer1_outputs(819) <= not a or b;
    layer1_outputs(820) <= b;
    layer1_outputs(821) <= 1'b1;
    layer1_outputs(822) <= not (a xor b);
    layer1_outputs(823) <= b and not a;
    layer1_outputs(824) <= b and not a;
    layer1_outputs(825) <= not a;
    layer1_outputs(826) <= a and b;
    layer1_outputs(827) <= a and not b;
    layer1_outputs(828) <= b;
    layer1_outputs(829) <= b and not a;
    layer1_outputs(830) <= not b;
    layer1_outputs(831) <= a and not b;
    layer1_outputs(832) <= not a or b;
    layer1_outputs(833) <= b;
    layer1_outputs(834) <= a or b;
    layer1_outputs(835) <= not (a or b);
    layer1_outputs(836) <= not (a and b);
    layer1_outputs(837) <= a xor b;
    layer1_outputs(838) <= 1'b0;
    layer1_outputs(839) <= not b;
    layer1_outputs(840) <= not b;
    layer1_outputs(841) <= not a;
    layer1_outputs(842) <= not (a and b);
    layer1_outputs(843) <= a or b;
    layer1_outputs(844) <= not a;
    layer1_outputs(845) <= not (a or b);
    layer1_outputs(846) <= not b;
    layer1_outputs(847) <= not a or b;
    layer1_outputs(848) <= a and not b;
    layer1_outputs(849) <= a or b;
    layer1_outputs(850) <= a;
    layer1_outputs(851) <= not (a xor b);
    layer1_outputs(852) <= a;
    layer1_outputs(853) <= b;
    layer1_outputs(854) <= not (a xor b);
    layer1_outputs(855) <= not a;
    layer1_outputs(856) <= not (a xor b);
    layer1_outputs(857) <= not (a and b);
    layer1_outputs(858) <= not (a xor b);
    layer1_outputs(859) <= not a;
    layer1_outputs(860) <= b;
    layer1_outputs(861) <= not (a and b);
    layer1_outputs(862) <= b and not a;
    layer1_outputs(863) <= not (a and b);
    layer1_outputs(864) <= a or b;
    layer1_outputs(865) <= b and not a;
    layer1_outputs(866) <= b;
    layer1_outputs(867) <= not (a and b);
    layer1_outputs(868) <= b and not a;
    layer1_outputs(869) <= not (a and b);
    layer1_outputs(870) <= a;
    layer1_outputs(871) <= a;
    layer1_outputs(872) <= not a or b;
    layer1_outputs(873) <= a xor b;
    layer1_outputs(874) <= a or b;
    layer1_outputs(875) <= not (a or b);
    layer1_outputs(876) <= not b;
    layer1_outputs(877) <= not (a and b);
    layer1_outputs(878) <= not (a xor b);
    layer1_outputs(879) <= a xor b;
    layer1_outputs(880) <= not (a xor b);
    layer1_outputs(881) <= a and not b;
    layer1_outputs(882) <= not b or a;
    layer1_outputs(883) <= not (a xor b);
    layer1_outputs(884) <= 1'b0;
    layer1_outputs(885) <= not b or a;
    layer1_outputs(886) <= a or b;
    layer1_outputs(887) <= not b;
    layer1_outputs(888) <= a xor b;
    layer1_outputs(889) <= not b;
    layer1_outputs(890) <= b;
    layer1_outputs(891) <= a;
    layer1_outputs(892) <= not a;
    layer1_outputs(893) <= not (a and b);
    layer1_outputs(894) <= not b or a;
    layer1_outputs(895) <= b;
    layer1_outputs(896) <= not a;
    layer1_outputs(897) <= not (a and b);
    layer1_outputs(898) <= a;
    layer1_outputs(899) <= not a;
    layer1_outputs(900) <= a xor b;
    layer1_outputs(901) <= a and b;
    layer1_outputs(902) <= a xor b;
    layer1_outputs(903) <= a and not b;
    layer1_outputs(904) <= not (a and b);
    layer1_outputs(905) <= 1'b0;
    layer1_outputs(906) <= not (a or b);
    layer1_outputs(907) <= a and b;
    layer1_outputs(908) <= b and not a;
    layer1_outputs(909) <= not (a xor b);
    layer1_outputs(910) <= not b or a;
    layer1_outputs(911) <= a;
    layer1_outputs(912) <= not (a xor b);
    layer1_outputs(913) <= not (a xor b);
    layer1_outputs(914) <= not (a xor b);
    layer1_outputs(915) <= not b;
    layer1_outputs(916) <= b and not a;
    layer1_outputs(917) <= not (a and b);
    layer1_outputs(918) <= b;
    layer1_outputs(919) <= not (a xor b);
    layer1_outputs(920) <= b and not a;
    layer1_outputs(921) <= not b or a;
    layer1_outputs(922) <= not (a xor b);
    layer1_outputs(923) <= b and not a;
    layer1_outputs(924) <= a and not b;
    layer1_outputs(925) <= b and not a;
    layer1_outputs(926) <= a xor b;
    layer1_outputs(927) <= not (a xor b);
    layer1_outputs(928) <= not b or a;
    layer1_outputs(929) <= a and not b;
    layer1_outputs(930) <= not b or a;
    layer1_outputs(931) <= a or b;
    layer1_outputs(932) <= a and b;
    layer1_outputs(933) <= a or b;
    layer1_outputs(934) <= not a;
    layer1_outputs(935) <= not (a or b);
    layer1_outputs(936) <= b and not a;
    layer1_outputs(937) <= b;
    layer1_outputs(938) <= not a;
    layer1_outputs(939) <= not b or a;
    layer1_outputs(940) <= a and b;
    layer1_outputs(941) <= not a;
    layer1_outputs(942) <= a and not b;
    layer1_outputs(943) <= not b or a;
    layer1_outputs(944) <= not b;
    layer1_outputs(945) <= not (a and b);
    layer1_outputs(946) <= a;
    layer1_outputs(947) <= not (a and b);
    layer1_outputs(948) <= a and not b;
    layer1_outputs(949) <= not (a xor b);
    layer1_outputs(950) <= a and not b;
    layer1_outputs(951) <= not b;
    layer1_outputs(952) <= b;
    layer1_outputs(953) <= not (a or b);
    layer1_outputs(954) <= a;
    layer1_outputs(955) <= a and not b;
    layer1_outputs(956) <= not b or a;
    layer1_outputs(957) <= not a or b;
    layer1_outputs(958) <= not (a and b);
    layer1_outputs(959) <= a and not b;
    layer1_outputs(960) <= not a;
    layer1_outputs(961) <= a and b;
    layer1_outputs(962) <= not b;
    layer1_outputs(963) <= a and not b;
    layer1_outputs(964) <= not a;
    layer1_outputs(965) <= b;
    layer1_outputs(966) <= b;
    layer1_outputs(967) <= not a;
    layer1_outputs(968) <= a xor b;
    layer1_outputs(969) <= b;
    layer1_outputs(970) <= a and not b;
    layer1_outputs(971) <= not b;
    layer1_outputs(972) <= not a or b;
    layer1_outputs(973) <= a or b;
    layer1_outputs(974) <= b and not a;
    layer1_outputs(975) <= not a;
    layer1_outputs(976) <= b and not a;
    layer1_outputs(977) <= not a or b;
    layer1_outputs(978) <= a;
    layer1_outputs(979) <= not b or a;
    layer1_outputs(980) <= a and b;
    layer1_outputs(981) <= a and not b;
    layer1_outputs(982) <= not b;
    layer1_outputs(983) <= not b;
    layer1_outputs(984) <= a and not b;
    layer1_outputs(985) <= a and not b;
    layer1_outputs(986) <= not (a xor b);
    layer1_outputs(987) <= a xor b;
    layer1_outputs(988) <= not (a or b);
    layer1_outputs(989) <= b and not a;
    layer1_outputs(990) <= not a;
    layer1_outputs(991) <= a xor b;
    layer1_outputs(992) <= not (a or b);
    layer1_outputs(993) <= not (a xor b);
    layer1_outputs(994) <= a and b;
    layer1_outputs(995) <= b;
    layer1_outputs(996) <= 1'b0;
    layer1_outputs(997) <= not (a xor b);
    layer1_outputs(998) <= not (a xor b);
    layer1_outputs(999) <= not a or b;
    layer1_outputs(1000) <= not (a xor b);
    layer1_outputs(1001) <= not b or a;
    layer1_outputs(1002) <= not b or a;
    layer1_outputs(1003) <= a xor b;
    layer1_outputs(1004) <= not a;
    layer1_outputs(1005) <= not b or a;
    layer1_outputs(1006) <= not a;
    layer1_outputs(1007) <= not b or a;
    layer1_outputs(1008) <= a and not b;
    layer1_outputs(1009) <= not (a xor b);
    layer1_outputs(1010) <= a;
    layer1_outputs(1011) <= a and b;
    layer1_outputs(1012) <= a and b;
    layer1_outputs(1013) <= not (a xor b);
    layer1_outputs(1014) <= b and not a;
    layer1_outputs(1015) <= a or b;
    layer1_outputs(1016) <= b and not a;
    layer1_outputs(1017) <= b and not a;
    layer1_outputs(1018) <= b and not a;
    layer1_outputs(1019) <= not a;
    layer1_outputs(1020) <= not a;
    layer1_outputs(1021) <= not a or b;
    layer1_outputs(1022) <= a or b;
    layer1_outputs(1023) <= a or b;
    layer1_outputs(1024) <= not (a or b);
    layer1_outputs(1025) <= not b or a;
    layer1_outputs(1026) <= not b or a;
    layer1_outputs(1027) <= not a;
    layer1_outputs(1028) <= a;
    layer1_outputs(1029) <= a xor b;
    layer1_outputs(1030) <= not a;
    layer1_outputs(1031) <= not a;
    layer1_outputs(1032) <= not a;
    layer1_outputs(1033) <= a or b;
    layer1_outputs(1034) <= not (a xor b);
    layer1_outputs(1035) <= not (a and b);
    layer1_outputs(1036) <= a and b;
    layer1_outputs(1037) <= a xor b;
    layer1_outputs(1038) <= b;
    layer1_outputs(1039) <= not b or a;
    layer1_outputs(1040) <= a;
    layer1_outputs(1041) <= a and not b;
    layer1_outputs(1042) <= a or b;
    layer1_outputs(1043) <= not a or b;
    layer1_outputs(1044) <= b;
    layer1_outputs(1045) <= a and not b;
    layer1_outputs(1046) <= a and not b;
    layer1_outputs(1047) <= not (a or b);
    layer1_outputs(1048) <= a;
    layer1_outputs(1049) <= a;
    layer1_outputs(1050) <= not b or a;
    layer1_outputs(1051) <= a and b;
    layer1_outputs(1052) <= not b or a;
    layer1_outputs(1053) <= b and not a;
    layer1_outputs(1054) <= not a;
    layer1_outputs(1055) <= not (a or b);
    layer1_outputs(1056) <= a and not b;
    layer1_outputs(1057) <= a xor b;
    layer1_outputs(1058) <= b;
    layer1_outputs(1059) <= not (a and b);
    layer1_outputs(1060) <= 1'b0;
    layer1_outputs(1061) <= not a;
    layer1_outputs(1062) <= a and not b;
    layer1_outputs(1063) <= not b;
    layer1_outputs(1064) <= a or b;
    layer1_outputs(1065) <= b and not a;
    layer1_outputs(1066) <= not a;
    layer1_outputs(1067) <= a and not b;
    layer1_outputs(1068) <= b and not a;
    layer1_outputs(1069) <= a and b;
    layer1_outputs(1070) <= a and b;
    layer1_outputs(1071) <= a and not b;
    layer1_outputs(1072) <= not b;
    layer1_outputs(1073) <= a xor b;
    layer1_outputs(1074) <= a;
    layer1_outputs(1075) <= not b or a;
    layer1_outputs(1076) <= not a;
    layer1_outputs(1077) <= b and not a;
    layer1_outputs(1078) <= b and not a;
    layer1_outputs(1079) <= b;
    layer1_outputs(1080) <= not a;
    layer1_outputs(1081) <= b;
    layer1_outputs(1082) <= not (a xor b);
    layer1_outputs(1083) <= a or b;
    layer1_outputs(1084) <= not a;
    layer1_outputs(1085) <= a;
    layer1_outputs(1086) <= not (a xor b);
    layer1_outputs(1087) <= not a or b;
    layer1_outputs(1088) <= a xor b;
    layer1_outputs(1089) <= not a;
    layer1_outputs(1090) <= not (a or b);
    layer1_outputs(1091) <= not (a and b);
    layer1_outputs(1092) <= not a or b;
    layer1_outputs(1093) <= a;
    layer1_outputs(1094) <= not (a and b);
    layer1_outputs(1095) <= not a;
    layer1_outputs(1096) <= not (a or b);
    layer1_outputs(1097) <= not (a and b);
    layer1_outputs(1098) <= a xor b;
    layer1_outputs(1099) <= not (a and b);
    layer1_outputs(1100) <= a xor b;
    layer1_outputs(1101) <= a and not b;
    layer1_outputs(1102) <= not b;
    layer1_outputs(1103) <= not a;
    layer1_outputs(1104) <= not a;
    layer1_outputs(1105) <= a and b;
    layer1_outputs(1106) <= not (a xor b);
    layer1_outputs(1107) <= b;
    layer1_outputs(1108) <= not (a xor b);
    layer1_outputs(1109) <= not b or a;
    layer1_outputs(1110) <= not (a xor b);
    layer1_outputs(1111) <= a or b;
    layer1_outputs(1112) <= a;
    layer1_outputs(1113) <= not b;
    layer1_outputs(1114) <= 1'b1;
    layer1_outputs(1115) <= a;
    layer1_outputs(1116) <= not b;
    layer1_outputs(1117) <= b;
    layer1_outputs(1118) <= 1'b1;
    layer1_outputs(1119) <= b and not a;
    layer1_outputs(1120) <= not b;
    layer1_outputs(1121) <= a and b;
    layer1_outputs(1122) <= not a or b;
    layer1_outputs(1123) <= not (a or b);
    layer1_outputs(1124) <= not a;
    layer1_outputs(1125) <= a;
    layer1_outputs(1126) <= not b;
    layer1_outputs(1127) <= not a;
    layer1_outputs(1128) <= a and not b;
    layer1_outputs(1129) <= 1'b1;
    layer1_outputs(1130) <= not b or a;
    layer1_outputs(1131) <= a;
    layer1_outputs(1132) <= not (a xor b);
    layer1_outputs(1133) <= a;
    layer1_outputs(1134) <= not (a xor b);
    layer1_outputs(1135) <= a or b;
    layer1_outputs(1136) <= not b or a;
    layer1_outputs(1137) <= not (a and b);
    layer1_outputs(1138) <= a and b;
    layer1_outputs(1139) <= a and not b;
    layer1_outputs(1140) <= a;
    layer1_outputs(1141) <= not a or b;
    layer1_outputs(1142) <= a and b;
    layer1_outputs(1143) <= 1'b1;
    layer1_outputs(1144) <= a;
    layer1_outputs(1145) <= not a or b;
    layer1_outputs(1146) <= a or b;
    layer1_outputs(1147) <= not (a or b);
    layer1_outputs(1148) <= not b or a;
    layer1_outputs(1149) <= b and not a;
    layer1_outputs(1150) <= a or b;
    layer1_outputs(1151) <= not a or b;
    layer1_outputs(1152) <= a;
    layer1_outputs(1153) <= a;
    layer1_outputs(1154) <= not a or b;
    layer1_outputs(1155) <= a and b;
    layer1_outputs(1156) <= not b;
    layer1_outputs(1157) <= not a;
    layer1_outputs(1158) <= not b or a;
    layer1_outputs(1159) <= not a;
    layer1_outputs(1160) <= a or b;
    layer1_outputs(1161) <= 1'b0;
    layer1_outputs(1162) <= not (a or b);
    layer1_outputs(1163) <= a xor b;
    layer1_outputs(1164) <= not b;
    layer1_outputs(1165) <= not b;
    layer1_outputs(1166) <= not b or a;
    layer1_outputs(1167) <= a xor b;
    layer1_outputs(1168) <= a;
    layer1_outputs(1169) <= a;
    layer1_outputs(1170) <= not (a xor b);
    layer1_outputs(1171) <= a and b;
    layer1_outputs(1172) <= a and not b;
    layer1_outputs(1173) <= not b;
    layer1_outputs(1174) <= not a or b;
    layer1_outputs(1175) <= not b;
    layer1_outputs(1176) <= a or b;
    layer1_outputs(1177) <= not b;
    layer1_outputs(1178) <= b;
    layer1_outputs(1179) <= not a or b;
    layer1_outputs(1180) <= a and not b;
    layer1_outputs(1181) <= a;
    layer1_outputs(1182) <= not (a xor b);
    layer1_outputs(1183) <= b;
    layer1_outputs(1184) <= a and b;
    layer1_outputs(1185) <= b;
    layer1_outputs(1186) <= b and not a;
    layer1_outputs(1187) <= not (a or b);
    layer1_outputs(1188) <= not b or a;
    layer1_outputs(1189) <= not a or b;
    layer1_outputs(1190) <= a xor b;
    layer1_outputs(1191) <= a or b;
    layer1_outputs(1192) <= a or b;
    layer1_outputs(1193) <= a and not b;
    layer1_outputs(1194) <= not a;
    layer1_outputs(1195) <= a;
    layer1_outputs(1196) <= a or b;
    layer1_outputs(1197) <= not a or b;
    layer1_outputs(1198) <= not b;
    layer1_outputs(1199) <= not a;
    layer1_outputs(1200) <= not b;
    layer1_outputs(1201) <= b;
    layer1_outputs(1202) <= not (a xor b);
    layer1_outputs(1203) <= b;
    layer1_outputs(1204) <= a and not b;
    layer1_outputs(1205) <= a xor b;
    layer1_outputs(1206) <= not a;
    layer1_outputs(1207) <= a and b;
    layer1_outputs(1208) <= not a;
    layer1_outputs(1209) <= not b;
    layer1_outputs(1210) <= b and not a;
    layer1_outputs(1211) <= not a;
    layer1_outputs(1212) <= a and not b;
    layer1_outputs(1213) <= not a;
    layer1_outputs(1214) <= a;
    layer1_outputs(1215) <= not a;
    layer1_outputs(1216) <= not a or b;
    layer1_outputs(1217) <= a;
    layer1_outputs(1218) <= a;
    layer1_outputs(1219) <= not a or b;
    layer1_outputs(1220) <= a and b;
    layer1_outputs(1221) <= a and not b;
    layer1_outputs(1222) <= a xor b;
    layer1_outputs(1223) <= not a;
    layer1_outputs(1224) <= not b;
    layer1_outputs(1225) <= not a;
    layer1_outputs(1226) <= a;
    layer1_outputs(1227) <= b and not a;
    layer1_outputs(1228) <= 1'b0;
    layer1_outputs(1229) <= a;
    layer1_outputs(1230) <= not b;
    layer1_outputs(1231) <= a and not b;
    layer1_outputs(1232) <= not (a and b);
    layer1_outputs(1233) <= not (a or b);
    layer1_outputs(1234) <= a;
    layer1_outputs(1235) <= a;
    layer1_outputs(1236) <= 1'b0;
    layer1_outputs(1237) <= not a;
    layer1_outputs(1238) <= not (a and b);
    layer1_outputs(1239) <= not b or a;
    layer1_outputs(1240) <= not b;
    layer1_outputs(1241) <= a and not b;
    layer1_outputs(1242) <= not b;
    layer1_outputs(1243) <= not (a or b);
    layer1_outputs(1244) <= not a or b;
    layer1_outputs(1245) <= a;
    layer1_outputs(1246) <= a and b;
    layer1_outputs(1247) <= a;
    layer1_outputs(1248) <= 1'b0;
    layer1_outputs(1249) <= not b;
    layer1_outputs(1250) <= a and b;
    layer1_outputs(1251) <= not b or a;
    layer1_outputs(1252) <= a xor b;
    layer1_outputs(1253) <= 1'b0;
    layer1_outputs(1254) <= not (a or b);
    layer1_outputs(1255) <= not (a xor b);
    layer1_outputs(1256) <= b;
    layer1_outputs(1257) <= a xor b;
    layer1_outputs(1258) <= a xor b;
    layer1_outputs(1259) <= not (a or b);
    layer1_outputs(1260) <= a xor b;
    layer1_outputs(1261) <= not (a or b);
    layer1_outputs(1262) <= a and not b;
    layer1_outputs(1263) <= not b;
    layer1_outputs(1264) <= a xor b;
    layer1_outputs(1265) <= not (a and b);
    layer1_outputs(1266) <= not a;
    layer1_outputs(1267) <= not a;
    layer1_outputs(1268) <= not (a xor b);
    layer1_outputs(1269) <= a;
    layer1_outputs(1270) <= not (a xor b);
    layer1_outputs(1271) <= not a;
    layer1_outputs(1272) <= a;
    layer1_outputs(1273) <= not b;
    layer1_outputs(1274) <= a;
    layer1_outputs(1275) <= a xor b;
    layer1_outputs(1276) <= b;
    layer1_outputs(1277) <= not (a and b);
    layer1_outputs(1278) <= a and b;
    layer1_outputs(1279) <= not b;
    layer1_outputs(1280) <= a xor b;
    layer1_outputs(1281) <= not b;
    layer1_outputs(1282) <= a and not b;
    layer1_outputs(1283) <= not a;
    layer1_outputs(1284) <= not b;
    layer1_outputs(1285) <= b and not a;
    layer1_outputs(1286) <= b;
    layer1_outputs(1287) <= not a;
    layer1_outputs(1288) <= not b;
    layer1_outputs(1289) <= b;
    layer1_outputs(1290) <= a;
    layer1_outputs(1291) <= b;
    layer1_outputs(1292) <= not (a xor b);
    layer1_outputs(1293) <= 1'b0;
    layer1_outputs(1294) <= not b or a;
    layer1_outputs(1295) <= a or b;
    layer1_outputs(1296) <= not b;
    layer1_outputs(1297) <= a;
    layer1_outputs(1298) <= b and not a;
    layer1_outputs(1299) <= not b or a;
    layer1_outputs(1300) <= b and not a;
    layer1_outputs(1301) <= not b;
    layer1_outputs(1302) <= b;
    layer1_outputs(1303) <= not b or a;
    layer1_outputs(1304) <= not (a and b);
    layer1_outputs(1305) <= not b;
    layer1_outputs(1306) <= not a;
    layer1_outputs(1307) <= not a or b;
    layer1_outputs(1308) <= not a or b;
    layer1_outputs(1309) <= not (a xor b);
    layer1_outputs(1310) <= not a or b;
    layer1_outputs(1311) <= not a;
    layer1_outputs(1312) <= b;
    layer1_outputs(1313) <= a;
    layer1_outputs(1314) <= not b;
    layer1_outputs(1315) <= b;
    layer1_outputs(1316) <= not a;
    layer1_outputs(1317) <= b and not a;
    layer1_outputs(1318) <= a;
    layer1_outputs(1319) <= not (a xor b);
    layer1_outputs(1320) <= not (a xor b);
    layer1_outputs(1321) <= not b;
    layer1_outputs(1322) <= not a or b;
    layer1_outputs(1323) <= a;
    layer1_outputs(1324) <= not b;
    layer1_outputs(1325) <= not a or b;
    layer1_outputs(1326) <= not (a xor b);
    layer1_outputs(1327) <= not (a or b);
    layer1_outputs(1328) <= not b;
    layer1_outputs(1329) <= b and not a;
    layer1_outputs(1330) <= not b;
    layer1_outputs(1331) <= not b;
    layer1_outputs(1332) <= b and not a;
    layer1_outputs(1333) <= not a;
    layer1_outputs(1334) <= a or b;
    layer1_outputs(1335) <= a or b;
    layer1_outputs(1336) <= not b or a;
    layer1_outputs(1337) <= not a or b;
    layer1_outputs(1338) <= not (a xor b);
    layer1_outputs(1339) <= a xor b;
    layer1_outputs(1340) <= a and b;
    layer1_outputs(1341) <= a;
    layer1_outputs(1342) <= not b or a;
    layer1_outputs(1343) <= not (a xor b);
    layer1_outputs(1344) <= not b or a;
    layer1_outputs(1345) <= not b or a;
    layer1_outputs(1346) <= not a;
    layer1_outputs(1347) <= not b;
    layer1_outputs(1348) <= not (a xor b);
    layer1_outputs(1349) <= a and not b;
    layer1_outputs(1350) <= b and not a;
    layer1_outputs(1351) <= not b or a;
    layer1_outputs(1352) <= not b;
    layer1_outputs(1353) <= not (a and b);
    layer1_outputs(1354) <= b;
    layer1_outputs(1355) <= b;
    layer1_outputs(1356) <= b and not a;
    layer1_outputs(1357) <= not a;
    layer1_outputs(1358) <= not (a and b);
    layer1_outputs(1359) <= not (a and b);
    layer1_outputs(1360) <= a and not b;
    layer1_outputs(1361) <= not b or a;
    layer1_outputs(1362) <= b and not a;
    layer1_outputs(1363) <= a or b;
    layer1_outputs(1364) <= a xor b;
    layer1_outputs(1365) <= a;
    layer1_outputs(1366) <= a;
    layer1_outputs(1367) <= not b or a;
    layer1_outputs(1368) <= not a;
    layer1_outputs(1369) <= b;
    layer1_outputs(1370) <= a;
    layer1_outputs(1371) <= b and not a;
    layer1_outputs(1372) <= not a;
    layer1_outputs(1373) <= not (a xor b);
    layer1_outputs(1374) <= not a;
    layer1_outputs(1375) <= b;
    layer1_outputs(1376) <= a and not b;
    layer1_outputs(1377) <= not b;
    layer1_outputs(1378) <= not b;
    layer1_outputs(1379) <= a and b;
    layer1_outputs(1380) <= not a;
    layer1_outputs(1381) <= b;
    layer1_outputs(1382) <= a and not b;
    layer1_outputs(1383) <= a and b;
    layer1_outputs(1384) <= not (a xor b);
    layer1_outputs(1385) <= b;
    layer1_outputs(1386) <= not b;
    layer1_outputs(1387) <= b and not a;
    layer1_outputs(1388) <= a and not b;
    layer1_outputs(1389) <= not b;
    layer1_outputs(1390) <= a xor b;
    layer1_outputs(1391) <= b;
    layer1_outputs(1392) <= not (a or b);
    layer1_outputs(1393) <= b and not a;
    layer1_outputs(1394) <= a xor b;
    layer1_outputs(1395) <= a xor b;
    layer1_outputs(1396) <= not b;
    layer1_outputs(1397) <= not b;
    layer1_outputs(1398) <= a or b;
    layer1_outputs(1399) <= not b;
    layer1_outputs(1400) <= not a or b;
    layer1_outputs(1401) <= b;
    layer1_outputs(1402) <= a or b;
    layer1_outputs(1403) <= b;
    layer1_outputs(1404) <= a and b;
    layer1_outputs(1405) <= a;
    layer1_outputs(1406) <= b and not a;
    layer1_outputs(1407) <= a;
    layer1_outputs(1408) <= b;
    layer1_outputs(1409) <= not b or a;
    layer1_outputs(1410) <= a;
    layer1_outputs(1411) <= not (a or b);
    layer1_outputs(1412) <= b and not a;
    layer1_outputs(1413) <= a and b;
    layer1_outputs(1414) <= not a or b;
    layer1_outputs(1415) <= not a or b;
    layer1_outputs(1416) <= a or b;
    layer1_outputs(1417) <= b and not a;
    layer1_outputs(1418) <= not a;
    layer1_outputs(1419) <= b and not a;
    layer1_outputs(1420) <= 1'b1;
    layer1_outputs(1421) <= a and b;
    layer1_outputs(1422) <= a xor b;
    layer1_outputs(1423) <= a and not b;
    layer1_outputs(1424) <= not (a or b);
    layer1_outputs(1425) <= a and not b;
    layer1_outputs(1426) <= 1'b1;
    layer1_outputs(1427) <= a and b;
    layer1_outputs(1428) <= a or b;
    layer1_outputs(1429) <= a;
    layer1_outputs(1430) <= a and b;
    layer1_outputs(1431) <= a or b;
    layer1_outputs(1432) <= a and not b;
    layer1_outputs(1433) <= a and b;
    layer1_outputs(1434) <= not (a xor b);
    layer1_outputs(1435) <= b;
    layer1_outputs(1436) <= not b;
    layer1_outputs(1437) <= a xor b;
    layer1_outputs(1438) <= b and not a;
    layer1_outputs(1439) <= not (a or b);
    layer1_outputs(1440) <= a and b;
    layer1_outputs(1441) <= not a or b;
    layer1_outputs(1442) <= b and not a;
    layer1_outputs(1443) <= not b or a;
    layer1_outputs(1444) <= not a or b;
    layer1_outputs(1445) <= b;
    layer1_outputs(1446) <= a and b;
    layer1_outputs(1447) <= a and b;
    layer1_outputs(1448) <= a;
    layer1_outputs(1449) <= a xor b;
    layer1_outputs(1450) <= 1'b0;
    layer1_outputs(1451) <= not a;
    layer1_outputs(1452) <= not a;
    layer1_outputs(1453) <= not (a and b);
    layer1_outputs(1454) <= not b;
    layer1_outputs(1455) <= b and not a;
    layer1_outputs(1456) <= b and not a;
    layer1_outputs(1457) <= not (a xor b);
    layer1_outputs(1458) <= not a;
    layer1_outputs(1459) <= not b;
    layer1_outputs(1460) <= a or b;
    layer1_outputs(1461) <= not b;
    layer1_outputs(1462) <= not (a xor b);
    layer1_outputs(1463) <= not b;
    layer1_outputs(1464) <= a and not b;
    layer1_outputs(1465) <= not (a or b);
    layer1_outputs(1466) <= not (a and b);
    layer1_outputs(1467) <= not a or b;
    layer1_outputs(1468) <= b;
    layer1_outputs(1469) <= a xor b;
    layer1_outputs(1470) <= not (a or b);
    layer1_outputs(1471) <= not a or b;
    layer1_outputs(1472) <= a and b;
    layer1_outputs(1473) <= b and not a;
    layer1_outputs(1474) <= a and b;
    layer1_outputs(1475) <= not b or a;
    layer1_outputs(1476) <= not a or b;
    layer1_outputs(1477) <= not (a xor b);
    layer1_outputs(1478) <= a xor b;
    layer1_outputs(1479) <= not (a xor b);
    layer1_outputs(1480) <= a;
    layer1_outputs(1481) <= not a or b;
    layer1_outputs(1482) <= b;
    layer1_outputs(1483) <= not b;
    layer1_outputs(1484) <= b;
    layer1_outputs(1485) <= not (a xor b);
    layer1_outputs(1486) <= not b;
    layer1_outputs(1487) <= b;
    layer1_outputs(1488) <= a and not b;
    layer1_outputs(1489) <= not (a or b);
    layer1_outputs(1490) <= not (a or b);
    layer1_outputs(1491) <= not b;
    layer1_outputs(1492) <= not b or a;
    layer1_outputs(1493) <= not (a and b);
    layer1_outputs(1494) <= not (a or b);
    layer1_outputs(1495) <= a and not b;
    layer1_outputs(1496) <= 1'b0;
    layer1_outputs(1497) <= not (a or b);
    layer1_outputs(1498) <= 1'b0;
    layer1_outputs(1499) <= a;
    layer1_outputs(1500) <= b and not a;
    layer1_outputs(1501) <= b and not a;
    layer1_outputs(1502) <= not (a xor b);
    layer1_outputs(1503) <= a xor b;
    layer1_outputs(1504) <= a xor b;
    layer1_outputs(1505) <= not (a or b);
    layer1_outputs(1506) <= b;
    layer1_outputs(1507) <= a;
    layer1_outputs(1508) <= not b;
    layer1_outputs(1509) <= b and not a;
    layer1_outputs(1510) <= a;
    layer1_outputs(1511) <= not b or a;
    layer1_outputs(1512) <= a;
    layer1_outputs(1513) <= not b;
    layer1_outputs(1514) <= not (a and b);
    layer1_outputs(1515) <= not b or a;
    layer1_outputs(1516) <= not b;
    layer1_outputs(1517) <= 1'b0;
    layer1_outputs(1518) <= not a or b;
    layer1_outputs(1519) <= not (a xor b);
    layer1_outputs(1520) <= not a or b;
    layer1_outputs(1521) <= not b;
    layer1_outputs(1522) <= not b;
    layer1_outputs(1523) <= not b;
    layer1_outputs(1524) <= a and not b;
    layer1_outputs(1525) <= not a;
    layer1_outputs(1526) <= not a or b;
    layer1_outputs(1527) <= a xor b;
    layer1_outputs(1528) <= not a or b;
    layer1_outputs(1529) <= b and not a;
    layer1_outputs(1530) <= b;
    layer1_outputs(1531) <= 1'b1;
    layer1_outputs(1532) <= a or b;
    layer1_outputs(1533) <= a and not b;
    layer1_outputs(1534) <= b;
    layer1_outputs(1535) <= not (a or b);
    layer1_outputs(1536) <= not b or a;
    layer1_outputs(1537) <= b and not a;
    layer1_outputs(1538) <= not b;
    layer1_outputs(1539) <= not b or a;
    layer1_outputs(1540) <= not b or a;
    layer1_outputs(1541) <= not (a and b);
    layer1_outputs(1542) <= not b;
    layer1_outputs(1543) <= not b;
    layer1_outputs(1544) <= a and not b;
    layer1_outputs(1545) <= not (a and b);
    layer1_outputs(1546) <= a or b;
    layer1_outputs(1547) <= a xor b;
    layer1_outputs(1548) <= a and b;
    layer1_outputs(1549) <= a;
    layer1_outputs(1550) <= a or b;
    layer1_outputs(1551) <= not (a or b);
    layer1_outputs(1552) <= not a;
    layer1_outputs(1553) <= not b or a;
    layer1_outputs(1554) <= a;
    layer1_outputs(1555) <= a xor b;
    layer1_outputs(1556) <= b;
    layer1_outputs(1557) <= not (a and b);
    layer1_outputs(1558) <= a;
    layer1_outputs(1559) <= b;
    layer1_outputs(1560) <= 1'b0;
    layer1_outputs(1561) <= not b or a;
    layer1_outputs(1562) <= not a or b;
    layer1_outputs(1563) <= not (a xor b);
    layer1_outputs(1564) <= a;
    layer1_outputs(1565) <= not a;
    layer1_outputs(1566) <= not b;
    layer1_outputs(1567) <= b;
    layer1_outputs(1568) <= not b;
    layer1_outputs(1569) <= not a or b;
    layer1_outputs(1570) <= a;
    layer1_outputs(1571) <= b;
    layer1_outputs(1572) <= a and b;
    layer1_outputs(1573) <= a and not b;
    layer1_outputs(1574) <= not a or b;
    layer1_outputs(1575) <= not a;
    layer1_outputs(1576) <= not b;
    layer1_outputs(1577) <= not b;
    layer1_outputs(1578) <= not (a and b);
    layer1_outputs(1579) <= not a;
    layer1_outputs(1580) <= a;
    layer1_outputs(1581) <= not a or b;
    layer1_outputs(1582) <= not (a xor b);
    layer1_outputs(1583) <= not (a xor b);
    layer1_outputs(1584) <= a and b;
    layer1_outputs(1585) <= b and not a;
    layer1_outputs(1586) <= not (a xor b);
    layer1_outputs(1587) <= 1'b1;
    layer1_outputs(1588) <= not b;
    layer1_outputs(1589) <= a and not b;
    layer1_outputs(1590) <= not a or b;
    layer1_outputs(1591) <= a xor b;
    layer1_outputs(1592) <= a and b;
    layer1_outputs(1593) <= a;
    layer1_outputs(1594) <= not a;
    layer1_outputs(1595) <= not (a or b);
    layer1_outputs(1596) <= b;
    layer1_outputs(1597) <= a or b;
    layer1_outputs(1598) <= b and not a;
    layer1_outputs(1599) <= a xor b;
    layer1_outputs(1600) <= a;
    layer1_outputs(1601) <= not b or a;
    layer1_outputs(1602) <= not a;
    layer1_outputs(1603) <= not a or b;
    layer1_outputs(1604) <= not (a and b);
    layer1_outputs(1605) <= a or b;
    layer1_outputs(1606) <= a xor b;
    layer1_outputs(1607) <= not (a and b);
    layer1_outputs(1608) <= not b;
    layer1_outputs(1609) <= a and not b;
    layer1_outputs(1610) <= a and b;
    layer1_outputs(1611) <= a or b;
    layer1_outputs(1612) <= not (a and b);
    layer1_outputs(1613) <= b;
    layer1_outputs(1614) <= not (a and b);
    layer1_outputs(1615) <= not (a and b);
    layer1_outputs(1616) <= b;
    layer1_outputs(1617) <= a or b;
    layer1_outputs(1618) <= b and not a;
    layer1_outputs(1619) <= a or b;
    layer1_outputs(1620) <= b;
    layer1_outputs(1621) <= not a;
    layer1_outputs(1622) <= a and b;
    layer1_outputs(1623) <= not b;
    layer1_outputs(1624) <= not a;
    layer1_outputs(1625) <= b;
    layer1_outputs(1626) <= not (a or b);
    layer1_outputs(1627) <= not (a and b);
    layer1_outputs(1628) <= not (a xor b);
    layer1_outputs(1629) <= not a or b;
    layer1_outputs(1630) <= a;
    layer1_outputs(1631) <= not a;
    layer1_outputs(1632) <= not (a xor b);
    layer1_outputs(1633) <= a;
    layer1_outputs(1634) <= a and b;
    layer1_outputs(1635) <= not (a and b);
    layer1_outputs(1636) <= b;
    layer1_outputs(1637) <= a and b;
    layer1_outputs(1638) <= a and not b;
    layer1_outputs(1639) <= not (a or b);
    layer1_outputs(1640) <= a or b;
    layer1_outputs(1641) <= a or b;
    layer1_outputs(1642) <= not b;
    layer1_outputs(1643) <= a and b;
    layer1_outputs(1644) <= a and not b;
    layer1_outputs(1645) <= a xor b;
    layer1_outputs(1646) <= a;
    layer1_outputs(1647) <= a;
    layer1_outputs(1648) <= not a;
    layer1_outputs(1649) <= not (a or b);
    layer1_outputs(1650) <= a;
    layer1_outputs(1651) <= b;
    layer1_outputs(1652) <= not a or b;
    layer1_outputs(1653) <= not (a and b);
    layer1_outputs(1654) <= not (a and b);
    layer1_outputs(1655) <= a;
    layer1_outputs(1656) <= not b or a;
    layer1_outputs(1657) <= a or b;
    layer1_outputs(1658) <= not a;
    layer1_outputs(1659) <= not b or a;
    layer1_outputs(1660) <= not (a xor b);
    layer1_outputs(1661) <= b;
    layer1_outputs(1662) <= a xor b;
    layer1_outputs(1663) <= not (a or b);
    layer1_outputs(1664) <= b and not a;
    layer1_outputs(1665) <= not a;
    layer1_outputs(1666) <= not a;
    layer1_outputs(1667) <= not a;
    layer1_outputs(1668) <= b and not a;
    layer1_outputs(1669) <= not a;
    layer1_outputs(1670) <= not a or b;
    layer1_outputs(1671) <= a;
    layer1_outputs(1672) <= not (a xor b);
    layer1_outputs(1673) <= a or b;
    layer1_outputs(1674) <= b;
    layer1_outputs(1675) <= not (a and b);
    layer1_outputs(1676) <= not a;
    layer1_outputs(1677) <= not a;
    layer1_outputs(1678) <= a and not b;
    layer1_outputs(1679) <= a xor b;
    layer1_outputs(1680) <= not b;
    layer1_outputs(1681) <= not (a xor b);
    layer1_outputs(1682) <= b and not a;
    layer1_outputs(1683) <= not b;
    layer1_outputs(1684) <= not a or b;
    layer1_outputs(1685) <= a and not b;
    layer1_outputs(1686) <= b and not a;
    layer1_outputs(1687) <= not a;
    layer1_outputs(1688) <= not b or a;
    layer1_outputs(1689) <= not b;
    layer1_outputs(1690) <= a;
    layer1_outputs(1691) <= a xor b;
    layer1_outputs(1692) <= not a;
    layer1_outputs(1693) <= a or b;
    layer1_outputs(1694) <= not (a and b);
    layer1_outputs(1695) <= b;
    layer1_outputs(1696) <= not b or a;
    layer1_outputs(1697) <= not b or a;
    layer1_outputs(1698) <= a xor b;
    layer1_outputs(1699) <= b;
    layer1_outputs(1700) <= not (a or b);
    layer1_outputs(1701) <= not a or b;
    layer1_outputs(1702) <= b and not a;
    layer1_outputs(1703) <= not (a xor b);
    layer1_outputs(1704) <= a;
    layer1_outputs(1705) <= a and b;
    layer1_outputs(1706) <= a;
    layer1_outputs(1707) <= not a;
    layer1_outputs(1708) <= a and not b;
    layer1_outputs(1709) <= a and b;
    layer1_outputs(1710) <= not a;
    layer1_outputs(1711) <= not a or b;
    layer1_outputs(1712) <= a xor b;
    layer1_outputs(1713) <= not b or a;
    layer1_outputs(1714) <= a and b;
    layer1_outputs(1715) <= a and b;
    layer1_outputs(1716) <= not a;
    layer1_outputs(1717) <= b and not a;
    layer1_outputs(1718) <= not b;
    layer1_outputs(1719) <= not (a or b);
    layer1_outputs(1720) <= a and b;
    layer1_outputs(1721) <= not b or a;
    layer1_outputs(1722) <= not a or b;
    layer1_outputs(1723) <= not b or a;
    layer1_outputs(1724) <= not a or b;
    layer1_outputs(1725) <= a;
    layer1_outputs(1726) <= not a or b;
    layer1_outputs(1727) <= a;
    layer1_outputs(1728) <= a;
    layer1_outputs(1729) <= not b;
    layer1_outputs(1730) <= a and b;
    layer1_outputs(1731) <= not b;
    layer1_outputs(1732) <= not a or b;
    layer1_outputs(1733) <= a or b;
    layer1_outputs(1734) <= b and not a;
    layer1_outputs(1735) <= a xor b;
    layer1_outputs(1736) <= b and not a;
    layer1_outputs(1737) <= not a;
    layer1_outputs(1738) <= a xor b;
    layer1_outputs(1739) <= not (a xor b);
    layer1_outputs(1740) <= not (a or b);
    layer1_outputs(1741) <= not b;
    layer1_outputs(1742) <= not a or b;
    layer1_outputs(1743) <= a and not b;
    layer1_outputs(1744) <= a;
    layer1_outputs(1745) <= a;
    layer1_outputs(1746) <= not a or b;
    layer1_outputs(1747) <= not a;
    layer1_outputs(1748) <= not a or b;
    layer1_outputs(1749) <= b;
    layer1_outputs(1750) <= a;
    layer1_outputs(1751) <= a or b;
    layer1_outputs(1752) <= a;
    layer1_outputs(1753) <= a;
    layer1_outputs(1754) <= not (a xor b);
    layer1_outputs(1755) <= a;
    layer1_outputs(1756) <= b and not a;
    layer1_outputs(1757) <= b and not a;
    layer1_outputs(1758) <= a;
    layer1_outputs(1759) <= not b;
    layer1_outputs(1760) <= a and not b;
    layer1_outputs(1761) <= not (a or b);
    layer1_outputs(1762) <= b;
    layer1_outputs(1763) <= b;
    layer1_outputs(1764) <= a and not b;
    layer1_outputs(1765) <= not b or a;
    layer1_outputs(1766) <= not a;
    layer1_outputs(1767) <= not (a or b);
    layer1_outputs(1768) <= a or b;
    layer1_outputs(1769) <= b;
    layer1_outputs(1770) <= not (a xor b);
    layer1_outputs(1771) <= a;
    layer1_outputs(1772) <= a or b;
    layer1_outputs(1773) <= not (a xor b);
    layer1_outputs(1774) <= a xor b;
    layer1_outputs(1775) <= not b;
    layer1_outputs(1776) <= not a;
    layer1_outputs(1777) <= a or b;
    layer1_outputs(1778) <= b;
    layer1_outputs(1779) <= b;
    layer1_outputs(1780) <= a and b;
    layer1_outputs(1781) <= not a;
    layer1_outputs(1782) <= not a;
    layer1_outputs(1783) <= a and not b;
    layer1_outputs(1784) <= not b or a;
    layer1_outputs(1785) <= a;
    layer1_outputs(1786) <= not b or a;
    layer1_outputs(1787) <= b;
    layer1_outputs(1788) <= a and b;
    layer1_outputs(1789) <= b and not a;
    layer1_outputs(1790) <= not a;
    layer1_outputs(1791) <= a and b;
    layer1_outputs(1792) <= not b;
    layer1_outputs(1793) <= b and not a;
    layer1_outputs(1794) <= not (a or b);
    layer1_outputs(1795) <= not (a xor b);
    layer1_outputs(1796) <= not a;
    layer1_outputs(1797) <= not (a xor b);
    layer1_outputs(1798) <= not (a or b);
    layer1_outputs(1799) <= b and not a;
    layer1_outputs(1800) <= not b;
    layer1_outputs(1801) <= a xor b;
    layer1_outputs(1802) <= a xor b;
    layer1_outputs(1803) <= not a;
    layer1_outputs(1804) <= b;
    layer1_outputs(1805) <= not b;
    layer1_outputs(1806) <= b and not a;
    layer1_outputs(1807) <= a;
    layer1_outputs(1808) <= not b or a;
    layer1_outputs(1809) <= not (a or b);
    layer1_outputs(1810) <= not a or b;
    layer1_outputs(1811) <= a xor b;
    layer1_outputs(1812) <= not (a and b);
    layer1_outputs(1813) <= not b or a;
    layer1_outputs(1814) <= a or b;
    layer1_outputs(1815) <= a xor b;
    layer1_outputs(1816) <= not a or b;
    layer1_outputs(1817) <= a or b;
    layer1_outputs(1818) <= b and not a;
    layer1_outputs(1819) <= a;
    layer1_outputs(1820) <= a;
    layer1_outputs(1821) <= a and not b;
    layer1_outputs(1822) <= not a or b;
    layer1_outputs(1823) <= a xor b;
    layer1_outputs(1824) <= a;
    layer1_outputs(1825) <= a and b;
    layer1_outputs(1826) <= a;
    layer1_outputs(1827) <= b;
    layer1_outputs(1828) <= a xor b;
    layer1_outputs(1829) <= b;
    layer1_outputs(1830) <= a xor b;
    layer1_outputs(1831) <= b;
    layer1_outputs(1832) <= a and b;
    layer1_outputs(1833) <= b and not a;
    layer1_outputs(1834) <= a and not b;
    layer1_outputs(1835) <= not a or b;
    layer1_outputs(1836) <= not a or b;
    layer1_outputs(1837) <= 1'b0;
    layer1_outputs(1838) <= not a;
    layer1_outputs(1839) <= not a;
    layer1_outputs(1840) <= a;
    layer1_outputs(1841) <= not (a xor b);
    layer1_outputs(1842) <= a xor b;
    layer1_outputs(1843) <= b and not a;
    layer1_outputs(1844) <= a xor b;
    layer1_outputs(1845) <= b and not a;
    layer1_outputs(1846) <= not b;
    layer1_outputs(1847) <= a xor b;
    layer1_outputs(1848) <= a;
    layer1_outputs(1849) <= a xor b;
    layer1_outputs(1850) <= a and not b;
    layer1_outputs(1851) <= not (a and b);
    layer1_outputs(1852) <= not (a xor b);
    layer1_outputs(1853) <= b;
    layer1_outputs(1854) <= not b or a;
    layer1_outputs(1855) <= b;
    layer1_outputs(1856) <= not a;
    layer1_outputs(1857) <= not b or a;
    layer1_outputs(1858) <= a;
    layer1_outputs(1859) <= not (a and b);
    layer1_outputs(1860) <= not a or b;
    layer1_outputs(1861) <= b;
    layer1_outputs(1862) <= a;
    layer1_outputs(1863) <= not a;
    layer1_outputs(1864) <= a and not b;
    layer1_outputs(1865) <= not b;
    layer1_outputs(1866) <= not (a and b);
    layer1_outputs(1867) <= a and b;
    layer1_outputs(1868) <= not (a xor b);
    layer1_outputs(1869) <= not b;
    layer1_outputs(1870) <= a;
    layer1_outputs(1871) <= not (a or b);
    layer1_outputs(1872) <= 1'b1;
    layer1_outputs(1873) <= not a;
    layer1_outputs(1874) <= a and b;
    layer1_outputs(1875) <= b;
    layer1_outputs(1876) <= a;
    layer1_outputs(1877) <= b and not a;
    layer1_outputs(1878) <= b;
    layer1_outputs(1879) <= not b or a;
    layer1_outputs(1880) <= not a or b;
    layer1_outputs(1881) <= not a or b;
    layer1_outputs(1882) <= not a or b;
    layer1_outputs(1883) <= not b;
    layer1_outputs(1884) <= not a;
    layer1_outputs(1885) <= not b;
    layer1_outputs(1886) <= not b or a;
    layer1_outputs(1887) <= not a;
    layer1_outputs(1888) <= a and b;
    layer1_outputs(1889) <= not a or b;
    layer1_outputs(1890) <= b;
    layer1_outputs(1891) <= b and not a;
    layer1_outputs(1892) <= a and not b;
    layer1_outputs(1893) <= a and not b;
    layer1_outputs(1894) <= not (a or b);
    layer1_outputs(1895) <= a xor b;
    layer1_outputs(1896) <= not b;
    layer1_outputs(1897) <= not a or b;
    layer1_outputs(1898) <= not a;
    layer1_outputs(1899) <= not (a and b);
    layer1_outputs(1900) <= a or b;
    layer1_outputs(1901) <= not a;
    layer1_outputs(1902) <= b;
    layer1_outputs(1903) <= not (a or b);
    layer1_outputs(1904) <= not b;
    layer1_outputs(1905) <= not b or a;
    layer1_outputs(1906) <= b;
    layer1_outputs(1907) <= not a or b;
    layer1_outputs(1908) <= a and b;
    layer1_outputs(1909) <= not a;
    layer1_outputs(1910) <= b;
    layer1_outputs(1911) <= not b or a;
    layer1_outputs(1912) <= a and b;
    layer1_outputs(1913) <= a or b;
    layer1_outputs(1914) <= a and not b;
    layer1_outputs(1915) <= b;
    layer1_outputs(1916) <= not (a and b);
    layer1_outputs(1917) <= a xor b;
    layer1_outputs(1918) <= b and not a;
    layer1_outputs(1919) <= b and not a;
    layer1_outputs(1920) <= not b;
    layer1_outputs(1921) <= not b or a;
    layer1_outputs(1922) <= a and b;
    layer1_outputs(1923) <= a or b;
    layer1_outputs(1924) <= not b or a;
    layer1_outputs(1925) <= not b;
    layer1_outputs(1926) <= a and b;
    layer1_outputs(1927) <= not b;
    layer1_outputs(1928) <= not (a and b);
    layer1_outputs(1929) <= not b or a;
    layer1_outputs(1930) <= a;
    layer1_outputs(1931) <= not b or a;
    layer1_outputs(1932) <= not a;
    layer1_outputs(1933) <= a and not b;
    layer1_outputs(1934) <= not (a or b);
    layer1_outputs(1935) <= a or b;
    layer1_outputs(1936) <= not (a and b);
    layer1_outputs(1937) <= not (a or b);
    layer1_outputs(1938) <= a;
    layer1_outputs(1939) <= a xor b;
    layer1_outputs(1940) <= not b;
    layer1_outputs(1941) <= a;
    layer1_outputs(1942) <= b;
    layer1_outputs(1943) <= a and not b;
    layer1_outputs(1944) <= not a or b;
    layer1_outputs(1945) <= not (a xor b);
    layer1_outputs(1946) <= not b;
    layer1_outputs(1947) <= not (a xor b);
    layer1_outputs(1948) <= a or b;
    layer1_outputs(1949) <= not b or a;
    layer1_outputs(1950) <= b;
    layer1_outputs(1951) <= a or b;
    layer1_outputs(1952) <= b and not a;
    layer1_outputs(1953) <= a or b;
    layer1_outputs(1954) <= a and not b;
    layer1_outputs(1955) <= not (a and b);
    layer1_outputs(1956) <= not a or b;
    layer1_outputs(1957) <= a xor b;
    layer1_outputs(1958) <= not a or b;
    layer1_outputs(1959) <= b;
    layer1_outputs(1960) <= b;
    layer1_outputs(1961) <= not a;
    layer1_outputs(1962) <= not b or a;
    layer1_outputs(1963) <= 1'b1;
    layer1_outputs(1964) <= b and not a;
    layer1_outputs(1965) <= not a or b;
    layer1_outputs(1966) <= not b or a;
    layer1_outputs(1967) <= a or b;
    layer1_outputs(1968) <= a xor b;
    layer1_outputs(1969) <= not a or b;
    layer1_outputs(1970) <= not b;
    layer1_outputs(1971) <= a or b;
    layer1_outputs(1972) <= a and b;
    layer1_outputs(1973) <= not a;
    layer1_outputs(1974) <= a and b;
    layer1_outputs(1975) <= a and not b;
    layer1_outputs(1976) <= a and b;
    layer1_outputs(1977) <= a and not b;
    layer1_outputs(1978) <= not a;
    layer1_outputs(1979) <= not a or b;
    layer1_outputs(1980) <= not (a xor b);
    layer1_outputs(1981) <= a or b;
    layer1_outputs(1982) <= a xor b;
    layer1_outputs(1983) <= not a;
    layer1_outputs(1984) <= not (a xor b);
    layer1_outputs(1985) <= not b or a;
    layer1_outputs(1986) <= b;
    layer1_outputs(1987) <= not (a or b);
    layer1_outputs(1988) <= a or b;
    layer1_outputs(1989) <= b;
    layer1_outputs(1990) <= a xor b;
    layer1_outputs(1991) <= not a;
    layer1_outputs(1992) <= a;
    layer1_outputs(1993) <= not (a xor b);
    layer1_outputs(1994) <= a and not b;
    layer1_outputs(1995) <= not b;
    layer1_outputs(1996) <= a and not b;
    layer1_outputs(1997) <= a xor b;
    layer1_outputs(1998) <= not b;
    layer1_outputs(1999) <= not (a or b);
    layer1_outputs(2000) <= not (a or b);
    layer1_outputs(2001) <= not (a xor b);
    layer1_outputs(2002) <= not b or a;
    layer1_outputs(2003) <= b and not a;
    layer1_outputs(2004) <= b;
    layer1_outputs(2005) <= a and b;
    layer1_outputs(2006) <= not (a and b);
    layer1_outputs(2007) <= a and b;
    layer1_outputs(2008) <= a and b;
    layer1_outputs(2009) <= not (a or b);
    layer1_outputs(2010) <= not a;
    layer1_outputs(2011) <= a or b;
    layer1_outputs(2012) <= a;
    layer1_outputs(2013) <= not (a xor b);
    layer1_outputs(2014) <= b;
    layer1_outputs(2015) <= not a or b;
    layer1_outputs(2016) <= not b or a;
    layer1_outputs(2017) <= not (a or b);
    layer1_outputs(2018) <= a and not b;
    layer1_outputs(2019) <= not a;
    layer1_outputs(2020) <= not b;
    layer1_outputs(2021) <= a;
    layer1_outputs(2022) <= b;
    layer1_outputs(2023) <= not a or b;
    layer1_outputs(2024) <= not a;
    layer1_outputs(2025) <= a or b;
    layer1_outputs(2026) <= b;
    layer1_outputs(2027) <= a xor b;
    layer1_outputs(2028) <= not a;
    layer1_outputs(2029) <= not a or b;
    layer1_outputs(2030) <= not b;
    layer1_outputs(2031) <= not (a or b);
    layer1_outputs(2032) <= not (a or b);
    layer1_outputs(2033) <= b;
    layer1_outputs(2034) <= a and not b;
    layer1_outputs(2035) <= a;
    layer1_outputs(2036) <= a;
    layer1_outputs(2037) <= a and b;
    layer1_outputs(2038) <= not a or b;
    layer1_outputs(2039) <= not (a xor b);
    layer1_outputs(2040) <= not b or a;
    layer1_outputs(2041) <= b;
    layer1_outputs(2042) <= a and b;
    layer1_outputs(2043) <= b;
    layer1_outputs(2044) <= not b;
    layer1_outputs(2045) <= a and not b;
    layer1_outputs(2046) <= not b or a;
    layer1_outputs(2047) <= a;
    layer1_outputs(2048) <= not (a xor b);
    layer1_outputs(2049) <= a xor b;
    layer1_outputs(2050) <= not b or a;
    layer1_outputs(2051) <= not a;
    layer1_outputs(2052) <= a;
    layer1_outputs(2053) <= a and b;
    layer1_outputs(2054) <= not b;
    layer1_outputs(2055) <= a and b;
    layer1_outputs(2056) <= not (a or b);
    layer1_outputs(2057) <= b and not a;
    layer1_outputs(2058) <= not (a and b);
    layer1_outputs(2059) <= a and b;
    layer1_outputs(2060) <= not a or b;
    layer1_outputs(2061) <= a and b;
    layer1_outputs(2062) <= b and not a;
    layer1_outputs(2063) <= a;
    layer1_outputs(2064) <= b;
    layer1_outputs(2065) <= not b or a;
    layer1_outputs(2066) <= a xor b;
    layer1_outputs(2067) <= not (a or b);
    layer1_outputs(2068) <= not b;
    layer1_outputs(2069) <= b and not a;
    layer1_outputs(2070) <= not b;
    layer1_outputs(2071) <= b;
    layer1_outputs(2072) <= not (a or b);
    layer1_outputs(2073) <= b;
    layer1_outputs(2074) <= b and not a;
    layer1_outputs(2075) <= a or b;
    layer1_outputs(2076) <= not (a or b);
    layer1_outputs(2077) <= not (a and b);
    layer1_outputs(2078) <= not b or a;
    layer1_outputs(2079) <= not a;
    layer1_outputs(2080) <= not (a or b);
    layer1_outputs(2081) <= not (a or b);
    layer1_outputs(2082) <= not a or b;
    layer1_outputs(2083) <= not a or b;
    layer1_outputs(2084) <= not a;
    layer1_outputs(2085) <= a;
    layer1_outputs(2086) <= a and not b;
    layer1_outputs(2087) <= a and not b;
    layer1_outputs(2088) <= not (a or b);
    layer1_outputs(2089) <= 1'b1;
    layer1_outputs(2090) <= a;
    layer1_outputs(2091) <= not (a or b);
    layer1_outputs(2092) <= not a or b;
    layer1_outputs(2093) <= not a;
    layer1_outputs(2094) <= 1'b0;
    layer1_outputs(2095) <= b;
    layer1_outputs(2096) <= not b;
    layer1_outputs(2097) <= not b or a;
    layer1_outputs(2098) <= not b;
    layer1_outputs(2099) <= not (a or b);
    layer1_outputs(2100) <= a and b;
    layer1_outputs(2101) <= not a or b;
    layer1_outputs(2102) <= a and b;
    layer1_outputs(2103) <= not a;
    layer1_outputs(2104) <= b;
    layer1_outputs(2105) <= a;
    layer1_outputs(2106) <= b;
    layer1_outputs(2107) <= a xor b;
    layer1_outputs(2108) <= not b;
    layer1_outputs(2109) <= not b;
    layer1_outputs(2110) <= a and b;
    layer1_outputs(2111) <= not b;
    layer1_outputs(2112) <= not (a xor b);
    layer1_outputs(2113) <= a and b;
    layer1_outputs(2114) <= not (a or b);
    layer1_outputs(2115) <= a and b;
    layer1_outputs(2116) <= b;
    layer1_outputs(2117) <= b;
    layer1_outputs(2118) <= b and not a;
    layer1_outputs(2119) <= not (a and b);
    layer1_outputs(2120) <= not a;
    layer1_outputs(2121) <= not a or b;
    layer1_outputs(2122) <= b and not a;
    layer1_outputs(2123) <= not a or b;
    layer1_outputs(2124) <= not b;
    layer1_outputs(2125) <= b;
    layer1_outputs(2126) <= a xor b;
    layer1_outputs(2127) <= not b or a;
    layer1_outputs(2128) <= b;
    layer1_outputs(2129) <= not b;
    layer1_outputs(2130) <= b;
    layer1_outputs(2131) <= 1'b0;
    layer1_outputs(2132) <= a and not b;
    layer1_outputs(2133) <= a or b;
    layer1_outputs(2134) <= a;
    layer1_outputs(2135) <= a and not b;
    layer1_outputs(2136) <= b;
    layer1_outputs(2137) <= b and not a;
    layer1_outputs(2138) <= not (a xor b);
    layer1_outputs(2139) <= not a;
    layer1_outputs(2140) <= a and not b;
    layer1_outputs(2141) <= a and b;
    layer1_outputs(2142) <= not a;
    layer1_outputs(2143) <= a and b;
    layer1_outputs(2144) <= not a or b;
    layer1_outputs(2145) <= a xor b;
    layer1_outputs(2146) <= not b;
    layer1_outputs(2147) <= not (a or b);
    layer1_outputs(2148) <= a or b;
    layer1_outputs(2149) <= not b;
    layer1_outputs(2150) <= a;
    layer1_outputs(2151) <= not b;
    layer1_outputs(2152) <= not a;
    layer1_outputs(2153) <= not b;
    layer1_outputs(2154) <= not (a xor b);
    layer1_outputs(2155) <= not (a xor b);
    layer1_outputs(2156) <= b;
    layer1_outputs(2157) <= a and b;
    layer1_outputs(2158) <= b;
    layer1_outputs(2159) <= not b;
    layer1_outputs(2160) <= not a or b;
    layer1_outputs(2161) <= b;
    layer1_outputs(2162) <= not a;
    layer1_outputs(2163) <= a and not b;
    layer1_outputs(2164) <= a and b;
    layer1_outputs(2165) <= 1'b1;
    layer1_outputs(2166) <= b;
    layer1_outputs(2167) <= not (a xor b);
    layer1_outputs(2168) <= b;
    layer1_outputs(2169) <= b and not a;
    layer1_outputs(2170) <= a and not b;
    layer1_outputs(2171) <= not b;
    layer1_outputs(2172) <= a xor b;
    layer1_outputs(2173) <= not a or b;
    layer1_outputs(2174) <= 1'b0;
    layer1_outputs(2175) <= a or b;
    layer1_outputs(2176) <= b;
    layer1_outputs(2177) <= b and not a;
    layer1_outputs(2178) <= b;
    layer1_outputs(2179) <= not a;
    layer1_outputs(2180) <= not a;
    layer1_outputs(2181) <= not (a xor b);
    layer1_outputs(2182) <= a;
    layer1_outputs(2183) <= not (a or b);
    layer1_outputs(2184) <= not b or a;
    layer1_outputs(2185) <= a xor b;
    layer1_outputs(2186) <= a and b;
    layer1_outputs(2187) <= not a or b;
    layer1_outputs(2188) <= not b;
    layer1_outputs(2189) <= not (a xor b);
    layer1_outputs(2190) <= a xor b;
    layer1_outputs(2191) <= not b;
    layer1_outputs(2192) <= not a or b;
    layer1_outputs(2193) <= b and not a;
    layer1_outputs(2194) <= not b or a;
    layer1_outputs(2195) <= not a;
    layer1_outputs(2196) <= not (a and b);
    layer1_outputs(2197) <= a xor b;
    layer1_outputs(2198) <= not b or a;
    layer1_outputs(2199) <= not a;
    layer1_outputs(2200) <= not a or b;
    layer1_outputs(2201) <= b;
    layer1_outputs(2202) <= b and not a;
    layer1_outputs(2203) <= a and b;
    layer1_outputs(2204) <= a and b;
    layer1_outputs(2205) <= not b or a;
    layer1_outputs(2206) <= a and b;
    layer1_outputs(2207) <= not a or b;
    layer1_outputs(2208) <= a and not b;
    layer1_outputs(2209) <= not b;
    layer1_outputs(2210) <= a and not b;
    layer1_outputs(2211) <= not (a or b);
    layer1_outputs(2212) <= a;
    layer1_outputs(2213) <= a;
    layer1_outputs(2214) <= b;
    layer1_outputs(2215) <= a and not b;
    layer1_outputs(2216) <= not b;
    layer1_outputs(2217) <= not b;
    layer1_outputs(2218) <= not (a or b);
    layer1_outputs(2219) <= not b or a;
    layer1_outputs(2220) <= not (a xor b);
    layer1_outputs(2221) <= not b or a;
    layer1_outputs(2222) <= not b or a;
    layer1_outputs(2223) <= a xor b;
    layer1_outputs(2224) <= a or b;
    layer1_outputs(2225) <= a;
    layer1_outputs(2226) <= a xor b;
    layer1_outputs(2227) <= a;
    layer1_outputs(2228) <= not (a xor b);
    layer1_outputs(2229) <= b and not a;
    layer1_outputs(2230) <= a;
    layer1_outputs(2231) <= b and not a;
    layer1_outputs(2232) <= not a;
    layer1_outputs(2233) <= a;
    layer1_outputs(2234) <= a and not b;
    layer1_outputs(2235) <= not (a or b);
    layer1_outputs(2236) <= a and b;
    layer1_outputs(2237) <= a and not b;
    layer1_outputs(2238) <= a and b;
    layer1_outputs(2239) <= not (a and b);
    layer1_outputs(2240) <= a;
    layer1_outputs(2241) <= a xor b;
    layer1_outputs(2242) <= not a;
    layer1_outputs(2243) <= a and not b;
    layer1_outputs(2244) <= a;
    layer1_outputs(2245) <= not b;
    layer1_outputs(2246) <= b and not a;
    layer1_outputs(2247) <= a or b;
    layer1_outputs(2248) <= not b;
    layer1_outputs(2249) <= not b or a;
    layer1_outputs(2250) <= not b or a;
    layer1_outputs(2251) <= a or b;
    layer1_outputs(2252) <= not a or b;
    layer1_outputs(2253) <= not b;
    layer1_outputs(2254) <= b;
    layer1_outputs(2255) <= not (a xor b);
    layer1_outputs(2256) <= not a;
    layer1_outputs(2257) <= not b;
    layer1_outputs(2258) <= a and b;
    layer1_outputs(2259) <= not b or a;
    layer1_outputs(2260) <= a or b;
    layer1_outputs(2261) <= b;
    layer1_outputs(2262) <= b and not a;
    layer1_outputs(2263) <= b;
    layer1_outputs(2264) <= not b;
    layer1_outputs(2265) <= not b or a;
    layer1_outputs(2266) <= a;
    layer1_outputs(2267) <= a or b;
    layer1_outputs(2268) <= 1'b1;
    layer1_outputs(2269) <= a;
    layer1_outputs(2270) <= a and not b;
    layer1_outputs(2271) <= b;
    layer1_outputs(2272) <= a and not b;
    layer1_outputs(2273) <= not (a or b);
    layer1_outputs(2274) <= a;
    layer1_outputs(2275) <= b;
    layer1_outputs(2276) <= a and not b;
    layer1_outputs(2277) <= b and not a;
    layer1_outputs(2278) <= a xor b;
    layer1_outputs(2279) <= not (a and b);
    layer1_outputs(2280) <= not (a xor b);
    layer1_outputs(2281) <= a xor b;
    layer1_outputs(2282) <= not a;
    layer1_outputs(2283) <= a or b;
    layer1_outputs(2284) <= a and b;
    layer1_outputs(2285) <= not (a or b);
    layer1_outputs(2286) <= not (a or b);
    layer1_outputs(2287) <= not a;
    layer1_outputs(2288) <= a or b;
    layer1_outputs(2289) <= a and b;
    layer1_outputs(2290) <= a or b;
    layer1_outputs(2291) <= a or b;
    layer1_outputs(2292) <= a and not b;
    layer1_outputs(2293) <= not a or b;
    layer1_outputs(2294) <= a and not b;
    layer1_outputs(2295) <= not b or a;
    layer1_outputs(2296) <= not (a xor b);
    layer1_outputs(2297) <= not a;
    layer1_outputs(2298) <= a and b;
    layer1_outputs(2299) <= a xor b;
    layer1_outputs(2300) <= b;
    layer1_outputs(2301) <= not b;
    layer1_outputs(2302) <= b;
    layer1_outputs(2303) <= not (a xor b);
    layer1_outputs(2304) <= a xor b;
    layer1_outputs(2305) <= not b or a;
    layer1_outputs(2306) <= b and not a;
    layer1_outputs(2307) <= 1'b1;
    layer1_outputs(2308) <= not b;
    layer1_outputs(2309) <= not a or b;
    layer1_outputs(2310) <= b;
    layer1_outputs(2311) <= b;
    layer1_outputs(2312) <= not (a and b);
    layer1_outputs(2313) <= a xor b;
    layer1_outputs(2314) <= a and b;
    layer1_outputs(2315) <= b and not a;
    layer1_outputs(2316) <= not a or b;
    layer1_outputs(2317) <= not b or a;
    layer1_outputs(2318) <= b;
    layer1_outputs(2319) <= a;
    layer1_outputs(2320) <= not (a and b);
    layer1_outputs(2321) <= not b or a;
    layer1_outputs(2322) <= not (a and b);
    layer1_outputs(2323) <= a and not b;
    layer1_outputs(2324) <= not b;
    layer1_outputs(2325) <= a xor b;
    layer1_outputs(2326) <= not (a or b);
    layer1_outputs(2327) <= a or b;
    layer1_outputs(2328) <= b;
    layer1_outputs(2329) <= a and not b;
    layer1_outputs(2330) <= a and not b;
    layer1_outputs(2331) <= a;
    layer1_outputs(2332) <= not (a or b);
    layer1_outputs(2333) <= a or b;
    layer1_outputs(2334) <= not b;
    layer1_outputs(2335) <= not b;
    layer1_outputs(2336) <= a xor b;
    layer1_outputs(2337) <= a and not b;
    layer1_outputs(2338) <= a;
    layer1_outputs(2339) <= a and b;
    layer1_outputs(2340) <= not a;
    layer1_outputs(2341) <= not b or a;
    layer1_outputs(2342) <= not (a or b);
    layer1_outputs(2343) <= b and not a;
    layer1_outputs(2344) <= b;
    layer1_outputs(2345) <= b;
    layer1_outputs(2346) <= not b or a;
    layer1_outputs(2347) <= not b;
    layer1_outputs(2348) <= not b or a;
    layer1_outputs(2349) <= a and not b;
    layer1_outputs(2350) <= not b or a;
    layer1_outputs(2351) <= not (a or b);
    layer1_outputs(2352) <= a;
    layer1_outputs(2353) <= not a;
    layer1_outputs(2354) <= b and not a;
    layer1_outputs(2355) <= a;
    layer1_outputs(2356) <= a and b;
    layer1_outputs(2357) <= not a;
    layer1_outputs(2358) <= not b;
    layer1_outputs(2359) <= a and not b;
    layer1_outputs(2360) <= a and not b;
    layer1_outputs(2361) <= not b;
    layer1_outputs(2362) <= b;
    layer1_outputs(2363) <= a and not b;
    layer1_outputs(2364) <= b;
    layer1_outputs(2365) <= not (a or b);
    layer1_outputs(2366) <= a and not b;
    layer1_outputs(2367) <= not (a xor b);
    layer1_outputs(2368) <= b;
    layer1_outputs(2369) <= a;
    layer1_outputs(2370) <= a or b;
    layer1_outputs(2371) <= not (a and b);
    layer1_outputs(2372) <= a or b;
    layer1_outputs(2373) <= not a;
    layer1_outputs(2374) <= a and not b;
    layer1_outputs(2375) <= a or b;
    layer1_outputs(2376) <= b;
    layer1_outputs(2377) <= a;
    layer1_outputs(2378) <= a xor b;
    layer1_outputs(2379) <= a or b;
    layer1_outputs(2380) <= not (a xor b);
    layer1_outputs(2381) <= a or b;
    layer1_outputs(2382) <= 1'b0;
    layer1_outputs(2383) <= a or b;
    layer1_outputs(2384) <= b and not a;
    layer1_outputs(2385) <= not b;
    layer1_outputs(2386) <= a or b;
    layer1_outputs(2387) <= b;
    layer1_outputs(2388) <= not b;
    layer1_outputs(2389) <= a;
    layer1_outputs(2390) <= not (a xor b);
    layer1_outputs(2391) <= b and not a;
    layer1_outputs(2392) <= not (a and b);
    layer1_outputs(2393) <= a;
    layer1_outputs(2394) <= not a;
    layer1_outputs(2395) <= b;
    layer1_outputs(2396) <= a and b;
    layer1_outputs(2397) <= not b or a;
    layer1_outputs(2398) <= b;
    layer1_outputs(2399) <= b;
    layer1_outputs(2400) <= a;
    layer1_outputs(2401) <= a xor b;
    layer1_outputs(2402) <= a or b;
    layer1_outputs(2403) <= not a;
    layer1_outputs(2404) <= b and not a;
    layer1_outputs(2405) <= not b;
    layer1_outputs(2406) <= not b or a;
    layer1_outputs(2407) <= not a;
    layer1_outputs(2408) <= not (a xor b);
    layer1_outputs(2409) <= not (a or b);
    layer1_outputs(2410) <= a and not b;
    layer1_outputs(2411) <= not b;
    layer1_outputs(2412) <= a or b;
    layer1_outputs(2413) <= 1'b1;
    layer1_outputs(2414) <= b and not a;
    layer1_outputs(2415) <= not a or b;
    layer1_outputs(2416) <= not b;
    layer1_outputs(2417) <= not (a xor b);
    layer1_outputs(2418) <= not (a and b);
    layer1_outputs(2419) <= b and not a;
    layer1_outputs(2420) <= a;
    layer1_outputs(2421) <= b and not a;
    layer1_outputs(2422) <= not (a xor b);
    layer1_outputs(2423) <= a and not b;
    layer1_outputs(2424) <= a or b;
    layer1_outputs(2425) <= not b;
    layer1_outputs(2426) <= not (a or b);
    layer1_outputs(2427) <= b;
    layer1_outputs(2428) <= a and not b;
    layer1_outputs(2429) <= not (a xor b);
    layer1_outputs(2430) <= a and not b;
    layer1_outputs(2431) <= b and not a;
    layer1_outputs(2432) <= 1'b0;
    layer1_outputs(2433) <= not b;
    layer1_outputs(2434) <= not a or b;
    layer1_outputs(2435) <= a;
    layer1_outputs(2436) <= not (a and b);
    layer1_outputs(2437) <= a and not b;
    layer1_outputs(2438) <= not (a or b);
    layer1_outputs(2439) <= a xor b;
    layer1_outputs(2440) <= a xor b;
    layer1_outputs(2441) <= not (a and b);
    layer1_outputs(2442) <= not b or a;
    layer1_outputs(2443) <= b;
    layer1_outputs(2444) <= a and b;
    layer1_outputs(2445) <= not a or b;
    layer1_outputs(2446) <= b and not a;
    layer1_outputs(2447) <= a xor b;
    layer1_outputs(2448) <= a and not b;
    layer1_outputs(2449) <= a;
    layer1_outputs(2450) <= not (a xor b);
    layer1_outputs(2451) <= a xor b;
    layer1_outputs(2452) <= a and not b;
    layer1_outputs(2453) <= b;
    layer1_outputs(2454) <= a or b;
    layer1_outputs(2455) <= a xor b;
    layer1_outputs(2456) <= a xor b;
    layer1_outputs(2457) <= a and b;
    layer1_outputs(2458) <= b;
    layer1_outputs(2459) <= b and not a;
    layer1_outputs(2460) <= not a or b;
    layer1_outputs(2461) <= b;
    layer1_outputs(2462) <= a and not b;
    layer1_outputs(2463) <= not (a or b);
    layer1_outputs(2464) <= a xor b;
    layer1_outputs(2465) <= not a;
    layer1_outputs(2466) <= not a or b;
    layer1_outputs(2467) <= not a;
    layer1_outputs(2468) <= b;
    layer1_outputs(2469) <= not (a and b);
    layer1_outputs(2470) <= not a;
    layer1_outputs(2471) <= a;
    layer1_outputs(2472) <= a xor b;
    layer1_outputs(2473) <= a xor b;
    layer1_outputs(2474) <= b and not a;
    layer1_outputs(2475) <= not a;
    layer1_outputs(2476) <= a or b;
    layer1_outputs(2477) <= not b or a;
    layer1_outputs(2478) <= a and not b;
    layer1_outputs(2479) <= a;
    layer1_outputs(2480) <= not (a xor b);
    layer1_outputs(2481) <= b and not a;
    layer1_outputs(2482) <= a or b;
    layer1_outputs(2483) <= not (a xor b);
    layer1_outputs(2484) <= b;
    layer1_outputs(2485) <= not (a xor b);
    layer1_outputs(2486) <= a xor b;
    layer1_outputs(2487) <= not (a xor b);
    layer1_outputs(2488) <= b;
    layer1_outputs(2489) <= 1'b0;
    layer1_outputs(2490) <= a and b;
    layer1_outputs(2491) <= not a;
    layer1_outputs(2492) <= not (a xor b);
    layer1_outputs(2493) <= a;
    layer1_outputs(2494) <= b;
    layer1_outputs(2495) <= b and not a;
    layer1_outputs(2496) <= a and b;
    layer1_outputs(2497) <= b;
    layer1_outputs(2498) <= not (a and b);
    layer1_outputs(2499) <= a and b;
    layer1_outputs(2500) <= not a or b;
    layer1_outputs(2501) <= not b;
    layer1_outputs(2502) <= b;
    layer1_outputs(2503) <= not b;
    layer1_outputs(2504) <= b and not a;
    layer1_outputs(2505) <= not a or b;
    layer1_outputs(2506) <= not (a and b);
    layer1_outputs(2507) <= a and not b;
    layer1_outputs(2508) <= not a;
    layer1_outputs(2509) <= 1'b1;
    layer1_outputs(2510) <= a;
    layer1_outputs(2511) <= 1'b1;
    layer1_outputs(2512) <= not (a or b);
    layer1_outputs(2513) <= a or b;
    layer1_outputs(2514) <= a and not b;
    layer1_outputs(2515) <= not b or a;
    layer1_outputs(2516) <= not a or b;
    layer1_outputs(2517) <= not a or b;
    layer1_outputs(2518) <= not a;
    layer1_outputs(2519) <= not b;
    layer1_outputs(2520) <= a and b;
    layer1_outputs(2521) <= not (a or b);
    layer1_outputs(2522) <= not (a or b);
    layer1_outputs(2523) <= b;
    layer1_outputs(2524) <= a xor b;
    layer1_outputs(2525) <= b;
    layer1_outputs(2526) <= not a;
    layer1_outputs(2527) <= a;
    layer1_outputs(2528) <= a and not b;
    layer1_outputs(2529) <= b;
    layer1_outputs(2530) <= a and b;
    layer1_outputs(2531) <= not (a or b);
    layer1_outputs(2532) <= a and not b;
    layer1_outputs(2533) <= b;
    layer1_outputs(2534) <= not a;
    layer1_outputs(2535) <= a and not b;
    layer1_outputs(2536) <= b and not a;
    layer1_outputs(2537) <= 1'b1;
    layer1_outputs(2538) <= a xor b;
    layer1_outputs(2539) <= not b or a;
    layer1_outputs(2540) <= b;
    layer1_outputs(2541) <= not b or a;
    layer1_outputs(2542) <= a and b;
    layer1_outputs(2543) <= not b or a;
    layer1_outputs(2544) <= a xor b;
    layer1_outputs(2545) <= b;
    layer1_outputs(2546) <= not b or a;
    layer1_outputs(2547) <= not b;
    layer1_outputs(2548) <= not b;
    layer1_outputs(2549) <= b;
    layer1_outputs(2550) <= a and b;
    layer1_outputs(2551) <= not b;
    layer1_outputs(2552) <= not a or b;
    layer1_outputs(2553) <= not (a xor b);
    layer1_outputs(2554) <= not (a or b);
    layer1_outputs(2555) <= not (a xor b);
    layer1_outputs(2556) <= a and not b;
    layer1_outputs(2557) <= a and not b;
    layer1_outputs(2558) <= a and not b;
    layer1_outputs(2559) <= not b or a;
    layer1_outputs(2560) <= not b;
    layer1_outputs(2561) <= not b;
    layer1_outputs(2562) <= a and b;
    layer1_outputs(2563) <= not a;
    layer1_outputs(2564) <= not (a xor b);
    layer1_outputs(2565) <= not (a and b);
    layer1_outputs(2566) <= not a;
    layer1_outputs(2567) <= not (a xor b);
    layer1_outputs(2568) <= not (a or b);
    layer1_outputs(2569) <= a or b;
    layer1_outputs(2570) <= 1'b0;
    layer1_outputs(2571) <= a;
    layer1_outputs(2572) <= a;
    layer1_outputs(2573) <= not (a xor b);
    layer1_outputs(2574) <= not (a xor b);
    layer1_outputs(2575) <= a and not b;
    layer1_outputs(2576) <= a;
    layer1_outputs(2577) <= not a or b;
    layer1_outputs(2578) <= not (a xor b);
    layer1_outputs(2579) <= a xor b;
    layer1_outputs(2580) <= not a;
    layer1_outputs(2581) <= a and not b;
    layer1_outputs(2582) <= a xor b;
    layer1_outputs(2583) <= not b or a;
    layer1_outputs(2584) <= not a or b;
    layer1_outputs(2585) <= not a;
    layer1_outputs(2586) <= not (a or b);
    layer1_outputs(2587) <= not (a xor b);
    layer1_outputs(2588) <= not (a and b);
    layer1_outputs(2589) <= b and not a;
    layer1_outputs(2590) <= not (a or b);
    layer1_outputs(2591) <= a and not b;
    layer1_outputs(2592) <= not b or a;
    layer1_outputs(2593) <= not (a or b);
    layer1_outputs(2594) <= b;
    layer1_outputs(2595) <= not (a and b);
    layer1_outputs(2596) <= not b or a;
    layer1_outputs(2597) <= not b;
    layer1_outputs(2598) <= a xor b;
    layer1_outputs(2599) <= a and b;
    layer1_outputs(2600) <= not (a or b);
    layer1_outputs(2601) <= a or b;
    layer1_outputs(2602) <= not (a xor b);
    layer1_outputs(2603) <= not b;
    layer1_outputs(2604) <= a and b;
    layer1_outputs(2605) <= a;
    layer1_outputs(2606) <= not a or b;
    layer1_outputs(2607) <= a xor b;
    layer1_outputs(2608) <= b;
    layer1_outputs(2609) <= a or b;
    layer1_outputs(2610) <= not (a or b);
    layer1_outputs(2611) <= not b;
    layer1_outputs(2612) <= not a or b;
    layer1_outputs(2613) <= b and not a;
    layer1_outputs(2614) <= not a or b;
    layer1_outputs(2615) <= a and b;
    layer1_outputs(2616) <= b and not a;
    layer1_outputs(2617) <= b;
    layer1_outputs(2618) <= not (a or b);
    layer1_outputs(2619) <= a;
    layer1_outputs(2620) <= not a or b;
    layer1_outputs(2621) <= a and b;
    layer1_outputs(2622) <= b;
    layer1_outputs(2623) <= a and not b;
    layer1_outputs(2624) <= not (a and b);
    layer1_outputs(2625) <= a xor b;
    layer1_outputs(2626) <= not (a xor b);
    layer1_outputs(2627) <= not (a and b);
    layer1_outputs(2628) <= a xor b;
    layer1_outputs(2629) <= not a or b;
    layer1_outputs(2630) <= a;
    layer1_outputs(2631) <= a or b;
    layer1_outputs(2632) <= a xor b;
    layer1_outputs(2633) <= a and b;
    layer1_outputs(2634) <= not (a xor b);
    layer1_outputs(2635) <= b and not a;
    layer1_outputs(2636) <= a and not b;
    layer1_outputs(2637) <= not b;
    layer1_outputs(2638) <= a xor b;
    layer1_outputs(2639) <= a and not b;
    layer1_outputs(2640) <= b;
    layer1_outputs(2641) <= a;
    layer1_outputs(2642) <= a or b;
    layer1_outputs(2643) <= not (a and b);
    layer1_outputs(2644) <= not (a and b);
    layer1_outputs(2645) <= not a or b;
    layer1_outputs(2646) <= not b;
    layer1_outputs(2647) <= not a or b;
    layer1_outputs(2648) <= b;
    layer1_outputs(2649) <= a or b;
    layer1_outputs(2650) <= not b;
    layer1_outputs(2651) <= a and b;
    layer1_outputs(2652) <= a;
    layer1_outputs(2653) <= not (a and b);
    layer1_outputs(2654) <= not (a or b);
    layer1_outputs(2655) <= a;
    layer1_outputs(2656) <= 1'b0;
    layer1_outputs(2657) <= not (a xor b);
    layer1_outputs(2658) <= 1'b1;
    layer1_outputs(2659) <= not (a xor b);
    layer1_outputs(2660) <= a or b;
    layer1_outputs(2661) <= b;
    layer1_outputs(2662) <= b;
    layer1_outputs(2663) <= a and not b;
    layer1_outputs(2664) <= not b or a;
    layer1_outputs(2665) <= a;
    layer1_outputs(2666) <= 1'b0;
    layer1_outputs(2667) <= a and b;
    layer1_outputs(2668) <= a and b;
    layer1_outputs(2669) <= not a;
    layer1_outputs(2670) <= a or b;
    layer1_outputs(2671) <= b and not a;
    layer1_outputs(2672) <= b;
    layer1_outputs(2673) <= a;
    layer1_outputs(2674) <= b and not a;
    layer1_outputs(2675) <= a and not b;
    layer1_outputs(2676) <= not a;
    layer1_outputs(2677) <= not (a xor b);
    layer1_outputs(2678) <= not b;
    layer1_outputs(2679) <= a;
    layer1_outputs(2680) <= not a;
    layer1_outputs(2681) <= not (a or b);
    layer1_outputs(2682) <= a and not b;
    layer1_outputs(2683) <= not (a or b);
    layer1_outputs(2684) <= not b;
    layer1_outputs(2685) <= not (a xor b);
    layer1_outputs(2686) <= not b or a;
    layer1_outputs(2687) <= not b or a;
    layer1_outputs(2688) <= not (a xor b);
    layer1_outputs(2689) <= a xor b;
    layer1_outputs(2690) <= b and not a;
    layer1_outputs(2691) <= a or b;
    layer1_outputs(2692) <= not a;
    layer1_outputs(2693) <= 1'b1;
    layer1_outputs(2694) <= not b or a;
    layer1_outputs(2695) <= not a;
    layer1_outputs(2696) <= a or b;
    layer1_outputs(2697) <= not a or b;
    layer1_outputs(2698) <= not (a or b);
    layer1_outputs(2699) <= not a;
    layer1_outputs(2700) <= not b;
    layer1_outputs(2701) <= a and not b;
    layer1_outputs(2702) <= not (a xor b);
    layer1_outputs(2703) <= not (a or b);
    layer1_outputs(2704) <= not a;
    layer1_outputs(2705) <= not b;
    layer1_outputs(2706) <= not b or a;
    layer1_outputs(2707) <= a or b;
    layer1_outputs(2708) <= b;
    layer1_outputs(2709) <= a;
    layer1_outputs(2710) <= not b;
    layer1_outputs(2711) <= not (a or b);
    layer1_outputs(2712) <= not b or a;
    layer1_outputs(2713) <= not b;
    layer1_outputs(2714) <= not (a or b);
    layer1_outputs(2715) <= a and b;
    layer1_outputs(2716) <= a and not b;
    layer1_outputs(2717) <= not (a xor b);
    layer1_outputs(2718) <= not (a and b);
    layer1_outputs(2719) <= not (a and b);
    layer1_outputs(2720) <= b and not a;
    layer1_outputs(2721) <= not (a and b);
    layer1_outputs(2722) <= not (a xor b);
    layer1_outputs(2723) <= not (a or b);
    layer1_outputs(2724) <= a and b;
    layer1_outputs(2725) <= not b;
    layer1_outputs(2726) <= 1'b0;
    layer1_outputs(2727) <= not b;
    layer1_outputs(2728) <= not a or b;
    layer1_outputs(2729) <= not a;
    layer1_outputs(2730) <= a;
    layer1_outputs(2731) <= a or b;
    layer1_outputs(2732) <= a and not b;
    layer1_outputs(2733) <= a;
    layer1_outputs(2734) <= not a;
    layer1_outputs(2735) <= a or b;
    layer1_outputs(2736) <= a;
    layer1_outputs(2737) <= a or b;
    layer1_outputs(2738) <= 1'b0;
    layer1_outputs(2739) <= b;
    layer1_outputs(2740) <= a xor b;
    layer1_outputs(2741) <= not a;
    layer1_outputs(2742) <= not (a and b);
    layer1_outputs(2743) <= b and not a;
    layer1_outputs(2744) <= b;
    layer1_outputs(2745) <= a;
    layer1_outputs(2746) <= not b;
    layer1_outputs(2747) <= not a;
    layer1_outputs(2748) <= not a;
    layer1_outputs(2749) <= not a or b;
    layer1_outputs(2750) <= a;
    layer1_outputs(2751) <= not b;
    layer1_outputs(2752) <= not b;
    layer1_outputs(2753) <= not b;
    layer1_outputs(2754) <= a xor b;
    layer1_outputs(2755) <= a;
    layer1_outputs(2756) <= not (a or b);
    layer1_outputs(2757) <= a xor b;
    layer1_outputs(2758) <= b;
    layer1_outputs(2759) <= a and not b;
    layer1_outputs(2760) <= a xor b;
    layer1_outputs(2761) <= a and b;
    layer1_outputs(2762) <= not (a xor b);
    layer1_outputs(2763) <= a and b;
    layer1_outputs(2764) <= not a;
    layer1_outputs(2765) <= not (a xor b);
    layer1_outputs(2766) <= a and not b;
    layer1_outputs(2767) <= not (a or b);
    layer1_outputs(2768) <= b;
    layer1_outputs(2769) <= not b;
    layer1_outputs(2770) <= not (a or b);
    layer1_outputs(2771) <= not b or a;
    layer1_outputs(2772) <= a and b;
    layer1_outputs(2773) <= a xor b;
    layer1_outputs(2774) <= b;
    layer1_outputs(2775) <= b and not a;
    layer1_outputs(2776) <= a or b;
    layer1_outputs(2777) <= not b;
    layer1_outputs(2778) <= not a;
    layer1_outputs(2779) <= a and b;
    layer1_outputs(2780) <= a or b;
    layer1_outputs(2781) <= not (a xor b);
    layer1_outputs(2782) <= not (a or b);
    layer1_outputs(2783) <= not b;
    layer1_outputs(2784) <= not a;
    layer1_outputs(2785) <= not a;
    layer1_outputs(2786) <= a;
    layer1_outputs(2787) <= not a;
    layer1_outputs(2788) <= not a;
    layer1_outputs(2789) <= a or b;
    layer1_outputs(2790) <= a;
    layer1_outputs(2791) <= b;
    layer1_outputs(2792) <= b;
    layer1_outputs(2793) <= b;
    layer1_outputs(2794) <= a or b;
    layer1_outputs(2795) <= not a or b;
    layer1_outputs(2796) <= not b;
    layer1_outputs(2797) <= a and b;
    layer1_outputs(2798) <= not (a or b);
    layer1_outputs(2799) <= not b;
    layer1_outputs(2800) <= a and b;
    layer1_outputs(2801) <= not (a xor b);
    layer1_outputs(2802) <= a xor b;
    layer1_outputs(2803) <= a xor b;
    layer1_outputs(2804) <= not b or a;
    layer1_outputs(2805) <= not b;
    layer1_outputs(2806) <= not (a xor b);
    layer1_outputs(2807) <= not a or b;
    layer1_outputs(2808) <= a xor b;
    layer1_outputs(2809) <= not (a or b);
    layer1_outputs(2810) <= not (a and b);
    layer1_outputs(2811) <= a and b;
    layer1_outputs(2812) <= b and not a;
    layer1_outputs(2813) <= not (a xor b);
    layer1_outputs(2814) <= not (a and b);
    layer1_outputs(2815) <= not (a or b);
    layer1_outputs(2816) <= b;
    layer1_outputs(2817) <= not b;
    layer1_outputs(2818) <= b and not a;
    layer1_outputs(2819) <= b;
    layer1_outputs(2820) <= a and b;
    layer1_outputs(2821) <= a xor b;
    layer1_outputs(2822) <= a xor b;
    layer1_outputs(2823) <= not (a and b);
    layer1_outputs(2824) <= not (a or b);
    layer1_outputs(2825) <= a and not b;
    layer1_outputs(2826) <= not b;
    layer1_outputs(2827) <= b;
    layer1_outputs(2828) <= not a or b;
    layer1_outputs(2829) <= a and b;
    layer1_outputs(2830) <= b;
    layer1_outputs(2831) <= not b or a;
    layer1_outputs(2832) <= a and b;
    layer1_outputs(2833) <= b;
    layer1_outputs(2834) <= a and not b;
    layer1_outputs(2835) <= a and not b;
    layer1_outputs(2836) <= a;
    layer1_outputs(2837) <= a xor b;
    layer1_outputs(2838) <= a or b;
    layer1_outputs(2839) <= a or b;
    layer1_outputs(2840) <= a and b;
    layer1_outputs(2841) <= not (a xor b);
    layer1_outputs(2842) <= a and b;
    layer1_outputs(2843) <= b;
    layer1_outputs(2844) <= not a;
    layer1_outputs(2845) <= not (a or b);
    layer1_outputs(2846) <= not a;
    layer1_outputs(2847) <= b and not a;
    layer1_outputs(2848) <= b and not a;
    layer1_outputs(2849) <= not (a and b);
    layer1_outputs(2850) <= b and not a;
    layer1_outputs(2851) <= b;
    layer1_outputs(2852) <= a;
    layer1_outputs(2853) <= a and b;
    layer1_outputs(2854) <= not (a or b);
    layer1_outputs(2855) <= not (a and b);
    layer1_outputs(2856) <= not (a or b);
    layer1_outputs(2857) <= b and not a;
    layer1_outputs(2858) <= not b or a;
    layer1_outputs(2859) <= a xor b;
    layer1_outputs(2860) <= 1'b1;
    layer1_outputs(2861) <= a or b;
    layer1_outputs(2862) <= a or b;
    layer1_outputs(2863) <= not (a xor b);
    layer1_outputs(2864) <= a or b;
    layer1_outputs(2865) <= not b;
    layer1_outputs(2866) <= b;
    layer1_outputs(2867) <= 1'b0;
    layer1_outputs(2868) <= a and b;
    layer1_outputs(2869) <= not (a and b);
    layer1_outputs(2870) <= a xor b;
    layer1_outputs(2871) <= a xor b;
    layer1_outputs(2872) <= not (a or b);
    layer1_outputs(2873) <= a;
    layer1_outputs(2874) <= b and not a;
    layer1_outputs(2875) <= not a;
    layer1_outputs(2876) <= not b or a;
    layer1_outputs(2877) <= not (a or b);
    layer1_outputs(2878) <= not (a and b);
    layer1_outputs(2879) <= not a or b;
    layer1_outputs(2880) <= not (a xor b);
    layer1_outputs(2881) <= not a or b;
    layer1_outputs(2882) <= not a;
    layer1_outputs(2883) <= a and not b;
    layer1_outputs(2884) <= not (a or b);
    layer1_outputs(2885) <= a;
    layer1_outputs(2886) <= not (a or b);
    layer1_outputs(2887) <= not a;
    layer1_outputs(2888) <= not (a or b);
    layer1_outputs(2889) <= not b or a;
    layer1_outputs(2890) <= a and not b;
    layer1_outputs(2891) <= not (a or b);
    layer1_outputs(2892) <= a or b;
    layer1_outputs(2893) <= a;
    layer1_outputs(2894) <= a xor b;
    layer1_outputs(2895) <= not a;
    layer1_outputs(2896) <= a or b;
    layer1_outputs(2897) <= a and not b;
    layer1_outputs(2898) <= a and not b;
    layer1_outputs(2899) <= a or b;
    layer1_outputs(2900) <= 1'b0;
    layer1_outputs(2901) <= not (a and b);
    layer1_outputs(2902) <= a or b;
    layer1_outputs(2903) <= a xor b;
    layer1_outputs(2904) <= not a;
    layer1_outputs(2905) <= not a;
    layer1_outputs(2906) <= a xor b;
    layer1_outputs(2907) <= a or b;
    layer1_outputs(2908) <= a and b;
    layer1_outputs(2909) <= a;
    layer1_outputs(2910) <= not a;
    layer1_outputs(2911) <= a and not b;
    layer1_outputs(2912) <= not a;
    layer1_outputs(2913) <= not (a or b);
    layer1_outputs(2914) <= not a or b;
    layer1_outputs(2915) <= b;
    layer1_outputs(2916) <= not (a xor b);
    layer1_outputs(2917) <= not b;
    layer1_outputs(2918) <= a or b;
    layer1_outputs(2919) <= not a or b;
    layer1_outputs(2920) <= not a;
    layer1_outputs(2921) <= a;
    layer1_outputs(2922) <= a;
    layer1_outputs(2923) <= not b or a;
    layer1_outputs(2924) <= not a;
    layer1_outputs(2925) <= not a or b;
    layer1_outputs(2926) <= a;
    layer1_outputs(2927) <= a or b;
    layer1_outputs(2928) <= b and not a;
    layer1_outputs(2929) <= a xor b;
    layer1_outputs(2930) <= not (a and b);
    layer1_outputs(2931) <= not b;
    layer1_outputs(2932) <= a;
    layer1_outputs(2933) <= a and b;
    layer1_outputs(2934) <= not b or a;
    layer1_outputs(2935) <= not b or a;
    layer1_outputs(2936) <= not a or b;
    layer1_outputs(2937) <= 1'b0;
    layer1_outputs(2938) <= not b;
    layer1_outputs(2939) <= not b;
    layer1_outputs(2940) <= a or b;
    layer1_outputs(2941) <= b;
    layer1_outputs(2942) <= not b;
    layer1_outputs(2943) <= not a or b;
    layer1_outputs(2944) <= a or b;
    layer1_outputs(2945) <= 1'b1;
    layer1_outputs(2946) <= not b;
    layer1_outputs(2947) <= not (a and b);
    layer1_outputs(2948) <= 1'b0;
    layer1_outputs(2949) <= not (a and b);
    layer1_outputs(2950) <= a xor b;
    layer1_outputs(2951) <= 1'b1;
    layer1_outputs(2952) <= not b;
    layer1_outputs(2953) <= not (a xor b);
    layer1_outputs(2954) <= a and b;
    layer1_outputs(2955) <= not a or b;
    layer1_outputs(2956) <= a xor b;
    layer1_outputs(2957) <= b and not a;
    layer1_outputs(2958) <= a;
    layer1_outputs(2959) <= not (a or b);
    layer1_outputs(2960) <= b;
    layer1_outputs(2961) <= b;
    layer1_outputs(2962) <= a;
    layer1_outputs(2963) <= not a;
    layer1_outputs(2964) <= not b or a;
    layer1_outputs(2965) <= a xor b;
    layer1_outputs(2966) <= b and not a;
    layer1_outputs(2967) <= not b or a;
    layer1_outputs(2968) <= not (a and b);
    layer1_outputs(2969) <= a and not b;
    layer1_outputs(2970) <= not b;
    layer1_outputs(2971) <= b and not a;
    layer1_outputs(2972) <= a;
    layer1_outputs(2973) <= a and not b;
    layer1_outputs(2974) <= not (a or b);
    layer1_outputs(2975) <= not (a and b);
    layer1_outputs(2976) <= a xor b;
    layer1_outputs(2977) <= b;
    layer1_outputs(2978) <= not (a or b);
    layer1_outputs(2979) <= not (a or b);
    layer1_outputs(2980) <= not (a and b);
    layer1_outputs(2981) <= not b;
    layer1_outputs(2982) <= a;
    layer1_outputs(2983) <= not (a or b);
    layer1_outputs(2984) <= a xor b;
    layer1_outputs(2985) <= not (a or b);
    layer1_outputs(2986) <= a and b;
    layer1_outputs(2987) <= a;
    layer1_outputs(2988) <= not a or b;
    layer1_outputs(2989) <= not a or b;
    layer1_outputs(2990) <= not b;
    layer1_outputs(2991) <= a and not b;
    layer1_outputs(2992) <= not a or b;
    layer1_outputs(2993) <= a and not b;
    layer1_outputs(2994) <= a and b;
    layer1_outputs(2995) <= not (a or b);
    layer1_outputs(2996) <= 1'b0;
    layer1_outputs(2997) <= a or b;
    layer1_outputs(2998) <= b;
    layer1_outputs(2999) <= a or b;
    layer1_outputs(3000) <= not a or b;
    layer1_outputs(3001) <= a and b;
    layer1_outputs(3002) <= a xor b;
    layer1_outputs(3003) <= not (a or b);
    layer1_outputs(3004) <= not b;
    layer1_outputs(3005) <= a;
    layer1_outputs(3006) <= not a or b;
    layer1_outputs(3007) <= not a or b;
    layer1_outputs(3008) <= not a;
    layer1_outputs(3009) <= not b;
    layer1_outputs(3010) <= a and not b;
    layer1_outputs(3011) <= not a;
    layer1_outputs(3012) <= not b or a;
    layer1_outputs(3013) <= b;
    layer1_outputs(3014) <= not b;
    layer1_outputs(3015) <= not a;
    layer1_outputs(3016) <= not a or b;
    layer1_outputs(3017) <= not b or a;
    layer1_outputs(3018) <= not b;
    layer1_outputs(3019) <= not (a and b);
    layer1_outputs(3020) <= a;
    layer1_outputs(3021) <= b and not a;
    layer1_outputs(3022) <= not a or b;
    layer1_outputs(3023) <= a or b;
    layer1_outputs(3024) <= b;
    layer1_outputs(3025) <= not (a or b);
    layer1_outputs(3026) <= not (a xor b);
    layer1_outputs(3027) <= not b;
    layer1_outputs(3028) <= a or b;
    layer1_outputs(3029) <= a and b;
    layer1_outputs(3030) <= a and not b;
    layer1_outputs(3031) <= b;
    layer1_outputs(3032) <= a;
    layer1_outputs(3033) <= not (a xor b);
    layer1_outputs(3034) <= a;
    layer1_outputs(3035) <= b;
    layer1_outputs(3036) <= not (a xor b);
    layer1_outputs(3037) <= not a;
    layer1_outputs(3038) <= not b;
    layer1_outputs(3039) <= not (a and b);
    layer1_outputs(3040) <= not a;
    layer1_outputs(3041) <= not (a or b);
    layer1_outputs(3042) <= not (a and b);
    layer1_outputs(3043) <= 1'b1;
    layer1_outputs(3044) <= a xor b;
    layer1_outputs(3045) <= not a;
    layer1_outputs(3046) <= a or b;
    layer1_outputs(3047) <= not (a or b);
    layer1_outputs(3048) <= a and b;
    layer1_outputs(3049) <= a;
    layer1_outputs(3050) <= a or b;
    layer1_outputs(3051) <= not (a and b);
    layer1_outputs(3052) <= b and not a;
    layer1_outputs(3053) <= a and not b;
    layer1_outputs(3054) <= not (a xor b);
    layer1_outputs(3055) <= a;
    layer1_outputs(3056) <= not (a or b);
    layer1_outputs(3057) <= not b or a;
    layer1_outputs(3058) <= not b;
    layer1_outputs(3059) <= not b or a;
    layer1_outputs(3060) <= a xor b;
    layer1_outputs(3061) <= a and b;
    layer1_outputs(3062) <= a or b;
    layer1_outputs(3063) <= not (a or b);
    layer1_outputs(3064) <= b and not a;
    layer1_outputs(3065) <= a or b;
    layer1_outputs(3066) <= not b or a;
    layer1_outputs(3067) <= not b or a;
    layer1_outputs(3068) <= a;
    layer1_outputs(3069) <= a and b;
    layer1_outputs(3070) <= b;
    layer1_outputs(3071) <= not b or a;
    layer1_outputs(3072) <= not b;
    layer1_outputs(3073) <= not a or b;
    layer1_outputs(3074) <= b;
    layer1_outputs(3075) <= b;
    layer1_outputs(3076) <= a or b;
    layer1_outputs(3077) <= a or b;
    layer1_outputs(3078) <= a;
    layer1_outputs(3079) <= a and not b;
    layer1_outputs(3080) <= not (a and b);
    layer1_outputs(3081) <= not a;
    layer1_outputs(3082) <= not b;
    layer1_outputs(3083) <= not b;
    layer1_outputs(3084) <= not a or b;
    layer1_outputs(3085) <= a xor b;
    layer1_outputs(3086) <= not b or a;
    layer1_outputs(3087) <= a xor b;
    layer1_outputs(3088) <= b;
    layer1_outputs(3089) <= a;
    layer1_outputs(3090) <= not (a xor b);
    layer1_outputs(3091) <= a or b;
    layer1_outputs(3092) <= not (a or b);
    layer1_outputs(3093) <= not (a and b);
    layer1_outputs(3094) <= 1'b1;
    layer1_outputs(3095) <= not (a or b);
    layer1_outputs(3096) <= a;
    layer1_outputs(3097) <= b and not a;
    layer1_outputs(3098) <= a or b;
    layer1_outputs(3099) <= 1'b0;
    layer1_outputs(3100) <= a xor b;
    layer1_outputs(3101) <= not a or b;
    layer1_outputs(3102) <= a xor b;
    layer1_outputs(3103) <= not b;
    layer1_outputs(3104) <= b;
    layer1_outputs(3105) <= b and not a;
    layer1_outputs(3106) <= b;
    layer1_outputs(3107) <= a xor b;
    layer1_outputs(3108) <= b;
    layer1_outputs(3109) <= a xor b;
    layer1_outputs(3110) <= not a or b;
    layer1_outputs(3111) <= not b;
    layer1_outputs(3112) <= b and not a;
    layer1_outputs(3113) <= not a;
    layer1_outputs(3114) <= not a;
    layer1_outputs(3115) <= a;
    layer1_outputs(3116) <= not b or a;
    layer1_outputs(3117) <= 1'b1;
    layer1_outputs(3118) <= not (a or b);
    layer1_outputs(3119) <= a xor b;
    layer1_outputs(3120) <= not (a xor b);
    layer1_outputs(3121) <= not (a or b);
    layer1_outputs(3122) <= not (a or b);
    layer1_outputs(3123) <= not (a and b);
    layer1_outputs(3124) <= a and not b;
    layer1_outputs(3125) <= a xor b;
    layer1_outputs(3126) <= not a or b;
    layer1_outputs(3127) <= not b;
    layer1_outputs(3128) <= not (a xor b);
    layer1_outputs(3129) <= a and b;
    layer1_outputs(3130) <= b;
    layer1_outputs(3131) <= not a;
    layer1_outputs(3132) <= b and not a;
    layer1_outputs(3133) <= b;
    layer1_outputs(3134) <= not b;
    layer1_outputs(3135) <= b and not a;
    layer1_outputs(3136) <= a and b;
    layer1_outputs(3137) <= a and not b;
    layer1_outputs(3138) <= not (a xor b);
    layer1_outputs(3139) <= not (a xor b);
    layer1_outputs(3140) <= a;
    layer1_outputs(3141) <= b;
    layer1_outputs(3142) <= a and not b;
    layer1_outputs(3143) <= not a or b;
    layer1_outputs(3144) <= not b or a;
    layer1_outputs(3145) <= not b;
    layer1_outputs(3146) <= not b;
    layer1_outputs(3147) <= a;
    layer1_outputs(3148) <= not (a and b);
    layer1_outputs(3149) <= not a or b;
    layer1_outputs(3150) <= b;
    layer1_outputs(3151) <= not a;
    layer1_outputs(3152) <= not a or b;
    layer1_outputs(3153) <= not (a xor b);
    layer1_outputs(3154) <= a xor b;
    layer1_outputs(3155) <= a and b;
    layer1_outputs(3156) <= b and not a;
    layer1_outputs(3157) <= not a or b;
    layer1_outputs(3158) <= 1'b0;
    layer1_outputs(3159) <= not (a and b);
    layer1_outputs(3160) <= a and not b;
    layer1_outputs(3161) <= a xor b;
    layer1_outputs(3162) <= b;
    layer1_outputs(3163) <= b;
    layer1_outputs(3164) <= not a;
    layer1_outputs(3165) <= not b;
    layer1_outputs(3166) <= b and not a;
    layer1_outputs(3167) <= not a or b;
    layer1_outputs(3168) <= not a or b;
    layer1_outputs(3169) <= a or b;
    layer1_outputs(3170) <= a;
    layer1_outputs(3171) <= a or b;
    layer1_outputs(3172) <= not (a or b);
    layer1_outputs(3173) <= a and b;
    layer1_outputs(3174) <= not (a xor b);
    layer1_outputs(3175) <= not (a or b);
    layer1_outputs(3176) <= not a or b;
    layer1_outputs(3177) <= not b;
    layer1_outputs(3178) <= b and not a;
    layer1_outputs(3179) <= not (a xor b);
    layer1_outputs(3180) <= 1'b0;
    layer1_outputs(3181) <= a and not b;
    layer1_outputs(3182) <= a and b;
    layer1_outputs(3183) <= not b;
    layer1_outputs(3184) <= a and not b;
    layer1_outputs(3185) <= not (a and b);
    layer1_outputs(3186) <= a;
    layer1_outputs(3187) <= not (a and b);
    layer1_outputs(3188) <= a and not b;
    layer1_outputs(3189) <= not (a xor b);
    layer1_outputs(3190) <= not a or b;
    layer1_outputs(3191) <= not a or b;
    layer1_outputs(3192) <= not a;
    layer1_outputs(3193) <= not (a or b);
    layer1_outputs(3194) <= not a or b;
    layer1_outputs(3195) <= not (a xor b);
    layer1_outputs(3196) <= not b;
    layer1_outputs(3197) <= b and not a;
    layer1_outputs(3198) <= not a;
    layer1_outputs(3199) <= not b or a;
    layer1_outputs(3200) <= a;
    layer1_outputs(3201) <= a;
    layer1_outputs(3202) <= a or b;
    layer1_outputs(3203) <= not (a xor b);
    layer1_outputs(3204) <= a and not b;
    layer1_outputs(3205) <= not b;
    layer1_outputs(3206) <= b;
    layer1_outputs(3207) <= not a or b;
    layer1_outputs(3208) <= not b or a;
    layer1_outputs(3209) <= not (a and b);
    layer1_outputs(3210) <= not (a and b);
    layer1_outputs(3211) <= not (a or b);
    layer1_outputs(3212) <= a xor b;
    layer1_outputs(3213) <= not (a and b);
    layer1_outputs(3214) <= not (a or b);
    layer1_outputs(3215) <= b and not a;
    layer1_outputs(3216) <= a and not b;
    layer1_outputs(3217) <= not a;
    layer1_outputs(3218) <= not (a and b);
    layer1_outputs(3219) <= not (a and b);
    layer1_outputs(3220) <= a or b;
    layer1_outputs(3221) <= a;
    layer1_outputs(3222) <= not a or b;
    layer1_outputs(3223) <= not (a xor b);
    layer1_outputs(3224) <= b and not a;
    layer1_outputs(3225) <= not a or b;
    layer1_outputs(3226) <= b and not a;
    layer1_outputs(3227) <= not b or a;
    layer1_outputs(3228) <= b;
    layer1_outputs(3229) <= b and not a;
    layer1_outputs(3230) <= a and b;
    layer1_outputs(3231) <= a xor b;
    layer1_outputs(3232) <= b;
    layer1_outputs(3233) <= not a;
    layer1_outputs(3234) <= b and not a;
    layer1_outputs(3235) <= b;
    layer1_outputs(3236) <= a;
    layer1_outputs(3237) <= a;
    layer1_outputs(3238) <= b;
    layer1_outputs(3239) <= not (a and b);
    layer1_outputs(3240) <= a or b;
    layer1_outputs(3241) <= a xor b;
    layer1_outputs(3242) <= a xor b;
    layer1_outputs(3243) <= b and not a;
    layer1_outputs(3244) <= a;
    layer1_outputs(3245) <= a;
    layer1_outputs(3246) <= a xor b;
    layer1_outputs(3247) <= not b or a;
    layer1_outputs(3248) <= a and not b;
    layer1_outputs(3249) <= a;
    layer1_outputs(3250) <= b;
    layer1_outputs(3251) <= not a;
    layer1_outputs(3252) <= not a or b;
    layer1_outputs(3253) <= a;
    layer1_outputs(3254) <= not b;
    layer1_outputs(3255) <= not (a xor b);
    layer1_outputs(3256) <= not a;
    layer1_outputs(3257) <= not b;
    layer1_outputs(3258) <= a and not b;
    layer1_outputs(3259) <= not a;
    layer1_outputs(3260) <= not a;
    layer1_outputs(3261) <= a or b;
    layer1_outputs(3262) <= not b;
    layer1_outputs(3263) <= a or b;
    layer1_outputs(3264) <= not b;
    layer1_outputs(3265) <= a or b;
    layer1_outputs(3266) <= not b;
    layer1_outputs(3267) <= not (a and b);
    layer1_outputs(3268) <= not (a or b);
    layer1_outputs(3269) <= a and b;
    layer1_outputs(3270) <= not b or a;
    layer1_outputs(3271) <= a or b;
    layer1_outputs(3272) <= not (a or b);
    layer1_outputs(3273) <= not (a and b);
    layer1_outputs(3274) <= b and not a;
    layer1_outputs(3275) <= a;
    layer1_outputs(3276) <= not a;
    layer1_outputs(3277) <= a;
    layer1_outputs(3278) <= not (a and b);
    layer1_outputs(3279) <= b and not a;
    layer1_outputs(3280) <= not (a and b);
    layer1_outputs(3281) <= not a or b;
    layer1_outputs(3282) <= not (a xor b);
    layer1_outputs(3283) <= a or b;
    layer1_outputs(3284) <= not (a xor b);
    layer1_outputs(3285) <= 1'b0;
    layer1_outputs(3286) <= not b or a;
    layer1_outputs(3287) <= not b or a;
    layer1_outputs(3288) <= a and b;
    layer1_outputs(3289) <= a and not b;
    layer1_outputs(3290) <= a;
    layer1_outputs(3291) <= b and not a;
    layer1_outputs(3292) <= not a or b;
    layer1_outputs(3293) <= b and not a;
    layer1_outputs(3294) <= not a or b;
    layer1_outputs(3295) <= not a or b;
    layer1_outputs(3296) <= b;
    layer1_outputs(3297) <= b;
    layer1_outputs(3298) <= not b;
    layer1_outputs(3299) <= not b or a;
    layer1_outputs(3300) <= a xor b;
    layer1_outputs(3301) <= not b or a;
    layer1_outputs(3302) <= not (a and b);
    layer1_outputs(3303) <= not a;
    layer1_outputs(3304) <= a xor b;
    layer1_outputs(3305) <= not a or b;
    layer1_outputs(3306) <= not (a xor b);
    layer1_outputs(3307) <= not (a or b);
    layer1_outputs(3308) <= not (a or b);
    layer1_outputs(3309) <= not b or a;
    layer1_outputs(3310) <= not (a xor b);
    layer1_outputs(3311) <= a and b;
    layer1_outputs(3312) <= b and not a;
    layer1_outputs(3313) <= a and b;
    layer1_outputs(3314) <= not (a xor b);
    layer1_outputs(3315) <= b;
    layer1_outputs(3316) <= not a or b;
    layer1_outputs(3317) <= b and not a;
    layer1_outputs(3318) <= not b;
    layer1_outputs(3319) <= a and b;
    layer1_outputs(3320) <= not b;
    layer1_outputs(3321) <= not (a or b);
    layer1_outputs(3322) <= not b;
    layer1_outputs(3323) <= a xor b;
    layer1_outputs(3324) <= not a or b;
    layer1_outputs(3325) <= b and not a;
    layer1_outputs(3326) <= not (a xor b);
    layer1_outputs(3327) <= not (a xor b);
    layer1_outputs(3328) <= not a;
    layer1_outputs(3329) <= a xor b;
    layer1_outputs(3330) <= a or b;
    layer1_outputs(3331) <= not b or a;
    layer1_outputs(3332) <= b;
    layer1_outputs(3333) <= b and not a;
    layer1_outputs(3334) <= not b;
    layer1_outputs(3335) <= a xor b;
    layer1_outputs(3336) <= not b;
    layer1_outputs(3337) <= b;
    layer1_outputs(3338) <= a and not b;
    layer1_outputs(3339) <= a or b;
    layer1_outputs(3340) <= a;
    layer1_outputs(3341) <= a and not b;
    layer1_outputs(3342) <= b;
    layer1_outputs(3343) <= a xor b;
    layer1_outputs(3344) <= a xor b;
    layer1_outputs(3345) <= not (a xor b);
    layer1_outputs(3346) <= not (a or b);
    layer1_outputs(3347) <= not (a and b);
    layer1_outputs(3348) <= not (a xor b);
    layer1_outputs(3349) <= not a or b;
    layer1_outputs(3350) <= not (a or b);
    layer1_outputs(3351) <= not (a xor b);
    layer1_outputs(3352) <= a or b;
    layer1_outputs(3353) <= not (a and b);
    layer1_outputs(3354) <= a and not b;
    layer1_outputs(3355) <= not (a xor b);
    layer1_outputs(3356) <= a and b;
    layer1_outputs(3357) <= not (a xor b);
    layer1_outputs(3358) <= a;
    layer1_outputs(3359) <= not (a or b);
    layer1_outputs(3360) <= not b or a;
    layer1_outputs(3361) <= not (a xor b);
    layer1_outputs(3362) <= a;
    layer1_outputs(3363) <= not b or a;
    layer1_outputs(3364) <= not b;
    layer1_outputs(3365) <= a xor b;
    layer1_outputs(3366) <= 1'b1;
    layer1_outputs(3367) <= not a or b;
    layer1_outputs(3368) <= a or b;
    layer1_outputs(3369) <= a and b;
    layer1_outputs(3370) <= a and b;
    layer1_outputs(3371) <= not (a and b);
    layer1_outputs(3372) <= not a;
    layer1_outputs(3373) <= a and b;
    layer1_outputs(3374) <= a xor b;
    layer1_outputs(3375) <= not b or a;
    layer1_outputs(3376) <= a and not b;
    layer1_outputs(3377) <= b and not a;
    layer1_outputs(3378) <= not (a xor b);
    layer1_outputs(3379) <= a xor b;
    layer1_outputs(3380) <= a and not b;
    layer1_outputs(3381) <= a xor b;
    layer1_outputs(3382) <= a and not b;
    layer1_outputs(3383) <= a or b;
    layer1_outputs(3384) <= not a or b;
    layer1_outputs(3385) <= a and b;
    layer1_outputs(3386) <= not (a and b);
    layer1_outputs(3387) <= not (a and b);
    layer1_outputs(3388) <= b;
    layer1_outputs(3389) <= a xor b;
    layer1_outputs(3390) <= not b;
    layer1_outputs(3391) <= a xor b;
    layer1_outputs(3392) <= not b;
    layer1_outputs(3393) <= a and b;
    layer1_outputs(3394) <= a;
    layer1_outputs(3395) <= b and not a;
    layer1_outputs(3396) <= a and b;
    layer1_outputs(3397) <= not a;
    layer1_outputs(3398) <= a xor b;
    layer1_outputs(3399) <= b;
    layer1_outputs(3400) <= b;
    layer1_outputs(3401) <= not (a or b);
    layer1_outputs(3402) <= a;
    layer1_outputs(3403) <= a and b;
    layer1_outputs(3404) <= a;
    layer1_outputs(3405) <= b and not a;
    layer1_outputs(3406) <= not a;
    layer1_outputs(3407) <= a or b;
    layer1_outputs(3408) <= b;
    layer1_outputs(3409) <= a and b;
    layer1_outputs(3410) <= a or b;
    layer1_outputs(3411) <= a and b;
    layer1_outputs(3412) <= not (a or b);
    layer1_outputs(3413) <= not a or b;
    layer1_outputs(3414) <= not a or b;
    layer1_outputs(3415) <= a or b;
    layer1_outputs(3416) <= not b or a;
    layer1_outputs(3417) <= not (a xor b);
    layer1_outputs(3418) <= not b or a;
    layer1_outputs(3419) <= not (a xor b);
    layer1_outputs(3420) <= not (a xor b);
    layer1_outputs(3421) <= a xor b;
    layer1_outputs(3422) <= not a;
    layer1_outputs(3423) <= not a;
    layer1_outputs(3424) <= not a or b;
    layer1_outputs(3425) <= not b;
    layer1_outputs(3426) <= b;
    layer1_outputs(3427) <= a and not b;
    layer1_outputs(3428) <= a and b;
    layer1_outputs(3429) <= b and not a;
    layer1_outputs(3430) <= not (a or b);
    layer1_outputs(3431) <= b and not a;
    layer1_outputs(3432) <= a and b;
    layer1_outputs(3433) <= a and b;
    layer1_outputs(3434) <= not b or a;
    layer1_outputs(3435) <= not (a and b);
    layer1_outputs(3436) <= not b;
    layer1_outputs(3437) <= 1'b1;
    layer1_outputs(3438) <= not (a or b);
    layer1_outputs(3439) <= not b;
    layer1_outputs(3440) <= a and b;
    layer1_outputs(3441) <= not b;
    layer1_outputs(3442) <= not (a and b);
    layer1_outputs(3443) <= not a;
    layer1_outputs(3444) <= a and b;
    layer1_outputs(3445) <= b;
    layer1_outputs(3446) <= a and not b;
    layer1_outputs(3447) <= b;
    layer1_outputs(3448) <= a and b;
    layer1_outputs(3449) <= not (a or b);
    layer1_outputs(3450) <= b;
    layer1_outputs(3451) <= not (a xor b);
    layer1_outputs(3452) <= not (a xor b);
    layer1_outputs(3453) <= not b;
    layer1_outputs(3454) <= not (a and b);
    layer1_outputs(3455) <= not (a and b);
    layer1_outputs(3456) <= not a;
    layer1_outputs(3457) <= b;
    layer1_outputs(3458) <= a;
    layer1_outputs(3459) <= not b;
    layer1_outputs(3460) <= not (a xor b);
    layer1_outputs(3461) <= a and b;
    layer1_outputs(3462) <= a;
    layer1_outputs(3463) <= not b;
    layer1_outputs(3464) <= a and b;
    layer1_outputs(3465) <= a xor b;
    layer1_outputs(3466) <= a and not b;
    layer1_outputs(3467) <= not a or b;
    layer1_outputs(3468) <= not (a and b);
    layer1_outputs(3469) <= b and not a;
    layer1_outputs(3470) <= 1'b0;
    layer1_outputs(3471) <= not a;
    layer1_outputs(3472) <= a;
    layer1_outputs(3473) <= a;
    layer1_outputs(3474) <= a and not b;
    layer1_outputs(3475) <= b;
    layer1_outputs(3476) <= not b;
    layer1_outputs(3477) <= b;
    layer1_outputs(3478) <= b;
    layer1_outputs(3479) <= not (a and b);
    layer1_outputs(3480) <= not (a xor b);
    layer1_outputs(3481) <= b;
    layer1_outputs(3482) <= not b or a;
    layer1_outputs(3483) <= a xor b;
    layer1_outputs(3484) <= a;
    layer1_outputs(3485) <= not a;
    layer1_outputs(3486) <= b and not a;
    layer1_outputs(3487) <= a;
    layer1_outputs(3488) <= b and not a;
    layer1_outputs(3489) <= b;
    layer1_outputs(3490) <= a and not b;
    layer1_outputs(3491) <= a and not b;
    layer1_outputs(3492) <= a and b;
    layer1_outputs(3493) <= not a;
    layer1_outputs(3494) <= b;
    layer1_outputs(3495) <= a;
    layer1_outputs(3496) <= not b;
    layer1_outputs(3497) <= a and b;
    layer1_outputs(3498) <= a;
    layer1_outputs(3499) <= not a;
    layer1_outputs(3500) <= b and not a;
    layer1_outputs(3501) <= a or b;
    layer1_outputs(3502) <= b;
    layer1_outputs(3503) <= a;
    layer1_outputs(3504) <= not b;
    layer1_outputs(3505) <= not (a xor b);
    layer1_outputs(3506) <= not (a or b);
    layer1_outputs(3507) <= a xor b;
    layer1_outputs(3508) <= not (a or b);
    layer1_outputs(3509) <= not (a and b);
    layer1_outputs(3510) <= b and not a;
    layer1_outputs(3511) <= a or b;
    layer1_outputs(3512) <= a;
    layer1_outputs(3513) <= not a;
    layer1_outputs(3514) <= b and not a;
    layer1_outputs(3515) <= not a or b;
    layer1_outputs(3516) <= a or b;
    layer1_outputs(3517) <= a or b;
    layer1_outputs(3518) <= not (a or b);
    layer1_outputs(3519) <= 1'b1;
    layer1_outputs(3520) <= not b;
    layer1_outputs(3521) <= not a or b;
    layer1_outputs(3522) <= not a or b;
    layer1_outputs(3523) <= a and b;
    layer1_outputs(3524) <= a xor b;
    layer1_outputs(3525) <= not (a or b);
    layer1_outputs(3526) <= 1'b0;
    layer1_outputs(3527) <= not a;
    layer1_outputs(3528) <= not (a and b);
    layer1_outputs(3529) <= not (a and b);
    layer1_outputs(3530) <= not b;
    layer1_outputs(3531) <= a xor b;
    layer1_outputs(3532) <= not (a and b);
    layer1_outputs(3533) <= not a;
    layer1_outputs(3534) <= a;
    layer1_outputs(3535) <= a and b;
    layer1_outputs(3536) <= not (a xor b);
    layer1_outputs(3537) <= not b or a;
    layer1_outputs(3538) <= not a;
    layer1_outputs(3539) <= not a or b;
    layer1_outputs(3540) <= b and not a;
    layer1_outputs(3541) <= b;
    layer1_outputs(3542) <= not (a and b);
    layer1_outputs(3543) <= not (a xor b);
    layer1_outputs(3544) <= not (a and b);
    layer1_outputs(3545) <= b;
    layer1_outputs(3546) <= not (a and b);
    layer1_outputs(3547) <= not (a or b);
    layer1_outputs(3548) <= a and b;
    layer1_outputs(3549) <= a or b;
    layer1_outputs(3550) <= a;
    layer1_outputs(3551) <= b;
    layer1_outputs(3552) <= not (a or b);
    layer1_outputs(3553) <= b and not a;
    layer1_outputs(3554) <= a or b;
    layer1_outputs(3555) <= not (a or b);
    layer1_outputs(3556) <= b;
    layer1_outputs(3557) <= a;
    layer1_outputs(3558) <= 1'b0;
    layer1_outputs(3559) <= b;
    layer1_outputs(3560) <= a;
    layer1_outputs(3561) <= not b;
    layer1_outputs(3562) <= not b;
    layer1_outputs(3563) <= not b or a;
    layer1_outputs(3564) <= b and not a;
    layer1_outputs(3565) <= a or b;
    layer1_outputs(3566) <= not a;
    layer1_outputs(3567) <= not a or b;
    layer1_outputs(3568) <= a and b;
    layer1_outputs(3569) <= a and not b;
    layer1_outputs(3570) <= not b or a;
    layer1_outputs(3571) <= b and not a;
    layer1_outputs(3572) <= a and b;
    layer1_outputs(3573) <= not b;
    layer1_outputs(3574) <= b and not a;
    layer1_outputs(3575) <= not a or b;
    layer1_outputs(3576) <= not a;
    layer1_outputs(3577) <= not (a or b);
    layer1_outputs(3578) <= b;
    layer1_outputs(3579) <= a or b;
    layer1_outputs(3580) <= a or b;
    layer1_outputs(3581) <= b and not a;
    layer1_outputs(3582) <= not b;
    layer1_outputs(3583) <= 1'b0;
    layer1_outputs(3584) <= not (a or b);
    layer1_outputs(3585) <= not b or a;
    layer1_outputs(3586) <= not (a and b);
    layer1_outputs(3587) <= not b;
    layer1_outputs(3588) <= not (a xor b);
    layer1_outputs(3589) <= a or b;
    layer1_outputs(3590) <= not a;
    layer1_outputs(3591) <= b;
    layer1_outputs(3592) <= not (a and b);
    layer1_outputs(3593) <= a;
    layer1_outputs(3594) <= a;
    layer1_outputs(3595) <= not a or b;
    layer1_outputs(3596) <= not (a and b);
    layer1_outputs(3597) <= 1'b1;
    layer1_outputs(3598) <= a and b;
    layer1_outputs(3599) <= not (a xor b);
    layer1_outputs(3600) <= not a;
    layer1_outputs(3601) <= 1'b1;
    layer1_outputs(3602) <= not a or b;
    layer1_outputs(3603) <= a and b;
    layer1_outputs(3604) <= not a or b;
    layer1_outputs(3605) <= not (a and b);
    layer1_outputs(3606) <= a xor b;
    layer1_outputs(3607) <= a or b;
    layer1_outputs(3608) <= not (a and b);
    layer1_outputs(3609) <= a;
    layer1_outputs(3610) <= not a or b;
    layer1_outputs(3611) <= not (a and b);
    layer1_outputs(3612) <= b;
    layer1_outputs(3613) <= not b or a;
    layer1_outputs(3614) <= not a;
    layer1_outputs(3615) <= a;
    layer1_outputs(3616) <= a;
    layer1_outputs(3617) <= not a;
    layer1_outputs(3618) <= b;
    layer1_outputs(3619) <= not b;
    layer1_outputs(3620) <= a and b;
    layer1_outputs(3621) <= a;
    layer1_outputs(3622) <= not a or b;
    layer1_outputs(3623) <= not (a xor b);
    layer1_outputs(3624) <= not a or b;
    layer1_outputs(3625) <= b and not a;
    layer1_outputs(3626) <= a and not b;
    layer1_outputs(3627) <= not b or a;
    layer1_outputs(3628) <= a xor b;
    layer1_outputs(3629) <= not b or a;
    layer1_outputs(3630) <= not (a xor b);
    layer1_outputs(3631) <= not (a and b);
    layer1_outputs(3632) <= not a;
    layer1_outputs(3633) <= not a or b;
    layer1_outputs(3634) <= a;
    layer1_outputs(3635) <= not (a and b);
    layer1_outputs(3636) <= not (a xor b);
    layer1_outputs(3637) <= not a;
    layer1_outputs(3638) <= not b;
    layer1_outputs(3639) <= not (a xor b);
    layer1_outputs(3640) <= a and b;
    layer1_outputs(3641) <= not a;
    layer1_outputs(3642) <= not (a or b);
    layer1_outputs(3643) <= b and not a;
    layer1_outputs(3644) <= not a;
    layer1_outputs(3645) <= a and b;
    layer1_outputs(3646) <= a or b;
    layer1_outputs(3647) <= a and b;
    layer1_outputs(3648) <= not b;
    layer1_outputs(3649) <= a;
    layer1_outputs(3650) <= a xor b;
    layer1_outputs(3651) <= a;
    layer1_outputs(3652) <= not a;
    layer1_outputs(3653) <= 1'b1;
    layer1_outputs(3654) <= b;
    layer1_outputs(3655) <= not (a and b);
    layer1_outputs(3656) <= not a or b;
    layer1_outputs(3657) <= b;
    layer1_outputs(3658) <= not (a or b);
    layer1_outputs(3659) <= not (a and b);
    layer1_outputs(3660) <= not (a and b);
    layer1_outputs(3661) <= b;
    layer1_outputs(3662) <= a or b;
    layer1_outputs(3663) <= not (a and b);
    layer1_outputs(3664) <= not b or a;
    layer1_outputs(3665) <= a and b;
    layer1_outputs(3666) <= a xor b;
    layer1_outputs(3667) <= not b or a;
    layer1_outputs(3668) <= not (a or b);
    layer1_outputs(3669) <= not b;
    layer1_outputs(3670) <= a and b;
    layer1_outputs(3671) <= a;
    layer1_outputs(3672) <= not b or a;
    layer1_outputs(3673) <= not a or b;
    layer1_outputs(3674) <= b;
    layer1_outputs(3675) <= not b;
    layer1_outputs(3676) <= b;
    layer1_outputs(3677) <= a and b;
    layer1_outputs(3678) <= a and not b;
    layer1_outputs(3679) <= not (a or b);
    layer1_outputs(3680) <= a and not b;
    layer1_outputs(3681) <= b;
    layer1_outputs(3682) <= not (a xor b);
    layer1_outputs(3683) <= b and not a;
    layer1_outputs(3684) <= not a or b;
    layer1_outputs(3685) <= b and not a;
    layer1_outputs(3686) <= not b or a;
    layer1_outputs(3687) <= a and b;
    layer1_outputs(3688) <= a;
    layer1_outputs(3689) <= not (a and b);
    layer1_outputs(3690) <= 1'b1;
    layer1_outputs(3691) <= not a;
    layer1_outputs(3692) <= b;
    layer1_outputs(3693) <= a and not b;
    layer1_outputs(3694) <= not b;
    layer1_outputs(3695) <= not (a xor b);
    layer1_outputs(3696) <= a and b;
    layer1_outputs(3697) <= a and not b;
    layer1_outputs(3698) <= not b;
    layer1_outputs(3699) <= not a or b;
    layer1_outputs(3700) <= not a or b;
    layer1_outputs(3701) <= a;
    layer1_outputs(3702) <= b;
    layer1_outputs(3703) <= not (a or b);
    layer1_outputs(3704) <= b;
    layer1_outputs(3705) <= 1'b0;
    layer1_outputs(3706) <= not b;
    layer1_outputs(3707) <= not (a xor b);
    layer1_outputs(3708) <= not (a or b);
    layer1_outputs(3709) <= not a;
    layer1_outputs(3710) <= a;
    layer1_outputs(3711) <= a and not b;
    layer1_outputs(3712) <= not (a or b);
    layer1_outputs(3713) <= not a or b;
    layer1_outputs(3714) <= b;
    layer1_outputs(3715) <= a;
    layer1_outputs(3716) <= not b or a;
    layer1_outputs(3717) <= not (a or b);
    layer1_outputs(3718) <= not a;
    layer1_outputs(3719) <= a;
    layer1_outputs(3720) <= not a or b;
    layer1_outputs(3721) <= a xor b;
    layer1_outputs(3722) <= 1'b1;
    layer1_outputs(3723) <= not (a or b);
    layer1_outputs(3724) <= not (a and b);
    layer1_outputs(3725) <= not (a or b);
    layer1_outputs(3726) <= a or b;
    layer1_outputs(3727) <= not a;
    layer1_outputs(3728) <= not b;
    layer1_outputs(3729) <= not a;
    layer1_outputs(3730) <= b;
    layer1_outputs(3731) <= not a or b;
    layer1_outputs(3732) <= not a;
    layer1_outputs(3733) <= b and not a;
    layer1_outputs(3734) <= not (a xor b);
    layer1_outputs(3735) <= a or b;
    layer1_outputs(3736) <= not (a xor b);
    layer1_outputs(3737) <= a and b;
    layer1_outputs(3738) <= not a or b;
    layer1_outputs(3739) <= not b or a;
    layer1_outputs(3740) <= a;
    layer1_outputs(3741) <= not (a xor b);
    layer1_outputs(3742) <= b;
    layer1_outputs(3743) <= not b or a;
    layer1_outputs(3744) <= not b or a;
    layer1_outputs(3745) <= not (a or b);
    layer1_outputs(3746) <= 1'b0;
    layer1_outputs(3747) <= not a or b;
    layer1_outputs(3748) <= a and not b;
    layer1_outputs(3749) <= not b;
    layer1_outputs(3750) <= a and b;
    layer1_outputs(3751) <= 1'b1;
    layer1_outputs(3752) <= not (a xor b);
    layer1_outputs(3753) <= a;
    layer1_outputs(3754) <= b;
    layer1_outputs(3755) <= not b;
    layer1_outputs(3756) <= b and not a;
    layer1_outputs(3757) <= b;
    layer1_outputs(3758) <= b;
    layer1_outputs(3759) <= b;
    layer1_outputs(3760) <= not b;
    layer1_outputs(3761) <= a;
    layer1_outputs(3762) <= a and b;
    layer1_outputs(3763) <= a or b;
    layer1_outputs(3764) <= not (a or b);
    layer1_outputs(3765) <= b;
    layer1_outputs(3766) <= a and not b;
    layer1_outputs(3767) <= a;
    layer1_outputs(3768) <= not (a or b);
    layer1_outputs(3769) <= a;
    layer1_outputs(3770) <= not (a xor b);
    layer1_outputs(3771) <= a or b;
    layer1_outputs(3772) <= a;
    layer1_outputs(3773) <= 1'b0;
    layer1_outputs(3774) <= a and not b;
    layer1_outputs(3775) <= not b or a;
    layer1_outputs(3776) <= not a or b;
    layer1_outputs(3777) <= a;
    layer1_outputs(3778) <= not (a or b);
    layer1_outputs(3779) <= not b;
    layer1_outputs(3780) <= a;
    layer1_outputs(3781) <= not a;
    layer1_outputs(3782) <= not (a or b);
    layer1_outputs(3783) <= a xor b;
    layer1_outputs(3784) <= not (a and b);
    layer1_outputs(3785) <= not a;
    layer1_outputs(3786) <= a;
    layer1_outputs(3787) <= a;
    layer1_outputs(3788) <= 1'b1;
    layer1_outputs(3789) <= not b or a;
    layer1_outputs(3790) <= a xor b;
    layer1_outputs(3791) <= not b or a;
    layer1_outputs(3792) <= a and b;
    layer1_outputs(3793) <= b;
    layer1_outputs(3794) <= not a;
    layer1_outputs(3795) <= a;
    layer1_outputs(3796) <= a or b;
    layer1_outputs(3797) <= not b;
    layer1_outputs(3798) <= not a or b;
    layer1_outputs(3799) <= 1'b1;
    layer1_outputs(3800) <= not b;
    layer1_outputs(3801) <= a and not b;
    layer1_outputs(3802) <= b;
    layer1_outputs(3803) <= b and not a;
    layer1_outputs(3804) <= a;
    layer1_outputs(3805) <= not a or b;
    layer1_outputs(3806) <= not a or b;
    layer1_outputs(3807) <= 1'b1;
    layer1_outputs(3808) <= not a or b;
    layer1_outputs(3809) <= a and not b;
    layer1_outputs(3810) <= a and b;
    layer1_outputs(3811) <= not a;
    layer1_outputs(3812) <= a and not b;
    layer1_outputs(3813) <= not (a or b);
    layer1_outputs(3814) <= not b or a;
    layer1_outputs(3815) <= not (a or b);
    layer1_outputs(3816) <= not a;
    layer1_outputs(3817) <= b;
    layer1_outputs(3818) <= not a;
    layer1_outputs(3819) <= not (a xor b);
    layer1_outputs(3820) <= b and not a;
    layer1_outputs(3821) <= a or b;
    layer1_outputs(3822) <= a;
    layer1_outputs(3823) <= not b;
    layer1_outputs(3824) <= b and not a;
    layer1_outputs(3825) <= a and b;
    layer1_outputs(3826) <= a xor b;
    layer1_outputs(3827) <= 1'b1;
    layer1_outputs(3828) <= b;
    layer1_outputs(3829) <= not a or b;
    layer1_outputs(3830) <= 1'b0;
    layer1_outputs(3831) <= not (a and b);
    layer1_outputs(3832) <= b;
    layer1_outputs(3833) <= a xor b;
    layer1_outputs(3834) <= not (a and b);
    layer1_outputs(3835) <= a;
    layer1_outputs(3836) <= b and not a;
    layer1_outputs(3837) <= a or b;
    layer1_outputs(3838) <= not a or b;
    layer1_outputs(3839) <= not (a and b);
    layer1_outputs(3840) <= not (a or b);
    layer1_outputs(3841) <= not (a xor b);
    layer1_outputs(3842) <= not b;
    layer1_outputs(3843) <= not b;
    layer1_outputs(3844) <= not b;
    layer1_outputs(3845) <= a and not b;
    layer1_outputs(3846) <= not a or b;
    layer1_outputs(3847) <= not b;
    layer1_outputs(3848) <= not b or a;
    layer1_outputs(3849) <= not (a and b);
    layer1_outputs(3850) <= not (a xor b);
    layer1_outputs(3851) <= a and b;
    layer1_outputs(3852) <= b;
    layer1_outputs(3853) <= not b or a;
    layer1_outputs(3854) <= a and b;
    layer1_outputs(3855) <= 1'b1;
    layer1_outputs(3856) <= b and not a;
    layer1_outputs(3857) <= not (a or b);
    layer1_outputs(3858) <= 1'b0;
    layer1_outputs(3859) <= a and b;
    layer1_outputs(3860) <= a;
    layer1_outputs(3861) <= not (a and b);
    layer1_outputs(3862) <= b;
    layer1_outputs(3863) <= not (a or b);
    layer1_outputs(3864) <= not a;
    layer1_outputs(3865) <= not b;
    layer1_outputs(3866) <= not (a or b);
    layer1_outputs(3867) <= 1'b1;
    layer1_outputs(3868) <= a and b;
    layer1_outputs(3869) <= b and not a;
    layer1_outputs(3870) <= not (a xor b);
    layer1_outputs(3871) <= not (a or b);
    layer1_outputs(3872) <= b and not a;
    layer1_outputs(3873) <= b and not a;
    layer1_outputs(3874) <= not a or b;
    layer1_outputs(3875) <= a and b;
    layer1_outputs(3876) <= not a;
    layer1_outputs(3877) <= b;
    layer1_outputs(3878) <= a;
    layer1_outputs(3879) <= a and b;
    layer1_outputs(3880) <= not (a and b);
    layer1_outputs(3881) <= not (a xor b);
    layer1_outputs(3882) <= not b;
    layer1_outputs(3883) <= a or b;
    layer1_outputs(3884) <= b and not a;
    layer1_outputs(3885) <= not (a or b);
    layer1_outputs(3886) <= not a;
    layer1_outputs(3887) <= not b;
    layer1_outputs(3888) <= not (a and b);
    layer1_outputs(3889) <= not (a xor b);
    layer1_outputs(3890) <= not b or a;
    layer1_outputs(3891) <= not a;
    layer1_outputs(3892) <= not b or a;
    layer1_outputs(3893) <= a and b;
    layer1_outputs(3894) <= not b or a;
    layer1_outputs(3895) <= not (a xor b);
    layer1_outputs(3896) <= a xor b;
    layer1_outputs(3897) <= b and not a;
    layer1_outputs(3898) <= not b or a;
    layer1_outputs(3899) <= b and not a;
    layer1_outputs(3900) <= a and b;
    layer1_outputs(3901) <= a and not b;
    layer1_outputs(3902) <= not a;
    layer1_outputs(3903) <= not a or b;
    layer1_outputs(3904) <= b and not a;
    layer1_outputs(3905) <= a and b;
    layer1_outputs(3906) <= b;
    layer1_outputs(3907) <= not (a and b);
    layer1_outputs(3908) <= not b;
    layer1_outputs(3909) <= a;
    layer1_outputs(3910) <= b;
    layer1_outputs(3911) <= b;
    layer1_outputs(3912) <= not b;
    layer1_outputs(3913) <= a;
    layer1_outputs(3914) <= a or b;
    layer1_outputs(3915) <= not (a xor b);
    layer1_outputs(3916) <= not b;
    layer1_outputs(3917) <= not b;
    layer1_outputs(3918) <= a and not b;
    layer1_outputs(3919) <= b;
    layer1_outputs(3920) <= not a or b;
    layer1_outputs(3921) <= not (a xor b);
    layer1_outputs(3922) <= not (a or b);
    layer1_outputs(3923) <= not a;
    layer1_outputs(3924) <= not b or a;
    layer1_outputs(3925) <= a xor b;
    layer1_outputs(3926) <= a and not b;
    layer1_outputs(3927) <= b;
    layer1_outputs(3928) <= a and not b;
    layer1_outputs(3929) <= not a or b;
    layer1_outputs(3930) <= b and not a;
    layer1_outputs(3931) <= not a;
    layer1_outputs(3932) <= a xor b;
    layer1_outputs(3933) <= not b;
    layer1_outputs(3934) <= a;
    layer1_outputs(3935) <= 1'b0;
    layer1_outputs(3936) <= not b;
    layer1_outputs(3937) <= not b;
    layer1_outputs(3938) <= not b;
    layer1_outputs(3939) <= a and b;
    layer1_outputs(3940) <= b;
    layer1_outputs(3941) <= 1'b0;
    layer1_outputs(3942) <= b and not a;
    layer1_outputs(3943) <= b and not a;
    layer1_outputs(3944) <= a and not b;
    layer1_outputs(3945) <= not a or b;
    layer1_outputs(3946) <= a or b;
    layer1_outputs(3947) <= not (a xor b);
    layer1_outputs(3948) <= b and not a;
    layer1_outputs(3949) <= not (a xor b);
    layer1_outputs(3950) <= not (a or b);
    layer1_outputs(3951) <= b and not a;
    layer1_outputs(3952) <= not (a or b);
    layer1_outputs(3953) <= not b;
    layer1_outputs(3954) <= not (a or b);
    layer1_outputs(3955) <= not (a or b);
    layer1_outputs(3956) <= a and b;
    layer1_outputs(3957) <= a;
    layer1_outputs(3958) <= a and not b;
    layer1_outputs(3959) <= not a or b;
    layer1_outputs(3960) <= b;
    layer1_outputs(3961) <= b and not a;
    layer1_outputs(3962) <= not a;
    layer1_outputs(3963) <= not a;
    layer1_outputs(3964) <= not b or a;
    layer1_outputs(3965) <= not (a xor b);
    layer1_outputs(3966) <= not (a xor b);
    layer1_outputs(3967) <= not a;
    layer1_outputs(3968) <= a and not b;
    layer1_outputs(3969) <= not a;
    layer1_outputs(3970) <= a or b;
    layer1_outputs(3971) <= not b or a;
    layer1_outputs(3972) <= a;
    layer1_outputs(3973) <= a;
    layer1_outputs(3974) <= not b;
    layer1_outputs(3975) <= not a;
    layer1_outputs(3976) <= not (a or b);
    layer1_outputs(3977) <= b and not a;
    layer1_outputs(3978) <= not a or b;
    layer1_outputs(3979) <= 1'b1;
    layer1_outputs(3980) <= a and b;
    layer1_outputs(3981) <= not (a and b);
    layer1_outputs(3982) <= not (a xor b);
    layer1_outputs(3983) <= not b or a;
    layer1_outputs(3984) <= a and b;
    layer1_outputs(3985) <= a;
    layer1_outputs(3986) <= not b;
    layer1_outputs(3987) <= not b;
    layer1_outputs(3988) <= a;
    layer1_outputs(3989) <= b;
    layer1_outputs(3990) <= a or b;
    layer1_outputs(3991) <= not (a or b);
    layer1_outputs(3992) <= not (a or b);
    layer1_outputs(3993) <= not (a xor b);
    layer1_outputs(3994) <= not b;
    layer1_outputs(3995) <= not a;
    layer1_outputs(3996) <= b;
    layer1_outputs(3997) <= a;
    layer1_outputs(3998) <= a or b;
    layer1_outputs(3999) <= not a;
    layer1_outputs(4000) <= a;
    layer1_outputs(4001) <= a or b;
    layer1_outputs(4002) <= b and not a;
    layer1_outputs(4003) <= b;
    layer1_outputs(4004) <= not b;
    layer1_outputs(4005) <= not b;
    layer1_outputs(4006) <= a or b;
    layer1_outputs(4007) <= not a or b;
    layer1_outputs(4008) <= not (a or b);
    layer1_outputs(4009) <= not (a or b);
    layer1_outputs(4010) <= not b or a;
    layer1_outputs(4011) <= not a;
    layer1_outputs(4012) <= not b or a;
    layer1_outputs(4013) <= a xor b;
    layer1_outputs(4014) <= not (a and b);
    layer1_outputs(4015) <= b;
    layer1_outputs(4016) <= a;
    layer1_outputs(4017) <= a and b;
    layer1_outputs(4018) <= b;
    layer1_outputs(4019) <= not a or b;
    layer1_outputs(4020) <= not (a and b);
    layer1_outputs(4021) <= not a;
    layer1_outputs(4022) <= not (a xor b);
    layer1_outputs(4023) <= not (a xor b);
    layer1_outputs(4024) <= not b or a;
    layer1_outputs(4025) <= a xor b;
    layer1_outputs(4026) <= a and b;
    layer1_outputs(4027) <= a;
    layer1_outputs(4028) <= a and not b;
    layer1_outputs(4029) <= b and not a;
    layer1_outputs(4030) <= 1'b1;
    layer1_outputs(4031) <= a;
    layer1_outputs(4032) <= not (a and b);
    layer1_outputs(4033) <= not a;
    layer1_outputs(4034) <= not a or b;
    layer1_outputs(4035) <= a or b;
    layer1_outputs(4036) <= a and b;
    layer1_outputs(4037) <= not a or b;
    layer1_outputs(4038) <= a xor b;
    layer1_outputs(4039) <= a and b;
    layer1_outputs(4040) <= not (a or b);
    layer1_outputs(4041) <= not a or b;
    layer1_outputs(4042) <= not (a xor b);
    layer1_outputs(4043) <= b;
    layer1_outputs(4044) <= b;
    layer1_outputs(4045) <= not a;
    layer1_outputs(4046) <= not a;
    layer1_outputs(4047) <= a and b;
    layer1_outputs(4048) <= not a;
    layer1_outputs(4049) <= not b;
    layer1_outputs(4050) <= not (a or b);
    layer1_outputs(4051) <= b and not a;
    layer1_outputs(4052) <= not (a xor b);
    layer1_outputs(4053) <= not (a or b);
    layer1_outputs(4054) <= b and not a;
    layer1_outputs(4055) <= not b;
    layer1_outputs(4056) <= not (a or b);
    layer1_outputs(4057) <= a;
    layer1_outputs(4058) <= not b;
    layer1_outputs(4059) <= not a or b;
    layer1_outputs(4060) <= not (a xor b);
    layer1_outputs(4061) <= a and not b;
    layer1_outputs(4062) <= not a;
    layer1_outputs(4063) <= not (a xor b);
    layer1_outputs(4064) <= not b;
    layer1_outputs(4065) <= a or b;
    layer1_outputs(4066) <= b;
    layer1_outputs(4067) <= not a;
    layer1_outputs(4068) <= a and b;
    layer1_outputs(4069) <= 1'b0;
    layer1_outputs(4070) <= b;
    layer1_outputs(4071) <= a xor b;
    layer1_outputs(4072) <= b;
    layer1_outputs(4073) <= a and not b;
    layer1_outputs(4074) <= not a;
    layer1_outputs(4075) <= b;
    layer1_outputs(4076) <= not (a and b);
    layer1_outputs(4077) <= not b;
    layer1_outputs(4078) <= b;
    layer1_outputs(4079) <= b and not a;
    layer1_outputs(4080) <= a or b;
    layer1_outputs(4081) <= a;
    layer1_outputs(4082) <= a xor b;
    layer1_outputs(4083) <= not (a or b);
    layer1_outputs(4084) <= not (a or b);
    layer1_outputs(4085) <= a and b;
    layer1_outputs(4086) <= a and b;
    layer1_outputs(4087) <= b and not a;
    layer1_outputs(4088) <= a;
    layer1_outputs(4089) <= not b;
    layer1_outputs(4090) <= not b or a;
    layer1_outputs(4091) <= not (a and b);
    layer1_outputs(4092) <= a and b;
    layer1_outputs(4093) <= a xor b;
    layer1_outputs(4094) <= a xor b;
    layer1_outputs(4095) <= a and b;
    layer1_outputs(4096) <= a or b;
    layer1_outputs(4097) <= not a or b;
    layer1_outputs(4098) <= b and not a;
    layer1_outputs(4099) <= not (a xor b);
    layer1_outputs(4100) <= a;
    layer1_outputs(4101) <= a;
    layer1_outputs(4102) <= not (a or b);
    layer1_outputs(4103) <= not a or b;
    layer1_outputs(4104) <= not (a and b);
    layer1_outputs(4105) <= 1'b1;
    layer1_outputs(4106) <= not b or a;
    layer1_outputs(4107) <= a and b;
    layer1_outputs(4108) <= not b;
    layer1_outputs(4109) <= a xor b;
    layer1_outputs(4110) <= not (a and b);
    layer1_outputs(4111) <= b;
    layer1_outputs(4112) <= b;
    layer1_outputs(4113) <= a;
    layer1_outputs(4114) <= b;
    layer1_outputs(4115) <= a xor b;
    layer1_outputs(4116) <= b and not a;
    layer1_outputs(4117) <= b;
    layer1_outputs(4118) <= a and b;
    layer1_outputs(4119) <= not b;
    layer1_outputs(4120) <= a and b;
    layer1_outputs(4121) <= not (a and b);
    layer1_outputs(4122) <= not (a or b);
    layer1_outputs(4123) <= not b;
    layer1_outputs(4124) <= a and b;
    layer1_outputs(4125) <= a and b;
    layer1_outputs(4126) <= b;
    layer1_outputs(4127) <= 1'b0;
    layer1_outputs(4128) <= not b or a;
    layer1_outputs(4129) <= not (a and b);
    layer1_outputs(4130) <= b;
    layer1_outputs(4131) <= not b;
    layer1_outputs(4132) <= a;
    layer1_outputs(4133) <= a and not b;
    layer1_outputs(4134) <= a;
    layer1_outputs(4135) <= not a;
    layer1_outputs(4136) <= a and b;
    layer1_outputs(4137) <= not a;
    layer1_outputs(4138) <= not (a and b);
    layer1_outputs(4139) <= not b;
    layer1_outputs(4140) <= 1'b1;
    layer1_outputs(4141) <= a and not b;
    layer1_outputs(4142) <= not b or a;
    layer1_outputs(4143) <= not (a and b);
    layer1_outputs(4144) <= b and not a;
    layer1_outputs(4145) <= not b or a;
    layer1_outputs(4146) <= not (a xor b);
    layer1_outputs(4147) <= not (a and b);
    layer1_outputs(4148) <= a;
    layer1_outputs(4149) <= a or b;
    layer1_outputs(4150) <= a;
    layer1_outputs(4151) <= not b;
    layer1_outputs(4152) <= b and not a;
    layer1_outputs(4153) <= not (a and b);
    layer1_outputs(4154) <= a;
    layer1_outputs(4155) <= not b;
    layer1_outputs(4156) <= a;
    layer1_outputs(4157) <= a and b;
    layer1_outputs(4158) <= b and not a;
    layer1_outputs(4159) <= not b or a;
    layer1_outputs(4160) <= not a;
    layer1_outputs(4161) <= a;
    layer1_outputs(4162) <= not (a or b);
    layer1_outputs(4163) <= not b or a;
    layer1_outputs(4164) <= not b or a;
    layer1_outputs(4165) <= a xor b;
    layer1_outputs(4166) <= b and not a;
    layer1_outputs(4167) <= a and b;
    layer1_outputs(4168) <= a or b;
    layer1_outputs(4169) <= not b or a;
    layer1_outputs(4170) <= not a;
    layer1_outputs(4171) <= not (a and b);
    layer1_outputs(4172) <= a xor b;
    layer1_outputs(4173) <= not b;
    layer1_outputs(4174) <= a xor b;
    layer1_outputs(4175) <= not (a xor b);
    layer1_outputs(4176) <= a and b;
    layer1_outputs(4177) <= a xor b;
    layer1_outputs(4178) <= not (a or b);
    layer1_outputs(4179) <= not b or a;
    layer1_outputs(4180) <= a;
    layer1_outputs(4181) <= not b or a;
    layer1_outputs(4182) <= not a or b;
    layer1_outputs(4183) <= a and not b;
    layer1_outputs(4184) <= a xor b;
    layer1_outputs(4185) <= not b;
    layer1_outputs(4186) <= not a;
    layer1_outputs(4187) <= a xor b;
    layer1_outputs(4188) <= not b;
    layer1_outputs(4189) <= a xor b;
    layer1_outputs(4190) <= not a;
    layer1_outputs(4191) <= not a;
    layer1_outputs(4192) <= not b or a;
    layer1_outputs(4193) <= not (a or b);
    layer1_outputs(4194) <= not a;
    layer1_outputs(4195) <= not a or b;
    layer1_outputs(4196) <= a or b;
    layer1_outputs(4197) <= not a;
    layer1_outputs(4198) <= a;
    layer1_outputs(4199) <= not (a and b);
    layer1_outputs(4200) <= b and not a;
    layer1_outputs(4201) <= not (a and b);
    layer1_outputs(4202) <= not (a and b);
    layer1_outputs(4203) <= a and not b;
    layer1_outputs(4204) <= a or b;
    layer1_outputs(4205) <= not a;
    layer1_outputs(4206) <= a or b;
    layer1_outputs(4207) <= a;
    layer1_outputs(4208) <= not a;
    layer1_outputs(4209) <= b;
    layer1_outputs(4210) <= a;
    layer1_outputs(4211) <= 1'b0;
    layer1_outputs(4212) <= not (a and b);
    layer1_outputs(4213) <= not b or a;
    layer1_outputs(4214) <= not a or b;
    layer1_outputs(4215) <= a;
    layer1_outputs(4216) <= not (a xor b);
    layer1_outputs(4217) <= not (a and b);
    layer1_outputs(4218) <= b and not a;
    layer1_outputs(4219) <= a or b;
    layer1_outputs(4220) <= a or b;
    layer1_outputs(4221) <= b;
    layer1_outputs(4222) <= 1'b1;
    layer1_outputs(4223) <= b;
    layer1_outputs(4224) <= a;
    layer1_outputs(4225) <= a;
    layer1_outputs(4226) <= 1'b1;
    layer1_outputs(4227) <= a and not b;
    layer1_outputs(4228) <= b;
    layer1_outputs(4229) <= not (a and b);
    layer1_outputs(4230) <= a and b;
    layer1_outputs(4231) <= a;
    layer1_outputs(4232) <= not b;
    layer1_outputs(4233) <= not b;
    layer1_outputs(4234) <= not a or b;
    layer1_outputs(4235) <= not a or b;
    layer1_outputs(4236) <= not a;
    layer1_outputs(4237) <= not a or b;
    layer1_outputs(4238) <= a xor b;
    layer1_outputs(4239) <= b;
    layer1_outputs(4240) <= not a or b;
    layer1_outputs(4241) <= b;
    layer1_outputs(4242) <= not b or a;
    layer1_outputs(4243) <= a or b;
    layer1_outputs(4244) <= a or b;
    layer1_outputs(4245) <= a and not b;
    layer1_outputs(4246) <= 1'b0;
    layer1_outputs(4247) <= a xor b;
    layer1_outputs(4248) <= a;
    layer1_outputs(4249) <= not a;
    layer1_outputs(4250) <= a and b;
    layer1_outputs(4251) <= not (a or b);
    layer1_outputs(4252) <= not a;
    layer1_outputs(4253) <= a;
    layer1_outputs(4254) <= a or b;
    layer1_outputs(4255) <= not a or b;
    layer1_outputs(4256) <= a and b;
    layer1_outputs(4257) <= b and not a;
    layer1_outputs(4258) <= a and b;
    layer1_outputs(4259) <= a and not b;
    layer1_outputs(4260) <= a;
    layer1_outputs(4261) <= not (a xor b);
    layer1_outputs(4262) <= b and not a;
    layer1_outputs(4263) <= not (a or b);
    layer1_outputs(4264) <= not (a xor b);
    layer1_outputs(4265) <= not (a xor b);
    layer1_outputs(4266) <= b;
    layer1_outputs(4267) <= a;
    layer1_outputs(4268) <= not b or a;
    layer1_outputs(4269) <= not a or b;
    layer1_outputs(4270) <= not (a or b);
    layer1_outputs(4271) <= a or b;
    layer1_outputs(4272) <= b;
    layer1_outputs(4273) <= not (a and b);
    layer1_outputs(4274) <= a and b;
    layer1_outputs(4275) <= a xor b;
    layer1_outputs(4276) <= a and b;
    layer1_outputs(4277) <= a xor b;
    layer1_outputs(4278) <= b and not a;
    layer1_outputs(4279) <= a;
    layer1_outputs(4280) <= not a or b;
    layer1_outputs(4281) <= not (a and b);
    layer1_outputs(4282) <= b;
    layer1_outputs(4283) <= not a or b;
    layer1_outputs(4284) <= not a or b;
    layer1_outputs(4285) <= a and b;
    layer1_outputs(4286) <= not (a and b);
    layer1_outputs(4287) <= b and not a;
    layer1_outputs(4288) <= a or b;
    layer1_outputs(4289) <= a and b;
    layer1_outputs(4290) <= not b or a;
    layer1_outputs(4291) <= not a;
    layer1_outputs(4292) <= not a;
    layer1_outputs(4293) <= not a;
    layer1_outputs(4294) <= not b or a;
    layer1_outputs(4295) <= a xor b;
    layer1_outputs(4296) <= not (a or b);
    layer1_outputs(4297) <= not b or a;
    layer1_outputs(4298) <= a;
    layer1_outputs(4299) <= not a;
    layer1_outputs(4300) <= b;
    layer1_outputs(4301) <= a and not b;
    layer1_outputs(4302) <= a;
    layer1_outputs(4303) <= not a or b;
    layer1_outputs(4304) <= not b;
    layer1_outputs(4305) <= not (a and b);
    layer1_outputs(4306) <= a;
    layer1_outputs(4307) <= b and not a;
    layer1_outputs(4308) <= b;
    layer1_outputs(4309) <= not a or b;
    layer1_outputs(4310) <= a or b;
    layer1_outputs(4311) <= a xor b;
    layer1_outputs(4312) <= not (a and b);
    layer1_outputs(4313) <= a;
    layer1_outputs(4314) <= a or b;
    layer1_outputs(4315) <= b;
    layer1_outputs(4316) <= a and not b;
    layer1_outputs(4317) <= a;
    layer1_outputs(4318) <= not a;
    layer1_outputs(4319) <= not a;
    layer1_outputs(4320) <= a;
    layer1_outputs(4321) <= a xor b;
    layer1_outputs(4322) <= not a;
    layer1_outputs(4323) <= b;
    layer1_outputs(4324) <= not (a xor b);
    layer1_outputs(4325) <= not (a xor b);
    layer1_outputs(4326) <= b;
    layer1_outputs(4327) <= a xor b;
    layer1_outputs(4328) <= not b or a;
    layer1_outputs(4329) <= a;
    layer1_outputs(4330) <= a xor b;
    layer1_outputs(4331) <= a or b;
    layer1_outputs(4332) <= not (a and b);
    layer1_outputs(4333) <= not b;
    layer1_outputs(4334) <= b;
    layer1_outputs(4335) <= not a or b;
    layer1_outputs(4336) <= not b;
    layer1_outputs(4337) <= a xor b;
    layer1_outputs(4338) <= b;
    layer1_outputs(4339) <= not a;
    layer1_outputs(4340) <= b;
    layer1_outputs(4341) <= a xor b;
    layer1_outputs(4342) <= a and b;
    layer1_outputs(4343) <= a and not b;
    layer1_outputs(4344) <= not (a or b);
    layer1_outputs(4345) <= b;
    layer1_outputs(4346) <= not (a and b);
    layer1_outputs(4347) <= not (a and b);
    layer1_outputs(4348) <= not b;
    layer1_outputs(4349) <= not a;
    layer1_outputs(4350) <= a;
    layer1_outputs(4351) <= not b or a;
    layer1_outputs(4352) <= b;
    layer1_outputs(4353) <= a xor b;
    layer1_outputs(4354) <= not b;
    layer1_outputs(4355) <= not b;
    layer1_outputs(4356) <= a;
    layer1_outputs(4357) <= b;
    layer1_outputs(4358) <= not b;
    layer1_outputs(4359) <= not a;
    layer1_outputs(4360) <= 1'b0;
    layer1_outputs(4361) <= not a;
    layer1_outputs(4362) <= a;
    layer1_outputs(4363) <= a and b;
    layer1_outputs(4364) <= not a or b;
    layer1_outputs(4365) <= not a or b;
    layer1_outputs(4366) <= a xor b;
    layer1_outputs(4367) <= not a;
    layer1_outputs(4368) <= a or b;
    layer1_outputs(4369) <= a;
    layer1_outputs(4370) <= 1'b1;
    layer1_outputs(4371) <= not a or b;
    layer1_outputs(4372) <= a;
    layer1_outputs(4373) <= a;
    layer1_outputs(4374) <= not a or b;
    layer1_outputs(4375) <= a and b;
    layer1_outputs(4376) <= not a or b;
    layer1_outputs(4377) <= a;
    layer1_outputs(4378) <= a and b;
    layer1_outputs(4379) <= a or b;
    layer1_outputs(4380) <= a;
    layer1_outputs(4381) <= not b;
    layer1_outputs(4382) <= not a or b;
    layer1_outputs(4383) <= b;
    layer1_outputs(4384) <= not b;
    layer1_outputs(4385) <= b and not a;
    layer1_outputs(4386) <= not b or a;
    layer1_outputs(4387) <= a or b;
    layer1_outputs(4388) <= not a or b;
    layer1_outputs(4389) <= not b or a;
    layer1_outputs(4390) <= a and not b;
    layer1_outputs(4391) <= not (a and b);
    layer1_outputs(4392) <= not (a or b);
    layer1_outputs(4393) <= not b or a;
    layer1_outputs(4394) <= not b or a;
    layer1_outputs(4395) <= not a;
    layer1_outputs(4396) <= not b;
    layer1_outputs(4397) <= not b or a;
    layer1_outputs(4398) <= a;
    layer1_outputs(4399) <= a and not b;
    layer1_outputs(4400) <= a xor b;
    layer1_outputs(4401) <= not (a xor b);
    layer1_outputs(4402) <= a or b;
    layer1_outputs(4403) <= a or b;
    layer1_outputs(4404) <= not (a or b);
    layer1_outputs(4405) <= not a;
    layer1_outputs(4406) <= b;
    layer1_outputs(4407) <= not b;
    layer1_outputs(4408) <= not a;
    layer1_outputs(4409) <= not (a or b);
    layer1_outputs(4410) <= b;
    layer1_outputs(4411) <= not (a and b);
    layer1_outputs(4412) <= a;
    layer1_outputs(4413) <= b;
    layer1_outputs(4414) <= not (a xor b);
    layer1_outputs(4415) <= a and not b;
    layer1_outputs(4416) <= not a or b;
    layer1_outputs(4417) <= a and b;
    layer1_outputs(4418) <= not (a and b);
    layer1_outputs(4419) <= a and not b;
    layer1_outputs(4420) <= not a;
    layer1_outputs(4421) <= not b;
    layer1_outputs(4422) <= not (a or b);
    layer1_outputs(4423) <= not b or a;
    layer1_outputs(4424) <= not a;
    layer1_outputs(4425) <= a and not b;
    layer1_outputs(4426) <= not (a or b);
    layer1_outputs(4427) <= not (a xor b);
    layer1_outputs(4428) <= a xor b;
    layer1_outputs(4429) <= a and b;
    layer1_outputs(4430) <= a and not b;
    layer1_outputs(4431) <= b and not a;
    layer1_outputs(4432) <= a;
    layer1_outputs(4433) <= 1'b1;
    layer1_outputs(4434) <= not b;
    layer1_outputs(4435) <= a or b;
    layer1_outputs(4436) <= 1'b0;
    layer1_outputs(4437) <= a;
    layer1_outputs(4438) <= b;
    layer1_outputs(4439) <= not (a and b);
    layer1_outputs(4440) <= not a or b;
    layer1_outputs(4441) <= b and not a;
    layer1_outputs(4442) <= not a or b;
    layer1_outputs(4443) <= a and b;
    layer1_outputs(4444) <= not (a or b);
    layer1_outputs(4445) <= b;
    layer1_outputs(4446) <= not (a and b);
    layer1_outputs(4447) <= 1'b1;
    layer1_outputs(4448) <= a and not b;
    layer1_outputs(4449) <= a and not b;
    layer1_outputs(4450) <= not a;
    layer1_outputs(4451) <= a and b;
    layer1_outputs(4452) <= a xor b;
    layer1_outputs(4453) <= a;
    layer1_outputs(4454) <= not b or a;
    layer1_outputs(4455) <= not b;
    layer1_outputs(4456) <= not a or b;
    layer1_outputs(4457) <= not b or a;
    layer1_outputs(4458) <= a and b;
    layer1_outputs(4459) <= not b;
    layer1_outputs(4460) <= not a or b;
    layer1_outputs(4461) <= b;
    layer1_outputs(4462) <= b;
    layer1_outputs(4463) <= a and b;
    layer1_outputs(4464) <= not (a xor b);
    layer1_outputs(4465) <= a and b;
    layer1_outputs(4466) <= not a or b;
    layer1_outputs(4467) <= not a or b;
    layer1_outputs(4468) <= not (a and b);
    layer1_outputs(4469) <= not (a or b);
    layer1_outputs(4470) <= b and not a;
    layer1_outputs(4471) <= not a;
    layer1_outputs(4472) <= not a;
    layer1_outputs(4473) <= b;
    layer1_outputs(4474) <= not (a and b);
    layer1_outputs(4475) <= not b or a;
    layer1_outputs(4476) <= a or b;
    layer1_outputs(4477) <= b and not a;
    layer1_outputs(4478) <= not a;
    layer1_outputs(4479) <= b;
    layer1_outputs(4480) <= a;
    layer1_outputs(4481) <= a;
    layer1_outputs(4482) <= a;
    layer1_outputs(4483) <= not (a and b);
    layer1_outputs(4484) <= a and b;
    layer1_outputs(4485) <= b;
    layer1_outputs(4486) <= a and not b;
    layer1_outputs(4487) <= a and b;
    layer1_outputs(4488) <= not (a and b);
    layer1_outputs(4489) <= a xor b;
    layer1_outputs(4490) <= not a or b;
    layer1_outputs(4491) <= b;
    layer1_outputs(4492) <= a and b;
    layer1_outputs(4493) <= not (a xor b);
    layer1_outputs(4494) <= a and b;
    layer1_outputs(4495) <= b and not a;
    layer1_outputs(4496) <= a and not b;
    layer1_outputs(4497) <= not (a and b);
    layer1_outputs(4498) <= not (a or b);
    layer1_outputs(4499) <= 1'b0;
    layer1_outputs(4500) <= not b or a;
    layer1_outputs(4501) <= not (a or b);
    layer1_outputs(4502) <= not b or a;
    layer1_outputs(4503) <= not (a or b);
    layer1_outputs(4504) <= not b or a;
    layer1_outputs(4505) <= b;
    layer1_outputs(4506) <= not (a and b);
    layer1_outputs(4507) <= b;
    layer1_outputs(4508) <= b;
    layer1_outputs(4509) <= not b;
    layer1_outputs(4510) <= not (a xor b);
    layer1_outputs(4511) <= a and b;
    layer1_outputs(4512) <= not b;
    layer1_outputs(4513) <= not b;
    layer1_outputs(4514) <= a or b;
    layer1_outputs(4515) <= not (a or b);
    layer1_outputs(4516) <= a;
    layer1_outputs(4517) <= 1'b1;
    layer1_outputs(4518) <= b;
    layer1_outputs(4519) <= not (a or b);
    layer1_outputs(4520) <= a or b;
    layer1_outputs(4521) <= a;
    layer1_outputs(4522) <= a and b;
    layer1_outputs(4523) <= b;
    layer1_outputs(4524) <= b;
    layer1_outputs(4525) <= 1'b0;
    layer1_outputs(4526) <= a and b;
    layer1_outputs(4527) <= 1'b0;
    layer1_outputs(4528) <= not a;
    layer1_outputs(4529) <= not b or a;
    layer1_outputs(4530) <= a;
    layer1_outputs(4531) <= not b;
    layer1_outputs(4532) <= a xor b;
    layer1_outputs(4533) <= not (a xor b);
    layer1_outputs(4534) <= not b;
    layer1_outputs(4535) <= a and not b;
    layer1_outputs(4536) <= not (a or b);
    layer1_outputs(4537) <= 1'b0;
    layer1_outputs(4538) <= b;
    layer1_outputs(4539) <= a;
    layer1_outputs(4540) <= not (a or b);
    layer1_outputs(4541) <= a and not b;
    layer1_outputs(4542) <= not b;
    layer1_outputs(4543) <= b;
    layer1_outputs(4544) <= a and not b;
    layer1_outputs(4545) <= not (a xor b);
    layer1_outputs(4546) <= not (a xor b);
    layer1_outputs(4547) <= a;
    layer1_outputs(4548) <= not b;
    layer1_outputs(4549) <= not (a xor b);
    layer1_outputs(4550) <= a or b;
    layer1_outputs(4551) <= a and not b;
    layer1_outputs(4552) <= a and b;
    layer1_outputs(4553) <= not (a or b);
    layer1_outputs(4554) <= not (a and b);
    layer1_outputs(4555) <= not b or a;
    layer1_outputs(4556) <= b;
    layer1_outputs(4557) <= a;
    layer1_outputs(4558) <= not (a and b);
    layer1_outputs(4559) <= a xor b;
    layer1_outputs(4560) <= a;
    layer1_outputs(4561) <= not b;
    layer1_outputs(4562) <= b and not a;
    layer1_outputs(4563) <= not a;
    layer1_outputs(4564) <= not b;
    layer1_outputs(4565) <= not (a and b);
    layer1_outputs(4566) <= a;
    layer1_outputs(4567) <= not (a or b);
    layer1_outputs(4568) <= b;
    layer1_outputs(4569) <= not (a and b);
    layer1_outputs(4570) <= a and b;
    layer1_outputs(4571) <= not (a xor b);
    layer1_outputs(4572) <= not (a xor b);
    layer1_outputs(4573) <= a and not b;
    layer1_outputs(4574) <= not (a or b);
    layer1_outputs(4575) <= a and not b;
    layer1_outputs(4576) <= a xor b;
    layer1_outputs(4577) <= a and not b;
    layer1_outputs(4578) <= b and not a;
    layer1_outputs(4579) <= not b;
    layer1_outputs(4580) <= a and not b;
    layer1_outputs(4581) <= not a;
    layer1_outputs(4582) <= not (a and b);
    layer1_outputs(4583) <= not a;
    layer1_outputs(4584) <= b;
    layer1_outputs(4585) <= not (a and b);
    layer1_outputs(4586) <= not b or a;
    layer1_outputs(4587) <= a and not b;
    layer1_outputs(4588) <= b and not a;
    layer1_outputs(4589) <= a or b;
    layer1_outputs(4590) <= b and not a;
    layer1_outputs(4591) <= not a;
    layer1_outputs(4592) <= not b;
    layer1_outputs(4593) <= not b;
    layer1_outputs(4594) <= b;
    layer1_outputs(4595) <= a and not b;
    layer1_outputs(4596) <= b;
    layer1_outputs(4597) <= not (a or b);
    layer1_outputs(4598) <= not b;
    layer1_outputs(4599) <= not (a and b);
    layer1_outputs(4600) <= a and not b;
    layer1_outputs(4601) <= a;
    layer1_outputs(4602) <= 1'b0;
    layer1_outputs(4603) <= not a;
    layer1_outputs(4604) <= a and not b;
    layer1_outputs(4605) <= not a;
    layer1_outputs(4606) <= not a or b;
    layer1_outputs(4607) <= not (a xor b);
    layer1_outputs(4608) <= b;
    layer1_outputs(4609) <= a and b;
    layer1_outputs(4610) <= not a;
    layer1_outputs(4611) <= not a;
    layer1_outputs(4612) <= not (a or b);
    layer1_outputs(4613) <= b;
    layer1_outputs(4614) <= a and not b;
    layer1_outputs(4615) <= a;
    layer1_outputs(4616) <= not b;
    layer1_outputs(4617) <= b;
    layer1_outputs(4618) <= b;
    layer1_outputs(4619) <= a and not b;
    layer1_outputs(4620) <= not (a or b);
    layer1_outputs(4621) <= b and not a;
    layer1_outputs(4622) <= b;
    layer1_outputs(4623) <= a;
    layer1_outputs(4624) <= b and not a;
    layer1_outputs(4625) <= not b;
    layer1_outputs(4626) <= not (a and b);
    layer1_outputs(4627) <= not b;
    layer1_outputs(4628) <= b;
    layer1_outputs(4629) <= not b;
    layer1_outputs(4630) <= not (a or b);
    layer1_outputs(4631) <= not b;
    layer1_outputs(4632) <= not b or a;
    layer1_outputs(4633) <= not a;
    layer1_outputs(4634) <= b;
    layer1_outputs(4635) <= a and b;
    layer1_outputs(4636) <= not (a xor b);
    layer1_outputs(4637) <= 1'b0;
    layer1_outputs(4638) <= a xor b;
    layer1_outputs(4639) <= not a or b;
    layer1_outputs(4640) <= b;
    layer1_outputs(4641) <= 1'b0;
    layer1_outputs(4642) <= a xor b;
    layer1_outputs(4643) <= a xor b;
    layer1_outputs(4644) <= not a or b;
    layer1_outputs(4645) <= not b;
    layer1_outputs(4646) <= a and b;
    layer1_outputs(4647) <= a;
    layer1_outputs(4648) <= a and not b;
    layer1_outputs(4649) <= a or b;
    layer1_outputs(4650) <= a or b;
    layer1_outputs(4651) <= not (a xor b);
    layer1_outputs(4652) <= a and b;
    layer1_outputs(4653) <= not (a or b);
    layer1_outputs(4654) <= not (a or b);
    layer1_outputs(4655) <= 1'b1;
    layer1_outputs(4656) <= not (a and b);
    layer1_outputs(4657) <= a or b;
    layer1_outputs(4658) <= not b;
    layer1_outputs(4659) <= 1'b1;
    layer1_outputs(4660) <= a and b;
    layer1_outputs(4661) <= a and b;
    layer1_outputs(4662) <= not (a or b);
    layer1_outputs(4663) <= a and b;
    layer1_outputs(4664) <= a;
    layer1_outputs(4665) <= not (a or b);
    layer1_outputs(4666) <= not b or a;
    layer1_outputs(4667) <= not b or a;
    layer1_outputs(4668) <= b;
    layer1_outputs(4669) <= not a or b;
    layer1_outputs(4670) <= b and not a;
    layer1_outputs(4671) <= not a;
    layer1_outputs(4672) <= b and not a;
    layer1_outputs(4673) <= not b;
    layer1_outputs(4674) <= a xor b;
    layer1_outputs(4675) <= a xor b;
    layer1_outputs(4676) <= not b or a;
    layer1_outputs(4677) <= a xor b;
    layer1_outputs(4678) <= not b or a;
    layer1_outputs(4679) <= not b;
    layer1_outputs(4680) <= a or b;
    layer1_outputs(4681) <= b and not a;
    layer1_outputs(4682) <= a xor b;
    layer1_outputs(4683) <= a and not b;
    layer1_outputs(4684) <= not (a xor b);
    layer1_outputs(4685) <= not (a and b);
    layer1_outputs(4686) <= a xor b;
    layer1_outputs(4687) <= not b;
    layer1_outputs(4688) <= a and not b;
    layer1_outputs(4689) <= b and not a;
    layer1_outputs(4690) <= a and not b;
    layer1_outputs(4691) <= a and b;
    layer1_outputs(4692) <= not a;
    layer1_outputs(4693) <= a xor b;
    layer1_outputs(4694) <= not (a and b);
    layer1_outputs(4695) <= b and not a;
    layer1_outputs(4696) <= not a;
    layer1_outputs(4697) <= a and b;
    layer1_outputs(4698) <= not a;
    layer1_outputs(4699) <= not b or a;
    layer1_outputs(4700) <= a;
    layer1_outputs(4701) <= a or b;
    layer1_outputs(4702) <= not b or a;
    layer1_outputs(4703) <= not a or b;
    layer1_outputs(4704) <= not b;
    layer1_outputs(4705) <= not a or b;
    layer1_outputs(4706) <= not b or a;
    layer1_outputs(4707) <= b and not a;
    layer1_outputs(4708) <= not b;
    layer1_outputs(4709) <= b;
    layer1_outputs(4710) <= a xor b;
    layer1_outputs(4711) <= b and not a;
    layer1_outputs(4712) <= not a or b;
    layer1_outputs(4713) <= b;
    layer1_outputs(4714) <= not a or b;
    layer1_outputs(4715) <= a and b;
    layer1_outputs(4716) <= a and b;
    layer1_outputs(4717) <= b;
    layer1_outputs(4718) <= a xor b;
    layer1_outputs(4719) <= b and not a;
    layer1_outputs(4720) <= a or b;
    layer1_outputs(4721) <= not (a xor b);
    layer1_outputs(4722) <= a;
    layer1_outputs(4723) <= a;
    layer1_outputs(4724) <= b and not a;
    layer1_outputs(4725) <= b and not a;
    layer1_outputs(4726) <= not (a or b);
    layer1_outputs(4727) <= not b;
    layer1_outputs(4728) <= a and not b;
    layer1_outputs(4729) <= not a or b;
    layer1_outputs(4730) <= not (a or b);
    layer1_outputs(4731) <= not b or a;
    layer1_outputs(4732) <= not a;
    layer1_outputs(4733) <= not a or b;
    layer1_outputs(4734) <= b;
    layer1_outputs(4735) <= b;
    layer1_outputs(4736) <= not (a xor b);
    layer1_outputs(4737) <= a xor b;
    layer1_outputs(4738) <= a and b;
    layer1_outputs(4739) <= not a;
    layer1_outputs(4740) <= a;
    layer1_outputs(4741) <= 1'b0;
    layer1_outputs(4742) <= not (a or b);
    layer1_outputs(4743) <= a and b;
    layer1_outputs(4744) <= a xor b;
    layer1_outputs(4745) <= b;
    layer1_outputs(4746) <= not (a xor b);
    layer1_outputs(4747) <= not a;
    layer1_outputs(4748) <= a or b;
    layer1_outputs(4749) <= not b;
    layer1_outputs(4750) <= a;
    layer1_outputs(4751) <= b and not a;
    layer1_outputs(4752) <= not a;
    layer1_outputs(4753) <= a xor b;
    layer1_outputs(4754) <= not a;
    layer1_outputs(4755) <= not a;
    layer1_outputs(4756) <= a xor b;
    layer1_outputs(4757) <= not (a or b);
    layer1_outputs(4758) <= a;
    layer1_outputs(4759) <= not a or b;
    layer1_outputs(4760) <= not b or a;
    layer1_outputs(4761) <= b;
    layer1_outputs(4762) <= not b or a;
    layer1_outputs(4763) <= a xor b;
    layer1_outputs(4764) <= a;
    layer1_outputs(4765) <= b;
    layer1_outputs(4766) <= not (a and b);
    layer1_outputs(4767) <= not b;
    layer1_outputs(4768) <= b;
    layer1_outputs(4769) <= a and not b;
    layer1_outputs(4770) <= b and not a;
    layer1_outputs(4771) <= a;
    layer1_outputs(4772) <= b and not a;
    layer1_outputs(4773) <= not b or a;
    layer1_outputs(4774) <= not (a xor b);
    layer1_outputs(4775) <= a;
    layer1_outputs(4776) <= not (a or b);
    layer1_outputs(4777) <= b and not a;
    layer1_outputs(4778) <= not a or b;
    layer1_outputs(4779) <= not b;
    layer1_outputs(4780) <= a and not b;
    layer1_outputs(4781) <= a and b;
    layer1_outputs(4782) <= not (a xor b);
    layer1_outputs(4783) <= not (a xor b);
    layer1_outputs(4784) <= not (a xor b);
    layer1_outputs(4785) <= not a;
    layer1_outputs(4786) <= not a;
    layer1_outputs(4787) <= not (a xor b);
    layer1_outputs(4788) <= a xor b;
    layer1_outputs(4789) <= a and b;
    layer1_outputs(4790) <= not b;
    layer1_outputs(4791) <= not (a xor b);
    layer1_outputs(4792) <= not a;
    layer1_outputs(4793) <= not b;
    layer1_outputs(4794) <= a xor b;
    layer1_outputs(4795) <= a;
    layer1_outputs(4796) <= a;
    layer1_outputs(4797) <= a and b;
    layer1_outputs(4798) <= a xor b;
    layer1_outputs(4799) <= a or b;
    layer1_outputs(4800) <= not (a or b);
    layer1_outputs(4801) <= a and not b;
    layer1_outputs(4802) <= not a;
    layer1_outputs(4803) <= a and not b;
    layer1_outputs(4804) <= a;
    layer1_outputs(4805) <= not (a or b);
    layer1_outputs(4806) <= not (a xor b);
    layer1_outputs(4807) <= not a;
    layer1_outputs(4808) <= b;
    layer1_outputs(4809) <= b and not a;
    layer1_outputs(4810) <= not (a xor b);
    layer1_outputs(4811) <= not (a or b);
    layer1_outputs(4812) <= a;
    layer1_outputs(4813) <= b;
    layer1_outputs(4814) <= not a or b;
    layer1_outputs(4815) <= a or b;
    layer1_outputs(4816) <= a and not b;
    layer1_outputs(4817) <= not b;
    layer1_outputs(4818) <= not b or a;
    layer1_outputs(4819) <= a xor b;
    layer1_outputs(4820) <= not b or a;
    layer1_outputs(4821) <= not b or a;
    layer1_outputs(4822) <= a xor b;
    layer1_outputs(4823) <= a and not b;
    layer1_outputs(4824) <= a;
    layer1_outputs(4825) <= a or b;
    layer1_outputs(4826) <= not (a xor b);
    layer1_outputs(4827) <= b;
    layer1_outputs(4828) <= a xor b;
    layer1_outputs(4829) <= not (a and b);
    layer1_outputs(4830) <= not b;
    layer1_outputs(4831) <= not (a or b);
    layer1_outputs(4832) <= a and b;
    layer1_outputs(4833) <= a or b;
    layer1_outputs(4834) <= b and not a;
    layer1_outputs(4835) <= not (a xor b);
    layer1_outputs(4836) <= not (a xor b);
    layer1_outputs(4837) <= not a;
    layer1_outputs(4838) <= not b;
    layer1_outputs(4839) <= a or b;
    layer1_outputs(4840) <= a or b;
    layer1_outputs(4841) <= 1'b1;
    layer1_outputs(4842) <= not (a or b);
    layer1_outputs(4843) <= not (a or b);
    layer1_outputs(4844) <= not b;
    layer1_outputs(4845) <= a or b;
    layer1_outputs(4846) <= not a;
    layer1_outputs(4847) <= not b;
    layer1_outputs(4848) <= a;
    layer1_outputs(4849) <= not b;
    layer1_outputs(4850) <= not b;
    layer1_outputs(4851) <= a or b;
    layer1_outputs(4852) <= a xor b;
    layer1_outputs(4853) <= not a or b;
    layer1_outputs(4854) <= not b or a;
    layer1_outputs(4855) <= not b or a;
    layer1_outputs(4856) <= a and not b;
    layer1_outputs(4857) <= a and not b;
    layer1_outputs(4858) <= a and b;
    layer1_outputs(4859) <= a and not b;
    layer1_outputs(4860) <= not (a or b);
    layer1_outputs(4861) <= a;
    layer1_outputs(4862) <= a and b;
    layer1_outputs(4863) <= a and b;
    layer1_outputs(4864) <= not b;
    layer1_outputs(4865) <= b;
    layer1_outputs(4866) <= a and b;
    layer1_outputs(4867) <= not b or a;
    layer1_outputs(4868) <= a or b;
    layer1_outputs(4869) <= b;
    layer1_outputs(4870) <= not a or b;
    layer1_outputs(4871) <= not a or b;
    layer1_outputs(4872) <= not a;
    layer1_outputs(4873) <= a;
    layer1_outputs(4874) <= a and not b;
    layer1_outputs(4875) <= a and not b;
    layer1_outputs(4876) <= not b;
    layer1_outputs(4877) <= not a or b;
    layer1_outputs(4878) <= not (a and b);
    layer1_outputs(4879) <= not b;
    layer1_outputs(4880) <= a or b;
    layer1_outputs(4881) <= a;
    layer1_outputs(4882) <= b and not a;
    layer1_outputs(4883) <= not b;
    layer1_outputs(4884) <= b;
    layer1_outputs(4885) <= b;
    layer1_outputs(4886) <= not (a xor b);
    layer1_outputs(4887) <= a;
    layer1_outputs(4888) <= not (a and b);
    layer1_outputs(4889) <= b;
    layer1_outputs(4890) <= not b or a;
    layer1_outputs(4891) <= a;
    layer1_outputs(4892) <= a or b;
    layer1_outputs(4893) <= not b;
    layer1_outputs(4894) <= not b or a;
    layer1_outputs(4895) <= a xor b;
    layer1_outputs(4896) <= not (a xor b);
    layer1_outputs(4897) <= b and not a;
    layer1_outputs(4898) <= a;
    layer1_outputs(4899) <= a xor b;
    layer1_outputs(4900) <= a and not b;
    layer1_outputs(4901) <= a and b;
    layer1_outputs(4902) <= not b;
    layer1_outputs(4903) <= a xor b;
    layer1_outputs(4904) <= not b;
    layer1_outputs(4905) <= a;
    layer1_outputs(4906) <= b;
    layer1_outputs(4907) <= 1'b0;
    layer1_outputs(4908) <= not a or b;
    layer1_outputs(4909) <= not (a or b);
    layer1_outputs(4910) <= not b or a;
    layer1_outputs(4911) <= b and not a;
    layer1_outputs(4912) <= a and not b;
    layer1_outputs(4913) <= a and b;
    layer1_outputs(4914) <= not (a or b);
    layer1_outputs(4915) <= not b;
    layer1_outputs(4916) <= not a or b;
    layer1_outputs(4917) <= a;
    layer1_outputs(4918) <= not a or b;
    layer1_outputs(4919) <= 1'b1;
    layer1_outputs(4920) <= a xor b;
    layer1_outputs(4921) <= a;
    layer1_outputs(4922) <= a or b;
    layer1_outputs(4923) <= a;
    layer1_outputs(4924) <= a;
    layer1_outputs(4925) <= a or b;
    layer1_outputs(4926) <= not b or a;
    layer1_outputs(4927) <= b and not a;
    layer1_outputs(4928) <= not (a or b);
    layer1_outputs(4929) <= not (a and b);
    layer1_outputs(4930) <= b;
    layer1_outputs(4931) <= a;
    layer1_outputs(4932) <= not b or a;
    layer1_outputs(4933) <= not (a xor b);
    layer1_outputs(4934) <= not a;
    layer1_outputs(4935) <= not (a and b);
    layer1_outputs(4936) <= a and not b;
    layer1_outputs(4937) <= not (a xor b);
    layer1_outputs(4938) <= a and not b;
    layer1_outputs(4939) <= not b or a;
    layer1_outputs(4940) <= a;
    layer1_outputs(4941) <= not a or b;
    layer1_outputs(4942) <= not b;
    layer1_outputs(4943) <= not (a xor b);
    layer1_outputs(4944) <= a and not b;
    layer1_outputs(4945) <= a and b;
    layer1_outputs(4946) <= not b;
    layer1_outputs(4947) <= a or b;
    layer1_outputs(4948) <= a and b;
    layer1_outputs(4949) <= not a or b;
    layer1_outputs(4950) <= not b;
    layer1_outputs(4951) <= not b;
    layer1_outputs(4952) <= b and not a;
    layer1_outputs(4953) <= 1'b1;
    layer1_outputs(4954) <= not (a or b);
    layer1_outputs(4955) <= not b;
    layer1_outputs(4956) <= not (a and b);
    layer1_outputs(4957) <= b;
    layer1_outputs(4958) <= a xor b;
    layer1_outputs(4959) <= not a or b;
    layer1_outputs(4960) <= b;
    layer1_outputs(4961) <= 1'b1;
    layer1_outputs(4962) <= not (a or b);
    layer1_outputs(4963) <= a;
    layer1_outputs(4964) <= not (a xor b);
    layer1_outputs(4965) <= not (a and b);
    layer1_outputs(4966) <= a xor b;
    layer1_outputs(4967) <= not (a and b);
    layer1_outputs(4968) <= not b;
    layer1_outputs(4969) <= not a;
    layer1_outputs(4970) <= not (a or b);
    layer1_outputs(4971) <= not a;
    layer1_outputs(4972) <= not b;
    layer1_outputs(4973) <= b;
    layer1_outputs(4974) <= not b or a;
    layer1_outputs(4975) <= 1'b0;
    layer1_outputs(4976) <= b;
    layer1_outputs(4977) <= a xor b;
    layer1_outputs(4978) <= not (a or b);
    layer1_outputs(4979) <= a xor b;
    layer1_outputs(4980) <= not a;
    layer1_outputs(4981) <= a or b;
    layer1_outputs(4982) <= not (a and b);
    layer1_outputs(4983) <= not b or a;
    layer1_outputs(4984) <= b and not a;
    layer1_outputs(4985) <= not b;
    layer1_outputs(4986) <= a;
    layer1_outputs(4987) <= not a;
    layer1_outputs(4988) <= a and not b;
    layer1_outputs(4989) <= not a;
    layer1_outputs(4990) <= a and not b;
    layer1_outputs(4991) <= not (a or b);
    layer1_outputs(4992) <= not b or a;
    layer1_outputs(4993) <= a and b;
    layer1_outputs(4994) <= not b or a;
    layer1_outputs(4995) <= not b;
    layer1_outputs(4996) <= a or b;
    layer1_outputs(4997) <= a and b;
    layer1_outputs(4998) <= b and not a;
    layer1_outputs(4999) <= a;
    layer1_outputs(5000) <= not a;
    layer1_outputs(5001) <= not a or b;
    layer1_outputs(5002) <= b and not a;
    layer1_outputs(5003) <= not a or b;
    layer1_outputs(5004) <= a and b;
    layer1_outputs(5005) <= a;
    layer1_outputs(5006) <= not b;
    layer1_outputs(5007) <= not a or b;
    layer1_outputs(5008) <= not (a xor b);
    layer1_outputs(5009) <= not (a and b);
    layer1_outputs(5010) <= not (a and b);
    layer1_outputs(5011) <= b;
    layer1_outputs(5012) <= a;
    layer1_outputs(5013) <= not (a xor b);
    layer1_outputs(5014) <= a or b;
    layer1_outputs(5015) <= not a;
    layer1_outputs(5016) <= b;
    layer1_outputs(5017) <= b and not a;
    layer1_outputs(5018) <= b;
    layer1_outputs(5019) <= not (a or b);
    layer1_outputs(5020) <= not a or b;
    layer1_outputs(5021) <= a xor b;
    layer1_outputs(5022) <= b;
    layer1_outputs(5023) <= not (a or b);
    layer1_outputs(5024) <= not (a or b);
    layer1_outputs(5025) <= a;
    layer1_outputs(5026) <= not b;
    layer1_outputs(5027) <= b and not a;
    layer1_outputs(5028) <= not (a and b);
    layer1_outputs(5029) <= not a or b;
    layer1_outputs(5030) <= a xor b;
    layer1_outputs(5031) <= a or b;
    layer1_outputs(5032) <= a or b;
    layer1_outputs(5033) <= a xor b;
    layer1_outputs(5034) <= not (a and b);
    layer1_outputs(5035) <= not (a xor b);
    layer1_outputs(5036) <= not (a or b);
    layer1_outputs(5037) <= b;
    layer1_outputs(5038) <= a and not b;
    layer1_outputs(5039) <= not b;
    layer1_outputs(5040) <= a and b;
    layer1_outputs(5041) <= not (a and b);
    layer1_outputs(5042) <= a and b;
    layer1_outputs(5043) <= not b;
    layer1_outputs(5044) <= not b or a;
    layer1_outputs(5045) <= b and not a;
    layer1_outputs(5046) <= a;
    layer1_outputs(5047) <= not b or a;
    layer1_outputs(5048) <= not a or b;
    layer1_outputs(5049) <= a and b;
    layer1_outputs(5050) <= not (a or b);
    layer1_outputs(5051) <= a xor b;
    layer1_outputs(5052) <= not b;
    layer1_outputs(5053) <= not (a or b);
    layer1_outputs(5054) <= b;
    layer1_outputs(5055) <= not (a or b);
    layer1_outputs(5056) <= a xor b;
    layer1_outputs(5057) <= not b or a;
    layer1_outputs(5058) <= b and not a;
    layer1_outputs(5059) <= a;
    layer1_outputs(5060) <= a;
    layer1_outputs(5061) <= b;
    layer1_outputs(5062) <= not b or a;
    layer1_outputs(5063) <= a or b;
    layer1_outputs(5064) <= not (a xor b);
    layer1_outputs(5065) <= not b or a;
    layer1_outputs(5066) <= b and not a;
    layer1_outputs(5067) <= not b;
    layer1_outputs(5068) <= a;
    layer1_outputs(5069) <= a and not b;
    layer1_outputs(5070) <= a and not b;
    layer1_outputs(5071) <= a or b;
    layer1_outputs(5072) <= not (a xor b);
    layer1_outputs(5073) <= b;
    layer1_outputs(5074) <= a or b;
    layer1_outputs(5075) <= b;
    layer1_outputs(5076) <= a and not b;
    layer1_outputs(5077) <= not b or a;
    layer1_outputs(5078) <= not b;
    layer1_outputs(5079) <= a;
    layer1_outputs(5080) <= a;
    layer1_outputs(5081) <= a xor b;
    layer1_outputs(5082) <= not (a or b);
    layer1_outputs(5083) <= a and b;
    layer1_outputs(5084) <= not b or a;
    layer1_outputs(5085) <= b and not a;
    layer1_outputs(5086) <= not a;
    layer1_outputs(5087) <= a or b;
    layer1_outputs(5088) <= a;
    layer1_outputs(5089) <= b and not a;
    layer1_outputs(5090) <= a and not b;
    layer1_outputs(5091) <= not b or a;
    layer1_outputs(5092) <= not a;
    layer1_outputs(5093) <= not (a and b);
    layer1_outputs(5094) <= b;
    layer1_outputs(5095) <= not (a xor b);
    layer1_outputs(5096) <= b and not a;
    layer1_outputs(5097) <= a;
    layer1_outputs(5098) <= not b;
    layer1_outputs(5099) <= a or b;
    layer1_outputs(5100) <= a xor b;
    layer1_outputs(5101) <= not a;
    layer1_outputs(5102) <= not b;
    layer1_outputs(5103) <= not (a or b);
    layer1_outputs(5104) <= a and not b;
    layer1_outputs(5105) <= a;
    layer1_outputs(5106) <= not (a or b);
    layer1_outputs(5107) <= not a or b;
    layer1_outputs(5108) <= a and not b;
    layer1_outputs(5109) <= a and b;
    layer1_outputs(5110) <= a and b;
    layer1_outputs(5111) <= a xor b;
    layer1_outputs(5112) <= not a or b;
    layer1_outputs(5113) <= not (a or b);
    layer1_outputs(5114) <= b;
    layer1_outputs(5115) <= not a;
    layer1_outputs(5116) <= not b or a;
    layer1_outputs(5117) <= b and not a;
    layer1_outputs(5118) <= not b;
    layer1_outputs(5119) <= 1'b1;
    layer1_outputs(5120) <= not a or b;
    layer1_outputs(5121) <= b and not a;
    layer1_outputs(5122) <= not (a xor b);
    layer1_outputs(5123) <= a and b;
    layer1_outputs(5124) <= a;
    layer1_outputs(5125) <= b and not a;
    layer1_outputs(5126) <= a or b;
    layer1_outputs(5127) <= b and not a;
    layer1_outputs(5128) <= a xor b;
    layer1_outputs(5129) <= not a or b;
    layer1_outputs(5130) <= b;
    layer1_outputs(5131) <= not b;
    layer1_outputs(5132) <= a xor b;
    layer1_outputs(5133) <= not a;
    layer1_outputs(5134) <= not a or b;
    layer1_outputs(5135) <= not (a and b);
    layer1_outputs(5136) <= a;
    layer1_outputs(5137) <= not (a and b);
    layer1_outputs(5138) <= b;
    layer1_outputs(5139) <= b;
    layer1_outputs(5140) <= a xor b;
    layer1_outputs(5141) <= not b or a;
    layer1_outputs(5142) <= not b;
    layer1_outputs(5143) <= a and b;
    layer1_outputs(5144) <= a;
    layer1_outputs(5145) <= not a or b;
    layer1_outputs(5146) <= a;
    layer1_outputs(5147) <= a and b;
    layer1_outputs(5148) <= b;
    layer1_outputs(5149) <= a;
    layer1_outputs(5150) <= not (a and b);
    layer1_outputs(5151) <= not a;
    layer1_outputs(5152) <= not a;
    layer1_outputs(5153) <= a and not b;
    layer1_outputs(5154) <= not a or b;
    layer1_outputs(5155) <= not (a xor b);
    layer1_outputs(5156) <= a;
    layer1_outputs(5157) <= not (a and b);
    layer1_outputs(5158) <= not b;
    layer1_outputs(5159) <= not a;
    layer1_outputs(5160) <= not b or a;
    layer1_outputs(5161) <= not (a xor b);
    layer1_outputs(5162) <= a;
    layer1_outputs(5163) <= not a;
    layer1_outputs(5164) <= b and not a;
    layer1_outputs(5165) <= b and not a;
    layer1_outputs(5166) <= a or b;
    layer1_outputs(5167) <= b and not a;
    layer1_outputs(5168) <= not b or a;
    layer1_outputs(5169) <= a;
    layer1_outputs(5170) <= not b or a;
    layer1_outputs(5171) <= 1'b1;
    layer1_outputs(5172) <= not b or a;
    layer1_outputs(5173) <= not b;
    layer1_outputs(5174) <= a and not b;
    layer1_outputs(5175) <= 1'b1;
    layer1_outputs(5176) <= not (a and b);
    layer1_outputs(5177) <= a xor b;
    layer1_outputs(5178) <= not b or a;
    layer1_outputs(5179) <= not (a or b);
    layer1_outputs(5180) <= a;
    layer1_outputs(5181) <= a xor b;
    layer1_outputs(5182) <= a and b;
    layer1_outputs(5183) <= b;
    layer1_outputs(5184) <= b;
    layer1_outputs(5185) <= b and not a;
    layer1_outputs(5186) <= b;
    layer1_outputs(5187) <= not b or a;
    layer1_outputs(5188) <= not a;
    layer1_outputs(5189) <= not (a or b);
    layer1_outputs(5190) <= not b or a;
    layer1_outputs(5191) <= not b;
    layer1_outputs(5192) <= not (a xor b);
    layer1_outputs(5193) <= b and not a;
    layer1_outputs(5194) <= not a;
    layer1_outputs(5195) <= b;
    layer1_outputs(5196) <= not b;
    layer1_outputs(5197) <= not b;
    layer1_outputs(5198) <= b;
    layer1_outputs(5199) <= 1'b1;
    layer1_outputs(5200) <= b;
    layer1_outputs(5201) <= a and b;
    layer1_outputs(5202) <= not (a or b);
    layer1_outputs(5203) <= not (a xor b);
    layer1_outputs(5204) <= a;
    layer1_outputs(5205) <= a and b;
    layer1_outputs(5206) <= not (a xor b);
    layer1_outputs(5207) <= not b or a;
    layer1_outputs(5208) <= not b;
    layer1_outputs(5209) <= not (a and b);
    layer1_outputs(5210) <= a or b;
    layer1_outputs(5211) <= not a or b;
    layer1_outputs(5212) <= a;
    layer1_outputs(5213) <= not (a and b);
    layer1_outputs(5214) <= not (a xor b);
    layer1_outputs(5215) <= not a;
    layer1_outputs(5216) <= 1'b1;
    layer1_outputs(5217) <= not (a xor b);
    layer1_outputs(5218) <= a;
    layer1_outputs(5219) <= a;
    layer1_outputs(5220) <= not b;
    layer1_outputs(5221) <= not a;
    layer1_outputs(5222) <= a and not b;
    layer1_outputs(5223) <= not (a and b);
    layer1_outputs(5224) <= not (a or b);
    layer1_outputs(5225) <= a;
    layer1_outputs(5226) <= a or b;
    layer1_outputs(5227) <= a xor b;
    layer1_outputs(5228) <= not (a and b);
    layer1_outputs(5229) <= b;
    layer1_outputs(5230) <= not (a xor b);
    layer1_outputs(5231) <= not b;
    layer1_outputs(5232) <= not a or b;
    layer1_outputs(5233) <= not b;
    layer1_outputs(5234) <= not b or a;
    layer1_outputs(5235) <= a;
    layer1_outputs(5236) <= not (a xor b);
    layer1_outputs(5237) <= a;
    layer1_outputs(5238) <= a;
    layer1_outputs(5239) <= a and b;
    layer1_outputs(5240) <= not a;
    layer1_outputs(5241) <= b and not a;
    layer1_outputs(5242) <= a and b;
    layer1_outputs(5243) <= b;
    layer1_outputs(5244) <= b;
    layer1_outputs(5245) <= a and not b;
    layer1_outputs(5246) <= b and not a;
    layer1_outputs(5247) <= not a or b;
    layer1_outputs(5248) <= a xor b;
    layer1_outputs(5249) <= not a;
    layer1_outputs(5250) <= b;
    layer1_outputs(5251) <= a and b;
    layer1_outputs(5252) <= a and b;
    layer1_outputs(5253) <= b and not a;
    layer1_outputs(5254) <= not (a or b);
    layer1_outputs(5255) <= a xor b;
    layer1_outputs(5256) <= a xor b;
    layer1_outputs(5257) <= not (a xor b);
    layer1_outputs(5258) <= not (a xor b);
    layer1_outputs(5259) <= not a or b;
    layer1_outputs(5260) <= not (a xor b);
    layer1_outputs(5261) <= a or b;
    layer1_outputs(5262) <= not a or b;
    layer1_outputs(5263) <= not b or a;
    layer1_outputs(5264) <= a xor b;
    layer1_outputs(5265) <= not a;
    layer1_outputs(5266) <= not (a or b);
    layer1_outputs(5267) <= b and not a;
    layer1_outputs(5268) <= not b or a;
    layer1_outputs(5269) <= not (a or b);
    layer1_outputs(5270) <= not b or a;
    layer1_outputs(5271) <= a xor b;
    layer1_outputs(5272) <= not a;
    layer1_outputs(5273) <= not b or a;
    layer1_outputs(5274) <= b;
    layer1_outputs(5275) <= not (a and b);
    layer1_outputs(5276) <= b;
    layer1_outputs(5277) <= not a;
    layer1_outputs(5278) <= b and not a;
    layer1_outputs(5279) <= a or b;
    layer1_outputs(5280) <= not a or b;
    layer1_outputs(5281) <= not a or b;
    layer1_outputs(5282) <= not b;
    layer1_outputs(5283) <= a or b;
    layer1_outputs(5284) <= b;
    layer1_outputs(5285) <= a;
    layer1_outputs(5286) <= a or b;
    layer1_outputs(5287) <= a or b;
    layer1_outputs(5288) <= not (a and b);
    layer1_outputs(5289) <= not (a and b);
    layer1_outputs(5290) <= b and not a;
    layer1_outputs(5291) <= not b;
    layer1_outputs(5292) <= a xor b;
    layer1_outputs(5293) <= a xor b;
    layer1_outputs(5294) <= not b or a;
    layer1_outputs(5295) <= b;
    layer1_outputs(5296) <= b and not a;
    layer1_outputs(5297) <= a xor b;
    layer1_outputs(5298) <= b;
    layer1_outputs(5299) <= a;
    layer1_outputs(5300) <= a xor b;
    layer1_outputs(5301) <= not (a and b);
    layer1_outputs(5302) <= a;
    layer1_outputs(5303) <= not b or a;
    layer1_outputs(5304) <= not b or a;
    layer1_outputs(5305) <= not b or a;
    layer1_outputs(5306) <= not (a or b);
    layer1_outputs(5307) <= a and not b;
    layer1_outputs(5308) <= b and not a;
    layer1_outputs(5309) <= not b;
    layer1_outputs(5310) <= not a;
    layer1_outputs(5311) <= b;
    layer1_outputs(5312) <= b and not a;
    layer1_outputs(5313) <= b and not a;
    layer1_outputs(5314) <= b;
    layer1_outputs(5315) <= not (a or b);
    layer1_outputs(5316) <= a xor b;
    layer1_outputs(5317) <= b;
    layer1_outputs(5318) <= not (a or b);
    layer1_outputs(5319) <= a and b;
    layer1_outputs(5320) <= not b;
    layer1_outputs(5321) <= not b or a;
    layer1_outputs(5322) <= b and not a;
    layer1_outputs(5323) <= not a or b;
    layer1_outputs(5324) <= a;
    layer1_outputs(5325) <= a or b;
    layer1_outputs(5326) <= not (a xor b);
    layer1_outputs(5327) <= a xor b;
    layer1_outputs(5328) <= not (a and b);
    layer1_outputs(5329) <= not b;
    layer1_outputs(5330) <= not (a or b);
    layer1_outputs(5331) <= not b or a;
    layer1_outputs(5332) <= not b;
    layer1_outputs(5333) <= a or b;
    layer1_outputs(5334) <= a and not b;
    layer1_outputs(5335) <= a and not b;
    layer1_outputs(5336) <= b and not a;
    layer1_outputs(5337) <= b;
    layer1_outputs(5338) <= not b;
    layer1_outputs(5339) <= a or b;
    layer1_outputs(5340) <= a xor b;
    layer1_outputs(5341) <= a and not b;
    layer1_outputs(5342) <= b and not a;
    layer1_outputs(5343) <= not (a and b);
    layer1_outputs(5344) <= a xor b;
    layer1_outputs(5345) <= b;
    layer1_outputs(5346) <= not (a or b);
    layer1_outputs(5347) <= b;
    layer1_outputs(5348) <= not (a xor b);
    layer1_outputs(5349) <= not a;
    layer1_outputs(5350) <= a;
    layer1_outputs(5351) <= not (a or b);
    layer1_outputs(5352) <= a and b;
    layer1_outputs(5353) <= a and not b;
    layer1_outputs(5354) <= b;
    layer1_outputs(5355) <= not (a or b);
    layer1_outputs(5356) <= not a;
    layer1_outputs(5357) <= not a;
    layer1_outputs(5358) <= 1'b1;
    layer1_outputs(5359) <= a and b;
    layer1_outputs(5360) <= not (a or b);
    layer1_outputs(5361) <= a or b;
    layer1_outputs(5362) <= a and not b;
    layer1_outputs(5363) <= not a;
    layer1_outputs(5364) <= not a;
    layer1_outputs(5365) <= not b;
    layer1_outputs(5366) <= a and b;
    layer1_outputs(5367) <= a and not b;
    layer1_outputs(5368) <= not b or a;
    layer1_outputs(5369) <= not b;
    layer1_outputs(5370) <= a and not b;
    layer1_outputs(5371) <= not b;
    layer1_outputs(5372) <= not (a and b);
    layer1_outputs(5373) <= a;
    layer1_outputs(5374) <= a xor b;
    layer1_outputs(5375) <= 1'b1;
    layer1_outputs(5376) <= a;
    layer1_outputs(5377) <= not a or b;
    layer1_outputs(5378) <= a xor b;
    layer1_outputs(5379) <= not (a and b);
    layer1_outputs(5380) <= not (a and b);
    layer1_outputs(5381) <= a xor b;
    layer1_outputs(5382) <= a;
    layer1_outputs(5383) <= not (a xor b);
    layer1_outputs(5384) <= a;
    layer1_outputs(5385) <= not b or a;
    layer1_outputs(5386) <= not a;
    layer1_outputs(5387) <= b and not a;
    layer1_outputs(5388) <= a;
    layer1_outputs(5389) <= not b;
    layer1_outputs(5390) <= a;
    layer1_outputs(5391) <= b and not a;
    layer1_outputs(5392) <= not a;
    layer1_outputs(5393) <= a;
    layer1_outputs(5394) <= b and not a;
    layer1_outputs(5395) <= 1'b1;
    layer1_outputs(5396) <= b and not a;
    layer1_outputs(5397) <= b;
    layer1_outputs(5398) <= not (a xor b);
    layer1_outputs(5399) <= not (a xor b);
    layer1_outputs(5400) <= not (a or b);
    layer1_outputs(5401) <= not a;
    layer1_outputs(5402) <= not a;
    layer1_outputs(5403) <= not (a or b);
    layer1_outputs(5404) <= a and not b;
    layer1_outputs(5405) <= not b;
    layer1_outputs(5406) <= not (a or b);
    layer1_outputs(5407) <= b and not a;
    layer1_outputs(5408) <= not a;
    layer1_outputs(5409) <= not b or a;
    layer1_outputs(5410) <= not (a and b);
    layer1_outputs(5411) <= b;
    layer1_outputs(5412) <= b;
    layer1_outputs(5413) <= a and b;
    layer1_outputs(5414) <= a or b;
    layer1_outputs(5415) <= a and b;
    layer1_outputs(5416) <= b and not a;
    layer1_outputs(5417) <= b and not a;
    layer1_outputs(5418) <= not b or a;
    layer1_outputs(5419) <= a xor b;
    layer1_outputs(5420) <= not b or a;
    layer1_outputs(5421) <= not b;
    layer1_outputs(5422) <= not (a xor b);
    layer1_outputs(5423) <= not (a or b);
    layer1_outputs(5424) <= not b;
    layer1_outputs(5425) <= not b;
    layer1_outputs(5426) <= a;
    layer1_outputs(5427) <= b and not a;
    layer1_outputs(5428) <= not a;
    layer1_outputs(5429) <= not (a xor b);
    layer1_outputs(5430) <= not b;
    layer1_outputs(5431) <= not b or a;
    layer1_outputs(5432) <= a and not b;
    layer1_outputs(5433) <= 1'b0;
    layer1_outputs(5434) <= 1'b1;
    layer1_outputs(5435) <= a;
    layer1_outputs(5436) <= not b;
    layer1_outputs(5437) <= a and not b;
    layer1_outputs(5438) <= not (a xor b);
    layer1_outputs(5439) <= a or b;
    layer1_outputs(5440) <= not a;
    layer1_outputs(5441) <= not b or a;
    layer1_outputs(5442) <= a xor b;
    layer1_outputs(5443) <= a;
    layer1_outputs(5444) <= not (a or b);
    layer1_outputs(5445) <= not b or a;
    layer1_outputs(5446) <= a xor b;
    layer1_outputs(5447) <= not (a and b);
    layer1_outputs(5448) <= not a;
    layer1_outputs(5449) <= a;
    layer1_outputs(5450) <= not b;
    layer1_outputs(5451) <= not b or a;
    layer1_outputs(5452) <= a xor b;
    layer1_outputs(5453) <= not (a xor b);
    layer1_outputs(5454) <= a and b;
    layer1_outputs(5455) <= a xor b;
    layer1_outputs(5456) <= not a or b;
    layer1_outputs(5457) <= not (a xor b);
    layer1_outputs(5458) <= 1'b0;
    layer1_outputs(5459) <= a;
    layer1_outputs(5460) <= not (a and b);
    layer1_outputs(5461) <= not a;
    layer1_outputs(5462) <= a;
    layer1_outputs(5463) <= not a or b;
    layer1_outputs(5464) <= a or b;
    layer1_outputs(5465) <= not a or b;
    layer1_outputs(5466) <= not (a and b);
    layer1_outputs(5467) <= not b or a;
    layer1_outputs(5468) <= not (a and b);
    layer1_outputs(5469) <= a and not b;
    layer1_outputs(5470) <= a xor b;
    layer1_outputs(5471) <= not a;
    layer1_outputs(5472) <= a or b;
    layer1_outputs(5473) <= not b;
    layer1_outputs(5474) <= not b;
    layer1_outputs(5475) <= a and b;
    layer1_outputs(5476) <= not (a or b);
    layer1_outputs(5477) <= a;
    layer1_outputs(5478) <= not (a or b);
    layer1_outputs(5479) <= a;
    layer1_outputs(5480) <= a and b;
    layer1_outputs(5481) <= a and not b;
    layer1_outputs(5482) <= 1'b1;
    layer1_outputs(5483) <= not (a xor b);
    layer1_outputs(5484) <= a and not b;
    layer1_outputs(5485) <= a and b;
    layer1_outputs(5486) <= not a;
    layer1_outputs(5487) <= not b or a;
    layer1_outputs(5488) <= not b or a;
    layer1_outputs(5489) <= not (a xor b);
    layer1_outputs(5490) <= a;
    layer1_outputs(5491) <= a;
    layer1_outputs(5492) <= b and not a;
    layer1_outputs(5493) <= not a;
    layer1_outputs(5494) <= a and not b;
    layer1_outputs(5495) <= a and not b;
    layer1_outputs(5496) <= b;
    layer1_outputs(5497) <= a;
    layer1_outputs(5498) <= a;
    layer1_outputs(5499) <= b;
    layer1_outputs(5500) <= a and b;
    layer1_outputs(5501) <= not a;
    layer1_outputs(5502) <= not (a and b);
    layer1_outputs(5503) <= not (a and b);
    layer1_outputs(5504) <= a;
    layer1_outputs(5505) <= a or b;
    layer1_outputs(5506) <= a or b;
    layer1_outputs(5507) <= not (a and b);
    layer1_outputs(5508) <= not b or a;
    layer1_outputs(5509) <= not (a xor b);
    layer1_outputs(5510) <= not a;
    layer1_outputs(5511) <= a and b;
    layer1_outputs(5512) <= not (a xor b);
    layer1_outputs(5513) <= b;
    layer1_outputs(5514) <= not b or a;
    layer1_outputs(5515) <= not (a and b);
    layer1_outputs(5516) <= a or b;
    layer1_outputs(5517) <= a and not b;
    layer1_outputs(5518) <= not b or a;
    layer1_outputs(5519) <= not a;
    layer1_outputs(5520) <= a or b;
    layer1_outputs(5521) <= not (a or b);
    layer1_outputs(5522) <= a xor b;
    layer1_outputs(5523) <= not b;
    layer1_outputs(5524) <= a;
    layer1_outputs(5525) <= not a or b;
    layer1_outputs(5526) <= not b;
    layer1_outputs(5527) <= 1'b1;
    layer1_outputs(5528) <= a and b;
    layer1_outputs(5529) <= a;
    layer1_outputs(5530) <= not a or b;
    layer1_outputs(5531) <= not b or a;
    layer1_outputs(5532) <= not b;
    layer1_outputs(5533) <= not (a or b);
    layer1_outputs(5534) <= not b;
    layer1_outputs(5535) <= not b or a;
    layer1_outputs(5536) <= a and not b;
    layer1_outputs(5537) <= not a;
    layer1_outputs(5538) <= not (a xor b);
    layer1_outputs(5539) <= not b;
    layer1_outputs(5540) <= b and not a;
    layer1_outputs(5541) <= a and not b;
    layer1_outputs(5542) <= not (a xor b);
    layer1_outputs(5543) <= not b;
    layer1_outputs(5544) <= 1'b0;
    layer1_outputs(5545) <= a xor b;
    layer1_outputs(5546) <= not a;
    layer1_outputs(5547) <= b;
    layer1_outputs(5548) <= not (a xor b);
    layer1_outputs(5549) <= not a or b;
    layer1_outputs(5550) <= a and b;
    layer1_outputs(5551) <= not (a or b);
    layer1_outputs(5552) <= b;
    layer1_outputs(5553) <= a and b;
    layer1_outputs(5554) <= not a;
    layer1_outputs(5555) <= a or b;
    layer1_outputs(5556) <= not (a and b);
    layer1_outputs(5557) <= a and b;
    layer1_outputs(5558) <= not a or b;
    layer1_outputs(5559) <= b;
    layer1_outputs(5560) <= not (a and b);
    layer1_outputs(5561) <= not (a xor b);
    layer1_outputs(5562) <= a and not b;
    layer1_outputs(5563) <= not b or a;
    layer1_outputs(5564) <= 1'b0;
    layer1_outputs(5565) <= not (a or b);
    layer1_outputs(5566) <= not a;
    layer1_outputs(5567) <= a xor b;
    layer1_outputs(5568) <= 1'b1;
    layer1_outputs(5569) <= b;
    layer1_outputs(5570) <= not (a xor b);
    layer1_outputs(5571) <= not a or b;
    layer1_outputs(5572) <= not a;
    layer1_outputs(5573) <= not a or b;
    layer1_outputs(5574) <= not (a xor b);
    layer1_outputs(5575) <= not a;
    layer1_outputs(5576) <= not a;
    layer1_outputs(5577) <= not a;
    layer1_outputs(5578) <= not b or a;
    layer1_outputs(5579) <= not (a and b);
    layer1_outputs(5580) <= not (a or b);
    layer1_outputs(5581) <= not b;
    layer1_outputs(5582) <= not (a and b);
    layer1_outputs(5583) <= a or b;
    layer1_outputs(5584) <= not (a or b);
    layer1_outputs(5585) <= not a;
    layer1_outputs(5586) <= a or b;
    layer1_outputs(5587) <= 1'b0;
    layer1_outputs(5588) <= a and not b;
    layer1_outputs(5589) <= a and b;
    layer1_outputs(5590) <= a and b;
    layer1_outputs(5591) <= not b or a;
    layer1_outputs(5592) <= a xor b;
    layer1_outputs(5593) <= not a;
    layer1_outputs(5594) <= b and not a;
    layer1_outputs(5595) <= a and not b;
    layer1_outputs(5596) <= not a;
    layer1_outputs(5597) <= not b;
    layer1_outputs(5598) <= not (a and b);
    layer1_outputs(5599) <= a;
    layer1_outputs(5600) <= b and not a;
    layer1_outputs(5601) <= a xor b;
    layer1_outputs(5602) <= a xor b;
    layer1_outputs(5603) <= not a;
    layer1_outputs(5604) <= b;
    layer1_outputs(5605) <= a or b;
    layer1_outputs(5606) <= not a;
    layer1_outputs(5607) <= not b;
    layer1_outputs(5608) <= not b or a;
    layer1_outputs(5609) <= a xor b;
    layer1_outputs(5610) <= not b or a;
    layer1_outputs(5611) <= a and b;
    layer1_outputs(5612) <= a xor b;
    layer1_outputs(5613) <= a and not b;
    layer1_outputs(5614) <= not (a and b);
    layer1_outputs(5615) <= not b;
    layer1_outputs(5616) <= a;
    layer1_outputs(5617) <= not (a xor b);
    layer1_outputs(5618) <= a xor b;
    layer1_outputs(5619) <= not b;
    layer1_outputs(5620) <= not b;
    layer1_outputs(5621) <= a and b;
    layer1_outputs(5622) <= not b;
    layer1_outputs(5623) <= not (a or b);
    layer1_outputs(5624) <= a;
    layer1_outputs(5625) <= b;
    layer1_outputs(5626) <= b;
    layer1_outputs(5627) <= a xor b;
    layer1_outputs(5628) <= a or b;
    layer1_outputs(5629) <= a xor b;
    layer1_outputs(5630) <= not a;
    layer1_outputs(5631) <= not b;
    layer1_outputs(5632) <= not a;
    layer1_outputs(5633) <= a or b;
    layer1_outputs(5634) <= not (a and b);
    layer1_outputs(5635) <= a and b;
    layer1_outputs(5636) <= not b;
    layer1_outputs(5637) <= not a or b;
    layer1_outputs(5638) <= not (a or b);
    layer1_outputs(5639) <= not (a or b);
    layer1_outputs(5640) <= not a or b;
    layer1_outputs(5641) <= not a;
    layer1_outputs(5642) <= a;
    layer1_outputs(5643) <= a and not b;
    layer1_outputs(5644) <= not b or a;
    layer1_outputs(5645) <= not a;
    layer1_outputs(5646) <= a;
    layer1_outputs(5647) <= a xor b;
    layer1_outputs(5648) <= a and b;
    layer1_outputs(5649) <= a xor b;
    layer1_outputs(5650) <= not (a or b);
    layer1_outputs(5651) <= b and not a;
    layer1_outputs(5652) <= not a or b;
    layer1_outputs(5653) <= not (a and b);
    layer1_outputs(5654) <= a xor b;
    layer1_outputs(5655) <= not (a and b);
    layer1_outputs(5656) <= b and not a;
    layer1_outputs(5657) <= b;
    layer1_outputs(5658) <= not a or b;
    layer1_outputs(5659) <= b;
    layer1_outputs(5660) <= a;
    layer1_outputs(5661) <= not (a or b);
    layer1_outputs(5662) <= a and not b;
    layer1_outputs(5663) <= not a;
    layer1_outputs(5664) <= a;
    layer1_outputs(5665) <= not (a xor b);
    layer1_outputs(5666) <= a or b;
    layer1_outputs(5667) <= b and not a;
    layer1_outputs(5668) <= a and b;
    layer1_outputs(5669) <= not (a or b);
    layer1_outputs(5670) <= b and not a;
    layer1_outputs(5671) <= a or b;
    layer1_outputs(5672) <= a or b;
    layer1_outputs(5673) <= not a;
    layer1_outputs(5674) <= not (a and b);
    layer1_outputs(5675) <= 1'b1;
    layer1_outputs(5676) <= not b;
    layer1_outputs(5677) <= a xor b;
    layer1_outputs(5678) <= not b or a;
    layer1_outputs(5679) <= a and b;
    layer1_outputs(5680) <= not b or a;
    layer1_outputs(5681) <= a and not b;
    layer1_outputs(5682) <= not a;
    layer1_outputs(5683) <= a and not b;
    layer1_outputs(5684) <= not (a xor b);
    layer1_outputs(5685) <= not (a or b);
    layer1_outputs(5686) <= not a or b;
    layer1_outputs(5687) <= not b;
    layer1_outputs(5688) <= not a;
    layer1_outputs(5689) <= a xor b;
    layer1_outputs(5690) <= not b;
    layer1_outputs(5691) <= b and not a;
    layer1_outputs(5692) <= not a;
    layer1_outputs(5693) <= a and b;
    layer1_outputs(5694) <= not a;
    layer1_outputs(5695) <= b and not a;
    layer1_outputs(5696) <= a and b;
    layer1_outputs(5697) <= not (a xor b);
    layer1_outputs(5698) <= a and not b;
    layer1_outputs(5699) <= b;
    layer1_outputs(5700) <= not b;
    layer1_outputs(5701) <= not b or a;
    layer1_outputs(5702) <= b and not a;
    layer1_outputs(5703) <= not a;
    layer1_outputs(5704) <= a;
    layer1_outputs(5705) <= b;
    layer1_outputs(5706) <= 1'b0;
    layer1_outputs(5707) <= a xor b;
    layer1_outputs(5708) <= b and not a;
    layer1_outputs(5709) <= not (a or b);
    layer1_outputs(5710) <= not (a xor b);
    layer1_outputs(5711) <= not b;
    layer1_outputs(5712) <= not a or b;
    layer1_outputs(5713) <= a;
    layer1_outputs(5714) <= not a;
    layer1_outputs(5715) <= b;
    layer1_outputs(5716) <= not b;
    layer1_outputs(5717) <= a;
    layer1_outputs(5718) <= not a;
    layer1_outputs(5719) <= a and b;
    layer1_outputs(5720) <= not b;
    layer1_outputs(5721) <= a;
    layer1_outputs(5722) <= a;
    layer1_outputs(5723) <= a and not b;
    layer1_outputs(5724) <= a xor b;
    layer1_outputs(5725) <= not b;
    layer1_outputs(5726) <= a and not b;
    layer1_outputs(5727) <= not (a or b);
    layer1_outputs(5728) <= not (a and b);
    layer1_outputs(5729) <= a or b;
    layer1_outputs(5730) <= not (a or b);
    layer1_outputs(5731) <= not a or b;
    layer1_outputs(5732) <= not a;
    layer1_outputs(5733) <= not b;
    layer1_outputs(5734) <= a and not b;
    layer1_outputs(5735) <= a and b;
    layer1_outputs(5736) <= not b;
    layer1_outputs(5737) <= 1'b0;
    layer1_outputs(5738) <= a xor b;
    layer1_outputs(5739) <= not (a xor b);
    layer1_outputs(5740) <= b;
    layer1_outputs(5741) <= not a or b;
    layer1_outputs(5742) <= a and not b;
    layer1_outputs(5743) <= a;
    layer1_outputs(5744) <= b;
    layer1_outputs(5745) <= a and b;
    layer1_outputs(5746) <= a or b;
    layer1_outputs(5747) <= b and not a;
    layer1_outputs(5748) <= a;
    layer1_outputs(5749) <= not a or b;
    layer1_outputs(5750) <= not a or b;
    layer1_outputs(5751) <= not b;
    layer1_outputs(5752) <= not b;
    layer1_outputs(5753) <= not a;
    layer1_outputs(5754) <= a;
    layer1_outputs(5755) <= not (a xor b);
    layer1_outputs(5756) <= a and not b;
    layer1_outputs(5757) <= a or b;
    layer1_outputs(5758) <= a and not b;
    layer1_outputs(5759) <= a or b;
    layer1_outputs(5760) <= not (a and b);
    layer1_outputs(5761) <= a;
    layer1_outputs(5762) <= not a;
    layer1_outputs(5763) <= a;
    layer1_outputs(5764) <= not b;
    layer1_outputs(5765) <= a;
    layer1_outputs(5766) <= a;
    layer1_outputs(5767) <= not b;
    layer1_outputs(5768) <= not b;
    layer1_outputs(5769) <= b;
    layer1_outputs(5770) <= not a;
    layer1_outputs(5771) <= a and b;
    layer1_outputs(5772) <= not (a and b);
    layer1_outputs(5773) <= 1'b0;
    layer1_outputs(5774) <= b and not a;
    layer1_outputs(5775) <= a and not b;
    layer1_outputs(5776) <= not (a xor b);
    layer1_outputs(5777) <= not (a xor b);
    layer1_outputs(5778) <= 1'b1;
    layer1_outputs(5779) <= a and b;
    layer1_outputs(5780) <= not b;
    layer1_outputs(5781) <= a and not b;
    layer1_outputs(5782) <= not b or a;
    layer1_outputs(5783) <= not (a and b);
    layer1_outputs(5784) <= a and not b;
    layer1_outputs(5785) <= not (a and b);
    layer1_outputs(5786) <= a;
    layer1_outputs(5787) <= not a or b;
    layer1_outputs(5788) <= not b;
    layer1_outputs(5789) <= not b;
    layer1_outputs(5790) <= a and not b;
    layer1_outputs(5791) <= not b or a;
    layer1_outputs(5792) <= a xor b;
    layer1_outputs(5793) <= b and not a;
    layer1_outputs(5794) <= not b;
    layer1_outputs(5795) <= b and not a;
    layer1_outputs(5796) <= 1'b1;
    layer1_outputs(5797) <= a;
    layer1_outputs(5798) <= not b;
    layer1_outputs(5799) <= not a;
    layer1_outputs(5800) <= not a;
    layer1_outputs(5801) <= b and not a;
    layer1_outputs(5802) <= a or b;
    layer1_outputs(5803) <= not (a xor b);
    layer1_outputs(5804) <= not b;
    layer1_outputs(5805) <= b and not a;
    layer1_outputs(5806) <= not (a or b);
    layer1_outputs(5807) <= 1'b1;
    layer1_outputs(5808) <= a xor b;
    layer1_outputs(5809) <= a and not b;
    layer1_outputs(5810) <= not (a xor b);
    layer1_outputs(5811) <= b;
    layer1_outputs(5812) <= not a;
    layer1_outputs(5813) <= a or b;
    layer1_outputs(5814) <= not (a xor b);
    layer1_outputs(5815) <= not a;
    layer1_outputs(5816) <= a or b;
    layer1_outputs(5817) <= not a or b;
    layer1_outputs(5818) <= not a;
    layer1_outputs(5819) <= b;
    layer1_outputs(5820) <= not (a and b);
    layer1_outputs(5821) <= not (a or b);
    layer1_outputs(5822) <= a;
    layer1_outputs(5823) <= not (a and b);
    layer1_outputs(5824) <= not (a xor b);
    layer1_outputs(5825) <= not (a or b);
    layer1_outputs(5826) <= a and not b;
    layer1_outputs(5827) <= b;
    layer1_outputs(5828) <= a;
    layer1_outputs(5829) <= not a or b;
    layer1_outputs(5830) <= not a or b;
    layer1_outputs(5831) <= not (a and b);
    layer1_outputs(5832) <= not a;
    layer1_outputs(5833) <= a or b;
    layer1_outputs(5834) <= a and not b;
    layer1_outputs(5835) <= b;
    layer1_outputs(5836) <= not a or b;
    layer1_outputs(5837) <= a xor b;
    layer1_outputs(5838) <= a xor b;
    layer1_outputs(5839) <= not b;
    layer1_outputs(5840) <= not a;
    layer1_outputs(5841) <= a xor b;
    layer1_outputs(5842) <= a and b;
    layer1_outputs(5843) <= not (a xor b);
    layer1_outputs(5844) <= not b;
    layer1_outputs(5845) <= a and not b;
    layer1_outputs(5846) <= a;
    layer1_outputs(5847) <= b;
    layer1_outputs(5848) <= a and b;
    layer1_outputs(5849) <= not (a xor b);
    layer1_outputs(5850) <= a and b;
    layer1_outputs(5851) <= not (a or b);
    layer1_outputs(5852) <= not b or a;
    layer1_outputs(5853) <= not b;
    layer1_outputs(5854) <= b;
    layer1_outputs(5855) <= a;
    layer1_outputs(5856) <= a or b;
    layer1_outputs(5857) <= a;
    layer1_outputs(5858) <= b;
    layer1_outputs(5859) <= b;
    layer1_outputs(5860) <= b;
    layer1_outputs(5861) <= not a or b;
    layer1_outputs(5862) <= a and b;
    layer1_outputs(5863) <= not a or b;
    layer1_outputs(5864) <= not (a xor b);
    layer1_outputs(5865) <= not a or b;
    layer1_outputs(5866) <= a or b;
    layer1_outputs(5867) <= not (a or b);
    layer1_outputs(5868) <= not (a xor b);
    layer1_outputs(5869) <= a or b;
    layer1_outputs(5870) <= not a;
    layer1_outputs(5871) <= a and b;
    layer1_outputs(5872) <= not (a xor b);
    layer1_outputs(5873) <= not b;
    layer1_outputs(5874) <= not (a or b);
    layer1_outputs(5875) <= a;
    layer1_outputs(5876) <= a;
    layer1_outputs(5877) <= not (a and b);
    layer1_outputs(5878) <= not a;
    layer1_outputs(5879) <= a and not b;
    layer1_outputs(5880) <= a;
    layer1_outputs(5881) <= not (a and b);
    layer1_outputs(5882) <= not (a xor b);
    layer1_outputs(5883) <= not a or b;
    layer1_outputs(5884) <= a xor b;
    layer1_outputs(5885) <= not (a or b);
    layer1_outputs(5886) <= a;
    layer1_outputs(5887) <= a xor b;
    layer1_outputs(5888) <= not (a xor b);
    layer1_outputs(5889) <= not (a xor b);
    layer1_outputs(5890) <= a xor b;
    layer1_outputs(5891) <= b;
    layer1_outputs(5892) <= not (a xor b);
    layer1_outputs(5893) <= a xor b;
    layer1_outputs(5894) <= not a;
    layer1_outputs(5895) <= a;
    layer1_outputs(5896) <= not b;
    layer1_outputs(5897) <= b;
    layer1_outputs(5898) <= a;
    layer1_outputs(5899) <= not b;
    layer1_outputs(5900) <= a and b;
    layer1_outputs(5901) <= not (a or b);
    layer1_outputs(5902) <= not a or b;
    layer1_outputs(5903) <= not b or a;
    layer1_outputs(5904) <= b and not a;
    layer1_outputs(5905) <= not a;
    layer1_outputs(5906) <= b and not a;
    layer1_outputs(5907) <= b and not a;
    layer1_outputs(5908) <= b and not a;
    layer1_outputs(5909) <= a and not b;
    layer1_outputs(5910) <= b and not a;
    layer1_outputs(5911) <= not (a and b);
    layer1_outputs(5912) <= b and not a;
    layer1_outputs(5913) <= not a or b;
    layer1_outputs(5914) <= a and not b;
    layer1_outputs(5915) <= b;
    layer1_outputs(5916) <= a;
    layer1_outputs(5917) <= b;
    layer1_outputs(5918) <= a and not b;
    layer1_outputs(5919) <= a;
    layer1_outputs(5920) <= a and not b;
    layer1_outputs(5921) <= b;
    layer1_outputs(5922) <= b;
    layer1_outputs(5923) <= a and b;
    layer1_outputs(5924) <= not a;
    layer1_outputs(5925) <= b;
    layer1_outputs(5926) <= not b;
    layer1_outputs(5927) <= not b or a;
    layer1_outputs(5928) <= a and b;
    layer1_outputs(5929) <= not (a xor b);
    layer1_outputs(5930) <= not b or a;
    layer1_outputs(5931) <= not b;
    layer1_outputs(5932) <= a and not b;
    layer1_outputs(5933) <= not (a or b);
    layer1_outputs(5934) <= a or b;
    layer1_outputs(5935) <= not b;
    layer1_outputs(5936) <= a xor b;
    layer1_outputs(5937) <= a or b;
    layer1_outputs(5938) <= a or b;
    layer1_outputs(5939) <= not (a and b);
    layer1_outputs(5940) <= a or b;
    layer1_outputs(5941) <= not (a xor b);
    layer1_outputs(5942) <= b;
    layer1_outputs(5943) <= not a or b;
    layer1_outputs(5944) <= b and not a;
    layer1_outputs(5945) <= not (a xor b);
    layer1_outputs(5946) <= not b;
    layer1_outputs(5947) <= a and b;
    layer1_outputs(5948) <= a or b;
    layer1_outputs(5949) <= b and not a;
    layer1_outputs(5950) <= b and not a;
    layer1_outputs(5951) <= not a;
    layer1_outputs(5952) <= not b;
    layer1_outputs(5953) <= 1'b0;
    layer1_outputs(5954) <= not (a or b);
    layer1_outputs(5955) <= not a or b;
    layer1_outputs(5956) <= not a or b;
    layer1_outputs(5957) <= not b;
    layer1_outputs(5958) <= not (a xor b);
    layer1_outputs(5959) <= a;
    layer1_outputs(5960) <= not (a or b);
    layer1_outputs(5961) <= a;
    layer1_outputs(5962) <= a;
    layer1_outputs(5963) <= not (a and b);
    layer1_outputs(5964) <= a and not b;
    layer1_outputs(5965) <= not (a and b);
    layer1_outputs(5966) <= a and not b;
    layer1_outputs(5967) <= a;
    layer1_outputs(5968) <= not (a or b);
    layer1_outputs(5969) <= not a;
    layer1_outputs(5970) <= not (a or b);
    layer1_outputs(5971) <= 1'b1;
    layer1_outputs(5972) <= not (a or b);
    layer1_outputs(5973) <= not b;
    layer1_outputs(5974) <= a and b;
    layer1_outputs(5975) <= a or b;
    layer1_outputs(5976) <= a or b;
    layer1_outputs(5977) <= b;
    layer1_outputs(5978) <= a xor b;
    layer1_outputs(5979) <= a and not b;
    layer1_outputs(5980) <= not a or b;
    layer1_outputs(5981) <= not (a and b);
    layer1_outputs(5982) <= not (a and b);
    layer1_outputs(5983) <= b and not a;
    layer1_outputs(5984) <= a and b;
    layer1_outputs(5985) <= not b or a;
    layer1_outputs(5986) <= not b;
    layer1_outputs(5987) <= a;
    layer1_outputs(5988) <= not a;
    layer1_outputs(5989) <= a and not b;
    layer1_outputs(5990) <= a or b;
    layer1_outputs(5991) <= b;
    layer1_outputs(5992) <= not a;
    layer1_outputs(5993) <= 1'b0;
    layer1_outputs(5994) <= not a;
    layer1_outputs(5995) <= 1'b1;
    layer1_outputs(5996) <= a and b;
    layer1_outputs(5997) <= a xor b;
    layer1_outputs(5998) <= a or b;
    layer1_outputs(5999) <= not (a and b);
    layer1_outputs(6000) <= not (a and b);
    layer1_outputs(6001) <= not b;
    layer1_outputs(6002) <= a and b;
    layer1_outputs(6003) <= not (a xor b);
    layer1_outputs(6004) <= b;
    layer1_outputs(6005) <= a and b;
    layer1_outputs(6006) <= not b;
    layer1_outputs(6007) <= not a;
    layer1_outputs(6008) <= a or b;
    layer1_outputs(6009) <= a and not b;
    layer1_outputs(6010) <= not a or b;
    layer1_outputs(6011) <= a and b;
    layer1_outputs(6012) <= not a or b;
    layer1_outputs(6013) <= b and not a;
    layer1_outputs(6014) <= not b or a;
    layer1_outputs(6015) <= a or b;
    layer1_outputs(6016) <= a and b;
    layer1_outputs(6017) <= not b;
    layer1_outputs(6018) <= not b;
    layer1_outputs(6019) <= b;
    layer1_outputs(6020) <= b;
    layer1_outputs(6021) <= b;
    layer1_outputs(6022) <= not b or a;
    layer1_outputs(6023) <= not b;
    layer1_outputs(6024) <= not a or b;
    layer1_outputs(6025) <= a and not b;
    layer1_outputs(6026) <= a and b;
    layer1_outputs(6027) <= a;
    layer1_outputs(6028) <= not (a and b);
    layer1_outputs(6029) <= a and b;
    layer1_outputs(6030) <= not a;
    layer1_outputs(6031) <= a and not b;
    layer1_outputs(6032) <= not a or b;
    layer1_outputs(6033) <= not a or b;
    layer1_outputs(6034) <= a and not b;
    layer1_outputs(6035) <= b;
    layer1_outputs(6036) <= a or b;
    layer1_outputs(6037) <= not (a or b);
    layer1_outputs(6038) <= not a or b;
    layer1_outputs(6039) <= b and not a;
    layer1_outputs(6040) <= not (a xor b);
    layer1_outputs(6041) <= a or b;
    layer1_outputs(6042) <= a;
    layer1_outputs(6043) <= not (a and b);
    layer1_outputs(6044) <= not b or a;
    layer1_outputs(6045) <= not (a or b);
    layer1_outputs(6046) <= b and not a;
    layer1_outputs(6047) <= not a or b;
    layer1_outputs(6048) <= a and b;
    layer1_outputs(6049) <= b and not a;
    layer1_outputs(6050) <= a or b;
    layer1_outputs(6051) <= not a;
    layer1_outputs(6052) <= a;
    layer1_outputs(6053) <= not (a or b);
    layer1_outputs(6054) <= not b;
    layer1_outputs(6055) <= b and not a;
    layer1_outputs(6056) <= not (a xor b);
    layer1_outputs(6057) <= not (a and b);
    layer1_outputs(6058) <= a xor b;
    layer1_outputs(6059) <= a and not b;
    layer1_outputs(6060) <= a and b;
    layer1_outputs(6061) <= not (a and b);
    layer1_outputs(6062) <= a xor b;
    layer1_outputs(6063) <= not a;
    layer1_outputs(6064) <= a and b;
    layer1_outputs(6065) <= 1'b1;
    layer1_outputs(6066) <= not b;
    layer1_outputs(6067) <= not b;
    layer1_outputs(6068) <= a and not b;
    layer1_outputs(6069) <= a and not b;
    layer1_outputs(6070) <= a;
    layer1_outputs(6071) <= a;
    layer1_outputs(6072) <= b and not a;
    layer1_outputs(6073) <= not b;
    layer1_outputs(6074) <= a and b;
    layer1_outputs(6075) <= b and not a;
    layer1_outputs(6076) <= not b;
    layer1_outputs(6077) <= not a;
    layer1_outputs(6078) <= b and not a;
    layer1_outputs(6079) <= a or b;
    layer1_outputs(6080) <= not (a and b);
    layer1_outputs(6081) <= a;
    layer1_outputs(6082) <= a and not b;
    layer1_outputs(6083) <= a xor b;
    layer1_outputs(6084) <= not b or a;
    layer1_outputs(6085) <= not b;
    layer1_outputs(6086) <= not a;
    layer1_outputs(6087) <= a or b;
    layer1_outputs(6088) <= a and b;
    layer1_outputs(6089) <= b and not a;
    layer1_outputs(6090) <= not b;
    layer1_outputs(6091) <= b;
    layer1_outputs(6092) <= not b;
    layer1_outputs(6093) <= not b;
    layer1_outputs(6094) <= 1'b0;
    layer1_outputs(6095) <= not b or a;
    layer1_outputs(6096) <= a xor b;
    layer1_outputs(6097) <= not b;
    layer1_outputs(6098) <= a xor b;
    layer1_outputs(6099) <= b and not a;
    layer1_outputs(6100) <= not b;
    layer1_outputs(6101) <= not (a or b);
    layer1_outputs(6102) <= a;
    layer1_outputs(6103) <= not a or b;
    layer1_outputs(6104) <= a;
    layer1_outputs(6105) <= not b or a;
    layer1_outputs(6106) <= a;
    layer1_outputs(6107) <= not (a or b);
    layer1_outputs(6108) <= a and b;
    layer1_outputs(6109) <= a or b;
    layer1_outputs(6110) <= a or b;
    layer1_outputs(6111) <= a and not b;
    layer1_outputs(6112) <= not (a or b);
    layer1_outputs(6113) <= not b or a;
    layer1_outputs(6114) <= not b;
    layer1_outputs(6115) <= not (a or b);
    layer1_outputs(6116) <= not (a and b);
    layer1_outputs(6117) <= 1'b0;
    layer1_outputs(6118) <= a and b;
    layer1_outputs(6119) <= not a;
    layer1_outputs(6120) <= a and b;
    layer1_outputs(6121) <= not (a and b);
    layer1_outputs(6122) <= not b or a;
    layer1_outputs(6123) <= not b or a;
    layer1_outputs(6124) <= a or b;
    layer1_outputs(6125) <= a and b;
    layer1_outputs(6126) <= a or b;
    layer1_outputs(6127) <= a;
    layer1_outputs(6128) <= a xor b;
    layer1_outputs(6129) <= a and b;
    layer1_outputs(6130) <= a xor b;
    layer1_outputs(6131) <= not a or b;
    layer1_outputs(6132) <= not (a xor b);
    layer1_outputs(6133) <= a;
    layer1_outputs(6134) <= a or b;
    layer1_outputs(6135) <= not b or a;
    layer1_outputs(6136) <= a;
    layer1_outputs(6137) <= a and not b;
    layer1_outputs(6138) <= not (a and b);
    layer1_outputs(6139) <= a and b;
    layer1_outputs(6140) <= b;
    layer1_outputs(6141) <= not (a and b);
    layer1_outputs(6142) <= not (a and b);
    layer1_outputs(6143) <= not (a xor b);
    layer1_outputs(6144) <= not b;
    layer1_outputs(6145) <= not b;
    layer1_outputs(6146) <= not a;
    layer1_outputs(6147) <= not b or a;
    layer1_outputs(6148) <= not a;
    layer1_outputs(6149) <= b;
    layer1_outputs(6150) <= not a or b;
    layer1_outputs(6151) <= a or b;
    layer1_outputs(6152) <= b;
    layer1_outputs(6153) <= not a or b;
    layer1_outputs(6154) <= not a;
    layer1_outputs(6155) <= not a;
    layer1_outputs(6156) <= not a;
    layer1_outputs(6157) <= a or b;
    layer1_outputs(6158) <= not b or a;
    layer1_outputs(6159) <= a and b;
    layer1_outputs(6160) <= b;
    layer1_outputs(6161) <= not b or a;
    layer1_outputs(6162) <= a xor b;
    layer1_outputs(6163) <= a;
    layer1_outputs(6164) <= 1'b1;
    layer1_outputs(6165) <= a or b;
    layer1_outputs(6166) <= not b;
    layer1_outputs(6167) <= not (a and b);
    layer1_outputs(6168) <= not (a and b);
    layer1_outputs(6169) <= b;
    layer1_outputs(6170) <= not (a xor b);
    layer1_outputs(6171) <= a xor b;
    layer1_outputs(6172) <= b;
    layer1_outputs(6173) <= b;
    layer1_outputs(6174) <= a;
    layer1_outputs(6175) <= a and b;
    layer1_outputs(6176) <= not a;
    layer1_outputs(6177) <= not (a or b);
    layer1_outputs(6178) <= a and b;
    layer1_outputs(6179) <= not (a or b);
    layer1_outputs(6180) <= not (a and b);
    layer1_outputs(6181) <= not (a or b);
    layer1_outputs(6182) <= b and not a;
    layer1_outputs(6183) <= a xor b;
    layer1_outputs(6184) <= not (a xor b);
    layer1_outputs(6185) <= a and not b;
    layer1_outputs(6186) <= not a or b;
    layer1_outputs(6187) <= not (a and b);
    layer1_outputs(6188) <= a and not b;
    layer1_outputs(6189) <= a and b;
    layer1_outputs(6190) <= not (a xor b);
    layer1_outputs(6191) <= a xor b;
    layer1_outputs(6192) <= a xor b;
    layer1_outputs(6193) <= a or b;
    layer1_outputs(6194) <= not b;
    layer1_outputs(6195) <= not b;
    layer1_outputs(6196) <= a;
    layer1_outputs(6197) <= a or b;
    layer1_outputs(6198) <= a or b;
    layer1_outputs(6199) <= 1'b0;
    layer1_outputs(6200) <= not b;
    layer1_outputs(6201) <= a and b;
    layer1_outputs(6202) <= a;
    layer1_outputs(6203) <= not (a or b);
    layer1_outputs(6204) <= a;
    layer1_outputs(6205) <= not (a xor b);
    layer1_outputs(6206) <= a and not b;
    layer1_outputs(6207) <= 1'b1;
    layer1_outputs(6208) <= b;
    layer1_outputs(6209) <= a;
    layer1_outputs(6210) <= not (a and b);
    layer1_outputs(6211) <= a or b;
    layer1_outputs(6212) <= not a or b;
    layer1_outputs(6213) <= not b or a;
    layer1_outputs(6214) <= b and not a;
    layer1_outputs(6215) <= a or b;
    layer1_outputs(6216) <= not a or b;
    layer1_outputs(6217) <= not b;
    layer1_outputs(6218) <= b and not a;
    layer1_outputs(6219) <= not a or b;
    layer1_outputs(6220) <= b;
    layer1_outputs(6221) <= a xor b;
    layer1_outputs(6222) <= a;
    layer1_outputs(6223) <= b;
    layer1_outputs(6224) <= b and not a;
    layer1_outputs(6225) <= not a or b;
    layer1_outputs(6226) <= a or b;
    layer1_outputs(6227) <= a;
    layer1_outputs(6228) <= b;
    layer1_outputs(6229) <= not a;
    layer1_outputs(6230) <= a xor b;
    layer1_outputs(6231) <= b;
    layer1_outputs(6232) <= a;
    layer1_outputs(6233) <= b and not a;
    layer1_outputs(6234) <= 1'b0;
    layer1_outputs(6235) <= not b or a;
    layer1_outputs(6236) <= b and not a;
    layer1_outputs(6237) <= a or b;
    layer1_outputs(6238) <= not a;
    layer1_outputs(6239) <= b and not a;
    layer1_outputs(6240) <= not b;
    layer1_outputs(6241) <= 1'b1;
    layer1_outputs(6242) <= not (a xor b);
    layer1_outputs(6243) <= not b or a;
    layer1_outputs(6244) <= not a;
    layer1_outputs(6245) <= b;
    layer1_outputs(6246) <= a and not b;
    layer1_outputs(6247) <= a xor b;
    layer1_outputs(6248) <= b;
    layer1_outputs(6249) <= a xor b;
    layer1_outputs(6250) <= b and not a;
    layer1_outputs(6251) <= not (a xor b);
    layer1_outputs(6252) <= not (a xor b);
    layer1_outputs(6253) <= not a;
    layer1_outputs(6254) <= a xor b;
    layer1_outputs(6255) <= a;
    layer1_outputs(6256) <= a and not b;
    layer1_outputs(6257) <= b and not a;
    layer1_outputs(6258) <= a or b;
    layer1_outputs(6259) <= not a or b;
    layer1_outputs(6260) <= not (a and b);
    layer1_outputs(6261) <= not (a and b);
    layer1_outputs(6262) <= a and not b;
    layer1_outputs(6263) <= not b;
    layer1_outputs(6264) <= not a;
    layer1_outputs(6265) <= not b or a;
    layer1_outputs(6266) <= a xor b;
    layer1_outputs(6267) <= a and b;
    layer1_outputs(6268) <= not (a and b);
    layer1_outputs(6269) <= a;
    layer1_outputs(6270) <= b and not a;
    layer1_outputs(6271) <= not b;
    layer1_outputs(6272) <= not (a or b);
    layer1_outputs(6273) <= not b;
    layer1_outputs(6274) <= not b;
    layer1_outputs(6275) <= 1'b0;
    layer1_outputs(6276) <= not b or a;
    layer1_outputs(6277) <= not (a xor b);
    layer1_outputs(6278) <= a and not b;
    layer1_outputs(6279) <= a and not b;
    layer1_outputs(6280) <= a and b;
    layer1_outputs(6281) <= a and b;
    layer1_outputs(6282) <= a and not b;
    layer1_outputs(6283) <= not b;
    layer1_outputs(6284) <= a;
    layer1_outputs(6285) <= not a or b;
    layer1_outputs(6286) <= not b;
    layer1_outputs(6287) <= a;
    layer1_outputs(6288) <= not a;
    layer1_outputs(6289) <= a xor b;
    layer1_outputs(6290) <= not (a or b);
    layer1_outputs(6291) <= not a;
    layer1_outputs(6292) <= not a or b;
    layer1_outputs(6293) <= a or b;
    layer1_outputs(6294) <= a;
    layer1_outputs(6295) <= not (a xor b);
    layer1_outputs(6296) <= a;
    layer1_outputs(6297) <= b and not a;
    layer1_outputs(6298) <= a and b;
    layer1_outputs(6299) <= a and b;
    layer1_outputs(6300) <= b;
    layer1_outputs(6301) <= not (a xor b);
    layer1_outputs(6302) <= b;
    layer1_outputs(6303) <= not b;
    layer1_outputs(6304) <= a;
    layer1_outputs(6305) <= not a or b;
    layer1_outputs(6306) <= a xor b;
    layer1_outputs(6307) <= a and b;
    layer1_outputs(6308) <= not (a and b);
    layer1_outputs(6309) <= not (a and b);
    layer1_outputs(6310) <= a and b;
    layer1_outputs(6311) <= a and not b;
    layer1_outputs(6312) <= b;
    layer1_outputs(6313) <= b;
    layer1_outputs(6314) <= not (a and b);
    layer1_outputs(6315) <= not b;
    layer1_outputs(6316) <= not b or a;
    layer1_outputs(6317) <= a and not b;
    layer1_outputs(6318) <= b;
    layer1_outputs(6319) <= a and b;
    layer1_outputs(6320) <= b and not a;
    layer1_outputs(6321) <= not b;
    layer1_outputs(6322) <= b;
    layer1_outputs(6323) <= a xor b;
    layer1_outputs(6324) <= b and not a;
    layer1_outputs(6325) <= not b or a;
    layer1_outputs(6326) <= not (a xor b);
    layer1_outputs(6327) <= a and not b;
    layer1_outputs(6328) <= a or b;
    layer1_outputs(6329) <= a xor b;
    layer1_outputs(6330) <= a and b;
    layer1_outputs(6331) <= not b;
    layer1_outputs(6332) <= a and not b;
    layer1_outputs(6333) <= not (a and b);
    layer1_outputs(6334) <= not a;
    layer1_outputs(6335) <= a xor b;
    layer1_outputs(6336) <= b and not a;
    layer1_outputs(6337) <= b and not a;
    layer1_outputs(6338) <= a and not b;
    layer1_outputs(6339) <= not b;
    layer1_outputs(6340) <= not a;
    layer1_outputs(6341) <= not a or b;
    layer1_outputs(6342) <= b and not a;
    layer1_outputs(6343) <= not b or a;
    layer1_outputs(6344) <= not a or b;
    layer1_outputs(6345) <= not b;
    layer1_outputs(6346) <= not (a or b);
    layer1_outputs(6347) <= not b or a;
    layer1_outputs(6348) <= not b;
    layer1_outputs(6349) <= not a or b;
    layer1_outputs(6350) <= not (a xor b);
    layer1_outputs(6351) <= a or b;
    layer1_outputs(6352) <= not (a or b);
    layer1_outputs(6353) <= not b or a;
    layer1_outputs(6354) <= b;
    layer1_outputs(6355) <= not b;
    layer1_outputs(6356) <= not (a xor b);
    layer1_outputs(6357) <= b;
    layer1_outputs(6358) <= not a;
    layer1_outputs(6359) <= not b;
    layer1_outputs(6360) <= not b or a;
    layer1_outputs(6361) <= not (a xor b);
    layer1_outputs(6362) <= a;
    layer1_outputs(6363) <= not (a and b);
    layer1_outputs(6364) <= not b or a;
    layer1_outputs(6365) <= a;
    layer1_outputs(6366) <= b;
    layer1_outputs(6367) <= not (a or b);
    layer1_outputs(6368) <= not b;
    layer1_outputs(6369) <= not (a or b);
    layer1_outputs(6370) <= not (a or b);
    layer1_outputs(6371) <= b;
    layer1_outputs(6372) <= a and b;
    layer1_outputs(6373) <= not b;
    layer1_outputs(6374) <= not (a and b);
    layer1_outputs(6375) <= not b;
    layer1_outputs(6376) <= not b;
    layer1_outputs(6377) <= a;
    layer1_outputs(6378) <= a and b;
    layer1_outputs(6379) <= not (a or b);
    layer1_outputs(6380) <= not b or a;
    layer1_outputs(6381) <= not a;
    layer1_outputs(6382) <= not a or b;
    layer1_outputs(6383) <= b and not a;
    layer1_outputs(6384) <= a and not b;
    layer1_outputs(6385) <= a;
    layer1_outputs(6386) <= b;
    layer1_outputs(6387) <= a xor b;
    layer1_outputs(6388) <= a and not b;
    layer1_outputs(6389) <= not b;
    layer1_outputs(6390) <= a and not b;
    layer1_outputs(6391) <= a;
    layer1_outputs(6392) <= not a;
    layer1_outputs(6393) <= a xor b;
    layer1_outputs(6394) <= not (a or b);
    layer1_outputs(6395) <= b;
    layer1_outputs(6396) <= b and not a;
    layer1_outputs(6397) <= 1'b0;
    layer1_outputs(6398) <= b;
    layer1_outputs(6399) <= not b;
    layer1_outputs(6400) <= not b or a;
    layer1_outputs(6401) <= not (a and b);
    layer1_outputs(6402) <= a xor b;
    layer1_outputs(6403) <= not (a or b);
    layer1_outputs(6404) <= not a;
    layer1_outputs(6405) <= b;
    layer1_outputs(6406) <= a and not b;
    layer1_outputs(6407) <= b;
    layer1_outputs(6408) <= b;
    layer1_outputs(6409) <= not (a and b);
    layer1_outputs(6410) <= not a;
    layer1_outputs(6411) <= a;
    layer1_outputs(6412) <= not (a or b);
    layer1_outputs(6413) <= a and b;
    layer1_outputs(6414) <= a and not b;
    layer1_outputs(6415) <= not a;
    layer1_outputs(6416) <= b and not a;
    layer1_outputs(6417) <= a xor b;
    layer1_outputs(6418) <= a and not b;
    layer1_outputs(6419) <= a and b;
    layer1_outputs(6420) <= a or b;
    layer1_outputs(6421) <= not a;
    layer1_outputs(6422) <= not b or a;
    layer1_outputs(6423) <= b;
    layer1_outputs(6424) <= a;
    layer1_outputs(6425) <= not a;
    layer1_outputs(6426) <= not a;
    layer1_outputs(6427) <= b;
    layer1_outputs(6428) <= 1'b0;
    layer1_outputs(6429) <= a xor b;
    layer1_outputs(6430) <= not b or a;
    layer1_outputs(6431) <= a or b;
    layer1_outputs(6432) <= a;
    layer1_outputs(6433) <= b;
    layer1_outputs(6434) <= a xor b;
    layer1_outputs(6435) <= a xor b;
    layer1_outputs(6436) <= not (a or b);
    layer1_outputs(6437) <= not b;
    layer1_outputs(6438) <= not a;
    layer1_outputs(6439) <= a and b;
    layer1_outputs(6440) <= a;
    layer1_outputs(6441) <= not b;
    layer1_outputs(6442) <= not (a or b);
    layer1_outputs(6443) <= a;
    layer1_outputs(6444) <= not b or a;
    layer1_outputs(6445) <= not a or b;
    layer1_outputs(6446) <= not b;
    layer1_outputs(6447) <= not (a and b);
    layer1_outputs(6448) <= b;
    layer1_outputs(6449) <= not a;
    layer1_outputs(6450) <= not (a xor b);
    layer1_outputs(6451) <= not (a or b);
    layer1_outputs(6452) <= a xor b;
    layer1_outputs(6453) <= b and not a;
    layer1_outputs(6454) <= a or b;
    layer1_outputs(6455) <= not (a or b);
    layer1_outputs(6456) <= not a or b;
    layer1_outputs(6457) <= b;
    layer1_outputs(6458) <= a and b;
    layer1_outputs(6459) <= a or b;
    layer1_outputs(6460) <= a xor b;
    layer1_outputs(6461) <= a xor b;
    layer1_outputs(6462) <= not (a and b);
    layer1_outputs(6463) <= not b;
    layer1_outputs(6464) <= not a;
    layer1_outputs(6465) <= a xor b;
    layer1_outputs(6466) <= b and not a;
    layer1_outputs(6467) <= 1'b0;
    layer1_outputs(6468) <= b and not a;
    layer1_outputs(6469) <= b;
    layer1_outputs(6470) <= not b;
    layer1_outputs(6471) <= not (a and b);
    layer1_outputs(6472) <= b and not a;
    layer1_outputs(6473) <= b and not a;
    layer1_outputs(6474) <= a or b;
    layer1_outputs(6475) <= a and not b;
    layer1_outputs(6476) <= 1'b0;
    layer1_outputs(6477) <= not b;
    layer1_outputs(6478) <= not a;
    layer1_outputs(6479) <= not b or a;
    layer1_outputs(6480) <= a;
    layer1_outputs(6481) <= not a or b;
    layer1_outputs(6482) <= not b or a;
    layer1_outputs(6483) <= not a or b;
    layer1_outputs(6484) <= b;
    layer1_outputs(6485) <= b;
    layer1_outputs(6486) <= not (a or b);
    layer1_outputs(6487) <= not b;
    layer1_outputs(6488) <= not b;
    layer1_outputs(6489) <= not a or b;
    layer1_outputs(6490) <= a;
    layer1_outputs(6491) <= a and b;
    layer1_outputs(6492) <= not b;
    layer1_outputs(6493) <= not a;
    layer1_outputs(6494) <= not a;
    layer1_outputs(6495) <= b;
    layer1_outputs(6496) <= not (a xor b);
    layer1_outputs(6497) <= a and not b;
    layer1_outputs(6498) <= not b;
    layer1_outputs(6499) <= a or b;
    layer1_outputs(6500) <= a;
    layer1_outputs(6501) <= a xor b;
    layer1_outputs(6502) <= not b;
    layer1_outputs(6503) <= not (a or b);
    layer1_outputs(6504) <= not b;
    layer1_outputs(6505) <= not (a or b);
    layer1_outputs(6506) <= not b or a;
    layer1_outputs(6507) <= a and not b;
    layer1_outputs(6508) <= not a;
    layer1_outputs(6509) <= not a or b;
    layer1_outputs(6510) <= b and not a;
    layer1_outputs(6511) <= a or b;
    layer1_outputs(6512) <= a xor b;
    layer1_outputs(6513) <= not b or a;
    layer1_outputs(6514) <= a xor b;
    layer1_outputs(6515) <= a xor b;
    layer1_outputs(6516) <= a and not b;
    layer1_outputs(6517) <= not b or a;
    layer1_outputs(6518) <= b;
    layer1_outputs(6519) <= not b or a;
    layer1_outputs(6520) <= b;
    layer1_outputs(6521) <= not a;
    layer1_outputs(6522) <= b;
    layer1_outputs(6523) <= not (a and b);
    layer1_outputs(6524) <= not a;
    layer1_outputs(6525) <= a or b;
    layer1_outputs(6526) <= not (a and b);
    layer1_outputs(6527) <= a xor b;
    layer1_outputs(6528) <= not (a and b);
    layer1_outputs(6529) <= not a or b;
    layer1_outputs(6530) <= a and b;
    layer1_outputs(6531) <= a and not b;
    layer1_outputs(6532) <= b;
    layer1_outputs(6533) <= not a;
    layer1_outputs(6534) <= not (a or b);
    layer1_outputs(6535) <= not b;
    layer1_outputs(6536) <= a xor b;
    layer1_outputs(6537) <= a;
    layer1_outputs(6538) <= not (a xor b);
    layer1_outputs(6539) <= a and not b;
    layer1_outputs(6540) <= b;
    layer1_outputs(6541) <= not b;
    layer1_outputs(6542) <= not (a or b);
    layer1_outputs(6543) <= not b or a;
    layer1_outputs(6544) <= not (a or b);
    layer1_outputs(6545) <= not (a xor b);
    layer1_outputs(6546) <= a or b;
    layer1_outputs(6547) <= a or b;
    layer1_outputs(6548) <= b and not a;
    layer1_outputs(6549) <= a xor b;
    layer1_outputs(6550) <= not a;
    layer1_outputs(6551) <= not (a xor b);
    layer1_outputs(6552) <= b and not a;
    layer1_outputs(6553) <= a xor b;
    layer1_outputs(6554) <= a and b;
    layer1_outputs(6555) <= not (a and b);
    layer1_outputs(6556) <= not b;
    layer1_outputs(6557) <= a and b;
    layer1_outputs(6558) <= not (a or b);
    layer1_outputs(6559) <= not b or a;
    layer1_outputs(6560) <= not (a and b);
    layer1_outputs(6561) <= not (a xor b);
    layer1_outputs(6562) <= a and b;
    layer1_outputs(6563) <= b and not a;
    layer1_outputs(6564) <= not a or b;
    layer1_outputs(6565) <= not a;
    layer1_outputs(6566) <= not (a xor b);
    layer1_outputs(6567) <= a xor b;
    layer1_outputs(6568) <= a;
    layer1_outputs(6569) <= a and not b;
    layer1_outputs(6570) <= a and not b;
    layer1_outputs(6571) <= b;
    layer1_outputs(6572) <= b;
    layer1_outputs(6573) <= b and not a;
    layer1_outputs(6574) <= b;
    layer1_outputs(6575) <= not a or b;
    layer1_outputs(6576) <= not a or b;
    layer1_outputs(6577) <= 1'b1;
    layer1_outputs(6578) <= a;
    layer1_outputs(6579) <= a;
    layer1_outputs(6580) <= a and b;
    layer1_outputs(6581) <= a and b;
    layer1_outputs(6582) <= b;
    layer1_outputs(6583) <= not b or a;
    layer1_outputs(6584) <= not a;
    layer1_outputs(6585) <= a and b;
    layer1_outputs(6586) <= b and not a;
    layer1_outputs(6587) <= not a or b;
    layer1_outputs(6588) <= a;
    layer1_outputs(6589) <= not b;
    layer1_outputs(6590) <= b and not a;
    layer1_outputs(6591) <= a or b;
    layer1_outputs(6592) <= not (a xor b);
    layer1_outputs(6593) <= not a;
    layer1_outputs(6594) <= not (a or b);
    layer1_outputs(6595) <= not a or b;
    layer1_outputs(6596) <= not (a and b);
    layer1_outputs(6597) <= a and not b;
    layer1_outputs(6598) <= not a or b;
    layer1_outputs(6599) <= not (a or b);
    layer1_outputs(6600) <= b;
    layer1_outputs(6601) <= not (a or b);
    layer1_outputs(6602) <= b;
    layer1_outputs(6603) <= a and not b;
    layer1_outputs(6604) <= not b;
    layer1_outputs(6605) <= not a or b;
    layer1_outputs(6606) <= not a or b;
    layer1_outputs(6607) <= not b or a;
    layer1_outputs(6608) <= not a;
    layer1_outputs(6609) <= not b;
    layer1_outputs(6610) <= a and not b;
    layer1_outputs(6611) <= not b or a;
    layer1_outputs(6612) <= a and not b;
    layer1_outputs(6613) <= not (a xor b);
    layer1_outputs(6614) <= not (a xor b);
    layer1_outputs(6615) <= not (a xor b);
    layer1_outputs(6616) <= not a;
    layer1_outputs(6617) <= a or b;
    layer1_outputs(6618) <= not a or b;
    layer1_outputs(6619) <= not a or b;
    layer1_outputs(6620) <= not a or b;
    layer1_outputs(6621) <= not a;
    layer1_outputs(6622) <= not b or a;
    layer1_outputs(6623) <= not a or b;
    layer1_outputs(6624) <= not a or b;
    layer1_outputs(6625) <= not b;
    layer1_outputs(6626) <= b;
    layer1_outputs(6627) <= b;
    layer1_outputs(6628) <= not (a xor b);
    layer1_outputs(6629) <= a or b;
    layer1_outputs(6630) <= b;
    layer1_outputs(6631) <= not a or b;
    layer1_outputs(6632) <= a or b;
    layer1_outputs(6633) <= b;
    layer1_outputs(6634) <= not a;
    layer1_outputs(6635) <= not b or a;
    layer1_outputs(6636) <= a;
    layer1_outputs(6637) <= not a or b;
    layer1_outputs(6638) <= b and not a;
    layer1_outputs(6639) <= b;
    layer1_outputs(6640) <= not b or a;
    layer1_outputs(6641) <= not (a or b);
    layer1_outputs(6642) <= not b;
    layer1_outputs(6643) <= not b or a;
    layer1_outputs(6644) <= not a or b;
    layer1_outputs(6645) <= not a;
    layer1_outputs(6646) <= a xor b;
    layer1_outputs(6647) <= not (a xor b);
    layer1_outputs(6648) <= b;
    layer1_outputs(6649) <= not (a xor b);
    layer1_outputs(6650) <= not a;
    layer1_outputs(6651) <= a and b;
    layer1_outputs(6652) <= b;
    layer1_outputs(6653) <= a;
    layer1_outputs(6654) <= not b or a;
    layer1_outputs(6655) <= not a;
    layer1_outputs(6656) <= a or b;
    layer1_outputs(6657) <= a;
    layer1_outputs(6658) <= b;
    layer1_outputs(6659) <= a;
    layer1_outputs(6660) <= not (a xor b);
    layer1_outputs(6661) <= not b;
    layer1_outputs(6662) <= not a or b;
    layer1_outputs(6663) <= not b;
    layer1_outputs(6664) <= not a;
    layer1_outputs(6665) <= not a;
    layer1_outputs(6666) <= a and b;
    layer1_outputs(6667) <= a xor b;
    layer1_outputs(6668) <= b;
    layer1_outputs(6669) <= not (a xor b);
    layer1_outputs(6670) <= not b or a;
    layer1_outputs(6671) <= a xor b;
    layer1_outputs(6672) <= a and b;
    layer1_outputs(6673) <= not (a and b);
    layer1_outputs(6674) <= not (a xor b);
    layer1_outputs(6675) <= not a;
    layer1_outputs(6676) <= not b;
    layer1_outputs(6677) <= not a or b;
    layer1_outputs(6678) <= a and not b;
    layer1_outputs(6679) <= b and not a;
    layer1_outputs(6680) <= not (a and b);
    layer1_outputs(6681) <= a xor b;
    layer1_outputs(6682) <= a;
    layer1_outputs(6683) <= 1'b1;
    layer1_outputs(6684) <= not a or b;
    layer1_outputs(6685) <= not a or b;
    layer1_outputs(6686) <= b;
    layer1_outputs(6687) <= a xor b;
    layer1_outputs(6688) <= b;
    layer1_outputs(6689) <= not (a and b);
    layer1_outputs(6690) <= a or b;
    layer1_outputs(6691) <= a and not b;
    layer1_outputs(6692) <= not a or b;
    layer1_outputs(6693) <= a;
    layer1_outputs(6694) <= a;
    layer1_outputs(6695) <= not b or a;
    layer1_outputs(6696) <= not a;
    layer1_outputs(6697) <= a and b;
    layer1_outputs(6698) <= not (a or b);
    layer1_outputs(6699) <= a xor b;
    layer1_outputs(6700) <= b and not a;
    layer1_outputs(6701) <= a or b;
    layer1_outputs(6702) <= not (a or b);
    layer1_outputs(6703) <= not (a or b);
    layer1_outputs(6704) <= not b;
    layer1_outputs(6705) <= a xor b;
    layer1_outputs(6706) <= not b or a;
    layer1_outputs(6707) <= a and not b;
    layer1_outputs(6708) <= not a or b;
    layer1_outputs(6709) <= not a;
    layer1_outputs(6710) <= not b;
    layer1_outputs(6711) <= not a;
    layer1_outputs(6712) <= a;
    layer1_outputs(6713) <= not a;
    layer1_outputs(6714) <= a or b;
    layer1_outputs(6715) <= a and not b;
    layer1_outputs(6716) <= not b or a;
    layer1_outputs(6717) <= b;
    layer1_outputs(6718) <= a;
    layer1_outputs(6719) <= not a;
    layer1_outputs(6720) <= not (a and b);
    layer1_outputs(6721) <= not b;
    layer1_outputs(6722) <= a and b;
    layer1_outputs(6723) <= a xor b;
    layer1_outputs(6724) <= a and b;
    layer1_outputs(6725) <= not a;
    layer1_outputs(6726) <= not (a xor b);
    layer1_outputs(6727) <= a and b;
    layer1_outputs(6728) <= not b or a;
    layer1_outputs(6729) <= a;
    layer1_outputs(6730) <= not a;
    layer1_outputs(6731) <= not (a or b);
    layer1_outputs(6732) <= not (a xor b);
    layer1_outputs(6733) <= 1'b1;
    layer1_outputs(6734) <= not (a xor b);
    layer1_outputs(6735) <= a and not b;
    layer1_outputs(6736) <= a and b;
    layer1_outputs(6737) <= a and not b;
    layer1_outputs(6738) <= not (a or b);
    layer1_outputs(6739) <= not b;
    layer1_outputs(6740) <= not b;
    layer1_outputs(6741) <= not b or a;
    layer1_outputs(6742) <= b and not a;
    layer1_outputs(6743) <= b;
    layer1_outputs(6744) <= not b;
    layer1_outputs(6745) <= not a;
    layer1_outputs(6746) <= a and b;
    layer1_outputs(6747) <= b and not a;
    layer1_outputs(6748) <= a and b;
    layer1_outputs(6749) <= b and not a;
    layer1_outputs(6750) <= not (a and b);
    layer1_outputs(6751) <= b and not a;
    layer1_outputs(6752) <= not b;
    layer1_outputs(6753) <= not a or b;
    layer1_outputs(6754) <= a and b;
    layer1_outputs(6755) <= not (a or b);
    layer1_outputs(6756) <= b;
    layer1_outputs(6757) <= not (a xor b);
    layer1_outputs(6758) <= a or b;
    layer1_outputs(6759) <= a and b;
    layer1_outputs(6760) <= not (a or b);
    layer1_outputs(6761) <= a xor b;
    layer1_outputs(6762) <= not b or a;
    layer1_outputs(6763) <= not b;
    layer1_outputs(6764) <= not (a xor b);
    layer1_outputs(6765) <= not a;
    layer1_outputs(6766) <= not b or a;
    layer1_outputs(6767) <= a;
    layer1_outputs(6768) <= not b;
    layer1_outputs(6769) <= not (a or b);
    layer1_outputs(6770) <= b;
    layer1_outputs(6771) <= a;
    layer1_outputs(6772) <= not (a and b);
    layer1_outputs(6773) <= not b or a;
    layer1_outputs(6774) <= a and not b;
    layer1_outputs(6775) <= a;
    layer1_outputs(6776) <= b and not a;
    layer1_outputs(6777) <= 1'b1;
    layer1_outputs(6778) <= a xor b;
    layer1_outputs(6779) <= b;
    layer1_outputs(6780) <= not (a or b);
    layer1_outputs(6781) <= not (a and b);
    layer1_outputs(6782) <= a and not b;
    layer1_outputs(6783) <= not (a and b);
    layer1_outputs(6784) <= a and b;
    layer1_outputs(6785) <= a or b;
    layer1_outputs(6786) <= a xor b;
    layer1_outputs(6787) <= a or b;
    layer1_outputs(6788) <= not (a xor b);
    layer1_outputs(6789) <= b;
    layer1_outputs(6790) <= not (a or b);
    layer1_outputs(6791) <= a and not b;
    layer1_outputs(6792) <= a xor b;
    layer1_outputs(6793) <= 1'b1;
    layer1_outputs(6794) <= b and not a;
    layer1_outputs(6795) <= a and not b;
    layer1_outputs(6796) <= not b;
    layer1_outputs(6797) <= b and not a;
    layer1_outputs(6798) <= not b;
    layer1_outputs(6799) <= a;
    layer1_outputs(6800) <= not a or b;
    layer1_outputs(6801) <= a and not b;
    layer1_outputs(6802) <= a;
    layer1_outputs(6803) <= b;
    layer1_outputs(6804) <= not (a and b);
    layer1_outputs(6805) <= not b;
    layer1_outputs(6806) <= not b or a;
    layer1_outputs(6807) <= b and not a;
    layer1_outputs(6808) <= not b;
    layer1_outputs(6809) <= not a;
    layer1_outputs(6810) <= not a or b;
    layer1_outputs(6811) <= a;
    layer1_outputs(6812) <= not b;
    layer1_outputs(6813) <= not b;
    layer1_outputs(6814) <= a and not b;
    layer1_outputs(6815) <= a and not b;
    layer1_outputs(6816) <= not a or b;
    layer1_outputs(6817) <= a;
    layer1_outputs(6818) <= a;
    layer1_outputs(6819) <= not (a xor b);
    layer1_outputs(6820) <= not b;
    layer1_outputs(6821) <= not (a xor b);
    layer1_outputs(6822) <= not (a and b);
    layer1_outputs(6823) <= a xor b;
    layer1_outputs(6824) <= a xor b;
    layer1_outputs(6825) <= not (a xor b);
    layer1_outputs(6826) <= a;
    layer1_outputs(6827) <= not a;
    layer1_outputs(6828) <= a and b;
    layer1_outputs(6829) <= not b;
    layer1_outputs(6830) <= not b;
    layer1_outputs(6831) <= a;
    layer1_outputs(6832) <= a;
    layer1_outputs(6833) <= a;
    layer1_outputs(6834) <= not a;
    layer1_outputs(6835) <= a xor b;
    layer1_outputs(6836) <= a xor b;
    layer1_outputs(6837) <= a and not b;
    layer1_outputs(6838) <= not a or b;
    layer1_outputs(6839) <= not (a or b);
    layer1_outputs(6840) <= b and not a;
    layer1_outputs(6841) <= a or b;
    layer1_outputs(6842) <= b and not a;
    layer1_outputs(6843) <= b and not a;
    layer1_outputs(6844) <= not b or a;
    layer1_outputs(6845) <= b;
    layer1_outputs(6846) <= b;
    layer1_outputs(6847) <= a or b;
    layer1_outputs(6848) <= a;
    layer1_outputs(6849) <= a or b;
    layer1_outputs(6850) <= b;
    layer1_outputs(6851) <= not b;
    layer1_outputs(6852) <= not a or b;
    layer1_outputs(6853) <= b;
    layer1_outputs(6854) <= 1'b1;
    layer1_outputs(6855) <= not (a and b);
    layer1_outputs(6856) <= not a;
    layer1_outputs(6857) <= b and not a;
    layer1_outputs(6858) <= a and not b;
    layer1_outputs(6859) <= a;
    layer1_outputs(6860) <= not b or a;
    layer1_outputs(6861) <= not a;
    layer1_outputs(6862) <= not b;
    layer1_outputs(6863) <= b and not a;
    layer1_outputs(6864) <= not (a or b);
    layer1_outputs(6865) <= not a;
    layer1_outputs(6866) <= b;
    layer1_outputs(6867) <= not (a or b);
    layer1_outputs(6868) <= a and not b;
    layer1_outputs(6869) <= a or b;
    layer1_outputs(6870) <= a and not b;
    layer1_outputs(6871) <= b and not a;
    layer1_outputs(6872) <= a or b;
    layer1_outputs(6873) <= not a or b;
    layer1_outputs(6874) <= a;
    layer1_outputs(6875) <= a and b;
    layer1_outputs(6876) <= not (a and b);
    layer1_outputs(6877) <= not (a and b);
    layer1_outputs(6878) <= not (a or b);
    layer1_outputs(6879) <= 1'b0;
    layer1_outputs(6880) <= not (a or b);
    layer1_outputs(6881) <= a or b;
    layer1_outputs(6882) <= a and b;
    layer1_outputs(6883) <= not b;
    layer1_outputs(6884) <= not (a xor b);
    layer1_outputs(6885) <= a;
    layer1_outputs(6886) <= a;
    layer1_outputs(6887) <= not b;
    layer1_outputs(6888) <= a and b;
    layer1_outputs(6889) <= not (a xor b);
    layer1_outputs(6890) <= a or b;
    layer1_outputs(6891) <= a or b;
    layer1_outputs(6892) <= b;
    layer1_outputs(6893) <= not (a xor b);
    layer1_outputs(6894) <= b;
    layer1_outputs(6895) <= b;
    layer1_outputs(6896) <= not (a and b);
    layer1_outputs(6897) <= b;
    layer1_outputs(6898) <= not a;
    layer1_outputs(6899) <= 1'b0;
    layer1_outputs(6900) <= a;
    layer1_outputs(6901) <= a or b;
    layer1_outputs(6902) <= a;
    layer1_outputs(6903) <= a;
    layer1_outputs(6904) <= not b or a;
    layer1_outputs(6905) <= a and b;
    layer1_outputs(6906) <= b;
    layer1_outputs(6907) <= a xor b;
    layer1_outputs(6908) <= not (a and b);
    layer1_outputs(6909) <= a or b;
    layer1_outputs(6910) <= a xor b;
    layer1_outputs(6911) <= b;
    layer1_outputs(6912) <= b and not a;
    layer1_outputs(6913) <= not b;
    layer1_outputs(6914) <= not b;
    layer1_outputs(6915) <= b;
    layer1_outputs(6916) <= not a;
    layer1_outputs(6917) <= not (a and b);
    layer1_outputs(6918) <= not b or a;
    layer1_outputs(6919) <= not b;
    layer1_outputs(6920) <= not b or a;
    layer1_outputs(6921) <= a and not b;
    layer1_outputs(6922) <= not (a or b);
    layer1_outputs(6923) <= not (a and b);
    layer1_outputs(6924) <= not a or b;
    layer1_outputs(6925) <= not (a or b);
    layer1_outputs(6926) <= b;
    layer1_outputs(6927) <= not a or b;
    layer1_outputs(6928) <= a;
    layer1_outputs(6929) <= not b;
    layer1_outputs(6930) <= b;
    layer1_outputs(6931) <= a and not b;
    layer1_outputs(6932) <= not b;
    layer1_outputs(6933) <= not b or a;
    layer1_outputs(6934) <= a xor b;
    layer1_outputs(6935) <= not a;
    layer1_outputs(6936) <= 1'b0;
    layer1_outputs(6937) <= not a;
    layer1_outputs(6938) <= a or b;
    layer1_outputs(6939) <= a and b;
    layer1_outputs(6940) <= b and not a;
    layer1_outputs(6941) <= a;
    layer1_outputs(6942) <= b;
    layer1_outputs(6943) <= not b;
    layer1_outputs(6944) <= a or b;
    layer1_outputs(6945) <= not (a or b);
    layer1_outputs(6946) <= a and b;
    layer1_outputs(6947) <= not a;
    layer1_outputs(6948) <= not (a or b);
    layer1_outputs(6949) <= b;
    layer1_outputs(6950) <= not (a or b);
    layer1_outputs(6951) <= not a or b;
    layer1_outputs(6952) <= a;
    layer1_outputs(6953) <= a;
    layer1_outputs(6954) <= not a;
    layer1_outputs(6955) <= b;
    layer1_outputs(6956) <= not (a xor b);
    layer1_outputs(6957) <= a and b;
    layer1_outputs(6958) <= b and not a;
    layer1_outputs(6959) <= a and b;
    layer1_outputs(6960) <= not b;
    layer1_outputs(6961) <= not a;
    layer1_outputs(6962) <= b;
    layer1_outputs(6963) <= not (a xor b);
    layer1_outputs(6964) <= a and b;
    layer1_outputs(6965) <= b;
    layer1_outputs(6966) <= not a or b;
    layer1_outputs(6967) <= not b or a;
    layer1_outputs(6968) <= a and not b;
    layer1_outputs(6969) <= not (a and b);
    layer1_outputs(6970) <= not a;
    layer1_outputs(6971) <= b;
    layer1_outputs(6972) <= b;
    layer1_outputs(6973) <= a xor b;
    layer1_outputs(6974) <= a and not b;
    layer1_outputs(6975) <= b;
    layer1_outputs(6976) <= a or b;
    layer1_outputs(6977) <= not b;
    layer1_outputs(6978) <= a and b;
    layer1_outputs(6979) <= not (a xor b);
    layer1_outputs(6980) <= not b;
    layer1_outputs(6981) <= not a;
    layer1_outputs(6982) <= not a;
    layer1_outputs(6983) <= not (a and b);
    layer1_outputs(6984) <= a and b;
    layer1_outputs(6985) <= b;
    layer1_outputs(6986) <= not a;
    layer1_outputs(6987) <= 1'b0;
    layer1_outputs(6988) <= not (a and b);
    layer1_outputs(6989) <= a xor b;
    layer1_outputs(6990) <= not (a or b);
    layer1_outputs(6991) <= not b;
    layer1_outputs(6992) <= a xor b;
    layer1_outputs(6993) <= not (a or b);
    layer1_outputs(6994) <= not (a xor b);
    layer1_outputs(6995) <= not a or b;
    layer1_outputs(6996) <= not (a xor b);
    layer1_outputs(6997) <= not a;
    layer1_outputs(6998) <= b and not a;
    layer1_outputs(6999) <= a and b;
    layer1_outputs(7000) <= not (a and b);
    layer1_outputs(7001) <= a and b;
    layer1_outputs(7002) <= not b;
    layer1_outputs(7003) <= a and not b;
    layer1_outputs(7004) <= b and not a;
    layer1_outputs(7005) <= not a;
    layer1_outputs(7006) <= not (a xor b);
    layer1_outputs(7007) <= b and not a;
    layer1_outputs(7008) <= not a or b;
    layer1_outputs(7009) <= not b;
    layer1_outputs(7010) <= not a or b;
    layer1_outputs(7011) <= a;
    layer1_outputs(7012) <= not b or a;
    layer1_outputs(7013) <= a and not b;
    layer1_outputs(7014) <= a or b;
    layer1_outputs(7015) <= not b or a;
    layer1_outputs(7016) <= b;
    layer1_outputs(7017) <= b and not a;
    layer1_outputs(7018) <= not b;
    layer1_outputs(7019) <= b;
    layer1_outputs(7020) <= a xor b;
    layer1_outputs(7021) <= not (a and b);
    layer1_outputs(7022) <= a xor b;
    layer1_outputs(7023) <= b and not a;
    layer1_outputs(7024) <= a;
    layer1_outputs(7025) <= a;
    layer1_outputs(7026) <= b and not a;
    layer1_outputs(7027) <= a;
    layer1_outputs(7028) <= not a;
    layer1_outputs(7029) <= not a or b;
    layer1_outputs(7030) <= a xor b;
    layer1_outputs(7031) <= not (a xor b);
    layer1_outputs(7032) <= not b;
    layer1_outputs(7033) <= not (a or b);
    layer1_outputs(7034) <= not b;
    layer1_outputs(7035) <= not a;
    layer1_outputs(7036) <= not a or b;
    layer1_outputs(7037) <= a;
    layer1_outputs(7038) <= not b or a;
    layer1_outputs(7039) <= not a or b;
    layer1_outputs(7040) <= a and not b;
    layer1_outputs(7041) <= b;
    layer1_outputs(7042) <= not a or b;
    layer1_outputs(7043) <= a xor b;
    layer1_outputs(7044) <= not (a or b);
    layer1_outputs(7045) <= 1'b0;
    layer1_outputs(7046) <= not a or b;
    layer1_outputs(7047) <= a and not b;
    layer1_outputs(7048) <= b;
    layer1_outputs(7049) <= not a;
    layer1_outputs(7050) <= a;
    layer1_outputs(7051) <= b;
    layer1_outputs(7052) <= not (a xor b);
    layer1_outputs(7053) <= a and b;
    layer1_outputs(7054) <= a;
    layer1_outputs(7055) <= not b;
    layer1_outputs(7056) <= not (a and b);
    layer1_outputs(7057) <= not a or b;
    layer1_outputs(7058) <= not a;
    layer1_outputs(7059) <= a;
    layer1_outputs(7060) <= a and not b;
    layer1_outputs(7061) <= a xor b;
    layer1_outputs(7062) <= b;
    layer1_outputs(7063) <= not b;
    layer1_outputs(7064) <= a xor b;
    layer1_outputs(7065) <= not (a and b);
    layer1_outputs(7066) <= not a;
    layer1_outputs(7067) <= not (a or b);
    layer1_outputs(7068) <= not a or b;
    layer1_outputs(7069) <= a and not b;
    layer1_outputs(7070) <= not b;
    layer1_outputs(7071) <= not b;
    layer1_outputs(7072) <= not (a and b);
    layer1_outputs(7073) <= not (a xor b);
    layer1_outputs(7074) <= a and b;
    layer1_outputs(7075) <= not (a xor b);
    layer1_outputs(7076) <= a and not b;
    layer1_outputs(7077) <= not (a xor b);
    layer1_outputs(7078) <= a or b;
    layer1_outputs(7079) <= not a;
    layer1_outputs(7080) <= a and not b;
    layer1_outputs(7081) <= not b;
    layer1_outputs(7082) <= not a;
    layer1_outputs(7083) <= a;
    layer1_outputs(7084) <= a or b;
    layer1_outputs(7085) <= not b;
    layer1_outputs(7086) <= not (a and b);
    layer1_outputs(7087) <= 1'b1;
    layer1_outputs(7088) <= not (a and b);
    layer1_outputs(7089) <= b;
    layer1_outputs(7090) <= a;
    layer1_outputs(7091) <= a and not b;
    layer1_outputs(7092) <= not (a or b);
    layer1_outputs(7093) <= b and not a;
    layer1_outputs(7094) <= a or b;
    layer1_outputs(7095) <= not a;
    layer1_outputs(7096) <= a and not b;
    layer1_outputs(7097) <= not a;
    layer1_outputs(7098) <= b;
    layer1_outputs(7099) <= a and not b;
    layer1_outputs(7100) <= a or b;
    layer1_outputs(7101) <= not a or b;
    layer1_outputs(7102) <= not (a xor b);
    layer1_outputs(7103) <= not (a xor b);
    layer1_outputs(7104) <= not a;
    layer1_outputs(7105) <= not b;
    layer1_outputs(7106) <= not a;
    layer1_outputs(7107) <= b and not a;
    layer1_outputs(7108) <= not a;
    layer1_outputs(7109) <= a or b;
    layer1_outputs(7110) <= not a or b;
    layer1_outputs(7111) <= not b;
    layer1_outputs(7112) <= not b;
    layer1_outputs(7113) <= not a or b;
    layer1_outputs(7114) <= not (a and b);
    layer1_outputs(7115) <= b;
    layer1_outputs(7116) <= a and b;
    layer1_outputs(7117) <= a;
    layer1_outputs(7118) <= not b;
    layer1_outputs(7119) <= not b or a;
    layer1_outputs(7120) <= not a or b;
    layer1_outputs(7121) <= not a;
    layer1_outputs(7122) <= not (a and b);
    layer1_outputs(7123) <= not a;
    layer1_outputs(7124) <= not (a xor b);
    layer1_outputs(7125) <= b and not a;
    layer1_outputs(7126) <= b;
    layer1_outputs(7127) <= not a or b;
    layer1_outputs(7128) <= a xor b;
    layer1_outputs(7129) <= not (a and b);
    layer1_outputs(7130) <= b and not a;
    layer1_outputs(7131) <= not (a xor b);
    layer1_outputs(7132) <= a xor b;
    layer1_outputs(7133) <= b;
    layer1_outputs(7134) <= b;
    layer1_outputs(7135) <= a;
    layer1_outputs(7136) <= b;
    layer1_outputs(7137) <= not b;
    layer1_outputs(7138) <= b;
    layer1_outputs(7139) <= not (a or b);
    layer1_outputs(7140) <= a;
    layer1_outputs(7141) <= not (a and b);
    layer1_outputs(7142) <= not b or a;
    layer1_outputs(7143) <= a or b;
    layer1_outputs(7144) <= not b or a;
    layer1_outputs(7145) <= a and b;
    layer1_outputs(7146) <= not a;
    layer1_outputs(7147) <= a and b;
    layer1_outputs(7148) <= a and b;
    layer1_outputs(7149) <= b;
    layer1_outputs(7150) <= a and b;
    layer1_outputs(7151) <= not (a and b);
    layer1_outputs(7152) <= a and b;
    layer1_outputs(7153) <= a;
    layer1_outputs(7154) <= not b;
    layer1_outputs(7155) <= 1'b0;
    layer1_outputs(7156) <= not a;
    layer1_outputs(7157) <= b;
    layer1_outputs(7158) <= not (a and b);
    layer1_outputs(7159) <= b;
    layer1_outputs(7160) <= a or b;
    layer1_outputs(7161) <= b and not a;
    layer1_outputs(7162) <= not b;
    layer1_outputs(7163) <= not b or a;
    layer1_outputs(7164) <= not b or a;
    layer1_outputs(7165) <= not a or b;
    layer1_outputs(7166) <= not b;
    layer1_outputs(7167) <= b and not a;
    layer1_outputs(7168) <= not (a or b);
    layer1_outputs(7169) <= not (a and b);
    layer1_outputs(7170) <= a;
    layer1_outputs(7171) <= not a;
    layer1_outputs(7172) <= not a;
    layer1_outputs(7173) <= not (a and b);
    layer1_outputs(7174) <= b;
    layer1_outputs(7175) <= not a or b;
    layer1_outputs(7176) <= a or b;
    layer1_outputs(7177) <= not a;
    layer1_outputs(7178) <= not (a or b);
    layer1_outputs(7179) <= not b;
    layer1_outputs(7180) <= 1'b0;
    layer1_outputs(7181) <= not a;
    layer1_outputs(7182) <= b;
    layer1_outputs(7183) <= not (a xor b);
    layer1_outputs(7184) <= 1'b1;
    layer1_outputs(7185) <= b and not a;
    layer1_outputs(7186) <= a or b;
    layer1_outputs(7187) <= a;
    layer1_outputs(7188) <= a and not b;
    layer1_outputs(7189) <= not (a and b);
    layer1_outputs(7190) <= not (a or b);
    layer1_outputs(7191) <= not a or b;
    layer1_outputs(7192) <= not a or b;
    layer1_outputs(7193) <= b;
    layer1_outputs(7194) <= not (a or b);
    layer1_outputs(7195) <= a and b;
    layer1_outputs(7196) <= not a or b;
    layer1_outputs(7197) <= a;
    layer1_outputs(7198) <= a;
    layer1_outputs(7199) <= not b;
    layer1_outputs(7200) <= a xor b;
    layer1_outputs(7201) <= not a or b;
    layer1_outputs(7202) <= not (a and b);
    layer1_outputs(7203) <= a and b;
    layer1_outputs(7204) <= a and b;
    layer1_outputs(7205) <= b and not a;
    layer1_outputs(7206) <= not (a and b);
    layer1_outputs(7207) <= 1'b0;
    layer1_outputs(7208) <= not b;
    layer1_outputs(7209) <= b;
    layer1_outputs(7210) <= a and b;
    layer1_outputs(7211) <= b and not a;
    layer1_outputs(7212) <= not b or a;
    layer1_outputs(7213) <= not b or a;
    layer1_outputs(7214) <= a and not b;
    layer1_outputs(7215) <= not (a xor b);
    layer1_outputs(7216) <= a;
    layer1_outputs(7217) <= a;
    layer1_outputs(7218) <= b;
    layer1_outputs(7219) <= not b;
    layer1_outputs(7220) <= not (a and b);
    layer1_outputs(7221) <= a;
    layer1_outputs(7222) <= a and b;
    layer1_outputs(7223) <= not a;
    layer1_outputs(7224) <= not (a and b);
    layer1_outputs(7225) <= a or b;
    layer1_outputs(7226) <= not (a or b);
    layer1_outputs(7227) <= not (a and b);
    layer1_outputs(7228) <= not (a or b);
    layer1_outputs(7229) <= a;
    layer1_outputs(7230) <= not a;
    layer1_outputs(7231) <= not b or a;
    layer1_outputs(7232) <= not a or b;
    layer1_outputs(7233) <= a and not b;
    layer1_outputs(7234) <= not b;
    layer1_outputs(7235) <= not b;
    layer1_outputs(7236) <= not b;
    layer1_outputs(7237) <= a;
    layer1_outputs(7238) <= b;
    layer1_outputs(7239) <= a and b;
    layer1_outputs(7240) <= a and b;
    layer1_outputs(7241) <= not b;
    layer1_outputs(7242) <= a and b;
    layer1_outputs(7243) <= a and b;
    layer1_outputs(7244) <= not a or b;
    layer1_outputs(7245) <= a xor b;
    layer1_outputs(7246) <= a and not b;
    layer1_outputs(7247) <= a;
    layer1_outputs(7248) <= not (a or b);
    layer1_outputs(7249) <= a or b;
    layer1_outputs(7250) <= not a or b;
    layer1_outputs(7251) <= not b;
    layer1_outputs(7252) <= b;
    layer1_outputs(7253) <= b and not a;
    layer1_outputs(7254) <= a;
    layer1_outputs(7255) <= a and b;
    layer1_outputs(7256) <= a;
    layer1_outputs(7257) <= not (a and b);
    layer1_outputs(7258) <= a;
    layer1_outputs(7259) <= not (a or b);
    layer1_outputs(7260) <= a or b;
    layer1_outputs(7261) <= 1'b1;
    layer1_outputs(7262) <= not a;
    layer1_outputs(7263) <= a;
    layer1_outputs(7264) <= a and not b;
    layer1_outputs(7265) <= a xor b;
    layer1_outputs(7266) <= b and not a;
    layer1_outputs(7267) <= a or b;
    layer1_outputs(7268) <= not (a xor b);
    layer1_outputs(7269) <= not (a xor b);
    layer1_outputs(7270) <= not b or a;
    layer1_outputs(7271) <= 1'b0;
    layer1_outputs(7272) <= not (a or b);
    layer1_outputs(7273) <= not (a xor b);
    layer1_outputs(7274) <= not (a and b);
    layer1_outputs(7275) <= not b;
    layer1_outputs(7276) <= a xor b;
    layer1_outputs(7277) <= b;
    layer1_outputs(7278) <= a xor b;
    layer1_outputs(7279) <= a xor b;
    layer1_outputs(7280) <= not a;
    layer1_outputs(7281) <= a xor b;
    layer1_outputs(7282) <= not (a xor b);
    layer1_outputs(7283) <= not a;
    layer1_outputs(7284) <= not b;
    layer1_outputs(7285) <= not a;
    layer1_outputs(7286) <= a and not b;
    layer1_outputs(7287) <= b and not a;
    layer1_outputs(7288) <= a;
    layer1_outputs(7289) <= b and not a;
    layer1_outputs(7290) <= not b;
    layer1_outputs(7291) <= a or b;
    layer1_outputs(7292) <= not a or b;
    layer1_outputs(7293) <= b;
    layer1_outputs(7294) <= b;
    layer1_outputs(7295) <= not (a xor b);
    layer1_outputs(7296) <= not b;
    layer1_outputs(7297) <= not (a xor b);
    layer1_outputs(7298) <= a or b;
    layer1_outputs(7299) <= a or b;
    layer1_outputs(7300) <= a and not b;
    layer1_outputs(7301) <= a and not b;
    layer1_outputs(7302) <= a xor b;
    layer1_outputs(7303) <= a or b;
    layer1_outputs(7304) <= b;
    layer1_outputs(7305) <= a and not b;
    layer1_outputs(7306) <= b and not a;
    layer1_outputs(7307) <= a;
    layer1_outputs(7308) <= not b;
    layer1_outputs(7309) <= not (a or b);
    layer1_outputs(7310) <= a and not b;
    layer1_outputs(7311) <= not a or b;
    layer1_outputs(7312) <= a xor b;
    layer1_outputs(7313) <= not b;
    layer1_outputs(7314) <= a or b;
    layer1_outputs(7315) <= a and not b;
    layer1_outputs(7316) <= b;
    layer1_outputs(7317) <= a and not b;
    layer1_outputs(7318) <= not (a or b);
    layer1_outputs(7319) <= a or b;
    layer1_outputs(7320) <= b;
    layer1_outputs(7321) <= not a or b;
    layer1_outputs(7322) <= not a;
    layer1_outputs(7323) <= not a;
    layer1_outputs(7324) <= not a;
    layer1_outputs(7325) <= not (a or b);
    layer1_outputs(7326) <= not a;
    layer1_outputs(7327) <= b and not a;
    layer1_outputs(7328) <= a or b;
    layer1_outputs(7329) <= not a;
    layer1_outputs(7330) <= not a or b;
    layer1_outputs(7331) <= 1'b0;
    layer1_outputs(7332) <= b;
    layer1_outputs(7333) <= b and not a;
    layer1_outputs(7334) <= a and b;
    layer1_outputs(7335) <= not (a and b);
    layer1_outputs(7336) <= not (a xor b);
    layer1_outputs(7337) <= a and b;
    layer1_outputs(7338) <= not b;
    layer1_outputs(7339) <= a and b;
    layer1_outputs(7340) <= a and b;
    layer1_outputs(7341) <= not (a xor b);
    layer1_outputs(7342) <= a and not b;
    layer1_outputs(7343) <= a;
    layer1_outputs(7344) <= not (a xor b);
    layer1_outputs(7345) <= b;
    layer1_outputs(7346) <= 1'b0;
    layer1_outputs(7347) <= b and not a;
    layer1_outputs(7348) <= a;
    layer1_outputs(7349) <= not (a and b);
    layer1_outputs(7350) <= not (a or b);
    layer1_outputs(7351) <= b and not a;
    layer1_outputs(7352) <= b and not a;
    layer1_outputs(7353) <= not b or a;
    layer1_outputs(7354) <= a and not b;
    layer1_outputs(7355) <= not b;
    layer1_outputs(7356) <= not a;
    layer1_outputs(7357) <= not a;
    layer1_outputs(7358) <= a;
    layer1_outputs(7359) <= not b;
    layer1_outputs(7360) <= b and not a;
    layer1_outputs(7361) <= a and b;
    layer1_outputs(7362) <= b;
    layer1_outputs(7363) <= not (a or b);
    layer1_outputs(7364) <= a xor b;
    layer1_outputs(7365) <= not b;
    layer1_outputs(7366) <= not a;
    layer1_outputs(7367) <= not (a or b);
    layer1_outputs(7368) <= not b;
    layer1_outputs(7369) <= a xor b;
    layer1_outputs(7370) <= not a;
    layer1_outputs(7371) <= not a;
    layer1_outputs(7372) <= not (a and b);
    layer1_outputs(7373) <= not (a xor b);
    layer1_outputs(7374) <= not (a and b);
    layer1_outputs(7375) <= a;
    layer1_outputs(7376) <= a and not b;
    layer1_outputs(7377) <= a and not b;
    layer1_outputs(7378) <= not (a xor b);
    layer1_outputs(7379) <= not b;
    layer1_outputs(7380) <= not a;
    layer1_outputs(7381) <= not a;
    layer1_outputs(7382) <= b;
    layer1_outputs(7383) <= not b or a;
    layer1_outputs(7384) <= not a or b;
    layer1_outputs(7385) <= a;
    layer1_outputs(7386) <= 1'b0;
    layer1_outputs(7387) <= b and not a;
    layer1_outputs(7388) <= not (a xor b);
    layer1_outputs(7389) <= not b or a;
    layer1_outputs(7390) <= a or b;
    layer1_outputs(7391) <= b;
    layer1_outputs(7392) <= a and not b;
    layer1_outputs(7393) <= not a;
    layer1_outputs(7394) <= 1'b1;
    layer1_outputs(7395) <= a xor b;
    layer1_outputs(7396) <= not a or b;
    layer1_outputs(7397) <= not a;
    layer1_outputs(7398) <= a or b;
    layer1_outputs(7399) <= not a;
    layer1_outputs(7400) <= not b;
    layer1_outputs(7401) <= a and not b;
    layer1_outputs(7402) <= not (a and b);
    layer1_outputs(7403) <= not a;
    layer1_outputs(7404) <= not (a or b);
    layer1_outputs(7405) <= not (a and b);
    layer1_outputs(7406) <= not (a or b);
    layer1_outputs(7407) <= not (a or b);
    layer1_outputs(7408) <= a and not b;
    layer1_outputs(7409) <= a;
    layer1_outputs(7410) <= 1'b1;
    layer1_outputs(7411) <= not b or a;
    layer1_outputs(7412) <= not b or a;
    layer1_outputs(7413) <= not a or b;
    layer1_outputs(7414) <= a and not b;
    layer1_outputs(7415) <= a and b;
    layer1_outputs(7416) <= not (a and b);
    layer1_outputs(7417) <= a and not b;
    layer1_outputs(7418) <= b;
    layer1_outputs(7419) <= b and not a;
    layer1_outputs(7420) <= a or b;
    layer1_outputs(7421) <= a;
    layer1_outputs(7422) <= a xor b;
    layer1_outputs(7423) <= not b or a;
    layer1_outputs(7424) <= a or b;
    layer1_outputs(7425) <= 1'b0;
    layer1_outputs(7426) <= not b;
    layer1_outputs(7427) <= b;
    layer1_outputs(7428) <= a;
    layer1_outputs(7429) <= a and b;
    layer1_outputs(7430) <= not (a xor b);
    layer1_outputs(7431) <= a and b;
    layer1_outputs(7432) <= 1'b1;
    layer1_outputs(7433) <= not (a and b);
    layer1_outputs(7434) <= not (a or b);
    layer1_outputs(7435) <= a and not b;
    layer1_outputs(7436) <= not (a xor b);
    layer1_outputs(7437) <= not (a xor b);
    layer1_outputs(7438) <= b and not a;
    layer1_outputs(7439) <= not a;
    layer1_outputs(7440) <= not b or a;
    layer1_outputs(7441) <= a;
    layer1_outputs(7442) <= not a or b;
    layer1_outputs(7443) <= not b or a;
    layer1_outputs(7444) <= a xor b;
    layer1_outputs(7445) <= b;
    layer1_outputs(7446) <= not (a or b);
    layer1_outputs(7447) <= not b;
    layer1_outputs(7448) <= not b or a;
    layer1_outputs(7449) <= a or b;
    layer1_outputs(7450) <= a xor b;
    layer1_outputs(7451) <= not b;
    layer1_outputs(7452) <= a or b;
    layer1_outputs(7453) <= not (a and b);
    layer1_outputs(7454) <= a;
    layer1_outputs(7455) <= a;
    layer1_outputs(7456) <= not a;
    layer1_outputs(7457) <= 1'b1;
    layer1_outputs(7458) <= not (a xor b);
    layer1_outputs(7459) <= 1'b0;
    layer1_outputs(7460) <= a xor b;
    layer1_outputs(7461) <= not b;
    layer1_outputs(7462) <= not (a xor b);
    layer1_outputs(7463) <= not b;
    layer1_outputs(7464) <= a or b;
    layer1_outputs(7465) <= b and not a;
    layer1_outputs(7466) <= a or b;
    layer1_outputs(7467) <= a and b;
    layer1_outputs(7468) <= a and b;
    layer1_outputs(7469) <= not b;
    layer1_outputs(7470) <= a and b;
    layer1_outputs(7471) <= 1'b1;
    layer1_outputs(7472) <= not a or b;
    layer1_outputs(7473) <= b and not a;
    layer1_outputs(7474) <= a;
    layer1_outputs(7475) <= b;
    layer1_outputs(7476) <= a or b;
    layer1_outputs(7477) <= a and not b;
    layer1_outputs(7478) <= not a;
    layer1_outputs(7479) <= not a;
    layer1_outputs(7480) <= b;
    layer1_outputs(7481) <= not b or a;
    layer1_outputs(7482) <= not b;
    layer1_outputs(7483) <= not b;
    layer1_outputs(7484) <= b and not a;
    layer1_outputs(7485) <= b;
    layer1_outputs(7486) <= a and b;
    layer1_outputs(7487) <= b and not a;
    layer1_outputs(7488) <= a or b;
    layer1_outputs(7489) <= not b;
    layer1_outputs(7490) <= not a;
    layer1_outputs(7491) <= 1'b0;
    layer1_outputs(7492) <= a and not b;
    layer1_outputs(7493) <= b and not a;
    layer1_outputs(7494) <= a and b;
    layer1_outputs(7495) <= 1'b0;
    layer1_outputs(7496) <= not a or b;
    layer1_outputs(7497) <= not b or a;
    layer1_outputs(7498) <= a and not b;
    layer1_outputs(7499) <= not a;
    layer1_outputs(7500) <= a;
    layer1_outputs(7501) <= a xor b;
    layer1_outputs(7502) <= not a;
    layer1_outputs(7503) <= a and b;
    layer1_outputs(7504) <= not (a and b);
    layer1_outputs(7505) <= a and not b;
    layer1_outputs(7506) <= not (a and b);
    layer1_outputs(7507) <= not (a xor b);
    layer1_outputs(7508) <= b;
    layer1_outputs(7509) <= a or b;
    layer1_outputs(7510) <= a and b;
    layer1_outputs(7511) <= not (a and b);
    layer1_outputs(7512) <= not b or a;
    layer1_outputs(7513) <= a xor b;
    layer1_outputs(7514) <= not (a and b);
    layer1_outputs(7515) <= a xor b;
    layer1_outputs(7516) <= not (a and b);
    layer1_outputs(7517) <= a or b;
    layer1_outputs(7518) <= not a or b;
    layer1_outputs(7519) <= a;
    layer1_outputs(7520) <= not a;
    layer1_outputs(7521) <= not (a xor b);
    layer1_outputs(7522) <= not a;
    layer1_outputs(7523) <= a and not b;
    layer1_outputs(7524) <= not (a and b);
    layer1_outputs(7525) <= not a;
    layer1_outputs(7526) <= b;
    layer1_outputs(7527) <= a and not b;
    layer1_outputs(7528) <= not a or b;
    layer1_outputs(7529) <= b and not a;
    layer1_outputs(7530) <= not a;
    layer1_outputs(7531) <= not a;
    layer1_outputs(7532) <= not b;
    layer1_outputs(7533) <= not a;
    layer1_outputs(7534) <= a;
    layer1_outputs(7535) <= not b or a;
    layer1_outputs(7536) <= not b;
    layer1_outputs(7537) <= b;
    layer1_outputs(7538) <= not a;
    layer1_outputs(7539) <= b and not a;
    layer1_outputs(7540) <= not (a or b);
    layer1_outputs(7541) <= not a;
    layer1_outputs(7542) <= not a;
    layer1_outputs(7543) <= not b or a;
    layer1_outputs(7544) <= a and not b;
    layer1_outputs(7545) <= b;
    layer1_outputs(7546) <= a and b;
    layer1_outputs(7547) <= not b;
    layer1_outputs(7548) <= not (a xor b);
    layer1_outputs(7549) <= not (a or b);
    layer1_outputs(7550) <= not b;
    layer1_outputs(7551) <= a;
    layer1_outputs(7552) <= 1'b0;
    layer1_outputs(7553) <= not b or a;
    layer1_outputs(7554) <= not (a and b);
    layer1_outputs(7555) <= a and b;
    layer1_outputs(7556) <= 1'b0;
    layer1_outputs(7557) <= a or b;
    layer1_outputs(7558) <= a and not b;
    layer1_outputs(7559) <= b;
    layer1_outputs(7560) <= a;
    layer1_outputs(7561) <= a and b;
    layer1_outputs(7562) <= a and b;
    layer1_outputs(7563) <= not b;
    layer1_outputs(7564) <= a xor b;
    layer1_outputs(7565) <= a xor b;
    layer1_outputs(7566) <= not b;
    layer1_outputs(7567) <= b;
    layer1_outputs(7568) <= not b or a;
    layer1_outputs(7569) <= not a or b;
    layer1_outputs(7570) <= b;
    layer1_outputs(7571) <= b;
    layer1_outputs(7572) <= b and not a;
    layer1_outputs(7573) <= a or b;
    layer1_outputs(7574) <= not b or a;
    layer1_outputs(7575) <= a;
    layer1_outputs(7576) <= not (a or b);
    layer1_outputs(7577) <= a;
    layer1_outputs(7578) <= a;
    layer1_outputs(7579) <= not (a xor b);
    layer1_outputs(7580) <= not (a or b);
    layer1_outputs(7581) <= a xor b;
    layer1_outputs(7582) <= a;
    layer1_outputs(7583) <= b and not a;
    layer1_outputs(7584) <= a or b;
    layer1_outputs(7585) <= not (a or b);
    layer1_outputs(7586) <= not b;
    layer1_outputs(7587) <= not b or a;
    layer1_outputs(7588) <= 1'b1;
    layer1_outputs(7589) <= a xor b;
    layer1_outputs(7590) <= a and not b;
    layer1_outputs(7591) <= a xor b;
    layer1_outputs(7592) <= not b;
    layer1_outputs(7593) <= not a;
    layer1_outputs(7594) <= not a;
    layer1_outputs(7595) <= a and b;
    layer1_outputs(7596) <= not (a and b);
    layer1_outputs(7597) <= a and not b;
    layer1_outputs(7598) <= a and not b;
    layer1_outputs(7599) <= not a;
    layer1_outputs(7600) <= a and b;
    layer1_outputs(7601) <= not b;
    layer1_outputs(7602) <= a xor b;
    layer1_outputs(7603) <= a or b;
    layer1_outputs(7604) <= a or b;
    layer1_outputs(7605) <= b and not a;
    layer1_outputs(7606) <= a and b;
    layer1_outputs(7607) <= a xor b;
    layer1_outputs(7608) <= b;
    layer1_outputs(7609) <= a;
    layer1_outputs(7610) <= not (a and b);
    layer1_outputs(7611) <= a;
    layer1_outputs(7612) <= b and not a;
    layer1_outputs(7613) <= not (a xor b);
    layer1_outputs(7614) <= not b;
    layer1_outputs(7615) <= a;
    layer1_outputs(7616) <= 1'b1;
    layer1_outputs(7617) <= not (a xor b);
    layer1_outputs(7618) <= b and not a;
    layer1_outputs(7619) <= a and b;
    layer1_outputs(7620) <= not a;
    layer1_outputs(7621) <= 1'b1;
    layer1_outputs(7622) <= b;
    layer1_outputs(7623) <= not (a and b);
    layer1_outputs(7624) <= not (a or b);
    layer1_outputs(7625) <= not a or b;
    layer1_outputs(7626) <= a;
    layer1_outputs(7627) <= b and not a;
    layer1_outputs(7628) <= not b;
    layer1_outputs(7629) <= not (a xor b);
    layer1_outputs(7630) <= a or b;
    layer1_outputs(7631) <= a and not b;
    layer1_outputs(7632) <= not (a or b);
    layer1_outputs(7633) <= b and not a;
    layer1_outputs(7634) <= b and not a;
    layer1_outputs(7635) <= 1'b0;
    layer1_outputs(7636) <= b and not a;
    layer1_outputs(7637) <= a xor b;
    layer1_outputs(7638) <= a xor b;
    layer1_outputs(7639) <= not (a or b);
    layer1_outputs(7640) <= a xor b;
    layer1_outputs(7641) <= b and not a;
    layer1_outputs(7642) <= not a or b;
    layer1_outputs(7643) <= not (a xor b);
    layer1_outputs(7644) <= not (a xor b);
    layer1_outputs(7645) <= not (a or b);
    layer1_outputs(7646) <= a;
    layer1_outputs(7647) <= not (a or b);
    layer1_outputs(7648) <= b;
    layer1_outputs(7649) <= a and not b;
    layer1_outputs(7650) <= b;
    layer1_outputs(7651) <= b;
    layer1_outputs(7652) <= not (a or b);
    layer1_outputs(7653) <= not (a or b);
    layer1_outputs(7654) <= not b or a;
    layer1_outputs(7655) <= a xor b;
    layer1_outputs(7656) <= b;
    layer1_outputs(7657) <= not b or a;
    layer1_outputs(7658) <= not (a or b);
    layer1_outputs(7659) <= 1'b1;
    layer1_outputs(7660) <= a and not b;
    layer1_outputs(7661) <= not a or b;
    layer1_outputs(7662) <= b and not a;
    layer1_outputs(7663) <= not a;
    layer1_outputs(7664) <= not b or a;
    layer1_outputs(7665) <= a xor b;
    layer1_outputs(7666) <= not a or b;
    layer1_outputs(7667) <= a xor b;
    layer1_outputs(7668) <= not a;
    layer1_outputs(7669) <= not (a or b);
    layer1_outputs(7670) <= not b or a;
    layer1_outputs(7671) <= a or b;
    layer1_outputs(7672) <= b and not a;
    layer1_outputs(7673) <= not (a or b);
    layer1_outputs(7674) <= a or b;
    layer1_outputs(7675) <= not a or b;
    layer1_outputs(7676) <= a;
    layer1_outputs(7677) <= not a;
    layer1_outputs(7678) <= not (a or b);
    layer1_outputs(7679) <= a;
    layer2_outputs(0) <= not (a or b);
    layer2_outputs(1) <= b;
    layer2_outputs(2) <= not b;
    layer2_outputs(3) <= not (a xor b);
    layer2_outputs(4) <= a or b;
    layer2_outputs(5) <= not a or b;
    layer2_outputs(6) <= a;
    layer2_outputs(7) <= a and not b;
    layer2_outputs(8) <= not (a xor b);
    layer2_outputs(9) <= not b;
    layer2_outputs(10) <= not (a xor b);
    layer2_outputs(11) <= b and not a;
    layer2_outputs(12) <= not a;
    layer2_outputs(13) <= not (a xor b);
    layer2_outputs(14) <= a and not b;
    layer2_outputs(15) <= not (a or b);
    layer2_outputs(16) <= not (a xor b);
    layer2_outputs(17) <= b and not a;
    layer2_outputs(18) <= not (a or b);
    layer2_outputs(19) <= not (a and b);
    layer2_outputs(20) <= 1'b1;
    layer2_outputs(21) <= a;
    layer2_outputs(22) <= b and not a;
    layer2_outputs(23) <= a xor b;
    layer2_outputs(24) <= not b;
    layer2_outputs(25) <= not a or b;
    layer2_outputs(26) <= not (a or b);
    layer2_outputs(27) <= a and b;
    layer2_outputs(28) <= not a;
    layer2_outputs(29) <= a or b;
    layer2_outputs(30) <= b;
    layer2_outputs(31) <= a and not b;
    layer2_outputs(32) <= a xor b;
    layer2_outputs(33) <= not a;
    layer2_outputs(34) <= a and not b;
    layer2_outputs(35) <= not b;
    layer2_outputs(36) <= a;
    layer2_outputs(37) <= a or b;
    layer2_outputs(38) <= not (a or b);
    layer2_outputs(39) <= b;
    layer2_outputs(40) <= not (a and b);
    layer2_outputs(41) <= a or b;
    layer2_outputs(42) <= not (a xor b);
    layer2_outputs(43) <= a xor b;
    layer2_outputs(44) <= not b or a;
    layer2_outputs(45) <= a;
    layer2_outputs(46) <= b and not a;
    layer2_outputs(47) <= b and not a;
    layer2_outputs(48) <= a or b;
    layer2_outputs(49) <= not (a xor b);
    layer2_outputs(50) <= b and not a;
    layer2_outputs(51) <= b;
    layer2_outputs(52) <= not (a or b);
    layer2_outputs(53) <= a and b;
    layer2_outputs(54) <= not (a xor b);
    layer2_outputs(55) <= not a or b;
    layer2_outputs(56) <= not (a xor b);
    layer2_outputs(57) <= a;
    layer2_outputs(58) <= not a;
    layer2_outputs(59) <= not a;
    layer2_outputs(60) <= not b;
    layer2_outputs(61) <= not a;
    layer2_outputs(62) <= not a or b;
    layer2_outputs(63) <= not (a and b);
    layer2_outputs(64) <= b;
    layer2_outputs(65) <= a and not b;
    layer2_outputs(66) <= a xor b;
    layer2_outputs(67) <= not a or b;
    layer2_outputs(68) <= a;
    layer2_outputs(69) <= a xor b;
    layer2_outputs(70) <= not (a xor b);
    layer2_outputs(71) <= not (a and b);
    layer2_outputs(72) <= not (a or b);
    layer2_outputs(73) <= not (a xor b);
    layer2_outputs(74) <= not b;
    layer2_outputs(75) <= not b or a;
    layer2_outputs(76) <= b and not a;
    layer2_outputs(77) <= b;
    layer2_outputs(78) <= a xor b;
    layer2_outputs(79) <= a or b;
    layer2_outputs(80) <= a and b;
    layer2_outputs(81) <= a;
    layer2_outputs(82) <= not b;
    layer2_outputs(83) <= not (a xor b);
    layer2_outputs(84) <= a;
    layer2_outputs(85) <= a or b;
    layer2_outputs(86) <= a or b;
    layer2_outputs(87) <= not (a xor b);
    layer2_outputs(88) <= not b;
    layer2_outputs(89) <= a;
    layer2_outputs(90) <= a or b;
    layer2_outputs(91) <= a or b;
    layer2_outputs(92) <= not a or b;
    layer2_outputs(93) <= not a;
    layer2_outputs(94) <= a and b;
    layer2_outputs(95) <= not a;
    layer2_outputs(96) <= not (a or b);
    layer2_outputs(97) <= not a or b;
    layer2_outputs(98) <= a and b;
    layer2_outputs(99) <= b and not a;
    layer2_outputs(100) <= not b;
    layer2_outputs(101) <= not b or a;
    layer2_outputs(102) <= not (a and b);
    layer2_outputs(103) <= not b;
    layer2_outputs(104) <= not b;
    layer2_outputs(105) <= not a;
    layer2_outputs(106) <= not (a xor b);
    layer2_outputs(107) <= a;
    layer2_outputs(108) <= b;
    layer2_outputs(109) <= b;
    layer2_outputs(110) <= a xor b;
    layer2_outputs(111) <= a;
    layer2_outputs(112) <= b;
    layer2_outputs(113) <= not a;
    layer2_outputs(114) <= b;
    layer2_outputs(115) <= not b;
    layer2_outputs(116) <= not b;
    layer2_outputs(117) <= a and not b;
    layer2_outputs(118) <= a and not b;
    layer2_outputs(119) <= a xor b;
    layer2_outputs(120) <= a;
    layer2_outputs(121) <= not a;
    layer2_outputs(122) <= a;
    layer2_outputs(123) <= a or b;
    layer2_outputs(124) <= a;
    layer2_outputs(125) <= not a;
    layer2_outputs(126) <= not a or b;
    layer2_outputs(127) <= b;
    layer2_outputs(128) <= a;
    layer2_outputs(129) <= a xor b;
    layer2_outputs(130) <= a xor b;
    layer2_outputs(131) <= b;
    layer2_outputs(132) <= not b or a;
    layer2_outputs(133) <= b;
    layer2_outputs(134) <= not b or a;
    layer2_outputs(135) <= a;
    layer2_outputs(136) <= not a;
    layer2_outputs(137) <= not b;
    layer2_outputs(138) <= not b;
    layer2_outputs(139) <= not (a or b);
    layer2_outputs(140) <= b and not a;
    layer2_outputs(141) <= a and b;
    layer2_outputs(142) <= a or b;
    layer2_outputs(143) <= b and not a;
    layer2_outputs(144) <= not (a and b);
    layer2_outputs(145) <= a;
    layer2_outputs(146) <= a and b;
    layer2_outputs(147) <= not (a xor b);
    layer2_outputs(148) <= a or b;
    layer2_outputs(149) <= b;
    layer2_outputs(150) <= not b;
    layer2_outputs(151) <= b;
    layer2_outputs(152) <= not (a or b);
    layer2_outputs(153) <= a and b;
    layer2_outputs(154) <= a xor b;
    layer2_outputs(155) <= not a;
    layer2_outputs(156) <= a;
    layer2_outputs(157) <= not a or b;
    layer2_outputs(158) <= not (a or b);
    layer2_outputs(159) <= b;
    layer2_outputs(160) <= not a;
    layer2_outputs(161) <= not b;
    layer2_outputs(162) <= a;
    layer2_outputs(163) <= not a or b;
    layer2_outputs(164) <= not b;
    layer2_outputs(165) <= not a;
    layer2_outputs(166) <= not (a or b);
    layer2_outputs(167) <= not b;
    layer2_outputs(168) <= a xor b;
    layer2_outputs(169) <= a and b;
    layer2_outputs(170) <= not b;
    layer2_outputs(171) <= a;
    layer2_outputs(172) <= a or b;
    layer2_outputs(173) <= not a;
    layer2_outputs(174) <= a or b;
    layer2_outputs(175) <= a and not b;
    layer2_outputs(176) <= not b or a;
    layer2_outputs(177) <= a;
    layer2_outputs(178) <= not (a or b);
    layer2_outputs(179) <= not a or b;
    layer2_outputs(180) <= a;
    layer2_outputs(181) <= not b or a;
    layer2_outputs(182) <= a;
    layer2_outputs(183) <= not (a xor b);
    layer2_outputs(184) <= a;
    layer2_outputs(185) <= not b;
    layer2_outputs(186) <= b;
    layer2_outputs(187) <= not a;
    layer2_outputs(188) <= 1'b1;
    layer2_outputs(189) <= not b;
    layer2_outputs(190) <= a xor b;
    layer2_outputs(191) <= b and not a;
    layer2_outputs(192) <= not a or b;
    layer2_outputs(193) <= b;
    layer2_outputs(194) <= a;
    layer2_outputs(195) <= a and not b;
    layer2_outputs(196) <= b;
    layer2_outputs(197) <= not a;
    layer2_outputs(198) <= a and b;
    layer2_outputs(199) <= not a;
    layer2_outputs(200) <= not (a or b);
    layer2_outputs(201) <= a and not b;
    layer2_outputs(202) <= not b or a;
    layer2_outputs(203) <= a and b;
    layer2_outputs(204) <= not (a xor b);
    layer2_outputs(205) <= b;
    layer2_outputs(206) <= a or b;
    layer2_outputs(207) <= a;
    layer2_outputs(208) <= a xor b;
    layer2_outputs(209) <= a;
    layer2_outputs(210) <= a;
    layer2_outputs(211) <= not (a xor b);
    layer2_outputs(212) <= a;
    layer2_outputs(213) <= a or b;
    layer2_outputs(214) <= b;
    layer2_outputs(215) <= a;
    layer2_outputs(216) <= b;
    layer2_outputs(217) <= not (a and b);
    layer2_outputs(218) <= not (a or b);
    layer2_outputs(219) <= not b or a;
    layer2_outputs(220) <= a and not b;
    layer2_outputs(221) <= a xor b;
    layer2_outputs(222) <= not (a xor b);
    layer2_outputs(223) <= not a or b;
    layer2_outputs(224) <= not (a xor b);
    layer2_outputs(225) <= a or b;
    layer2_outputs(226) <= not (a and b);
    layer2_outputs(227) <= b and not a;
    layer2_outputs(228) <= a or b;
    layer2_outputs(229) <= not (a xor b);
    layer2_outputs(230) <= not (a and b);
    layer2_outputs(231) <= not b;
    layer2_outputs(232) <= not (a and b);
    layer2_outputs(233) <= a and b;
    layer2_outputs(234) <= not (a and b);
    layer2_outputs(235) <= not b;
    layer2_outputs(236) <= not (a and b);
    layer2_outputs(237) <= not b;
    layer2_outputs(238) <= not a;
    layer2_outputs(239) <= not (a xor b);
    layer2_outputs(240) <= not a;
    layer2_outputs(241) <= b and not a;
    layer2_outputs(242) <= not a;
    layer2_outputs(243) <= b;
    layer2_outputs(244) <= b;
    layer2_outputs(245) <= a or b;
    layer2_outputs(246) <= a and not b;
    layer2_outputs(247) <= a and b;
    layer2_outputs(248) <= a;
    layer2_outputs(249) <= 1'b1;
    layer2_outputs(250) <= not b;
    layer2_outputs(251) <= b;
    layer2_outputs(252) <= not (a or b);
    layer2_outputs(253) <= a or b;
    layer2_outputs(254) <= a xor b;
    layer2_outputs(255) <= b and not a;
    layer2_outputs(256) <= not a or b;
    layer2_outputs(257) <= not (a xor b);
    layer2_outputs(258) <= not b;
    layer2_outputs(259) <= not b or a;
    layer2_outputs(260) <= not b;
    layer2_outputs(261) <= a xor b;
    layer2_outputs(262) <= a xor b;
    layer2_outputs(263) <= not b;
    layer2_outputs(264) <= not b;
    layer2_outputs(265) <= a and b;
    layer2_outputs(266) <= not b or a;
    layer2_outputs(267) <= not (a and b);
    layer2_outputs(268) <= not b or a;
    layer2_outputs(269) <= a and not b;
    layer2_outputs(270) <= not (a xor b);
    layer2_outputs(271) <= a xor b;
    layer2_outputs(272) <= a xor b;
    layer2_outputs(273) <= not (a and b);
    layer2_outputs(274) <= not a;
    layer2_outputs(275) <= not (a and b);
    layer2_outputs(276) <= a;
    layer2_outputs(277) <= a;
    layer2_outputs(278) <= b;
    layer2_outputs(279) <= not a;
    layer2_outputs(280) <= not b;
    layer2_outputs(281) <= a and b;
    layer2_outputs(282) <= not b;
    layer2_outputs(283) <= a;
    layer2_outputs(284) <= not a;
    layer2_outputs(285) <= not b;
    layer2_outputs(286) <= a xor b;
    layer2_outputs(287) <= not b or a;
    layer2_outputs(288) <= not (a and b);
    layer2_outputs(289) <= not b or a;
    layer2_outputs(290) <= not (a xor b);
    layer2_outputs(291) <= a xor b;
    layer2_outputs(292) <= a;
    layer2_outputs(293) <= a;
    layer2_outputs(294) <= b and not a;
    layer2_outputs(295) <= a and not b;
    layer2_outputs(296) <= not (a and b);
    layer2_outputs(297) <= a;
    layer2_outputs(298) <= not (a or b);
    layer2_outputs(299) <= not a;
    layer2_outputs(300) <= a;
    layer2_outputs(301) <= a;
    layer2_outputs(302) <= b;
    layer2_outputs(303) <= b;
    layer2_outputs(304) <= a and b;
    layer2_outputs(305) <= a;
    layer2_outputs(306) <= not (a xor b);
    layer2_outputs(307) <= a;
    layer2_outputs(308) <= not a;
    layer2_outputs(309) <= not b;
    layer2_outputs(310) <= a or b;
    layer2_outputs(311) <= not (a and b);
    layer2_outputs(312) <= not a or b;
    layer2_outputs(313) <= not b;
    layer2_outputs(314) <= b;
    layer2_outputs(315) <= a;
    layer2_outputs(316) <= a;
    layer2_outputs(317) <= not b;
    layer2_outputs(318) <= b and not a;
    layer2_outputs(319) <= not a or b;
    layer2_outputs(320) <= b;
    layer2_outputs(321) <= a xor b;
    layer2_outputs(322) <= a and not b;
    layer2_outputs(323) <= a xor b;
    layer2_outputs(324) <= a;
    layer2_outputs(325) <= not (a xor b);
    layer2_outputs(326) <= not b;
    layer2_outputs(327) <= not (a and b);
    layer2_outputs(328) <= not a;
    layer2_outputs(329) <= not a;
    layer2_outputs(330) <= not (a and b);
    layer2_outputs(331) <= not b or a;
    layer2_outputs(332) <= b and not a;
    layer2_outputs(333) <= a xor b;
    layer2_outputs(334) <= not b;
    layer2_outputs(335) <= not a or b;
    layer2_outputs(336) <= not a;
    layer2_outputs(337) <= a and b;
    layer2_outputs(338) <= not (a or b);
    layer2_outputs(339) <= not b;
    layer2_outputs(340) <= not b or a;
    layer2_outputs(341) <= not a;
    layer2_outputs(342) <= not (a and b);
    layer2_outputs(343) <= a and b;
    layer2_outputs(344) <= b;
    layer2_outputs(345) <= not a or b;
    layer2_outputs(346) <= a;
    layer2_outputs(347) <= a and b;
    layer2_outputs(348) <= not a or b;
    layer2_outputs(349) <= b and not a;
    layer2_outputs(350) <= not a;
    layer2_outputs(351) <= a and not b;
    layer2_outputs(352) <= a or b;
    layer2_outputs(353) <= a xor b;
    layer2_outputs(354) <= a and not b;
    layer2_outputs(355) <= a and b;
    layer2_outputs(356) <= not a or b;
    layer2_outputs(357) <= not b;
    layer2_outputs(358) <= not (a or b);
    layer2_outputs(359) <= a and b;
    layer2_outputs(360) <= not b;
    layer2_outputs(361) <= a and not b;
    layer2_outputs(362) <= not b or a;
    layer2_outputs(363) <= a and b;
    layer2_outputs(364) <= not a or b;
    layer2_outputs(365) <= b;
    layer2_outputs(366) <= not a or b;
    layer2_outputs(367) <= not a;
    layer2_outputs(368) <= a xor b;
    layer2_outputs(369) <= a and b;
    layer2_outputs(370) <= not a;
    layer2_outputs(371) <= b;
    layer2_outputs(372) <= not (a and b);
    layer2_outputs(373) <= not a;
    layer2_outputs(374) <= a and b;
    layer2_outputs(375) <= b;
    layer2_outputs(376) <= b;
    layer2_outputs(377) <= 1'b1;
    layer2_outputs(378) <= a and not b;
    layer2_outputs(379) <= a xor b;
    layer2_outputs(380) <= not b;
    layer2_outputs(381) <= not (a xor b);
    layer2_outputs(382) <= a;
    layer2_outputs(383) <= a xor b;
    layer2_outputs(384) <= a xor b;
    layer2_outputs(385) <= not b or a;
    layer2_outputs(386) <= not (a and b);
    layer2_outputs(387) <= not a;
    layer2_outputs(388) <= not (a xor b);
    layer2_outputs(389) <= not (a xor b);
    layer2_outputs(390) <= not b;
    layer2_outputs(391) <= not b;
    layer2_outputs(392) <= not (a and b);
    layer2_outputs(393) <= not b;
    layer2_outputs(394) <= a xor b;
    layer2_outputs(395) <= not (a or b);
    layer2_outputs(396) <= not (a xor b);
    layer2_outputs(397) <= b;
    layer2_outputs(398) <= not a or b;
    layer2_outputs(399) <= a xor b;
    layer2_outputs(400) <= b and not a;
    layer2_outputs(401) <= not b or a;
    layer2_outputs(402) <= a xor b;
    layer2_outputs(403) <= a and not b;
    layer2_outputs(404) <= b and not a;
    layer2_outputs(405) <= a xor b;
    layer2_outputs(406) <= not a;
    layer2_outputs(407) <= not b;
    layer2_outputs(408) <= not (a xor b);
    layer2_outputs(409) <= a and b;
    layer2_outputs(410) <= not a or b;
    layer2_outputs(411) <= not (a and b);
    layer2_outputs(412) <= not b;
    layer2_outputs(413) <= not b or a;
    layer2_outputs(414) <= a and b;
    layer2_outputs(415) <= a xor b;
    layer2_outputs(416) <= not (a or b);
    layer2_outputs(417) <= not b;
    layer2_outputs(418) <= b;
    layer2_outputs(419) <= not b;
    layer2_outputs(420) <= b;
    layer2_outputs(421) <= not b;
    layer2_outputs(422) <= not a;
    layer2_outputs(423) <= not (a and b);
    layer2_outputs(424) <= not (a xor b);
    layer2_outputs(425) <= not a;
    layer2_outputs(426) <= not (a and b);
    layer2_outputs(427) <= not (a xor b);
    layer2_outputs(428) <= not b;
    layer2_outputs(429) <= a;
    layer2_outputs(430) <= not a or b;
    layer2_outputs(431) <= not b;
    layer2_outputs(432) <= a;
    layer2_outputs(433) <= not (a or b);
    layer2_outputs(434) <= a;
    layer2_outputs(435) <= not b or a;
    layer2_outputs(436) <= not b;
    layer2_outputs(437) <= a and b;
    layer2_outputs(438) <= not a or b;
    layer2_outputs(439) <= not (a xor b);
    layer2_outputs(440) <= a;
    layer2_outputs(441) <= not a;
    layer2_outputs(442) <= a;
    layer2_outputs(443) <= a xor b;
    layer2_outputs(444) <= not (a xor b);
    layer2_outputs(445) <= a and not b;
    layer2_outputs(446) <= not (a xor b);
    layer2_outputs(447) <= a;
    layer2_outputs(448) <= a xor b;
    layer2_outputs(449) <= not (a or b);
    layer2_outputs(450) <= b;
    layer2_outputs(451) <= a xor b;
    layer2_outputs(452) <= b;
    layer2_outputs(453) <= not (a or b);
    layer2_outputs(454) <= not a or b;
    layer2_outputs(455) <= a and b;
    layer2_outputs(456) <= a;
    layer2_outputs(457) <= b;
    layer2_outputs(458) <= a and b;
    layer2_outputs(459) <= not b;
    layer2_outputs(460) <= not a;
    layer2_outputs(461) <= not a;
    layer2_outputs(462) <= not (a or b);
    layer2_outputs(463) <= a;
    layer2_outputs(464) <= a and b;
    layer2_outputs(465) <= not a or b;
    layer2_outputs(466) <= a and b;
    layer2_outputs(467) <= a;
    layer2_outputs(468) <= b;
    layer2_outputs(469) <= not (a xor b);
    layer2_outputs(470) <= a;
    layer2_outputs(471) <= a xor b;
    layer2_outputs(472) <= a;
    layer2_outputs(473) <= b and not a;
    layer2_outputs(474) <= not b;
    layer2_outputs(475) <= not (a and b);
    layer2_outputs(476) <= not (a and b);
    layer2_outputs(477) <= not a or b;
    layer2_outputs(478) <= not a;
    layer2_outputs(479) <= not b or a;
    layer2_outputs(480) <= not (a and b);
    layer2_outputs(481) <= not (a or b);
    layer2_outputs(482) <= b;
    layer2_outputs(483) <= not b;
    layer2_outputs(484) <= not a;
    layer2_outputs(485) <= a and b;
    layer2_outputs(486) <= a and b;
    layer2_outputs(487) <= a and not b;
    layer2_outputs(488) <= not (a xor b);
    layer2_outputs(489) <= not b;
    layer2_outputs(490) <= a or b;
    layer2_outputs(491) <= not (a or b);
    layer2_outputs(492) <= a;
    layer2_outputs(493) <= not (a and b);
    layer2_outputs(494) <= a and b;
    layer2_outputs(495) <= 1'b1;
    layer2_outputs(496) <= not a or b;
    layer2_outputs(497) <= not a;
    layer2_outputs(498) <= not a;
    layer2_outputs(499) <= not a;
    layer2_outputs(500) <= not a;
    layer2_outputs(501) <= not b;
    layer2_outputs(502) <= not b;
    layer2_outputs(503) <= not b;
    layer2_outputs(504) <= b;
    layer2_outputs(505) <= a and not b;
    layer2_outputs(506) <= a;
    layer2_outputs(507) <= 1'b0;
    layer2_outputs(508) <= b;
    layer2_outputs(509) <= b;
    layer2_outputs(510) <= a and not b;
    layer2_outputs(511) <= a or b;
    layer2_outputs(512) <= not b;
    layer2_outputs(513) <= not (a or b);
    layer2_outputs(514) <= a and not b;
    layer2_outputs(515) <= not (a or b);
    layer2_outputs(516) <= not (a or b);
    layer2_outputs(517) <= b;
    layer2_outputs(518) <= not a;
    layer2_outputs(519) <= a and not b;
    layer2_outputs(520) <= a xor b;
    layer2_outputs(521) <= not a or b;
    layer2_outputs(522) <= a and not b;
    layer2_outputs(523) <= not (a and b);
    layer2_outputs(524) <= not b;
    layer2_outputs(525) <= a or b;
    layer2_outputs(526) <= not (a xor b);
    layer2_outputs(527) <= not a or b;
    layer2_outputs(528) <= a and not b;
    layer2_outputs(529) <= not a;
    layer2_outputs(530) <= a xor b;
    layer2_outputs(531) <= b;
    layer2_outputs(532) <= not (a xor b);
    layer2_outputs(533) <= not (a xor b);
    layer2_outputs(534) <= a xor b;
    layer2_outputs(535) <= not a or b;
    layer2_outputs(536) <= a and b;
    layer2_outputs(537) <= a xor b;
    layer2_outputs(538) <= a and b;
    layer2_outputs(539) <= b;
    layer2_outputs(540) <= a;
    layer2_outputs(541) <= not a;
    layer2_outputs(542) <= not (a or b);
    layer2_outputs(543) <= b;
    layer2_outputs(544) <= not (a and b);
    layer2_outputs(545) <= b;
    layer2_outputs(546) <= not b or a;
    layer2_outputs(547) <= a;
    layer2_outputs(548) <= not (a and b);
    layer2_outputs(549) <= not b or a;
    layer2_outputs(550) <= a;
    layer2_outputs(551) <= a or b;
    layer2_outputs(552) <= a xor b;
    layer2_outputs(553) <= a;
    layer2_outputs(554) <= not b;
    layer2_outputs(555) <= b;
    layer2_outputs(556) <= not (a xor b);
    layer2_outputs(557) <= a xor b;
    layer2_outputs(558) <= a and not b;
    layer2_outputs(559) <= a;
    layer2_outputs(560) <= not a;
    layer2_outputs(561) <= a;
    layer2_outputs(562) <= not b;
    layer2_outputs(563) <= a;
    layer2_outputs(564) <= not a or b;
    layer2_outputs(565) <= not a or b;
    layer2_outputs(566) <= a xor b;
    layer2_outputs(567) <= not (a xor b);
    layer2_outputs(568) <= not (a and b);
    layer2_outputs(569) <= not a or b;
    layer2_outputs(570) <= b;
    layer2_outputs(571) <= b;
    layer2_outputs(572) <= a xor b;
    layer2_outputs(573) <= not (a or b);
    layer2_outputs(574) <= b and not a;
    layer2_outputs(575) <= not (a and b);
    layer2_outputs(576) <= a;
    layer2_outputs(577) <= not a;
    layer2_outputs(578) <= not (a and b);
    layer2_outputs(579) <= not a or b;
    layer2_outputs(580) <= not a;
    layer2_outputs(581) <= a and b;
    layer2_outputs(582) <= b;
    layer2_outputs(583) <= a;
    layer2_outputs(584) <= a and not b;
    layer2_outputs(585) <= not b;
    layer2_outputs(586) <= not a;
    layer2_outputs(587) <= not b;
    layer2_outputs(588) <= not b;
    layer2_outputs(589) <= a and b;
    layer2_outputs(590) <= not b or a;
    layer2_outputs(591) <= not a;
    layer2_outputs(592) <= not b;
    layer2_outputs(593) <= b and not a;
    layer2_outputs(594) <= a;
    layer2_outputs(595) <= a or b;
    layer2_outputs(596) <= a;
    layer2_outputs(597) <= not (a xor b);
    layer2_outputs(598) <= not b;
    layer2_outputs(599) <= a;
    layer2_outputs(600) <= a or b;
    layer2_outputs(601) <= a or b;
    layer2_outputs(602) <= not (a and b);
    layer2_outputs(603) <= not (a or b);
    layer2_outputs(604) <= not (a xor b);
    layer2_outputs(605) <= a;
    layer2_outputs(606) <= a and not b;
    layer2_outputs(607) <= b;
    layer2_outputs(608) <= not (a xor b);
    layer2_outputs(609) <= not b;
    layer2_outputs(610) <= b;
    layer2_outputs(611) <= a;
    layer2_outputs(612) <= b;
    layer2_outputs(613) <= not b;
    layer2_outputs(614) <= a xor b;
    layer2_outputs(615) <= b;
    layer2_outputs(616) <= a;
    layer2_outputs(617) <= not (a or b);
    layer2_outputs(618) <= not (a and b);
    layer2_outputs(619) <= not (a or b);
    layer2_outputs(620) <= not (a or b);
    layer2_outputs(621) <= a;
    layer2_outputs(622) <= b;
    layer2_outputs(623) <= not a;
    layer2_outputs(624) <= not (a or b);
    layer2_outputs(625) <= a;
    layer2_outputs(626) <= not a or b;
    layer2_outputs(627) <= not b or a;
    layer2_outputs(628) <= not b;
    layer2_outputs(629) <= a xor b;
    layer2_outputs(630) <= not b;
    layer2_outputs(631) <= a;
    layer2_outputs(632) <= a and not b;
    layer2_outputs(633) <= not b or a;
    layer2_outputs(634) <= not a or b;
    layer2_outputs(635) <= 1'b1;
    layer2_outputs(636) <= not (a and b);
    layer2_outputs(637) <= not (a xor b);
    layer2_outputs(638) <= not b;
    layer2_outputs(639) <= a xor b;
    layer2_outputs(640) <= a;
    layer2_outputs(641) <= a;
    layer2_outputs(642) <= not (a or b);
    layer2_outputs(643) <= not a;
    layer2_outputs(644) <= not (a or b);
    layer2_outputs(645) <= not a;
    layer2_outputs(646) <= b;
    layer2_outputs(647) <= a;
    layer2_outputs(648) <= b and not a;
    layer2_outputs(649) <= not b;
    layer2_outputs(650) <= not b or a;
    layer2_outputs(651) <= a and not b;
    layer2_outputs(652) <= a and not b;
    layer2_outputs(653) <= not (a or b);
    layer2_outputs(654) <= a or b;
    layer2_outputs(655) <= not (a or b);
    layer2_outputs(656) <= not b;
    layer2_outputs(657) <= b;
    layer2_outputs(658) <= a;
    layer2_outputs(659) <= a;
    layer2_outputs(660) <= a and not b;
    layer2_outputs(661) <= not a;
    layer2_outputs(662) <= not a;
    layer2_outputs(663) <= a xor b;
    layer2_outputs(664) <= a xor b;
    layer2_outputs(665) <= not (a or b);
    layer2_outputs(666) <= a or b;
    layer2_outputs(667) <= not a;
    layer2_outputs(668) <= not b or a;
    layer2_outputs(669) <= not (a and b);
    layer2_outputs(670) <= a;
    layer2_outputs(671) <= b and not a;
    layer2_outputs(672) <= a;
    layer2_outputs(673) <= a;
    layer2_outputs(674) <= a;
    layer2_outputs(675) <= b and not a;
    layer2_outputs(676) <= a or b;
    layer2_outputs(677) <= a and not b;
    layer2_outputs(678) <= a and not b;
    layer2_outputs(679) <= a or b;
    layer2_outputs(680) <= 1'b1;
    layer2_outputs(681) <= not b or a;
    layer2_outputs(682) <= not a;
    layer2_outputs(683) <= a xor b;
    layer2_outputs(684) <= a and b;
    layer2_outputs(685) <= b and not a;
    layer2_outputs(686) <= b and not a;
    layer2_outputs(687) <= not (a and b);
    layer2_outputs(688) <= a xor b;
    layer2_outputs(689) <= a and not b;
    layer2_outputs(690) <= a or b;
    layer2_outputs(691) <= not a or b;
    layer2_outputs(692) <= not a;
    layer2_outputs(693) <= a and not b;
    layer2_outputs(694) <= not (a or b);
    layer2_outputs(695) <= not (a xor b);
    layer2_outputs(696) <= 1'b0;
    layer2_outputs(697) <= not b;
    layer2_outputs(698) <= a or b;
    layer2_outputs(699) <= not a;
    layer2_outputs(700) <= not a or b;
    layer2_outputs(701) <= a;
    layer2_outputs(702) <= not b;
    layer2_outputs(703) <= not b;
    layer2_outputs(704) <= not b;
    layer2_outputs(705) <= a and b;
    layer2_outputs(706) <= a xor b;
    layer2_outputs(707) <= not b or a;
    layer2_outputs(708) <= not b;
    layer2_outputs(709) <= a or b;
    layer2_outputs(710) <= not (a xor b);
    layer2_outputs(711) <= a and b;
    layer2_outputs(712) <= not a;
    layer2_outputs(713) <= not a;
    layer2_outputs(714) <= a and not b;
    layer2_outputs(715) <= b;
    layer2_outputs(716) <= not b;
    layer2_outputs(717) <= not a;
    layer2_outputs(718) <= not b or a;
    layer2_outputs(719) <= a xor b;
    layer2_outputs(720) <= b and not a;
    layer2_outputs(721) <= not b or a;
    layer2_outputs(722) <= a xor b;
    layer2_outputs(723) <= not b or a;
    layer2_outputs(724) <= not b or a;
    layer2_outputs(725) <= a and b;
    layer2_outputs(726) <= a;
    layer2_outputs(727) <= not (a xor b);
    layer2_outputs(728) <= not (a or b);
    layer2_outputs(729) <= b and not a;
    layer2_outputs(730) <= not a or b;
    layer2_outputs(731) <= b;
    layer2_outputs(732) <= not b;
    layer2_outputs(733) <= b;
    layer2_outputs(734) <= not a;
    layer2_outputs(735) <= not a or b;
    layer2_outputs(736) <= not b;
    layer2_outputs(737) <= a or b;
    layer2_outputs(738) <= a;
    layer2_outputs(739) <= not (a xor b);
    layer2_outputs(740) <= 1'b1;
    layer2_outputs(741) <= b and not a;
    layer2_outputs(742) <= b and not a;
    layer2_outputs(743) <= a and not b;
    layer2_outputs(744) <= not b;
    layer2_outputs(745) <= a and not b;
    layer2_outputs(746) <= not b or a;
    layer2_outputs(747) <= a;
    layer2_outputs(748) <= b;
    layer2_outputs(749) <= not b;
    layer2_outputs(750) <= b and not a;
    layer2_outputs(751) <= 1'b1;
    layer2_outputs(752) <= a and not b;
    layer2_outputs(753) <= not a;
    layer2_outputs(754) <= a;
    layer2_outputs(755) <= a;
    layer2_outputs(756) <= not b;
    layer2_outputs(757) <= a and b;
    layer2_outputs(758) <= a xor b;
    layer2_outputs(759) <= 1'b0;
    layer2_outputs(760) <= a;
    layer2_outputs(761) <= not a;
    layer2_outputs(762) <= b;
    layer2_outputs(763) <= a;
    layer2_outputs(764) <= a;
    layer2_outputs(765) <= a and b;
    layer2_outputs(766) <= not (a xor b);
    layer2_outputs(767) <= b;
    layer2_outputs(768) <= not a;
    layer2_outputs(769) <= a and not b;
    layer2_outputs(770) <= not a;
    layer2_outputs(771) <= 1'b0;
    layer2_outputs(772) <= not b;
    layer2_outputs(773) <= a xor b;
    layer2_outputs(774) <= a and not b;
    layer2_outputs(775) <= not (a or b);
    layer2_outputs(776) <= b;
    layer2_outputs(777) <= not (a and b);
    layer2_outputs(778) <= not a;
    layer2_outputs(779) <= a;
    layer2_outputs(780) <= a or b;
    layer2_outputs(781) <= b;
    layer2_outputs(782) <= a;
    layer2_outputs(783) <= not a or b;
    layer2_outputs(784) <= not (a xor b);
    layer2_outputs(785) <= not a;
    layer2_outputs(786) <= not b;
    layer2_outputs(787) <= not b or a;
    layer2_outputs(788) <= not a;
    layer2_outputs(789) <= not b;
    layer2_outputs(790) <= not a;
    layer2_outputs(791) <= not a;
    layer2_outputs(792) <= not b;
    layer2_outputs(793) <= a or b;
    layer2_outputs(794) <= not (a or b);
    layer2_outputs(795) <= a xor b;
    layer2_outputs(796) <= a xor b;
    layer2_outputs(797) <= not (a or b);
    layer2_outputs(798) <= not a;
    layer2_outputs(799) <= b and not a;
    layer2_outputs(800) <= a and b;
    layer2_outputs(801) <= b;
    layer2_outputs(802) <= a and b;
    layer2_outputs(803) <= not (a and b);
    layer2_outputs(804) <= not a;
    layer2_outputs(805) <= not (a xor b);
    layer2_outputs(806) <= a xor b;
    layer2_outputs(807) <= 1'b0;
    layer2_outputs(808) <= b;
    layer2_outputs(809) <= not a;
    layer2_outputs(810) <= not b;
    layer2_outputs(811) <= not (a xor b);
    layer2_outputs(812) <= not (a xor b);
    layer2_outputs(813) <= a and not b;
    layer2_outputs(814) <= a xor b;
    layer2_outputs(815) <= a and b;
    layer2_outputs(816) <= a and b;
    layer2_outputs(817) <= a and not b;
    layer2_outputs(818) <= not b;
    layer2_outputs(819) <= not (a and b);
    layer2_outputs(820) <= b and not a;
    layer2_outputs(821) <= not b;
    layer2_outputs(822) <= not b;
    layer2_outputs(823) <= not a or b;
    layer2_outputs(824) <= not b;
    layer2_outputs(825) <= not a or b;
    layer2_outputs(826) <= b;
    layer2_outputs(827) <= not (a xor b);
    layer2_outputs(828) <= a and b;
    layer2_outputs(829) <= not b;
    layer2_outputs(830) <= not (a and b);
    layer2_outputs(831) <= b;
    layer2_outputs(832) <= not a or b;
    layer2_outputs(833) <= not a;
    layer2_outputs(834) <= a and not b;
    layer2_outputs(835) <= a;
    layer2_outputs(836) <= not b or a;
    layer2_outputs(837) <= a xor b;
    layer2_outputs(838) <= not b;
    layer2_outputs(839) <= not a or b;
    layer2_outputs(840) <= a and not b;
    layer2_outputs(841) <= not (a xor b);
    layer2_outputs(842) <= not (a xor b);
    layer2_outputs(843) <= a and b;
    layer2_outputs(844) <= b and not a;
    layer2_outputs(845) <= b;
    layer2_outputs(846) <= not (a and b);
    layer2_outputs(847) <= a;
    layer2_outputs(848) <= not b or a;
    layer2_outputs(849) <= a and not b;
    layer2_outputs(850) <= b;
    layer2_outputs(851) <= not (a xor b);
    layer2_outputs(852) <= not a or b;
    layer2_outputs(853) <= a;
    layer2_outputs(854) <= a xor b;
    layer2_outputs(855) <= not (a or b);
    layer2_outputs(856) <= not b or a;
    layer2_outputs(857) <= b;
    layer2_outputs(858) <= not (a or b);
    layer2_outputs(859) <= not b;
    layer2_outputs(860) <= a xor b;
    layer2_outputs(861) <= not b;
    layer2_outputs(862) <= a or b;
    layer2_outputs(863) <= a and not b;
    layer2_outputs(864) <= a;
    layer2_outputs(865) <= not b or a;
    layer2_outputs(866) <= a and not b;
    layer2_outputs(867) <= not (a and b);
    layer2_outputs(868) <= a;
    layer2_outputs(869) <= a xor b;
    layer2_outputs(870) <= not b or a;
    layer2_outputs(871) <= not (a xor b);
    layer2_outputs(872) <= a;
    layer2_outputs(873) <= not a or b;
    layer2_outputs(874) <= b;
    layer2_outputs(875) <= not (a and b);
    layer2_outputs(876) <= not (a or b);
    layer2_outputs(877) <= a and b;
    layer2_outputs(878) <= a;
    layer2_outputs(879) <= not b or a;
    layer2_outputs(880) <= a;
    layer2_outputs(881) <= not b or a;
    layer2_outputs(882) <= a xor b;
    layer2_outputs(883) <= a and b;
    layer2_outputs(884) <= a;
    layer2_outputs(885) <= a;
    layer2_outputs(886) <= a and not b;
    layer2_outputs(887) <= b and not a;
    layer2_outputs(888) <= not (a xor b);
    layer2_outputs(889) <= not a or b;
    layer2_outputs(890) <= not a or b;
    layer2_outputs(891) <= a;
    layer2_outputs(892) <= a;
    layer2_outputs(893) <= b;
    layer2_outputs(894) <= a xor b;
    layer2_outputs(895) <= not a or b;
    layer2_outputs(896) <= a xor b;
    layer2_outputs(897) <= a and not b;
    layer2_outputs(898) <= not (a xor b);
    layer2_outputs(899) <= not (a or b);
    layer2_outputs(900) <= not (a and b);
    layer2_outputs(901) <= b;
    layer2_outputs(902) <= not b;
    layer2_outputs(903) <= a and b;
    layer2_outputs(904) <= not (a xor b);
    layer2_outputs(905) <= not a or b;
    layer2_outputs(906) <= not a or b;
    layer2_outputs(907) <= not a or b;
    layer2_outputs(908) <= a and b;
    layer2_outputs(909) <= a;
    layer2_outputs(910) <= b;
    layer2_outputs(911) <= a xor b;
    layer2_outputs(912) <= a and not b;
    layer2_outputs(913) <= a;
    layer2_outputs(914) <= not (a xor b);
    layer2_outputs(915) <= b;
    layer2_outputs(916) <= not (a xor b);
    layer2_outputs(917) <= not b;
    layer2_outputs(918) <= not (a xor b);
    layer2_outputs(919) <= not a;
    layer2_outputs(920) <= not (a and b);
    layer2_outputs(921) <= not a or b;
    layer2_outputs(922) <= not a;
    layer2_outputs(923) <= a;
    layer2_outputs(924) <= a or b;
    layer2_outputs(925) <= not a;
    layer2_outputs(926) <= a and b;
    layer2_outputs(927) <= not (a and b);
    layer2_outputs(928) <= a and not b;
    layer2_outputs(929) <= b;
    layer2_outputs(930) <= not (a or b);
    layer2_outputs(931) <= b;
    layer2_outputs(932) <= not b;
    layer2_outputs(933) <= a and not b;
    layer2_outputs(934) <= not a;
    layer2_outputs(935) <= not (a xor b);
    layer2_outputs(936) <= a xor b;
    layer2_outputs(937) <= a and not b;
    layer2_outputs(938) <= a xor b;
    layer2_outputs(939) <= a and not b;
    layer2_outputs(940) <= a xor b;
    layer2_outputs(941) <= a or b;
    layer2_outputs(942) <= a and b;
    layer2_outputs(943) <= not b;
    layer2_outputs(944) <= a;
    layer2_outputs(945) <= a;
    layer2_outputs(946) <= not a;
    layer2_outputs(947) <= a;
    layer2_outputs(948) <= not b;
    layer2_outputs(949) <= not b or a;
    layer2_outputs(950) <= a xor b;
    layer2_outputs(951) <= not b;
    layer2_outputs(952) <= a or b;
    layer2_outputs(953) <= b and not a;
    layer2_outputs(954) <= a and b;
    layer2_outputs(955) <= b and not a;
    layer2_outputs(956) <= not (a and b);
    layer2_outputs(957) <= not b or a;
    layer2_outputs(958) <= not (a xor b);
    layer2_outputs(959) <= not a or b;
    layer2_outputs(960) <= not (a or b);
    layer2_outputs(961) <= a or b;
    layer2_outputs(962) <= a and b;
    layer2_outputs(963) <= a xor b;
    layer2_outputs(964) <= b;
    layer2_outputs(965) <= not (a or b);
    layer2_outputs(966) <= a;
    layer2_outputs(967) <= 1'b0;
    layer2_outputs(968) <= not a;
    layer2_outputs(969) <= not (a and b);
    layer2_outputs(970) <= b;
    layer2_outputs(971) <= not (a and b);
    layer2_outputs(972) <= a;
    layer2_outputs(973) <= not (a and b);
    layer2_outputs(974) <= a;
    layer2_outputs(975) <= not b;
    layer2_outputs(976) <= not a;
    layer2_outputs(977) <= b and not a;
    layer2_outputs(978) <= not (a or b);
    layer2_outputs(979) <= a or b;
    layer2_outputs(980) <= a xor b;
    layer2_outputs(981) <= a and not b;
    layer2_outputs(982) <= a;
    layer2_outputs(983) <= not b;
    layer2_outputs(984) <= not (a xor b);
    layer2_outputs(985) <= not a;
    layer2_outputs(986) <= not b;
    layer2_outputs(987) <= a;
    layer2_outputs(988) <= not (a xor b);
    layer2_outputs(989) <= a and b;
    layer2_outputs(990) <= not b or a;
    layer2_outputs(991) <= b and not a;
    layer2_outputs(992) <= not b;
    layer2_outputs(993) <= not (a or b);
    layer2_outputs(994) <= not b;
    layer2_outputs(995) <= b and not a;
    layer2_outputs(996) <= not a;
    layer2_outputs(997) <= a xor b;
    layer2_outputs(998) <= b;
    layer2_outputs(999) <= a and not b;
    layer2_outputs(1000) <= not a or b;
    layer2_outputs(1001) <= not (a or b);
    layer2_outputs(1002) <= not a;
    layer2_outputs(1003) <= a and b;
    layer2_outputs(1004) <= not (a and b);
    layer2_outputs(1005) <= not a;
    layer2_outputs(1006) <= a and not b;
    layer2_outputs(1007) <= b;
    layer2_outputs(1008) <= not (a and b);
    layer2_outputs(1009) <= a and not b;
    layer2_outputs(1010) <= b;
    layer2_outputs(1011) <= not a or b;
    layer2_outputs(1012) <= not (a and b);
    layer2_outputs(1013) <= a;
    layer2_outputs(1014) <= a or b;
    layer2_outputs(1015) <= not b or a;
    layer2_outputs(1016) <= not a;
    layer2_outputs(1017) <= b;
    layer2_outputs(1018) <= a and not b;
    layer2_outputs(1019) <= 1'b0;
    layer2_outputs(1020) <= not a;
    layer2_outputs(1021) <= a;
    layer2_outputs(1022) <= not (a or b);
    layer2_outputs(1023) <= not b or a;
    layer2_outputs(1024) <= a and not b;
    layer2_outputs(1025) <= not (a xor b);
    layer2_outputs(1026) <= a xor b;
    layer2_outputs(1027) <= not a or b;
    layer2_outputs(1028) <= b and not a;
    layer2_outputs(1029) <= a or b;
    layer2_outputs(1030) <= a;
    layer2_outputs(1031) <= a;
    layer2_outputs(1032) <= a or b;
    layer2_outputs(1033) <= a xor b;
    layer2_outputs(1034) <= a and not b;
    layer2_outputs(1035) <= a and not b;
    layer2_outputs(1036) <= b;
    layer2_outputs(1037) <= b;
    layer2_outputs(1038) <= b;
    layer2_outputs(1039) <= a and b;
    layer2_outputs(1040) <= b;
    layer2_outputs(1041) <= not a or b;
    layer2_outputs(1042) <= 1'b1;
    layer2_outputs(1043) <= a;
    layer2_outputs(1044) <= a and b;
    layer2_outputs(1045) <= not a;
    layer2_outputs(1046) <= not a;
    layer2_outputs(1047) <= a xor b;
    layer2_outputs(1048) <= not b;
    layer2_outputs(1049) <= a or b;
    layer2_outputs(1050) <= 1'b1;
    layer2_outputs(1051) <= not b or a;
    layer2_outputs(1052) <= a and b;
    layer2_outputs(1053) <= not b or a;
    layer2_outputs(1054) <= b and not a;
    layer2_outputs(1055) <= not a or b;
    layer2_outputs(1056) <= b and not a;
    layer2_outputs(1057) <= not b;
    layer2_outputs(1058) <= not a or b;
    layer2_outputs(1059) <= not a or b;
    layer2_outputs(1060) <= a and not b;
    layer2_outputs(1061) <= a and b;
    layer2_outputs(1062) <= a;
    layer2_outputs(1063) <= not (a and b);
    layer2_outputs(1064) <= not (a and b);
    layer2_outputs(1065) <= b;
    layer2_outputs(1066) <= not a;
    layer2_outputs(1067) <= not (a xor b);
    layer2_outputs(1068) <= not (a or b);
    layer2_outputs(1069) <= not b;
    layer2_outputs(1070) <= not (a xor b);
    layer2_outputs(1071) <= not a or b;
    layer2_outputs(1072) <= a or b;
    layer2_outputs(1073) <= a xor b;
    layer2_outputs(1074) <= not (a or b);
    layer2_outputs(1075) <= not (a and b);
    layer2_outputs(1076) <= b and not a;
    layer2_outputs(1077) <= b;
    layer2_outputs(1078) <= not (a or b);
    layer2_outputs(1079) <= not b;
    layer2_outputs(1080) <= not b or a;
    layer2_outputs(1081) <= a or b;
    layer2_outputs(1082) <= not b or a;
    layer2_outputs(1083) <= not (a and b);
    layer2_outputs(1084) <= a and not b;
    layer2_outputs(1085) <= not a;
    layer2_outputs(1086) <= a;
    layer2_outputs(1087) <= b;
    layer2_outputs(1088) <= a;
    layer2_outputs(1089) <= a and b;
    layer2_outputs(1090) <= a or b;
    layer2_outputs(1091) <= not a;
    layer2_outputs(1092) <= b;
    layer2_outputs(1093) <= not (a and b);
    layer2_outputs(1094) <= a xor b;
    layer2_outputs(1095) <= b and not a;
    layer2_outputs(1096) <= b;
    layer2_outputs(1097) <= not b or a;
    layer2_outputs(1098) <= a or b;
    layer2_outputs(1099) <= not a or b;
    layer2_outputs(1100) <= not (a xor b);
    layer2_outputs(1101) <= not (a and b);
    layer2_outputs(1102) <= a;
    layer2_outputs(1103) <= not a or b;
    layer2_outputs(1104) <= not (a and b);
    layer2_outputs(1105) <= not b;
    layer2_outputs(1106) <= a and not b;
    layer2_outputs(1107) <= 1'b1;
    layer2_outputs(1108) <= not b or a;
    layer2_outputs(1109) <= not b;
    layer2_outputs(1110) <= a;
    layer2_outputs(1111) <= not (a or b);
    layer2_outputs(1112) <= not (a and b);
    layer2_outputs(1113) <= a and not b;
    layer2_outputs(1114) <= a xor b;
    layer2_outputs(1115) <= not b;
    layer2_outputs(1116) <= not b or a;
    layer2_outputs(1117) <= a and b;
    layer2_outputs(1118) <= not a or b;
    layer2_outputs(1119) <= a;
    layer2_outputs(1120) <= a xor b;
    layer2_outputs(1121) <= not (a xor b);
    layer2_outputs(1122) <= not a or b;
    layer2_outputs(1123) <= not (a or b);
    layer2_outputs(1124) <= b;
    layer2_outputs(1125) <= a and b;
    layer2_outputs(1126) <= a or b;
    layer2_outputs(1127) <= not a or b;
    layer2_outputs(1128) <= not b;
    layer2_outputs(1129) <= a;
    layer2_outputs(1130) <= not a or b;
    layer2_outputs(1131) <= a or b;
    layer2_outputs(1132) <= not a or b;
    layer2_outputs(1133) <= not a or b;
    layer2_outputs(1134) <= b;
    layer2_outputs(1135) <= a or b;
    layer2_outputs(1136) <= not (a xor b);
    layer2_outputs(1137) <= b;
    layer2_outputs(1138) <= b and not a;
    layer2_outputs(1139) <= not a or b;
    layer2_outputs(1140) <= not (a or b);
    layer2_outputs(1141) <= b;
    layer2_outputs(1142) <= a or b;
    layer2_outputs(1143) <= b;
    layer2_outputs(1144) <= not b;
    layer2_outputs(1145) <= a;
    layer2_outputs(1146) <= a and b;
    layer2_outputs(1147) <= b and not a;
    layer2_outputs(1148) <= not (a and b);
    layer2_outputs(1149) <= a xor b;
    layer2_outputs(1150) <= not (a and b);
    layer2_outputs(1151) <= not b;
    layer2_outputs(1152) <= a xor b;
    layer2_outputs(1153) <= not b;
    layer2_outputs(1154) <= b and not a;
    layer2_outputs(1155) <= a and not b;
    layer2_outputs(1156) <= not b or a;
    layer2_outputs(1157) <= a or b;
    layer2_outputs(1158) <= not a;
    layer2_outputs(1159) <= not b;
    layer2_outputs(1160) <= b;
    layer2_outputs(1161) <= not (a xor b);
    layer2_outputs(1162) <= b and not a;
    layer2_outputs(1163) <= not (a and b);
    layer2_outputs(1164) <= a xor b;
    layer2_outputs(1165) <= a xor b;
    layer2_outputs(1166) <= a xor b;
    layer2_outputs(1167) <= not a;
    layer2_outputs(1168) <= b;
    layer2_outputs(1169) <= not b;
    layer2_outputs(1170) <= not (a xor b);
    layer2_outputs(1171) <= a;
    layer2_outputs(1172) <= a or b;
    layer2_outputs(1173) <= a;
    layer2_outputs(1174) <= a and b;
    layer2_outputs(1175) <= not (a and b);
    layer2_outputs(1176) <= not b or a;
    layer2_outputs(1177) <= not b or a;
    layer2_outputs(1178) <= b;
    layer2_outputs(1179) <= a xor b;
    layer2_outputs(1180) <= a xor b;
    layer2_outputs(1181) <= not a;
    layer2_outputs(1182) <= b and not a;
    layer2_outputs(1183) <= not b;
    layer2_outputs(1184) <= b;
    layer2_outputs(1185) <= a and not b;
    layer2_outputs(1186) <= b;
    layer2_outputs(1187) <= not b or a;
    layer2_outputs(1188) <= a;
    layer2_outputs(1189) <= not (a and b);
    layer2_outputs(1190) <= not a or b;
    layer2_outputs(1191) <= not (a or b);
    layer2_outputs(1192) <= a and not b;
    layer2_outputs(1193) <= a and b;
    layer2_outputs(1194) <= a xor b;
    layer2_outputs(1195) <= a and b;
    layer2_outputs(1196) <= not b;
    layer2_outputs(1197) <= not b;
    layer2_outputs(1198) <= not (a xor b);
    layer2_outputs(1199) <= b;
    layer2_outputs(1200) <= b and not a;
    layer2_outputs(1201) <= not (a or b);
    layer2_outputs(1202) <= not a;
    layer2_outputs(1203) <= not b;
    layer2_outputs(1204) <= not b or a;
    layer2_outputs(1205) <= not b or a;
    layer2_outputs(1206) <= b and not a;
    layer2_outputs(1207) <= a;
    layer2_outputs(1208) <= a and not b;
    layer2_outputs(1209) <= not (a xor b);
    layer2_outputs(1210) <= not b;
    layer2_outputs(1211) <= a and not b;
    layer2_outputs(1212) <= a and not b;
    layer2_outputs(1213) <= not a or b;
    layer2_outputs(1214) <= a or b;
    layer2_outputs(1215) <= not b or a;
    layer2_outputs(1216) <= not (a and b);
    layer2_outputs(1217) <= not (a xor b);
    layer2_outputs(1218) <= b;
    layer2_outputs(1219) <= not a or b;
    layer2_outputs(1220) <= a xor b;
    layer2_outputs(1221) <= not b or a;
    layer2_outputs(1222) <= not (a or b);
    layer2_outputs(1223) <= a xor b;
    layer2_outputs(1224) <= b;
    layer2_outputs(1225) <= not b or a;
    layer2_outputs(1226) <= a or b;
    layer2_outputs(1227) <= b;
    layer2_outputs(1228) <= not (a xor b);
    layer2_outputs(1229) <= a or b;
    layer2_outputs(1230) <= not (a and b);
    layer2_outputs(1231) <= not b;
    layer2_outputs(1232) <= a;
    layer2_outputs(1233) <= b;
    layer2_outputs(1234) <= not b;
    layer2_outputs(1235) <= not b or a;
    layer2_outputs(1236) <= a or b;
    layer2_outputs(1237) <= not a;
    layer2_outputs(1238) <= 1'b0;
    layer2_outputs(1239) <= not a;
    layer2_outputs(1240) <= a xor b;
    layer2_outputs(1241) <= not b;
    layer2_outputs(1242) <= a or b;
    layer2_outputs(1243) <= not (a or b);
    layer2_outputs(1244) <= a;
    layer2_outputs(1245) <= not b;
    layer2_outputs(1246) <= not b;
    layer2_outputs(1247) <= a and b;
    layer2_outputs(1248) <= a;
    layer2_outputs(1249) <= not b or a;
    layer2_outputs(1250) <= not (a and b);
    layer2_outputs(1251) <= a or b;
    layer2_outputs(1252) <= a;
    layer2_outputs(1253) <= not b;
    layer2_outputs(1254) <= a;
    layer2_outputs(1255) <= a;
    layer2_outputs(1256) <= not a or b;
    layer2_outputs(1257) <= a;
    layer2_outputs(1258) <= b;
    layer2_outputs(1259) <= not (a and b);
    layer2_outputs(1260) <= b;
    layer2_outputs(1261) <= not (a or b);
    layer2_outputs(1262) <= not a;
    layer2_outputs(1263) <= a;
    layer2_outputs(1264) <= not (a xor b);
    layer2_outputs(1265) <= a and not b;
    layer2_outputs(1266) <= a and b;
    layer2_outputs(1267) <= not (a xor b);
    layer2_outputs(1268) <= not a;
    layer2_outputs(1269) <= a and not b;
    layer2_outputs(1270) <= b;
    layer2_outputs(1271) <= b;
    layer2_outputs(1272) <= b and not a;
    layer2_outputs(1273) <= a or b;
    layer2_outputs(1274) <= a and not b;
    layer2_outputs(1275) <= 1'b1;
    layer2_outputs(1276) <= a xor b;
    layer2_outputs(1277) <= b;
    layer2_outputs(1278) <= not a;
    layer2_outputs(1279) <= not b;
    layer2_outputs(1280) <= not a;
    layer2_outputs(1281) <= not (a xor b);
    layer2_outputs(1282) <= a and b;
    layer2_outputs(1283) <= b;
    layer2_outputs(1284) <= a xor b;
    layer2_outputs(1285) <= b;
    layer2_outputs(1286) <= a or b;
    layer2_outputs(1287) <= not (a and b);
    layer2_outputs(1288) <= not b;
    layer2_outputs(1289) <= a;
    layer2_outputs(1290) <= a;
    layer2_outputs(1291) <= a and b;
    layer2_outputs(1292) <= a and b;
    layer2_outputs(1293) <= not (a xor b);
    layer2_outputs(1294) <= b;
    layer2_outputs(1295) <= not b;
    layer2_outputs(1296) <= a;
    layer2_outputs(1297) <= a and b;
    layer2_outputs(1298) <= not (a or b);
    layer2_outputs(1299) <= not a or b;
    layer2_outputs(1300) <= not b;
    layer2_outputs(1301) <= not (a or b);
    layer2_outputs(1302) <= b;
    layer2_outputs(1303) <= not (a and b);
    layer2_outputs(1304) <= not b;
    layer2_outputs(1305) <= not (a or b);
    layer2_outputs(1306) <= a;
    layer2_outputs(1307) <= not (a xor b);
    layer2_outputs(1308) <= 1'b0;
    layer2_outputs(1309) <= not (a or b);
    layer2_outputs(1310) <= b;
    layer2_outputs(1311) <= b;
    layer2_outputs(1312) <= not a or b;
    layer2_outputs(1313) <= not (a or b);
    layer2_outputs(1314) <= not (a xor b);
    layer2_outputs(1315) <= not b;
    layer2_outputs(1316) <= b;
    layer2_outputs(1317) <= not (a xor b);
    layer2_outputs(1318) <= b and not a;
    layer2_outputs(1319) <= a or b;
    layer2_outputs(1320) <= not (a or b);
    layer2_outputs(1321) <= a and b;
    layer2_outputs(1322) <= not (a and b);
    layer2_outputs(1323) <= a xor b;
    layer2_outputs(1324) <= not a;
    layer2_outputs(1325) <= a and not b;
    layer2_outputs(1326) <= not b or a;
    layer2_outputs(1327) <= b;
    layer2_outputs(1328) <= a and b;
    layer2_outputs(1329) <= not (a or b);
    layer2_outputs(1330) <= 1'b0;
    layer2_outputs(1331) <= not (a and b);
    layer2_outputs(1332) <= a and b;
    layer2_outputs(1333) <= b and not a;
    layer2_outputs(1334) <= not b;
    layer2_outputs(1335) <= not (a xor b);
    layer2_outputs(1336) <= a and not b;
    layer2_outputs(1337) <= not b or a;
    layer2_outputs(1338) <= a and not b;
    layer2_outputs(1339) <= not (a or b);
    layer2_outputs(1340) <= a and b;
    layer2_outputs(1341) <= a and not b;
    layer2_outputs(1342) <= not b or a;
    layer2_outputs(1343) <= a;
    layer2_outputs(1344) <= not a;
    layer2_outputs(1345) <= not (a xor b);
    layer2_outputs(1346) <= a;
    layer2_outputs(1347) <= not b;
    layer2_outputs(1348) <= not (a or b);
    layer2_outputs(1349) <= not b;
    layer2_outputs(1350) <= a;
    layer2_outputs(1351) <= not b;
    layer2_outputs(1352) <= not (a and b);
    layer2_outputs(1353) <= a or b;
    layer2_outputs(1354) <= b;
    layer2_outputs(1355) <= b;
    layer2_outputs(1356) <= not a or b;
    layer2_outputs(1357) <= b;
    layer2_outputs(1358) <= b and not a;
    layer2_outputs(1359) <= a;
    layer2_outputs(1360) <= not (a or b);
    layer2_outputs(1361) <= not (a and b);
    layer2_outputs(1362) <= a and not b;
    layer2_outputs(1363) <= b;
    layer2_outputs(1364) <= not (a or b);
    layer2_outputs(1365) <= not a;
    layer2_outputs(1366) <= not (a and b);
    layer2_outputs(1367) <= not (a xor b);
    layer2_outputs(1368) <= not b;
    layer2_outputs(1369) <= not (a or b);
    layer2_outputs(1370) <= not (a and b);
    layer2_outputs(1371) <= b;
    layer2_outputs(1372) <= a or b;
    layer2_outputs(1373) <= not b or a;
    layer2_outputs(1374) <= a and not b;
    layer2_outputs(1375) <= a;
    layer2_outputs(1376) <= b;
    layer2_outputs(1377) <= not b;
    layer2_outputs(1378) <= a;
    layer2_outputs(1379) <= not b;
    layer2_outputs(1380) <= not a;
    layer2_outputs(1381) <= a;
    layer2_outputs(1382) <= not (a and b);
    layer2_outputs(1383) <= a and not b;
    layer2_outputs(1384) <= not (a and b);
    layer2_outputs(1385) <= not a;
    layer2_outputs(1386) <= a xor b;
    layer2_outputs(1387) <= not a;
    layer2_outputs(1388) <= not a;
    layer2_outputs(1389) <= not a;
    layer2_outputs(1390) <= b;
    layer2_outputs(1391) <= a and not b;
    layer2_outputs(1392) <= not (a xor b);
    layer2_outputs(1393) <= not (a or b);
    layer2_outputs(1394) <= not (a xor b);
    layer2_outputs(1395) <= b and not a;
    layer2_outputs(1396) <= a and b;
    layer2_outputs(1397) <= not a;
    layer2_outputs(1398) <= not b;
    layer2_outputs(1399) <= b and not a;
    layer2_outputs(1400) <= a or b;
    layer2_outputs(1401) <= a;
    layer2_outputs(1402) <= a;
    layer2_outputs(1403) <= a and not b;
    layer2_outputs(1404) <= not (a xor b);
    layer2_outputs(1405) <= not (a and b);
    layer2_outputs(1406) <= not (a or b);
    layer2_outputs(1407) <= not a;
    layer2_outputs(1408) <= a and not b;
    layer2_outputs(1409) <= a and b;
    layer2_outputs(1410) <= not a or b;
    layer2_outputs(1411) <= b and not a;
    layer2_outputs(1412) <= not b;
    layer2_outputs(1413) <= not (a xor b);
    layer2_outputs(1414) <= a;
    layer2_outputs(1415) <= not a;
    layer2_outputs(1416) <= a and not b;
    layer2_outputs(1417) <= not (a xor b);
    layer2_outputs(1418) <= not (a xor b);
    layer2_outputs(1419) <= not (a and b);
    layer2_outputs(1420) <= a xor b;
    layer2_outputs(1421) <= not (a xor b);
    layer2_outputs(1422) <= not a;
    layer2_outputs(1423) <= not (a or b);
    layer2_outputs(1424) <= b and not a;
    layer2_outputs(1425) <= b;
    layer2_outputs(1426) <= a or b;
    layer2_outputs(1427) <= not (a or b);
    layer2_outputs(1428) <= a or b;
    layer2_outputs(1429) <= not b or a;
    layer2_outputs(1430) <= b and not a;
    layer2_outputs(1431) <= a;
    layer2_outputs(1432) <= not a or b;
    layer2_outputs(1433) <= not (a or b);
    layer2_outputs(1434) <= not b;
    layer2_outputs(1435) <= not (a or b);
    layer2_outputs(1436) <= not (a and b);
    layer2_outputs(1437) <= a;
    layer2_outputs(1438) <= a and not b;
    layer2_outputs(1439) <= not a;
    layer2_outputs(1440) <= a or b;
    layer2_outputs(1441) <= not b or a;
    layer2_outputs(1442) <= b;
    layer2_outputs(1443) <= not b or a;
    layer2_outputs(1444) <= not (a and b);
    layer2_outputs(1445) <= b;
    layer2_outputs(1446) <= not (a xor b);
    layer2_outputs(1447) <= not a or b;
    layer2_outputs(1448) <= not b;
    layer2_outputs(1449) <= a;
    layer2_outputs(1450) <= b and not a;
    layer2_outputs(1451) <= not a;
    layer2_outputs(1452) <= not b or a;
    layer2_outputs(1453) <= b and not a;
    layer2_outputs(1454) <= not (a and b);
    layer2_outputs(1455) <= b;
    layer2_outputs(1456) <= a;
    layer2_outputs(1457) <= not b;
    layer2_outputs(1458) <= a xor b;
    layer2_outputs(1459) <= not b;
    layer2_outputs(1460) <= not b;
    layer2_outputs(1461) <= a;
    layer2_outputs(1462) <= b and not a;
    layer2_outputs(1463) <= not (a xor b);
    layer2_outputs(1464) <= 1'b0;
    layer2_outputs(1465) <= not (a xor b);
    layer2_outputs(1466) <= a or b;
    layer2_outputs(1467) <= b;
    layer2_outputs(1468) <= not a;
    layer2_outputs(1469) <= a and not b;
    layer2_outputs(1470) <= b and not a;
    layer2_outputs(1471) <= a and not b;
    layer2_outputs(1472) <= not (a or b);
    layer2_outputs(1473) <= not b;
    layer2_outputs(1474) <= a and b;
    layer2_outputs(1475) <= not b or a;
    layer2_outputs(1476) <= a xor b;
    layer2_outputs(1477) <= not (a and b);
    layer2_outputs(1478) <= not (a xor b);
    layer2_outputs(1479) <= a;
    layer2_outputs(1480) <= not (a xor b);
    layer2_outputs(1481) <= a and not b;
    layer2_outputs(1482) <= not (a xor b);
    layer2_outputs(1483) <= not a;
    layer2_outputs(1484) <= a and not b;
    layer2_outputs(1485) <= not b;
    layer2_outputs(1486) <= not b;
    layer2_outputs(1487) <= not (a xor b);
    layer2_outputs(1488) <= not a or b;
    layer2_outputs(1489) <= a xor b;
    layer2_outputs(1490) <= not a;
    layer2_outputs(1491) <= a or b;
    layer2_outputs(1492) <= a;
    layer2_outputs(1493) <= a;
    layer2_outputs(1494) <= b;
    layer2_outputs(1495) <= a;
    layer2_outputs(1496) <= not a;
    layer2_outputs(1497) <= a or b;
    layer2_outputs(1498) <= a and b;
    layer2_outputs(1499) <= b;
    layer2_outputs(1500) <= a or b;
    layer2_outputs(1501) <= a and not b;
    layer2_outputs(1502) <= b;
    layer2_outputs(1503) <= a;
    layer2_outputs(1504) <= not b or a;
    layer2_outputs(1505) <= a;
    layer2_outputs(1506) <= not b;
    layer2_outputs(1507) <= not b or a;
    layer2_outputs(1508) <= a or b;
    layer2_outputs(1509) <= not (a or b);
    layer2_outputs(1510) <= not (a and b);
    layer2_outputs(1511) <= a xor b;
    layer2_outputs(1512) <= not b;
    layer2_outputs(1513) <= not a;
    layer2_outputs(1514) <= not b;
    layer2_outputs(1515) <= not (a or b);
    layer2_outputs(1516) <= not b or a;
    layer2_outputs(1517) <= not b or a;
    layer2_outputs(1518) <= not (a and b);
    layer2_outputs(1519) <= a and b;
    layer2_outputs(1520) <= not b or a;
    layer2_outputs(1521) <= a xor b;
    layer2_outputs(1522) <= b;
    layer2_outputs(1523) <= not (a xor b);
    layer2_outputs(1524) <= a or b;
    layer2_outputs(1525) <= a and not b;
    layer2_outputs(1526) <= not b;
    layer2_outputs(1527) <= not b;
    layer2_outputs(1528) <= b and not a;
    layer2_outputs(1529) <= not a or b;
    layer2_outputs(1530) <= not (a and b);
    layer2_outputs(1531) <= a and not b;
    layer2_outputs(1532) <= a or b;
    layer2_outputs(1533) <= b;
    layer2_outputs(1534) <= not b;
    layer2_outputs(1535) <= not (a xor b);
    layer2_outputs(1536) <= not b;
    layer2_outputs(1537) <= not a;
    layer2_outputs(1538) <= a;
    layer2_outputs(1539) <= not b;
    layer2_outputs(1540) <= not a or b;
    layer2_outputs(1541) <= not b;
    layer2_outputs(1542) <= b;
    layer2_outputs(1543) <= a or b;
    layer2_outputs(1544) <= not b;
    layer2_outputs(1545) <= b and not a;
    layer2_outputs(1546) <= a;
    layer2_outputs(1547) <= a xor b;
    layer2_outputs(1548) <= b;
    layer2_outputs(1549) <= not b;
    layer2_outputs(1550) <= not (a xor b);
    layer2_outputs(1551) <= not b;
    layer2_outputs(1552) <= b and not a;
    layer2_outputs(1553) <= not b;
    layer2_outputs(1554) <= not (a and b);
    layer2_outputs(1555) <= not a;
    layer2_outputs(1556) <= not b or a;
    layer2_outputs(1557) <= not a;
    layer2_outputs(1558) <= a and not b;
    layer2_outputs(1559) <= not b or a;
    layer2_outputs(1560) <= not (a xor b);
    layer2_outputs(1561) <= not b or a;
    layer2_outputs(1562) <= a and b;
    layer2_outputs(1563) <= not a or b;
    layer2_outputs(1564) <= a xor b;
    layer2_outputs(1565) <= a;
    layer2_outputs(1566) <= b and not a;
    layer2_outputs(1567) <= not (a and b);
    layer2_outputs(1568) <= b;
    layer2_outputs(1569) <= a or b;
    layer2_outputs(1570) <= not (a and b);
    layer2_outputs(1571) <= not (a xor b);
    layer2_outputs(1572) <= not (a or b);
    layer2_outputs(1573) <= b;
    layer2_outputs(1574) <= not b or a;
    layer2_outputs(1575) <= not (a xor b);
    layer2_outputs(1576) <= not (a xor b);
    layer2_outputs(1577) <= not a;
    layer2_outputs(1578) <= a xor b;
    layer2_outputs(1579) <= 1'b0;
    layer2_outputs(1580) <= a and not b;
    layer2_outputs(1581) <= b;
    layer2_outputs(1582) <= not (a xor b);
    layer2_outputs(1583) <= not b;
    layer2_outputs(1584) <= a xor b;
    layer2_outputs(1585) <= not (a or b);
    layer2_outputs(1586) <= not a;
    layer2_outputs(1587) <= a and not b;
    layer2_outputs(1588) <= b and not a;
    layer2_outputs(1589) <= not (a xor b);
    layer2_outputs(1590) <= 1'b0;
    layer2_outputs(1591) <= a or b;
    layer2_outputs(1592) <= not b or a;
    layer2_outputs(1593) <= a or b;
    layer2_outputs(1594) <= not a or b;
    layer2_outputs(1595) <= a;
    layer2_outputs(1596) <= not (a xor b);
    layer2_outputs(1597) <= 1'b1;
    layer2_outputs(1598) <= a and b;
    layer2_outputs(1599) <= b and not a;
    layer2_outputs(1600) <= not a;
    layer2_outputs(1601) <= not b;
    layer2_outputs(1602) <= b;
    layer2_outputs(1603) <= a or b;
    layer2_outputs(1604) <= b;
    layer2_outputs(1605) <= a and b;
    layer2_outputs(1606) <= 1'b1;
    layer2_outputs(1607) <= b and not a;
    layer2_outputs(1608) <= a xor b;
    layer2_outputs(1609) <= b;
    layer2_outputs(1610) <= not (a and b);
    layer2_outputs(1611) <= not b;
    layer2_outputs(1612) <= not (a xor b);
    layer2_outputs(1613) <= not (a and b);
    layer2_outputs(1614) <= not (a xor b);
    layer2_outputs(1615) <= b;
    layer2_outputs(1616) <= a and not b;
    layer2_outputs(1617) <= a xor b;
    layer2_outputs(1618) <= not (a xor b);
    layer2_outputs(1619) <= not (a or b);
    layer2_outputs(1620) <= not a;
    layer2_outputs(1621) <= not b;
    layer2_outputs(1622) <= not (a xor b);
    layer2_outputs(1623) <= not b;
    layer2_outputs(1624) <= not b;
    layer2_outputs(1625) <= b;
    layer2_outputs(1626) <= a and b;
    layer2_outputs(1627) <= not (a xor b);
    layer2_outputs(1628) <= not a;
    layer2_outputs(1629) <= not a;
    layer2_outputs(1630) <= a and b;
    layer2_outputs(1631) <= not b;
    layer2_outputs(1632) <= b;
    layer2_outputs(1633) <= not (a and b);
    layer2_outputs(1634) <= b and not a;
    layer2_outputs(1635) <= not a or b;
    layer2_outputs(1636) <= a xor b;
    layer2_outputs(1637) <= not (a or b);
    layer2_outputs(1638) <= a or b;
    layer2_outputs(1639) <= not (a or b);
    layer2_outputs(1640) <= not (a and b);
    layer2_outputs(1641) <= not (a xor b);
    layer2_outputs(1642) <= a and not b;
    layer2_outputs(1643) <= not b;
    layer2_outputs(1644) <= a;
    layer2_outputs(1645) <= a and b;
    layer2_outputs(1646) <= not (a xor b);
    layer2_outputs(1647) <= not a;
    layer2_outputs(1648) <= b;
    layer2_outputs(1649) <= not a or b;
    layer2_outputs(1650) <= not (a xor b);
    layer2_outputs(1651) <= not b;
    layer2_outputs(1652) <= a xor b;
    layer2_outputs(1653) <= not b;
    layer2_outputs(1654) <= b;
    layer2_outputs(1655) <= b;
    layer2_outputs(1656) <= b;
    layer2_outputs(1657) <= not a;
    layer2_outputs(1658) <= a xor b;
    layer2_outputs(1659) <= a xor b;
    layer2_outputs(1660) <= not b;
    layer2_outputs(1661) <= a or b;
    layer2_outputs(1662) <= a;
    layer2_outputs(1663) <= not (a xor b);
    layer2_outputs(1664) <= not b;
    layer2_outputs(1665) <= not b;
    layer2_outputs(1666) <= not a;
    layer2_outputs(1667) <= not (a xor b);
    layer2_outputs(1668) <= not (a and b);
    layer2_outputs(1669) <= not b or a;
    layer2_outputs(1670) <= a;
    layer2_outputs(1671) <= b;
    layer2_outputs(1672) <= a;
    layer2_outputs(1673) <= a and not b;
    layer2_outputs(1674) <= a xor b;
    layer2_outputs(1675) <= b and not a;
    layer2_outputs(1676) <= not b or a;
    layer2_outputs(1677) <= a xor b;
    layer2_outputs(1678) <= a and not b;
    layer2_outputs(1679) <= a xor b;
    layer2_outputs(1680) <= a;
    layer2_outputs(1681) <= b and not a;
    layer2_outputs(1682) <= b;
    layer2_outputs(1683) <= not a;
    layer2_outputs(1684) <= a;
    layer2_outputs(1685) <= not b;
    layer2_outputs(1686) <= b;
    layer2_outputs(1687) <= not b or a;
    layer2_outputs(1688) <= not a or b;
    layer2_outputs(1689) <= not a;
    layer2_outputs(1690) <= a xor b;
    layer2_outputs(1691) <= not a;
    layer2_outputs(1692) <= b and not a;
    layer2_outputs(1693) <= a or b;
    layer2_outputs(1694) <= not b or a;
    layer2_outputs(1695) <= not b or a;
    layer2_outputs(1696) <= not (a and b);
    layer2_outputs(1697) <= not (a or b);
    layer2_outputs(1698) <= a;
    layer2_outputs(1699) <= b and not a;
    layer2_outputs(1700) <= not (a or b);
    layer2_outputs(1701) <= not (a or b);
    layer2_outputs(1702) <= a;
    layer2_outputs(1703) <= b;
    layer2_outputs(1704) <= a and b;
    layer2_outputs(1705) <= not (a xor b);
    layer2_outputs(1706) <= a and b;
    layer2_outputs(1707) <= b and not a;
    layer2_outputs(1708) <= not b or a;
    layer2_outputs(1709) <= a and b;
    layer2_outputs(1710) <= not b or a;
    layer2_outputs(1711) <= not (a xor b);
    layer2_outputs(1712) <= not b;
    layer2_outputs(1713) <= not a;
    layer2_outputs(1714) <= not a or b;
    layer2_outputs(1715) <= a or b;
    layer2_outputs(1716) <= not a;
    layer2_outputs(1717) <= a xor b;
    layer2_outputs(1718) <= b;
    layer2_outputs(1719) <= b and not a;
    layer2_outputs(1720) <= not (a xor b);
    layer2_outputs(1721) <= not b or a;
    layer2_outputs(1722) <= b;
    layer2_outputs(1723) <= b;
    layer2_outputs(1724) <= a xor b;
    layer2_outputs(1725) <= not a;
    layer2_outputs(1726) <= b and not a;
    layer2_outputs(1727) <= not a;
    layer2_outputs(1728) <= a;
    layer2_outputs(1729) <= a;
    layer2_outputs(1730) <= not a;
    layer2_outputs(1731) <= not a;
    layer2_outputs(1732) <= b;
    layer2_outputs(1733) <= not a;
    layer2_outputs(1734) <= not a or b;
    layer2_outputs(1735) <= a or b;
    layer2_outputs(1736) <= not b or a;
    layer2_outputs(1737) <= a or b;
    layer2_outputs(1738) <= a xor b;
    layer2_outputs(1739) <= not a or b;
    layer2_outputs(1740) <= a and not b;
    layer2_outputs(1741) <= not a or b;
    layer2_outputs(1742) <= a;
    layer2_outputs(1743) <= b and not a;
    layer2_outputs(1744) <= b;
    layer2_outputs(1745) <= not (a and b);
    layer2_outputs(1746) <= b and not a;
    layer2_outputs(1747) <= b;
    layer2_outputs(1748) <= not (a or b);
    layer2_outputs(1749) <= a and b;
    layer2_outputs(1750) <= not b or a;
    layer2_outputs(1751) <= not b or a;
    layer2_outputs(1752) <= not (a and b);
    layer2_outputs(1753) <= a and not b;
    layer2_outputs(1754) <= 1'b0;
    layer2_outputs(1755) <= a or b;
    layer2_outputs(1756) <= not a or b;
    layer2_outputs(1757) <= b and not a;
    layer2_outputs(1758) <= a;
    layer2_outputs(1759) <= not b;
    layer2_outputs(1760) <= not b;
    layer2_outputs(1761) <= not (a or b);
    layer2_outputs(1762) <= a;
    layer2_outputs(1763) <= a and not b;
    layer2_outputs(1764) <= not (a and b);
    layer2_outputs(1765) <= a or b;
    layer2_outputs(1766) <= not b;
    layer2_outputs(1767) <= not (a xor b);
    layer2_outputs(1768) <= not b;
    layer2_outputs(1769) <= not b;
    layer2_outputs(1770) <= not a;
    layer2_outputs(1771) <= a xor b;
    layer2_outputs(1772) <= a and b;
    layer2_outputs(1773) <= not b;
    layer2_outputs(1774) <= not a or b;
    layer2_outputs(1775) <= not (a or b);
    layer2_outputs(1776) <= not a;
    layer2_outputs(1777) <= not b;
    layer2_outputs(1778) <= a xor b;
    layer2_outputs(1779) <= a xor b;
    layer2_outputs(1780) <= not a;
    layer2_outputs(1781) <= a;
    layer2_outputs(1782) <= a;
    layer2_outputs(1783) <= not b;
    layer2_outputs(1784) <= a xor b;
    layer2_outputs(1785) <= not (a and b);
    layer2_outputs(1786) <= a;
    layer2_outputs(1787) <= not b;
    layer2_outputs(1788) <= not (a xor b);
    layer2_outputs(1789) <= a xor b;
    layer2_outputs(1790) <= not (a or b);
    layer2_outputs(1791) <= not b or a;
    layer2_outputs(1792) <= b;
    layer2_outputs(1793) <= a xor b;
    layer2_outputs(1794) <= not b or a;
    layer2_outputs(1795) <= b and not a;
    layer2_outputs(1796) <= a;
    layer2_outputs(1797) <= a and b;
    layer2_outputs(1798) <= not b;
    layer2_outputs(1799) <= a;
    layer2_outputs(1800) <= not b;
    layer2_outputs(1801) <= b and not a;
    layer2_outputs(1802) <= not a;
    layer2_outputs(1803) <= b;
    layer2_outputs(1804) <= not (a or b);
    layer2_outputs(1805) <= a and not b;
    layer2_outputs(1806) <= a xor b;
    layer2_outputs(1807) <= not (a or b);
    layer2_outputs(1808) <= a xor b;
    layer2_outputs(1809) <= a;
    layer2_outputs(1810) <= a and b;
    layer2_outputs(1811) <= not b;
    layer2_outputs(1812) <= a and not b;
    layer2_outputs(1813) <= b;
    layer2_outputs(1814) <= not b or a;
    layer2_outputs(1815) <= not (a xor b);
    layer2_outputs(1816) <= a or b;
    layer2_outputs(1817) <= a xor b;
    layer2_outputs(1818) <= a xor b;
    layer2_outputs(1819) <= a and not b;
    layer2_outputs(1820) <= b;
    layer2_outputs(1821) <= not b;
    layer2_outputs(1822) <= not (a or b);
    layer2_outputs(1823) <= 1'b1;
    layer2_outputs(1824) <= a and not b;
    layer2_outputs(1825) <= a xor b;
    layer2_outputs(1826) <= not (a or b);
    layer2_outputs(1827) <= not a;
    layer2_outputs(1828) <= a;
    layer2_outputs(1829) <= b;
    layer2_outputs(1830) <= not b;
    layer2_outputs(1831) <= not (a and b);
    layer2_outputs(1832) <= a and not b;
    layer2_outputs(1833) <= b;
    layer2_outputs(1834) <= b and not a;
    layer2_outputs(1835) <= not b;
    layer2_outputs(1836) <= not a;
    layer2_outputs(1837) <= not a or b;
    layer2_outputs(1838) <= a xor b;
    layer2_outputs(1839) <= not b or a;
    layer2_outputs(1840) <= not (a and b);
    layer2_outputs(1841) <= a and b;
    layer2_outputs(1842) <= not a;
    layer2_outputs(1843) <= b;
    layer2_outputs(1844) <= not (a xor b);
    layer2_outputs(1845) <= not b;
    layer2_outputs(1846) <= not a or b;
    layer2_outputs(1847) <= not b;
    layer2_outputs(1848) <= not b;
    layer2_outputs(1849) <= a;
    layer2_outputs(1850) <= not a;
    layer2_outputs(1851) <= b and not a;
    layer2_outputs(1852) <= not b;
    layer2_outputs(1853) <= a xor b;
    layer2_outputs(1854) <= a;
    layer2_outputs(1855) <= not (a xor b);
    layer2_outputs(1856) <= not (a or b);
    layer2_outputs(1857) <= not b;
    layer2_outputs(1858) <= a and b;
    layer2_outputs(1859) <= a;
    layer2_outputs(1860) <= a;
    layer2_outputs(1861) <= b;
    layer2_outputs(1862) <= a;
    layer2_outputs(1863) <= a xor b;
    layer2_outputs(1864) <= b and not a;
    layer2_outputs(1865) <= a and b;
    layer2_outputs(1866) <= not b;
    layer2_outputs(1867) <= not (a or b);
    layer2_outputs(1868) <= not a or b;
    layer2_outputs(1869) <= a or b;
    layer2_outputs(1870) <= a or b;
    layer2_outputs(1871) <= a or b;
    layer2_outputs(1872) <= b and not a;
    layer2_outputs(1873) <= not b;
    layer2_outputs(1874) <= a or b;
    layer2_outputs(1875) <= not a;
    layer2_outputs(1876) <= b;
    layer2_outputs(1877) <= a or b;
    layer2_outputs(1878) <= not (a xor b);
    layer2_outputs(1879) <= not b;
    layer2_outputs(1880) <= not (a or b);
    layer2_outputs(1881) <= b;
    layer2_outputs(1882) <= not b;
    layer2_outputs(1883) <= not (a xor b);
    layer2_outputs(1884) <= not a;
    layer2_outputs(1885) <= not b;
    layer2_outputs(1886) <= a;
    layer2_outputs(1887) <= not a;
    layer2_outputs(1888) <= not (a xor b);
    layer2_outputs(1889) <= not b or a;
    layer2_outputs(1890) <= a xor b;
    layer2_outputs(1891) <= not a;
    layer2_outputs(1892) <= not (a and b);
    layer2_outputs(1893) <= not (a or b);
    layer2_outputs(1894) <= not b or a;
    layer2_outputs(1895) <= not a or b;
    layer2_outputs(1896) <= b and not a;
    layer2_outputs(1897) <= not b;
    layer2_outputs(1898) <= a xor b;
    layer2_outputs(1899) <= b and not a;
    layer2_outputs(1900) <= not (a or b);
    layer2_outputs(1901) <= b and not a;
    layer2_outputs(1902) <= a;
    layer2_outputs(1903) <= a and b;
    layer2_outputs(1904) <= not (a or b);
    layer2_outputs(1905) <= not b;
    layer2_outputs(1906) <= b;
    layer2_outputs(1907) <= b;
    layer2_outputs(1908) <= b;
    layer2_outputs(1909) <= not b;
    layer2_outputs(1910) <= b;
    layer2_outputs(1911) <= not (a or b);
    layer2_outputs(1912) <= not a or b;
    layer2_outputs(1913) <= not a;
    layer2_outputs(1914) <= a;
    layer2_outputs(1915) <= b and not a;
    layer2_outputs(1916) <= a or b;
    layer2_outputs(1917) <= b;
    layer2_outputs(1918) <= b;
    layer2_outputs(1919) <= a xor b;
    layer2_outputs(1920) <= not (a and b);
    layer2_outputs(1921) <= not b or a;
    layer2_outputs(1922) <= b;
    layer2_outputs(1923) <= not (a xor b);
    layer2_outputs(1924) <= b;
    layer2_outputs(1925) <= not b or a;
    layer2_outputs(1926) <= not a;
    layer2_outputs(1927) <= not (a and b);
    layer2_outputs(1928) <= a;
    layer2_outputs(1929) <= not (a xor b);
    layer2_outputs(1930) <= b;
    layer2_outputs(1931) <= not (a and b);
    layer2_outputs(1932) <= not b;
    layer2_outputs(1933) <= not b;
    layer2_outputs(1934) <= not a;
    layer2_outputs(1935) <= not a;
    layer2_outputs(1936) <= not (a or b);
    layer2_outputs(1937) <= a;
    layer2_outputs(1938) <= a and b;
    layer2_outputs(1939) <= a and b;
    layer2_outputs(1940) <= not (a xor b);
    layer2_outputs(1941) <= a;
    layer2_outputs(1942) <= b;
    layer2_outputs(1943) <= a and not b;
    layer2_outputs(1944) <= a and not b;
    layer2_outputs(1945) <= not (a or b);
    layer2_outputs(1946) <= not b;
    layer2_outputs(1947) <= not (a and b);
    layer2_outputs(1948) <= not b or a;
    layer2_outputs(1949) <= not a;
    layer2_outputs(1950) <= b;
    layer2_outputs(1951) <= not (a or b);
    layer2_outputs(1952) <= b;
    layer2_outputs(1953) <= not (a and b);
    layer2_outputs(1954) <= not a;
    layer2_outputs(1955) <= not b;
    layer2_outputs(1956) <= not b;
    layer2_outputs(1957) <= b and not a;
    layer2_outputs(1958) <= not (a and b);
    layer2_outputs(1959) <= a and not b;
    layer2_outputs(1960) <= not (a or b);
    layer2_outputs(1961) <= not a;
    layer2_outputs(1962) <= a;
    layer2_outputs(1963) <= b;
    layer2_outputs(1964) <= not (a xor b);
    layer2_outputs(1965) <= not a or b;
    layer2_outputs(1966) <= a;
    layer2_outputs(1967) <= not a;
    layer2_outputs(1968) <= not a;
    layer2_outputs(1969) <= a;
    layer2_outputs(1970) <= not b or a;
    layer2_outputs(1971) <= b and not a;
    layer2_outputs(1972) <= b;
    layer2_outputs(1973) <= not a;
    layer2_outputs(1974) <= not b;
    layer2_outputs(1975) <= a and not b;
    layer2_outputs(1976) <= a and not b;
    layer2_outputs(1977) <= a and not b;
    layer2_outputs(1978) <= not a;
    layer2_outputs(1979) <= not (a xor b);
    layer2_outputs(1980) <= not a;
    layer2_outputs(1981) <= a;
    layer2_outputs(1982) <= not b;
    layer2_outputs(1983) <= not a;
    layer2_outputs(1984) <= a;
    layer2_outputs(1985) <= not a;
    layer2_outputs(1986) <= not a;
    layer2_outputs(1987) <= not b;
    layer2_outputs(1988) <= a or b;
    layer2_outputs(1989) <= not b;
    layer2_outputs(1990) <= not b or a;
    layer2_outputs(1991) <= a and b;
    layer2_outputs(1992) <= a xor b;
    layer2_outputs(1993) <= not (a xor b);
    layer2_outputs(1994) <= not a;
    layer2_outputs(1995) <= b;
    layer2_outputs(1996) <= not (a xor b);
    layer2_outputs(1997) <= a;
    layer2_outputs(1998) <= not (a xor b);
    layer2_outputs(1999) <= b and not a;
    layer2_outputs(2000) <= a or b;
    layer2_outputs(2001) <= not (a and b);
    layer2_outputs(2002) <= a;
    layer2_outputs(2003) <= not (a xor b);
    layer2_outputs(2004) <= not a or b;
    layer2_outputs(2005) <= not (a and b);
    layer2_outputs(2006) <= not (a or b);
    layer2_outputs(2007) <= b;
    layer2_outputs(2008) <= not b;
    layer2_outputs(2009) <= b;
    layer2_outputs(2010) <= a;
    layer2_outputs(2011) <= not b;
    layer2_outputs(2012) <= b;
    layer2_outputs(2013) <= b and not a;
    layer2_outputs(2014) <= a and b;
    layer2_outputs(2015) <= not b;
    layer2_outputs(2016) <= a and not b;
    layer2_outputs(2017) <= not a;
    layer2_outputs(2018) <= a;
    layer2_outputs(2019) <= not a or b;
    layer2_outputs(2020) <= not (a or b);
    layer2_outputs(2021) <= a or b;
    layer2_outputs(2022) <= not a;
    layer2_outputs(2023) <= b;
    layer2_outputs(2024) <= b;
    layer2_outputs(2025) <= a and not b;
    layer2_outputs(2026) <= not a;
    layer2_outputs(2027) <= not (a xor b);
    layer2_outputs(2028) <= not b or a;
    layer2_outputs(2029) <= not (a and b);
    layer2_outputs(2030) <= b;
    layer2_outputs(2031) <= not (a xor b);
    layer2_outputs(2032) <= a and b;
    layer2_outputs(2033) <= not a or b;
    layer2_outputs(2034) <= a xor b;
    layer2_outputs(2035) <= not (a xor b);
    layer2_outputs(2036) <= not a or b;
    layer2_outputs(2037) <= b;
    layer2_outputs(2038) <= not a;
    layer2_outputs(2039) <= not a;
    layer2_outputs(2040) <= 1'b1;
    layer2_outputs(2041) <= not b or a;
    layer2_outputs(2042) <= b;
    layer2_outputs(2043) <= a;
    layer2_outputs(2044) <= b and not a;
    layer2_outputs(2045) <= a;
    layer2_outputs(2046) <= a xor b;
    layer2_outputs(2047) <= a or b;
    layer2_outputs(2048) <= not a;
    layer2_outputs(2049) <= a and not b;
    layer2_outputs(2050) <= not b;
    layer2_outputs(2051) <= not a;
    layer2_outputs(2052) <= not (a or b);
    layer2_outputs(2053) <= not (a xor b);
    layer2_outputs(2054) <= not a;
    layer2_outputs(2055) <= not (a and b);
    layer2_outputs(2056) <= b and not a;
    layer2_outputs(2057) <= not a;
    layer2_outputs(2058) <= b;
    layer2_outputs(2059) <= a;
    layer2_outputs(2060) <= a;
    layer2_outputs(2061) <= not (a and b);
    layer2_outputs(2062) <= not (a or b);
    layer2_outputs(2063) <= a and b;
    layer2_outputs(2064) <= b;
    layer2_outputs(2065) <= not a;
    layer2_outputs(2066) <= not (a and b);
    layer2_outputs(2067) <= not (a xor b);
    layer2_outputs(2068) <= not b or a;
    layer2_outputs(2069) <= not b;
    layer2_outputs(2070) <= not b or a;
    layer2_outputs(2071) <= not b or a;
    layer2_outputs(2072) <= not b;
    layer2_outputs(2073) <= a;
    layer2_outputs(2074) <= a and b;
    layer2_outputs(2075) <= b and not a;
    layer2_outputs(2076) <= a and not b;
    layer2_outputs(2077) <= b;
    layer2_outputs(2078) <= a or b;
    layer2_outputs(2079) <= a;
    layer2_outputs(2080) <= not (a and b);
    layer2_outputs(2081) <= not b;
    layer2_outputs(2082) <= not (a xor b);
    layer2_outputs(2083) <= b and not a;
    layer2_outputs(2084) <= a;
    layer2_outputs(2085) <= not b or a;
    layer2_outputs(2086) <= not b;
    layer2_outputs(2087) <= a;
    layer2_outputs(2088) <= a and b;
    layer2_outputs(2089) <= not (a or b);
    layer2_outputs(2090) <= not b;
    layer2_outputs(2091) <= not b;
    layer2_outputs(2092) <= a;
    layer2_outputs(2093) <= 1'b1;
    layer2_outputs(2094) <= a xor b;
    layer2_outputs(2095) <= a;
    layer2_outputs(2096) <= not b or a;
    layer2_outputs(2097) <= b;
    layer2_outputs(2098) <= not (a xor b);
    layer2_outputs(2099) <= not a;
    layer2_outputs(2100) <= not a;
    layer2_outputs(2101) <= not a;
    layer2_outputs(2102) <= b;
    layer2_outputs(2103) <= not (a and b);
    layer2_outputs(2104) <= b;
    layer2_outputs(2105) <= not (a xor b);
    layer2_outputs(2106) <= a or b;
    layer2_outputs(2107) <= a xor b;
    layer2_outputs(2108) <= not (a and b);
    layer2_outputs(2109) <= b;
    layer2_outputs(2110) <= not b;
    layer2_outputs(2111) <= not (a and b);
    layer2_outputs(2112) <= a and not b;
    layer2_outputs(2113) <= a;
    layer2_outputs(2114) <= not b or a;
    layer2_outputs(2115) <= not a or b;
    layer2_outputs(2116) <= not (a or b);
    layer2_outputs(2117) <= not (a and b);
    layer2_outputs(2118) <= not (a or b);
    layer2_outputs(2119) <= not a or b;
    layer2_outputs(2120) <= not b;
    layer2_outputs(2121) <= a and b;
    layer2_outputs(2122) <= not (a and b);
    layer2_outputs(2123) <= a and not b;
    layer2_outputs(2124) <= a;
    layer2_outputs(2125) <= not b;
    layer2_outputs(2126) <= not (a or b);
    layer2_outputs(2127) <= not a;
    layer2_outputs(2128) <= a and not b;
    layer2_outputs(2129) <= a;
    layer2_outputs(2130) <= not b or a;
    layer2_outputs(2131) <= a and b;
    layer2_outputs(2132) <= not a;
    layer2_outputs(2133) <= a and b;
    layer2_outputs(2134) <= not (a and b);
    layer2_outputs(2135) <= a and not b;
    layer2_outputs(2136) <= b and not a;
    layer2_outputs(2137) <= not (a or b);
    layer2_outputs(2138) <= not (a xor b);
    layer2_outputs(2139) <= a xor b;
    layer2_outputs(2140) <= b and not a;
    layer2_outputs(2141) <= not a or b;
    layer2_outputs(2142) <= a and b;
    layer2_outputs(2143) <= a or b;
    layer2_outputs(2144) <= not b;
    layer2_outputs(2145) <= a;
    layer2_outputs(2146) <= not (a and b);
    layer2_outputs(2147) <= not a;
    layer2_outputs(2148) <= not b;
    layer2_outputs(2149) <= a or b;
    layer2_outputs(2150) <= not (a xor b);
    layer2_outputs(2151) <= a or b;
    layer2_outputs(2152) <= a;
    layer2_outputs(2153) <= a;
    layer2_outputs(2154) <= not b;
    layer2_outputs(2155) <= not a;
    layer2_outputs(2156) <= not b;
    layer2_outputs(2157) <= not a or b;
    layer2_outputs(2158) <= not (a or b);
    layer2_outputs(2159) <= not b;
    layer2_outputs(2160) <= a and not b;
    layer2_outputs(2161) <= a;
    layer2_outputs(2162) <= b;
    layer2_outputs(2163) <= a and not b;
    layer2_outputs(2164) <= not a or b;
    layer2_outputs(2165) <= a and b;
    layer2_outputs(2166) <= a and b;
    layer2_outputs(2167) <= a xor b;
    layer2_outputs(2168) <= not a;
    layer2_outputs(2169) <= not (a or b);
    layer2_outputs(2170) <= not a;
    layer2_outputs(2171) <= a or b;
    layer2_outputs(2172) <= a xor b;
    layer2_outputs(2173) <= a xor b;
    layer2_outputs(2174) <= a;
    layer2_outputs(2175) <= not b;
    layer2_outputs(2176) <= not b;
    layer2_outputs(2177) <= not (a xor b);
    layer2_outputs(2178) <= b;
    layer2_outputs(2179) <= not (a and b);
    layer2_outputs(2180) <= a or b;
    layer2_outputs(2181) <= not (a xor b);
    layer2_outputs(2182) <= a xor b;
    layer2_outputs(2183) <= b;
    layer2_outputs(2184) <= not (a or b);
    layer2_outputs(2185) <= not b;
    layer2_outputs(2186) <= a;
    layer2_outputs(2187) <= not a;
    layer2_outputs(2188) <= not a;
    layer2_outputs(2189) <= not a or b;
    layer2_outputs(2190) <= not (a xor b);
    layer2_outputs(2191) <= a and b;
    layer2_outputs(2192) <= a;
    layer2_outputs(2193) <= not b;
    layer2_outputs(2194) <= not b or a;
    layer2_outputs(2195) <= a or b;
    layer2_outputs(2196) <= not a;
    layer2_outputs(2197) <= a and not b;
    layer2_outputs(2198) <= not a or b;
    layer2_outputs(2199) <= b and not a;
    layer2_outputs(2200) <= not (a and b);
    layer2_outputs(2201) <= not b;
    layer2_outputs(2202) <= b;
    layer2_outputs(2203) <= a;
    layer2_outputs(2204) <= b;
    layer2_outputs(2205) <= not a;
    layer2_outputs(2206) <= a or b;
    layer2_outputs(2207) <= a and not b;
    layer2_outputs(2208) <= a and not b;
    layer2_outputs(2209) <= not a;
    layer2_outputs(2210) <= b;
    layer2_outputs(2211) <= b and not a;
    layer2_outputs(2212) <= a;
    layer2_outputs(2213) <= not b;
    layer2_outputs(2214) <= not a;
    layer2_outputs(2215) <= not a;
    layer2_outputs(2216) <= b;
    layer2_outputs(2217) <= a;
    layer2_outputs(2218) <= not a or b;
    layer2_outputs(2219) <= not (a or b);
    layer2_outputs(2220) <= not (a and b);
    layer2_outputs(2221) <= not (a xor b);
    layer2_outputs(2222) <= not a;
    layer2_outputs(2223) <= b;
    layer2_outputs(2224) <= a and b;
    layer2_outputs(2225) <= a and b;
    layer2_outputs(2226) <= a or b;
    layer2_outputs(2227) <= a xor b;
    layer2_outputs(2228) <= not a;
    layer2_outputs(2229) <= not b;
    layer2_outputs(2230) <= not b or a;
    layer2_outputs(2231) <= not (a or b);
    layer2_outputs(2232) <= a and not b;
    layer2_outputs(2233) <= not a or b;
    layer2_outputs(2234) <= not a;
    layer2_outputs(2235) <= not (a or b);
    layer2_outputs(2236) <= not b or a;
    layer2_outputs(2237) <= not a;
    layer2_outputs(2238) <= b;
    layer2_outputs(2239) <= not a;
    layer2_outputs(2240) <= not b or a;
    layer2_outputs(2241) <= not b;
    layer2_outputs(2242) <= a;
    layer2_outputs(2243) <= a and not b;
    layer2_outputs(2244) <= b;
    layer2_outputs(2245) <= not (a or b);
    layer2_outputs(2246) <= not (a xor b);
    layer2_outputs(2247) <= not a or b;
    layer2_outputs(2248) <= not (a or b);
    layer2_outputs(2249) <= not b;
    layer2_outputs(2250) <= b and not a;
    layer2_outputs(2251) <= a;
    layer2_outputs(2252) <= a;
    layer2_outputs(2253) <= not b;
    layer2_outputs(2254) <= not (a xor b);
    layer2_outputs(2255) <= not b;
    layer2_outputs(2256) <= b;
    layer2_outputs(2257) <= b;
    layer2_outputs(2258) <= not a;
    layer2_outputs(2259) <= not b or a;
    layer2_outputs(2260) <= not a;
    layer2_outputs(2261) <= not (a xor b);
    layer2_outputs(2262) <= not a;
    layer2_outputs(2263) <= a;
    layer2_outputs(2264) <= not a or b;
    layer2_outputs(2265) <= b and not a;
    layer2_outputs(2266) <= not b or a;
    layer2_outputs(2267) <= not a;
    layer2_outputs(2268) <= not b;
    layer2_outputs(2269) <= a xor b;
    layer2_outputs(2270) <= not b;
    layer2_outputs(2271) <= not (a xor b);
    layer2_outputs(2272) <= a xor b;
    layer2_outputs(2273) <= b and not a;
    layer2_outputs(2274) <= a;
    layer2_outputs(2275) <= not b or a;
    layer2_outputs(2276) <= b;
    layer2_outputs(2277) <= b and not a;
    layer2_outputs(2278) <= a and not b;
    layer2_outputs(2279) <= a;
    layer2_outputs(2280) <= a and not b;
    layer2_outputs(2281) <= not b;
    layer2_outputs(2282) <= b;
    layer2_outputs(2283) <= not (a or b);
    layer2_outputs(2284) <= b;
    layer2_outputs(2285) <= not a;
    layer2_outputs(2286) <= not (a xor b);
    layer2_outputs(2287) <= not a or b;
    layer2_outputs(2288) <= a;
    layer2_outputs(2289) <= a and not b;
    layer2_outputs(2290) <= not b or a;
    layer2_outputs(2291) <= a;
    layer2_outputs(2292) <= not (a xor b);
    layer2_outputs(2293) <= not b or a;
    layer2_outputs(2294) <= b;
    layer2_outputs(2295) <= not b or a;
    layer2_outputs(2296) <= not a or b;
    layer2_outputs(2297) <= not b;
    layer2_outputs(2298) <= not (a or b);
    layer2_outputs(2299) <= b and not a;
    layer2_outputs(2300) <= not a;
    layer2_outputs(2301) <= b;
    layer2_outputs(2302) <= a xor b;
    layer2_outputs(2303) <= not b or a;
    layer2_outputs(2304) <= a;
    layer2_outputs(2305) <= not (a and b);
    layer2_outputs(2306) <= not b;
    layer2_outputs(2307) <= a xor b;
    layer2_outputs(2308) <= not b;
    layer2_outputs(2309) <= not (a and b);
    layer2_outputs(2310) <= a xor b;
    layer2_outputs(2311) <= b and not a;
    layer2_outputs(2312) <= not b;
    layer2_outputs(2313) <= a or b;
    layer2_outputs(2314) <= b and not a;
    layer2_outputs(2315) <= a and not b;
    layer2_outputs(2316) <= not b;
    layer2_outputs(2317) <= not a;
    layer2_outputs(2318) <= not b;
    layer2_outputs(2319) <= b;
    layer2_outputs(2320) <= not b;
    layer2_outputs(2321) <= a and not b;
    layer2_outputs(2322) <= a and b;
    layer2_outputs(2323) <= not b or a;
    layer2_outputs(2324) <= not b or a;
    layer2_outputs(2325) <= not b;
    layer2_outputs(2326) <= not b or a;
    layer2_outputs(2327) <= b and not a;
    layer2_outputs(2328) <= not a or b;
    layer2_outputs(2329) <= b;
    layer2_outputs(2330) <= not b;
    layer2_outputs(2331) <= not (a xor b);
    layer2_outputs(2332) <= not a;
    layer2_outputs(2333) <= not b;
    layer2_outputs(2334) <= b;
    layer2_outputs(2335) <= a;
    layer2_outputs(2336) <= not (a xor b);
    layer2_outputs(2337) <= a xor b;
    layer2_outputs(2338) <= a xor b;
    layer2_outputs(2339) <= not a or b;
    layer2_outputs(2340) <= a;
    layer2_outputs(2341) <= not b;
    layer2_outputs(2342) <= a or b;
    layer2_outputs(2343) <= not (a and b);
    layer2_outputs(2344) <= a and b;
    layer2_outputs(2345) <= 1'b1;
    layer2_outputs(2346) <= not b;
    layer2_outputs(2347) <= a and b;
    layer2_outputs(2348) <= not b;
    layer2_outputs(2349) <= a and b;
    layer2_outputs(2350) <= not (a xor b);
    layer2_outputs(2351) <= a;
    layer2_outputs(2352) <= a;
    layer2_outputs(2353) <= not a;
    layer2_outputs(2354) <= not (a xor b);
    layer2_outputs(2355) <= a and not b;
    layer2_outputs(2356) <= a or b;
    layer2_outputs(2357) <= not b;
    layer2_outputs(2358) <= b;
    layer2_outputs(2359) <= not (a xor b);
    layer2_outputs(2360) <= b;
    layer2_outputs(2361) <= not a;
    layer2_outputs(2362) <= a and not b;
    layer2_outputs(2363) <= not (a or b);
    layer2_outputs(2364) <= not b;
    layer2_outputs(2365) <= not b or a;
    layer2_outputs(2366) <= not a;
    layer2_outputs(2367) <= b;
    layer2_outputs(2368) <= not (a or b);
    layer2_outputs(2369) <= not a;
    layer2_outputs(2370) <= not b;
    layer2_outputs(2371) <= b and not a;
    layer2_outputs(2372) <= not (a xor b);
    layer2_outputs(2373) <= b and not a;
    layer2_outputs(2374) <= b;
    layer2_outputs(2375) <= not b or a;
    layer2_outputs(2376) <= b;
    layer2_outputs(2377) <= not a or b;
    layer2_outputs(2378) <= b;
    layer2_outputs(2379) <= a;
    layer2_outputs(2380) <= a;
    layer2_outputs(2381) <= a and not b;
    layer2_outputs(2382) <= a xor b;
    layer2_outputs(2383) <= a or b;
    layer2_outputs(2384) <= not (a and b);
    layer2_outputs(2385) <= not a;
    layer2_outputs(2386) <= not b;
    layer2_outputs(2387) <= not a;
    layer2_outputs(2388) <= not a or b;
    layer2_outputs(2389) <= not (a or b);
    layer2_outputs(2390) <= not (a and b);
    layer2_outputs(2391) <= not a;
    layer2_outputs(2392) <= not a;
    layer2_outputs(2393) <= not a or b;
    layer2_outputs(2394) <= b;
    layer2_outputs(2395) <= not (a and b);
    layer2_outputs(2396) <= a and b;
    layer2_outputs(2397) <= a xor b;
    layer2_outputs(2398) <= not b;
    layer2_outputs(2399) <= not b or a;
    layer2_outputs(2400) <= b;
    layer2_outputs(2401) <= not (a and b);
    layer2_outputs(2402) <= not a;
    layer2_outputs(2403) <= b;
    layer2_outputs(2404) <= a;
    layer2_outputs(2405) <= not b or a;
    layer2_outputs(2406) <= a and b;
    layer2_outputs(2407) <= not a;
    layer2_outputs(2408) <= not a;
    layer2_outputs(2409) <= not a;
    layer2_outputs(2410) <= a;
    layer2_outputs(2411) <= not (a or b);
    layer2_outputs(2412) <= not (a or b);
    layer2_outputs(2413) <= not b;
    layer2_outputs(2414) <= not a or b;
    layer2_outputs(2415) <= a and not b;
    layer2_outputs(2416) <= not b;
    layer2_outputs(2417) <= a and not b;
    layer2_outputs(2418) <= not (a or b);
    layer2_outputs(2419) <= not (a and b);
    layer2_outputs(2420) <= not a;
    layer2_outputs(2421) <= not a;
    layer2_outputs(2422) <= a and b;
    layer2_outputs(2423) <= not (a or b);
    layer2_outputs(2424) <= b;
    layer2_outputs(2425) <= not b or a;
    layer2_outputs(2426) <= not b or a;
    layer2_outputs(2427) <= a;
    layer2_outputs(2428) <= a or b;
    layer2_outputs(2429) <= not a or b;
    layer2_outputs(2430) <= a and not b;
    layer2_outputs(2431) <= not a;
    layer2_outputs(2432) <= b and not a;
    layer2_outputs(2433) <= not a;
    layer2_outputs(2434) <= a and not b;
    layer2_outputs(2435) <= b;
    layer2_outputs(2436) <= a;
    layer2_outputs(2437) <= a;
    layer2_outputs(2438) <= b;
    layer2_outputs(2439) <= not a or b;
    layer2_outputs(2440) <= not a;
    layer2_outputs(2441) <= not b;
    layer2_outputs(2442) <= b;
    layer2_outputs(2443) <= not b;
    layer2_outputs(2444) <= not (a or b);
    layer2_outputs(2445) <= a xor b;
    layer2_outputs(2446) <= a xor b;
    layer2_outputs(2447) <= a or b;
    layer2_outputs(2448) <= not a;
    layer2_outputs(2449) <= a and b;
    layer2_outputs(2450) <= b and not a;
    layer2_outputs(2451) <= a and b;
    layer2_outputs(2452) <= not b or a;
    layer2_outputs(2453) <= not (a and b);
    layer2_outputs(2454) <= not b or a;
    layer2_outputs(2455) <= not a or b;
    layer2_outputs(2456) <= not (a or b);
    layer2_outputs(2457) <= a and not b;
    layer2_outputs(2458) <= not a;
    layer2_outputs(2459) <= not b;
    layer2_outputs(2460) <= not a;
    layer2_outputs(2461) <= a;
    layer2_outputs(2462) <= b and not a;
    layer2_outputs(2463) <= a;
    layer2_outputs(2464) <= b and not a;
    layer2_outputs(2465) <= not b;
    layer2_outputs(2466) <= not a or b;
    layer2_outputs(2467) <= not b;
    layer2_outputs(2468) <= a;
    layer2_outputs(2469) <= not b;
    layer2_outputs(2470) <= a;
    layer2_outputs(2471) <= b;
    layer2_outputs(2472) <= not (a and b);
    layer2_outputs(2473) <= not b;
    layer2_outputs(2474) <= not b;
    layer2_outputs(2475) <= a and b;
    layer2_outputs(2476) <= not b;
    layer2_outputs(2477) <= b;
    layer2_outputs(2478) <= not a;
    layer2_outputs(2479) <= a;
    layer2_outputs(2480) <= a;
    layer2_outputs(2481) <= 1'b1;
    layer2_outputs(2482) <= not a;
    layer2_outputs(2483) <= not (a or b);
    layer2_outputs(2484) <= not (a and b);
    layer2_outputs(2485) <= not (a or b);
    layer2_outputs(2486) <= a and not b;
    layer2_outputs(2487) <= a and not b;
    layer2_outputs(2488) <= not a;
    layer2_outputs(2489) <= not b or a;
    layer2_outputs(2490) <= not (a or b);
    layer2_outputs(2491) <= a or b;
    layer2_outputs(2492) <= b and not a;
    layer2_outputs(2493) <= not a;
    layer2_outputs(2494) <= not b;
    layer2_outputs(2495) <= a and b;
    layer2_outputs(2496) <= a and b;
    layer2_outputs(2497) <= not b or a;
    layer2_outputs(2498) <= not b;
    layer2_outputs(2499) <= not b;
    layer2_outputs(2500) <= a;
    layer2_outputs(2501) <= b and not a;
    layer2_outputs(2502) <= a and not b;
    layer2_outputs(2503) <= not a;
    layer2_outputs(2504) <= not b;
    layer2_outputs(2505) <= b;
    layer2_outputs(2506) <= a and b;
    layer2_outputs(2507) <= not (a or b);
    layer2_outputs(2508) <= not a or b;
    layer2_outputs(2509) <= a;
    layer2_outputs(2510) <= not (a or b);
    layer2_outputs(2511) <= not a or b;
    layer2_outputs(2512) <= a and b;
    layer2_outputs(2513) <= b;
    layer2_outputs(2514) <= b and not a;
    layer2_outputs(2515) <= not (a xor b);
    layer2_outputs(2516) <= a xor b;
    layer2_outputs(2517) <= b;
    layer2_outputs(2518) <= b;
    layer2_outputs(2519) <= not b or a;
    layer2_outputs(2520) <= b and not a;
    layer2_outputs(2521) <= not b;
    layer2_outputs(2522) <= not b;
    layer2_outputs(2523) <= not (a and b);
    layer2_outputs(2524) <= not a or b;
    layer2_outputs(2525) <= not (a or b);
    layer2_outputs(2526) <= not b;
    layer2_outputs(2527) <= not (a and b);
    layer2_outputs(2528) <= a or b;
    layer2_outputs(2529) <= a xor b;
    layer2_outputs(2530) <= a xor b;
    layer2_outputs(2531) <= a xor b;
    layer2_outputs(2532) <= not a;
    layer2_outputs(2533) <= not b or a;
    layer2_outputs(2534) <= not a or b;
    layer2_outputs(2535) <= not a;
    layer2_outputs(2536) <= not (a or b);
    layer2_outputs(2537) <= not (a xor b);
    layer2_outputs(2538) <= not b or a;
    layer2_outputs(2539) <= not b;
    layer2_outputs(2540) <= a or b;
    layer2_outputs(2541) <= a or b;
    layer2_outputs(2542) <= a and b;
    layer2_outputs(2543) <= not a or b;
    layer2_outputs(2544) <= not a;
    layer2_outputs(2545) <= a or b;
    layer2_outputs(2546) <= not a;
    layer2_outputs(2547) <= not a;
    layer2_outputs(2548) <= a;
    layer2_outputs(2549) <= b;
    layer2_outputs(2550) <= not a;
    layer2_outputs(2551) <= not a;
    layer2_outputs(2552) <= b;
    layer2_outputs(2553) <= a and not b;
    layer2_outputs(2554) <= a and not b;
    layer2_outputs(2555) <= a xor b;
    layer2_outputs(2556) <= a;
    layer2_outputs(2557) <= b;
    layer2_outputs(2558) <= not (a and b);
    layer2_outputs(2559) <= not b;
    layer2_outputs(2560) <= not b or a;
    layer2_outputs(2561) <= a xor b;
    layer2_outputs(2562) <= not a;
    layer2_outputs(2563) <= a or b;
    layer2_outputs(2564) <= not (a and b);
    layer2_outputs(2565) <= not (a xor b);
    layer2_outputs(2566) <= not (a xor b);
    layer2_outputs(2567) <= a xor b;
    layer2_outputs(2568) <= not a;
    layer2_outputs(2569) <= not (a or b);
    layer2_outputs(2570) <= not a;
    layer2_outputs(2571) <= not a or b;
    layer2_outputs(2572) <= a and b;
    layer2_outputs(2573) <= not a;
    layer2_outputs(2574) <= not (a and b);
    layer2_outputs(2575) <= not (a xor b);
    layer2_outputs(2576) <= not b;
    layer2_outputs(2577) <= not (a or b);
    layer2_outputs(2578) <= not (a or b);
    layer2_outputs(2579) <= not a;
    layer2_outputs(2580) <= not a or b;
    layer2_outputs(2581) <= a xor b;
    layer2_outputs(2582) <= not a;
    layer2_outputs(2583) <= not (a or b);
    layer2_outputs(2584) <= not b;
    layer2_outputs(2585) <= not (a and b);
    layer2_outputs(2586) <= a;
    layer2_outputs(2587) <= not b or a;
    layer2_outputs(2588) <= not (a xor b);
    layer2_outputs(2589) <= not b or a;
    layer2_outputs(2590) <= not b or a;
    layer2_outputs(2591) <= not (a and b);
    layer2_outputs(2592) <= not b;
    layer2_outputs(2593) <= not a;
    layer2_outputs(2594) <= not b;
    layer2_outputs(2595) <= b;
    layer2_outputs(2596) <= not b;
    layer2_outputs(2597) <= not (a or b);
    layer2_outputs(2598) <= b;
    layer2_outputs(2599) <= a;
    layer2_outputs(2600) <= b;
    layer2_outputs(2601) <= not (a xor b);
    layer2_outputs(2602) <= a;
    layer2_outputs(2603) <= not (a xor b);
    layer2_outputs(2604) <= b and not a;
    layer2_outputs(2605) <= a xor b;
    layer2_outputs(2606) <= a or b;
    layer2_outputs(2607) <= a and b;
    layer2_outputs(2608) <= b;
    layer2_outputs(2609) <= a and not b;
    layer2_outputs(2610) <= b;
    layer2_outputs(2611) <= not a or b;
    layer2_outputs(2612) <= a xor b;
    layer2_outputs(2613) <= not b;
    layer2_outputs(2614) <= not a;
    layer2_outputs(2615) <= not a or b;
    layer2_outputs(2616) <= b;
    layer2_outputs(2617) <= b;
    layer2_outputs(2618) <= a;
    layer2_outputs(2619) <= not (a xor b);
    layer2_outputs(2620) <= not (a or b);
    layer2_outputs(2621) <= b;
    layer2_outputs(2622) <= a xor b;
    layer2_outputs(2623) <= not (a or b);
    layer2_outputs(2624) <= not a;
    layer2_outputs(2625) <= a xor b;
    layer2_outputs(2626) <= a and b;
    layer2_outputs(2627) <= b and not a;
    layer2_outputs(2628) <= a or b;
    layer2_outputs(2629) <= not (a xor b);
    layer2_outputs(2630) <= b;
    layer2_outputs(2631) <= not b or a;
    layer2_outputs(2632) <= a and b;
    layer2_outputs(2633) <= not b;
    layer2_outputs(2634) <= b and not a;
    layer2_outputs(2635) <= b;
    layer2_outputs(2636) <= not (a xor b);
    layer2_outputs(2637) <= not b or a;
    layer2_outputs(2638) <= not (a xor b);
    layer2_outputs(2639) <= b;
    layer2_outputs(2640) <= not a;
    layer2_outputs(2641) <= a or b;
    layer2_outputs(2642) <= b and not a;
    layer2_outputs(2643) <= a or b;
    layer2_outputs(2644) <= a or b;
    layer2_outputs(2645) <= not (a xor b);
    layer2_outputs(2646) <= not a or b;
    layer2_outputs(2647) <= not (a or b);
    layer2_outputs(2648) <= not b;
    layer2_outputs(2649) <= not (a xor b);
    layer2_outputs(2650) <= not (a and b);
    layer2_outputs(2651) <= 1'b1;
    layer2_outputs(2652) <= not (a or b);
    layer2_outputs(2653) <= not (a xor b);
    layer2_outputs(2654) <= b;
    layer2_outputs(2655) <= not b;
    layer2_outputs(2656) <= not a or b;
    layer2_outputs(2657) <= not (a xor b);
    layer2_outputs(2658) <= not b;
    layer2_outputs(2659) <= b and not a;
    layer2_outputs(2660) <= not a;
    layer2_outputs(2661) <= not a or b;
    layer2_outputs(2662) <= b;
    layer2_outputs(2663) <= a;
    layer2_outputs(2664) <= a or b;
    layer2_outputs(2665) <= b;
    layer2_outputs(2666) <= a or b;
    layer2_outputs(2667) <= b and not a;
    layer2_outputs(2668) <= a;
    layer2_outputs(2669) <= not (a xor b);
    layer2_outputs(2670) <= not b;
    layer2_outputs(2671) <= a and not b;
    layer2_outputs(2672) <= a and b;
    layer2_outputs(2673) <= not (a or b);
    layer2_outputs(2674) <= not b;
    layer2_outputs(2675) <= not (a and b);
    layer2_outputs(2676) <= a xor b;
    layer2_outputs(2677) <= a and not b;
    layer2_outputs(2678) <= not (a and b);
    layer2_outputs(2679) <= a;
    layer2_outputs(2680) <= b;
    layer2_outputs(2681) <= not a;
    layer2_outputs(2682) <= not a;
    layer2_outputs(2683) <= a and not b;
    layer2_outputs(2684) <= a and b;
    layer2_outputs(2685) <= b;
    layer2_outputs(2686) <= not a;
    layer2_outputs(2687) <= b;
    layer2_outputs(2688) <= a;
    layer2_outputs(2689) <= a or b;
    layer2_outputs(2690) <= not (a or b);
    layer2_outputs(2691) <= a xor b;
    layer2_outputs(2692) <= not b or a;
    layer2_outputs(2693) <= not b;
    layer2_outputs(2694) <= not a;
    layer2_outputs(2695) <= not a;
    layer2_outputs(2696) <= b;
    layer2_outputs(2697) <= not a;
    layer2_outputs(2698) <= a and b;
    layer2_outputs(2699) <= a xor b;
    layer2_outputs(2700) <= not a;
    layer2_outputs(2701) <= a or b;
    layer2_outputs(2702) <= a or b;
    layer2_outputs(2703) <= not (a xor b);
    layer2_outputs(2704) <= not a or b;
    layer2_outputs(2705) <= a and b;
    layer2_outputs(2706) <= not (a and b);
    layer2_outputs(2707) <= not a;
    layer2_outputs(2708) <= not a;
    layer2_outputs(2709) <= not a or b;
    layer2_outputs(2710) <= not a or b;
    layer2_outputs(2711) <= a and not b;
    layer2_outputs(2712) <= not (a or b);
    layer2_outputs(2713) <= not (a xor b);
    layer2_outputs(2714) <= b;
    layer2_outputs(2715) <= not b;
    layer2_outputs(2716) <= not b;
    layer2_outputs(2717) <= a xor b;
    layer2_outputs(2718) <= a and b;
    layer2_outputs(2719) <= a xor b;
    layer2_outputs(2720) <= not (a xor b);
    layer2_outputs(2721) <= not (a or b);
    layer2_outputs(2722) <= b and not a;
    layer2_outputs(2723) <= not (a xor b);
    layer2_outputs(2724) <= not b;
    layer2_outputs(2725) <= b and not a;
    layer2_outputs(2726) <= b and not a;
    layer2_outputs(2727) <= 1'b0;
    layer2_outputs(2728) <= not (a and b);
    layer2_outputs(2729) <= a and not b;
    layer2_outputs(2730) <= a and b;
    layer2_outputs(2731) <= b;
    layer2_outputs(2732) <= not a or b;
    layer2_outputs(2733) <= not (a or b);
    layer2_outputs(2734) <= b;
    layer2_outputs(2735) <= a or b;
    layer2_outputs(2736) <= b;
    layer2_outputs(2737) <= a or b;
    layer2_outputs(2738) <= a or b;
    layer2_outputs(2739) <= not b or a;
    layer2_outputs(2740) <= a xor b;
    layer2_outputs(2741) <= not a;
    layer2_outputs(2742) <= a and b;
    layer2_outputs(2743) <= a or b;
    layer2_outputs(2744) <= b;
    layer2_outputs(2745) <= not a;
    layer2_outputs(2746) <= not b;
    layer2_outputs(2747) <= not (a xor b);
    layer2_outputs(2748) <= not (a or b);
    layer2_outputs(2749) <= not b or a;
    layer2_outputs(2750) <= a or b;
    layer2_outputs(2751) <= not a or b;
    layer2_outputs(2752) <= not a or b;
    layer2_outputs(2753) <= not (a xor b);
    layer2_outputs(2754) <= a or b;
    layer2_outputs(2755) <= not (a and b);
    layer2_outputs(2756) <= a;
    layer2_outputs(2757) <= a;
    layer2_outputs(2758) <= not a;
    layer2_outputs(2759) <= not a;
    layer2_outputs(2760) <= not a;
    layer2_outputs(2761) <= not b;
    layer2_outputs(2762) <= a and not b;
    layer2_outputs(2763) <= not a;
    layer2_outputs(2764) <= not a;
    layer2_outputs(2765) <= a xor b;
    layer2_outputs(2766) <= a or b;
    layer2_outputs(2767) <= b;
    layer2_outputs(2768) <= not b;
    layer2_outputs(2769) <= not a;
    layer2_outputs(2770) <= a and not b;
    layer2_outputs(2771) <= not a or b;
    layer2_outputs(2772) <= a;
    layer2_outputs(2773) <= not (a and b);
    layer2_outputs(2774) <= a or b;
    layer2_outputs(2775) <= not a or b;
    layer2_outputs(2776) <= not b or a;
    layer2_outputs(2777) <= b and not a;
    layer2_outputs(2778) <= not (a xor b);
    layer2_outputs(2779) <= a or b;
    layer2_outputs(2780) <= not a;
    layer2_outputs(2781) <= not a;
    layer2_outputs(2782) <= not b;
    layer2_outputs(2783) <= not (a and b);
    layer2_outputs(2784) <= a and b;
    layer2_outputs(2785) <= a and not b;
    layer2_outputs(2786) <= not b or a;
    layer2_outputs(2787) <= a xor b;
    layer2_outputs(2788) <= not b;
    layer2_outputs(2789) <= b and not a;
    layer2_outputs(2790) <= b;
    layer2_outputs(2791) <= a;
    layer2_outputs(2792) <= a;
    layer2_outputs(2793) <= a xor b;
    layer2_outputs(2794) <= a;
    layer2_outputs(2795) <= not a or b;
    layer2_outputs(2796) <= not (a xor b);
    layer2_outputs(2797) <= a;
    layer2_outputs(2798) <= not b;
    layer2_outputs(2799) <= b and not a;
    layer2_outputs(2800) <= not (a xor b);
    layer2_outputs(2801) <= a;
    layer2_outputs(2802) <= b;
    layer2_outputs(2803) <= a;
    layer2_outputs(2804) <= b and not a;
    layer2_outputs(2805) <= not a;
    layer2_outputs(2806) <= a or b;
    layer2_outputs(2807) <= not (a and b);
    layer2_outputs(2808) <= a;
    layer2_outputs(2809) <= not (a or b);
    layer2_outputs(2810) <= b;
    layer2_outputs(2811) <= a;
    layer2_outputs(2812) <= a;
    layer2_outputs(2813) <= a xor b;
    layer2_outputs(2814) <= not b;
    layer2_outputs(2815) <= a xor b;
    layer2_outputs(2816) <= not b;
    layer2_outputs(2817) <= a xor b;
    layer2_outputs(2818) <= not a or b;
    layer2_outputs(2819) <= not (a xor b);
    layer2_outputs(2820) <= not (a or b);
    layer2_outputs(2821) <= a xor b;
    layer2_outputs(2822) <= not a;
    layer2_outputs(2823) <= not b;
    layer2_outputs(2824) <= b;
    layer2_outputs(2825) <= not b;
    layer2_outputs(2826) <= a or b;
    layer2_outputs(2827) <= not (a and b);
    layer2_outputs(2828) <= 1'b0;
    layer2_outputs(2829) <= a;
    layer2_outputs(2830) <= b;
    layer2_outputs(2831) <= a or b;
    layer2_outputs(2832) <= a;
    layer2_outputs(2833) <= not b;
    layer2_outputs(2834) <= a xor b;
    layer2_outputs(2835) <= b;
    layer2_outputs(2836) <= not a or b;
    layer2_outputs(2837) <= not (a xor b);
    layer2_outputs(2838) <= a;
    layer2_outputs(2839) <= b and not a;
    layer2_outputs(2840) <= not a;
    layer2_outputs(2841) <= a;
    layer2_outputs(2842) <= not b;
    layer2_outputs(2843) <= b;
    layer2_outputs(2844) <= a xor b;
    layer2_outputs(2845) <= 1'b0;
    layer2_outputs(2846) <= a;
    layer2_outputs(2847) <= b;
    layer2_outputs(2848) <= not (a and b);
    layer2_outputs(2849) <= b;
    layer2_outputs(2850) <= not (a and b);
    layer2_outputs(2851) <= not (a or b);
    layer2_outputs(2852) <= not a;
    layer2_outputs(2853) <= a and not b;
    layer2_outputs(2854) <= a and not b;
    layer2_outputs(2855) <= not a or b;
    layer2_outputs(2856) <= a or b;
    layer2_outputs(2857) <= not (a and b);
    layer2_outputs(2858) <= a or b;
    layer2_outputs(2859) <= b;
    layer2_outputs(2860) <= not (a and b);
    layer2_outputs(2861) <= not a;
    layer2_outputs(2862) <= a or b;
    layer2_outputs(2863) <= not b or a;
    layer2_outputs(2864) <= b;
    layer2_outputs(2865) <= b;
    layer2_outputs(2866) <= not (a or b);
    layer2_outputs(2867) <= a xor b;
    layer2_outputs(2868) <= a;
    layer2_outputs(2869) <= a;
    layer2_outputs(2870) <= not b or a;
    layer2_outputs(2871) <= not b;
    layer2_outputs(2872) <= not a;
    layer2_outputs(2873) <= a or b;
    layer2_outputs(2874) <= not b;
    layer2_outputs(2875) <= not a or b;
    layer2_outputs(2876) <= a xor b;
    layer2_outputs(2877) <= b and not a;
    layer2_outputs(2878) <= not (a xor b);
    layer2_outputs(2879) <= not (a and b);
    layer2_outputs(2880) <= not (a and b);
    layer2_outputs(2881) <= not a or b;
    layer2_outputs(2882) <= not a;
    layer2_outputs(2883) <= b;
    layer2_outputs(2884) <= a;
    layer2_outputs(2885) <= b;
    layer2_outputs(2886) <= a or b;
    layer2_outputs(2887) <= not b or a;
    layer2_outputs(2888) <= not (a or b);
    layer2_outputs(2889) <= not b or a;
    layer2_outputs(2890) <= not a or b;
    layer2_outputs(2891) <= a xor b;
    layer2_outputs(2892) <= not b or a;
    layer2_outputs(2893) <= not b or a;
    layer2_outputs(2894) <= not b;
    layer2_outputs(2895) <= a and not b;
    layer2_outputs(2896) <= a xor b;
    layer2_outputs(2897) <= a or b;
    layer2_outputs(2898) <= not a;
    layer2_outputs(2899) <= not b;
    layer2_outputs(2900) <= not (a or b);
    layer2_outputs(2901) <= not (a xor b);
    layer2_outputs(2902) <= not a or b;
    layer2_outputs(2903) <= not b;
    layer2_outputs(2904) <= not b;
    layer2_outputs(2905) <= a and not b;
    layer2_outputs(2906) <= not (a or b);
    layer2_outputs(2907) <= not a;
    layer2_outputs(2908) <= not a or b;
    layer2_outputs(2909) <= a xor b;
    layer2_outputs(2910) <= not a;
    layer2_outputs(2911) <= a and b;
    layer2_outputs(2912) <= a xor b;
    layer2_outputs(2913) <= a and b;
    layer2_outputs(2914) <= not (a xor b);
    layer2_outputs(2915) <= b;
    layer2_outputs(2916) <= a xor b;
    layer2_outputs(2917) <= not (a or b);
    layer2_outputs(2918) <= a xor b;
    layer2_outputs(2919) <= not a;
    layer2_outputs(2920) <= b and not a;
    layer2_outputs(2921) <= a or b;
    layer2_outputs(2922) <= not a;
    layer2_outputs(2923) <= not a;
    layer2_outputs(2924) <= a and not b;
    layer2_outputs(2925) <= not (a or b);
    layer2_outputs(2926) <= not a or b;
    layer2_outputs(2927) <= a or b;
    layer2_outputs(2928) <= not a;
    layer2_outputs(2929) <= a or b;
    layer2_outputs(2930) <= not b;
    layer2_outputs(2931) <= not a;
    layer2_outputs(2932) <= a and not b;
    layer2_outputs(2933) <= not a;
    layer2_outputs(2934) <= not (a xor b);
    layer2_outputs(2935) <= not a;
    layer2_outputs(2936) <= not (a xor b);
    layer2_outputs(2937) <= a and b;
    layer2_outputs(2938) <= b;
    layer2_outputs(2939) <= not (a xor b);
    layer2_outputs(2940) <= a;
    layer2_outputs(2941) <= a and not b;
    layer2_outputs(2942) <= b and not a;
    layer2_outputs(2943) <= not (a or b);
    layer2_outputs(2944) <= not (a or b);
    layer2_outputs(2945) <= not a;
    layer2_outputs(2946) <= not b;
    layer2_outputs(2947) <= a and not b;
    layer2_outputs(2948) <= a or b;
    layer2_outputs(2949) <= not b or a;
    layer2_outputs(2950) <= a;
    layer2_outputs(2951) <= a and b;
    layer2_outputs(2952) <= a;
    layer2_outputs(2953) <= b;
    layer2_outputs(2954) <= not b or a;
    layer2_outputs(2955) <= a;
    layer2_outputs(2956) <= a and b;
    layer2_outputs(2957) <= a and b;
    layer2_outputs(2958) <= b and not a;
    layer2_outputs(2959) <= not a;
    layer2_outputs(2960) <= b;
    layer2_outputs(2961) <= a and not b;
    layer2_outputs(2962) <= not a;
    layer2_outputs(2963) <= a xor b;
    layer2_outputs(2964) <= not (a or b);
    layer2_outputs(2965) <= not a;
    layer2_outputs(2966) <= a and not b;
    layer2_outputs(2967) <= a;
    layer2_outputs(2968) <= a;
    layer2_outputs(2969) <= not b;
    layer2_outputs(2970) <= a;
    layer2_outputs(2971) <= not b;
    layer2_outputs(2972) <= not a or b;
    layer2_outputs(2973) <= not b or a;
    layer2_outputs(2974) <= not a or b;
    layer2_outputs(2975) <= a;
    layer2_outputs(2976) <= not a;
    layer2_outputs(2977) <= b;
    layer2_outputs(2978) <= a and b;
    layer2_outputs(2979) <= not b;
    layer2_outputs(2980) <= a xor b;
    layer2_outputs(2981) <= a and b;
    layer2_outputs(2982) <= a;
    layer2_outputs(2983) <= a and b;
    layer2_outputs(2984) <= b and not a;
    layer2_outputs(2985) <= not b or a;
    layer2_outputs(2986) <= not a or b;
    layer2_outputs(2987) <= a or b;
    layer2_outputs(2988) <= not b;
    layer2_outputs(2989) <= not (a xor b);
    layer2_outputs(2990) <= a or b;
    layer2_outputs(2991) <= not b;
    layer2_outputs(2992) <= a and b;
    layer2_outputs(2993) <= not a or b;
    layer2_outputs(2994) <= not b or a;
    layer2_outputs(2995) <= not b;
    layer2_outputs(2996) <= b and not a;
    layer2_outputs(2997) <= not a;
    layer2_outputs(2998) <= not a or b;
    layer2_outputs(2999) <= not (a xor b);
    layer2_outputs(3000) <= a;
    layer2_outputs(3001) <= a and not b;
    layer2_outputs(3002) <= not b;
    layer2_outputs(3003) <= not b or a;
    layer2_outputs(3004) <= a and not b;
    layer2_outputs(3005) <= b and not a;
    layer2_outputs(3006) <= not b;
    layer2_outputs(3007) <= not (a xor b);
    layer2_outputs(3008) <= not b;
    layer2_outputs(3009) <= b;
    layer2_outputs(3010) <= not a;
    layer2_outputs(3011) <= not (a or b);
    layer2_outputs(3012) <= not (a or b);
    layer2_outputs(3013) <= not a or b;
    layer2_outputs(3014) <= not b;
    layer2_outputs(3015) <= not a;
    layer2_outputs(3016) <= not b or a;
    layer2_outputs(3017) <= not b or a;
    layer2_outputs(3018) <= a and b;
    layer2_outputs(3019) <= not a;
    layer2_outputs(3020) <= a and b;
    layer2_outputs(3021) <= a xor b;
    layer2_outputs(3022) <= not a;
    layer2_outputs(3023) <= not a;
    layer2_outputs(3024) <= a xor b;
    layer2_outputs(3025) <= a;
    layer2_outputs(3026) <= a or b;
    layer2_outputs(3027) <= not (a and b);
    layer2_outputs(3028) <= a;
    layer2_outputs(3029) <= not (a or b);
    layer2_outputs(3030) <= not (a or b);
    layer2_outputs(3031) <= not a or b;
    layer2_outputs(3032) <= a;
    layer2_outputs(3033) <= not (a and b);
    layer2_outputs(3034) <= a;
    layer2_outputs(3035) <= a and not b;
    layer2_outputs(3036) <= a;
    layer2_outputs(3037) <= not (a xor b);
    layer2_outputs(3038) <= not (a or b);
    layer2_outputs(3039) <= not a or b;
    layer2_outputs(3040) <= a or b;
    layer2_outputs(3041) <= not a or b;
    layer2_outputs(3042) <= not (a and b);
    layer2_outputs(3043) <= not a or b;
    layer2_outputs(3044) <= not b or a;
    layer2_outputs(3045) <= not (a or b);
    layer2_outputs(3046) <= a or b;
    layer2_outputs(3047) <= a;
    layer2_outputs(3048) <= b;
    layer2_outputs(3049) <= not (a xor b);
    layer2_outputs(3050) <= not b;
    layer2_outputs(3051) <= not b or a;
    layer2_outputs(3052) <= b and not a;
    layer2_outputs(3053) <= not b;
    layer2_outputs(3054) <= a xor b;
    layer2_outputs(3055) <= a and not b;
    layer2_outputs(3056) <= not (a xor b);
    layer2_outputs(3057) <= b and not a;
    layer2_outputs(3058) <= not (a xor b);
    layer2_outputs(3059) <= a and not b;
    layer2_outputs(3060) <= b;
    layer2_outputs(3061) <= not (a and b);
    layer2_outputs(3062) <= b and not a;
    layer2_outputs(3063) <= not b or a;
    layer2_outputs(3064) <= not a;
    layer2_outputs(3065) <= not (a xor b);
    layer2_outputs(3066) <= a;
    layer2_outputs(3067) <= not (a or b);
    layer2_outputs(3068) <= not a or b;
    layer2_outputs(3069) <= a xor b;
    layer2_outputs(3070) <= not (a xor b);
    layer2_outputs(3071) <= not a;
    layer2_outputs(3072) <= not (a or b);
    layer2_outputs(3073) <= a xor b;
    layer2_outputs(3074) <= a xor b;
    layer2_outputs(3075) <= not a;
    layer2_outputs(3076) <= not a;
    layer2_outputs(3077) <= not a;
    layer2_outputs(3078) <= a;
    layer2_outputs(3079) <= not (a and b);
    layer2_outputs(3080) <= a;
    layer2_outputs(3081) <= a xor b;
    layer2_outputs(3082) <= not b;
    layer2_outputs(3083) <= not a or b;
    layer2_outputs(3084) <= not (a and b);
    layer2_outputs(3085) <= not (a or b);
    layer2_outputs(3086) <= b;
    layer2_outputs(3087) <= not (a xor b);
    layer2_outputs(3088) <= a xor b;
    layer2_outputs(3089) <= not b;
    layer2_outputs(3090) <= not (a or b);
    layer2_outputs(3091) <= a xor b;
    layer2_outputs(3092) <= not (a xor b);
    layer2_outputs(3093) <= not b or a;
    layer2_outputs(3094) <= a;
    layer2_outputs(3095) <= not a;
    layer2_outputs(3096) <= a xor b;
    layer2_outputs(3097) <= not b or a;
    layer2_outputs(3098) <= a;
    layer2_outputs(3099) <= a and not b;
    layer2_outputs(3100) <= b;
    layer2_outputs(3101) <= b and not a;
    layer2_outputs(3102) <= not b;
    layer2_outputs(3103) <= a xor b;
    layer2_outputs(3104) <= a xor b;
    layer2_outputs(3105) <= not a;
    layer2_outputs(3106) <= a;
    layer2_outputs(3107) <= not (a and b);
    layer2_outputs(3108) <= not a;
    layer2_outputs(3109) <= not (a and b);
    layer2_outputs(3110) <= a and b;
    layer2_outputs(3111) <= not b or a;
    layer2_outputs(3112) <= a and not b;
    layer2_outputs(3113) <= b;
    layer2_outputs(3114) <= a and not b;
    layer2_outputs(3115) <= not (a xor b);
    layer2_outputs(3116) <= not (a or b);
    layer2_outputs(3117) <= a xor b;
    layer2_outputs(3118) <= a;
    layer2_outputs(3119) <= a or b;
    layer2_outputs(3120) <= a or b;
    layer2_outputs(3121) <= not (a xor b);
    layer2_outputs(3122) <= not (a or b);
    layer2_outputs(3123) <= a;
    layer2_outputs(3124) <= not b or a;
    layer2_outputs(3125) <= b;
    layer2_outputs(3126) <= a;
    layer2_outputs(3127) <= a or b;
    layer2_outputs(3128) <= not a or b;
    layer2_outputs(3129) <= a or b;
    layer2_outputs(3130) <= not a;
    layer2_outputs(3131) <= a or b;
    layer2_outputs(3132) <= not a or b;
    layer2_outputs(3133) <= a;
    layer2_outputs(3134) <= a xor b;
    layer2_outputs(3135) <= not b or a;
    layer2_outputs(3136) <= not (a and b);
    layer2_outputs(3137) <= b;
    layer2_outputs(3138) <= b and not a;
    layer2_outputs(3139) <= a;
    layer2_outputs(3140) <= a;
    layer2_outputs(3141) <= a and not b;
    layer2_outputs(3142) <= not (a xor b);
    layer2_outputs(3143) <= not (a or b);
    layer2_outputs(3144) <= b and not a;
    layer2_outputs(3145) <= b and not a;
    layer2_outputs(3146) <= not b or a;
    layer2_outputs(3147) <= b;
    layer2_outputs(3148) <= b;
    layer2_outputs(3149) <= not (a and b);
    layer2_outputs(3150) <= not b;
    layer2_outputs(3151) <= not (a xor b);
    layer2_outputs(3152) <= not b;
    layer2_outputs(3153) <= a or b;
    layer2_outputs(3154) <= b and not a;
    layer2_outputs(3155) <= 1'b1;
    layer2_outputs(3156) <= not b or a;
    layer2_outputs(3157) <= b;
    layer2_outputs(3158) <= not b or a;
    layer2_outputs(3159) <= b;
    layer2_outputs(3160) <= not a or b;
    layer2_outputs(3161) <= a and b;
    layer2_outputs(3162) <= not (a and b);
    layer2_outputs(3163) <= not a;
    layer2_outputs(3164) <= not (a or b);
    layer2_outputs(3165) <= a xor b;
    layer2_outputs(3166) <= a and b;
    layer2_outputs(3167) <= not a;
    layer2_outputs(3168) <= a;
    layer2_outputs(3169) <= not b or a;
    layer2_outputs(3170) <= not a;
    layer2_outputs(3171) <= not a;
    layer2_outputs(3172) <= a;
    layer2_outputs(3173) <= not b;
    layer2_outputs(3174) <= a or b;
    layer2_outputs(3175) <= a and not b;
    layer2_outputs(3176) <= not a or b;
    layer2_outputs(3177) <= a;
    layer2_outputs(3178) <= a and b;
    layer2_outputs(3179) <= not b;
    layer2_outputs(3180) <= not a;
    layer2_outputs(3181) <= not a;
    layer2_outputs(3182) <= a and b;
    layer2_outputs(3183) <= not (a and b);
    layer2_outputs(3184) <= a and b;
    layer2_outputs(3185) <= b;
    layer2_outputs(3186) <= b;
    layer2_outputs(3187) <= a and b;
    layer2_outputs(3188) <= not (a xor b);
    layer2_outputs(3189) <= a and b;
    layer2_outputs(3190) <= a xor b;
    layer2_outputs(3191) <= a and b;
    layer2_outputs(3192) <= b and not a;
    layer2_outputs(3193) <= b and not a;
    layer2_outputs(3194) <= b;
    layer2_outputs(3195) <= a;
    layer2_outputs(3196) <= a and b;
    layer2_outputs(3197) <= not b or a;
    layer2_outputs(3198) <= a;
    layer2_outputs(3199) <= b;
    layer2_outputs(3200) <= not b;
    layer2_outputs(3201) <= a xor b;
    layer2_outputs(3202) <= not a;
    layer2_outputs(3203) <= b and not a;
    layer2_outputs(3204) <= not a or b;
    layer2_outputs(3205) <= not (a and b);
    layer2_outputs(3206) <= a and not b;
    layer2_outputs(3207) <= not b;
    layer2_outputs(3208) <= a xor b;
    layer2_outputs(3209) <= a and not b;
    layer2_outputs(3210) <= not a;
    layer2_outputs(3211) <= not b;
    layer2_outputs(3212) <= a;
    layer2_outputs(3213) <= not (a xor b);
    layer2_outputs(3214) <= not a or b;
    layer2_outputs(3215) <= not a;
    layer2_outputs(3216) <= a xor b;
    layer2_outputs(3217) <= a;
    layer2_outputs(3218) <= a or b;
    layer2_outputs(3219) <= b;
    layer2_outputs(3220) <= not a;
    layer2_outputs(3221) <= a;
    layer2_outputs(3222) <= not a;
    layer2_outputs(3223) <= not b or a;
    layer2_outputs(3224) <= a xor b;
    layer2_outputs(3225) <= a and b;
    layer2_outputs(3226) <= not a;
    layer2_outputs(3227) <= a;
    layer2_outputs(3228) <= a and b;
    layer2_outputs(3229) <= not a;
    layer2_outputs(3230) <= not b;
    layer2_outputs(3231) <= a;
    layer2_outputs(3232) <= b and not a;
    layer2_outputs(3233) <= a;
    layer2_outputs(3234) <= a and not b;
    layer2_outputs(3235) <= not a or b;
    layer2_outputs(3236) <= b;
    layer2_outputs(3237) <= b;
    layer2_outputs(3238) <= b and not a;
    layer2_outputs(3239) <= not b;
    layer2_outputs(3240) <= a xor b;
    layer2_outputs(3241) <= not b or a;
    layer2_outputs(3242) <= a or b;
    layer2_outputs(3243) <= b;
    layer2_outputs(3244) <= not (a and b);
    layer2_outputs(3245) <= a;
    layer2_outputs(3246) <= not b or a;
    layer2_outputs(3247) <= not b;
    layer2_outputs(3248) <= not b or a;
    layer2_outputs(3249) <= a xor b;
    layer2_outputs(3250) <= not (a or b);
    layer2_outputs(3251) <= not (a and b);
    layer2_outputs(3252) <= not b;
    layer2_outputs(3253) <= a and not b;
    layer2_outputs(3254) <= a and b;
    layer2_outputs(3255) <= not a or b;
    layer2_outputs(3256) <= b and not a;
    layer2_outputs(3257) <= a and b;
    layer2_outputs(3258) <= a;
    layer2_outputs(3259) <= a xor b;
    layer2_outputs(3260) <= not (a and b);
    layer2_outputs(3261) <= b;
    layer2_outputs(3262) <= not b or a;
    layer2_outputs(3263) <= not b;
    layer2_outputs(3264) <= not a;
    layer2_outputs(3265) <= not b;
    layer2_outputs(3266) <= not (a or b);
    layer2_outputs(3267) <= not b;
    layer2_outputs(3268) <= a xor b;
    layer2_outputs(3269) <= not b;
    layer2_outputs(3270) <= a;
    layer2_outputs(3271) <= not a;
    layer2_outputs(3272) <= b;
    layer2_outputs(3273) <= a or b;
    layer2_outputs(3274) <= not (a and b);
    layer2_outputs(3275) <= a and not b;
    layer2_outputs(3276) <= b;
    layer2_outputs(3277) <= not (a or b);
    layer2_outputs(3278) <= a and b;
    layer2_outputs(3279) <= a xor b;
    layer2_outputs(3280) <= not (a xor b);
    layer2_outputs(3281) <= not a;
    layer2_outputs(3282) <= a xor b;
    layer2_outputs(3283) <= a or b;
    layer2_outputs(3284) <= a and b;
    layer2_outputs(3285) <= b;
    layer2_outputs(3286) <= not a;
    layer2_outputs(3287) <= not b;
    layer2_outputs(3288) <= not (a or b);
    layer2_outputs(3289) <= not b or a;
    layer2_outputs(3290) <= a xor b;
    layer2_outputs(3291) <= a;
    layer2_outputs(3292) <= not a;
    layer2_outputs(3293) <= not (a or b);
    layer2_outputs(3294) <= not a;
    layer2_outputs(3295) <= b;
    layer2_outputs(3296) <= a or b;
    layer2_outputs(3297) <= not a or b;
    layer2_outputs(3298) <= a xor b;
    layer2_outputs(3299) <= a or b;
    layer2_outputs(3300) <= a xor b;
    layer2_outputs(3301) <= not (a and b);
    layer2_outputs(3302) <= not (a xor b);
    layer2_outputs(3303) <= not a;
    layer2_outputs(3304) <= not a;
    layer2_outputs(3305) <= a and b;
    layer2_outputs(3306) <= b and not a;
    layer2_outputs(3307) <= a and b;
    layer2_outputs(3308) <= not b;
    layer2_outputs(3309) <= not a;
    layer2_outputs(3310) <= a and not b;
    layer2_outputs(3311) <= a and b;
    layer2_outputs(3312) <= not (a and b);
    layer2_outputs(3313) <= b;
    layer2_outputs(3314) <= a;
    layer2_outputs(3315) <= not a;
    layer2_outputs(3316) <= a and b;
    layer2_outputs(3317) <= not (a and b);
    layer2_outputs(3318) <= b;
    layer2_outputs(3319) <= not b;
    layer2_outputs(3320) <= a xor b;
    layer2_outputs(3321) <= not b or a;
    layer2_outputs(3322) <= a and b;
    layer2_outputs(3323) <= not a or b;
    layer2_outputs(3324) <= a xor b;
    layer2_outputs(3325) <= a;
    layer2_outputs(3326) <= a xor b;
    layer2_outputs(3327) <= a or b;
    layer2_outputs(3328) <= a and not b;
    layer2_outputs(3329) <= not b;
    layer2_outputs(3330) <= b and not a;
    layer2_outputs(3331) <= b and not a;
    layer2_outputs(3332) <= not a or b;
    layer2_outputs(3333) <= a xor b;
    layer2_outputs(3334) <= b;
    layer2_outputs(3335) <= a;
    layer2_outputs(3336) <= not a or b;
    layer2_outputs(3337) <= not (a or b);
    layer2_outputs(3338) <= a or b;
    layer2_outputs(3339) <= a and b;
    layer2_outputs(3340) <= a or b;
    layer2_outputs(3341) <= not a or b;
    layer2_outputs(3342) <= a xor b;
    layer2_outputs(3343) <= a or b;
    layer2_outputs(3344) <= not a or b;
    layer2_outputs(3345) <= b and not a;
    layer2_outputs(3346) <= b;
    layer2_outputs(3347) <= not b or a;
    layer2_outputs(3348) <= b and not a;
    layer2_outputs(3349) <= a and b;
    layer2_outputs(3350) <= not (a xor b);
    layer2_outputs(3351) <= not a;
    layer2_outputs(3352) <= not b;
    layer2_outputs(3353) <= 1'b0;
    layer2_outputs(3354) <= b;
    layer2_outputs(3355) <= not (a or b);
    layer2_outputs(3356) <= not (a or b);
    layer2_outputs(3357) <= a and b;
    layer2_outputs(3358) <= a;
    layer2_outputs(3359) <= b and not a;
    layer2_outputs(3360) <= 1'b0;
    layer2_outputs(3361) <= b and not a;
    layer2_outputs(3362) <= not b;
    layer2_outputs(3363) <= not (a or b);
    layer2_outputs(3364) <= b;
    layer2_outputs(3365) <= b and not a;
    layer2_outputs(3366) <= b;
    layer2_outputs(3367) <= 1'b1;
    layer2_outputs(3368) <= not (a and b);
    layer2_outputs(3369) <= a xor b;
    layer2_outputs(3370) <= a or b;
    layer2_outputs(3371) <= not b;
    layer2_outputs(3372) <= a and not b;
    layer2_outputs(3373) <= not a;
    layer2_outputs(3374) <= not (a and b);
    layer2_outputs(3375) <= a;
    layer2_outputs(3376) <= not (a xor b);
    layer2_outputs(3377) <= a;
    layer2_outputs(3378) <= not a;
    layer2_outputs(3379) <= not (a and b);
    layer2_outputs(3380) <= not (a and b);
    layer2_outputs(3381) <= not a;
    layer2_outputs(3382) <= a xor b;
    layer2_outputs(3383) <= a xor b;
    layer2_outputs(3384) <= b;
    layer2_outputs(3385) <= not a or b;
    layer2_outputs(3386) <= not b or a;
    layer2_outputs(3387) <= a or b;
    layer2_outputs(3388) <= b;
    layer2_outputs(3389) <= not a;
    layer2_outputs(3390) <= a and b;
    layer2_outputs(3391) <= b and not a;
    layer2_outputs(3392) <= a and not b;
    layer2_outputs(3393) <= b and not a;
    layer2_outputs(3394) <= b;
    layer2_outputs(3395) <= not (a and b);
    layer2_outputs(3396) <= a and not b;
    layer2_outputs(3397) <= not a or b;
    layer2_outputs(3398) <= not b;
    layer2_outputs(3399) <= not a;
    layer2_outputs(3400) <= not a;
    layer2_outputs(3401) <= a;
    layer2_outputs(3402) <= a;
    layer2_outputs(3403) <= not b or a;
    layer2_outputs(3404) <= b and not a;
    layer2_outputs(3405) <= a and b;
    layer2_outputs(3406) <= b;
    layer2_outputs(3407) <= not (a xor b);
    layer2_outputs(3408) <= b;
    layer2_outputs(3409) <= not b;
    layer2_outputs(3410) <= not a or b;
    layer2_outputs(3411) <= a xor b;
    layer2_outputs(3412) <= not a;
    layer2_outputs(3413) <= not (a and b);
    layer2_outputs(3414) <= not a;
    layer2_outputs(3415) <= not a or b;
    layer2_outputs(3416) <= a xor b;
    layer2_outputs(3417) <= a or b;
    layer2_outputs(3418) <= b;
    layer2_outputs(3419) <= not a;
    layer2_outputs(3420) <= a;
    layer2_outputs(3421) <= not b;
    layer2_outputs(3422) <= a xor b;
    layer2_outputs(3423) <= a;
    layer2_outputs(3424) <= not a;
    layer2_outputs(3425) <= not (a or b);
    layer2_outputs(3426) <= b and not a;
    layer2_outputs(3427) <= not b or a;
    layer2_outputs(3428) <= b and not a;
    layer2_outputs(3429) <= b;
    layer2_outputs(3430) <= a xor b;
    layer2_outputs(3431) <= a or b;
    layer2_outputs(3432) <= a or b;
    layer2_outputs(3433) <= not b or a;
    layer2_outputs(3434) <= a xor b;
    layer2_outputs(3435) <= b and not a;
    layer2_outputs(3436) <= a xor b;
    layer2_outputs(3437) <= not a or b;
    layer2_outputs(3438) <= not (a and b);
    layer2_outputs(3439) <= a;
    layer2_outputs(3440) <= a and not b;
    layer2_outputs(3441) <= not (a or b);
    layer2_outputs(3442) <= not a;
    layer2_outputs(3443) <= a and b;
    layer2_outputs(3444) <= b and not a;
    layer2_outputs(3445) <= a;
    layer2_outputs(3446) <= 1'b0;
    layer2_outputs(3447) <= not b;
    layer2_outputs(3448) <= not (a or b);
    layer2_outputs(3449) <= b;
    layer2_outputs(3450) <= a xor b;
    layer2_outputs(3451) <= a and not b;
    layer2_outputs(3452) <= not b;
    layer2_outputs(3453) <= a;
    layer2_outputs(3454) <= not a;
    layer2_outputs(3455) <= not b;
    layer2_outputs(3456) <= a xor b;
    layer2_outputs(3457) <= a;
    layer2_outputs(3458) <= a;
    layer2_outputs(3459) <= a and not b;
    layer2_outputs(3460) <= a;
    layer2_outputs(3461) <= b and not a;
    layer2_outputs(3462) <= a and not b;
    layer2_outputs(3463) <= not (a or b);
    layer2_outputs(3464) <= b;
    layer2_outputs(3465) <= not b;
    layer2_outputs(3466) <= not (a or b);
    layer2_outputs(3467) <= a and not b;
    layer2_outputs(3468) <= b and not a;
    layer2_outputs(3469) <= not (a xor b);
    layer2_outputs(3470) <= a or b;
    layer2_outputs(3471) <= a;
    layer2_outputs(3472) <= not (a or b);
    layer2_outputs(3473) <= not b;
    layer2_outputs(3474) <= not b;
    layer2_outputs(3475) <= a xor b;
    layer2_outputs(3476) <= not a;
    layer2_outputs(3477) <= b;
    layer2_outputs(3478) <= a xor b;
    layer2_outputs(3479) <= a;
    layer2_outputs(3480) <= a;
    layer2_outputs(3481) <= not a;
    layer2_outputs(3482) <= a;
    layer2_outputs(3483) <= a xor b;
    layer2_outputs(3484) <= a;
    layer2_outputs(3485) <= a and b;
    layer2_outputs(3486) <= not (a and b);
    layer2_outputs(3487) <= b and not a;
    layer2_outputs(3488) <= not b or a;
    layer2_outputs(3489) <= not (a xor b);
    layer2_outputs(3490) <= not (a or b);
    layer2_outputs(3491) <= a;
    layer2_outputs(3492) <= a or b;
    layer2_outputs(3493) <= not (a or b);
    layer2_outputs(3494) <= b;
    layer2_outputs(3495) <= a;
    layer2_outputs(3496) <= not b;
    layer2_outputs(3497) <= a and b;
    layer2_outputs(3498) <= a;
    layer2_outputs(3499) <= not b;
    layer2_outputs(3500) <= not a;
    layer2_outputs(3501) <= not b;
    layer2_outputs(3502) <= a;
    layer2_outputs(3503) <= not (a xor b);
    layer2_outputs(3504) <= a and not b;
    layer2_outputs(3505) <= a and not b;
    layer2_outputs(3506) <= not b;
    layer2_outputs(3507) <= a or b;
    layer2_outputs(3508) <= not a or b;
    layer2_outputs(3509) <= not b or a;
    layer2_outputs(3510) <= b;
    layer2_outputs(3511) <= a;
    layer2_outputs(3512) <= not a;
    layer2_outputs(3513) <= not a;
    layer2_outputs(3514) <= not (a xor b);
    layer2_outputs(3515) <= a xor b;
    layer2_outputs(3516) <= a or b;
    layer2_outputs(3517) <= not b or a;
    layer2_outputs(3518) <= a and b;
    layer2_outputs(3519) <= not a or b;
    layer2_outputs(3520) <= b;
    layer2_outputs(3521) <= a;
    layer2_outputs(3522) <= b and not a;
    layer2_outputs(3523) <= b and not a;
    layer2_outputs(3524) <= a;
    layer2_outputs(3525) <= a xor b;
    layer2_outputs(3526) <= not a or b;
    layer2_outputs(3527) <= a and not b;
    layer2_outputs(3528) <= b and not a;
    layer2_outputs(3529) <= a;
    layer2_outputs(3530) <= b and not a;
    layer2_outputs(3531) <= not (a or b);
    layer2_outputs(3532) <= not (a xor b);
    layer2_outputs(3533) <= a;
    layer2_outputs(3534) <= a xor b;
    layer2_outputs(3535) <= b;
    layer2_outputs(3536) <= a xor b;
    layer2_outputs(3537) <= a and b;
    layer2_outputs(3538) <= a xor b;
    layer2_outputs(3539) <= not b;
    layer2_outputs(3540) <= a xor b;
    layer2_outputs(3541) <= not b or a;
    layer2_outputs(3542) <= b and not a;
    layer2_outputs(3543) <= a or b;
    layer2_outputs(3544) <= a and not b;
    layer2_outputs(3545) <= b;
    layer2_outputs(3546) <= not (a xor b);
    layer2_outputs(3547) <= b;
    layer2_outputs(3548) <= not b or a;
    layer2_outputs(3549) <= a;
    layer2_outputs(3550) <= a and b;
    layer2_outputs(3551) <= a;
    layer2_outputs(3552) <= not a;
    layer2_outputs(3553) <= b;
    layer2_outputs(3554) <= not a;
    layer2_outputs(3555) <= b;
    layer2_outputs(3556) <= not b;
    layer2_outputs(3557) <= a;
    layer2_outputs(3558) <= a and b;
    layer2_outputs(3559) <= a or b;
    layer2_outputs(3560) <= a and b;
    layer2_outputs(3561) <= not a;
    layer2_outputs(3562) <= b and not a;
    layer2_outputs(3563) <= a;
    layer2_outputs(3564) <= a or b;
    layer2_outputs(3565) <= a or b;
    layer2_outputs(3566) <= not b;
    layer2_outputs(3567) <= 1'b1;
    layer2_outputs(3568) <= b;
    layer2_outputs(3569) <= b;
    layer2_outputs(3570) <= a xor b;
    layer2_outputs(3571) <= a;
    layer2_outputs(3572) <= not (a xor b);
    layer2_outputs(3573) <= b;
    layer2_outputs(3574) <= not a;
    layer2_outputs(3575) <= b;
    layer2_outputs(3576) <= a and b;
    layer2_outputs(3577) <= not (a xor b);
    layer2_outputs(3578) <= b and not a;
    layer2_outputs(3579) <= not (a or b);
    layer2_outputs(3580) <= not b;
    layer2_outputs(3581) <= a xor b;
    layer2_outputs(3582) <= a and b;
    layer2_outputs(3583) <= not b;
    layer2_outputs(3584) <= not (a or b);
    layer2_outputs(3585) <= a and not b;
    layer2_outputs(3586) <= b;
    layer2_outputs(3587) <= a;
    layer2_outputs(3588) <= not b;
    layer2_outputs(3589) <= not a;
    layer2_outputs(3590) <= not (a xor b);
    layer2_outputs(3591) <= a or b;
    layer2_outputs(3592) <= not b;
    layer2_outputs(3593) <= not (a and b);
    layer2_outputs(3594) <= not (a or b);
    layer2_outputs(3595) <= b and not a;
    layer2_outputs(3596) <= a xor b;
    layer2_outputs(3597) <= not b or a;
    layer2_outputs(3598) <= not (a or b);
    layer2_outputs(3599) <= a xor b;
    layer2_outputs(3600) <= not a or b;
    layer2_outputs(3601) <= a and b;
    layer2_outputs(3602) <= a xor b;
    layer2_outputs(3603) <= not a or b;
    layer2_outputs(3604) <= not (a or b);
    layer2_outputs(3605) <= a xor b;
    layer2_outputs(3606) <= not b;
    layer2_outputs(3607) <= a;
    layer2_outputs(3608) <= not (a or b);
    layer2_outputs(3609) <= a;
    layer2_outputs(3610) <= a and b;
    layer2_outputs(3611) <= a;
    layer2_outputs(3612) <= a and b;
    layer2_outputs(3613) <= not (a or b);
    layer2_outputs(3614) <= a;
    layer2_outputs(3615) <= not a or b;
    layer2_outputs(3616) <= not b or a;
    layer2_outputs(3617) <= a xor b;
    layer2_outputs(3618) <= not (a xor b);
    layer2_outputs(3619) <= not a or b;
    layer2_outputs(3620) <= not (a or b);
    layer2_outputs(3621) <= not b;
    layer2_outputs(3622) <= a or b;
    layer2_outputs(3623) <= b and not a;
    layer2_outputs(3624) <= not b;
    layer2_outputs(3625) <= not (a and b);
    layer2_outputs(3626) <= a or b;
    layer2_outputs(3627) <= a xor b;
    layer2_outputs(3628) <= not a;
    layer2_outputs(3629) <= not (a xor b);
    layer2_outputs(3630) <= not b;
    layer2_outputs(3631) <= a or b;
    layer2_outputs(3632) <= a or b;
    layer2_outputs(3633) <= a and not b;
    layer2_outputs(3634) <= a;
    layer2_outputs(3635) <= a and not b;
    layer2_outputs(3636) <= b and not a;
    layer2_outputs(3637) <= not (a xor b);
    layer2_outputs(3638) <= b and not a;
    layer2_outputs(3639) <= b and not a;
    layer2_outputs(3640) <= not (a xor b);
    layer2_outputs(3641) <= b;
    layer2_outputs(3642) <= not a;
    layer2_outputs(3643) <= not b;
    layer2_outputs(3644) <= not a or b;
    layer2_outputs(3645) <= not (a xor b);
    layer2_outputs(3646) <= not a;
    layer2_outputs(3647) <= not a or b;
    layer2_outputs(3648) <= not b;
    layer2_outputs(3649) <= not b;
    layer2_outputs(3650) <= b;
    layer2_outputs(3651) <= b and not a;
    layer2_outputs(3652) <= not a;
    layer2_outputs(3653) <= not a or b;
    layer2_outputs(3654) <= a and b;
    layer2_outputs(3655) <= b and not a;
    layer2_outputs(3656) <= not b or a;
    layer2_outputs(3657) <= a and b;
    layer2_outputs(3658) <= not b;
    layer2_outputs(3659) <= not b or a;
    layer2_outputs(3660) <= a and b;
    layer2_outputs(3661) <= not b;
    layer2_outputs(3662) <= not (a xor b);
    layer2_outputs(3663) <= not (a xor b);
    layer2_outputs(3664) <= not b;
    layer2_outputs(3665) <= not a;
    layer2_outputs(3666) <= not (a or b);
    layer2_outputs(3667) <= a;
    layer2_outputs(3668) <= not (a xor b);
    layer2_outputs(3669) <= a and not b;
    layer2_outputs(3670) <= not a or b;
    layer2_outputs(3671) <= b and not a;
    layer2_outputs(3672) <= not (a or b);
    layer2_outputs(3673) <= not a;
    layer2_outputs(3674) <= a and b;
    layer2_outputs(3675) <= not b or a;
    layer2_outputs(3676) <= b;
    layer2_outputs(3677) <= a or b;
    layer2_outputs(3678) <= a xor b;
    layer2_outputs(3679) <= not (a or b);
    layer2_outputs(3680) <= a and not b;
    layer2_outputs(3681) <= b;
    layer2_outputs(3682) <= not b;
    layer2_outputs(3683) <= not b;
    layer2_outputs(3684) <= a and b;
    layer2_outputs(3685) <= a and not b;
    layer2_outputs(3686) <= a and b;
    layer2_outputs(3687) <= a and not b;
    layer2_outputs(3688) <= not a or b;
    layer2_outputs(3689) <= not (a or b);
    layer2_outputs(3690) <= not b;
    layer2_outputs(3691) <= a xor b;
    layer2_outputs(3692) <= b and not a;
    layer2_outputs(3693) <= not b;
    layer2_outputs(3694) <= a and b;
    layer2_outputs(3695) <= b and not a;
    layer2_outputs(3696) <= a;
    layer2_outputs(3697) <= not (a xor b);
    layer2_outputs(3698) <= a or b;
    layer2_outputs(3699) <= 1'b0;
    layer2_outputs(3700) <= b;
    layer2_outputs(3701) <= not (a xor b);
    layer2_outputs(3702) <= b;
    layer2_outputs(3703) <= a and not b;
    layer2_outputs(3704) <= not (a or b);
    layer2_outputs(3705) <= a xor b;
    layer2_outputs(3706) <= not (a and b);
    layer2_outputs(3707) <= not b;
    layer2_outputs(3708) <= a;
    layer2_outputs(3709) <= a and b;
    layer2_outputs(3710) <= not b or a;
    layer2_outputs(3711) <= b;
    layer2_outputs(3712) <= a;
    layer2_outputs(3713) <= not a;
    layer2_outputs(3714) <= b and not a;
    layer2_outputs(3715) <= not (a xor b);
    layer2_outputs(3716) <= b;
    layer2_outputs(3717) <= not (a or b);
    layer2_outputs(3718) <= not b;
    layer2_outputs(3719) <= a;
    layer2_outputs(3720) <= not b;
    layer2_outputs(3721) <= not b or a;
    layer2_outputs(3722) <= not a;
    layer2_outputs(3723) <= not a or b;
    layer2_outputs(3724) <= a and not b;
    layer2_outputs(3725) <= a xor b;
    layer2_outputs(3726) <= b and not a;
    layer2_outputs(3727) <= not a;
    layer2_outputs(3728) <= not b;
    layer2_outputs(3729) <= not a;
    layer2_outputs(3730) <= not a;
    layer2_outputs(3731) <= a or b;
    layer2_outputs(3732) <= not a;
    layer2_outputs(3733) <= a or b;
    layer2_outputs(3734) <= b;
    layer2_outputs(3735) <= b;
    layer2_outputs(3736) <= a;
    layer2_outputs(3737) <= a or b;
    layer2_outputs(3738) <= a and b;
    layer2_outputs(3739) <= b;
    layer2_outputs(3740) <= not (a xor b);
    layer2_outputs(3741) <= a xor b;
    layer2_outputs(3742) <= not a or b;
    layer2_outputs(3743) <= a;
    layer2_outputs(3744) <= a;
    layer2_outputs(3745) <= not b or a;
    layer2_outputs(3746) <= b and not a;
    layer2_outputs(3747) <= not (a xor b);
    layer2_outputs(3748) <= not (a xor b);
    layer2_outputs(3749) <= not a;
    layer2_outputs(3750) <= not b;
    layer2_outputs(3751) <= not b;
    layer2_outputs(3752) <= not (a and b);
    layer2_outputs(3753) <= not (a or b);
    layer2_outputs(3754) <= a;
    layer2_outputs(3755) <= not b or a;
    layer2_outputs(3756) <= not a or b;
    layer2_outputs(3757) <= not b;
    layer2_outputs(3758) <= a or b;
    layer2_outputs(3759) <= not b or a;
    layer2_outputs(3760) <= a or b;
    layer2_outputs(3761) <= not b or a;
    layer2_outputs(3762) <= a;
    layer2_outputs(3763) <= b;
    layer2_outputs(3764) <= not a or b;
    layer2_outputs(3765) <= a;
    layer2_outputs(3766) <= a and b;
    layer2_outputs(3767) <= not a;
    layer2_outputs(3768) <= not a or b;
    layer2_outputs(3769) <= not (a or b);
    layer2_outputs(3770) <= a;
    layer2_outputs(3771) <= not b or a;
    layer2_outputs(3772) <= b;
    layer2_outputs(3773) <= not (a and b);
    layer2_outputs(3774) <= a xor b;
    layer2_outputs(3775) <= not a or b;
    layer2_outputs(3776) <= a xor b;
    layer2_outputs(3777) <= a and b;
    layer2_outputs(3778) <= a or b;
    layer2_outputs(3779) <= a and b;
    layer2_outputs(3780) <= a;
    layer2_outputs(3781) <= not b or a;
    layer2_outputs(3782) <= not (a and b);
    layer2_outputs(3783) <= a;
    layer2_outputs(3784) <= a and not b;
    layer2_outputs(3785) <= b;
    layer2_outputs(3786) <= b and not a;
    layer2_outputs(3787) <= b;
    layer2_outputs(3788) <= not b;
    layer2_outputs(3789) <= a xor b;
    layer2_outputs(3790) <= not (a and b);
    layer2_outputs(3791) <= a or b;
    layer2_outputs(3792) <= b;
    layer2_outputs(3793) <= b;
    layer2_outputs(3794) <= not (a and b);
    layer2_outputs(3795) <= not (a or b);
    layer2_outputs(3796) <= not a or b;
    layer2_outputs(3797) <= a xor b;
    layer2_outputs(3798) <= a;
    layer2_outputs(3799) <= not (a xor b);
    layer2_outputs(3800) <= not a or b;
    layer2_outputs(3801) <= not b;
    layer2_outputs(3802) <= a;
    layer2_outputs(3803) <= a and b;
    layer2_outputs(3804) <= not b or a;
    layer2_outputs(3805) <= not (a and b);
    layer2_outputs(3806) <= not b or a;
    layer2_outputs(3807) <= a and not b;
    layer2_outputs(3808) <= not a or b;
    layer2_outputs(3809) <= not a;
    layer2_outputs(3810) <= not a or b;
    layer2_outputs(3811) <= not (a xor b);
    layer2_outputs(3812) <= a and not b;
    layer2_outputs(3813) <= a;
    layer2_outputs(3814) <= not (a xor b);
    layer2_outputs(3815) <= not a;
    layer2_outputs(3816) <= not (a or b);
    layer2_outputs(3817) <= not b;
    layer2_outputs(3818) <= a and not b;
    layer2_outputs(3819) <= not a;
    layer2_outputs(3820) <= a;
    layer2_outputs(3821) <= not (a xor b);
    layer2_outputs(3822) <= not a or b;
    layer2_outputs(3823) <= not b;
    layer2_outputs(3824) <= a and b;
    layer2_outputs(3825) <= not a;
    layer2_outputs(3826) <= not b;
    layer2_outputs(3827) <= not (a and b);
    layer2_outputs(3828) <= a or b;
    layer2_outputs(3829) <= not a;
    layer2_outputs(3830) <= a xor b;
    layer2_outputs(3831) <= b;
    layer2_outputs(3832) <= not (a xor b);
    layer2_outputs(3833) <= a and not b;
    layer2_outputs(3834) <= not (a or b);
    layer2_outputs(3835) <= not a or b;
    layer2_outputs(3836) <= not a;
    layer2_outputs(3837) <= not a;
    layer2_outputs(3838) <= not a;
    layer2_outputs(3839) <= a;
    layer2_outputs(3840) <= b;
    layer2_outputs(3841) <= a and b;
    layer2_outputs(3842) <= a;
    layer2_outputs(3843) <= b;
    layer2_outputs(3844) <= not (a and b);
    layer2_outputs(3845) <= not b;
    layer2_outputs(3846) <= not b;
    layer2_outputs(3847) <= a or b;
    layer2_outputs(3848) <= 1'b0;
    layer2_outputs(3849) <= a or b;
    layer2_outputs(3850) <= not (a xor b);
    layer2_outputs(3851) <= a or b;
    layer2_outputs(3852) <= not a or b;
    layer2_outputs(3853) <= not a;
    layer2_outputs(3854) <= a;
    layer2_outputs(3855) <= a;
    layer2_outputs(3856) <= not b;
    layer2_outputs(3857) <= not b;
    layer2_outputs(3858) <= b and not a;
    layer2_outputs(3859) <= not (a and b);
    layer2_outputs(3860) <= a;
    layer2_outputs(3861) <= a and not b;
    layer2_outputs(3862) <= a or b;
    layer2_outputs(3863) <= not b;
    layer2_outputs(3864) <= not b;
    layer2_outputs(3865) <= not b or a;
    layer2_outputs(3866) <= not a;
    layer2_outputs(3867) <= not b;
    layer2_outputs(3868) <= not b or a;
    layer2_outputs(3869) <= not (a xor b);
    layer2_outputs(3870) <= not (a xor b);
    layer2_outputs(3871) <= b;
    layer2_outputs(3872) <= not (a and b);
    layer2_outputs(3873) <= a and b;
    layer2_outputs(3874) <= a or b;
    layer2_outputs(3875) <= not b;
    layer2_outputs(3876) <= not b or a;
    layer2_outputs(3877) <= not b;
    layer2_outputs(3878) <= b;
    layer2_outputs(3879) <= not b;
    layer2_outputs(3880) <= b and not a;
    layer2_outputs(3881) <= b and not a;
    layer2_outputs(3882) <= a or b;
    layer2_outputs(3883) <= a;
    layer2_outputs(3884) <= not a;
    layer2_outputs(3885) <= a xor b;
    layer2_outputs(3886) <= a and b;
    layer2_outputs(3887) <= not (a xor b);
    layer2_outputs(3888) <= not a;
    layer2_outputs(3889) <= not a;
    layer2_outputs(3890) <= not (a or b);
    layer2_outputs(3891) <= a xor b;
    layer2_outputs(3892) <= not a or b;
    layer2_outputs(3893) <= a and not b;
    layer2_outputs(3894) <= a xor b;
    layer2_outputs(3895) <= not b;
    layer2_outputs(3896) <= b and not a;
    layer2_outputs(3897) <= not a;
    layer2_outputs(3898) <= b and not a;
    layer2_outputs(3899) <= b and not a;
    layer2_outputs(3900) <= not (a or b);
    layer2_outputs(3901) <= b and not a;
    layer2_outputs(3902) <= not (a or b);
    layer2_outputs(3903) <= not b or a;
    layer2_outputs(3904) <= b and not a;
    layer2_outputs(3905) <= a;
    layer2_outputs(3906) <= 1'b0;
    layer2_outputs(3907) <= a and not b;
    layer2_outputs(3908) <= not (a and b);
    layer2_outputs(3909) <= a xor b;
    layer2_outputs(3910) <= a xor b;
    layer2_outputs(3911) <= b;
    layer2_outputs(3912) <= b;
    layer2_outputs(3913) <= not a or b;
    layer2_outputs(3914) <= not b;
    layer2_outputs(3915) <= 1'b0;
    layer2_outputs(3916) <= not (a xor b);
    layer2_outputs(3917) <= not b;
    layer2_outputs(3918) <= not b;
    layer2_outputs(3919) <= a or b;
    layer2_outputs(3920) <= not (a and b);
    layer2_outputs(3921) <= not a or b;
    layer2_outputs(3922) <= not a;
    layer2_outputs(3923) <= not b or a;
    layer2_outputs(3924) <= a xor b;
    layer2_outputs(3925) <= not (a or b);
    layer2_outputs(3926) <= b;
    layer2_outputs(3927) <= not (a or b);
    layer2_outputs(3928) <= not a;
    layer2_outputs(3929) <= not (a xor b);
    layer2_outputs(3930) <= not (a and b);
    layer2_outputs(3931) <= a and b;
    layer2_outputs(3932) <= not (a and b);
    layer2_outputs(3933) <= a xor b;
    layer2_outputs(3934) <= a;
    layer2_outputs(3935) <= not b or a;
    layer2_outputs(3936) <= not a;
    layer2_outputs(3937) <= a;
    layer2_outputs(3938) <= not b;
    layer2_outputs(3939) <= not b;
    layer2_outputs(3940) <= not b or a;
    layer2_outputs(3941) <= not a;
    layer2_outputs(3942) <= a xor b;
    layer2_outputs(3943) <= a or b;
    layer2_outputs(3944) <= a;
    layer2_outputs(3945) <= not (a or b);
    layer2_outputs(3946) <= not b or a;
    layer2_outputs(3947) <= not b or a;
    layer2_outputs(3948) <= not a or b;
    layer2_outputs(3949) <= b;
    layer2_outputs(3950) <= a xor b;
    layer2_outputs(3951) <= a or b;
    layer2_outputs(3952) <= not (a xor b);
    layer2_outputs(3953) <= not b;
    layer2_outputs(3954) <= b and not a;
    layer2_outputs(3955) <= not a;
    layer2_outputs(3956) <= a or b;
    layer2_outputs(3957) <= a and not b;
    layer2_outputs(3958) <= not (a or b);
    layer2_outputs(3959) <= a xor b;
    layer2_outputs(3960) <= not a or b;
    layer2_outputs(3961) <= not a or b;
    layer2_outputs(3962) <= not b;
    layer2_outputs(3963) <= a;
    layer2_outputs(3964) <= not (a xor b);
    layer2_outputs(3965) <= not (a xor b);
    layer2_outputs(3966) <= a and b;
    layer2_outputs(3967) <= not a;
    layer2_outputs(3968) <= a or b;
    layer2_outputs(3969) <= a or b;
    layer2_outputs(3970) <= not a or b;
    layer2_outputs(3971) <= not b or a;
    layer2_outputs(3972) <= a;
    layer2_outputs(3973) <= a xor b;
    layer2_outputs(3974) <= not a or b;
    layer2_outputs(3975) <= not b;
    layer2_outputs(3976) <= a and b;
    layer2_outputs(3977) <= not a or b;
    layer2_outputs(3978) <= a;
    layer2_outputs(3979) <= b;
    layer2_outputs(3980) <= not (a or b);
    layer2_outputs(3981) <= not (a xor b);
    layer2_outputs(3982) <= not b;
    layer2_outputs(3983) <= not b;
    layer2_outputs(3984) <= a xor b;
    layer2_outputs(3985) <= b and not a;
    layer2_outputs(3986) <= not (a xor b);
    layer2_outputs(3987) <= a;
    layer2_outputs(3988) <= not b;
    layer2_outputs(3989) <= not b;
    layer2_outputs(3990) <= not a;
    layer2_outputs(3991) <= not a;
    layer2_outputs(3992) <= not a;
    layer2_outputs(3993) <= not a;
    layer2_outputs(3994) <= not b;
    layer2_outputs(3995) <= a and b;
    layer2_outputs(3996) <= a xor b;
    layer2_outputs(3997) <= not (a and b);
    layer2_outputs(3998) <= not a;
    layer2_outputs(3999) <= a xor b;
    layer2_outputs(4000) <= not a;
    layer2_outputs(4001) <= a xor b;
    layer2_outputs(4002) <= not (a xor b);
    layer2_outputs(4003) <= a xor b;
    layer2_outputs(4004) <= b and not a;
    layer2_outputs(4005) <= 1'b1;
    layer2_outputs(4006) <= a and b;
    layer2_outputs(4007) <= a;
    layer2_outputs(4008) <= a and b;
    layer2_outputs(4009) <= not a;
    layer2_outputs(4010) <= not (a xor b);
    layer2_outputs(4011) <= b;
    layer2_outputs(4012) <= not b or a;
    layer2_outputs(4013) <= not (a or b);
    layer2_outputs(4014) <= a and not b;
    layer2_outputs(4015) <= b;
    layer2_outputs(4016) <= not b;
    layer2_outputs(4017) <= b and not a;
    layer2_outputs(4018) <= a or b;
    layer2_outputs(4019) <= b and not a;
    layer2_outputs(4020) <= a;
    layer2_outputs(4021) <= not (a and b);
    layer2_outputs(4022) <= b;
    layer2_outputs(4023) <= not b;
    layer2_outputs(4024) <= not a;
    layer2_outputs(4025) <= a or b;
    layer2_outputs(4026) <= a and b;
    layer2_outputs(4027) <= not (a xor b);
    layer2_outputs(4028) <= a or b;
    layer2_outputs(4029) <= a or b;
    layer2_outputs(4030) <= not a or b;
    layer2_outputs(4031) <= a and b;
    layer2_outputs(4032) <= a;
    layer2_outputs(4033) <= b and not a;
    layer2_outputs(4034) <= b;
    layer2_outputs(4035) <= a or b;
    layer2_outputs(4036) <= not (a xor b);
    layer2_outputs(4037) <= a or b;
    layer2_outputs(4038) <= not (a and b);
    layer2_outputs(4039) <= not a;
    layer2_outputs(4040) <= b and not a;
    layer2_outputs(4041) <= a and not b;
    layer2_outputs(4042) <= not (a or b);
    layer2_outputs(4043) <= not b;
    layer2_outputs(4044) <= not (a and b);
    layer2_outputs(4045) <= not b;
    layer2_outputs(4046) <= a and b;
    layer2_outputs(4047) <= a xor b;
    layer2_outputs(4048) <= a;
    layer2_outputs(4049) <= a xor b;
    layer2_outputs(4050) <= a;
    layer2_outputs(4051) <= a and b;
    layer2_outputs(4052) <= not a;
    layer2_outputs(4053) <= not b or a;
    layer2_outputs(4054) <= a xor b;
    layer2_outputs(4055) <= a xor b;
    layer2_outputs(4056) <= b;
    layer2_outputs(4057) <= b;
    layer2_outputs(4058) <= a and b;
    layer2_outputs(4059) <= not (a and b);
    layer2_outputs(4060) <= not (a or b);
    layer2_outputs(4061) <= not a or b;
    layer2_outputs(4062) <= not (a xor b);
    layer2_outputs(4063) <= not (a xor b);
    layer2_outputs(4064) <= b;
    layer2_outputs(4065) <= a;
    layer2_outputs(4066) <= not (a or b);
    layer2_outputs(4067) <= a or b;
    layer2_outputs(4068) <= not (a and b);
    layer2_outputs(4069) <= a xor b;
    layer2_outputs(4070) <= b and not a;
    layer2_outputs(4071) <= not b or a;
    layer2_outputs(4072) <= a;
    layer2_outputs(4073) <= not b;
    layer2_outputs(4074) <= not b or a;
    layer2_outputs(4075) <= not (a xor b);
    layer2_outputs(4076) <= not b;
    layer2_outputs(4077) <= a;
    layer2_outputs(4078) <= not b or a;
    layer2_outputs(4079) <= a or b;
    layer2_outputs(4080) <= not a or b;
    layer2_outputs(4081) <= a;
    layer2_outputs(4082) <= not (a and b);
    layer2_outputs(4083) <= b;
    layer2_outputs(4084) <= not b;
    layer2_outputs(4085) <= not a or b;
    layer2_outputs(4086) <= b and not a;
    layer2_outputs(4087) <= not b;
    layer2_outputs(4088) <= not (a or b);
    layer2_outputs(4089) <= not b or a;
    layer2_outputs(4090) <= a;
    layer2_outputs(4091) <= b and not a;
    layer2_outputs(4092) <= not (a or b);
    layer2_outputs(4093) <= not b;
    layer2_outputs(4094) <= not (a and b);
    layer2_outputs(4095) <= b;
    layer2_outputs(4096) <= a;
    layer2_outputs(4097) <= a;
    layer2_outputs(4098) <= b and not a;
    layer2_outputs(4099) <= not a or b;
    layer2_outputs(4100) <= a and b;
    layer2_outputs(4101) <= a and b;
    layer2_outputs(4102) <= a and not b;
    layer2_outputs(4103) <= a;
    layer2_outputs(4104) <= b and not a;
    layer2_outputs(4105) <= b and not a;
    layer2_outputs(4106) <= not a or b;
    layer2_outputs(4107) <= not a;
    layer2_outputs(4108) <= not b;
    layer2_outputs(4109) <= b and not a;
    layer2_outputs(4110) <= not (a and b);
    layer2_outputs(4111) <= not a or b;
    layer2_outputs(4112) <= not b;
    layer2_outputs(4113) <= not (a xor b);
    layer2_outputs(4114) <= not a or b;
    layer2_outputs(4115) <= not b or a;
    layer2_outputs(4116) <= a xor b;
    layer2_outputs(4117) <= a and not b;
    layer2_outputs(4118) <= b and not a;
    layer2_outputs(4119) <= not b;
    layer2_outputs(4120) <= a;
    layer2_outputs(4121) <= not b;
    layer2_outputs(4122) <= a;
    layer2_outputs(4123) <= not a;
    layer2_outputs(4124) <= a;
    layer2_outputs(4125) <= not (a xor b);
    layer2_outputs(4126) <= a or b;
    layer2_outputs(4127) <= not (a and b);
    layer2_outputs(4128) <= a;
    layer2_outputs(4129) <= not b or a;
    layer2_outputs(4130) <= a or b;
    layer2_outputs(4131) <= not (a and b);
    layer2_outputs(4132) <= not (a xor b);
    layer2_outputs(4133) <= not (a or b);
    layer2_outputs(4134) <= not (a or b);
    layer2_outputs(4135) <= b;
    layer2_outputs(4136) <= not a;
    layer2_outputs(4137) <= a xor b;
    layer2_outputs(4138) <= a;
    layer2_outputs(4139) <= a and b;
    layer2_outputs(4140) <= not (a and b);
    layer2_outputs(4141) <= a xor b;
    layer2_outputs(4142) <= a;
    layer2_outputs(4143) <= a;
    layer2_outputs(4144) <= not a;
    layer2_outputs(4145) <= not b;
    layer2_outputs(4146) <= a or b;
    layer2_outputs(4147) <= b;
    layer2_outputs(4148) <= a xor b;
    layer2_outputs(4149) <= not a;
    layer2_outputs(4150) <= a and b;
    layer2_outputs(4151) <= a;
    layer2_outputs(4152) <= b;
    layer2_outputs(4153) <= not a;
    layer2_outputs(4154) <= not (a or b);
    layer2_outputs(4155) <= not b;
    layer2_outputs(4156) <= a and not b;
    layer2_outputs(4157) <= a and b;
    layer2_outputs(4158) <= a;
    layer2_outputs(4159) <= not a;
    layer2_outputs(4160) <= not (a and b);
    layer2_outputs(4161) <= not a;
    layer2_outputs(4162) <= not b;
    layer2_outputs(4163) <= b;
    layer2_outputs(4164) <= a and b;
    layer2_outputs(4165) <= a xor b;
    layer2_outputs(4166) <= not b or a;
    layer2_outputs(4167) <= b;
    layer2_outputs(4168) <= not (a xor b);
    layer2_outputs(4169) <= b and not a;
    layer2_outputs(4170) <= not a;
    layer2_outputs(4171) <= not b;
    layer2_outputs(4172) <= b;
    layer2_outputs(4173) <= not a or b;
    layer2_outputs(4174) <= not a;
    layer2_outputs(4175) <= not b or a;
    layer2_outputs(4176) <= b;
    layer2_outputs(4177) <= not (a xor b);
    layer2_outputs(4178) <= not a;
    layer2_outputs(4179) <= not b;
    layer2_outputs(4180) <= not b;
    layer2_outputs(4181) <= not (a and b);
    layer2_outputs(4182) <= not b;
    layer2_outputs(4183) <= a;
    layer2_outputs(4184) <= a or b;
    layer2_outputs(4185) <= not (a xor b);
    layer2_outputs(4186) <= not a;
    layer2_outputs(4187) <= not b;
    layer2_outputs(4188) <= not a or b;
    layer2_outputs(4189) <= a;
    layer2_outputs(4190) <= not (a and b);
    layer2_outputs(4191) <= not b;
    layer2_outputs(4192) <= not (a or b);
    layer2_outputs(4193) <= not (a or b);
    layer2_outputs(4194) <= b;
    layer2_outputs(4195) <= not a;
    layer2_outputs(4196) <= a and not b;
    layer2_outputs(4197) <= a and not b;
    layer2_outputs(4198) <= b;
    layer2_outputs(4199) <= not b;
    layer2_outputs(4200) <= not a or b;
    layer2_outputs(4201) <= not (a xor b);
    layer2_outputs(4202) <= not (a xor b);
    layer2_outputs(4203) <= not a or b;
    layer2_outputs(4204) <= b;
    layer2_outputs(4205) <= b;
    layer2_outputs(4206) <= not (a xor b);
    layer2_outputs(4207) <= a or b;
    layer2_outputs(4208) <= not a;
    layer2_outputs(4209) <= a;
    layer2_outputs(4210) <= not (a xor b);
    layer2_outputs(4211) <= b;
    layer2_outputs(4212) <= not (a xor b);
    layer2_outputs(4213) <= a;
    layer2_outputs(4214) <= not b or a;
    layer2_outputs(4215) <= a xor b;
    layer2_outputs(4216) <= not a or b;
    layer2_outputs(4217) <= not a;
    layer2_outputs(4218) <= b;
    layer2_outputs(4219) <= a xor b;
    layer2_outputs(4220) <= not a or b;
    layer2_outputs(4221) <= not a;
    layer2_outputs(4222) <= a and not b;
    layer2_outputs(4223) <= a and b;
    layer2_outputs(4224) <= a and b;
    layer2_outputs(4225) <= not a or b;
    layer2_outputs(4226) <= not a or b;
    layer2_outputs(4227) <= not a;
    layer2_outputs(4228) <= not a;
    layer2_outputs(4229) <= a xor b;
    layer2_outputs(4230) <= a;
    layer2_outputs(4231) <= not (a or b);
    layer2_outputs(4232) <= not b;
    layer2_outputs(4233) <= a or b;
    layer2_outputs(4234) <= b;
    layer2_outputs(4235) <= not a;
    layer2_outputs(4236) <= not b or a;
    layer2_outputs(4237) <= a and not b;
    layer2_outputs(4238) <= a and b;
    layer2_outputs(4239) <= not b or a;
    layer2_outputs(4240) <= not (a or b);
    layer2_outputs(4241) <= a;
    layer2_outputs(4242) <= b;
    layer2_outputs(4243) <= a;
    layer2_outputs(4244) <= not a;
    layer2_outputs(4245) <= a and b;
    layer2_outputs(4246) <= not a or b;
    layer2_outputs(4247) <= a;
    layer2_outputs(4248) <= a or b;
    layer2_outputs(4249) <= not (a xor b);
    layer2_outputs(4250) <= a xor b;
    layer2_outputs(4251) <= not (a and b);
    layer2_outputs(4252) <= not (a and b);
    layer2_outputs(4253) <= not b;
    layer2_outputs(4254) <= not (a and b);
    layer2_outputs(4255) <= not b;
    layer2_outputs(4256) <= b and not a;
    layer2_outputs(4257) <= not a or b;
    layer2_outputs(4258) <= a and not b;
    layer2_outputs(4259) <= b and not a;
    layer2_outputs(4260) <= a or b;
    layer2_outputs(4261) <= a and not b;
    layer2_outputs(4262) <= a;
    layer2_outputs(4263) <= not a;
    layer2_outputs(4264) <= a;
    layer2_outputs(4265) <= a;
    layer2_outputs(4266) <= b;
    layer2_outputs(4267) <= a or b;
    layer2_outputs(4268) <= a and not b;
    layer2_outputs(4269) <= not b or a;
    layer2_outputs(4270) <= a or b;
    layer2_outputs(4271) <= a;
    layer2_outputs(4272) <= b and not a;
    layer2_outputs(4273) <= not b;
    layer2_outputs(4274) <= b and not a;
    layer2_outputs(4275) <= not a;
    layer2_outputs(4276) <= b and not a;
    layer2_outputs(4277) <= not b or a;
    layer2_outputs(4278) <= b and not a;
    layer2_outputs(4279) <= not b or a;
    layer2_outputs(4280) <= not b or a;
    layer2_outputs(4281) <= b and not a;
    layer2_outputs(4282) <= not b;
    layer2_outputs(4283) <= not a or b;
    layer2_outputs(4284) <= not a;
    layer2_outputs(4285) <= not b;
    layer2_outputs(4286) <= a and not b;
    layer2_outputs(4287) <= not (a xor b);
    layer2_outputs(4288) <= not a;
    layer2_outputs(4289) <= not (a or b);
    layer2_outputs(4290) <= not a or b;
    layer2_outputs(4291) <= a;
    layer2_outputs(4292) <= not b;
    layer2_outputs(4293) <= not b;
    layer2_outputs(4294) <= not a or b;
    layer2_outputs(4295) <= b;
    layer2_outputs(4296) <= not a;
    layer2_outputs(4297) <= not a;
    layer2_outputs(4298) <= b and not a;
    layer2_outputs(4299) <= b and not a;
    layer2_outputs(4300) <= a and not b;
    layer2_outputs(4301) <= a and b;
    layer2_outputs(4302) <= b;
    layer2_outputs(4303) <= a and not b;
    layer2_outputs(4304) <= a xor b;
    layer2_outputs(4305) <= a xor b;
    layer2_outputs(4306) <= b;
    layer2_outputs(4307) <= not b;
    layer2_outputs(4308) <= not b;
    layer2_outputs(4309) <= b;
    layer2_outputs(4310) <= a and not b;
    layer2_outputs(4311) <= a;
    layer2_outputs(4312) <= b;
    layer2_outputs(4313) <= not (a and b);
    layer2_outputs(4314) <= b;
    layer2_outputs(4315) <= a;
    layer2_outputs(4316) <= not b;
    layer2_outputs(4317) <= b and not a;
    layer2_outputs(4318) <= b;
    layer2_outputs(4319) <= not b or a;
    layer2_outputs(4320) <= not a;
    layer2_outputs(4321) <= not (a or b);
    layer2_outputs(4322) <= not a;
    layer2_outputs(4323) <= a xor b;
    layer2_outputs(4324) <= not a;
    layer2_outputs(4325) <= a xor b;
    layer2_outputs(4326) <= not a;
    layer2_outputs(4327) <= b;
    layer2_outputs(4328) <= not b;
    layer2_outputs(4329) <= b and not a;
    layer2_outputs(4330) <= a;
    layer2_outputs(4331) <= a or b;
    layer2_outputs(4332) <= not b;
    layer2_outputs(4333) <= not (a or b);
    layer2_outputs(4334) <= a;
    layer2_outputs(4335) <= a xor b;
    layer2_outputs(4336) <= not (a and b);
    layer2_outputs(4337) <= b;
    layer2_outputs(4338) <= b;
    layer2_outputs(4339) <= a and not b;
    layer2_outputs(4340) <= not (a xor b);
    layer2_outputs(4341) <= b;
    layer2_outputs(4342) <= not b or a;
    layer2_outputs(4343) <= not (a and b);
    layer2_outputs(4344) <= b;
    layer2_outputs(4345) <= a;
    layer2_outputs(4346) <= not a or b;
    layer2_outputs(4347) <= b;
    layer2_outputs(4348) <= a and not b;
    layer2_outputs(4349) <= not b;
    layer2_outputs(4350) <= not a;
    layer2_outputs(4351) <= not a or b;
    layer2_outputs(4352) <= b;
    layer2_outputs(4353) <= not b;
    layer2_outputs(4354) <= a and not b;
    layer2_outputs(4355) <= b;
    layer2_outputs(4356) <= a xor b;
    layer2_outputs(4357) <= b;
    layer2_outputs(4358) <= b;
    layer2_outputs(4359) <= a or b;
    layer2_outputs(4360) <= not b;
    layer2_outputs(4361) <= a;
    layer2_outputs(4362) <= not b;
    layer2_outputs(4363) <= b and not a;
    layer2_outputs(4364) <= not a;
    layer2_outputs(4365) <= not b or a;
    layer2_outputs(4366) <= a;
    layer2_outputs(4367) <= b;
    layer2_outputs(4368) <= b;
    layer2_outputs(4369) <= not a or b;
    layer2_outputs(4370) <= a and not b;
    layer2_outputs(4371) <= b;
    layer2_outputs(4372) <= a and not b;
    layer2_outputs(4373) <= not a or b;
    layer2_outputs(4374) <= not (a and b);
    layer2_outputs(4375) <= not b or a;
    layer2_outputs(4376) <= not a;
    layer2_outputs(4377) <= b and not a;
    layer2_outputs(4378) <= a and not b;
    layer2_outputs(4379) <= a xor b;
    layer2_outputs(4380) <= a and b;
    layer2_outputs(4381) <= not b;
    layer2_outputs(4382) <= not (a and b);
    layer2_outputs(4383) <= not (a xor b);
    layer2_outputs(4384) <= b;
    layer2_outputs(4385) <= not a or b;
    layer2_outputs(4386) <= not (a or b);
    layer2_outputs(4387) <= a and not b;
    layer2_outputs(4388) <= not b or a;
    layer2_outputs(4389) <= not b or a;
    layer2_outputs(4390) <= a;
    layer2_outputs(4391) <= a;
    layer2_outputs(4392) <= a;
    layer2_outputs(4393) <= not (a xor b);
    layer2_outputs(4394) <= not b or a;
    layer2_outputs(4395) <= not a;
    layer2_outputs(4396) <= not a or b;
    layer2_outputs(4397) <= a xor b;
    layer2_outputs(4398) <= b;
    layer2_outputs(4399) <= a and not b;
    layer2_outputs(4400) <= a and b;
    layer2_outputs(4401) <= not a;
    layer2_outputs(4402) <= a;
    layer2_outputs(4403) <= a and not b;
    layer2_outputs(4404) <= a;
    layer2_outputs(4405) <= not b;
    layer2_outputs(4406) <= a;
    layer2_outputs(4407) <= b;
    layer2_outputs(4408) <= b and not a;
    layer2_outputs(4409) <= not (a or b);
    layer2_outputs(4410) <= not b;
    layer2_outputs(4411) <= a;
    layer2_outputs(4412) <= b;
    layer2_outputs(4413) <= b and not a;
    layer2_outputs(4414) <= not b;
    layer2_outputs(4415) <= a and b;
    layer2_outputs(4416) <= not b;
    layer2_outputs(4417) <= b and not a;
    layer2_outputs(4418) <= b;
    layer2_outputs(4419) <= b;
    layer2_outputs(4420) <= not a;
    layer2_outputs(4421) <= b;
    layer2_outputs(4422) <= b and not a;
    layer2_outputs(4423) <= b;
    layer2_outputs(4424) <= not b or a;
    layer2_outputs(4425) <= b;
    layer2_outputs(4426) <= not a;
    layer2_outputs(4427) <= not (a xor b);
    layer2_outputs(4428) <= not a or b;
    layer2_outputs(4429) <= a xor b;
    layer2_outputs(4430) <= a and b;
    layer2_outputs(4431) <= not a or b;
    layer2_outputs(4432) <= 1'b1;
    layer2_outputs(4433) <= a;
    layer2_outputs(4434) <= not b or a;
    layer2_outputs(4435) <= not (a and b);
    layer2_outputs(4436) <= not (a or b);
    layer2_outputs(4437) <= 1'b0;
    layer2_outputs(4438) <= not b or a;
    layer2_outputs(4439) <= not b;
    layer2_outputs(4440) <= b and not a;
    layer2_outputs(4441) <= not (a xor b);
    layer2_outputs(4442) <= not b or a;
    layer2_outputs(4443) <= not a or b;
    layer2_outputs(4444) <= a;
    layer2_outputs(4445) <= a;
    layer2_outputs(4446) <= not b;
    layer2_outputs(4447) <= a;
    layer2_outputs(4448) <= a xor b;
    layer2_outputs(4449) <= a and b;
    layer2_outputs(4450) <= not b;
    layer2_outputs(4451) <= b;
    layer2_outputs(4452) <= a xor b;
    layer2_outputs(4453) <= a and b;
    layer2_outputs(4454) <= not (a and b);
    layer2_outputs(4455) <= not (a or b);
    layer2_outputs(4456) <= b;
    layer2_outputs(4457) <= not (a and b);
    layer2_outputs(4458) <= b;
    layer2_outputs(4459) <= a xor b;
    layer2_outputs(4460) <= not a;
    layer2_outputs(4461) <= not (a xor b);
    layer2_outputs(4462) <= not a;
    layer2_outputs(4463) <= a and b;
    layer2_outputs(4464) <= a and not b;
    layer2_outputs(4465) <= not b or a;
    layer2_outputs(4466) <= a and b;
    layer2_outputs(4467) <= not b or a;
    layer2_outputs(4468) <= a;
    layer2_outputs(4469) <= a xor b;
    layer2_outputs(4470) <= not (a or b);
    layer2_outputs(4471) <= a and not b;
    layer2_outputs(4472) <= not b;
    layer2_outputs(4473) <= a;
    layer2_outputs(4474) <= not (a xor b);
    layer2_outputs(4475) <= a or b;
    layer2_outputs(4476) <= a;
    layer2_outputs(4477) <= a xor b;
    layer2_outputs(4478) <= a or b;
    layer2_outputs(4479) <= not a;
    layer2_outputs(4480) <= a xor b;
    layer2_outputs(4481) <= not a;
    layer2_outputs(4482) <= not (a xor b);
    layer2_outputs(4483) <= not (a xor b);
    layer2_outputs(4484) <= not (a or b);
    layer2_outputs(4485) <= not a or b;
    layer2_outputs(4486) <= a;
    layer2_outputs(4487) <= a or b;
    layer2_outputs(4488) <= not a;
    layer2_outputs(4489) <= not (a xor b);
    layer2_outputs(4490) <= b and not a;
    layer2_outputs(4491) <= b and not a;
    layer2_outputs(4492) <= not b;
    layer2_outputs(4493) <= not (a xor b);
    layer2_outputs(4494) <= not (a or b);
    layer2_outputs(4495) <= a;
    layer2_outputs(4496) <= not b or a;
    layer2_outputs(4497) <= not b or a;
    layer2_outputs(4498) <= 1'b1;
    layer2_outputs(4499) <= not (a and b);
    layer2_outputs(4500) <= not (a xor b);
    layer2_outputs(4501) <= a;
    layer2_outputs(4502) <= not (a xor b);
    layer2_outputs(4503) <= a;
    layer2_outputs(4504) <= not a or b;
    layer2_outputs(4505) <= not b or a;
    layer2_outputs(4506) <= b and not a;
    layer2_outputs(4507) <= not b or a;
    layer2_outputs(4508) <= not (a xor b);
    layer2_outputs(4509) <= a;
    layer2_outputs(4510) <= not (a xor b);
    layer2_outputs(4511) <= not b;
    layer2_outputs(4512) <= not (a or b);
    layer2_outputs(4513) <= not (a or b);
    layer2_outputs(4514) <= not b;
    layer2_outputs(4515) <= b;
    layer2_outputs(4516) <= a;
    layer2_outputs(4517) <= b and not a;
    layer2_outputs(4518) <= not (a xor b);
    layer2_outputs(4519) <= not a;
    layer2_outputs(4520) <= not b;
    layer2_outputs(4521) <= not a;
    layer2_outputs(4522) <= a xor b;
    layer2_outputs(4523) <= a and b;
    layer2_outputs(4524) <= not b;
    layer2_outputs(4525) <= a;
    layer2_outputs(4526) <= not (a or b);
    layer2_outputs(4527) <= b;
    layer2_outputs(4528) <= not b;
    layer2_outputs(4529) <= b and not a;
    layer2_outputs(4530) <= not a;
    layer2_outputs(4531) <= not a;
    layer2_outputs(4532) <= not a;
    layer2_outputs(4533) <= b;
    layer2_outputs(4534) <= a or b;
    layer2_outputs(4535) <= not (a or b);
    layer2_outputs(4536) <= b and not a;
    layer2_outputs(4537) <= b;
    layer2_outputs(4538) <= not a or b;
    layer2_outputs(4539) <= not (a xor b);
    layer2_outputs(4540) <= a and not b;
    layer2_outputs(4541) <= a xor b;
    layer2_outputs(4542) <= a and b;
    layer2_outputs(4543) <= b;
    layer2_outputs(4544) <= a or b;
    layer2_outputs(4545) <= not (a xor b);
    layer2_outputs(4546) <= not a;
    layer2_outputs(4547) <= not b;
    layer2_outputs(4548) <= not b or a;
    layer2_outputs(4549) <= not (a xor b);
    layer2_outputs(4550) <= not b or a;
    layer2_outputs(4551) <= a and b;
    layer2_outputs(4552) <= not b or a;
    layer2_outputs(4553) <= not a;
    layer2_outputs(4554) <= not b;
    layer2_outputs(4555) <= not (a or b);
    layer2_outputs(4556) <= not (a and b);
    layer2_outputs(4557) <= a or b;
    layer2_outputs(4558) <= not b;
    layer2_outputs(4559) <= a or b;
    layer2_outputs(4560) <= 1'b0;
    layer2_outputs(4561) <= not a;
    layer2_outputs(4562) <= b;
    layer2_outputs(4563) <= b;
    layer2_outputs(4564) <= not (a or b);
    layer2_outputs(4565) <= a;
    layer2_outputs(4566) <= b;
    layer2_outputs(4567) <= a xor b;
    layer2_outputs(4568) <= a xor b;
    layer2_outputs(4569) <= a and not b;
    layer2_outputs(4570) <= a and not b;
    layer2_outputs(4571) <= a;
    layer2_outputs(4572) <= b and not a;
    layer2_outputs(4573) <= not b;
    layer2_outputs(4574) <= not (a xor b);
    layer2_outputs(4575) <= a and not b;
    layer2_outputs(4576) <= not (a xor b);
    layer2_outputs(4577) <= b and not a;
    layer2_outputs(4578) <= not b or a;
    layer2_outputs(4579) <= a;
    layer2_outputs(4580) <= not a;
    layer2_outputs(4581) <= a and not b;
    layer2_outputs(4582) <= a and b;
    layer2_outputs(4583) <= b and not a;
    layer2_outputs(4584) <= b;
    layer2_outputs(4585) <= a xor b;
    layer2_outputs(4586) <= not b;
    layer2_outputs(4587) <= not b or a;
    layer2_outputs(4588) <= not b;
    layer2_outputs(4589) <= not a;
    layer2_outputs(4590) <= a;
    layer2_outputs(4591) <= not (a xor b);
    layer2_outputs(4592) <= a;
    layer2_outputs(4593) <= b and not a;
    layer2_outputs(4594) <= a and not b;
    layer2_outputs(4595) <= a and b;
    layer2_outputs(4596) <= a;
    layer2_outputs(4597) <= a and not b;
    layer2_outputs(4598) <= not a;
    layer2_outputs(4599) <= not b;
    layer2_outputs(4600) <= b;
    layer2_outputs(4601) <= a;
    layer2_outputs(4602) <= a and not b;
    layer2_outputs(4603) <= not a or b;
    layer2_outputs(4604) <= not a or b;
    layer2_outputs(4605) <= a and not b;
    layer2_outputs(4606) <= not b;
    layer2_outputs(4607) <= not (a or b);
    layer2_outputs(4608) <= b;
    layer2_outputs(4609) <= a;
    layer2_outputs(4610) <= not b or a;
    layer2_outputs(4611) <= a xor b;
    layer2_outputs(4612) <= not (a and b);
    layer2_outputs(4613) <= a or b;
    layer2_outputs(4614) <= b;
    layer2_outputs(4615) <= a and not b;
    layer2_outputs(4616) <= a xor b;
    layer2_outputs(4617) <= a xor b;
    layer2_outputs(4618) <= a and b;
    layer2_outputs(4619) <= not (a xor b);
    layer2_outputs(4620) <= not a;
    layer2_outputs(4621) <= not b;
    layer2_outputs(4622) <= not b;
    layer2_outputs(4623) <= not a or b;
    layer2_outputs(4624) <= b and not a;
    layer2_outputs(4625) <= b and not a;
    layer2_outputs(4626) <= a;
    layer2_outputs(4627) <= b and not a;
    layer2_outputs(4628) <= b and not a;
    layer2_outputs(4629) <= a or b;
    layer2_outputs(4630) <= not (a or b);
    layer2_outputs(4631) <= not (a or b);
    layer2_outputs(4632) <= a;
    layer2_outputs(4633) <= not (a xor b);
    layer2_outputs(4634) <= a xor b;
    layer2_outputs(4635) <= b;
    layer2_outputs(4636) <= not a;
    layer2_outputs(4637) <= a and not b;
    layer2_outputs(4638) <= not a or b;
    layer2_outputs(4639) <= a xor b;
    layer2_outputs(4640) <= not b;
    layer2_outputs(4641) <= not (a and b);
    layer2_outputs(4642) <= not a;
    layer2_outputs(4643) <= not (a and b);
    layer2_outputs(4644) <= a and not b;
    layer2_outputs(4645) <= a;
    layer2_outputs(4646) <= not b or a;
    layer2_outputs(4647) <= not (a xor b);
    layer2_outputs(4648) <= not (a xor b);
    layer2_outputs(4649) <= not a;
    layer2_outputs(4650) <= not a or b;
    layer2_outputs(4651) <= a or b;
    layer2_outputs(4652) <= not b or a;
    layer2_outputs(4653) <= a;
    layer2_outputs(4654) <= not b or a;
    layer2_outputs(4655) <= a;
    layer2_outputs(4656) <= not (a xor b);
    layer2_outputs(4657) <= not (a xor b);
    layer2_outputs(4658) <= a and b;
    layer2_outputs(4659) <= not a or b;
    layer2_outputs(4660) <= a and b;
    layer2_outputs(4661) <= b;
    layer2_outputs(4662) <= not a;
    layer2_outputs(4663) <= not (a or b);
    layer2_outputs(4664) <= b and not a;
    layer2_outputs(4665) <= 1'b0;
    layer2_outputs(4666) <= a;
    layer2_outputs(4667) <= not a or b;
    layer2_outputs(4668) <= not (a xor b);
    layer2_outputs(4669) <= a and b;
    layer2_outputs(4670) <= a or b;
    layer2_outputs(4671) <= not (a xor b);
    layer2_outputs(4672) <= a and b;
    layer2_outputs(4673) <= a or b;
    layer2_outputs(4674) <= a;
    layer2_outputs(4675) <= not b;
    layer2_outputs(4676) <= not (a xor b);
    layer2_outputs(4677) <= not b or a;
    layer2_outputs(4678) <= a;
    layer2_outputs(4679) <= a xor b;
    layer2_outputs(4680) <= not (a xor b);
    layer2_outputs(4681) <= b and not a;
    layer2_outputs(4682) <= not (a and b);
    layer2_outputs(4683) <= a xor b;
    layer2_outputs(4684) <= not (a xor b);
    layer2_outputs(4685) <= not a;
    layer2_outputs(4686) <= not (a or b);
    layer2_outputs(4687) <= b and not a;
    layer2_outputs(4688) <= not a;
    layer2_outputs(4689) <= not (a xor b);
    layer2_outputs(4690) <= not a or b;
    layer2_outputs(4691) <= b;
    layer2_outputs(4692) <= not b;
    layer2_outputs(4693) <= not b;
    layer2_outputs(4694) <= a;
    layer2_outputs(4695) <= a or b;
    layer2_outputs(4696) <= b and not a;
    layer2_outputs(4697) <= not a;
    layer2_outputs(4698) <= a or b;
    layer2_outputs(4699) <= a or b;
    layer2_outputs(4700) <= not b;
    layer2_outputs(4701) <= b and not a;
    layer2_outputs(4702) <= b;
    layer2_outputs(4703) <= not (a xor b);
    layer2_outputs(4704) <= not (a and b);
    layer2_outputs(4705) <= b and not a;
    layer2_outputs(4706) <= a and not b;
    layer2_outputs(4707) <= a;
    layer2_outputs(4708) <= 1'b1;
    layer2_outputs(4709) <= b;
    layer2_outputs(4710) <= not b;
    layer2_outputs(4711) <= a;
    layer2_outputs(4712) <= not a or b;
    layer2_outputs(4713) <= not a or b;
    layer2_outputs(4714) <= not b;
    layer2_outputs(4715) <= a and b;
    layer2_outputs(4716) <= a and not b;
    layer2_outputs(4717) <= not (a or b);
    layer2_outputs(4718) <= b;
    layer2_outputs(4719) <= not (a and b);
    layer2_outputs(4720) <= a and not b;
    layer2_outputs(4721) <= not (a and b);
    layer2_outputs(4722) <= not b;
    layer2_outputs(4723) <= not (a xor b);
    layer2_outputs(4724) <= not b;
    layer2_outputs(4725) <= a and b;
    layer2_outputs(4726) <= not a;
    layer2_outputs(4727) <= not (a and b);
    layer2_outputs(4728) <= b and not a;
    layer2_outputs(4729) <= not a;
    layer2_outputs(4730) <= not b or a;
    layer2_outputs(4731) <= not a;
    layer2_outputs(4732) <= not b;
    layer2_outputs(4733) <= a and not b;
    layer2_outputs(4734) <= not (a xor b);
    layer2_outputs(4735) <= not (a and b);
    layer2_outputs(4736) <= a or b;
    layer2_outputs(4737) <= b and not a;
    layer2_outputs(4738) <= b and not a;
    layer2_outputs(4739) <= not a or b;
    layer2_outputs(4740) <= a;
    layer2_outputs(4741) <= not (a xor b);
    layer2_outputs(4742) <= a and not b;
    layer2_outputs(4743) <= a;
    layer2_outputs(4744) <= not (a xor b);
    layer2_outputs(4745) <= not b;
    layer2_outputs(4746) <= a xor b;
    layer2_outputs(4747) <= a;
    layer2_outputs(4748) <= not a;
    layer2_outputs(4749) <= not b or a;
    layer2_outputs(4750) <= a or b;
    layer2_outputs(4751) <= not a;
    layer2_outputs(4752) <= a;
    layer2_outputs(4753) <= a and b;
    layer2_outputs(4754) <= 1'b1;
    layer2_outputs(4755) <= not b;
    layer2_outputs(4756) <= a xor b;
    layer2_outputs(4757) <= a or b;
    layer2_outputs(4758) <= a or b;
    layer2_outputs(4759) <= not b or a;
    layer2_outputs(4760) <= a xor b;
    layer2_outputs(4761) <= a and not b;
    layer2_outputs(4762) <= a xor b;
    layer2_outputs(4763) <= not b or a;
    layer2_outputs(4764) <= a;
    layer2_outputs(4765) <= not b;
    layer2_outputs(4766) <= not b;
    layer2_outputs(4767) <= not (a xor b);
    layer2_outputs(4768) <= not (a xor b);
    layer2_outputs(4769) <= not (a or b);
    layer2_outputs(4770) <= a and b;
    layer2_outputs(4771) <= not b;
    layer2_outputs(4772) <= b;
    layer2_outputs(4773) <= not b;
    layer2_outputs(4774) <= not b;
    layer2_outputs(4775) <= not b or a;
    layer2_outputs(4776) <= not a or b;
    layer2_outputs(4777) <= not b;
    layer2_outputs(4778) <= not (a or b);
    layer2_outputs(4779) <= not a or b;
    layer2_outputs(4780) <= not (a and b);
    layer2_outputs(4781) <= b and not a;
    layer2_outputs(4782) <= a or b;
    layer2_outputs(4783) <= not b;
    layer2_outputs(4784) <= not (a and b);
    layer2_outputs(4785) <= a and not b;
    layer2_outputs(4786) <= not b or a;
    layer2_outputs(4787) <= not b;
    layer2_outputs(4788) <= a xor b;
    layer2_outputs(4789) <= not a;
    layer2_outputs(4790) <= not (a and b);
    layer2_outputs(4791) <= not b;
    layer2_outputs(4792) <= not a;
    layer2_outputs(4793) <= not (a xor b);
    layer2_outputs(4794) <= not a or b;
    layer2_outputs(4795) <= not (a or b);
    layer2_outputs(4796) <= b;
    layer2_outputs(4797) <= a xor b;
    layer2_outputs(4798) <= not a;
    layer2_outputs(4799) <= b;
    layer2_outputs(4800) <= not b;
    layer2_outputs(4801) <= b;
    layer2_outputs(4802) <= a;
    layer2_outputs(4803) <= a and b;
    layer2_outputs(4804) <= b and not a;
    layer2_outputs(4805) <= b;
    layer2_outputs(4806) <= not (a xor b);
    layer2_outputs(4807) <= a and b;
    layer2_outputs(4808) <= not a;
    layer2_outputs(4809) <= a and not b;
    layer2_outputs(4810) <= a xor b;
    layer2_outputs(4811) <= not a or b;
    layer2_outputs(4812) <= not (a or b);
    layer2_outputs(4813) <= not a;
    layer2_outputs(4814) <= b;
    layer2_outputs(4815) <= b and not a;
    layer2_outputs(4816) <= a;
    layer2_outputs(4817) <= not b;
    layer2_outputs(4818) <= not (a xor b);
    layer2_outputs(4819) <= not b or a;
    layer2_outputs(4820) <= a and not b;
    layer2_outputs(4821) <= not a;
    layer2_outputs(4822) <= not (a or b);
    layer2_outputs(4823) <= a xor b;
    layer2_outputs(4824) <= not (a xor b);
    layer2_outputs(4825) <= not a;
    layer2_outputs(4826) <= b;
    layer2_outputs(4827) <= a and b;
    layer2_outputs(4828) <= not a;
    layer2_outputs(4829) <= not a or b;
    layer2_outputs(4830) <= not a or b;
    layer2_outputs(4831) <= not a or b;
    layer2_outputs(4832) <= a or b;
    layer2_outputs(4833) <= a;
    layer2_outputs(4834) <= not (a xor b);
    layer2_outputs(4835) <= not a or b;
    layer2_outputs(4836) <= not b;
    layer2_outputs(4837) <= not (a or b);
    layer2_outputs(4838) <= not (a or b);
    layer2_outputs(4839) <= not b;
    layer2_outputs(4840) <= not (a xor b);
    layer2_outputs(4841) <= not a or b;
    layer2_outputs(4842) <= a;
    layer2_outputs(4843) <= not (a and b);
    layer2_outputs(4844) <= not b;
    layer2_outputs(4845) <= not b or a;
    layer2_outputs(4846) <= b and not a;
    layer2_outputs(4847) <= a xor b;
    layer2_outputs(4848) <= not a;
    layer2_outputs(4849) <= not b or a;
    layer2_outputs(4850) <= a;
    layer2_outputs(4851) <= not a or b;
    layer2_outputs(4852) <= b and not a;
    layer2_outputs(4853) <= not a;
    layer2_outputs(4854) <= not b;
    layer2_outputs(4855) <= not a or b;
    layer2_outputs(4856) <= not b or a;
    layer2_outputs(4857) <= not b;
    layer2_outputs(4858) <= a xor b;
    layer2_outputs(4859) <= a and not b;
    layer2_outputs(4860) <= a and not b;
    layer2_outputs(4861) <= a;
    layer2_outputs(4862) <= not a;
    layer2_outputs(4863) <= not b or a;
    layer2_outputs(4864) <= b and not a;
    layer2_outputs(4865) <= not b or a;
    layer2_outputs(4866) <= not b;
    layer2_outputs(4867) <= a;
    layer2_outputs(4868) <= a xor b;
    layer2_outputs(4869) <= not b;
    layer2_outputs(4870) <= not (a xor b);
    layer2_outputs(4871) <= not (a and b);
    layer2_outputs(4872) <= not (a xor b);
    layer2_outputs(4873) <= a or b;
    layer2_outputs(4874) <= not (a xor b);
    layer2_outputs(4875) <= b;
    layer2_outputs(4876) <= a xor b;
    layer2_outputs(4877) <= a or b;
    layer2_outputs(4878) <= not a;
    layer2_outputs(4879) <= not b or a;
    layer2_outputs(4880) <= not (a or b);
    layer2_outputs(4881) <= not b or a;
    layer2_outputs(4882) <= b and not a;
    layer2_outputs(4883) <= not (a or b);
    layer2_outputs(4884) <= not (a xor b);
    layer2_outputs(4885) <= a xor b;
    layer2_outputs(4886) <= not b or a;
    layer2_outputs(4887) <= b;
    layer2_outputs(4888) <= not (a or b);
    layer2_outputs(4889) <= a and b;
    layer2_outputs(4890) <= a and b;
    layer2_outputs(4891) <= not (a and b);
    layer2_outputs(4892) <= a;
    layer2_outputs(4893) <= a and b;
    layer2_outputs(4894) <= not b;
    layer2_outputs(4895) <= not (a and b);
    layer2_outputs(4896) <= not (a or b);
    layer2_outputs(4897) <= 1'b1;
    layer2_outputs(4898) <= a or b;
    layer2_outputs(4899) <= a and b;
    layer2_outputs(4900) <= not (a and b);
    layer2_outputs(4901) <= not b;
    layer2_outputs(4902) <= not (a or b);
    layer2_outputs(4903) <= a and not b;
    layer2_outputs(4904) <= not b;
    layer2_outputs(4905) <= not b;
    layer2_outputs(4906) <= a;
    layer2_outputs(4907) <= b;
    layer2_outputs(4908) <= not (a xor b);
    layer2_outputs(4909) <= not b;
    layer2_outputs(4910) <= a;
    layer2_outputs(4911) <= a and b;
    layer2_outputs(4912) <= a xor b;
    layer2_outputs(4913) <= b and not a;
    layer2_outputs(4914) <= a and b;
    layer2_outputs(4915) <= not b or a;
    layer2_outputs(4916) <= b and not a;
    layer2_outputs(4917) <= not a;
    layer2_outputs(4918) <= b;
    layer2_outputs(4919) <= a and b;
    layer2_outputs(4920) <= not (a and b);
    layer2_outputs(4921) <= 1'b0;
    layer2_outputs(4922) <= a xor b;
    layer2_outputs(4923) <= a and not b;
    layer2_outputs(4924) <= not a;
    layer2_outputs(4925) <= not (a or b);
    layer2_outputs(4926) <= b;
    layer2_outputs(4927) <= b;
    layer2_outputs(4928) <= a xor b;
    layer2_outputs(4929) <= not (a and b);
    layer2_outputs(4930) <= b and not a;
    layer2_outputs(4931) <= b;
    layer2_outputs(4932) <= a xor b;
    layer2_outputs(4933) <= not b;
    layer2_outputs(4934) <= not a or b;
    layer2_outputs(4935) <= a and not b;
    layer2_outputs(4936) <= not a or b;
    layer2_outputs(4937) <= not a or b;
    layer2_outputs(4938) <= a and b;
    layer2_outputs(4939) <= not (a and b);
    layer2_outputs(4940) <= not b or a;
    layer2_outputs(4941) <= not b or a;
    layer2_outputs(4942) <= b;
    layer2_outputs(4943) <= a;
    layer2_outputs(4944) <= b and not a;
    layer2_outputs(4945) <= not (a or b);
    layer2_outputs(4946) <= b and not a;
    layer2_outputs(4947) <= not (a xor b);
    layer2_outputs(4948) <= a;
    layer2_outputs(4949) <= not (a xor b);
    layer2_outputs(4950) <= not b or a;
    layer2_outputs(4951) <= a or b;
    layer2_outputs(4952) <= b;
    layer2_outputs(4953) <= not b or a;
    layer2_outputs(4954) <= not a or b;
    layer2_outputs(4955) <= not b;
    layer2_outputs(4956) <= a and b;
    layer2_outputs(4957) <= a and not b;
    layer2_outputs(4958) <= not b;
    layer2_outputs(4959) <= b;
    layer2_outputs(4960) <= not a;
    layer2_outputs(4961) <= a;
    layer2_outputs(4962) <= a or b;
    layer2_outputs(4963) <= a xor b;
    layer2_outputs(4964) <= not (a xor b);
    layer2_outputs(4965) <= not b;
    layer2_outputs(4966) <= a;
    layer2_outputs(4967) <= a or b;
    layer2_outputs(4968) <= b;
    layer2_outputs(4969) <= not (a xor b);
    layer2_outputs(4970) <= not (a xor b);
    layer2_outputs(4971) <= a and not b;
    layer2_outputs(4972) <= b and not a;
    layer2_outputs(4973) <= not b or a;
    layer2_outputs(4974) <= a and not b;
    layer2_outputs(4975) <= not b;
    layer2_outputs(4976) <= not (a and b);
    layer2_outputs(4977) <= not b;
    layer2_outputs(4978) <= a xor b;
    layer2_outputs(4979) <= not (a xor b);
    layer2_outputs(4980) <= not b;
    layer2_outputs(4981) <= 1'b1;
    layer2_outputs(4982) <= a;
    layer2_outputs(4983) <= a;
    layer2_outputs(4984) <= not (a xor b);
    layer2_outputs(4985) <= not a or b;
    layer2_outputs(4986) <= a;
    layer2_outputs(4987) <= a and b;
    layer2_outputs(4988) <= a xor b;
    layer2_outputs(4989) <= a or b;
    layer2_outputs(4990) <= not b or a;
    layer2_outputs(4991) <= b and not a;
    layer2_outputs(4992) <= b;
    layer2_outputs(4993) <= not (a or b);
    layer2_outputs(4994) <= not b;
    layer2_outputs(4995) <= not b or a;
    layer2_outputs(4996) <= not b;
    layer2_outputs(4997) <= b and not a;
    layer2_outputs(4998) <= b;
    layer2_outputs(4999) <= not a;
    layer2_outputs(5000) <= not (a or b);
    layer2_outputs(5001) <= a;
    layer2_outputs(5002) <= a xor b;
    layer2_outputs(5003) <= a and not b;
    layer2_outputs(5004) <= not b;
    layer2_outputs(5005) <= a and b;
    layer2_outputs(5006) <= not (a and b);
    layer2_outputs(5007) <= a or b;
    layer2_outputs(5008) <= b;
    layer2_outputs(5009) <= not (a and b);
    layer2_outputs(5010) <= a or b;
    layer2_outputs(5011) <= b and not a;
    layer2_outputs(5012) <= a and not b;
    layer2_outputs(5013) <= not (a xor b);
    layer2_outputs(5014) <= a or b;
    layer2_outputs(5015) <= not b or a;
    layer2_outputs(5016) <= a and not b;
    layer2_outputs(5017) <= a xor b;
    layer2_outputs(5018) <= a or b;
    layer2_outputs(5019) <= not (a and b);
    layer2_outputs(5020) <= not b or a;
    layer2_outputs(5021) <= not (a and b);
    layer2_outputs(5022) <= a and b;
    layer2_outputs(5023) <= not a;
    layer2_outputs(5024) <= not a;
    layer2_outputs(5025) <= a xor b;
    layer2_outputs(5026) <= a and b;
    layer2_outputs(5027) <= not (a xor b);
    layer2_outputs(5028) <= b;
    layer2_outputs(5029) <= not a or b;
    layer2_outputs(5030) <= a and b;
    layer2_outputs(5031) <= not (a or b);
    layer2_outputs(5032) <= b;
    layer2_outputs(5033) <= not b;
    layer2_outputs(5034) <= a and b;
    layer2_outputs(5035) <= not (a xor b);
    layer2_outputs(5036) <= a or b;
    layer2_outputs(5037) <= not b;
    layer2_outputs(5038) <= not (a and b);
    layer2_outputs(5039) <= not a;
    layer2_outputs(5040) <= not b or a;
    layer2_outputs(5041) <= not (a xor b);
    layer2_outputs(5042) <= a;
    layer2_outputs(5043) <= not a;
    layer2_outputs(5044) <= not a;
    layer2_outputs(5045) <= a and not b;
    layer2_outputs(5046) <= not a;
    layer2_outputs(5047) <= a;
    layer2_outputs(5048) <= a;
    layer2_outputs(5049) <= a xor b;
    layer2_outputs(5050) <= not a;
    layer2_outputs(5051) <= not b or a;
    layer2_outputs(5052) <= b;
    layer2_outputs(5053) <= a and b;
    layer2_outputs(5054) <= not (a or b);
    layer2_outputs(5055) <= not (a xor b);
    layer2_outputs(5056) <= not (a and b);
    layer2_outputs(5057) <= not b;
    layer2_outputs(5058) <= not (a or b);
    layer2_outputs(5059) <= a or b;
    layer2_outputs(5060) <= b and not a;
    layer2_outputs(5061) <= a and b;
    layer2_outputs(5062) <= a;
    layer2_outputs(5063) <= not b or a;
    layer2_outputs(5064) <= not (a and b);
    layer2_outputs(5065) <= not (a and b);
    layer2_outputs(5066) <= a xor b;
    layer2_outputs(5067) <= not b or a;
    layer2_outputs(5068) <= a and not b;
    layer2_outputs(5069) <= a;
    layer2_outputs(5070) <= not b;
    layer2_outputs(5071) <= not (a or b);
    layer2_outputs(5072) <= not a;
    layer2_outputs(5073) <= b;
    layer2_outputs(5074) <= not (a or b);
    layer2_outputs(5075) <= not (a and b);
    layer2_outputs(5076) <= a or b;
    layer2_outputs(5077) <= a and not b;
    layer2_outputs(5078) <= b and not a;
    layer2_outputs(5079) <= not a;
    layer2_outputs(5080) <= not a;
    layer2_outputs(5081) <= b and not a;
    layer2_outputs(5082) <= a or b;
    layer2_outputs(5083) <= b;
    layer2_outputs(5084) <= not b or a;
    layer2_outputs(5085) <= not b or a;
    layer2_outputs(5086) <= a;
    layer2_outputs(5087) <= not (a xor b);
    layer2_outputs(5088) <= not a;
    layer2_outputs(5089) <= not b or a;
    layer2_outputs(5090) <= b and not a;
    layer2_outputs(5091) <= not a;
    layer2_outputs(5092) <= not b;
    layer2_outputs(5093) <= a xor b;
    layer2_outputs(5094) <= a or b;
    layer2_outputs(5095) <= not a or b;
    layer2_outputs(5096) <= b and not a;
    layer2_outputs(5097) <= a or b;
    layer2_outputs(5098) <= b;
    layer2_outputs(5099) <= a and not b;
    layer2_outputs(5100) <= a and not b;
    layer2_outputs(5101) <= b;
    layer2_outputs(5102) <= not b;
    layer2_outputs(5103) <= a and not b;
    layer2_outputs(5104) <= not (a and b);
    layer2_outputs(5105) <= a and b;
    layer2_outputs(5106) <= not b or a;
    layer2_outputs(5107) <= b;
    layer2_outputs(5108) <= a or b;
    layer2_outputs(5109) <= not a or b;
    layer2_outputs(5110) <= a or b;
    layer2_outputs(5111) <= a xor b;
    layer2_outputs(5112) <= a;
    layer2_outputs(5113) <= not a;
    layer2_outputs(5114) <= a xor b;
    layer2_outputs(5115) <= not a or b;
    layer2_outputs(5116) <= b;
    layer2_outputs(5117) <= not a or b;
    layer2_outputs(5118) <= not b;
    layer2_outputs(5119) <= a xor b;
    layer2_outputs(5120) <= a xor b;
    layer2_outputs(5121) <= b and not a;
    layer2_outputs(5122) <= not (a xor b);
    layer2_outputs(5123) <= a;
    layer2_outputs(5124) <= not (a xor b);
    layer2_outputs(5125) <= 1'b0;
    layer2_outputs(5126) <= not (a xor b);
    layer2_outputs(5127) <= not (a and b);
    layer2_outputs(5128) <= a;
    layer2_outputs(5129) <= not (a xor b);
    layer2_outputs(5130) <= a;
    layer2_outputs(5131) <= a and not b;
    layer2_outputs(5132) <= not a or b;
    layer2_outputs(5133) <= 1'b1;
    layer2_outputs(5134) <= b;
    layer2_outputs(5135) <= a xor b;
    layer2_outputs(5136) <= a and not b;
    layer2_outputs(5137) <= not b or a;
    layer2_outputs(5138) <= b and not a;
    layer2_outputs(5139) <= b and not a;
    layer2_outputs(5140) <= not b;
    layer2_outputs(5141) <= b and not a;
    layer2_outputs(5142) <= b and not a;
    layer2_outputs(5143) <= not a or b;
    layer2_outputs(5144) <= not a or b;
    layer2_outputs(5145) <= not (a xor b);
    layer2_outputs(5146) <= a and b;
    layer2_outputs(5147) <= b and not a;
    layer2_outputs(5148) <= not b;
    layer2_outputs(5149) <= not b;
    layer2_outputs(5150) <= a;
    layer2_outputs(5151) <= b and not a;
    layer2_outputs(5152) <= not (a xor b);
    layer2_outputs(5153) <= a and not b;
    layer2_outputs(5154) <= a or b;
    layer2_outputs(5155) <= not (a and b);
    layer2_outputs(5156) <= not b;
    layer2_outputs(5157) <= a or b;
    layer2_outputs(5158) <= not b;
    layer2_outputs(5159) <= not b;
    layer2_outputs(5160) <= a and b;
    layer2_outputs(5161) <= a;
    layer2_outputs(5162) <= a or b;
    layer2_outputs(5163) <= not (a xor b);
    layer2_outputs(5164) <= not a;
    layer2_outputs(5165) <= not (a or b);
    layer2_outputs(5166) <= not a or b;
    layer2_outputs(5167) <= b;
    layer2_outputs(5168) <= not b;
    layer2_outputs(5169) <= not b;
    layer2_outputs(5170) <= b and not a;
    layer2_outputs(5171) <= a;
    layer2_outputs(5172) <= a or b;
    layer2_outputs(5173) <= b and not a;
    layer2_outputs(5174) <= not b;
    layer2_outputs(5175) <= a or b;
    layer2_outputs(5176) <= b and not a;
    layer2_outputs(5177) <= not a;
    layer2_outputs(5178) <= not (a xor b);
    layer2_outputs(5179) <= not (a or b);
    layer2_outputs(5180) <= 1'b0;
    layer2_outputs(5181) <= not (a and b);
    layer2_outputs(5182) <= a or b;
    layer2_outputs(5183) <= not a or b;
    layer2_outputs(5184) <= not (a or b);
    layer2_outputs(5185) <= not (a xor b);
    layer2_outputs(5186) <= not a or b;
    layer2_outputs(5187) <= not (a and b);
    layer2_outputs(5188) <= a or b;
    layer2_outputs(5189) <= a xor b;
    layer2_outputs(5190) <= not b;
    layer2_outputs(5191) <= a or b;
    layer2_outputs(5192) <= not a;
    layer2_outputs(5193) <= not (a or b);
    layer2_outputs(5194) <= a xor b;
    layer2_outputs(5195) <= a and b;
    layer2_outputs(5196) <= not b;
    layer2_outputs(5197) <= not (a and b);
    layer2_outputs(5198) <= b and not a;
    layer2_outputs(5199) <= not (a xor b);
    layer2_outputs(5200) <= a xor b;
    layer2_outputs(5201) <= not a;
    layer2_outputs(5202) <= b;
    layer2_outputs(5203) <= a xor b;
    layer2_outputs(5204) <= a;
    layer2_outputs(5205) <= a;
    layer2_outputs(5206) <= a;
    layer2_outputs(5207) <= b;
    layer2_outputs(5208) <= not (a and b);
    layer2_outputs(5209) <= not (a and b);
    layer2_outputs(5210) <= b;
    layer2_outputs(5211) <= not a;
    layer2_outputs(5212) <= a;
    layer2_outputs(5213) <= a and b;
    layer2_outputs(5214) <= not a or b;
    layer2_outputs(5215) <= not a or b;
    layer2_outputs(5216) <= b and not a;
    layer2_outputs(5217) <= a and b;
    layer2_outputs(5218) <= not (a xor b);
    layer2_outputs(5219) <= not a or b;
    layer2_outputs(5220) <= not a;
    layer2_outputs(5221) <= b and not a;
    layer2_outputs(5222) <= not (a and b);
    layer2_outputs(5223) <= a;
    layer2_outputs(5224) <= b and not a;
    layer2_outputs(5225) <= not b;
    layer2_outputs(5226) <= not b or a;
    layer2_outputs(5227) <= b and not a;
    layer2_outputs(5228) <= not b;
    layer2_outputs(5229) <= a;
    layer2_outputs(5230) <= a;
    layer2_outputs(5231) <= a or b;
    layer2_outputs(5232) <= a or b;
    layer2_outputs(5233) <= not b;
    layer2_outputs(5234) <= not a;
    layer2_outputs(5235) <= a xor b;
    layer2_outputs(5236) <= not (a and b);
    layer2_outputs(5237) <= not b;
    layer2_outputs(5238) <= not a;
    layer2_outputs(5239) <= not b;
    layer2_outputs(5240) <= not (a xor b);
    layer2_outputs(5241) <= not a;
    layer2_outputs(5242) <= b;
    layer2_outputs(5243) <= not a or b;
    layer2_outputs(5244) <= a and b;
    layer2_outputs(5245) <= not b or a;
    layer2_outputs(5246) <= not a;
    layer2_outputs(5247) <= a;
    layer2_outputs(5248) <= b;
    layer2_outputs(5249) <= b;
    layer2_outputs(5250) <= a and b;
    layer2_outputs(5251) <= not (a and b);
    layer2_outputs(5252) <= not (a or b);
    layer2_outputs(5253) <= a and b;
    layer2_outputs(5254) <= not (a or b);
    layer2_outputs(5255) <= not b;
    layer2_outputs(5256) <= b;
    layer2_outputs(5257) <= b;
    layer2_outputs(5258) <= not (a xor b);
    layer2_outputs(5259) <= a;
    layer2_outputs(5260) <= a and b;
    layer2_outputs(5261) <= b;
    layer2_outputs(5262) <= not a or b;
    layer2_outputs(5263) <= not b;
    layer2_outputs(5264) <= a and not b;
    layer2_outputs(5265) <= a xor b;
    layer2_outputs(5266) <= not b;
    layer2_outputs(5267) <= a and b;
    layer2_outputs(5268) <= b;
    layer2_outputs(5269) <= 1'b0;
    layer2_outputs(5270) <= a and b;
    layer2_outputs(5271) <= a xor b;
    layer2_outputs(5272) <= not b;
    layer2_outputs(5273) <= b;
    layer2_outputs(5274) <= a or b;
    layer2_outputs(5275) <= not (a and b);
    layer2_outputs(5276) <= a;
    layer2_outputs(5277) <= a and b;
    layer2_outputs(5278) <= b;
    layer2_outputs(5279) <= not (a xor b);
    layer2_outputs(5280) <= not (a xor b);
    layer2_outputs(5281) <= a and not b;
    layer2_outputs(5282) <= a xor b;
    layer2_outputs(5283) <= 1'b1;
    layer2_outputs(5284) <= b;
    layer2_outputs(5285) <= b;
    layer2_outputs(5286) <= not (a and b);
    layer2_outputs(5287) <= a and not b;
    layer2_outputs(5288) <= not (a or b);
    layer2_outputs(5289) <= a and not b;
    layer2_outputs(5290) <= a xor b;
    layer2_outputs(5291) <= not (a xor b);
    layer2_outputs(5292) <= a;
    layer2_outputs(5293) <= not a or b;
    layer2_outputs(5294) <= b;
    layer2_outputs(5295) <= not a or b;
    layer2_outputs(5296) <= not b;
    layer2_outputs(5297) <= not a;
    layer2_outputs(5298) <= a and b;
    layer2_outputs(5299) <= not a;
    layer2_outputs(5300) <= a or b;
    layer2_outputs(5301) <= b;
    layer2_outputs(5302) <= not b or a;
    layer2_outputs(5303) <= a and b;
    layer2_outputs(5304) <= not a;
    layer2_outputs(5305) <= a;
    layer2_outputs(5306) <= not (a and b);
    layer2_outputs(5307) <= not (a and b);
    layer2_outputs(5308) <= a and not b;
    layer2_outputs(5309) <= a xor b;
    layer2_outputs(5310) <= a or b;
    layer2_outputs(5311) <= a xor b;
    layer2_outputs(5312) <= a;
    layer2_outputs(5313) <= not a;
    layer2_outputs(5314) <= b and not a;
    layer2_outputs(5315) <= not b;
    layer2_outputs(5316) <= not (a and b);
    layer2_outputs(5317) <= not a;
    layer2_outputs(5318) <= not (a or b);
    layer2_outputs(5319) <= not (a and b);
    layer2_outputs(5320) <= not (a or b);
    layer2_outputs(5321) <= a xor b;
    layer2_outputs(5322) <= not a or b;
    layer2_outputs(5323) <= not b;
    layer2_outputs(5324) <= b;
    layer2_outputs(5325) <= 1'b0;
    layer2_outputs(5326) <= a and not b;
    layer2_outputs(5327) <= a and b;
    layer2_outputs(5328) <= a and not b;
    layer2_outputs(5329) <= a or b;
    layer2_outputs(5330) <= a xor b;
    layer2_outputs(5331) <= b;
    layer2_outputs(5332) <= a xor b;
    layer2_outputs(5333) <= a and not b;
    layer2_outputs(5334) <= b;
    layer2_outputs(5335) <= a xor b;
    layer2_outputs(5336) <= not (a xor b);
    layer2_outputs(5337) <= not b;
    layer2_outputs(5338) <= not b;
    layer2_outputs(5339) <= not (a xor b);
    layer2_outputs(5340) <= not a or b;
    layer2_outputs(5341) <= b and not a;
    layer2_outputs(5342) <= not b or a;
    layer2_outputs(5343) <= not a or b;
    layer2_outputs(5344) <= not (a xor b);
    layer2_outputs(5345) <= b;
    layer2_outputs(5346) <= not a or b;
    layer2_outputs(5347) <= a xor b;
    layer2_outputs(5348) <= a xor b;
    layer2_outputs(5349) <= not a;
    layer2_outputs(5350) <= a and b;
    layer2_outputs(5351) <= not (a xor b);
    layer2_outputs(5352) <= b and not a;
    layer2_outputs(5353) <= not a;
    layer2_outputs(5354) <= not (a or b);
    layer2_outputs(5355) <= not (a and b);
    layer2_outputs(5356) <= b and not a;
    layer2_outputs(5357) <= not (a or b);
    layer2_outputs(5358) <= not (a and b);
    layer2_outputs(5359) <= b and not a;
    layer2_outputs(5360) <= not b or a;
    layer2_outputs(5361) <= a and not b;
    layer2_outputs(5362) <= a;
    layer2_outputs(5363) <= not (a and b);
    layer2_outputs(5364) <= b and not a;
    layer2_outputs(5365) <= b;
    layer2_outputs(5366) <= not (a or b);
    layer2_outputs(5367) <= not a or b;
    layer2_outputs(5368) <= not (a xor b);
    layer2_outputs(5369) <= not b;
    layer2_outputs(5370) <= a;
    layer2_outputs(5371) <= not a or b;
    layer2_outputs(5372) <= not (a xor b);
    layer2_outputs(5373) <= 1'b0;
    layer2_outputs(5374) <= b;
    layer2_outputs(5375) <= not (a and b);
    layer2_outputs(5376) <= not b or a;
    layer2_outputs(5377) <= not a or b;
    layer2_outputs(5378) <= a and b;
    layer2_outputs(5379) <= b;
    layer2_outputs(5380) <= not b;
    layer2_outputs(5381) <= not b or a;
    layer2_outputs(5382) <= not (a or b);
    layer2_outputs(5383) <= not b;
    layer2_outputs(5384) <= b;
    layer2_outputs(5385) <= a;
    layer2_outputs(5386) <= not (a and b);
    layer2_outputs(5387) <= not b;
    layer2_outputs(5388) <= not a;
    layer2_outputs(5389) <= a or b;
    layer2_outputs(5390) <= not (a xor b);
    layer2_outputs(5391) <= not a;
    layer2_outputs(5392) <= b;
    layer2_outputs(5393) <= a and not b;
    layer2_outputs(5394) <= a and not b;
    layer2_outputs(5395) <= not a;
    layer2_outputs(5396) <= not (a and b);
    layer2_outputs(5397) <= not (a or b);
    layer2_outputs(5398) <= not a or b;
    layer2_outputs(5399) <= not a;
    layer2_outputs(5400) <= a or b;
    layer2_outputs(5401) <= not b;
    layer2_outputs(5402) <= not a;
    layer2_outputs(5403) <= not a;
    layer2_outputs(5404) <= a or b;
    layer2_outputs(5405) <= not b;
    layer2_outputs(5406) <= b;
    layer2_outputs(5407) <= not (a xor b);
    layer2_outputs(5408) <= not b;
    layer2_outputs(5409) <= b and not a;
    layer2_outputs(5410) <= not a or b;
    layer2_outputs(5411) <= a or b;
    layer2_outputs(5412) <= a and not b;
    layer2_outputs(5413) <= a or b;
    layer2_outputs(5414) <= a xor b;
    layer2_outputs(5415) <= not b;
    layer2_outputs(5416) <= not (a and b);
    layer2_outputs(5417) <= not (a xor b);
    layer2_outputs(5418) <= a;
    layer2_outputs(5419) <= a and b;
    layer2_outputs(5420) <= not a;
    layer2_outputs(5421) <= not a;
    layer2_outputs(5422) <= not (a and b);
    layer2_outputs(5423) <= a and b;
    layer2_outputs(5424) <= not (a or b);
    layer2_outputs(5425) <= not (a xor b);
    layer2_outputs(5426) <= a and b;
    layer2_outputs(5427) <= a or b;
    layer2_outputs(5428) <= a and b;
    layer2_outputs(5429) <= a and b;
    layer2_outputs(5430) <= not a;
    layer2_outputs(5431) <= b and not a;
    layer2_outputs(5432) <= not (a or b);
    layer2_outputs(5433) <= not (a or b);
    layer2_outputs(5434) <= not (a and b);
    layer2_outputs(5435) <= a and not b;
    layer2_outputs(5436) <= not a or b;
    layer2_outputs(5437) <= not a;
    layer2_outputs(5438) <= not b;
    layer2_outputs(5439) <= not (a xor b);
    layer2_outputs(5440) <= not a;
    layer2_outputs(5441) <= not a;
    layer2_outputs(5442) <= b;
    layer2_outputs(5443) <= b and not a;
    layer2_outputs(5444) <= b;
    layer2_outputs(5445) <= a xor b;
    layer2_outputs(5446) <= not a;
    layer2_outputs(5447) <= not b;
    layer2_outputs(5448) <= not (a xor b);
    layer2_outputs(5449) <= not a;
    layer2_outputs(5450) <= a and not b;
    layer2_outputs(5451) <= not a;
    layer2_outputs(5452) <= not (a and b);
    layer2_outputs(5453) <= a;
    layer2_outputs(5454) <= a and b;
    layer2_outputs(5455) <= a xor b;
    layer2_outputs(5456) <= not b or a;
    layer2_outputs(5457) <= not (a and b);
    layer2_outputs(5458) <= a and not b;
    layer2_outputs(5459) <= a;
    layer2_outputs(5460) <= b and not a;
    layer2_outputs(5461) <= not a;
    layer2_outputs(5462) <= a and b;
    layer2_outputs(5463) <= not a;
    layer2_outputs(5464) <= not a;
    layer2_outputs(5465) <= not (a xor b);
    layer2_outputs(5466) <= a;
    layer2_outputs(5467) <= not a;
    layer2_outputs(5468) <= not b;
    layer2_outputs(5469) <= not a;
    layer2_outputs(5470) <= not (a xor b);
    layer2_outputs(5471) <= not b;
    layer2_outputs(5472) <= b;
    layer2_outputs(5473) <= not (a xor b);
    layer2_outputs(5474) <= b;
    layer2_outputs(5475) <= not (a xor b);
    layer2_outputs(5476) <= a xor b;
    layer2_outputs(5477) <= not b;
    layer2_outputs(5478) <= a xor b;
    layer2_outputs(5479) <= not b;
    layer2_outputs(5480) <= a or b;
    layer2_outputs(5481) <= not (a and b);
    layer2_outputs(5482) <= a;
    layer2_outputs(5483) <= b;
    layer2_outputs(5484) <= a xor b;
    layer2_outputs(5485) <= not (a and b);
    layer2_outputs(5486) <= not a or b;
    layer2_outputs(5487) <= not a;
    layer2_outputs(5488) <= a;
    layer2_outputs(5489) <= a;
    layer2_outputs(5490) <= a;
    layer2_outputs(5491) <= not b or a;
    layer2_outputs(5492) <= a and not b;
    layer2_outputs(5493) <= a;
    layer2_outputs(5494) <= a or b;
    layer2_outputs(5495) <= not a or b;
    layer2_outputs(5496) <= not a;
    layer2_outputs(5497) <= not (a or b);
    layer2_outputs(5498) <= not (a and b);
    layer2_outputs(5499) <= not b;
    layer2_outputs(5500) <= a and b;
    layer2_outputs(5501) <= b;
    layer2_outputs(5502) <= a xor b;
    layer2_outputs(5503) <= a and not b;
    layer2_outputs(5504) <= a or b;
    layer2_outputs(5505) <= a;
    layer2_outputs(5506) <= a;
    layer2_outputs(5507) <= not (a or b);
    layer2_outputs(5508) <= not b or a;
    layer2_outputs(5509) <= not a;
    layer2_outputs(5510) <= 1'b1;
    layer2_outputs(5511) <= not b;
    layer2_outputs(5512) <= b and not a;
    layer2_outputs(5513) <= a and not b;
    layer2_outputs(5514) <= b;
    layer2_outputs(5515) <= not b;
    layer2_outputs(5516) <= b and not a;
    layer2_outputs(5517) <= not (a and b);
    layer2_outputs(5518) <= not a or b;
    layer2_outputs(5519) <= a or b;
    layer2_outputs(5520) <= not (a xor b);
    layer2_outputs(5521) <= not a;
    layer2_outputs(5522) <= not (a xor b);
    layer2_outputs(5523) <= not (a and b);
    layer2_outputs(5524) <= not (a xor b);
    layer2_outputs(5525) <= a xor b;
    layer2_outputs(5526) <= not b;
    layer2_outputs(5527) <= a;
    layer2_outputs(5528) <= not b;
    layer2_outputs(5529) <= not (a xor b);
    layer2_outputs(5530) <= not a;
    layer2_outputs(5531) <= a and b;
    layer2_outputs(5532) <= b;
    layer2_outputs(5533) <= a or b;
    layer2_outputs(5534) <= not (a and b);
    layer2_outputs(5535) <= a and b;
    layer2_outputs(5536) <= not a;
    layer2_outputs(5537) <= a xor b;
    layer2_outputs(5538) <= not (a and b);
    layer2_outputs(5539) <= not (a and b);
    layer2_outputs(5540) <= not (a xor b);
    layer2_outputs(5541) <= a and b;
    layer2_outputs(5542) <= not (a xor b);
    layer2_outputs(5543) <= not b or a;
    layer2_outputs(5544) <= a;
    layer2_outputs(5545) <= not a;
    layer2_outputs(5546) <= a and not b;
    layer2_outputs(5547) <= not a or b;
    layer2_outputs(5548) <= b;
    layer2_outputs(5549) <= b and not a;
    layer2_outputs(5550) <= a xor b;
    layer2_outputs(5551) <= not (a and b);
    layer2_outputs(5552) <= b;
    layer2_outputs(5553) <= not a;
    layer2_outputs(5554) <= a;
    layer2_outputs(5555) <= not a;
    layer2_outputs(5556) <= b;
    layer2_outputs(5557) <= b and not a;
    layer2_outputs(5558) <= b and not a;
    layer2_outputs(5559) <= 1'b0;
    layer2_outputs(5560) <= a;
    layer2_outputs(5561) <= not (a and b);
    layer2_outputs(5562) <= not (a xor b);
    layer2_outputs(5563) <= not b or a;
    layer2_outputs(5564) <= a and not b;
    layer2_outputs(5565) <= a and b;
    layer2_outputs(5566) <= a and b;
    layer2_outputs(5567) <= not (a xor b);
    layer2_outputs(5568) <= a or b;
    layer2_outputs(5569) <= a xor b;
    layer2_outputs(5570) <= a xor b;
    layer2_outputs(5571) <= a xor b;
    layer2_outputs(5572) <= a xor b;
    layer2_outputs(5573) <= a;
    layer2_outputs(5574) <= not (a or b);
    layer2_outputs(5575) <= a and not b;
    layer2_outputs(5576) <= not b;
    layer2_outputs(5577) <= not a;
    layer2_outputs(5578) <= b;
    layer2_outputs(5579) <= a;
    layer2_outputs(5580) <= a and not b;
    layer2_outputs(5581) <= not b or a;
    layer2_outputs(5582) <= b and not a;
    layer2_outputs(5583) <= not (a and b);
    layer2_outputs(5584) <= b and not a;
    layer2_outputs(5585) <= not b or a;
    layer2_outputs(5586) <= not (a and b);
    layer2_outputs(5587) <= not (a and b);
    layer2_outputs(5588) <= b;
    layer2_outputs(5589) <= a;
    layer2_outputs(5590) <= not (a and b);
    layer2_outputs(5591) <= a and b;
    layer2_outputs(5592) <= a;
    layer2_outputs(5593) <= a and not b;
    layer2_outputs(5594) <= a and not b;
    layer2_outputs(5595) <= not b or a;
    layer2_outputs(5596) <= a xor b;
    layer2_outputs(5597) <= b;
    layer2_outputs(5598) <= a or b;
    layer2_outputs(5599) <= b;
    layer2_outputs(5600) <= not a;
    layer2_outputs(5601) <= a xor b;
    layer2_outputs(5602) <= not (a or b);
    layer2_outputs(5603) <= not (a and b);
    layer2_outputs(5604) <= a or b;
    layer2_outputs(5605) <= b;
    layer2_outputs(5606) <= b and not a;
    layer2_outputs(5607) <= a;
    layer2_outputs(5608) <= not b or a;
    layer2_outputs(5609) <= a and not b;
    layer2_outputs(5610) <= not (a xor b);
    layer2_outputs(5611) <= a;
    layer2_outputs(5612) <= not a;
    layer2_outputs(5613) <= not a;
    layer2_outputs(5614) <= not (a or b);
    layer2_outputs(5615) <= b;
    layer2_outputs(5616) <= not b;
    layer2_outputs(5617) <= not b;
    layer2_outputs(5618) <= a;
    layer2_outputs(5619) <= not a or b;
    layer2_outputs(5620) <= b and not a;
    layer2_outputs(5621) <= not b;
    layer2_outputs(5622) <= a and not b;
    layer2_outputs(5623) <= not a;
    layer2_outputs(5624) <= not (a and b);
    layer2_outputs(5625) <= a and not b;
    layer2_outputs(5626) <= not (a and b);
    layer2_outputs(5627) <= b;
    layer2_outputs(5628) <= b;
    layer2_outputs(5629) <= not b;
    layer2_outputs(5630) <= not (a or b);
    layer2_outputs(5631) <= not (a xor b);
    layer2_outputs(5632) <= not b;
    layer2_outputs(5633) <= not a;
    layer2_outputs(5634) <= a;
    layer2_outputs(5635) <= 1'b1;
    layer2_outputs(5636) <= not a;
    layer2_outputs(5637) <= b;
    layer2_outputs(5638) <= b;
    layer2_outputs(5639) <= a and b;
    layer2_outputs(5640) <= not (a or b);
    layer2_outputs(5641) <= not a or b;
    layer2_outputs(5642) <= a;
    layer2_outputs(5643) <= not (a or b);
    layer2_outputs(5644) <= not (a or b);
    layer2_outputs(5645) <= a xor b;
    layer2_outputs(5646) <= b;
    layer2_outputs(5647) <= not b;
    layer2_outputs(5648) <= not b;
    layer2_outputs(5649) <= a xor b;
    layer2_outputs(5650) <= a and b;
    layer2_outputs(5651) <= b;
    layer2_outputs(5652) <= not (a xor b);
    layer2_outputs(5653) <= not b or a;
    layer2_outputs(5654) <= a or b;
    layer2_outputs(5655) <= not a;
    layer2_outputs(5656) <= a;
    layer2_outputs(5657) <= not (a xor b);
    layer2_outputs(5658) <= not a;
    layer2_outputs(5659) <= b;
    layer2_outputs(5660) <= a;
    layer2_outputs(5661) <= not (a and b);
    layer2_outputs(5662) <= not b;
    layer2_outputs(5663) <= a or b;
    layer2_outputs(5664) <= b;
    layer2_outputs(5665) <= a;
    layer2_outputs(5666) <= a and not b;
    layer2_outputs(5667) <= b;
    layer2_outputs(5668) <= not b or a;
    layer2_outputs(5669) <= not b;
    layer2_outputs(5670) <= a and not b;
    layer2_outputs(5671) <= not a;
    layer2_outputs(5672) <= a;
    layer2_outputs(5673) <= not a;
    layer2_outputs(5674) <= b and not a;
    layer2_outputs(5675) <= not a;
    layer2_outputs(5676) <= a and not b;
    layer2_outputs(5677) <= not a or b;
    layer2_outputs(5678) <= not a;
    layer2_outputs(5679) <= a or b;
    layer2_outputs(5680) <= not b;
    layer2_outputs(5681) <= b;
    layer2_outputs(5682) <= a;
    layer2_outputs(5683) <= 1'b0;
    layer2_outputs(5684) <= not (a or b);
    layer2_outputs(5685) <= a;
    layer2_outputs(5686) <= not a;
    layer2_outputs(5687) <= not a or b;
    layer2_outputs(5688) <= not b;
    layer2_outputs(5689) <= b and not a;
    layer2_outputs(5690) <= b and not a;
    layer2_outputs(5691) <= not (a and b);
    layer2_outputs(5692) <= not a;
    layer2_outputs(5693) <= not (a xor b);
    layer2_outputs(5694) <= not b;
    layer2_outputs(5695) <= not (a and b);
    layer2_outputs(5696) <= a and not b;
    layer2_outputs(5697) <= a;
    layer2_outputs(5698) <= a xor b;
    layer2_outputs(5699) <= not a or b;
    layer2_outputs(5700) <= not a;
    layer2_outputs(5701) <= b and not a;
    layer2_outputs(5702) <= not a or b;
    layer2_outputs(5703) <= not a;
    layer2_outputs(5704) <= a xor b;
    layer2_outputs(5705) <= not a or b;
    layer2_outputs(5706) <= a and not b;
    layer2_outputs(5707) <= b;
    layer2_outputs(5708) <= a or b;
    layer2_outputs(5709) <= not b;
    layer2_outputs(5710) <= not (a or b);
    layer2_outputs(5711) <= not a;
    layer2_outputs(5712) <= not a or b;
    layer2_outputs(5713) <= a;
    layer2_outputs(5714) <= not (a and b);
    layer2_outputs(5715) <= not (a xor b);
    layer2_outputs(5716) <= a xor b;
    layer2_outputs(5717) <= a and b;
    layer2_outputs(5718) <= not b;
    layer2_outputs(5719) <= not (a xor b);
    layer2_outputs(5720) <= a and not b;
    layer2_outputs(5721) <= b and not a;
    layer2_outputs(5722) <= not a;
    layer2_outputs(5723) <= b;
    layer2_outputs(5724) <= a and not b;
    layer2_outputs(5725) <= a;
    layer2_outputs(5726) <= not (a xor b);
    layer2_outputs(5727) <= not b or a;
    layer2_outputs(5728) <= not (a and b);
    layer2_outputs(5729) <= not (a or b);
    layer2_outputs(5730) <= b and not a;
    layer2_outputs(5731) <= b and not a;
    layer2_outputs(5732) <= not (a xor b);
    layer2_outputs(5733) <= not (a and b);
    layer2_outputs(5734) <= a xor b;
    layer2_outputs(5735) <= b;
    layer2_outputs(5736) <= not b or a;
    layer2_outputs(5737) <= not b or a;
    layer2_outputs(5738) <= b and not a;
    layer2_outputs(5739) <= not (a and b);
    layer2_outputs(5740) <= a and not b;
    layer2_outputs(5741) <= not b;
    layer2_outputs(5742) <= a and b;
    layer2_outputs(5743) <= not a;
    layer2_outputs(5744) <= not (a and b);
    layer2_outputs(5745) <= not (a or b);
    layer2_outputs(5746) <= a and not b;
    layer2_outputs(5747) <= not a or b;
    layer2_outputs(5748) <= b;
    layer2_outputs(5749) <= b;
    layer2_outputs(5750) <= a;
    layer2_outputs(5751) <= a and b;
    layer2_outputs(5752) <= b;
    layer2_outputs(5753) <= a;
    layer2_outputs(5754) <= b;
    layer2_outputs(5755) <= a or b;
    layer2_outputs(5756) <= not a;
    layer2_outputs(5757) <= b;
    layer2_outputs(5758) <= not (a and b);
    layer2_outputs(5759) <= b and not a;
    layer2_outputs(5760) <= b;
    layer2_outputs(5761) <= not (a and b);
    layer2_outputs(5762) <= not b or a;
    layer2_outputs(5763) <= not (a xor b);
    layer2_outputs(5764) <= not b;
    layer2_outputs(5765) <= b and not a;
    layer2_outputs(5766) <= not (a xor b);
    layer2_outputs(5767) <= a and b;
    layer2_outputs(5768) <= not b;
    layer2_outputs(5769) <= a and b;
    layer2_outputs(5770) <= not (a or b);
    layer2_outputs(5771) <= b;
    layer2_outputs(5772) <= not (a xor b);
    layer2_outputs(5773) <= not a or b;
    layer2_outputs(5774) <= b;
    layer2_outputs(5775) <= not (a and b);
    layer2_outputs(5776) <= a xor b;
    layer2_outputs(5777) <= not (a xor b);
    layer2_outputs(5778) <= not a;
    layer2_outputs(5779) <= not a or b;
    layer2_outputs(5780) <= b;
    layer2_outputs(5781) <= not (a xor b);
    layer2_outputs(5782) <= a and b;
    layer2_outputs(5783) <= b and not a;
    layer2_outputs(5784) <= not b or a;
    layer2_outputs(5785) <= not (a xor b);
    layer2_outputs(5786) <= not (a or b);
    layer2_outputs(5787) <= a or b;
    layer2_outputs(5788) <= a or b;
    layer2_outputs(5789) <= not (a or b);
    layer2_outputs(5790) <= not a or b;
    layer2_outputs(5791) <= not a;
    layer2_outputs(5792) <= not b or a;
    layer2_outputs(5793) <= a;
    layer2_outputs(5794) <= a;
    layer2_outputs(5795) <= b;
    layer2_outputs(5796) <= not (a or b);
    layer2_outputs(5797) <= a and not b;
    layer2_outputs(5798) <= a xor b;
    layer2_outputs(5799) <= a xor b;
    layer2_outputs(5800) <= not a;
    layer2_outputs(5801) <= not (a xor b);
    layer2_outputs(5802) <= not b;
    layer2_outputs(5803) <= not a or b;
    layer2_outputs(5804) <= a or b;
    layer2_outputs(5805) <= b;
    layer2_outputs(5806) <= a xor b;
    layer2_outputs(5807) <= not (a and b);
    layer2_outputs(5808) <= not (a or b);
    layer2_outputs(5809) <= a;
    layer2_outputs(5810) <= not (a or b);
    layer2_outputs(5811) <= a and b;
    layer2_outputs(5812) <= a;
    layer2_outputs(5813) <= not (a and b);
    layer2_outputs(5814) <= not (a and b);
    layer2_outputs(5815) <= not b;
    layer2_outputs(5816) <= a;
    layer2_outputs(5817) <= not b or a;
    layer2_outputs(5818) <= not b or a;
    layer2_outputs(5819) <= a and not b;
    layer2_outputs(5820) <= a;
    layer2_outputs(5821) <= b;
    layer2_outputs(5822) <= 1'b0;
    layer2_outputs(5823) <= not b;
    layer2_outputs(5824) <= not a;
    layer2_outputs(5825) <= not (a and b);
    layer2_outputs(5826) <= b;
    layer2_outputs(5827) <= not (a xor b);
    layer2_outputs(5828) <= not a or b;
    layer2_outputs(5829) <= a;
    layer2_outputs(5830) <= not b;
    layer2_outputs(5831) <= not (a or b);
    layer2_outputs(5832) <= not a;
    layer2_outputs(5833) <= not a or b;
    layer2_outputs(5834) <= a xor b;
    layer2_outputs(5835) <= a;
    layer2_outputs(5836) <= a or b;
    layer2_outputs(5837) <= b;
    layer2_outputs(5838) <= a and b;
    layer2_outputs(5839) <= b and not a;
    layer2_outputs(5840) <= not b;
    layer2_outputs(5841) <= not b;
    layer2_outputs(5842) <= a and not b;
    layer2_outputs(5843) <= not a;
    layer2_outputs(5844) <= not (a or b);
    layer2_outputs(5845) <= b;
    layer2_outputs(5846) <= b;
    layer2_outputs(5847) <= b;
    layer2_outputs(5848) <= not b or a;
    layer2_outputs(5849) <= a;
    layer2_outputs(5850) <= a or b;
    layer2_outputs(5851) <= not (a and b);
    layer2_outputs(5852) <= not b or a;
    layer2_outputs(5853) <= a xor b;
    layer2_outputs(5854) <= not (a or b);
    layer2_outputs(5855) <= a and not b;
    layer2_outputs(5856) <= a and not b;
    layer2_outputs(5857) <= not b;
    layer2_outputs(5858) <= a and b;
    layer2_outputs(5859) <= a xor b;
    layer2_outputs(5860) <= a or b;
    layer2_outputs(5861) <= not a;
    layer2_outputs(5862) <= a xor b;
    layer2_outputs(5863) <= a;
    layer2_outputs(5864) <= a;
    layer2_outputs(5865) <= a;
    layer2_outputs(5866) <= not b;
    layer2_outputs(5867) <= not (a and b);
    layer2_outputs(5868) <= a xor b;
    layer2_outputs(5869) <= a or b;
    layer2_outputs(5870) <= not a;
    layer2_outputs(5871) <= not b or a;
    layer2_outputs(5872) <= a xor b;
    layer2_outputs(5873) <= not b or a;
    layer2_outputs(5874) <= not a;
    layer2_outputs(5875) <= not a or b;
    layer2_outputs(5876) <= a and b;
    layer2_outputs(5877) <= not (a and b);
    layer2_outputs(5878) <= b and not a;
    layer2_outputs(5879) <= a xor b;
    layer2_outputs(5880) <= a and b;
    layer2_outputs(5881) <= a;
    layer2_outputs(5882) <= a xor b;
    layer2_outputs(5883) <= b;
    layer2_outputs(5884) <= a or b;
    layer2_outputs(5885) <= b;
    layer2_outputs(5886) <= a;
    layer2_outputs(5887) <= b;
    layer2_outputs(5888) <= not (a xor b);
    layer2_outputs(5889) <= not b or a;
    layer2_outputs(5890) <= not b;
    layer2_outputs(5891) <= not a;
    layer2_outputs(5892) <= b and not a;
    layer2_outputs(5893) <= 1'b0;
    layer2_outputs(5894) <= not b;
    layer2_outputs(5895) <= not (a or b);
    layer2_outputs(5896) <= a;
    layer2_outputs(5897) <= a;
    layer2_outputs(5898) <= a and not b;
    layer2_outputs(5899) <= a;
    layer2_outputs(5900) <= a;
    layer2_outputs(5901) <= b and not a;
    layer2_outputs(5902) <= b and not a;
    layer2_outputs(5903) <= a xor b;
    layer2_outputs(5904) <= b and not a;
    layer2_outputs(5905) <= a and b;
    layer2_outputs(5906) <= not a;
    layer2_outputs(5907) <= a or b;
    layer2_outputs(5908) <= a;
    layer2_outputs(5909) <= not (a or b);
    layer2_outputs(5910) <= a or b;
    layer2_outputs(5911) <= a and b;
    layer2_outputs(5912) <= not b or a;
    layer2_outputs(5913) <= not a;
    layer2_outputs(5914) <= not a;
    layer2_outputs(5915) <= not a;
    layer2_outputs(5916) <= b;
    layer2_outputs(5917) <= a;
    layer2_outputs(5918) <= not (a or b);
    layer2_outputs(5919) <= not b;
    layer2_outputs(5920) <= not (a and b);
    layer2_outputs(5921) <= not a;
    layer2_outputs(5922) <= a and b;
    layer2_outputs(5923) <= a;
    layer2_outputs(5924) <= a or b;
    layer2_outputs(5925) <= a and not b;
    layer2_outputs(5926) <= a or b;
    layer2_outputs(5927) <= b;
    layer2_outputs(5928) <= not (a xor b);
    layer2_outputs(5929) <= not (a xor b);
    layer2_outputs(5930) <= not a or b;
    layer2_outputs(5931) <= a xor b;
    layer2_outputs(5932) <= not b or a;
    layer2_outputs(5933) <= a xor b;
    layer2_outputs(5934) <= not b or a;
    layer2_outputs(5935) <= not (a and b);
    layer2_outputs(5936) <= not a;
    layer2_outputs(5937) <= a and b;
    layer2_outputs(5938) <= a and not b;
    layer2_outputs(5939) <= not (a and b);
    layer2_outputs(5940) <= not a;
    layer2_outputs(5941) <= a xor b;
    layer2_outputs(5942) <= not b;
    layer2_outputs(5943) <= not b;
    layer2_outputs(5944) <= not a;
    layer2_outputs(5945) <= a and b;
    layer2_outputs(5946) <= a and not b;
    layer2_outputs(5947) <= b;
    layer2_outputs(5948) <= not b or a;
    layer2_outputs(5949) <= not a or b;
    layer2_outputs(5950) <= not (a xor b);
    layer2_outputs(5951) <= not b;
    layer2_outputs(5952) <= a xor b;
    layer2_outputs(5953) <= a or b;
    layer2_outputs(5954) <= not b or a;
    layer2_outputs(5955) <= not a;
    layer2_outputs(5956) <= not (a and b);
    layer2_outputs(5957) <= b and not a;
    layer2_outputs(5958) <= not a or b;
    layer2_outputs(5959) <= not a;
    layer2_outputs(5960) <= not (a xor b);
    layer2_outputs(5961) <= a;
    layer2_outputs(5962) <= not a;
    layer2_outputs(5963) <= b and not a;
    layer2_outputs(5964) <= not b or a;
    layer2_outputs(5965) <= a xor b;
    layer2_outputs(5966) <= not a;
    layer2_outputs(5967) <= not a;
    layer2_outputs(5968) <= not b;
    layer2_outputs(5969) <= not b or a;
    layer2_outputs(5970) <= b;
    layer2_outputs(5971) <= 1'b1;
    layer2_outputs(5972) <= b;
    layer2_outputs(5973) <= not (a xor b);
    layer2_outputs(5974) <= b and not a;
    layer2_outputs(5975) <= not b;
    layer2_outputs(5976) <= a and not b;
    layer2_outputs(5977) <= not (a and b);
    layer2_outputs(5978) <= not b or a;
    layer2_outputs(5979) <= a xor b;
    layer2_outputs(5980) <= not a;
    layer2_outputs(5981) <= not b;
    layer2_outputs(5982) <= not a or b;
    layer2_outputs(5983) <= b and not a;
    layer2_outputs(5984) <= not a;
    layer2_outputs(5985) <= a or b;
    layer2_outputs(5986) <= a xor b;
    layer2_outputs(5987) <= a;
    layer2_outputs(5988) <= not a;
    layer2_outputs(5989) <= not (a and b);
    layer2_outputs(5990) <= a xor b;
    layer2_outputs(5991) <= not (a and b);
    layer2_outputs(5992) <= not b;
    layer2_outputs(5993) <= not a or b;
    layer2_outputs(5994) <= not b or a;
    layer2_outputs(5995) <= not (a and b);
    layer2_outputs(5996) <= b and not a;
    layer2_outputs(5997) <= a;
    layer2_outputs(5998) <= not a;
    layer2_outputs(5999) <= not a or b;
    layer2_outputs(6000) <= b;
    layer2_outputs(6001) <= not a or b;
    layer2_outputs(6002) <= not (a and b);
    layer2_outputs(6003) <= not a;
    layer2_outputs(6004) <= a and b;
    layer2_outputs(6005) <= a and b;
    layer2_outputs(6006) <= a and not b;
    layer2_outputs(6007) <= a xor b;
    layer2_outputs(6008) <= not (a xor b);
    layer2_outputs(6009) <= a xor b;
    layer2_outputs(6010) <= a xor b;
    layer2_outputs(6011) <= not b;
    layer2_outputs(6012) <= not (a and b);
    layer2_outputs(6013) <= not a;
    layer2_outputs(6014) <= not (a and b);
    layer2_outputs(6015) <= not b;
    layer2_outputs(6016) <= a and b;
    layer2_outputs(6017) <= not (a or b);
    layer2_outputs(6018) <= not a or b;
    layer2_outputs(6019) <= b;
    layer2_outputs(6020) <= a xor b;
    layer2_outputs(6021) <= b;
    layer2_outputs(6022) <= b and not a;
    layer2_outputs(6023) <= a xor b;
    layer2_outputs(6024) <= a and not b;
    layer2_outputs(6025) <= not a;
    layer2_outputs(6026) <= not a;
    layer2_outputs(6027) <= a and b;
    layer2_outputs(6028) <= a and not b;
    layer2_outputs(6029) <= a or b;
    layer2_outputs(6030) <= b and not a;
    layer2_outputs(6031) <= not b;
    layer2_outputs(6032) <= not (a or b);
    layer2_outputs(6033) <= b and not a;
    layer2_outputs(6034) <= not b or a;
    layer2_outputs(6035) <= a and not b;
    layer2_outputs(6036) <= not a;
    layer2_outputs(6037) <= b;
    layer2_outputs(6038) <= not (a xor b);
    layer2_outputs(6039) <= not b;
    layer2_outputs(6040) <= b;
    layer2_outputs(6041) <= a and not b;
    layer2_outputs(6042) <= not a;
    layer2_outputs(6043) <= a;
    layer2_outputs(6044) <= b;
    layer2_outputs(6045) <= b;
    layer2_outputs(6046) <= not a or b;
    layer2_outputs(6047) <= not a;
    layer2_outputs(6048) <= not (a xor b);
    layer2_outputs(6049) <= b;
    layer2_outputs(6050) <= a or b;
    layer2_outputs(6051) <= not b or a;
    layer2_outputs(6052) <= not a or b;
    layer2_outputs(6053) <= not a;
    layer2_outputs(6054) <= b and not a;
    layer2_outputs(6055) <= not a or b;
    layer2_outputs(6056) <= not a;
    layer2_outputs(6057) <= b;
    layer2_outputs(6058) <= not a;
    layer2_outputs(6059) <= not b;
    layer2_outputs(6060) <= b and not a;
    layer2_outputs(6061) <= not (a and b);
    layer2_outputs(6062) <= a;
    layer2_outputs(6063) <= not a;
    layer2_outputs(6064) <= a xor b;
    layer2_outputs(6065) <= b;
    layer2_outputs(6066) <= a and not b;
    layer2_outputs(6067) <= a and not b;
    layer2_outputs(6068) <= not b;
    layer2_outputs(6069) <= not a;
    layer2_outputs(6070) <= a and not b;
    layer2_outputs(6071) <= not a or b;
    layer2_outputs(6072) <= not b;
    layer2_outputs(6073) <= a or b;
    layer2_outputs(6074) <= b;
    layer2_outputs(6075) <= not a or b;
    layer2_outputs(6076) <= b;
    layer2_outputs(6077) <= a or b;
    layer2_outputs(6078) <= a and b;
    layer2_outputs(6079) <= not (a xor b);
    layer2_outputs(6080) <= not (a xor b);
    layer2_outputs(6081) <= b;
    layer2_outputs(6082) <= not a;
    layer2_outputs(6083) <= not (a or b);
    layer2_outputs(6084) <= not a or b;
    layer2_outputs(6085) <= not (a and b);
    layer2_outputs(6086) <= b and not a;
    layer2_outputs(6087) <= a and b;
    layer2_outputs(6088) <= not a;
    layer2_outputs(6089) <= a or b;
    layer2_outputs(6090) <= a;
    layer2_outputs(6091) <= not a;
    layer2_outputs(6092) <= not (a xor b);
    layer2_outputs(6093) <= not a;
    layer2_outputs(6094) <= not (a xor b);
    layer2_outputs(6095) <= not b;
    layer2_outputs(6096) <= not b;
    layer2_outputs(6097) <= a;
    layer2_outputs(6098) <= not (a xor b);
    layer2_outputs(6099) <= not a;
    layer2_outputs(6100) <= a;
    layer2_outputs(6101) <= not a;
    layer2_outputs(6102) <= a xor b;
    layer2_outputs(6103) <= a and b;
    layer2_outputs(6104) <= not (a and b);
    layer2_outputs(6105) <= not a;
    layer2_outputs(6106) <= a and b;
    layer2_outputs(6107) <= not b;
    layer2_outputs(6108) <= not (a and b);
    layer2_outputs(6109) <= not (a xor b);
    layer2_outputs(6110) <= a and not b;
    layer2_outputs(6111) <= not a or b;
    layer2_outputs(6112) <= a;
    layer2_outputs(6113) <= not b;
    layer2_outputs(6114) <= b and not a;
    layer2_outputs(6115) <= not (a or b);
    layer2_outputs(6116) <= not a or b;
    layer2_outputs(6117) <= not b or a;
    layer2_outputs(6118) <= b;
    layer2_outputs(6119) <= a and not b;
    layer2_outputs(6120) <= b;
    layer2_outputs(6121) <= not a or b;
    layer2_outputs(6122) <= not a;
    layer2_outputs(6123) <= b;
    layer2_outputs(6124) <= b;
    layer2_outputs(6125) <= a or b;
    layer2_outputs(6126) <= b and not a;
    layer2_outputs(6127) <= not a or b;
    layer2_outputs(6128) <= not a or b;
    layer2_outputs(6129) <= a or b;
    layer2_outputs(6130) <= b;
    layer2_outputs(6131) <= a xor b;
    layer2_outputs(6132) <= not a;
    layer2_outputs(6133) <= b and not a;
    layer2_outputs(6134) <= not (a xor b);
    layer2_outputs(6135) <= not a;
    layer2_outputs(6136) <= not (a and b);
    layer2_outputs(6137) <= a or b;
    layer2_outputs(6138) <= a xor b;
    layer2_outputs(6139) <= a;
    layer2_outputs(6140) <= a or b;
    layer2_outputs(6141) <= a and not b;
    layer2_outputs(6142) <= 1'b1;
    layer2_outputs(6143) <= not (a and b);
    layer2_outputs(6144) <= not b or a;
    layer2_outputs(6145) <= not (a xor b);
    layer2_outputs(6146) <= not b or a;
    layer2_outputs(6147) <= b and not a;
    layer2_outputs(6148) <= a;
    layer2_outputs(6149) <= not a or b;
    layer2_outputs(6150) <= not b or a;
    layer2_outputs(6151) <= not a;
    layer2_outputs(6152) <= not a;
    layer2_outputs(6153) <= not (a and b);
    layer2_outputs(6154) <= not a or b;
    layer2_outputs(6155) <= not b or a;
    layer2_outputs(6156) <= not b;
    layer2_outputs(6157) <= 1'b1;
    layer2_outputs(6158) <= not (a or b);
    layer2_outputs(6159) <= a and b;
    layer2_outputs(6160) <= a;
    layer2_outputs(6161) <= not a;
    layer2_outputs(6162) <= not b;
    layer2_outputs(6163) <= not b;
    layer2_outputs(6164) <= a or b;
    layer2_outputs(6165) <= a;
    layer2_outputs(6166) <= not (a xor b);
    layer2_outputs(6167) <= not (a or b);
    layer2_outputs(6168) <= not (a xor b);
    layer2_outputs(6169) <= b;
    layer2_outputs(6170) <= a and b;
    layer2_outputs(6171) <= a and not b;
    layer2_outputs(6172) <= not (a and b);
    layer2_outputs(6173) <= a and b;
    layer2_outputs(6174) <= not (a xor b);
    layer2_outputs(6175) <= not a or b;
    layer2_outputs(6176) <= a;
    layer2_outputs(6177) <= b;
    layer2_outputs(6178) <= a and b;
    layer2_outputs(6179) <= not (a or b);
    layer2_outputs(6180) <= not a;
    layer2_outputs(6181) <= 1'b1;
    layer2_outputs(6182) <= not a;
    layer2_outputs(6183) <= a;
    layer2_outputs(6184) <= not b or a;
    layer2_outputs(6185) <= not a or b;
    layer2_outputs(6186) <= not (a or b);
    layer2_outputs(6187) <= not b;
    layer2_outputs(6188) <= a xor b;
    layer2_outputs(6189) <= a and b;
    layer2_outputs(6190) <= a and b;
    layer2_outputs(6191) <= not b;
    layer2_outputs(6192) <= not a;
    layer2_outputs(6193) <= a or b;
    layer2_outputs(6194) <= a and not b;
    layer2_outputs(6195) <= not (a and b);
    layer2_outputs(6196) <= not (a or b);
    layer2_outputs(6197) <= not b or a;
    layer2_outputs(6198) <= a;
    layer2_outputs(6199) <= not (a and b);
    layer2_outputs(6200) <= a;
    layer2_outputs(6201) <= not a;
    layer2_outputs(6202) <= a;
    layer2_outputs(6203) <= a and b;
    layer2_outputs(6204) <= a xor b;
    layer2_outputs(6205) <= not b;
    layer2_outputs(6206) <= not (a xor b);
    layer2_outputs(6207) <= not a;
    layer2_outputs(6208) <= not a or b;
    layer2_outputs(6209) <= not a or b;
    layer2_outputs(6210) <= not b;
    layer2_outputs(6211) <= not (a or b);
    layer2_outputs(6212) <= not b or a;
    layer2_outputs(6213) <= b;
    layer2_outputs(6214) <= a xor b;
    layer2_outputs(6215) <= a and not b;
    layer2_outputs(6216) <= not (a and b);
    layer2_outputs(6217) <= a;
    layer2_outputs(6218) <= a and b;
    layer2_outputs(6219) <= not (a and b);
    layer2_outputs(6220) <= b and not a;
    layer2_outputs(6221) <= a or b;
    layer2_outputs(6222) <= a;
    layer2_outputs(6223) <= b;
    layer2_outputs(6224) <= not (a xor b);
    layer2_outputs(6225) <= not (a and b);
    layer2_outputs(6226) <= not b;
    layer2_outputs(6227) <= not (a xor b);
    layer2_outputs(6228) <= not b;
    layer2_outputs(6229) <= a;
    layer2_outputs(6230) <= a or b;
    layer2_outputs(6231) <= not (a xor b);
    layer2_outputs(6232) <= not (a xor b);
    layer2_outputs(6233) <= a;
    layer2_outputs(6234) <= not (a xor b);
    layer2_outputs(6235) <= b and not a;
    layer2_outputs(6236) <= b and not a;
    layer2_outputs(6237) <= not (a or b);
    layer2_outputs(6238) <= not b;
    layer2_outputs(6239) <= not (a or b);
    layer2_outputs(6240) <= not b or a;
    layer2_outputs(6241) <= a and b;
    layer2_outputs(6242) <= a;
    layer2_outputs(6243) <= a and not b;
    layer2_outputs(6244) <= a or b;
    layer2_outputs(6245) <= not (a or b);
    layer2_outputs(6246) <= not b;
    layer2_outputs(6247) <= a or b;
    layer2_outputs(6248) <= not (a and b);
    layer2_outputs(6249) <= not b;
    layer2_outputs(6250) <= a xor b;
    layer2_outputs(6251) <= a xor b;
    layer2_outputs(6252) <= not (a or b);
    layer2_outputs(6253) <= a;
    layer2_outputs(6254) <= not b;
    layer2_outputs(6255) <= not (a or b);
    layer2_outputs(6256) <= not b;
    layer2_outputs(6257) <= not (a or b);
    layer2_outputs(6258) <= a and b;
    layer2_outputs(6259) <= not b or a;
    layer2_outputs(6260) <= not (a xor b);
    layer2_outputs(6261) <= a and b;
    layer2_outputs(6262) <= a xor b;
    layer2_outputs(6263) <= not b or a;
    layer2_outputs(6264) <= b and not a;
    layer2_outputs(6265) <= not b;
    layer2_outputs(6266) <= not (a or b);
    layer2_outputs(6267) <= not (a and b);
    layer2_outputs(6268) <= not a;
    layer2_outputs(6269) <= not (a xor b);
    layer2_outputs(6270) <= b;
    layer2_outputs(6271) <= not (a and b);
    layer2_outputs(6272) <= a xor b;
    layer2_outputs(6273) <= a;
    layer2_outputs(6274) <= not b or a;
    layer2_outputs(6275) <= not (a or b);
    layer2_outputs(6276) <= not (a xor b);
    layer2_outputs(6277) <= not a or b;
    layer2_outputs(6278) <= a;
    layer2_outputs(6279) <= not b;
    layer2_outputs(6280) <= not a;
    layer2_outputs(6281) <= not (a or b);
    layer2_outputs(6282) <= not (a and b);
    layer2_outputs(6283) <= b and not a;
    layer2_outputs(6284) <= not (a or b);
    layer2_outputs(6285) <= a;
    layer2_outputs(6286) <= not b or a;
    layer2_outputs(6287) <= not (a or b);
    layer2_outputs(6288) <= a;
    layer2_outputs(6289) <= a xor b;
    layer2_outputs(6290) <= not b;
    layer2_outputs(6291) <= a;
    layer2_outputs(6292) <= a or b;
    layer2_outputs(6293) <= b and not a;
    layer2_outputs(6294) <= b;
    layer2_outputs(6295) <= a;
    layer2_outputs(6296) <= not a or b;
    layer2_outputs(6297) <= not b;
    layer2_outputs(6298) <= not b or a;
    layer2_outputs(6299) <= a and not b;
    layer2_outputs(6300) <= a xor b;
    layer2_outputs(6301) <= not b or a;
    layer2_outputs(6302) <= not b;
    layer2_outputs(6303) <= not (a xor b);
    layer2_outputs(6304) <= a;
    layer2_outputs(6305) <= not (a or b);
    layer2_outputs(6306) <= not b;
    layer2_outputs(6307) <= not (a xor b);
    layer2_outputs(6308) <= not (a xor b);
    layer2_outputs(6309) <= b;
    layer2_outputs(6310) <= a xor b;
    layer2_outputs(6311) <= not (a xor b);
    layer2_outputs(6312) <= not (a or b);
    layer2_outputs(6313) <= not (a xor b);
    layer2_outputs(6314) <= 1'b1;
    layer2_outputs(6315) <= a xor b;
    layer2_outputs(6316) <= a xor b;
    layer2_outputs(6317) <= b;
    layer2_outputs(6318) <= not b or a;
    layer2_outputs(6319) <= not b;
    layer2_outputs(6320) <= a;
    layer2_outputs(6321) <= not b;
    layer2_outputs(6322) <= b and not a;
    layer2_outputs(6323) <= not (a xor b);
    layer2_outputs(6324) <= a or b;
    layer2_outputs(6325) <= not (a xor b);
    layer2_outputs(6326) <= a or b;
    layer2_outputs(6327) <= b;
    layer2_outputs(6328) <= not b or a;
    layer2_outputs(6329) <= a xor b;
    layer2_outputs(6330) <= not b;
    layer2_outputs(6331) <= not (a and b);
    layer2_outputs(6332) <= a and b;
    layer2_outputs(6333) <= b and not a;
    layer2_outputs(6334) <= not a;
    layer2_outputs(6335) <= a xor b;
    layer2_outputs(6336) <= not (a or b);
    layer2_outputs(6337) <= not b or a;
    layer2_outputs(6338) <= not b;
    layer2_outputs(6339) <= not a;
    layer2_outputs(6340) <= not b or a;
    layer2_outputs(6341) <= not (a or b);
    layer2_outputs(6342) <= not b;
    layer2_outputs(6343) <= a xor b;
    layer2_outputs(6344) <= not a;
    layer2_outputs(6345) <= not a;
    layer2_outputs(6346) <= not a or b;
    layer2_outputs(6347) <= not a;
    layer2_outputs(6348) <= b;
    layer2_outputs(6349) <= b and not a;
    layer2_outputs(6350) <= not a;
    layer2_outputs(6351) <= not b or a;
    layer2_outputs(6352) <= not (a xor b);
    layer2_outputs(6353) <= a;
    layer2_outputs(6354) <= not a or b;
    layer2_outputs(6355) <= not (a and b);
    layer2_outputs(6356) <= b and not a;
    layer2_outputs(6357) <= a;
    layer2_outputs(6358) <= not a;
    layer2_outputs(6359) <= a;
    layer2_outputs(6360) <= a xor b;
    layer2_outputs(6361) <= a and b;
    layer2_outputs(6362) <= b;
    layer2_outputs(6363) <= not b or a;
    layer2_outputs(6364) <= not b or a;
    layer2_outputs(6365) <= a xor b;
    layer2_outputs(6366) <= a xor b;
    layer2_outputs(6367) <= a or b;
    layer2_outputs(6368) <= not a or b;
    layer2_outputs(6369) <= not a;
    layer2_outputs(6370) <= a;
    layer2_outputs(6371) <= b;
    layer2_outputs(6372) <= not a or b;
    layer2_outputs(6373) <= not b;
    layer2_outputs(6374) <= b;
    layer2_outputs(6375) <= a;
    layer2_outputs(6376) <= not a;
    layer2_outputs(6377) <= not b or a;
    layer2_outputs(6378) <= not (a or b);
    layer2_outputs(6379) <= a and b;
    layer2_outputs(6380) <= a xor b;
    layer2_outputs(6381) <= not (a and b);
    layer2_outputs(6382) <= a xor b;
    layer2_outputs(6383) <= not b;
    layer2_outputs(6384) <= a and b;
    layer2_outputs(6385) <= b and not a;
    layer2_outputs(6386) <= not (a or b);
    layer2_outputs(6387) <= a xor b;
    layer2_outputs(6388) <= not a;
    layer2_outputs(6389) <= 1'b1;
    layer2_outputs(6390) <= not (a and b);
    layer2_outputs(6391) <= not (a or b);
    layer2_outputs(6392) <= a;
    layer2_outputs(6393) <= a;
    layer2_outputs(6394) <= b and not a;
    layer2_outputs(6395) <= not (a or b);
    layer2_outputs(6396) <= a and not b;
    layer2_outputs(6397) <= not b or a;
    layer2_outputs(6398) <= a;
    layer2_outputs(6399) <= a and not b;
    layer2_outputs(6400) <= a and b;
    layer2_outputs(6401) <= not a or b;
    layer2_outputs(6402) <= not (a xor b);
    layer2_outputs(6403) <= not b;
    layer2_outputs(6404) <= b;
    layer2_outputs(6405) <= not a;
    layer2_outputs(6406) <= a or b;
    layer2_outputs(6407) <= a xor b;
    layer2_outputs(6408) <= not b;
    layer2_outputs(6409) <= b and not a;
    layer2_outputs(6410) <= b;
    layer2_outputs(6411) <= a or b;
    layer2_outputs(6412) <= a and not b;
    layer2_outputs(6413) <= not a;
    layer2_outputs(6414) <= not a;
    layer2_outputs(6415) <= b;
    layer2_outputs(6416) <= not a or b;
    layer2_outputs(6417) <= a;
    layer2_outputs(6418) <= not a;
    layer2_outputs(6419) <= b;
    layer2_outputs(6420) <= not (a xor b);
    layer2_outputs(6421) <= b;
    layer2_outputs(6422) <= a and not b;
    layer2_outputs(6423) <= a or b;
    layer2_outputs(6424) <= not b;
    layer2_outputs(6425) <= not b;
    layer2_outputs(6426) <= not (a xor b);
    layer2_outputs(6427) <= not a or b;
    layer2_outputs(6428) <= a or b;
    layer2_outputs(6429) <= a and not b;
    layer2_outputs(6430) <= not (a or b);
    layer2_outputs(6431) <= a and b;
    layer2_outputs(6432) <= not b;
    layer2_outputs(6433) <= not (a and b);
    layer2_outputs(6434) <= a or b;
    layer2_outputs(6435) <= a xor b;
    layer2_outputs(6436) <= not (a xor b);
    layer2_outputs(6437) <= b;
    layer2_outputs(6438) <= b;
    layer2_outputs(6439) <= not a;
    layer2_outputs(6440) <= a;
    layer2_outputs(6441) <= not a;
    layer2_outputs(6442) <= a;
    layer2_outputs(6443) <= a xor b;
    layer2_outputs(6444) <= not a;
    layer2_outputs(6445) <= a xor b;
    layer2_outputs(6446) <= a xor b;
    layer2_outputs(6447) <= not a;
    layer2_outputs(6448) <= a;
    layer2_outputs(6449) <= not a;
    layer2_outputs(6450) <= a or b;
    layer2_outputs(6451) <= not (a or b);
    layer2_outputs(6452) <= a and not b;
    layer2_outputs(6453) <= a or b;
    layer2_outputs(6454) <= a and not b;
    layer2_outputs(6455) <= not a;
    layer2_outputs(6456) <= not a or b;
    layer2_outputs(6457) <= not a;
    layer2_outputs(6458) <= not a;
    layer2_outputs(6459) <= not b;
    layer2_outputs(6460) <= not b;
    layer2_outputs(6461) <= a and b;
    layer2_outputs(6462) <= b;
    layer2_outputs(6463) <= not a;
    layer2_outputs(6464) <= a xor b;
    layer2_outputs(6465) <= a and b;
    layer2_outputs(6466) <= not a;
    layer2_outputs(6467) <= not b or a;
    layer2_outputs(6468) <= b;
    layer2_outputs(6469) <= not b;
    layer2_outputs(6470) <= a;
    layer2_outputs(6471) <= a and not b;
    layer2_outputs(6472) <= not (a and b);
    layer2_outputs(6473) <= not (a and b);
    layer2_outputs(6474) <= not a;
    layer2_outputs(6475) <= not a;
    layer2_outputs(6476) <= not a;
    layer2_outputs(6477) <= not (a and b);
    layer2_outputs(6478) <= not b;
    layer2_outputs(6479) <= a and b;
    layer2_outputs(6480) <= a xor b;
    layer2_outputs(6481) <= not a or b;
    layer2_outputs(6482) <= 1'b0;
    layer2_outputs(6483) <= not b or a;
    layer2_outputs(6484) <= a;
    layer2_outputs(6485) <= b and not a;
    layer2_outputs(6486) <= 1'b0;
    layer2_outputs(6487) <= b and not a;
    layer2_outputs(6488) <= a;
    layer2_outputs(6489) <= b and not a;
    layer2_outputs(6490) <= not a;
    layer2_outputs(6491) <= not a;
    layer2_outputs(6492) <= a and not b;
    layer2_outputs(6493) <= a xor b;
    layer2_outputs(6494) <= not b;
    layer2_outputs(6495) <= b;
    layer2_outputs(6496) <= not a or b;
    layer2_outputs(6497) <= a and not b;
    layer2_outputs(6498) <= not b;
    layer2_outputs(6499) <= not (a or b);
    layer2_outputs(6500) <= a xor b;
    layer2_outputs(6501) <= not a;
    layer2_outputs(6502) <= not (a and b);
    layer2_outputs(6503) <= a and b;
    layer2_outputs(6504) <= not b;
    layer2_outputs(6505) <= a;
    layer2_outputs(6506) <= not (a xor b);
    layer2_outputs(6507) <= not (a xor b);
    layer2_outputs(6508) <= not a;
    layer2_outputs(6509) <= b and not a;
    layer2_outputs(6510) <= not b;
    layer2_outputs(6511) <= a and b;
    layer2_outputs(6512) <= b;
    layer2_outputs(6513) <= not (a and b);
    layer2_outputs(6514) <= b;
    layer2_outputs(6515) <= a or b;
    layer2_outputs(6516) <= not (a or b);
    layer2_outputs(6517) <= not (a and b);
    layer2_outputs(6518) <= b and not a;
    layer2_outputs(6519) <= b;
    layer2_outputs(6520) <= a xor b;
    layer2_outputs(6521) <= not b;
    layer2_outputs(6522) <= a or b;
    layer2_outputs(6523) <= a and b;
    layer2_outputs(6524) <= not a or b;
    layer2_outputs(6525) <= not (a xor b);
    layer2_outputs(6526) <= not b;
    layer2_outputs(6527) <= not a or b;
    layer2_outputs(6528) <= b and not a;
    layer2_outputs(6529) <= not (a xor b);
    layer2_outputs(6530) <= not (a or b);
    layer2_outputs(6531) <= not (a or b);
    layer2_outputs(6532) <= a xor b;
    layer2_outputs(6533) <= b and not a;
    layer2_outputs(6534) <= not a or b;
    layer2_outputs(6535) <= not (a or b);
    layer2_outputs(6536) <= b;
    layer2_outputs(6537) <= a and b;
    layer2_outputs(6538) <= not (a xor b);
    layer2_outputs(6539) <= 1'b1;
    layer2_outputs(6540) <= not b or a;
    layer2_outputs(6541) <= a and b;
    layer2_outputs(6542) <= not a;
    layer2_outputs(6543) <= not a;
    layer2_outputs(6544) <= a;
    layer2_outputs(6545) <= not (a xor b);
    layer2_outputs(6546) <= not (a or b);
    layer2_outputs(6547) <= not (a and b);
    layer2_outputs(6548) <= a xor b;
    layer2_outputs(6549) <= not a or b;
    layer2_outputs(6550) <= a;
    layer2_outputs(6551) <= not a;
    layer2_outputs(6552) <= not (a xor b);
    layer2_outputs(6553) <= a;
    layer2_outputs(6554) <= not a;
    layer2_outputs(6555) <= b;
    layer2_outputs(6556) <= not (a or b);
    layer2_outputs(6557) <= not (a or b);
    layer2_outputs(6558) <= a and b;
    layer2_outputs(6559) <= a;
    layer2_outputs(6560) <= not (a or b);
    layer2_outputs(6561) <= not (a and b);
    layer2_outputs(6562) <= b and not a;
    layer2_outputs(6563) <= a and b;
    layer2_outputs(6564) <= b;
    layer2_outputs(6565) <= not b or a;
    layer2_outputs(6566) <= not (a and b);
    layer2_outputs(6567) <= not b;
    layer2_outputs(6568) <= a xor b;
    layer2_outputs(6569) <= not a;
    layer2_outputs(6570) <= not b or a;
    layer2_outputs(6571) <= not a;
    layer2_outputs(6572) <= a and not b;
    layer2_outputs(6573) <= a;
    layer2_outputs(6574) <= b;
    layer2_outputs(6575) <= not a;
    layer2_outputs(6576) <= a and b;
    layer2_outputs(6577) <= a and b;
    layer2_outputs(6578) <= not a;
    layer2_outputs(6579) <= not a;
    layer2_outputs(6580) <= not a or b;
    layer2_outputs(6581) <= b and not a;
    layer2_outputs(6582) <= a;
    layer2_outputs(6583) <= b;
    layer2_outputs(6584) <= b;
    layer2_outputs(6585) <= b;
    layer2_outputs(6586) <= b and not a;
    layer2_outputs(6587) <= a and not b;
    layer2_outputs(6588) <= b;
    layer2_outputs(6589) <= b;
    layer2_outputs(6590) <= not (a xor b);
    layer2_outputs(6591) <= not b;
    layer2_outputs(6592) <= b and not a;
    layer2_outputs(6593) <= a;
    layer2_outputs(6594) <= a and b;
    layer2_outputs(6595) <= not b or a;
    layer2_outputs(6596) <= b;
    layer2_outputs(6597) <= a xor b;
    layer2_outputs(6598) <= b and not a;
    layer2_outputs(6599) <= 1'b1;
    layer2_outputs(6600) <= not (a xor b);
    layer2_outputs(6601) <= b;
    layer2_outputs(6602) <= not (a and b);
    layer2_outputs(6603) <= b;
    layer2_outputs(6604) <= a;
    layer2_outputs(6605) <= b and not a;
    layer2_outputs(6606) <= not (a or b);
    layer2_outputs(6607) <= not b;
    layer2_outputs(6608) <= a;
    layer2_outputs(6609) <= not (a and b);
    layer2_outputs(6610) <= a;
    layer2_outputs(6611) <= b;
    layer2_outputs(6612) <= b and not a;
    layer2_outputs(6613) <= b;
    layer2_outputs(6614) <= not a or b;
    layer2_outputs(6615) <= not b;
    layer2_outputs(6616) <= a xor b;
    layer2_outputs(6617) <= not (a or b);
    layer2_outputs(6618) <= a and b;
    layer2_outputs(6619) <= b and not a;
    layer2_outputs(6620) <= a;
    layer2_outputs(6621) <= a xor b;
    layer2_outputs(6622) <= not a;
    layer2_outputs(6623) <= not b;
    layer2_outputs(6624) <= a or b;
    layer2_outputs(6625) <= not b;
    layer2_outputs(6626) <= a and not b;
    layer2_outputs(6627) <= not (a xor b);
    layer2_outputs(6628) <= not a;
    layer2_outputs(6629) <= a and b;
    layer2_outputs(6630) <= a or b;
    layer2_outputs(6631) <= not (a or b);
    layer2_outputs(6632) <= a xor b;
    layer2_outputs(6633) <= a or b;
    layer2_outputs(6634) <= a and not b;
    layer2_outputs(6635) <= b and not a;
    layer2_outputs(6636) <= b;
    layer2_outputs(6637) <= not (a and b);
    layer2_outputs(6638) <= a;
    layer2_outputs(6639) <= a xor b;
    layer2_outputs(6640) <= not (a xor b);
    layer2_outputs(6641) <= a and not b;
    layer2_outputs(6642) <= a;
    layer2_outputs(6643) <= a;
    layer2_outputs(6644) <= not a;
    layer2_outputs(6645) <= a or b;
    layer2_outputs(6646) <= not b;
    layer2_outputs(6647) <= a and not b;
    layer2_outputs(6648) <= a and b;
    layer2_outputs(6649) <= b and not a;
    layer2_outputs(6650) <= not a or b;
    layer2_outputs(6651) <= b;
    layer2_outputs(6652) <= b;
    layer2_outputs(6653) <= a xor b;
    layer2_outputs(6654) <= not b;
    layer2_outputs(6655) <= not (a and b);
    layer2_outputs(6656) <= not b;
    layer2_outputs(6657) <= not (a xor b);
    layer2_outputs(6658) <= b;
    layer2_outputs(6659) <= a xor b;
    layer2_outputs(6660) <= not a or b;
    layer2_outputs(6661) <= not b;
    layer2_outputs(6662) <= b and not a;
    layer2_outputs(6663) <= not a;
    layer2_outputs(6664) <= b and not a;
    layer2_outputs(6665) <= a and not b;
    layer2_outputs(6666) <= not a;
    layer2_outputs(6667) <= not b;
    layer2_outputs(6668) <= not a;
    layer2_outputs(6669) <= b and not a;
    layer2_outputs(6670) <= a or b;
    layer2_outputs(6671) <= b;
    layer2_outputs(6672) <= not b or a;
    layer2_outputs(6673) <= b and not a;
    layer2_outputs(6674) <= b;
    layer2_outputs(6675) <= not (a or b);
    layer2_outputs(6676) <= a xor b;
    layer2_outputs(6677) <= a and not b;
    layer2_outputs(6678) <= not a;
    layer2_outputs(6679) <= a;
    layer2_outputs(6680) <= b and not a;
    layer2_outputs(6681) <= not b or a;
    layer2_outputs(6682) <= a xor b;
    layer2_outputs(6683) <= not (a xor b);
    layer2_outputs(6684) <= a and not b;
    layer2_outputs(6685) <= a and b;
    layer2_outputs(6686) <= not b or a;
    layer2_outputs(6687) <= not a;
    layer2_outputs(6688) <= b;
    layer2_outputs(6689) <= not b;
    layer2_outputs(6690) <= not b or a;
    layer2_outputs(6691) <= a xor b;
    layer2_outputs(6692) <= not b;
    layer2_outputs(6693) <= not a;
    layer2_outputs(6694) <= 1'b0;
    layer2_outputs(6695) <= not (a xor b);
    layer2_outputs(6696) <= b;
    layer2_outputs(6697) <= not b;
    layer2_outputs(6698) <= b;
    layer2_outputs(6699) <= a;
    layer2_outputs(6700) <= a;
    layer2_outputs(6701) <= b and not a;
    layer2_outputs(6702) <= not a or b;
    layer2_outputs(6703) <= not a;
    layer2_outputs(6704) <= b and not a;
    layer2_outputs(6705) <= not (a or b);
    layer2_outputs(6706) <= a;
    layer2_outputs(6707) <= a and b;
    layer2_outputs(6708) <= not a;
    layer2_outputs(6709) <= b;
    layer2_outputs(6710) <= a and not b;
    layer2_outputs(6711) <= b;
    layer2_outputs(6712) <= a and b;
    layer2_outputs(6713) <= b and not a;
    layer2_outputs(6714) <= b;
    layer2_outputs(6715) <= a xor b;
    layer2_outputs(6716) <= a;
    layer2_outputs(6717) <= not (a and b);
    layer2_outputs(6718) <= a xor b;
    layer2_outputs(6719) <= b;
    layer2_outputs(6720) <= a and not b;
    layer2_outputs(6721) <= a or b;
    layer2_outputs(6722) <= not (a and b);
    layer2_outputs(6723) <= not (a or b);
    layer2_outputs(6724) <= not b;
    layer2_outputs(6725) <= not (a or b);
    layer2_outputs(6726) <= a or b;
    layer2_outputs(6727) <= not (a xor b);
    layer2_outputs(6728) <= b;
    layer2_outputs(6729) <= 1'b1;
    layer2_outputs(6730) <= a and b;
    layer2_outputs(6731) <= not (a and b);
    layer2_outputs(6732) <= a;
    layer2_outputs(6733) <= not a;
    layer2_outputs(6734) <= b;
    layer2_outputs(6735) <= not b or a;
    layer2_outputs(6736) <= a;
    layer2_outputs(6737) <= b and not a;
    layer2_outputs(6738) <= a and not b;
    layer2_outputs(6739) <= not a;
    layer2_outputs(6740) <= b and not a;
    layer2_outputs(6741) <= b;
    layer2_outputs(6742) <= not a;
    layer2_outputs(6743) <= not a or b;
    layer2_outputs(6744) <= a and b;
    layer2_outputs(6745) <= b;
    layer2_outputs(6746) <= a and b;
    layer2_outputs(6747) <= a xor b;
    layer2_outputs(6748) <= a xor b;
    layer2_outputs(6749) <= a xor b;
    layer2_outputs(6750) <= not (a or b);
    layer2_outputs(6751) <= a;
    layer2_outputs(6752) <= not b;
    layer2_outputs(6753) <= a;
    layer2_outputs(6754) <= not (a xor b);
    layer2_outputs(6755) <= a or b;
    layer2_outputs(6756) <= a xor b;
    layer2_outputs(6757) <= b and not a;
    layer2_outputs(6758) <= not (a and b);
    layer2_outputs(6759) <= not a;
    layer2_outputs(6760) <= not b;
    layer2_outputs(6761) <= not (a and b);
    layer2_outputs(6762) <= not b or a;
    layer2_outputs(6763) <= a or b;
    layer2_outputs(6764) <= a;
    layer2_outputs(6765) <= a;
    layer2_outputs(6766) <= a and b;
    layer2_outputs(6767) <= b;
    layer2_outputs(6768) <= not a;
    layer2_outputs(6769) <= a and not b;
    layer2_outputs(6770) <= not a;
    layer2_outputs(6771) <= not (a xor b);
    layer2_outputs(6772) <= not (a xor b);
    layer2_outputs(6773) <= not b;
    layer2_outputs(6774) <= not a;
    layer2_outputs(6775) <= not a;
    layer2_outputs(6776) <= a and b;
    layer2_outputs(6777) <= not a;
    layer2_outputs(6778) <= a xor b;
    layer2_outputs(6779) <= b and not a;
    layer2_outputs(6780) <= a xor b;
    layer2_outputs(6781) <= a or b;
    layer2_outputs(6782) <= b;
    layer2_outputs(6783) <= not (a and b);
    layer2_outputs(6784) <= a or b;
    layer2_outputs(6785) <= not (a and b);
    layer2_outputs(6786) <= a xor b;
    layer2_outputs(6787) <= a and b;
    layer2_outputs(6788) <= not (a and b);
    layer2_outputs(6789) <= b;
    layer2_outputs(6790) <= not a or b;
    layer2_outputs(6791) <= a xor b;
    layer2_outputs(6792) <= not (a xor b);
    layer2_outputs(6793) <= b and not a;
    layer2_outputs(6794) <= not (a or b);
    layer2_outputs(6795) <= not b or a;
    layer2_outputs(6796) <= not b or a;
    layer2_outputs(6797) <= a and not b;
    layer2_outputs(6798) <= not (a xor b);
    layer2_outputs(6799) <= not a;
    layer2_outputs(6800) <= not (a and b);
    layer2_outputs(6801) <= not b;
    layer2_outputs(6802) <= not (a xor b);
    layer2_outputs(6803) <= b;
    layer2_outputs(6804) <= not b or a;
    layer2_outputs(6805) <= a and b;
    layer2_outputs(6806) <= not b or a;
    layer2_outputs(6807) <= a and b;
    layer2_outputs(6808) <= a or b;
    layer2_outputs(6809) <= a or b;
    layer2_outputs(6810) <= a xor b;
    layer2_outputs(6811) <= b;
    layer2_outputs(6812) <= not b;
    layer2_outputs(6813) <= a or b;
    layer2_outputs(6814) <= a or b;
    layer2_outputs(6815) <= 1'b1;
    layer2_outputs(6816) <= a;
    layer2_outputs(6817) <= not a;
    layer2_outputs(6818) <= not b or a;
    layer2_outputs(6819) <= not b or a;
    layer2_outputs(6820) <= not b or a;
    layer2_outputs(6821) <= not (a xor b);
    layer2_outputs(6822) <= a and b;
    layer2_outputs(6823) <= a and not b;
    layer2_outputs(6824) <= not a or b;
    layer2_outputs(6825) <= not b;
    layer2_outputs(6826) <= not (a xor b);
    layer2_outputs(6827) <= b;
    layer2_outputs(6828) <= not b;
    layer2_outputs(6829) <= a xor b;
    layer2_outputs(6830) <= not a or b;
    layer2_outputs(6831) <= a;
    layer2_outputs(6832) <= not b;
    layer2_outputs(6833) <= a and b;
    layer2_outputs(6834) <= not (a or b);
    layer2_outputs(6835) <= a or b;
    layer2_outputs(6836) <= a;
    layer2_outputs(6837) <= not a or b;
    layer2_outputs(6838) <= not (a xor b);
    layer2_outputs(6839) <= not (a xor b);
    layer2_outputs(6840) <= a and b;
    layer2_outputs(6841) <= a;
    layer2_outputs(6842) <= not b;
    layer2_outputs(6843) <= not a;
    layer2_outputs(6844) <= a and b;
    layer2_outputs(6845) <= not b;
    layer2_outputs(6846) <= a;
    layer2_outputs(6847) <= a or b;
    layer2_outputs(6848) <= a;
    layer2_outputs(6849) <= not b;
    layer2_outputs(6850) <= not b or a;
    layer2_outputs(6851) <= a;
    layer2_outputs(6852) <= not (a xor b);
    layer2_outputs(6853) <= not (a and b);
    layer2_outputs(6854) <= a;
    layer2_outputs(6855) <= not a or b;
    layer2_outputs(6856) <= a;
    layer2_outputs(6857) <= b;
    layer2_outputs(6858) <= not (a or b);
    layer2_outputs(6859) <= not a;
    layer2_outputs(6860) <= 1'b1;
    layer2_outputs(6861) <= not b;
    layer2_outputs(6862) <= b and not a;
    layer2_outputs(6863) <= not b;
    layer2_outputs(6864) <= b and not a;
    layer2_outputs(6865) <= a xor b;
    layer2_outputs(6866) <= b and not a;
    layer2_outputs(6867) <= not b;
    layer2_outputs(6868) <= not b;
    layer2_outputs(6869) <= not b;
    layer2_outputs(6870) <= not (a and b);
    layer2_outputs(6871) <= not (a or b);
    layer2_outputs(6872) <= a xor b;
    layer2_outputs(6873) <= a xor b;
    layer2_outputs(6874) <= a or b;
    layer2_outputs(6875) <= a xor b;
    layer2_outputs(6876) <= not a;
    layer2_outputs(6877) <= b;
    layer2_outputs(6878) <= b;
    layer2_outputs(6879) <= not (a xor b);
    layer2_outputs(6880) <= not (a and b);
    layer2_outputs(6881) <= a xor b;
    layer2_outputs(6882) <= not (a or b);
    layer2_outputs(6883) <= not (a and b);
    layer2_outputs(6884) <= not (a and b);
    layer2_outputs(6885) <= not b or a;
    layer2_outputs(6886) <= not b;
    layer2_outputs(6887) <= not a or b;
    layer2_outputs(6888) <= not (a xor b);
    layer2_outputs(6889) <= 1'b0;
    layer2_outputs(6890) <= not a or b;
    layer2_outputs(6891) <= not b;
    layer2_outputs(6892) <= not (a and b);
    layer2_outputs(6893) <= not a;
    layer2_outputs(6894) <= not a or b;
    layer2_outputs(6895) <= b and not a;
    layer2_outputs(6896) <= b;
    layer2_outputs(6897) <= a;
    layer2_outputs(6898) <= not a or b;
    layer2_outputs(6899) <= not b;
    layer2_outputs(6900) <= a xor b;
    layer2_outputs(6901) <= a;
    layer2_outputs(6902) <= not a;
    layer2_outputs(6903) <= a and b;
    layer2_outputs(6904) <= not (a and b);
    layer2_outputs(6905) <= not (a xor b);
    layer2_outputs(6906) <= not a or b;
    layer2_outputs(6907) <= a or b;
    layer2_outputs(6908) <= a;
    layer2_outputs(6909) <= not b;
    layer2_outputs(6910) <= not (a and b);
    layer2_outputs(6911) <= not a or b;
    layer2_outputs(6912) <= a or b;
    layer2_outputs(6913) <= not (a or b);
    layer2_outputs(6914) <= a;
    layer2_outputs(6915) <= a and not b;
    layer2_outputs(6916) <= a;
    layer2_outputs(6917) <= not a;
    layer2_outputs(6918) <= a or b;
    layer2_outputs(6919) <= a xor b;
    layer2_outputs(6920) <= not a;
    layer2_outputs(6921) <= a xor b;
    layer2_outputs(6922) <= not (a or b);
    layer2_outputs(6923) <= not a;
    layer2_outputs(6924) <= not b or a;
    layer2_outputs(6925) <= a and b;
    layer2_outputs(6926) <= a;
    layer2_outputs(6927) <= a;
    layer2_outputs(6928) <= not (a xor b);
    layer2_outputs(6929) <= a or b;
    layer2_outputs(6930) <= a xor b;
    layer2_outputs(6931) <= not b;
    layer2_outputs(6932) <= a;
    layer2_outputs(6933) <= a and not b;
    layer2_outputs(6934) <= a and b;
    layer2_outputs(6935) <= not (a or b);
    layer2_outputs(6936) <= not (a xor b);
    layer2_outputs(6937) <= a xor b;
    layer2_outputs(6938) <= not a or b;
    layer2_outputs(6939) <= a or b;
    layer2_outputs(6940) <= not a or b;
    layer2_outputs(6941) <= not (a xor b);
    layer2_outputs(6942) <= a and b;
    layer2_outputs(6943) <= b;
    layer2_outputs(6944) <= a or b;
    layer2_outputs(6945) <= not b or a;
    layer2_outputs(6946) <= a;
    layer2_outputs(6947) <= not a;
    layer2_outputs(6948) <= b;
    layer2_outputs(6949) <= not (a or b);
    layer2_outputs(6950) <= a or b;
    layer2_outputs(6951) <= not b or a;
    layer2_outputs(6952) <= not (a and b);
    layer2_outputs(6953) <= not (a and b);
    layer2_outputs(6954) <= b;
    layer2_outputs(6955) <= not b;
    layer2_outputs(6956) <= not b or a;
    layer2_outputs(6957) <= b;
    layer2_outputs(6958) <= a;
    layer2_outputs(6959) <= a and b;
    layer2_outputs(6960) <= not b;
    layer2_outputs(6961) <= not a;
    layer2_outputs(6962) <= a or b;
    layer2_outputs(6963) <= not a or b;
    layer2_outputs(6964) <= not b;
    layer2_outputs(6965) <= not a or b;
    layer2_outputs(6966) <= a and b;
    layer2_outputs(6967) <= not b;
    layer2_outputs(6968) <= a;
    layer2_outputs(6969) <= not (a xor b);
    layer2_outputs(6970) <= a and not b;
    layer2_outputs(6971) <= not a;
    layer2_outputs(6972) <= not b or a;
    layer2_outputs(6973) <= not (a or b);
    layer2_outputs(6974) <= not (a or b);
    layer2_outputs(6975) <= not b;
    layer2_outputs(6976) <= not b or a;
    layer2_outputs(6977) <= not a;
    layer2_outputs(6978) <= not b;
    layer2_outputs(6979) <= not a;
    layer2_outputs(6980) <= a or b;
    layer2_outputs(6981) <= not b;
    layer2_outputs(6982) <= a xor b;
    layer2_outputs(6983) <= b;
    layer2_outputs(6984) <= a and not b;
    layer2_outputs(6985) <= a or b;
    layer2_outputs(6986) <= not (a or b);
    layer2_outputs(6987) <= not (a and b);
    layer2_outputs(6988) <= not a;
    layer2_outputs(6989) <= not b;
    layer2_outputs(6990) <= not b;
    layer2_outputs(6991) <= not (a xor b);
    layer2_outputs(6992) <= not (a and b);
    layer2_outputs(6993) <= not b;
    layer2_outputs(6994) <= not b or a;
    layer2_outputs(6995) <= not (a xor b);
    layer2_outputs(6996) <= a or b;
    layer2_outputs(6997) <= a xor b;
    layer2_outputs(6998) <= not (a and b);
    layer2_outputs(6999) <= not b or a;
    layer2_outputs(7000) <= 1'b0;
    layer2_outputs(7001) <= not b or a;
    layer2_outputs(7002) <= a and b;
    layer2_outputs(7003) <= a or b;
    layer2_outputs(7004) <= not a;
    layer2_outputs(7005) <= b;
    layer2_outputs(7006) <= not b;
    layer2_outputs(7007) <= a xor b;
    layer2_outputs(7008) <= a and not b;
    layer2_outputs(7009) <= b;
    layer2_outputs(7010) <= not (a or b);
    layer2_outputs(7011) <= a or b;
    layer2_outputs(7012) <= a and not b;
    layer2_outputs(7013) <= b;
    layer2_outputs(7014) <= a;
    layer2_outputs(7015) <= a and b;
    layer2_outputs(7016) <= not b or a;
    layer2_outputs(7017) <= a xor b;
    layer2_outputs(7018) <= not a;
    layer2_outputs(7019) <= not b;
    layer2_outputs(7020) <= not a;
    layer2_outputs(7021) <= b;
    layer2_outputs(7022) <= a and b;
    layer2_outputs(7023) <= not b or a;
    layer2_outputs(7024) <= not b;
    layer2_outputs(7025) <= not b;
    layer2_outputs(7026) <= not a or b;
    layer2_outputs(7027) <= not (a xor b);
    layer2_outputs(7028) <= not a;
    layer2_outputs(7029) <= a;
    layer2_outputs(7030) <= a and not b;
    layer2_outputs(7031) <= not (a or b);
    layer2_outputs(7032) <= a;
    layer2_outputs(7033) <= not a;
    layer2_outputs(7034) <= a and not b;
    layer2_outputs(7035) <= a;
    layer2_outputs(7036) <= not a;
    layer2_outputs(7037) <= a;
    layer2_outputs(7038) <= a xor b;
    layer2_outputs(7039) <= b;
    layer2_outputs(7040) <= not (a or b);
    layer2_outputs(7041) <= not b;
    layer2_outputs(7042) <= not a;
    layer2_outputs(7043) <= not (a and b);
    layer2_outputs(7044) <= a xor b;
    layer2_outputs(7045) <= a and b;
    layer2_outputs(7046) <= b;
    layer2_outputs(7047) <= a and b;
    layer2_outputs(7048) <= b;
    layer2_outputs(7049) <= not b or a;
    layer2_outputs(7050) <= b;
    layer2_outputs(7051) <= a or b;
    layer2_outputs(7052) <= a;
    layer2_outputs(7053) <= a or b;
    layer2_outputs(7054) <= not b;
    layer2_outputs(7055) <= not a or b;
    layer2_outputs(7056) <= not (a and b);
    layer2_outputs(7057) <= not b;
    layer2_outputs(7058) <= not a;
    layer2_outputs(7059) <= b;
    layer2_outputs(7060) <= a;
    layer2_outputs(7061) <= a and b;
    layer2_outputs(7062) <= not b;
    layer2_outputs(7063) <= a and not b;
    layer2_outputs(7064) <= not a or b;
    layer2_outputs(7065) <= a xor b;
    layer2_outputs(7066) <= a and not b;
    layer2_outputs(7067) <= a;
    layer2_outputs(7068) <= not (a or b);
    layer2_outputs(7069) <= a;
    layer2_outputs(7070) <= b;
    layer2_outputs(7071) <= not a or b;
    layer2_outputs(7072) <= not (a or b);
    layer2_outputs(7073) <= a xor b;
    layer2_outputs(7074) <= not b or a;
    layer2_outputs(7075) <= a xor b;
    layer2_outputs(7076) <= not b;
    layer2_outputs(7077) <= a;
    layer2_outputs(7078) <= not b or a;
    layer2_outputs(7079) <= not (a or b);
    layer2_outputs(7080) <= not (a or b);
    layer2_outputs(7081) <= not (a and b);
    layer2_outputs(7082) <= a xor b;
    layer2_outputs(7083) <= a;
    layer2_outputs(7084) <= a;
    layer2_outputs(7085) <= a or b;
    layer2_outputs(7086) <= a or b;
    layer2_outputs(7087) <= not (a or b);
    layer2_outputs(7088) <= not b or a;
    layer2_outputs(7089) <= b;
    layer2_outputs(7090) <= a or b;
    layer2_outputs(7091) <= not b or a;
    layer2_outputs(7092) <= a or b;
    layer2_outputs(7093) <= not b;
    layer2_outputs(7094) <= not (a xor b);
    layer2_outputs(7095) <= not a or b;
    layer2_outputs(7096) <= a or b;
    layer2_outputs(7097) <= b and not a;
    layer2_outputs(7098) <= b and not a;
    layer2_outputs(7099) <= a;
    layer2_outputs(7100) <= b and not a;
    layer2_outputs(7101) <= a and not b;
    layer2_outputs(7102) <= 1'b0;
    layer2_outputs(7103) <= a and b;
    layer2_outputs(7104) <= a and b;
    layer2_outputs(7105) <= not (a xor b);
    layer2_outputs(7106) <= not b or a;
    layer2_outputs(7107) <= not a or b;
    layer2_outputs(7108) <= a and b;
    layer2_outputs(7109) <= a;
    layer2_outputs(7110) <= not a;
    layer2_outputs(7111) <= a or b;
    layer2_outputs(7112) <= b and not a;
    layer2_outputs(7113) <= not (a xor b);
    layer2_outputs(7114) <= b;
    layer2_outputs(7115) <= not a or b;
    layer2_outputs(7116) <= not b;
    layer2_outputs(7117) <= a and b;
    layer2_outputs(7118) <= a and b;
    layer2_outputs(7119) <= not a;
    layer2_outputs(7120) <= b;
    layer2_outputs(7121) <= a and not b;
    layer2_outputs(7122) <= not a;
    layer2_outputs(7123) <= not (a xor b);
    layer2_outputs(7124) <= a;
    layer2_outputs(7125) <= b and not a;
    layer2_outputs(7126) <= not b or a;
    layer2_outputs(7127) <= a or b;
    layer2_outputs(7128) <= a and b;
    layer2_outputs(7129) <= not b or a;
    layer2_outputs(7130) <= not b;
    layer2_outputs(7131) <= a;
    layer2_outputs(7132) <= 1'b1;
    layer2_outputs(7133) <= a;
    layer2_outputs(7134) <= not a or b;
    layer2_outputs(7135) <= not b;
    layer2_outputs(7136) <= not (a xor b);
    layer2_outputs(7137) <= not b;
    layer2_outputs(7138) <= a or b;
    layer2_outputs(7139) <= not (a or b);
    layer2_outputs(7140) <= not a;
    layer2_outputs(7141) <= a and not b;
    layer2_outputs(7142) <= not (a and b);
    layer2_outputs(7143) <= b and not a;
    layer2_outputs(7144) <= a;
    layer2_outputs(7145) <= b;
    layer2_outputs(7146) <= b;
    layer2_outputs(7147) <= a or b;
    layer2_outputs(7148) <= not b;
    layer2_outputs(7149) <= not (a or b);
    layer2_outputs(7150) <= not b;
    layer2_outputs(7151) <= a xor b;
    layer2_outputs(7152) <= b and not a;
    layer2_outputs(7153) <= a;
    layer2_outputs(7154) <= not b;
    layer2_outputs(7155) <= not (a xor b);
    layer2_outputs(7156) <= a and b;
    layer2_outputs(7157) <= b;
    layer2_outputs(7158) <= a and not b;
    layer2_outputs(7159) <= 1'b0;
    layer2_outputs(7160) <= not b or a;
    layer2_outputs(7161) <= not a or b;
    layer2_outputs(7162) <= not (a xor b);
    layer2_outputs(7163) <= a xor b;
    layer2_outputs(7164) <= not b;
    layer2_outputs(7165) <= b;
    layer2_outputs(7166) <= a xor b;
    layer2_outputs(7167) <= not b;
    layer2_outputs(7168) <= not b or a;
    layer2_outputs(7169) <= a xor b;
    layer2_outputs(7170) <= a xor b;
    layer2_outputs(7171) <= b and not a;
    layer2_outputs(7172) <= a and b;
    layer2_outputs(7173) <= a or b;
    layer2_outputs(7174) <= a or b;
    layer2_outputs(7175) <= not (a xor b);
    layer2_outputs(7176) <= b and not a;
    layer2_outputs(7177) <= not (a or b);
    layer2_outputs(7178) <= not b or a;
    layer2_outputs(7179) <= not a or b;
    layer2_outputs(7180) <= not a;
    layer2_outputs(7181) <= not b;
    layer2_outputs(7182) <= b;
    layer2_outputs(7183) <= a and not b;
    layer2_outputs(7184) <= a;
    layer2_outputs(7185) <= not (a or b);
    layer2_outputs(7186) <= b;
    layer2_outputs(7187) <= a and not b;
    layer2_outputs(7188) <= a and b;
    layer2_outputs(7189) <= a or b;
    layer2_outputs(7190) <= not b or a;
    layer2_outputs(7191) <= not a;
    layer2_outputs(7192) <= not (a xor b);
    layer2_outputs(7193) <= not b;
    layer2_outputs(7194) <= not (a or b);
    layer2_outputs(7195) <= a and not b;
    layer2_outputs(7196) <= not b;
    layer2_outputs(7197) <= not a;
    layer2_outputs(7198) <= not b or a;
    layer2_outputs(7199) <= a;
    layer2_outputs(7200) <= a xor b;
    layer2_outputs(7201) <= not a;
    layer2_outputs(7202) <= a;
    layer2_outputs(7203) <= not b;
    layer2_outputs(7204) <= b;
    layer2_outputs(7205) <= a or b;
    layer2_outputs(7206) <= a and not b;
    layer2_outputs(7207) <= b and not a;
    layer2_outputs(7208) <= a xor b;
    layer2_outputs(7209) <= a and b;
    layer2_outputs(7210) <= a;
    layer2_outputs(7211) <= a or b;
    layer2_outputs(7212) <= not b;
    layer2_outputs(7213) <= not b or a;
    layer2_outputs(7214) <= not a;
    layer2_outputs(7215) <= not (a xor b);
    layer2_outputs(7216) <= a or b;
    layer2_outputs(7217) <= not (a and b);
    layer2_outputs(7218) <= a;
    layer2_outputs(7219) <= not (a and b);
    layer2_outputs(7220) <= a;
    layer2_outputs(7221) <= not a or b;
    layer2_outputs(7222) <= a and b;
    layer2_outputs(7223) <= b;
    layer2_outputs(7224) <= not a;
    layer2_outputs(7225) <= not a or b;
    layer2_outputs(7226) <= not b;
    layer2_outputs(7227) <= not (a and b);
    layer2_outputs(7228) <= not (a and b);
    layer2_outputs(7229) <= b and not a;
    layer2_outputs(7230) <= not b or a;
    layer2_outputs(7231) <= not b or a;
    layer2_outputs(7232) <= b;
    layer2_outputs(7233) <= not a or b;
    layer2_outputs(7234) <= a xor b;
    layer2_outputs(7235) <= not (a xor b);
    layer2_outputs(7236) <= not b;
    layer2_outputs(7237) <= a;
    layer2_outputs(7238) <= b;
    layer2_outputs(7239) <= not b;
    layer2_outputs(7240) <= b;
    layer2_outputs(7241) <= a xor b;
    layer2_outputs(7242) <= not b;
    layer2_outputs(7243) <= not a;
    layer2_outputs(7244) <= not (a xor b);
    layer2_outputs(7245) <= a xor b;
    layer2_outputs(7246) <= a;
    layer2_outputs(7247) <= not b;
    layer2_outputs(7248) <= a;
    layer2_outputs(7249) <= not (a or b);
    layer2_outputs(7250) <= not b;
    layer2_outputs(7251) <= a xor b;
    layer2_outputs(7252) <= not (a xor b);
    layer2_outputs(7253) <= b;
    layer2_outputs(7254) <= a;
    layer2_outputs(7255) <= b;
    layer2_outputs(7256) <= not a;
    layer2_outputs(7257) <= not a;
    layer2_outputs(7258) <= not b;
    layer2_outputs(7259) <= not (a and b);
    layer2_outputs(7260) <= b and not a;
    layer2_outputs(7261) <= a xor b;
    layer2_outputs(7262) <= not b or a;
    layer2_outputs(7263) <= not (a xor b);
    layer2_outputs(7264) <= not (a or b);
    layer2_outputs(7265) <= not b;
    layer2_outputs(7266) <= not b or a;
    layer2_outputs(7267) <= not a or b;
    layer2_outputs(7268) <= b;
    layer2_outputs(7269) <= a xor b;
    layer2_outputs(7270) <= a or b;
    layer2_outputs(7271) <= b and not a;
    layer2_outputs(7272) <= not (a xor b);
    layer2_outputs(7273) <= b and not a;
    layer2_outputs(7274) <= not b or a;
    layer2_outputs(7275) <= b;
    layer2_outputs(7276) <= not (a xor b);
    layer2_outputs(7277) <= a and b;
    layer2_outputs(7278) <= a xor b;
    layer2_outputs(7279) <= not (a and b);
    layer2_outputs(7280) <= not b;
    layer2_outputs(7281) <= not b;
    layer2_outputs(7282) <= not a;
    layer2_outputs(7283) <= not a or b;
    layer2_outputs(7284) <= not (a xor b);
    layer2_outputs(7285) <= a;
    layer2_outputs(7286) <= not (a xor b);
    layer2_outputs(7287) <= not a;
    layer2_outputs(7288) <= not (a and b);
    layer2_outputs(7289) <= not b;
    layer2_outputs(7290) <= a;
    layer2_outputs(7291) <= not b or a;
    layer2_outputs(7292) <= not a;
    layer2_outputs(7293) <= b;
    layer2_outputs(7294) <= not a or b;
    layer2_outputs(7295) <= not (a and b);
    layer2_outputs(7296) <= a and b;
    layer2_outputs(7297) <= not (a and b);
    layer2_outputs(7298) <= a and b;
    layer2_outputs(7299) <= a;
    layer2_outputs(7300) <= not b;
    layer2_outputs(7301) <= a xor b;
    layer2_outputs(7302) <= a and b;
    layer2_outputs(7303) <= b;
    layer2_outputs(7304) <= not b;
    layer2_outputs(7305) <= not a;
    layer2_outputs(7306) <= a or b;
    layer2_outputs(7307) <= a xor b;
    layer2_outputs(7308) <= not a or b;
    layer2_outputs(7309) <= not a;
    layer2_outputs(7310) <= b;
    layer2_outputs(7311) <= a and not b;
    layer2_outputs(7312) <= a xor b;
    layer2_outputs(7313) <= b;
    layer2_outputs(7314) <= 1'b0;
    layer2_outputs(7315) <= a and not b;
    layer2_outputs(7316) <= a;
    layer2_outputs(7317) <= b;
    layer2_outputs(7318) <= a;
    layer2_outputs(7319) <= not (a and b);
    layer2_outputs(7320) <= a and not b;
    layer2_outputs(7321) <= not (a and b);
    layer2_outputs(7322) <= not a or b;
    layer2_outputs(7323) <= not a;
    layer2_outputs(7324) <= not a or b;
    layer2_outputs(7325) <= not (a and b);
    layer2_outputs(7326) <= not a;
    layer2_outputs(7327) <= not a;
    layer2_outputs(7328) <= b and not a;
    layer2_outputs(7329) <= a xor b;
    layer2_outputs(7330) <= a or b;
    layer2_outputs(7331) <= b;
    layer2_outputs(7332) <= a;
    layer2_outputs(7333) <= a;
    layer2_outputs(7334) <= not (a or b);
    layer2_outputs(7335) <= not (a or b);
    layer2_outputs(7336) <= not b;
    layer2_outputs(7337) <= a or b;
    layer2_outputs(7338) <= not (a or b);
    layer2_outputs(7339) <= not b;
    layer2_outputs(7340) <= not b;
    layer2_outputs(7341) <= a and not b;
    layer2_outputs(7342) <= not (a or b);
    layer2_outputs(7343) <= a and b;
    layer2_outputs(7344) <= not b or a;
    layer2_outputs(7345) <= a or b;
    layer2_outputs(7346) <= a and b;
    layer2_outputs(7347) <= b;
    layer2_outputs(7348) <= not b;
    layer2_outputs(7349) <= not b or a;
    layer2_outputs(7350) <= a and not b;
    layer2_outputs(7351) <= a;
    layer2_outputs(7352) <= not a;
    layer2_outputs(7353) <= a xor b;
    layer2_outputs(7354) <= not (a xor b);
    layer2_outputs(7355) <= b;
    layer2_outputs(7356) <= not (a or b);
    layer2_outputs(7357) <= a or b;
    layer2_outputs(7358) <= a or b;
    layer2_outputs(7359) <= not (a xor b);
    layer2_outputs(7360) <= not a;
    layer2_outputs(7361) <= a or b;
    layer2_outputs(7362) <= a or b;
    layer2_outputs(7363) <= not a;
    layer2_outputs(7364) <= not a;
    layer2_outputs(7365) <= b;
    layer2_outputs(7366) <= a;
    layer2_outputs(7367) <= not (a xor b);
    layer2_outputs(7368) <= a or b;
    layer2_outputs(7369) <= not a;
    layer2_outputs(7370) <= a and not b;
    layer2_outputs(7371) <= b;
    layer2_outputs(7372) <= b;
    layer2_outputs(7373) <= b and not a;
    layer2_outputs(7374) <= b and not a;
    layer2_outputs(7375) <= not (a xor b);
    layer2_outputs(7376) <= a or b;
    layer2_outputs(7377) <= a xor b;
    layer2_outputs(7378) <= a xor b;
    layer2_outputs(7379) <= a and not b;
    layer2_outputs(7380) <= a;
    layer2_outputs(7381) <= not a;
    layer2_outputs(7382) <= not (a xor b);
    layer2_outputs(7383) <= a;
    layer2_outputs(7384) <= not a or b;
    layer2_outputs(7385) <= a and not b;
    layer2_outputs(7386) <= not a;
    layer2_outputs(7387) <= a and not b;
    layer2_outputs(7388) <= a and b;
    layer2_outputs(7389) <= a xor b;
    layer2_outputs(7390) <= not (a and b);
    layer2_outputs(7391) <= not (a and b);
    layer2_outputs(7392) <= not (a and b);
    layer2_outputs(7393) <= not b;
    layer2_outputs(7394) <= b;
    layer2_outputs(7395) <= not a;
    layer2_outputs(7396) <= not (a or b);
    layer2_outputs(7397) <= a xor b;
    layer2_outputs(7398) <= a or b;
    layer2_outputs(7399) <= a xor b;
    layer2_outputs(7400) <= not b;
    layer2_outputs(7401) <= a xor b;
    layer2_outputs(7402) <= a and not b;
    layer2_outputs(7403) <= not b or a;
    layer2_outputs(7404) <= a;
    layer2_outputs(7405) <= a;
    layer2_outputs(7406) <= not (a or b);
    layer2_outputs(7407) <= a and b;
    layer2_outputs(7408) <= a xor b;
    layer2_outputs(7409) <= a or b;
    layer2_outputs(7410) <= not (a and b);
    layer2_outputs(7411) <= not b;
    layer2_outputs(7412) <= not b;
    layer2_outputs(7413) <= not (a and b);
    layer2_outputs(7414) <= a;
    layer2_outputs(7415) <= not a;
    layer2_outputs(7416) <= 1'b0;
    layer2_outputs(7417) <= b;
    layer2_outputs(7418) <= a xor b;
    layer2_outputs(7419) <= a xor b;
    layer2_outputs(7420) <= not (a xor b);
    layer2_outputs(7421) <= a xor b;
    layer2_outputs(7422) <= a;
    layer2_outputs(7423) <= a;
    layer2_outputs(7424) <= not (a or b);
    layer2_outputs(7425) <= not (a and b);
    layer2_outputs(7426) <= not (a and b);
    layer2_outputs(7427) <= not (a xor b);
    layer2_outputs(7428) <= not b or a;
    layer2_outputs(7429) <= a and not b;
    layer2_outputs(7430) <= not b;
    layer2_outputs(7431) <= a and b;
    layer2_outputs(7432) <= not a or b;
    layer2_outputs(7433) <= a xor b;
    layer2_outputs(7434) <= b and not a;
    layer2_outputs(7435) <= b;
    layer2_outputs(7436) <= a;
    layer2_outputs(7437) <= a and not b;
    layer2_outputs(7438) <= not b or a;
    layer2_outputs(7439) <= not (a or b);
    layer2_outputs(7440) <= not (a xor b);
    layer2_outputs(7441) <= a;
    layer2_outputs(7442) <= 1'b0;
    layer2_outputs(7443) <= not (a xor b);
    layer2_outputs(7444) <= not b or a;
    layer2_outputs(7445) <= a;
    layer2_outputs(7446) <= not (a xor b);
    layer2_outputs(7447) <= not b or a;
    layer2_outputs(7448) <= not a or b;
    layer2_outputs(7449) <= not b or a;
    layer2_outputs(7450) <= not (a xor b);
    layer2_outputs(7451) <= a and b;
    layer2_outputs(7452) <= b and not a;
    layer2_outputs(7453) <= not b;
    layer2_outputs(7454) <= not (a xor b);
    layer2_outputs(7455) <= not (a and b);
    layer2_outputs(7456) <= not (a xor b);
    layer2_outputs(7457) <= a and not b;
    layer2_outputs(7458) <= a and b;
    layer2_outputs(7459) <= not (a and b);
    layer2_outputs(7460) <= a or b;
    layer2_outputs(7461) <= b and not a;
    layer2_outputs(7462) <= not (a or b);
    layer2_outputs(7463) <= not b;
    layer2_outputs(7464) <= b;
    layer2_outputs(7465) <= a and b;
    layer2_outputs(7466) <= a and not b;
    layer2_outputs(7467) <= not (a xor b);
    layer2_outputs(7468) <= b;
    layer2_outputs(7469) <= a;
    layer2_outputs(7470) <= a;
    layer2_outputs(7471) <= a;
    layer2_outputs(7472) <= b;
    layer2_outputs(7473) <= not (a and b);
    layer2_outputs(7474) <= a and not b;
    layer2_outputs(7475) <= not b;
    layer2_outputs(7476) <= not b;
    layer2_outputs(7477) <= not (a or b);
    layer2_outputs(7478) <= not b;
    layer2_outputs(7479) <= not a;
    layer2_outputs(7480) <= not a;
    layer2_outputs(7481) <= not b;
    layer2_outputs(7482) <= a;
    layer2_outputs(7483) <= not (a and b);
    layer2_outputs(7484) <= not b or a;
    layer2_outputs(7485) <= not a;
    layer2_outputs(7486) <= a and not b;
    layer2_outputs(7487) <= a or b;
    layer2_outputs(7488) <= a;
    layer2_outputs(7489) <= not a;
    layer2_outputs(7490) <= a and b;
    layer2_outputs(7491) <= b and not a;
    layer2_outputs(7492) <= not b;
    layer2_outputs(7493) <= not (a and b);
    layer2_outputs(7494) <= b;
    layer2_outputs(7495) <= not a;
    layer2_outputs(7496) <= 1'b0;
    layer2_outputs(7497) <= b;
    layer2_outputs(7498) <= not b;
    layer2_outputs(7499) <= a;
    layer2_outputs(7500) <= b;
    layer2_outputs(7501) <= a;
    layer2_outputs(7502) <= not (a xor b);
    layer2_outputs(7503) <= not a or b;
    layer2_outputs(7504) <= a xor b;
    layer2_outputs(7505) <= a xor b;
    layer2_outputs(7506) <= a xor b;
    layer2_outputs(7507) <= 1'b0;
    layer2_outputs(7508) <= not a;
    layer2_outputs(7509) <= not a;
    layer2_outputs(7510) <= a and b;
    layer2_outputs(7511) <= not b;
    layer2_outputs(7512) <= not b;
    layer2_outputs(7513) <= not (a and b);
    layer2_outputs(7514) <= not a;
    layer2_outputs(7515) <= not b;
    layer2_outputs(7516) <= a or b;
    layer2_outputs(7517) <= not b;
    layer2_outputs(7518) <= not (a and b);
    layer2_outputs(7519) <= b;
    layer2_outputs(7520) <= a;
    layer2_outputs(7521) <= a xor b;
    layer2_outputs(7522) <= b and not a;
    layer2_outputs(7523) <= not (a or b);
    layer2_outputs(7524) <= a;
    layer2_outputs(7525) <= a and not b;
    layer2_outputs(7526) <= b and not a;
    layer2_outputs(7527) <= not (a xor b);
    layer2_outputs(7528) <= a and not b;
    layer2_outputs(7529) <= not a;
    layer2_outputs(7530) <= not (a and b);
    layer2_outputs(7531) <= b;
    layer2_outputs(7532) <= not (a and b);
    layer2_outputs(7533) <= not a or b;
    layer2_outputs(7534) <= a or b;
    layer2_outputs(7535) <= not (a xor b);
    layer2_outputs(7536) <= not b;
    layer2_outputs(7537) <= b and not a;
    layer2_outputs(7538) <= a and b;
    layer2_outputs(7539) <= not a;
    layer2_outputs(7540) <= not a;
    layer2_outputs(7541) <= not (a or b);
    layer2_outputs(7542) <= not (a xor b);
    layer2_outputs(7543) <= not b;
    layer2_outputs(7544) <= not a;
    layer2_outputs(7545) <= b;
    layer2_outputs(7546) <= not (a xor b);
    layer2_outputs(7547) <= not a;
    layer2_outputs(7548) <= a and not b;
    layer2_outputs(7549) <= a xor b;
    layer2_outputs(7550) <= b and not a;
    layer2_outputs(7551) <= not a;
    layer2_outputs(7552) <= b;
    layer2_outputs(7553) <= not a;
    layer2_outputs(7554) <= a;
    layer2_outputs(7555) <= not b;
    layer2_outputs(7556) <= not a or b;
    layer2_outputs(7557) <= b and not a;
    layer2_outputs(7558) <= a or b;
    layer2_outputs(7559) <= not a;
    layer2_outputs(7560) <= not a;
    layer2_outputs(7561) <= not b;
    layer2_outputs(7562) <= a and b;
    layer2_outputs(7563) <= a xor b;
    layer2_outputs(7564) <= not b;
    layer2_outputs(7565) <= b;
    layer2_outputs(7566) <= b;
    layer2_outputs(7567) <= a and not b;
    layer2_outputs(7568) <= b;
    layer2_outputs(7569) <= not b;
    layer2_outputs(7570) <= not a;
    layer2_outputs(7571) <= not (a and b);
    layer2_outputs(7572) <= b and not a;
    layer2_outputs(7573) <= not (a xor b);
    layer2_outputs(7574) <= not (a and b);
    layer2_outputs(7575) <= not a;
    layer2_outputs(7576) <= a and b;
    layer2_outputs(7577) <= not b;
    layer2_outputs(7578) <= not (a xor b);
    layer2_outputs(7579) <= not (a and b);
    layer2_outputs(7580) <= b;
    layer2_outputs(7581) <= b;
    layer2_outputs(7582) <= not b;
    layer2_outputs(7583) <= not b;
    layer2_outputs(7584) <= not a;
    layer2_outputs(7585) <= not (a and b);
    layer2_outputs(7586) <= not (a and b);
    layer2_outputs(7587) <= not (a or b);
    layer2_outputs(7588) <= a;
    layer2_outputs(7589) <= not (a xor b);
    layer2_outputs(7590) <= not a;
    layer2_outputs(7591) <= not a or b;
    layer2_outputs(7592) <= a xor b;
    layer2_outputs(7593) <= b;
    layer2_outputs(7594) <= a or b;
    layer2_outputs(7595) <= not a or b;
    layer2_outputs(7596) <= a or b;
    layer2_outputs(7597) <= not b or a;
    layer2_outputs(7598) <= not a;
    layer2_outputs(7599) <= not b or a;
    layer2_outputs(7600) <= a or b;
    layer2_outputs(7601) <= not (a xor b);
    layer2_outputs(7602) <= not a;
    layer2_outputs(7603) <= a;
    layer2_outputs(7604) <= b;
    layer2_outputs(7605) <= not b or a;
    layer2_outputs(7606) <= not (a or b);
    layer2_outputs(7607) <= not (a and b);
    layer2_outputs(7608) <= b;
    layer2_outputs(7609) <= not (a and b);
    layer2_outputs(7610) <= a and b;
    layer2_outputs(7611) <= not (a and b);
    layer2_outputs(7612) <= a;
    layer2_outputs(7613) <= not (a xor b);
    layer2_outputs(7614) <= not (a or b);
    layer2_outputs(7615) <= not (a and b);
    layer2_outputs(7616) <= not a or b;
    layer2_outputs(7617) <= not b or a;
    layer2_outputs(7618) <= a xor b;
    layer2_outputs(7619) <= a and not b;
    layer2_outputs(7620) <= a and not b;
    layer2_outputs(7621) <= b;
    layer2_outputs(7622) <= not (a or b);
    layer2_outputs(7623) <= a xor b;
    layer2_outputs(7624) <= a and b;
    layer2_outputs(7625) <= a or b;
    layer2_outputs(7626) <= not a;
    layer2_outputs(7627) <= not b;
    layer2_outputs(7628) <= not a;
    layer2_outputs(7629) <= a and not b;
    layer2_outputs(7630) <= not (a or b);
    layer2_outputs(7631) <= a xor b;
    layer2_outputs(7632) <= a and b;
    layer2_outputs(7633) <= a xor b;
    layer2_outputs(7634) <= a;
    layer2_outputs(7635) <= b;
    layer2_outputs(7636) <= not (a and b);
    layer2_outputs(7637) <= a and b;
    layer2_outputs(7638) <= b;
    layer2_outputs(7639) <= a and not b;
    layer2_outputs(7640) <= not (a and b);
    layer2_outputs(7641) <= not a or b;
    layer2_outputs(7642) <= a and not b;
    layer2_outputs(7643) <= a;
    layer2_outputs(7644) <= a or b;
    layer2_outputs(7645) <= b;
    layer2_outputs(7646) <= not a;
    layer2_outputs(7647) <= a and b;
    layer2_outputs(7648) <= b;
    layer2_outputs(7649) <= not a;
    layer2_outputs(7650) <= not (a or b);
    layer2_outputs(7651) <= not b;
    layer2_outputs(7652) <= a;
    layer2_outputs(7653) <= a or b;
    layer2_outputs(7654) <= b;
    layer2_outputs(7655) <= not b;
    layer2_outputs(7656) <= b;
    layer2_outputs(7657) <= b and not a;
    layer2_outputs(7658) <= a xor b;
    layer2_outputs(7659) <= not a;
    layer2_outputs(7660) <= a or b;
    layer2_outputs(7661) <= a and not b;
    layer2_outputs(7662) <= not (a xor b);
    layer2_outputs(7663) <= a and not b;
    layer2_outputs(7664) <= not a;
    layer2_outputs(7665) <= a;
    layer2_outputs(7666) <= a xor b;
    layer2_outputs(7667) <= b;
    layer2_outputs(7668) <= a or b;
    layer2_outputs(7669) <= a and b;
    layer2_outputs(7670) <= a or b;
    layer2_outputs(7671) <= a and not b;
    layer2_outputs(7672) <= a;
    layer2_outputs(7673) <= not b or a;
    layer2_outputs(7674) <= not b or a;
    layer2_outputs(7675) <= a;
    layer2_outputs(7676) <= not b or a;
    layer2_outputs(7677) <= a and b;
    layer2_outputs(7678) <= a or b;
    layer2_outputs(7679) <= a and not b;
    outputs(0) <= not (a and b);
    outputs(1) <= not a;
    outputs(2) <= not b;
    outputs(3) <= not a;
    outputs(4) <= not b;
    outputs(5) <= a xor b;
    outputs(6) <= a xor b;
    outputs(7) <= not a;
    outputs(8) <= not b;
    outputs(9) <= not b;
    outputs(10) <= a and not b;
    outputs(11) <= b;
    outputs(12) <= not (a xor b);
    outputs(13) <= not b;
    outputs(14) <= not (a xor b);
    outputs(15) <= not b;
    outputs(16) <= b;
    outputs(17) <= not (a xor b);
    outputs(18) <= b and not a;
    outputs(19) <= not (a or b);
    outputs(20) <= not b or a;
    outputs(21) <= not a;
    outputs(22) <= not b;
    outputs(23) <= b;
    outputs(24) <= not b;
    outputs(25) <= not a;
    outputs(26) <= not b;
    outputs(27) <= not b;
    outputs(28) <= not b;
    outputs(29) <= a and not b;
    outputs(30) <= not b;
    outputs(31) <= not b;
    outputs(32) <= not a;
    outputs(33) <= a xor b;
    outputs(34) <= not b;
    outputs(35) <= a xor b;
    outputs(36) <= not (a or b);
    outputs(37) <= b and not a;
    outputs(38) <= not a;
    outputs(39) <= a and b;
    outputs(40) <= a xor b;
    outputs(41) <= a and b;
    outputs(42) <= not a;
    outputs(43) <= a;
    outputs(44) <= not b;
    outputs(45) <= a xor b;
    outputs(46) <= not (a xor b);
    outputs(47) <= not (a and b);
    outputs(48) <= b and not a;
    outputs(49) <= not (a or b);
    outputs(50) <= b;
    outputs(51) <= a and b;
    outputs(52) <= not (a and b);
    outputs(53) <= a;
    outputs(54) <= b;
    outputs(55) <= a and not b;
    outputs(56) <= a;
    outputs(57) <= a xor b;
    outputs(58) <= a and b;
    outputs(59) <= a;
    outputs(60) <= a and not b;
    outputs(61) <= a and not b;
    outputs(62) <= not (a or b);
    outputs(63) <= a xor b;
    outputs(64) <= not a or b;
    outputs(65) <= a and not b;
    outputs(66) <= not b;
    outputs(67) <= a and not b;
    outputs(68) <= a;
    outputs(69) <= not (a and b);
    outputs(70) <= not a;
    outputs(71) <= not (a xor b);
    outputs(72) <= a;
    outputs(73) <= b;
    outputs(74) <= not (a or b);
    outputs(75) <= not b;
    outputs(76) <= a and b;
    outputs(77) <= a or b;
    outputs(78) <= not b;
    outputs(79) <= not (a xor b);
    outputs(80) <= not a or b;
    outputs(81) <= a;
    outputs(82) <= b and not a;
    outputs(83) <= a and b;
    outputs(84) <= a and not b;
    outputs(85) <= a xor b;
    outputs(86) <= a;
    outputs(87) <= not (a and b);
    outputs(88) <= b and not a;
    outputs(89) <= not (a xor b);
    outputs(90) <= not a;
    outputs(91) <= not (a xor b);
    outputs(92) <= not b;
    outputs(93) <= not a;
    outputs(94) <= a xor b;
    outputs(95) <= a or b;
    outputs(96) <= not (a xor b);
    outputs(97) <= not (a xor b);
    outputs(98) <= not a;
    outputs(99) <= not b;
    outputs(100) <= b;
    outputs(101) <= not a;
    outputs(102) <= b;
    outputs(103) <= not a;
    outputs(104) <= a and not b;
    outputs(105) <= b;
    outputs(106) <= b;
    outputs(107) <= not (a or b);
    outputs(108) <= not (a or b);
    outputs(109) <= b and not a;
    outputs(110) <= not a or b;
    outputs(111) <= not (a or b);
    outputs(112) <= b;
    outputs(113) <= b;
    outputs(114) <= a;
    outputs(115) <= not b or a;
    outputs(116) <= b;
    outputs(117) <= b and not a;
    outputs(118) <= a;
    outputs(119) <= a and not b;
    outputs(120) <= a and b;
    outputs(121) <= a;
    outputs(122) <= not (a xor b);
    outputs(123) <= b;
    outputs(124) <= not b or a;
    outputs(125) <= b and not a;
    outputs(126) <= not (a or b);
    outputs(127) <= not a;
    outputs(128) <= not (a xor b);
    outputs(129) <= not (a xor b);
    outputs(130) <= a and b;
    outputs(131) <= a;
    outputs(132) <= not (a or b);
    outputs(133) <= not a;
    outputs(134) <= b;
    outputs(135) <= not b;
    outputs(136) <= b;
    outputs(137) <= a and b;
    outputs(138) <= not a;
    outputs(139) <= not (a or b);
    outputs(140) <= not (a and b);
    outputs(141) <= a;
    outputs(142) <= not b or a;
    outputs(143) <= b and not a;
    outputs(144) <= a;
    outputs(145) <= not b;
    outputs(146) <= b;
    outputs(147) <= not b;
    outputs(148) <= a xor b;
    outputs(149) <= not a;
    outputs(150) <= a and not b;
    outputs(151) <= a;
    outputs(152) <= not b;
    outputs(153) <= a;
    outputs(154) <= b;
    outputs(155) <= not a or b;
    outputs(156) <= not b;
    outputs(157) <= a and not b;
    outputs(158) <= not (a and b);
    outputs(159) <= a and b;
    outputs(160) <= not a or b;
    outputs(161) <= a xor b;
    outputs(162) <= b and not a;
    outputs(163) <= b and not a;
    outputs(164) <= b;
    outputs(165) <= b;
    outputs(166) <= a xor b;
    outputs(167) <= not a;
    outputs(168) <= a and not b;
    outputs(169) <= a xor b;
    outputs(170) <= not b;
    outputs(171) <= a and not b;
    outputs(172) <= not a;
    outputs(173) <= a;
    outputs(174) <= not b or a;
    outputs(175) <= b and not a;
    outputs(176) <= not a;
    outputs(177) <= not (a xor b);
    outputs(178) <= a;
    outputs(179) <= a xor b;
    outputs(180) <= a or b;
    outputs(181) <= not (a xor b);
    outputs(182) <= not b;
    outputs(183) <= not a;
    outputs(184) <= not b;
    outputs(185) <= a and b;
    outputs(186) <= a xor b;
    outputs(187) <= a or b;
    outputs(188) <= a;
    outputs(189) <= not b;
    outputs(190) <= not (a xor b);
    outputs(191) <= b and not a;
    outputs(192) <= a;
    outputs(193) <= b and not a;
    outputs(194) <= b;
    outputs(195) <= not b;
    outputs(196) <= a;
    outputs(197) <= a;
    outputs(198) <= not b;
    outputs(199) <= a xor b;
    outputs(200) <= a;
    outputs(201) <= a or b;
    outputs(202) <= b;
    outputs(203) <= b;
    outputs(204) <= not (a and b);
    outputs(205) <= a and b;
    outputs(206) <= not a;
    outputs(207) <= a or b;
    outputs(208) <= not a;
    outputs(209) <= a and not b;
    outputs(210) <= b;
    outputs(211) <= a;
    outputs(212) <= not (a and b);
    outputs(213) <= a and not b;
    outputs(214) <= not (a or b);
    outputs(215) <= not (a and b);
    outputs(216) <= a;
    outputs(217) <= a;
    outputs(218) <= b;
    outputs(219) <= a and not b;
    outputs(220) <= not (a and b);
    outputs(221) <= not b;
    outputs(222) <= 1'b0;
    outputs(223) <= not (a xor b);
    outputs(224) <= a;
    outputs(225) <= a xor b;
    outputs(226) <= b;
    outputs(227) <= a and not b;
    outputs(228) <= not a;
    outputs(229) <= not b or a;
    outputs(230) <= a xor b;
    outputs(231) <= a xor b;
    outputs(232) <= not b;
    outputs(233) <= b;
    outputs(234) <= b and not a;
    outputs(235) <= a xor b;
    outputs(236) <= b;
    outputs(237) <= not b;
    outputs(238) <= not a;
    outputs(239) <= a;
    outputs(240) <= a and b;
    outputs(241) <= not b;
    outputs(242) <= not b or a;
    outputs(243) <= not (a or b);
    outputs(244) <= a and not b;
    outputs(245) <= not b;
    outputs(246) <= a or b;
    outputs(247) <= b;
    outputs(248) <= a and not b;
    outputs(249) <= b and not a;
    outputs(250) <= not (a xor b);
    outputs(251) <= a xor b;
    outputs(252) <= not a or b;
    outputs(253) <= not (a or b);
    outputs(254) <= b;
    outputs(255) <= not b;
    outputs(256) <= not a;
    outputs(257) <= b;
    outputs(258) <= not a;
    outputs(259) <= not b;
    outputs(260) <= not (a or b);
    outputs(261) <= a xor b;
    outputs(262) <= not (a xor b);
    outputs(263) <= b and not a;
    outputs(264) <= a;
    outputs(265) <= b;
    outputs(266) <= not (a and b);
    outputs(267) <= a and b;
    outputs(268) <= a;
    outputs(269) <= not a;
    outputs(270) <= not a;
    outputs(271) <= not b or a;
    outputs(272) <= a;
    outputs(273) <= not b;
    outputs(274) <= not a;
    outputs(275) <= a xor b;
    outputs(276) <= not (a and b);
    outputs(277) <= a and not b;
    outputs(278) <= a;
    outputs(279) <= not (a and b);
    outputs(280) <= not b or a;
    outputs(281) <= a and b;
    outputs(282) <= b;
    outputs(283) <= a and not b;
    outputs(284) <= b;
    outputs(285) <= not b;
    outputs(286) <= not b;
    outputs(287) <= a xor b;
    outputs(288) <= not b;
    outputs(289) <= a;
    outputs(290) <= a and not b;
    outputs(291) <= a and b;
    outputs(292) <= not a;
    outputs(293) <= not (a or b);
    outputs(294) <= a;
    outputs(295) <= a;
    outputs(296) <= not (a xor b);
    outputs(297) <= b;
    outputs(298) <= b;
    outputs(299) <= a xor b;
    outputs(300) <= b;
    outputs(301) <= a;
    outputs(302) <= not (a or b);
    outputs(303) <= not (a or b);
    outputs(304) <= a and b;
    outputs(305) <= a xor b;
    outputs(306) <= not a;
    outputs(307) <= a;
    outputs(308) <= not b;
    outputs(309) <= b and not a;
    outputs(310) <= a;
    outputs(311) <= not a or b;
    outputs(312) <= not (a or b);
    outputs(313) <= a xor b;
    outputs(314) <= not b or a;
    outputs(315) <= not b;
    outputs(316) <= a and b;
    outputs(317) <= not b;
    outputs(318) <= b;
    outputs(319) <= b;
    outputs(320) <= not (a xor b);
    outputs(321) <= a and not b;
    outputs(322) <= a;
    outputs(323) <= b;
    outputs(324) <= b;
    outputs(325) <= not b;
    outputs(326) <= a xor b;
    outputs(327) <= a;
    outputs(328) <= b;
    outputs(329) <= not b;
    outputs(330) <= a and not b;
    outputs(331) <= a and not b;
    outputs(332) <= b;
    outputs(333) <= not a;
    outputs(334) <= not a;
    outputs(335) <= a;
    outputs(336) <= a or b;
    outputs(337) <= not (a xor b);
    outputs(338) <= a and b;
    outputs(339) <= a;
    outputs(340) <= not (a xor b);
    outputs(341) <= b and not a;
    outputs(342) <= a and not b;
    outputs(343) <= not a;
    outputs(344) <= a xor b;
    outputs(345) <= not b;
    outputs(346) <= a and not b;
    outputs(347) <= a or b;
    outputs(348) <= b and not a;
    outputs(349) <= a;
    outputs(350) <= b and not a;
    outputs(351) <= not (a or b);
    outputs(352) <= not (a xor b);
    outputs(353) <= a;
    outputs(354) <= not b;
    outputs(355) <= a xor b;
    outputs(356) <= b;
    outputs(357) <= not (a and b);
    outputs(358) <= not (a xor b);
    outputs(359) <= not (a xor b);
    outputs(360) <= a xor b;
    outputs(361) <= not b;
    outputs(362) <= not b or a;
    outputs(363) <= not a;
    outputs(364) <= not a or b;
    outputs(365) <= not b;
    outputs(366) <= a xor b;
    outputs(367) <= b and not a;
    outputs(368) <= b and not a;
    outputs(369) <= not b;
    outputs(370) <= a xor b;
    outputs(371) <= not b;
    outputs(372) <= a xor b;
    outputs(373) <= not b;
    outputs(374) <= a;
    outputs(375) <= a;
    outputs(376) <= not b;
    outputs(377) <= a and b;
    outputs(378) <= a and b;
    outputs(379) <= not a;
    outputs(380) <= a xor b;
    outputs(381) <= a xor b;
    outputs(382) <= a or b;
    outputs(383) <= a and not b;
    outputs(384) <= a;
    outputs(385) <= a xor b;
    outputs(386) <= b;
    outputs(387) <= not b;
    outputs(388) <= not (a xor b);
    outputs(389) <= a and b;
    outputs(390) <= a xor b;
    outputs(391) <= a;
    outputs(392) <= a;
    outputs(393) <= not a;
    outputs(394) <= not (a and b);
    outputs(395) <= not a;
    outputs(396) <= b;
    outputs(397) <= a xor b;
    outputs(398) <= a xor b;
    outputs(399) <= not a or b;
    outputs(400) <= not a;
    outputs(401) <= a or b;
    outputs(402) <= b;
    outputs(403) <= a;
    outputs(404) <= not (a xor b);
    outputs(405) <= not (a xor b);
    outputs(406) <= not b;
    outputs(407) <= b;
    outputs(408) <= a and not b;
    outputs(409) <= not (a or b);
    outputs(410) <= not (a xor b);
    outputs(411) <= not (a and b);
    outputs(412) <= not b or a;
    outputs(413) <= a;
    outputs(414) <= a;
    outputs(415) <= not a;
    outputs(416) <= a and b;
    outputs(417) <= a and b;
    outputs(418) <= a xor b;
    outputs(419) <= a and not b;
    outputs(420) <= a xor b;
    outputs(421) <= b;
    outputs(422) <= b;
    outputs(423) <= not (a and b);
    outputs(424) <= not a;
    outputs(425) <= not a;
    outputs(426) <= a and b;
    outputs(427) <= a;
    outputs(428) <= not a;
    outputs(429) <= not (a or b);
    outputs(430) <= a;
    outputs(431) <= not b;
    outputs(432) <= b and not a;
    outputs(433) <= not (a xor b);
    outputs(434) <= not (a or b);
    outputs(435) <= not (a or b);
    outputs(436) <= a;
    outputs(437) <= a xor b;
    outputs(438) <= b and not a;
    outputs(439) <= a and not b;
    outputs(440) <= not a;
    outputs(441) <= not (a xor b);
    outputs(442) <= not (a or b);
    outputs(443) <= not (a or b);
    outputs(444) <= not b;
    outputs(445) <= a and b;
    outputs(446) <= a;
    outputs(447) <= a and b;
    outputs(448) <= a xor b;
    outputs(449) <= b;
    outputs(450) <= a and not b;
    outputs(451) <= b;
    outputs(452) <= not (a xor b);
    outputs(453) <= a and b;
    outputs(454) <= a or b;
    outputs(455) <= not b;
    outputs(456) <= a xor b;
    outputs(457) <= a and not b;
    outputs(458) <= not b;
    outputs(459) <= not b or a;
    outputs(460) <= not (a or b);
    outputs(461) <= not b;
    outputs(462) <= b and not a;
    outputs(463) <= a xor b;
    outputs(464) <= a;
    outputs(465) <= not b;
    outputs(466) <= a;
    outputs(467) <= a and b;
    outputs(468) <= a or b;
    outputs(469) <= a;
    outputs(470) <= a and b;
    outputs(471) <= not (a or b);
    outputs(472) <= not a;
    outputs(473) <= b;
    outputs(474) <= a xor b;
    outputs(475) <= not b;
    outputs(476) <= a and b;
    outputs(477) <= a and b;
    outputs(478) <= b;
    outputs(479) <= a and b;
    outputs(480) <= a;
    outputs(481) <= not a or b;
    outputs(482) <= a xor b;
    outputs(483) <= b;
    outputs(484) <= not a;
    outputs(485) <= not (a or b);
    outputs(486) <= not a;
    outputs(487) <= not a;
    outputs(488) <= not (a and b);
    outputs(489) <= not (a xor b);
    outputs(490) <= a xor b;
    outputs(491) <= not a or b;
    outputs(492) <= b;
    outputs(493) <= a;
    outputs(494) <= a xor b;
    outputs(495) <= not b;
    outputs(496) <= a and not b;
    outputs(497) <= a;
    outputs(498) <= a;
    outputs(499) <= a and b;
    outputs(500) <= b;
    outputs(501) <= a or b;
    outputs(502) <= not (a xor b);
    outputs(503) <= a xor b;
    outputs(504) <= not (a xor b);
    outputs(505) <= not (a xor b);
    outputs(506) <= not (a xor b);
    outputs(507) <= a;
    outputs(508) <= a xor b;
    outputs(509) <= not (a xor b);
    outputs(510) <= b;
    outputs(511) <= not b;
    outputs(512) <= a or b;
    outputs(513) <= not b;
    outputs(514) <= b and not a;
    outputs(515) <= not (a or b);
    outputs(516) <= a xor b;
    outputs(517) <= not (a and b);
    outputs(518) <= a;
    outputs(519) <= not b;
    outputs(520) <= not a or b;
    outputs(521) <= not a;
    outputs(522) <= a;
    outputs(523) <= not b or a;
    outputs(524) <= not (a or b);
    outputs(525) <= a xor b;
    outputs(526) <= not b or a;
    outputs(527) <= b;
    outputs(528) <= not a;
    outputs(529) <= not a;
    outputs(530) <= not b or a;
    outputs(531) <= not b;
    outputs(532) <= b and not a;
    outputs(533) <= a and not b;
    outputs(534) <= a or b;
    outputs(535) <= b;
    outputs(536) <= a;
    outputs(537) <= not a;
    outputs(538) <= not (a xor b);
    outputs(539) <= a and b;
    outputs(540) <= a;
    outputs(541) <= b and not a;
    outputs(542) <= a or b;
    outputs(543) <= not a;
    outputs(544) <= a;
    outputs(545) <= not (a or b);
    outputs(546) <= b;
    outputs(547) <= a and b;
    outputs(548) <= not a or b;
    outputs(549) <= b;
    outputs(550) <= not b;
    outputs(551) <= a;
    outputs(552) <= not b;
    outputs(553) <= b;
    outputs(554) <= not (a or b);
    outputs(555) <= not b;
    outputs(556) <= not (a or b);
    outputs(557) <= b;
    outputs(558) <= b;
    outputs(559) <= not a;
    outputs(560) <= not b;
    outputs(561) <= a xor b;
    outputs(562) <= a;
    outputs(563) <= a xor b;
    outputs(564) <= not a;
    outputs(565) <= a;
    outputs(566) <= not b or a;
    outputs(567) <= not a;
    outputs(568) <= not (a xor b);
    outputs(569) <= not a;
    outputs(570) <= not b;
    outputs(571) <= b;
    outputs(572) <= not (a xor b);
    outputs(573) <= not b;
    outputs(574) <= a or b;
    outputs(575) <= b and not a;
    outputs(576) <= a;
    outputs(577) <= not (a xor b);
    outputs(578) <= not a;
    outputs(579) <= b and not a;
    outputs(580) <= not b or a;
    outputs(581) <= a xor b;
    outputs(582) <= b;
    outputs(583) <= b and not a;
    outputs(584) <= not b;
    outputs(585) <= not (a or b);
    outputs(586) <= a and b;
    outputs(587) <= not a;
    outputs(588) <= b;
    outputs(589) <= b;
    outputs(590) <= a xor b;
    outputs(591) <= a;
    outputs(592) <= not b;
    outputs(593) <= not (a and b);
    outputs(594) <= not (a or b);
    outputs(595) <= not a;
    outputs(596) <= a xor b;
    outputs(597) <= not a;
    outputs(598) <= not b;
    outputs(599) <= not a;
    outputs(600) <= a;
    outputs(601) <= not b;
    outputs(602) <= a xor b;
    outputs(603) <= a xor b;
    outputs(604) <= not a;
    outputs(605) <= a and not b;
    outputs(606) <= not b or a;
    outputs(607) <= not (a and b);
    outputs(608) <= a xor b;
    outputs(609) <= b and not a;
    outputs(610) <= not (a or b);
    outputs(611) <= not (a or b);
    outputs(612) <= not (a xor b);
    outputs(613) <= b and not a;
    outputs(614) <= not b;
    outputs(615) <= a and not b;
    outputs(616) <= b and not a;
    outputs(617) <= a xor b;
    outputs(618) <= not a;
    outputs(619) <= a;
    outputs(620) <= a xor b;
    outputs(621) <= not b;
    outputs(622) <= not (a or b);
    outputs(623) <= not (a or b);
    outputs(624) <= not (a xor b);
    outputs(625) <= not b or a;
    outputs(626) <= a;
    outputs(627) <= a or b;
    outputs(628) <= not a;
    outputs(629) <= not (a or b);
    outputs(630) <= b;
    outputs(631) <= not b or a;
    outputs(632) <= a and not b;
    outputs(633) <= a and b;
    outputs(634) <= a xor b;
    outputs(635) <= b;
    outputs(636) <= a;
    outputs(637) <= not b;
    outputs(638) <= a xor b;
    outputs(639) <= not (a xor b);
    outputs(640) <= a;
    outputs(641) <= not b;
    outputs(642) <= not (a or b);
    outputs(643) <= a xor b;
    outputs(644) <= not (a xor b);
    outputs(645) <= not b;
    outputs(646) <= a;
    outputs(647) <= not b or a;
    outputs(648) <= b;
    outputs(649) <= not b;
    outputs(650) <= not a or b;
    outputs(651) <= not b;
    outputs(652) <= not (a xor b);
    outputs(653) <= b;
    outputs(654) <= a;
    outputs(655) <= not (a xor b);
    outputs(656) <= a;
    outputs(657) <= not a or b;
    outputs(658) <= a;
    outputs(659) <= not (a xor b);
    outputs(660) <= not b;
    outputs(661) <= b and not a;
    outputs(662) <= b;
    outputs(663) <= a;
    outputs(664) <= not (a and b);
    outputs(665) <= not (a and b);
    outputs(666) <= b and not a;
    outputs(667) <= not a;
    outputs(668) <= b;
    outputs(669) <= not b;
    outputs(670) <= not (a or b);
    outputs(671) <= b and not a;
    outputs(672) <= not (a xor b);
    outputs(673) <= a;
    outputs(674) <= not (a xor b);
    outputs(675) <= a;
    outputs(676) <= a and b;
    outputs(677) <= not b or a;
    outputs(678) <= not a or b;
    outputs(679) <= not b;
    outputs(680) <= a;
    outputs(681) <= a and not b;
    outputs(682) <= b;
    outputs(683) <= a xor b;
    outputs(684) <= a xor b;
    outputs(685) <= a and b;
    outputs(686) <= not a or b;
    outputs(687) <= not a;
    outputs(688) <= not b;
    outputs(689) <= not b;
    outputs(690) <= not (a and b);
    outputs(691) <= a xor b;
    outputs(692) <= not (a xor b);
    outputs(693) <= not b;
    outputs(694) <= a xor b;
    outputs(695) <= b;
    outputs(696) <= not a;
    outputs(697) <= a;
    outputs(698) <= not b or a;
    outputs(699) <= a;
    outputs(700) <= not (a xor b);
    outputs(701) <= not b;
    outputs(702) <= not (a xor b);
    outputs(703) <= b and not a;
    outputs(704) <= not b or a;
    outputs(705) <= not (a and b);
    outputs(706) <= a xor b;
    outputs(707) <= a xor b;
    outputs(708) <= not a or b;
    outputs(709) <= a and b;
    outputs(710) <= not b;
    outputs(711) <= not b;
    outputs(712) <= not (a xor b);
    outputs(713) <= b;
    outputs(714) <= a;
    outputs(715) <= a and b;
    outputs(716) <= not a;
    outputs(717) <= not b or a;
    outputs(718) <= b and not a;
    outputs(719) <= a;
    outputs(720) <= a and not b;
    outputs(721) <= not b;
    outputs(722) <= not b;
    outputs(723) <= not (a and b);
    outputs(724) <= b;
    outputs(725) <= not a or b;
    outputs(726) <= a xor b;
    outputs(727) <= a;
    outputs(728) <= not (a or b);
    outputs(729) <= not b or a;
    outputs(730) <= b and not a;
    outputs(731) <= b and not a;
    outputs(732) <= a and not b;
    outputs(733) <= a;
    outputs(734) <= b;
    outputs(735) <= not a;
    outputs(736) <= not (a xor b);
    outputs(737) <= not b;
    outputs(738) <= not a;
    outputs(739) <= a and b;
    outputs(740) <= not a;
    outputs(741) <= b and not a;
    outputs(742) <= b and not a;
    outputs(743) <= a;
    outputs(744) <= not b;
    outputs(745) <= not a;
    outputs(746) <= not a;
    outputs(747) <= b;
    outputs(748) <= not b;
    outputs(749) <= not b;
    outputs(750) <= not b;
    outputs(751) <= a xor b;
    outputs(752) <= a;
    outputs(753) <= a;
    outputs(754) <= not (a and b);
    outputs(755) <= not b;
    outputs(756) <= not (a and b);
    outputs(757) <= a and not b;
    outputs(758) <= not b or a;
    outputs(759) <= not a or b;
    outputs(760) <= a;
    outputs(761) <= a;
    outputs(762) <= a xor b;
    outputs(763) <= not b;
    outputs(764) <= not (a or b);
    outputs(765) <= not (a xor b);
    outputs(766) <= a and b;
    outputs(767) <= b;
    outputs(768) <= a and b;
    outputs(769) <= not a;
    outputs(770) <= a xor b;
    outputs(771) <= a xor b;
    outputs(772) <= b and not a;
    outputs(773) <= a;
    outputs(774) <= a xor b;
    outputs(775) <= not (a or b);
    outputs(776) <= not (a or b);
    outputs(777) <= a and not b;
    outputs(778) <= not (a xor b);
    outputs(779) <= a and b;
    outputs(780) <= b and not a;
    outputs(781) <= a;
    outputs(782) <= b and not a;
    outputs(783) <= a;
    outputs(784) <= not a;
    outputs(785) <= not a;
    outputs(786) <= b and not a;
    outputs(787) <= a and b;
    outputs(788) <= a xor b;
    outputs(789) <= a xor b;
    outputs(790) <= not (a xor b);
    outputs(791) <= b and not a;
    outputs(792) <= a and b;
    outputs(793) <= not (a or b);
    outputs(794) <= a;
    outputs(795) <= a and b;
    outputs(796) <= not (a and b);
    outputs(797) <= not a;
    outputs(798) <= not (a xor b);
    outputs(799) <= b and not a;
    outputs(800) <= b and not a;
    outputs(801) <= a and not b;
    outputs(802) <= b and not a;
    outputs(803) <= not a;
    outputs(804) <= b and not a;
    outputs(805) <= a;
    outputs(806) <= b;
    outputs(807) <= 1'b0;
    outputs(808) <= not (a or b);
    outputs(809) <= a xor b;
    outputs(810) <= not (a or b);
    outputs(811) <= a and not b;
    outputs(812) <= a and not b;
    outputs(813) <= b and not a;
    outputs(814) <= not (a xor b);
    outputs(815) <= b;
    outputs(816) <= a;
    outputs(817) <= not b;
    outputs(818) <= b and not a;
    outputs(819) <= not b;
    outputs(820) <= a;
    outputs(821) <= b and not a;
    outputs(822) <= b;
    outputs(823) <= a and not b;
    outputs(824) <= not (a or b);
    outputs(825) <= a xor b;
    outputs(826) <= not a;
    outputs(827) <= b and not a;
    outputs(828) <= a;
    outputs(829) <= 1'b0;
    outputs(830) <= not (a or b);
    outputs(831) <= not b;
    outputs(832) <= b and not a;
    outputs(833) <= b and not a;
    outputs(834) <= not (a xor b);
    outputs(835) <= not (a or b);
    outputs(836) <= a and b;
    outputs(837) <= b and not a;
    outputs(838) <= a and b;
    outputs(839) <= b and not a;
    outputs(840) <= b and not a;
    outputs(841) <= not (a or b);
    outputs(842) <= not (a or b);
    outputs(843) <= a and b;
    outputs(844) <= a and not b;
    outputs(845) <= 1'b0;
    outputs(846) <= a and not b;
    outputs(847) <= not (a xor b);
    outputs(848) <= not a;
    outputs(849) <= a and b;
    outputs(850) <= a and not b;
    outputs(851) <= a xor b;
    outputs(852) <= a xor b;
    outputs(853) <= not b or a;
    outputs(854) <= not a;
    outputs(855) <= a xor b;
    outputs(856) <= not (a and b);
    outputs(857) <= not b;
    outputs(858) <= not b;
    outputs(859) <= not b;
    outputs(860) <= b;
    outputs(861) <= a;
    outputs(862) <= not a;
    outputs(863) <= not a or b;
    outputs(864) <= a and not b;
    outputs(865) <= not (a or b);
    outputs(866) <= b;
    outputs(867) <= not (a or b);
    outputs(868) <= a and not b;
    outputs(869) <= a and not b;
    outputs(870) <= a and not b;
    outputs(871) <= not (a xor b);
    outputs(872) <= a and not b;
    outputs(873) <= b;
    outputs(874) <= b;
    outputs(875) <= b and not a;
    outputs(876) <= a and not b;
    outputs(877) <= not (a or b);
    outputs(878) <= a xor b;
    outputs(879) <= a;
    outputs(880) <= not a;
    outputs(881) <= a and not b;
    outputs(882) <= a xor b;
    outputs(883) <= not (a and b);
    outputs(884) <= not b;
    outputs(885) <= a xor b;
    outputs(886) <= not (a xor b);
    outputs(887) <= a and b;
    outputs(888) <= not (a or b);
    outputs(889) <= a and b;
    outputs(890) <= a xor b;
    outputs(891) <= b and not a;
    outputs(892) <= a and not b;
    outputs(893) <= not (a xor b);
    outputs(894) <= not b;
    outputs(895) <= not (a xor b);
    outputs(896) <= not (a xor b);
    outputs(897) <= 1'b0;
    outputs(898) <= not a;
    outputs(899) <= a and b;
    outputs(900) <= a and b;
    outputs(901) <= not (a xor b);
    outputs(902) <= not (a xor b);
    outputs(903) <= not b;
    outputs(904) <= not b;
    outputs(905) <= not (a or b);
    outputs(906) <= b;
    outputs(907) <= a and b;
    outputs(908) <= not (a or b);
    outputs(909) <= a and not b;
    outputs(910) <= 1'b0;
    outputs(911) <= a xor b;
    outputs(912) <= a and b;
    outputs(913) <= not (a or b);
    outputs(914) <= a and b;
    outputs(915) <= not (a or b);
    outputs(916) <= a and not b;
    outputs(917) <= b;
    outputs(918) <= a and not b;
    outputs(919) <= not (a or b);
    outputs(920) <= b and not a;
    outputs(921) <= a and b;
    outputs(922) <= b;
    outputs(923) <= b;
    outputs(924) <= not (a or b);
    outputs(925) <= a and b;
    outputs(926) <= not (a xor b);
    outputs(927) <= not a;
    outputs(928) <= not (a or b);
    outputs(929) <= b and not a;
    outputs(930) <= not b;
    outputs(931) <= a and not b;
    outputs(932) <= b and not a;
    outputs(933) <= b and not a;
    outputs(934) <= a xor b;
    outputs(935) <= a xor b;
    outputs(936) <= b;
    outputs(937) <= b and not a;
    outputs(938) <= a and not b;
    outputs(939) <= not (a or b);
    outputs(940) <= b and not a;
    outputs(941) <= a and not b;
    outputs(942) <= a and not b;
    outputs(943) <= not a or b;
    outputs(944) <= a xor b;
    outputs(945) <= not b;
    outputs(946) <= b and not a;
    outputs(947) <= a and not b;
    outputs(948) <= not (a or b);
    outputs(949) <= a and not b;
    outputs(950) <= b and not a;
    outputs(951) <= b and not a;
    outputs(952) <= b;
    outputs(953) <= b and not a;
    outputs(954) <= a;
    outputs(955) <= b;
    outputs(956) <= not (a or b);
    outputs(957) <= a and b;
    outputs(958) <= not b;
    outputs(959) <= b and not a;
    outputs(960) <= not b;
    outputs(961) <= a xor b;
    outputs(962) <= b and not a;
    outputs(963) <= not (a or b);
    outputs(964) <= a and not b;
    outputs(965) <= a;
    outputs(966) <= not (a xor b);
    outputs(967) <= not a;
    outputs(968) <= not a;
    outputs(969) <= a;
    outputs(970) <= not (a or b);
    outputs(971) <= not (a or b);
    outputs(972) <= b and not a;
    outputs(973) <= a xor b;
    outputs(974) <= b;
    outputs(975) <= not a;
    outputs(976) <= a and not b;
    outputs(977) <= a xor b;
    outputs(978) <= a and b;
    outputs(979) <= not b or a;
    outputs(980) <= a and not b;
    outputs(981) <= not a;
    outputs(982) <= a and not b;
    outputs(983) <= a and not b;
    outputs(984) <= a xor b;
    outputs(985) <= not (a or b);
    outputs(986) <= not (a xor b);
    outputs(987) <= not b;
    outputs(988) <= a;
    outputs(989) <= a xor b;
    outputs(990) <= a and b;
    outputs(991) <= a xor b;
    outputs(992) <= a and not b;
    outputs(993) <= a and not b;
    outputs(994) <= a xor b;
    outputs(995) <= 1'b0;
    outputs(996) <= a and not b;
    outputs(997) <= not (a or b);
    outputs(998) <= b and not a;
    outputs(999) <= b and not a;
    outputs(1000) <= b and not a;
    outputs(1001) <= not (a or b);
    outputs(1002) <= a and not b;
    outputs(1003) <= a and b;
    outputs(1004) <= not (a xor b);
    outputs(1005) <= not (a xor b);
    outputs(1006) <= a and b;
    outputs(1007) <= not (a or b);
    outputs(1008) <= b;
    outputs(1009) <= a and b;
    outputs(1010) <= a and not b;
    outputs(1011) <= not a;
    outputs(1012) <= not (a or b);
    outputs(1013) <= b and not a;
    outputs(1014) <= b and not a;
    outputs(1015) <= a and b;
    outputs(1016) <= not b;
    outputs(1017) <= b and not a;
    outputs(1018) <= not (a xor b);
    outputs(1019) <= a;
    outputs(1020) <= a and b;
    outputs(1021) <= a and not b;
    outputs(1022) <= a xor b;
    outputs(1023) <= b and not a;
    outputs(1024) <= not a;
    outputs(1025) <= a and not b;
    outputs(1026) <= b and not a;
    outputs(1027) <= not b;
    outputs(1028) <= not b;
    outputs(1029) <= a xor b;
    outputs(1030) <= not (a or b);
    outputs(1031) <= not (a or b);
    outputs(1032) <= not (a xor b);
    outputs(1033) <= b;
    outputs(1034) <= not (a xor b);
    outputs(1035) <= not (a or b);
    outputs(1036) <= not (a xor b);
    outputs(1037) <= a;
    outputs(1038) <= b and not a;
    outputs(1039) <= not (a xor b);
    outputs(1040) <= b and not a;
    outputs(1041) <= a xor b;
    outputs(1042) <= b and not a;
    outputs(1043) <= a and not b;
    outputs(1044) <= b and not a;
    outputs(1045) <= b;
    outputs(1046) <= not (a or b);
    outputs(1047) <= a and not b;
    outputs(1048) <= b and not a;
    outputs(1049) <= a;
    outputs(1050) <= a and not b;
    outputs(1051) <= a and not b;
    outputs(1052) <= not b;
    outputs(1053) <= a and not b;
    outputs(1054) <= a and not b;
    outputs(1055) <= a and not b;
    outputs(1056) <= b and not a;
    outputs(1057) <= a;
    outputs(1058) <= a and not b;
    outputs(1059) <= b and not a;
    outputs(1060) <= a and b;
    outputs(1061) <= b and not a;
    outputs(1062) <= not a;
    outputs(1063) <= not b;
    outputs(1064) <= not b;
    outputs(1065) <= a and not b;
    outputs(1066) <= not (a or b);
    outputs(1067) <= a xor b;
    outputs(1068) <= not b;
    outputs(1069) <= b;
    outputs(1070) <= not (a xor b);
    outputs(1071) <= a xor b;
    outputs(1072) <= a and b;
    outputs(1073) <= b and not a;
    outputs(1074) <= not (a or b);
    outputs(1075) <= not a;
    outputs(1076) <= a and b;
    outputs(1077) <= a xor b;
    outputs(1078) <= not a;
    outputs(1079) <= b;
    outputs(1080) <= b and not a;
    outputs(1081) <= a and b;
    outputs(1082) <= b and not a;
    outputs(1083) <= not (a or b);
    outputs(1084) <= b and not a;
    outputs(1085) <= a and b;
    outputs(1086) <= a and b;
    outputs(1087) <= a;
    outputs(1088) <= b and not a;
    outputs(1089) <= a and b;
    outputs(1090) <= a;
    outputs(1091) <= b;
    outputs(1092) <= a and b;
    outputs(1093) <= a;
    outputs(1094) <= a;
    outputs(1095) <= b;
    outputs(1096) <= not (a or b);
    outputs(1097) <= not b;
    outputs(1098) <= b;
    outputs(1099) <= not (a or b);
    outputs(1100) <= a and b;
    outputs(1101) <= not (a xor b);
    outputs(1102) <= a xor b;
    outputs(1103) <= not (a xor b);
    outputs(1104) <= not b;
    outputs(1105) <= not (a xor b);
    outputs(1106) <= not b;
    outputs(1107) <= a and b;
    outputs(1108) <= a and b;
    outputs(1109) <= a and not b;
    outputs(1110) <= not a or b;
    outputs(1111) <= a and not b;
    outputs(1112) <= a and b;
    outputs(1113) <= a xor b;
    outputs(1114) <= not (a xor b);
    outputs(1115) <= a and not b;
    outputs(1116) <= b and not a;
    outputs(1117) <= a and b;
    outputs(1118) <= a and not b;
    outputs(1119) <= b and not a;
    outputs(1120) <= b and not a;
    outputs(1121) <= a and b;
    outputs(1122) <= not (a xor b);
    outputs(1123) <= b;
    outputs(1124) <= not (a or b);
    outputs(1125) <= a;
    outputs(1126) <= a and b;
    outputs(1127) <= b and not a;
    outputs(1128) <= b and not a;
    outputs(1129) <= a;
    outputs(1130) <= b;
    outputs(1131) <= not b;
    outputs(1132) <= a and not b;
    outputs(1133) <= not b or a;
    outputs(1134) <= not (a or b);
    outputs(1135) <= not b;
    outputs(1136) <= not b;
    outputs(1137) <= a and not b;
    outputs(1138) <= a and b;
    outputs(1139) <= not (a or b);
    outputs(1140) <= not b;
    outputs(1141) <= a;
    outputs(1142) <= a and not b;
    outputs(1143) <= not (a xor b);
    outputs(1144) <= not (a xor b);
    outputs(1145) <= not a;
    outputs(1146) <= a and b;
    outputs(1147) <= a xor b;
    outputs(1148) <= not (a or b);
    outputs(1149) <= a and b;
    outputs(1150) <= not (a or b);
    outputs(1151) <= a and b;
    outputs(1152) <= not a;
    outputs(1153) <= not (a xor b);
    outputs(1154) <= a xor b;
    outputs(1155) <= a xor b;
    outputs(1156) <= not a;
    outputs(1157) <= a and not b;
    outputs(1158) <= a xor b;
    outputs(1159) <= a and b;
    outputs(1160) <= not a;
    outputs(1161) <= a and not b;
    outputs(1162) <= not a;
    outputs(1163) <= b;
    outputs(1164) <= a and not b;
    outputs(1165) <= a and not b;
    outputs(1166) <= a;
    outputs(1167) <= not (a or b);
    outputs(1168) <= a xor b;
    outputs(1169) <= not (a or b);
    outputs(1170) <= b and not a;
    outputs(1171) <= not (a xor b);
    outputs(1172) <= a and not b;
    outputs(1173) <= not (a xor b);
    outputs(1174) <= not b;
    outputs(1175) <= not (a or b);
    outputs(1176) <= not b or a;
    outputs(1177) <= b and not a;
    outputs(1178) <= a xor b;
    outputs(1179) <= a xor b;
    outputs(1180) <= not a;
    outputs(1181) <= a and b;
    outputs(1182) <= not (a xor b);
    outputs(1183) <= a and b;
    outputs(1184) <= b;
    outputs(1185) <= a xor b;
    outputs(1186) <= a and not b;
    outputs(1187) <= not a or b;
    outputs(1188) <= b and not a;
    outputs(1189) <= a and not b;
    outputs(1190) <= a;
    outputs(1191) <= b;
    outputs(1192) <= not (a or b);
    outputs(1193) <= a;
    outputs(1194) <= not (a xor b);
    outputs(1195) <= not (a or b);
    outputs(1196) <= b and not a;
    outputs(1197) <= a and not b;
    outputs(1198) <= not (a or b);
    outputs(1199) <= b and not a;
    outputs(1200) <= a xor b;
    outputs(1201) <= not (a and b);
    outputs(1202) <= not (a or b);
    outputs(1203) <= a and not b;
    outputs(1204) <= not b or a;
    outputs(1205) <= a and b;
    outputs(1206) <= b;
    outputs(1207) <= a and b;
    outputs(1208) <= not (a or b);
    outputs(1209) <= a;
    outputs(1210) <= a and not b;
    outputs(1211) <= not (a or b);
    outputs(1212) <= a and b;
    outputs(1213) <= not a or b;
    outputs(1214) <= not b;
    outputs(1215) <= a;
    outputs(1216) <= a;
    outputs(1217) <= a and b;
    outputs(1218) <= not (a xor b);
    outputs(1219) <= not (a xor b);
    outputs(1220) <= a and not b;
    outputs(1221) <= not (a xor b);
    outputs(1222) <= a and b;
    outputs(1223) <= a and b;
    outputs(1224) <= a;
    outputs(1225) <= b and not a;
    outputs(1226) <= not (a or b);
    outputs(1227) <= b and not a;
    outputs(1228) <= a and b;
    outputs(1229) <= a and not b;
    outputs(1230) <= b;
    outputs(1231) <= b and not a;
    outputs(1232) <= a xor b;
    outputs(1233) <= a and not b;
    outputs(1234) <= a and b;
    outputs(1235) <= b and not a;
    outputs(1236) <= not (a xor b);
    outputs(1237) <= not b;
    outputs(1238) <= a xor b;
    outputs(1239) <= a and not b;
    outputs(1240) <= not a;
    outputs(1241) <= not (a or b);
    outputs(1242) <= a and not b;
    outputs(1243) <= a;
    outputs(1244) <= not (a or b);
    outputs(1245) <= a;
    outputs(1246) <= a xor b;
    outputs(1247) <= 1'b0;
    outputs(1248) <= not (a or b);
    outputs(1249) <= b;
    outputs(1250) <= b and not a;
    outputs(1251) <= not (a or b);
    outputs(1252) <= not (a xor b);
    outputs(1253) <= b and not a;
    outputs(1254) <= a xor b;
    outputs(1255) <= a xor b;
    outputs(1256) <= not b;
    outputs(1257) <= a and b;
    outputs(1258) <= a and b;
    outputs(1259) <= not b;
    outputs(1260) <= b;
    outputs(1261) <= not a;
    outputs(1262) <= a and b;
    outputs(1263) <= b;
    outputs(1264) <= not a;
    outputs(1265) <= a and not b;
    outputs(1266) <= b and not a;
    outputs(1267) <= b and not a;
    outputs(1268) <= not (a xor b);
    outputs(1269) <= a and not b;
    outputs(1270) <= b and not a;
    outputs(1271) <= a xor b;
    outputs(1272) <= a;
    outputs(1273) <= b and not a;
    outputs(1274) <= b and not a;
    outputs(1275) <= not a;
    outputs(1276) <= not b;
    outputs(1277) <= a and b;
    outputs(1278) <= not (a or b);
    outputs(1279) <= not b;
    outputs(1280) <= a and b;
    outputs(1281) <= a xor b;
    outputs(1282) <= a and not b;
    outputs(1283) <= a and b;
    outputs(1284) <= a xor b;
    outputs(1285) <= a;
    outputs(1286) <= a and b;
    outputs(1287) <= not b;
    outputs(1288) <= a xor b;
    outputs(1289) <= not (a xor b);
    outputs(1290) <= b;
    outputs(1291) <= a and b;
    outputs(1292) <= not (a xor b);
    outputs(1293) <= a;
    outputs(1294) <= not b;
    outputs(1295) <= not (a or b);
    outputs(1296) <= a xor b;
    outputs(1297) <= not (a xor b);
    outputs(1298) <= a and b;
    outputs(1299) <= b and not a;
    outputs(1300) <= a xor b;
    outputs(1301) <= a xor b;
    outputs(1302) <= b and not a;
    outputs(1303) <= a and not b;
    outputs(1304) <= not (a or b);
    outputs(1305) <= a and not b;
    outputs(1306) <= not a;
    outputs(1307) <= a and b;
    outputs(1308) <= a xor b;
    outputs(1309) <= not a;
    outputs(1310) <= not (a xor b);
    outputs(1311) <= not (a or b);
    outputs(1312) <= not (a or b);
    outputs(1313) <= not a;
    outputs(1314) <= b;
    outputs(1315) <= not (a or b);
    outputs(1316) <= not b;
    outputs(1317) <= a xor b;
    outputs(1318) <= not (a xor b);
    outputs(1319) <= not b;
    outputs(1320) <= not b;
    outputs(1321) <= a;
    outputs(1322) <= not a;
    outputs(1323) <= b;
    outputs(1324) <= not a or b;
    outputs(1325) <= not (a xor b);
    outputs(1326) <= a and b;
    outputs(1327) <= a and not b;
    outputs(1328) <= b and not a;
    outputs(1329) <= not (a or b);
    outputs(1330) <= a xor b;
    outputs(1331) <= not a;
    outputs(1332) <= not a;
    outputs(1333) <= b and not a;
    outputs(1334) <= a xor b;
    outputs(1335) <= a;
    outputs(1336) <= a xor b;
    outputs(1337) <= not (a xor b);
    outputs(1338) <= not (a or b);
    outputs(1339) <= not a;
    outputs(1340) <= b;
    outputs(1341) <= a and b;
    outputs(1342) <= a and b;
    outputs(1343) <= a;
    outputs(1344) <= b;
    outputs(1345) <= not (a or b);
    outputs(1346) <= a and not b;
    outputs(1347) <= a;
    outputs(1348) <= not a or b;
    outputs(1349) <= a and b;
    outputs(1350) <= a xor b;
    outputs(1351) <= a and not b;
    outputs(1352) <= not (a or b);
    outputs(1353) <= not (a xor b);
    outputs(1354) <= not (a or b);
    outputs(1355) <= a and b;
    outputs(1356) <= a and b;
    outputs(1357) <= not b;
    outputs(1358) <= not (a xor b);
    outputs(1359) <= a and not b;
    outputs(1360) <= a and not b;
    outputs(1361) <= a and not b;
    outputs(1362) <= not a;
    outputs(1363) <= b and not a;
    outputs(1364) <= not (a xor b);
    outputs(1365) <= b and not a;
    outputs(1366) <= b and not a;
    outputs(1367) <= not (a or b);
    outputs(1368) <= b;
    outputs(1369) <= b and not a;
    outputs(1370) <= b;
    outputs(1371) <= b;
    outputs(1372) <= not (a or b);
    outputs(1373) <= not a;
    outputs(1374) <= not a;
    outputs(1375) <= not a;
    outputs(1376) <= a and not b;
    outputs(1377) <= not b;
    outputs(1378) <= 1'b0;
    outputs(1379) <= a and not b;
    outputs(1380) <= not (a or b);
    outputs(1381) <= a and b;
    outputs(1382) <= not b or a;
    outputs(1383) <= not (a xor b);
    outputs(1384) <= a and b;
    outputs(1385) <= a and not b;
    outputs(1386) <= a xor b;
    outputs(1387) <= a and b;
    outputs(1388) <= a and not b;
    outputs(1389) <= a xor b;
    outputs(1390) <= a and b;
    outputs(1391) <= a and b;
    outputs(1392) <= not a;
    outputs(1393) <= a;
    outputs(1394) <= a and not b;
    outputs(1395) <= b and not a;
    outputs(1396) <= a and b;
    outputs(1397) <= a and not b;
    outputs(1398) <= a and b;
    outputs(1399) <= b;
    outputs(1400) <= not (a or b);
    outputs(1401) <= a xor b;
    outputs(1402) <= not b;
    outputs(1403) <= b;
    outputs(1404) <= 1'b0;
    outputs(1405) <= b and not a;
    outputs(1406) <= b;
    outputs(1407) <= b and not a;
    outputs(1408) <= a and not b;
    outputs(1409) <= a and b;
    outputs(1410) <= a xor b;
    outputs(1411) <= a and not b;
    outputs(1412) <= a xor b;
    outputs(1413) <= a xor b;
    outputs(1414) <= b;
    outputs(1415) <= not a;
    outputs(1416) <= not (a xor b);
    outputs(1417) <= not a;
    outputs(1418) <= a and b;
    outputs(1419) <= a and b;
    outputs(1420) <= a and b;
    outputs(1421) <= a and not b;
    outputs(1422) <= b and not a;
    outputs(1423) <= not (a xor b);
    outputs(1424) <= b;
    outputs(1425) <= b and not a;
    outputs(1426) <= not b;
    outputs(1427) <= b and not a;
    outputs(1428) <= b and not a;
    outputs(1429) <= not (a xor b);
    outputs(1430) <= a and b;
    outputs(1431) <= a xor b;
    outputs(1432) <= a and not b;
    outputs(1433) <= a xor b;
    outputs(1434) <= b and not a;
    outputs(1435) <= a and b;
    outputs(1436) <= not (a or b);
    outputs(1437) <= not (a or b);
    outputs(1438) <= a and b;
    outputs(1439) <= not b;
    outputs(1440) <= not (a or b);
    outputs(1441) <= a and not b;
    outputs(1442) <= a and not b;
    outputs(1443) <= not (a or b);
    outputs(1444) <= a and b;
    outputs(1445) <= b;
    outputs(1446) <= not (a or b);
    outputs(1447) <= not b;
    outputs(1448) <= a and not b;
    outputs(1449) <= a and not b;
    outputs(1450) <= not a;
    outputs(1451) <= not (a or b);
    outputs(1452) <= not (a or b);
    outputs(1453) <= a xor b;
    outputs(1454) <= a and not b;
    outputs(1455) <= a and b;
    outputs(1456) <= not b;
    outputs(1457) <= b;
    outputs(1458) <= not (a xor b);
    outputs(1459) <= not (a xor b);
    outputs(1460) <= a;
    outputs(1461) <= b and not a;
    outputs(1462) <= not a;
    outputs(1463) <= not (a or b);
    outputs(1464) <= b and not a;
    outputs(1465) <= a and not b;
    outputs(1466) <= not b;
    outputs(1467) <= a;
    outputs(1468) <= a and not b;
    outputs(1469) <= a;
    outputs(1470) <= b;
    outputs(1471) <= a xor b;
    outputs(1472) <= b and not a;
    outputs(1473) <= not b;
    outputs(1474) <= not (a or b);
    outputs(1475) <= a and b;
    outputs(1476) <= a and not b;
    outputs(1477) <= a and b;
    outputs(1478) <= a xor b;
    outputs(1479) <= a xor b;
    outputs(1480) <= not (a or b);
    outputs(1481) <= a;
    outputs(1482) <= a;
    outputs(1483) <= b and not a;
    outputs(1484) <= b and not a;
    outputs(1485) <= a and not b;
    outputs(1486) <= a and b;
    outputs(1487) <= a xor b;
    outputs(1488) <= a and not b;
    outputs(1489) <= a and not b;
    outputs(1490) <= a and not b;
    outputs(1491) <= a and not b;
    outputs(1492) <= 1'b0;
    outputs(1493) <= a and not b;
    outputs(1494) <= a and b;
    outputs(1495) <= not (a or b);
    outputs(1496) <= a and not b;
    outputs(1497) <= a and b;
    outputs(1498) <= a and not b;
    outputs(1499) <= not (a xor b);
    outputs(1500) <= b and not a;
    outputs(1501) <= a and not b;
    outputs(1502) <= a and not b;
    outputs(1503) <= b;
    outputs(1504) <= b and not a;
    outputs(1505) <= a and not b;
    outputs(1506) <= not b;
    outputs(1507) <= not (a xor b);
    outputs(1508) <= not (a or b);
    outputs(1509) <= not (a xor b);
    outputs(1510) <= not (a or b);
    outputs(1511) <= b;
    outputs(1512) <= not b;
    outputs(1513) <= not (a or b);
    outputs(1514) <= a and b;
    outputs(1515) <= a xor b;
    outputs(1516) <= not (a xor b);
    outputs(1517) <= not a or b;
    outputs(1518) <= a xor b;
    outputs(1519) <= not a or b;
    outputs(1520) <= b and not a;
    outputs(1521) <= b;
    outputs(1522) <= not (a or b);
    outputs(1523) <= b and not a;
    outputs(1524) <= not (a xor b);
    outputs(1525) <= a and b;
    outputs(1526) <= a and b;
    outputs(1527) <= a xor b;
    outputs(1528) <= a;
    outputs(1529) <= not a;
    outputs(1530) <= not a;
    outputs(1531) <= a;
    outputs(1532) <= b and not a;
    outputs(1533) <= not b;
    outputs(1534) <= not (a or b);
    outputs(1535) <= not a;
    outputs(1536) <= not (a and b);
    outputs(1537) <= not a;
    outputs(1538) <= not b or a;
    outputs(1539) <= not a;
    outputs(1540) <= not b;
    outputs(1541) <= not (a or b);
    outputs(1542) <= b;
    outputs(1543) <= b;
    outputs(1544) <= a xor b;
    outputs(1545) <= not b;
    outputs(1546) <= b;
    outputs(1547) <= a;
    outputs(1548) <= not (a or b);
    outputs(1549) <= b;
    outputs(1550) <= b;
    outputs(1551) <= not a;
    outputs(1552) <= a and b;
    outputs(1553) <= not b or a;
    outputs(1554) <= a xor b;
    outputs(1555) <= b and not a;
    outputs(1556) <= a and not b;
    outputs(1557) <= not a;
    outputs(1558) <= not (a or b);
    outputs(1559) <= a xor b;
    outputs(1560) <= a xor b;
    outputs(1561) <= a and b;
    outputs(1562) <= not b;
    outputs(1563) <= a or b;
    outputs(1564) <= b and not a;
    outputs(1565) <= b and not a;
    outputs(1566) <= b and not a;
    outputs(1567) <= not a;
    outputs(1568) <= a;
    outputs(1569) <= a or b;
    outputs(1570) <= not (a xor b);
    outputs(1571) <= not a;
    outputs(1572) <= a and not b;
    outputs(1573) <= not b;
    outputs(1574) <= a;
    outputs(1575) <= a and b;
    outputs(1576) <= not (a xor b);
    outputs(1577) <= a;
    outputs(1578) <= not (a xor b);
    outputs(1579) <= b;
    outputs(1580) <= a or b;
    outputs(1581) <= b;
    outputs(1582) <= not b;
    outputs(1583) <= b;
    outputs(1584) <= a or b;
    outputs(1585) <= a xor b;
    outputs(1586) <= a;
    outputs(1587) <= a and not b;
    outputs(1588) <= b and not a;
    outputs(1589) <= a xor b;
    outputs(1590) <= not (a or b);
    outputs(1591) <= a and not b;
    outputs(1592) <= a or b;
    outputs(1593) <= not (a and b);
    outputs(1594) <= not b;
    outputs(1595) <= not (a and b);
    outputs(1596) <= not a or b;
    outputs(1597) <= not (a or b);
    outputs(1598) <= b;
    outputs(1599) <= b;
    outputs(1600) <= not a or b;
    outputs(1601) <= a xor b;
    outputs(1602) <= not (a xor b);
    outputs(1603) <= not b or a;
    outputs(1604) <= b;
    outputs(1605) <= not a or b;
    outputs(1606) <= b;
    outputs(1607) <= not b or a;
    outputs(1608) <= a xor b;
    outputs(1609) <= a and not b;
    outputs(1610) <= not a;
    outputs(1611) <= a xor b;
    outputs(1612) <= not (a and b);
    outputs(1613) <= not (a xor b);
    outputs(1614) <= a;
    outputs(1615) <= a;
    outputs(1616) <= a or b;
    outputs(1617) <= a and b;
    outputs(1618) <= b;
    outputs(1619) <= not a;
    outputs(1620) <= not (a xor b);
    outputs(1621) <= a;
    outputs(1622) <= b and not a;
    outputs(1623) <= a;
    outputs(1624) <= not b;
    outputs(1625) <= not a;
    outputs(1626) <= a and b;
    outputs(1627) <= not (a xor b);
    outputs(1628) <= a and not b;
    outputs(1629) <= not (a and b);
    outputs(1630) <= not a;
    outputs(1631) <= not (a or b);
    outputs(1632) <= a;
    outputs(1633) <= not (a xor b);
    outputs(1634) <= not a;
    outputs(1635) <= not b;
    outputs(1636) <= not b;
    outputs(1637) <= b;
    outputs(1638) <= not b;
    outputs(1639) <= not b or a;
    outputs(1640) <= a xor b;
    outputs(1641) <= a xor b;
    outputs(1642) <= not a;
    outputs(1643) <= not a;
    outputs(1644) <= not a;
    outputs(1645) <= not (a xor b);
    outputs(1646) <= b;
    outputs(1647) <= b;
    outputs(1648) <= not (a xor b);
    outputs(1649) <= a xor b;
    outputs(1650) <= not (a xor b);
    outputs(1651) <= not a;
    outputs(1652) <= a;
    outputs(1653) <= not b;
    outputs(1654) <= a;
    outputs(1655) <= not (a xor b);
    outputs(1656) <= not (a xor b);
    outputs(1657) <= a;
    outputs(1658) <= not (a xor b);
    outputs(1659) <= not (a or b);
    outputs(1660) <= not b;
    outputs(1661) <= b;
    outputs(1662) <= a;
    outputs(1663) <= b and not a;
    outputs(1664) <= not (a xor b);
    outputs(1665) <= not a;
    outputs(1666) <= not a;
    outputs(1667) <= a or b;
    outputs(1668) <= not b;
    outputs(1669) <= a xor b;
    outputs(1670) <= a xor b;
    outputs(1671) <= b;
    outputs(1672) <= a or b;
    outputs(1673) <= a or b;
    outputs(1674) <= b and not a;
    outputs(1675) <= not b or a;
    outputs(1676) <= a xor b;
    outputs(1677) <= a;
    outputs(1678) <= not (a or b);
    outputs(1679) <= not b;
    outputs(1680) <= a;
    outputs(1681) <= not b;
    outputs(1682) <= not (a and b);
    outputs(1683) <= a;
    outputs(1684) <= not b or a;
    outputs(1685) <= b and not a;
    outputs(1686) <= a or b;
    outputs(1687) <= not (a and b);
    outputs(1688) <= b and not a;
    outputs(1689) <= not a or b;
    outputs(1690) <= b and not a;
    outputs(1691) <= not b;
    outputs(1692) <= b;
    outputs(1693) <= b and not a;
    outputs(1694) <= not b;
    outputs(1695) <= not (a or b);
    outputs(1696) <= a and not b;
    outputs(1697) <= a;
    outputs(1698) <= not (a xor b);
    outputs(1699) <= not (a xor b);
    outputs(1700) <= b;
    outputs(1701) <= a and not b;
    outputs(1702) <= a;
    outputs(1703) <= not (a and b);
    outputs(1704) <= a xor b;
    outputs(1705) <= b;
    outputs(1706) <= a;
    outputs(1707) <= not (a and b);
    outputs(1708) <= b;
    outputs(1709) <= b;
    outputs(1710) <= a and not b;
    outputs(1711) <= not a;
    outputs(1712) <= not a;
    outputs(1713) <= a;
    outputs(1714) <= not a;
    outputs(1715) <= b;
    outputs(1716) <= not (a and b);
    outputs(1717) <= not a;
    outputs(1718) <= not (a xor b);
    outputs(1719) <= not (a or b);
    outputs(1720) <= a or b;
    outputs(1721) <= not b;
    outputs(1722) <= a and not b;
    outputs(1723) <= a or b;
    outputs(1724) <= not (a xor b);
    outputs(1725) <= not b;
    outputs(1726) <= b;
    outputs(1727) <= b and not a;
    outputs(1728) <= not (a xor b);
    outputs(1729) <= a and b;
    outputs(1730) <= not b;
    outputs(1731) <= not a;
    outputs(1732) <= not a;
    outputs(1733) <= a or b;
    outputs(1734) <= b;
    outputs(1735) <= a or b;
    outputs(1736) <= a xor b;
    outputs(1737) <= a xor b;
    outputs(1738) <= a or b;
    outputs(1739) <= a and b;
    outputs(1740) <= not (a or b);
    outputs(1741) <= a;
    outputs(1742) <= b;
    outputs(1743) <= not (a and b);
    outputs(1744) <= a xor b;
    outputs(1745) <= not a or b;
    outputs(1746) <= not a;
    outputs(1747) <= not a;
    outputs(1748) <= not (a or b);
    outputs(1749) <= a xor b;
    outputs(1750) <= b;
    outputs(1751) <= not b;
    outputs(1752) <= a;
    outputs(1753) <= not a;
    outputs(1754) <= not b;
    outputs(1755) <= not (a xor b);
    outputs(1756) <= not a;
    outputs(1757) <= a xor b;
    outputs(1758) <= a and b;
    outputs(1759) <= not a or b;
    outputs(1760) <= b;
    outputs(1761) <= a and not b;
    outputs(1762) <= a or b;
    outputs(1763) <= not (a xor b);
    outputs(1764) <= a xor b;
    outputs(1765) <= a;
    outputs(1766) <= not (a xor b);
    outputs(1767) <= b;
    outputs(1768) <= a;
    outputs(1769) <= b;
    outputs(1770) <= not (a xor b);
    outputs(1771) <= not a;
    outputs(1772) <= a and b;
    outputs(1773) <= not a;
    outputs(1774) <= not a;
    outputs(1775) <= not b;
    outputs(1776) <= b and not a;
    outputs(1777) <= b and not a;
    outputs(1778) <= a xor b;
    outputs(1779) <= b;
    outputs(1780) <= a and not b;
    outputs(1781) <= not b;
    outputs(1782) <= not b;
    outputs(1783) <= not a or b;
    outputs(1784) <= not a;
    outputs(1785) <= b and not a;
    outputs(1786) <= a or b;
    outputs(1787) <= not (a or b);
    outputs(1788) <= not (a xor b);
    outputs(1789) <= not b;
    outputs(1790) <= not b;
    outputs(1791) <= not b;
    outputs(1792) <= a;
    outputs(1793) <= a and not b;
    outputs(1794) <= not a;
    outputs(1795) <= a or b;
    outputs(1796) <= b;
    outputs(1797) <= a xor b;
    outputs(1798) <= not (a and b);
    outputs(1799) <= a and b;
    outputs(1800) <= not (a or b);
    outputs(1801) <= not (a xor b);
    outputs(1802) <= b;
    outputs(1803) <= a and not b;
    outputs(1804) <= not (a and b);
    outputs(1805) <= not (a xor b);
    outputs(1806) <= a xor b;
    outputs(1807) <= not (a xor b);
    outputs(1808) <= a and b;
    outputs(1809) <= a and not b;
    outputs(1810) <= not (a or b);
    outputs(1811) <= not b or a;
    outputs(1812) <= a;
    outputs(1813) <= not a or b;
    outputs(1814) <= not b;
    outputs(1815) <= b;
    outputs(1816) <= b and not a;
    outputs(1817) <= a;
    outputs(1818) <= not a or b;
    outputs(1819) <= b;
    outputs(1820) <= not b;
    outputs(1821) <= a xor b;
    outputs(1822) <= a and not b;
    outputs(1823) <= not a;
    outputs(1824) <= a;
    outputs(1825) <= b and not a;
    outputs(1826) <= b;
    outputs(1827) <= not a or b;
    outputs(1828) <= a and b;
    outputs(1829) <= not (a xor b);
    outputs(1830) <= a and b;
    outputs(1831) <= not b or a;
    outputs(1832) <= not b;
    outputs(1833) <= not (a xor b);
    outputs(1834) <= a xor b;
    outputs(1835) <= not (a xor b);
    outputs(1836) <= a or b;
    outputs(1837) <= a;
    outputs(1838) <= not (a xor b);
    outputs(1839) <= b;
    outputs(1840) <= a and not b;
    outputs(1841) <= not (a xor b);
    outputs(1842) <= a;
    outputs(1843) <= not a;
    outputs(1844) <= a;
    outputs(1845) <= not (a or b);
    outputs(1846) <= a and b;
    outputs(1847) <= a;
    outputs(1848) <= b;
    outputs(1849) <= b;
    outputs(1850) <= not a;
    outputs(1851) <= a or b;
    outputs(1852) <= a or b;
    outputs(1853) <= b and not a;
    outputs(1854) <= a;
    outputs(1855) <= not (a or b);
    outputs(1856) <= not b or a;
    outputs(1857) <= not b;
    outputs(1858) <= a xor b;
    outputs(1859) <= not (a xor b);
    outputs(1860) <= a;
    outputs(1861) <= a xor b;
    outputs(1862) <= not a or b;
    outputs(1863) <= not b or a;
    outputs(1864) <= not (a and b);
    outputs(1865) <= a and b;
    outputs(1866) <= a;
    outputs(1867) <= not a;
    outputs(1868) <= not b or a;
    outputs(1869) <= b;
    outputs(1870) <= a;
    outputs(1871) <= a xor b;
    outputs(1872) <= a xor b;
    outputs(1873) <= not (a or b);
    outputs(1874) <= not b or a;
    outputs(1875) <= b and not a;
    outputs(1876) <= not b;
    outputs(1877) <= not a or b;
    outputs(1878) <= not (a xor b);
    outputs(1879) <= a and not b;
    outputs(1880) <= a;
    outputs(1881) <= a xor b;
    outputs(1882) <= b;
    outputs(1883) <= not (a and b);
    outputs(1884) <= a xor b;
    outputs(1885) <= a;
    outputs(1886) <= b and not a;
    outputs(1887) <= not (a xor b);
    outputs(1888) <= not b or a;
    outputs(1889) <= not (a or b);
    outputs(1890) <= not a or b;
    outputs(1891) <= not a or b;
    outputs(1892) <= b;
    outputs(1893) <= a;
    outputs(1894) <= a or b;
    outputs(1895) <= not a;
    outputs(1896) <= not a or b;
    outputs(1897) <= a and not b;
    outputs(1898) <= not (a and b);
    outputs(1899) <= not a;
    outputs(1900) <= a xor b;
    outputs(1901) <= not a or b;
    outputs(1902) <= not b;
    outputs(1903) <= b and not a;
    outputs(1904) <= b;
    outputs(1905) <= not (a and b);
    outputs(1906) <= not (a or b);
    outputs(1907) <= not (a and b);
    outputs(1908) <= b;
    outputs(1909) <= a or b;
    outputs(1910) <= a;
    outputs(1911) <= b;
    outputs(1912) <= a xor b;
    outputs(1913) <= not b;
    outputs(1914) <= a;
    outputs(1915) <= not (a xor b);
    outputs(1916) <= a xor b;
    outputs(1917) <= a;
    outputs(1918) <= a and not b;
    outputs(1919) <= a and b;
    outputs(1920) <= not (a or b);
    outputs(1921) <= a xor b;
    outputs(1922) <= not b;
    outputs(1923) <= a xor b;
    outputs(1924) <= a;
    outputs(1925) <= a and not b;
    outputs(1926) <= not b;
    outputs(1927) <= not (a or b);
    outputs(1928) <= not a;
    outputs(1929) <= a;
    outputs(1930) <= not a;
    outputs(1931) <= not a;
    outputs(1932) <= a xor b;
    outputs(1933) <= a xor b;
    outputs(1934) <= a xor b;
    outputs(1935) <= not a or b;
    outputs(1936) <= not b;
    outputs(1937) <= a or b;
    outputs(1938) <= not (a and b);
    outputs(1939) <= not b;
    outputs(1940) <= a or b;
    outputs(1941) <= b;
    outputs(1942) <= not a or b;
    outputs(1943) <= b;
    outputs(1944) <= a;
    outputs(1945) <= not (a xor b);
    outputs(1946) <= b and not a;
    outputs(1947) <= not (a and b);
    outputs(1948) <= b;
    outputs(1949) <= not a;
    outputs(1950) <= not b;
    outputs(1951) <= b and not a;
    outputs(1952) <= a;
    outputs(1953) <= a xor b;
    outputs(1954) <= a xor b;
    outputs(1955) <= not b;
    outputs(1956) <= not (a or b);
    outputs(1957) <= not (a or b);
    outputs(1958) <= a and b;
    outputs(1959) <= a and b;
    outputs(1960) <= b;
    outputs(1961) <= not a or b;
    outputs(1962) <= a xor b;
    outputs(1963) <= not a;
    outputs(1964) <= not (a xor b);
    outputs(1965) <= a and b;
    outputs(1966) <= not b;
    outputs(1967) <= not a;
    outputs(1968) <= not a;
    outputs(1969) <= a and b;
    outputs(1970) <= not (a or b);
    outputs(1971) <= not a;
    outputs(1972) <= not b;
    outputs(1973) <= not a or b;
    outputs(1974) <= b;
    outputs(1975) <= a and b;
    outputs(1976) <= a or b;
    outputs(1977) <= not a or b;
    outputs(1978) <= not (a xor b);
    outputs(1979) <= not a or b;
    outputs(1980) <= b and not a;
    outputs(1981) <= b and not a;
    outputs(1982) <= b;
    outputs(1983) <= a or b;
    outputs(1984) <= b;
    outputs(1985) <= not a;
    outputs(1986) <= b and not a;
    outputs(1987) <= not b;
    outputs(1988) <= a and b;
    outputs(1989) <= a and b;
    outputs(1990) <= a;
    outputs(1991) <= b;
    outputs(1992) <= not b;
    outputs(1993) <= not b;
    outputs(1994) <= not b or a;
    outputs(1995) <= a xor b;
    outputs(1996) <= not b or a;
    outputs(1997) <= b and not a;
    outputs(1998) <= not a;
    outputs(1999) <= b;
    outputs(2000) <= a;
    outputs(2001) <= not (a xor b);
    outputs(2002) <= a;
    outputs(2003) <= not b or a;
    outputs(2004) <= a;
    outputs(2005) <= a;
    outputs(2006) <= not (a xor b);
    outputs(2007) <= a;
    outputs(2008) <= a and b;
    outputs(2009) <= not a or b;
    outputs(2010) <= not a;
    outputs(2011) <= not (a and b);
    outputs(2012) <= not (a xor b);
    outputs(2013) <= not (a xor b);
    outputs(2014) <= not b;
    outputs(2015) <= not (a and b);
    outputs(2016) <= a;
    outputs(2017) <= a;
    outputs(2018) <= not b;
    outputs(2019) <= not (a or b);
    outputs(2020) <= a and not b;
    outputs(2021) <= a or b;
    outputs(2022) <= b;
    outputs(2023) <= b;
    outputs(2024) <= not b;
    outputs(2025) <= not (a or b);
    outputs(2026) <= not (a xor b);
    outputs(2027) <= a or b;
    outputs(2028) <= not a or b;
    outputs(2029) <= not (a and b);
    outputs(2030) <= not a;
    outputs(2031) <= b;
    outputs(2032) <= not (a xor b);
    outputs(2033) <= a;
    outputs(2034) <= b and not a;
    outputs(2035) <= a xor b;
    outputs(2036) <= not a;
    outputs(2037) <= a xor b;
    outputs(2038) <= not b;
    outputs(2039) <= a xor b;
    outputs(2040) <= not a;
    outputs(2041) <= a;
    outputs(2042) <= not b or a;
    outputs(2043) <= not a;
    outputs(2044) <= a xor b;
    outputs(2045) <= a;
    outputs(2046) <= a;
    outputs(2047) <= a or b;
    outputs(2048) <= not a;
    outputs(2049) <= not a or b;
    outputs(2050) <= a and not b;
    outputs(2051) <= not b or a;
    outputs(2052) <= not a or b;
    outputs(2053) <= not a;
    outputs(2054) <= a xor b;
    outputs(2055) <= not (a and b);
    outputs(2056) <= not a;
    outputs(2057) <= b;
    outputs(2058) <= a xor b;
    outputs(2059) <= not b;
    outputs(2060) <= not b;
    outputs(2061) <= not (a or b);
    outputs(2062) <= not (a xor b);
    outputs(2063) <= b and not a;
    outputs(2064) <= not b;
    outputs(2065) <= a;
    outputs(2066) <= not (a xor b);
    outputs(2067) <= not (a or b);
    outputs(2068) <= a xor b;
    outputs(2069) <= b;
    outputs(2070) <= b;
    outputs(2071) <= a xor b;
    outputs(2072) <= not b or a;
    outputs(2073) <= b;
    outputs(2074) <= not b;
    outputs(2075) <= not (a xor b);
    outputs(2076) <= a;
    outputs(2077) <= a xor b;
    outputs(2078) <= not a;
    outputs(2079) <= a;
    outputs(2080) <= not b or a;
    outputs(2081) <= not b;
    outputs(2082) <= not (a xor b);
    outputs(2083) <= not a;
    outputs(2084) <= not a or b;
    outputs(2085) <= not a;
    outputs(2086) <= not b or a;
    outputs(2087) <= a or b;
    outputs(2088) <= a and not b;
    outputs(2089) <= not (a or b);
    outputs(2090) <= a;
    outputs(2091) <= not b or a;
    outputs(2092) <= not b;
    outputs(2093) <= not (a xor b);
    outputs(2094) <= a xor b;
    outputs(2095) <= a xor b;
    outputs(2096) <= not a;
    outputs(2097) <= not (a xor b);
    outputs(2098) <= not b;
    outputs(2099) <= not b;
    outputs(2100) <= a xor b;
    outputs(2101) <= not (a or b);
    outputs(2102) <= a and not b;
    outputs(2103) <= a and not b;
    outputs(2104) <= not (a and b);
    outputs(2105) <= not b;
    outputs(2106) <= b and not a;
    outputs(2107) <= a xor b;
    outputs(2108) <= a or b;
    outputs(2109) <= not a;
    outputs(2110) <= not (a xor b);
    outputs(2111) <= b;
    outputs(2112) <= not (a xor b);
    outputs(2113) <= not a;
    outputs(2114) <= not b;
    outputs(2115) <= not (a or b);
    outputs(2116) <= not (a or b);
    outputs(2117) <= b;
    outputs(2118) <= b;
    outputs(2119) <= a and not b;
    outputs(2120) <= not b;
    outputs(2121) <= a;
    outputs(2122) <= a xor b;
    outputs(2123) <= b;
    outputs(2124) <= not (a xor b);
    outputs(2125) <= not a;
    outputs(2126) <= not a or b;
    outputs(2127) <= not (a xor b);
    outputs(2128) <= not (a xor b);
    outputs(2129) <= a xor b;
    outputs(2130) <= a xor b;
    outputs(2131) <= a;
    outputs(2132) <= a;
    outputs(2133) <= not (a and b);
    outputs(2134) <= not a or b;
    outputs(2135) <= not (a xor b);
    outputs(2136) <= a xor b;
    outputs(2137) <= b and not a;
    outputs(2138) <= not (a and b);
    outputs(2139) <= a;
    outputs(2140) <= not b or a;
    outputs(2141) <= not b;
    outputs(2142) <= a and b;
    outputs(2143) <= a or b;
    outputs(2144) <= a;
    outputs(2145) <= not b or a;
    outputs(2146) <= a;
    outputs(2147) <= not b;
    outputs(2148) <= a and b;
    outputs(2149) <= a;
    outputs(2150) <= a or b;
    outputs(2151) <= not (a xor b);
    outputs(2152) <= not (a xor b);
    outputs(2153) <= not (a and b);
    outputs(2154) <= a or b;
    outputs(2155) <= not b or a;
    outputs(2156) <= a xor b;
    outputs(2157) <= a and b;
    outputs(2158) <= not (a xor b);
    outputs(2159) <= b;
    outputs(2160) <= a or b;
    outputs(2161) <= a xor b;
    outputs(2162) <= not b or a;
    outputs(2163) <= a and not b;
    outputs(2164) <= not (a and b);
    outputs(2165) <= a xor b;
    outputs(2166) <= not (a xor b);
    outputs(2167) <= not (a and b);
    outputs(2168) <= a or b;
    outputs(2169) <= not (a xor b);
    outputs(2170) <= not (a xor b);
    outputs(2171) <= not a or b;
    outputs(2172) <= a;
    outputs(2173) <= b;
    outputs(2174) <= not (a xor b);
    outputs(2175) <= not a or b;
    outputs(2176) <= not b;
    outputs(2177) <= not b;
    outputs(2178) <= a xor b;
    outputs(2179) <= b and not a;
    outputs(2180) <= a xor b;
    outputs(2181) <= a or b;
    outputs(2182) <= not a;
    outputs(2183) <= not (a and b);
    outputs(2184) <= a;
    outputs(2185) <= a or b;
    outputs(2186) <= a or b;
    outputs(2187) <= not b;
    outputs(2188) <= not a;
    outputs(2189) <= not b or a;
    outputs(2190) <= not b or a;
    outputs(2191) <= not (a xor b);
    outputs(2192) <= b;
    outputs(2193) <= a and b;
    outputs(2194) <= a;
    outputs(2195) <= a;
    outputs(2196) <= not (a or b);
    outputs(2197) <= a and b;
    outputs(2198) <= not (a xor b);
    outputs(2199) <= not a;
    outputs(2200) <= not b;
    outputs(2201) <= b and not a;
    outputs(2202) <= not a;
    outputs(2203) <= not b;
    outputs(2204) <= a and b;
    outputs(2205) <= a;
    outputs(2206) <= not (a xor b);
    outputs(2207) <= not b;
    outputs(2208) <= not a;
    outputs(2209) <= not b or a;
    outputs(2210) <= b;
    outputs(2211) <= not a or b;
    outputs(2212) <= b;
    outputs(2213) <= not b;
    outputs(2214) <= a;
    outputs(2215) <= a;
    outputs(2216) <= a and b;
    outputs(2217) <= b;
    outputs(2218) <= not b;
    outputs(2219) <= not a or b;
    outputs(2220) <= a;
    outputs(2221) <= a or b;
    outputs(2222) <= not b or a;
    outputs(2223) <= a xor b;
    outputs(2224) <= not (a xor b);
    outputs(2225) <= not (a and b);
    outputs(2226) <= a and not b;
    outputs(2227) <= a;
    outputs(2228) <= not (a and b);
    outputs(2229) <= not (a xor b);
    outputs(2230) <= not (a xor b);
    outputs(2231) <= a;
    outputs(2232) <= not (a xor b);
    outputs(2233) <= b;
    outputs(2234) <= not a;
    outputs(2235) <= a;
    outputs(2236) <= not b or a;
    outputs(2237) <= a xor b;
    outputs(2238) <= a xor b;
    outputs(2239) <= a or b;
    outputs(2240) <= not b;
    outputs(2241) <= a;
    outputs(2242) <= a and b;
    outputs(2243) <= not a or b;
    outputs(2244) <= b and not a;
    outputs(2245) <= a;
    outputs(2246) <= not (a or b);
    outputs(2247) <= not (a and b);
    outputs(2248) <= a;
    outputs(2249) <= not a;
    outputs(2250) <= a;
    outputs(2251) <= b;
    outputs(2252) <= a xor b;
    outputs(2253) <= a xor b;
    outputs(2254) <= a;
    outputs(2255) <= a;
    outputs(2256) <= not (a or b);
    outputs(2257) <= a and b;
    outputs(2258) <= a xor b;
    outputs(2259) <= a or b;
    outputs(2260) <= a xor b;
    outputs(2261) <= a xor b;
    outputs(2262) <= not a;
    outputs(2263) <= a or b;
    outputs(2264) <= not b or a;
    outputs(2265) <= a;
    outputs(2266) <= a xor b;
    outputs(2267) <= not b or a;
    outputs(2268) <= b and not a;
    outputs(2269) <= a xor b;
    outputs(2270) <= b;
    outputs(2271) <= not a;
    outputs(2272) <= not a;
    outputs(2273) <= b;
    outputs(2274) <= not (a or b);
    outputs(2275) <= b;
    outputs(2276) <= b;
    outputs(2277) <= not a;
    outputs(2278) <= b;
    outputs(2279) <= not (a or b);
    outputs(2280) <= not (a and b);
    outputs(2281) <= a;
    outputs(2282) <= not b;
    outputs(2283) <= a;
    outputs(2284) <= a and b;
    outputs(2285) <= not (a xor b);
    outputs(2286) <= a xor b;
    outputs(2287) <= b;
    outputs(2288) <= a;
    outputs(2289) <= not a;
    outputs(2290) <= not a;
    outputs(2291) <= b;
    outputs(2292) <= a or b;
    outputs(2293) <= a;
    outputs(2294) <= a and b;
    outputs(2295) <= b;
    outputs(2296) <= a;
    outputs(2297) <= a and b;
    outputs(2298) <= a xor b;
    outputs(2299) <= not (a xor b);
    outputs(2300) <= a;
    outputs(2301) <= a or b;
    outputs(2302) <= b and not a;
    outputs(2303) <= b;
    outputs(2304) <= not (a or b);
    outputs(2305) <= a or b;
    outputs(2306) <= b and not a;
    outputs(2307) <= a and not b;
    outputs(2308) <= not (a or b);
    outputs(2309) <= not b or a;
    outputs(2310) <= a;
    outputs(2311) <= not a;
    outputs(2312) <= b;
    outputs(2313) <= a and b;
    outputs(2314) <= a;
    outputs(2315) <= a;
    outputs(2316) <= not (a or b);
    outputs(2317) <= not b;
    outputs(2318) <= a and not b;
    outputs(2319) <= a or b;
    outputs(2320) <= not (a xor b);
    outputs(2321) <= a or b;
    outputs(2322) <= a;
    outputs(2323) <= not a or b;
    outputs(2324) <= not (a xor b);
    outputs(2325) <= b;
    outputs(2326) <= not (a xor b);
    outputs(2327) <= a or b;
    outputs(2328) <= not a;
    outputs(2329) <= a and not b;
    outputs(2330) <= b;
    outputs(2331) <= not (a xor b);
    outputs(2332) <= a;
    outputs(2333) <= b and not a;
    outputs(2334) <= a or b;
    outputs(2335) <= not b;
    outputs(2336) <= not (a xor b);
    outputs(2337) <= not b;
    outputs(2338) <= not a or b;
    outputs(2339) <= a xor b;
    outputs(2340) <= not b;
    outputs(2341) <= not (a or b);
    outputs(2342) <= not (a and b);
    outputs(2343) <= b;
    outputs(2344) <= a xor b;
    outputs(2345) <= not (a or b);
    outputs(2346) <= a and not b;
    outputs(2347) <= a or b;
    outputs(2348) <= not (a xor b);
    outputs(2349) <= not a;
    outputs(2350) <= b;
    outputs(2351) <= not (a or b);
    outputs(2352) <= not (a and b);
    outputs(2353) <= not (a xor b);
    outputs(2354) <= a;
    outputs(2355) <= not (a xor b);
    outputs(2356) <= a;
    outputs(2357) <= not a or b;
    outputs(2358) <= not a;
    outputs(2359) <= a and b;
    outputs(2360) <= not a;
    outputs(2361) <= b;
    outputs(2362) <= not b;
    outputs(2363) <= not a;
    outputs(2364) <= not a;
    outputs(2365) <= a xor b;
    outputs(2366) <= not (a and b);
    outputs(2367) <= a;
    outputs(2368) <= not b or a;
    outputs(2369) <= b and not a;
    outputs(2370) <= not b;
    outputs(2371) <= a;
    outputs(2372) <= a or b;
    outputs(2373) <= a and b;
    outputs(2374) <= not b;
    outputs(2375) <= not b;
    outputs(2376) <= not (a and b);
    outputs(2377) <= not (a xor b);
    outputs(2378) <= not (a and b);
    outputs(2379) <= a or b;
    outputs(2380) <= not (a xor b);
    outputs(2381) <= not b or a;
    outputs(2382) <= not b;
    outputs(2383) <= not a;
    outputs(2384) <= not (a and b);
    outputs(2385) <= not (a xor b);
    outputs(2386) <= not a;
    outputs(2387) <= b;
    outputs(2388) <= not b;
    outputs(2389) <= a and b;
    outputs(2390) <= a xor b;
    outputs(2391) <= not a;
    outputs(2392) <= not a;
    outputs(2393) <= a or b;
    outputs(2394) <= not (a or b);
    outputs(2395) <= b and not a;
    outputs(2396) <= a xor b;
    outputs(2397) <= not b or a;
    outputs(2398) <= not b;
    outputs(2399) <= b and not a;
    outputs(2400) <= not a or b;
    outputs(2401) <= not a;
    outputs(2402) <= not (a or b);
    outputs(2403) <= not b or a;
    outputs(2404) <= not b;
    outputs(2405) <= a xor b;
    outputs(2406) <= not a;
    outputs(2407) <= b;
    outputs(2408) <= a and b;
    outputs(2409) <= not (a and b);
    outputs(2410) <= not b;
    outputs(2411) <= a;
    outputs(2412) <= a;
    outputs(2413) <= b;
    outputs(2414) <= not (a xor b);
    outputs(2415) <= not (a or b);
    outputs(2416) <= b;
    outputs(2417) <= not a;
    outputs(2418) <= not (a xor b);
    outputs(2419) <= a and not b;
    outputs(2420) <= a;
    outputs(2421) <= not a;
    outputs(2422) <= a and b;
    outputs(2423) <= not a;
    outputs(2424) <= b;
    outputs(2425) <= not a;
    outputs(2426) <= a and not b;
    outputs(2427) <= a xor b;
    outputs(2428) <= not a;
    outputs(2429) <= not b or a;
    outputs(2430) <= a and not b;
    outputs(2431) <= not (a or b);
    outputs(2432) <= not (a xor b);
    outputs(2433) <= a xor b;
    outputs(2434) <= not a;
    outputs(2435) <= not (a xor b);
    outputs(2436) <= not (a or b);
    outputs(2437) <= a;
    outputs(2438) <= a;
    outputs(2439) <= not (a xor b);
    outputs(2440) <= a xor b;
    outputs(2441) <= not (a xor b);
    outputs(2442) <= not (a and b);
    outputs(2443) <= not a;
    outputs(2444) <= b;
    outputs(2445) <= b;
    outputs(2446) <= not b or a;
    outputs(2447) <= a and not b;
    outputs(2448) <= not b or a;
    outputs(2449) <= not b or a;
    outputs(2450) <= b;
    outputs(2451) <= not (a or b);
    outputs(2452) <= a and not b;
    outputs(2453) <= not a;
    outputs(2454) <= a;
    outputs(2455) <= not b;
    outputs(2456) <= a;
    outputs(2457) <= b and not a;
    outputs(2458) <= not a or b;
    outputs(2459) <= not a or b;
    outputs(2460) <= b and not a;
    outputs(2461) <= not (a xor b);
    outputs(2462) <= a xor b;
    outputs(2463) <= a or b;
    outputs(2464) <= a and not b;
    outputs(2465) <= a;
    outputs(2466) <= not a or b;
    outputs(2467) <= b and not a;
    outputs(2468) <= a xor b;
    outputs(2469) <= b;
    outputs(2470) <= b;
    outputs(2471) <= b and not a;
    outputs(2472) <= not (a or b);
    outputs(2473) <= not a;
    outputs(2474) <= not (a xor b);
    outputs(2475) <= b;
    outputs(2476) <= a;
    outputs(2477) <= a;
    outputs(2478) <= b;
    outputs(2479) <= not (a xor b);
    outputs(2480) <= a;
    outputs(2481) <= not b;
    outputs(2482) <= a;
    outputs(2483) <= a xor b;
    outputs(2484) <= a xor b;
    outputs(2485) <= not a;
    outputs(2486) <= not a or b;
    outputs(2487) <= not (a or b);
    outputs(2488) <= a xor b;
    outputs(2489) <= not (a xor b);
    outputs(2490) <= a xor b;
    outputs(2491) <= not b or a;
    outputs(2492) <= not b or a;
    outputs(2493) <= not (a xor b);
    outputs(2494) <= not b;
    outputs(2495) <= not b;
    outputs(2496) <= not b;
    outputs(2497) <= not (a xor b);
    outputs(2498) <= not b or a;
    outputs(2499) <= not (a and b);
    outputs(2500) <= not b;
    outputs(2501) <= a;
    outputs(2502) <= not (a xor b);
    outputs(2503) <= not (a and b);
    outputs(2504) <= b;
    outputs(2505) <= b;
    outputs(2506) <= not (a xor b);
    outputs(2507) <= a;
    outputs(2508) <= not b;
    outputs(2509) <= not (a xor b);
    outputs(2510) <= a;
    outputs(2511) <= a;
    outputs(2512) <= a and b;
    outputs(2513) <= a;
    outputs(2514) <= a;
    outputs(2515) <= not (a xor b);
    outputs(2516) <= a;
    outputs(2517) <= a and not b;
    outputs(2518) <= a and b;
    outputs(2519) <= b;
    outputs(2520) <= not b;
    outputs(2521) <= not a;
    outputs(2522) <= b;
    outputs(2523) <= a;
    outputs(2524) <= not b or a;
    outputs(2525) <= a and b;
    outputs(2526) <= a;
    outputs(2527) <= a;
    outputs(2528) <= not b or a;
    outputs(2529) <= not (a or b);
    outputs(2530) <= not b or a;
    outputs(2531) <= a and b;
    outputs(2532) <= not (a xor b);
    outputs(2533) <= a;
    outputs(2534) <= not (a xor b);
    outputs(2535) <= not (a xor b);
    outputs(2536) <= a;
    outputs(2537) <= b;
    outputs(2538) <= not (a xor b);
    outputs(2539) <= not b;
    outputs(2540) <= a and b;
    outputs(2541) <= b;
    outputs(2542) <= a;
    outputs(2543) <= a xor b;
    outputs(2544) <= b and not a;
    outputs(2545) <= a xor b;
    outputs(2546) <= not (a and b);
    outputs(2547) <= a or b;
    outputs(2548) <= a;
    outputs(2549) <= not (a xor b);
    outputs(2550) <= not (a xor b);
    outputs(2551) <= a;
    outputs(2552) <= b;
    outputs(2553) <= not a;
    outputs(2554) <= a xor b;
    outputs(2555) <= a;
    outputs(2556) <= a xor b;
    outputs(2557) <= not a;
    outputs(2558) <= not a;
    outputs(2559) <= not a or b;
    outputs(2560) <= a and not b;
    outputs(2561) <= not (a xor b);
    outputs(2562) <= a xor b;
    outputs(2563) <= not (a or b);
    outputs(2564) <= b;
    outputs(2565) <= a;
    outputs(2566) <= not (a xor b);
    outputs(2567) <= not (a xor b);
    outputs(2568) <= not b or a;
    outputs(2569) <= not a or b;
    outputs(2570) <= b;
    outputs(2571) <= not a;
    outputs(2572) <= not (a xor b);
    outputs(2573) <= a xor b;
    outputs(2574) <= not (a xor b);
    outputs(2575) <= not (a and b);
    outputs(2576) <= a xor b;
    outputs(2577) <= b;
    outputs(2578) <= b;
    outputs(2579) <= a;
    outputs(2580) <= not b;
    outputs(2581) <= not (a xor b);
    outputs(2582) <= not (a xor b);
    outputs(2583) <= not (a or b);
    outputs(2584) <= not (a xor b);
    outputs(2585) <= a;
    outputs(2586) <= not a or b;
    outputs(2587) <= a;
    outputs(2588) <= b;
    outputs(2589) <= not b;
    outputs(2590) <= a;
    outputs(2591) <= not (a or b);
    outputs(2592) <= a or b;
    outputs(2593) <= not b or a;
    outputs(2594) <= b and not a;
    outputs(2595) <= not (a xor b);
    outputs(2596) <= not b;
    outputs(2597) <= not (a xor b);
    outputs(2598) <= a or b;
    outputs(2599) <= a xor b;
    outputs(2600) <= not (a and b);
    outputs(2601) <= not a;
    outputs(2602) <= a and b;
    outputs(2603) <= a;
    outputs(2604) <= a and b;
    outputs(2605) <= a and not b;
    outputs(2606) <= b;
    outputs(2607) <= a and b;
    outputs(2608) <= not (a and b);
    outputs(2609) <= not (a xor b);
    outputs(2610) <= not a or b;
    outputs(2611) <= b and not a;
    outputs(2612) <= not (a xor b);
    outputs(2613) <= b;
    outputs(2614) <= a;
    outputs(2615) <= not a;
    outputs(2616) <= b;
    outputs(2617) <= not (a or b);
    outputs(2618) <= a xor b;
    outputs(2619) <= a and not b;
    outputs(2620) <= a;
    outputs(2621) <= not b;
    outputs(2622) <= not a;
    outputs(2623) <= a;
    outputs(2624) <= not b;
    outputs(2625) <= not b;
    outputs(2626) <= b;
    outputs(2627) <= not (a or b);
    outputs(2628) <= a and not b;
    outputs(2629) <= not b;
    outputs(2630) <= not b;
    outputs(2631) <= not (a xor b);
    outputs(2632) <= a and not b;
    outputs(2633) <= not a;
    outputs(2634) <= b;
    outputs(2635) <= not b;
    outputs(2636) <= not a;
    outputs(2637) <= a;
    outputs(2638) <= a;
    outputs(2639) <= b and not a;
    outputs(2640) <= not b;
    outputs(2641) <= not (a xor b);
    outputs(2642) <= a or b;
    outputs(2643) <= not (a and b);
    outputs(2644) <= b;
    outputs(2645) <= a xor b;
    outputs(2646) <= not b or a;
    outputs(2647) <= b;
    outputs(2648) <= not a;
    outputs(2649) <= b;
    outputs(2650) <= not a;
    outputs(2651) <= a;
    outputs(2652) <= not b;
    outputs(2653) <= b;
    outputs(2654) <= not a;
    outputs(2655) <= not (a xor b);
    outputs(2656) <= not a;
    outputs(2657) <= not a;
    outputs(2658) <= not a;
    outputs(2659) <= not a;
    outputs(2660) <= a and b;
    outputs(2661) <= not b or a;
    outputs(2662) <= b;
    outputs(2663) <= a xor b;
    outputs(2664) <= not (a or b);
    outputs(2665) <= not b;
    outputs(2666) <= a and not b;
    outputs(2667) <= b and not a;
    outputs(2668) <= not a or b;
    outputs(2669) <= not a;
    outputs(2670) <= b and not a;
    outputs(2671) <= a xor b;
    outputs(2672) <= not a;
    outputs(2673) <= a and b;
    outputs(2674) <= not (a xor b);
    outputs(2675) <= not b;
    outputs(2676) <= not (a xor b);
    outputs(2677) <= b;
    outputs(2678) <= not (a xor b);
    outputs(2679) <= not a;
    outputs(2680) <= not (a xor b);
    outputs(2681) <= not a;
    outputs(2682) <= b;
    outputs(2683) <= not b;
    outputs(2684) <= a or b;
    outputs(2685) <= b;
    outputs(2686) <= a;
    outputs(2687) <= not (a xor b);
    outputs(2688) <= not a;
    outputs(2689) <= a;
    outputs(2690) <= a and not b;
    outputs(2691) <= a;
    outputs(2692) <= a and not b;
    outputs(2693) <= b;
    outputs(2694) <= b;
    outputs(2695) <= not a;
    outputs(2696) <= a xor b;
    outputs(2697) <= b;
    outputs(2698) <= a;
    outputs(2699) <= b;
    outputs(2700) <= b and not a;
    outputs(2701) <= not (a xor b);
    outputs(2702) <= b;
    outputs(2703) <= not a or b;
    outputs(2704) <= not a;
    outputs(2705) <= a and not b;
    outputs(2706) <= not a;
    outputs(2707) <= a xor b;
    outputs(2708) <= not b;
    outputs(2709) <= not (a xor b);
    outputs(2710) <= b;
    outputs(2711) <= not (a xor b);
    outputs(2712) <= b and not a;
    outputs(2713) <= not a;
    outputs(2714) <= b;
    outputs(2715) <= a and b;
    outputs(2716) <= a and not b;
    outputs(2717) <= b;
    outputs(2718) <= not a;
    outputs(2719) <= not (a xor b);
    outputs(2720) <= b;
    outputs(2721) <= a xor b;
    outputs(2722) <= a and b;
    outputs(2723) <= b;
    outputs(2724) <= not (a xor b);
    outputs(2725) <= not a;
    outputs(2726) <= not b;
    outputs(2727) <= not (a and b);
    outputs(2728) <= not (a or b);
    outputs(2729) <= a;
    outputs(2730) <= a and b;
    outputs(2731) <= not a;
    outputs(2732) <= not b or a;
    outputs(2733) <= b;
    outputs(2734) <= not a;
    outputs(2735) <= a xor b;
    outputs(2736) <= not a;
    outputs(2737) <= a xor b;
    outputs(2738) <= b and not a;
    outputs(2739) <= b and not a;
    outputs(2740) <= not b;
    outputs(2741) <= a or b;
    outputs(2742) <= not (a and b);
    outputs(2743) <= not (a xor b);
    outputs(2744) <= a xor b;
    outputs(2745) <= not a;
    outputs(2746) <= b and not a;
    outputs(2747) <= a xor b;
    outputs(2748) <= a xor b;
    outputs(2749) <= not a;
    outputs(2750) <= a xor b;
    outputs(2751) <= b and not a;
    outputs(2752) <= b;
    outputs(2753) <= a xor b;
    outputs(2754) <= not a;
    outputs(2755) <= b and not a;
    outputs(2756) <= a;
    outputs(2757) <= a xor b;
    outputs(2758) <= a;
    outputs(2759) <= a xor b;
    outputs(2760) <= not (a xor b);
    outputs(2761) <= b and not a;
    outputs(2762) <= a xor b;
    outputs(2763) <= not b;
    outputs(2764) <= a;
    outputs(2765) <= not (a xor b);
    outputs(2766) <= a xor b;
    outputs(2767) <= a xor b;
    outputs(2768) <= not (a xor b);
    outputs(2769) <= a xor b;
    outputs(2770) <= a and b;
    outputs(2771) <= b;
    outputs(2772) <= not (a xor b);
    outputs(2773) <= not b or a;
    outputs(2774) <= a xor b;
    outputs(2775) <= not a;
    outputs(2776) <= not b;
    outputs(2777) <= not a;
    outputs(2778) <= not (a xor b);
    outputs(2779) <= not b;
    outputs(2780) <= not a;
    outputs(2781) <= not b;
    outputs(2782) <= not (a xor b);
    outputs(2783) <= not a;
    outputs(2784) <= not (a and b);
    outputs(2785) <= not a;
    outputs(2786) <= a and not b;
    outputs(2787) <= not (a xor b);
    outputs(2788) <= b and not a;
    outputs(2789) <= not (a xor b);
    outputs(2790) <= not b;
    outputs(2791) <= not b;
    outputs(2792) <= a or b;
    outputs(2793) <= not (a xor b);
    outputs(2794) <= not (a xor b);
    outputs(2795) <= a;
    outputs(2796) <= a;
    outputs(2797) <= not b;
    outputs(2798) <= not (a xor b);
    outputs(2799) <= not (a and b);
    outputs(2800) <= not (a or b);
    outputs(2801) <= not b or a;
    outputs(2802) <= not a;
    outputs(2803) <= not b;
    outputs(2804) <= not (a and b);
    outputs(2805) <= b;
    outputs(2806) <= a and b;
    outputs(2807) <= not b;
    outputs(2808) <= a or b;
    outputs(2809) <= not (a and b);
    outputs(2810) <= b;
    outputs(2811) <= a;
    outputs(2812) <= a and not b;
    outputs(2813) <= not a;
    outputs(2814) <= a and b;
    outputs(2815) <= not a;
    outputs(2816) <= a or b;
    outputs(2817) <= b;
    outputs(2818) <= not a;
    outputs(2819) <= not a;
    outputs(2820) <= b;
    outputs(2821) <= a and b;
    outputs(2822) <= not a or b;
    outputs(2823) <= b;
    outputs(2824) <= not a or b;
    outputs(2825) <= a xor b;
    outputs(2826) <= b and not a;
    outputs(2827) <= a and not b;
    outputs(2828) <= a xor b;
    outputs(2829) <= b;
    outputs(2830) <= not b;
    outputs(2831) <= b and not a;
    outputs(2832) <= not (a and b);
    outputs(2833) <= not b;
    outputs(2834) <= a and not b;
    outputs(2835) <= not (a xor b);
    outputs(2836) <= not (a xor b);
    outputs(2837) <= a and b;
    outputs(2838) <= not b;
    outputs(2839) <= not (a or b);
    outputs(2840) <= b and not a;
    outputs(2841) <= not (a and b);
    outputs(2842) <= a xor b;
    outputs(2843) <= not a;
    outputs(2844) <= a xor b;
    outputs(2845) <= not (a xor b);
    outputs(2846) <= b and not a;
    outputs(2847) <= a or b;
    outputs(2848) <= b;
    outputs(2849) <= a xor b;
    outputs(2850) <= not (a xor b);
    outputs(2851) <= a;
    outputs(2852) <= b;
    outputs(2853) <= b;
    outputs(2854) <= not (a xor b);
    outputs(2855) <= not a;
    outputs(2856) <= not (a xor b);
    outputs(2857) <= not (a or b);
    outputs(2858) <= a and not b;
    outputs(2859) <= a and b;
    outputs(2860) <= not (a xor b);
    outputs(2861) <= not b;
    outputs(2862) <= not (a xor b);
    outputs(2863) <= a xor b;
    outputs(2864) <= a or b;
    outputs(2865) <= not b or a;
    outputs(2866) <= not (a xor b);
    outputs(2867) <= b and not a;
    outputs(2868) <= not b;
    outputs(2869) <= a or b;
    outputs(2870) <= b and not a;
    outputs(2871) <= b;
    outputs(2872) <= not a or b;
    outputs(2873) <= not b;
    outputs(2874) <= not a;
    outputs(2875) <= a;
    outputs(2876) <= not (a xor b);
    outputs(2877) <= not (a xor b);
    outputs(2878) <= not (a xor b);
    outputs(2879) <= not (a xor b);
    outputs(2880) <= not (a xor b);
    outputs(2881) <= not a;
    outputs(2882) <= a and not b;
    outputs(2883) <= not a;
    outputs(2884) <= a;
    outputs(2885) <= a;
    outputs(2886) <= b;
    outputs(2887) <= not a or b;
    outputs(2888) <= b;
    outputs(2889) <= b and not a;
    outputs(2890) <= a and b;
    outputs(2891) <= not a;
    outputs(2892) <= not (a xor b);
    outputs(2893) <= not a;
    outputs(2894) <= a and b;
    outputs(2895) <= b;
    outputs(2896) <= not (a and b);
    outputs(2897) <= not a;
    outputs(2898) <= not a;
    outputs(2899) <= a or b;
    outputs(2900) <= a;
    outputs(2901) <= not (a or b);
    outputs(2902) <= a xor b;
    outputs(2903) <= a xor b;
    outputs(2904) <= a xor b;
    outputs(2905) <= b;
    outputs(2906) <= not (a and b);
    outputs(2907) <= not b;
    outputs(2908) <= a;
    outputs(2909) <= a;
    outputs(2910) <= not a or b;
    outputs(2911) <= b;
    outputs(2912) <= a;
    outputs(2913) <= a xor b;
    outputs(2914) <= a and b;
    outputs(2915) <= not b;
    outputs(2916) <= not b or a;
    outputs(2917) <= not b or a;
    outputs(2918) <= a or b;
    outputs(2919) <= b and not a;
    outputs(2920) <= not b;
    outputs(2921) <= a xor b;
    outputs(2922) <= not a;
    outputs(2923) <= b;
    outputs(2924) <= not (a xor b);
    outputs(2925) <= a or b;
    outputs(2926) <= a;
    outputs(2927) <= b and not a;
    outputs(2928) <= a or b;
    outputs(2929) <= not (a xor b);
    outputs(2930) <= not a;
    outputs(2931) <= a xor b;
    outputs(2932) <= a xor b;
    outputs(2933) <= a xor b;
    outputs(2934) <= not a;
    outputs(2935) <= a xor b;
    outputs(2936) <= not (a xor b);
    outputs(2937) <= a;
    outputs(2938) <= a xor b;
    outputs(2939) <= a xor b;
    outputs(2940) <= not b;
    outputs(2941) <= a and b;
    outputs(2942) <= not (a and b);
    outputs(2943) <= a;
    outputs(2944) <= a xor b;
    outputs(2945) <= not (a xor b);
    outputs(2946) <= not (a or b);
    outputs(2947) <= not a;
    outputs(2948) <= b;
    outputs(2949) <= a xor b;
    outputs(2950) <= b;
    outputs(2951) <= not (a and b);
    outputs(2952) <= a xor b;
    outputs(2953) <= b;
    outputs(2954) <= not a;
    outputs(2955) <= a and b;
    outputs(2956) <= a xor b;
    outputs(2957) <= a and b;
    outputs(2958) <= a;
    outputs(2959) <= a or b;
    outputs(2960) <= not (a xor b);
    outputs(2961) <= b;
    outputs(2962) <= a xor b;
    outputs(2963) <= a;
    outputs(2964) <= not b or a;
    outputs(2965) <= not a;
    outputs(2966) <= not a;
    outputs(2967) <= a and not b;
    outputs(2968) <= not (a and b);
    outputs(2969) <= a and b;
    outputs(2970) <= a;
    outputs(2971) <= not (a or b);
    outputs(2972) <= not (a xor b);
    outputs(2973) <= a xor b;
    outputs(2974) <= a;
    outputs(2975) <= a or b;
    outputs(2976) <= not (a and b);
    outputs(2977) <= not a;
    outputs(2978) <= not b;
    outputs(2979) <= a;
    outputs(2980) <= not (a and b);
    outputs(2981) <= a and not b;
    outputs(2982) <= not (a or b);
    outputs(2983) <= b;
    outputs(2984) <= not (a and b);
    outputs(2985) <= not a;
    outputs(2986) <= a and not b;
    outputs(2987) <= not (a and b);
    outputs(2988) <= b and not a;
    outputs(2989) <= b;
    outputs(2990) <= a;
    outputs(2991) <= a;
    outputs(2992) <= not a;
    outputs(2993) <= a or b;
    outputs(2994) <= b;
    outputs(2995) <= not a;
    outputs(2996) <= a xor b;
    outputs(2997) <= not (a and b);
    outputs(2998) <= a xor b;
    outputs(2999) <= b;
    outputs(3000) <= not b;
    outputs(3001) <= a;
    outputs(3002) <= not b;
    outputs(3003) <= a or b;
    outputs(3004) <= a;
    outputs(3005) <= not a;
    outputs(3006) <= not a or b;
    outputs(3007) <= a;
    outputs(3008) <= b and not a;
    outputs(3009) <= a;
    outputs(3010) <= not a;
    outputs(3011) <= not a;
    outputs(3012) <= not b or a;
    outputs(3013) <= b and not a;
    outputs(3014) <= not a;
    outputs(3015) <= not (a and b);
    outputs(3016) <= a;
    outputs(3017) <= a and b;
    outputs(3018) <= not b;
    outputs(3019) <= a or b;
    outputs(3020) <= b and not a;
    outputs(3021) <= not b;
    outputs(3022) <= not a;
    outputs(3023) <= not b;
    outputs(3024) <= a and not b;
    outputs(3025) <= a or b;
    outputs(3026) <= not b;
    outputs(3027) <= a xor b;
    outputs(3028) <= not (a or b);
    outputs(3029) <= a and b;
    outputs(3030) <= not b;
    outputs(3031) <= not (a xor b);
    outputs(3032) <= b and not a;
    outputs(3033) <= not a or b;
    outputs(3034) <= a;
    outputs(3035) <= not (a or b);
    outputs(3036) <= not b or a;
    outputs(3037) <= not (a xor b);
    outputs(3038) <= a xor b;
    outputs(3039) <= a;
    outputs(3040) <= not a;
    outputs(3041) <= a and not b;
    outputs(3042) <= not (a xor b);
    outputs(3043) <= a and b;
    outputs(3044) <= a;
    outputs(3045) <= a;
    outputs(3046) <= not a;
    outputs(3047) <= a xor b;
    outputs(3048) <= a and not b;
    outputs(3049) <= not b;
    outputs(3050) <= not (a and b);
    outputs(3051) <= a or b;
    outputs(3052) <= a xor b;
    outputs(3053) <= b;
    outputs(3054) <= not a;
    outputs(3055) <= not (a xor b);
    outputs(3056) <= not (a and b);
    outputs(3057) <= not b;
    outputs(3058) <= a and not b;
    outputs(3059) <= not (a xor b);
    outputs(3060) <= not b;
    outputs(3061) <= a;
    outputs(3062) <= not (a xor b);
    outputs(3063) <= not b or a;
    outputs(3064) <= b;
    outputs(3065) <= b;
    outputs(3066) <= not a;
    outputs(3067) <= not (a xor b);
    outputs(3068) <= a xor b;
    outputs(3069) <= b and not a;
    outputs(3070) <= b;
    outputs(3071) <= not (a xor b);
    outputs(3072) <= a xor b;
    outputs(3073) <= not (a xor b);
    outputs(3074) <= not (a xor b);
    outputs(3075) <= a and not b;
    outputs(3076) <= b and not a;
    outputs(3077) <= a;
    outputs(3078) <= b and not a;
    outputs(3079) <= not a;
    outputs(3080) <= not (a xor b);
    outputs(3081) <= a;
    outputs(3082) <= not b;
    outputs(3083) <= a and b;
    outputs(3084) <= not b;
    outputs(3085) <= not b;
    outputs(3086) <= b;
    outputs(3087) <= not b;
    outputs(3088) <= b;
    outputs(3089) <= a and b;
    outputs(3090) <= b;
    outputs(3091) <= not a;
    outputs(3092) <= b and not a;
    outputs(3093) <= a;
    outputs(3094) <= not (a xor b);
    outputs(3095) <= b;
    outputs(3096) <= not (a and b);
    outputs(3097) <= not a;
    outputs(3098) <= not (a and b);
    outputs(3099) <= not b;
    outputs(3100) <= not a;
    outputs(3101) <= b and not a;
    outputs(3102) <= a;
    outputs(3103) <= b and not a;
    outputs(3104) <= not (a or b);
    outputs(3105) <= b and not a;
    outputs(3106) <= a xor b;
    outputs(3107) <= a xor b;
    outputs(3108) <= b;
    outputs(3109) <= not a;
    outputs(3110) <= a;
    outputs(3111) <= b;
    outputs(3112) <= b;
    outputs(3113) <= a and b;
    outputs(3114) <= a xor b;
    outputs(3115) <= not a;
    outputs(3116) <= not a;
    outputs(3117) <= a;
    outputs(3118) <= not (a or b);
    outputs(3119) <= not b;
    outputs(3120) <= b;
    outputs(3121) <= not (a xor b);
    outputs(3122) <= a;
    outputs(3123) <= not a;
    outputs(3124) <= a;
    outputs(3125) <= a;
    outputs(3126) <= a or b;
    outputs(3127) <= a;
    outputs(3128) <= not a;
    outputs(3129) <= a and not b;
    outputs(3130) <= a and b;
    outputs(3131) <= not (a and b);
    outputs(3132) <= b;
    outputs(3133) <= not a;
    outputs(3134) <= a xor b;
    outputs(3135) <= a and b;
    outputs(3136) <= not a or b;
    outputs(3137) <= not b;
    outputs(3138) <= a or b;
    outputs(3139) <= not (a xor b);
    outputs(3140) <= not b;
    outputs(3141) <= not (a xor b);
    outputs(3142) <= b;
    outputs(3143) <= not (a or b);
    outputs(3144) <= not b;
    outputs(3145) <= a and b;
    outputs(3146) <= not b;
    outputs(3147) <= a xor b;
    outputs(3148) <= b and not a;
    outputs(3149) <= not a;
    outputs(3150) <= a;
    outputs(3151) <= not a;
    outputs(3152) <= not (a xor b);
    outputs(3153) <= b;
    outputs(3154) <= not a;
    outputs(3155) <= not b or a;
    outputs(3156) <= a;
    outputs(3157) <= not (a xor b);
    outputs(3158) <= not (a xor b);
    outputs(3159) <= b;
    outputs(3160) <= not (a or b);
    outputs(3161) <= a xor b;
    outputs(3162) <= not (a or b);
    outputs(3163) <= not b;
    outputs(3164) <= not (a or b);
    outputs(3165) <= not a;
    outputs(3166) <= b and not a;
    outputs(3167) <= b and not a;
    outputs(3168) <= b and not a;
    outputs(3169) <= b and not a;
    outputs(3170) <= b;
    outputs(3171) <= not a;
    outputs(3172) <= b and not a;
    outputs(3173) <= a;
    outputs(3174) <= not b;
    outputs(3175) <= not b or a;
    outputs(3176) <= a xor b;
    outputs(3177) <= not a;
    outputs(3178) <= not a or b;
    outputs(3179) <= a and not b;
    outputs(3180) <= a and b;
    outputs(3181) <= a xor b;
    outputs(3182) <= not (a or b);
    outputs(3183) <= a xor b;
    outputs(3184) <= a or b;
    outputs(3185) <= a;
    outputs(3186) <= not a;
    outputs(3187) <= a and b;
    outputs(3188) <= b;
    outputs(3189) <= not (a xor b);
    outputs(3190) <= not (a or b);
    outputs(3191) <= not (a xor b);
    outputs(3192) <= not b;
    outputs(3193) <= a xor b;
    outputs(3194) <= not a;
    outputs(3195) <= not (a or b);
    outputs(3196) <= a;
    outputs(3197) <= a and not b;
    outputs(3198) <= a and not b;
    outputs(3199) <= not b or a;
    outputs(3200) <= a xor b;
    outputs(3201) <= a and not b;
    outputs(3202) <= not b;
    outputs(3203) <= a or b;
    outputs(3204) <= b;
    outputs(3205) <= not b;
    outputs(3206) <= not b;
    outputs(3207) <= not b;
    outputs(3208) <= a;
    outputs(3209) <= not a or b;
    outputs(3210) <= a xor b;
    outputs(3211) <= a xor b;
    outputs(3212) <= not b;
    outputs(3213) <= not (a or b);
    outputs(3214) <= a and not b;
    outputs(3215) <= not b;
    outputs(3216) <= b;
    outputs(3217) <= not b;
    outputs(3218) <= not (a and b);
    outputs(3219) <= b and not a;
    outputs(3220) <= not b;
    outputs(3221) <= a and b;
    outputs(3222) <= a xor b;
    outputs(3223) <= not (a xor b);
    outputs(3224) <= not (a or b);
    outputs(3225) <= b;
    outputs(3226) <= a and b;
    outputs(3227) <= not (a and b);
    outputs(3228) <= not b or a;
    outputs(3229) <= b;
    outputs(3230) <= a and b;
    outputs(3231) <= not a or b;
    outputs(3232) <= a;
    outputs(3233) <= b and not a;
    outputs(3234) <= not a;
    outputs(3235) <= not a or b;
    outputs(3236) <= not (a xor b);
    outputs(3237) <= not b or a;
    outputs(3238) <= not (a or b);
    outputs(3239) <= a and not b;
    outputs(3240) <= a and b;
    outputs(3241) <= b and not a;
    outputs(3242) <= not (a or b);
    outputs(3243) <= not a;
    outputs(3244) <= a and b;
    outputs(3245) <= not (a or b);
    outputs(3246) <= not b;
    outputs(3247) <= not b;
    outputs(3248) <= not (a or b);
    outputs(3249) <= not a;
    outputs(3250) <= not b;
    outputs(3251) <= not a;
    outputs(3252) <= a and not b;
    outputs(3253) <= not b;
    outputs(3254) <= not b;
    outputs(3255) <= not (a or b);
    outputs(3256) <= not a;
    outputs(3257) <= not a;
    outputs(3258) <= not a;
    outputs(3259) <= b;
    outputs(3260) <= a and not b;
    outputs(3261) <= not b or a;
    outputs(3262) <= a xor b;
    outputs(3263) <= b and not a;
    outputs(3264) <= not a;
    outputs(3265) <= a or b;
    outputs(3266) <= a xor b;
    outputs(3267) <= a and b;
    outputs(3268) <= b and not a;
    outputs(3269) <= a;
    outputs(3270) <= b;
    outputs(3271) <= not (a or b);
    outputs(3272) <= a xor b;
    outputs(3273) <= a and not b;
    outputs(3274) <= not a or b;
    outputs(3275) <= a xor b;
    outputs(3276) <= not (a and b);
    outputs(3277) <= not (a or b);
    outputs(3278) <= not b;
    outputs(3279) <= a and not b;
    outputs(3280) <= a and not b;
    outputs(3281) <= a and b;
    outputs(3282) <= a;
    outputs(3283) <= a xor b;
    outputs(3284) <= a xor b;
    outputs(3285) <= a and b;
    outputs(3286) <= a;
    outputs(3287) <= not (a xor b);
    outputs(3288) <= a;
    outputs(3289) <= b;
    outputs(3290) <= not (a xor b);
    outputs(3291) <= a and not b;
    outputs(3292) <= b and not a;
    outputs(3293) <= b;
    outputs(3294) <= b;
    outputs(3295) <= a;
    outputs(3296) <= not b or a;
    outputs(3297) <= not (a xor b);
    outputs(3298) <= not (a and b);
    outputs(3299) <= not b;
    outputs(3300) <= a and not b;
    outputs(3301) <= not (a or b);
    outputs(3302) <= b and not a;
    outputs(3303) <= b;
    outputs(3304) <= b;
    outputs(3305) <= a and b;
    outputs(3306) <= a;
    outputs(3307) <= a and b;
    outputs(3308) <= not (a or b);
    outputs(3309) <= a;
    outputs(3310) <= b and not a;
    outputs(3311) <= a;
    outputs(3312) <= not (a xor b);
    outputs(3313) <= not (a xor b);
    outputs(3314) <= not b;
    outputs(3315) <= b;
    outputs(3316) <= not a or b;
    outputs(3317) <= not (a xor b);
    outputs(3318) <= not b;
    outputs(3319) <= not b;
    outputs(3320) <= b;
    outputs(3321) <= not (a xor b);
    outputs(3322) <= not b;
    outputs(3323) <= a;
    outputs(3324) <= not (a xor b);
    outputs(3325) <= a and b;
    outputs(3326) <= not a;
    outputs(3327) <= not b;
    outputs(3328) <= a and not b;
    outputs(3329) <= a xor b;
    outputs(3330) <= not b;
    outputs(3331) <= a;
    outputs(3332) <= not (a xor b);
    outputs(3333) <= a and b;
    outputs(3334) <= a;
    outputs(3335) <= not (a or b);
    outputs(3336) <= a and not b;
    outputs(3337) <= a or b;
    outputs(3338) <= b and not a;
    outputs(3339) <= not (a or b);
    outputs(3340) <= not b or a;
    outputs(3341) <= not (a or b);
    outputs(3342) <= b;
    outputs(3343) <= not (a xor b);
    outputs(3344) <= not a;
    outputs(3345) <= not b;
    outputs(3346) <= not b;
    outputs(3347) <= b;
    outputs(3348) <= a;
    outputs(3349) <= a and not b;
    outputs(3350) <= b;
    outputs(3351) <= a;
    outputs(3352) <= a and b;
    outputs(3353) <= not (a xor b);
    outputs(3354) <= not (a or b);
    outputs(3355) <= b;
    outputs(3356) <= a and not b;
    outputs(3357) <= b;
    outputs(3358) <= a;
    outputs(3359) <= not (a and b);
    outputs(3360) <= b and not a;
    outputs(3361) <= b;
    outputs(3362) <= not b;
    outputs(3363) <= not b;
    outputs(3364) <= a;
    outputs(3365) <= a;
    outputs(3366) <= not b;
    outputs(3367) <= a or b;
    outputs(3368) <= a xor b;
    outputs(3369) <= a;
    outputs(3370) <= a;
    outputs(3371) <= b;
    outputs(3372) <= not b;
    outputs(3373) <= not b;
    outputs(3374) <= not (a or b);
    outputs(3375) <= a or b;
    outputs(3376) <= a and not b;
    outputs(3377) <= a and not b;
    outputs(3378) <= b and not a;
    outputs(3379) <= a;
    outputs(3380) <= b;
    outputs(3381) <= b;
    outputs(3382) <= not b;
    outputs(3383) <= b;
    outputs(3384) <= not b;
    outputs(3385) <= a;
    outputs(3386) <= a and b;
    outputs(3387) <= not (a xor b);
    outputs(3388) <= not b;
    outputs(3389) <= b and not a;
    outputs(3390) <= a;
    outputs(3391) <= a xor b;
    outputs(3392) <= not (a or b);
    outputs(3393) <= a xor b;
    outputs(3394) <= not a;
    outputs(3395) <= not a;
    outputs(3396) <= a or b;
    outputs(3397) <= not (a or b);
    outputs(3398) <= not (a or b);
    outputs(3399) <= a xor b;
    outputs(3400) <= b;
    outputs(3401) <= not (a or b);
    outputs(3402) <= not a;
    outputs(3403) <= not (a and b);
    outputs(3404) <= not (a xor b);
    outputs(3405) <= a;
    outputs(3406) <= not a;
    outputs(3407) <= not a or b;
    outputs(3408) <= not (a and b);
    outputs(3409) <= a xor b;
    outputs(3410) <= b;
    outputs(3411) <= not b;
    outputs(3412) <= not a;
    outputs(3413) <= not (a xor b);
    outputs(3414) <= not a;
    outputs(3415) <= not (a or b);
    outputs(3416) <= not a or b;
    outputs(3417) <= not a;
    outputs(3418) <= not a;
    outputs(3419) <= not (a xor b);
    outputs(3420) <= a and b;
    outputs(3421) <= not b or a;
    outputs(3422) <= not a;
    outputs(3423) <= not a;
    outputs(3424) <= a;
    outputs(3425) <= b;
    outputs(3426) <= a and not b;
    outputs(3427) <= not a or b;
    outputs(3428) <= a;
    outputs(3429) <= not (a or b);
    outputs(3430) <= not a or b;
    outputs(3431) <= not (a or b);
    outputs(3432) <= not b;
    outputs(3433) <= not (a or b);
    outputs(3434) <= b;
    outputs(3435) <= not (a xor b);
    outputs(3436) <= b;
    outputs(3437) <= not a;
    outputs(3438) <= b and not a;
    outputs(3439) <= b;
    outputs(3440) <= b;
    outputs(3441) <= b;
    outputs(3442) <= not b or a;
    outputs(3443) <= a xor b;
    outputs(3444) <= not (a or b);
    outputs(3445) <= not b;
    outputs(3446) <= not a;
    outputs(3447) <= not a;
    outputs(3448) <= a and b;
    outputs(3449) <= not (a xor b);
    outputs(3450) <= not b;
    outputs(3451) <= b;
    outputs(3452) <= a;
    outputs(3453) <= a;
    outputs(3454) <= a and not b;
    outputs(3455) <= a xor b;
    outputs(3456) <= b;
    outputs(3457) <= b;
    outputs(3458) <= not b;
    outputs(3459) <= not (a and b);
    outputs(3460) <= not b;
    outputs(3461) <= not (a xor b);
    outputs(3462) <= a xor b;
    outputs(3463) <= a and b;
    outputs(3464) <= b and not a;
    outputs(3465) <= b and not a;
    outputs(3466) <= a and not b;
    outputs(3467) <= a or b;
    outputs(3468) <= a;
    outputs(3469) <= not b or a;
    outputs(3470) <= a and not b;
    outputs(3471) <= b and not a;
    outputs(3472) <= not a;
    outputs(3473) <= a xor b;
    outputs(3474) <= not (a xor b);
    outputs(3475) <= b and not a;
    outputs(3476) <= not (a xor b);
    outputs(3477) <= a;
    outputs(3478) <= not (a xor b);
    outputs(3479) <= b and not a;
    outputs(3480) <= b;
    outputs(3481) <= a and not b;
    outputs(3482) <= not a;
    outputs(3483) <= b;
    outputs(3484) <= a xor b;
    outputs(3485) <= not a;
    outputs(3486) <= not (a and b);
    outputs(3487) <= not (a xor b);
    outputs(3488) <= not b or a;
    outputs(3489) <= a xor b;
    outputs(3490) <= not a;
    outputs(3491) <= not b;
    outputs(3492) <= a or b;
    outputs(3493) <= b and not a;
    outputs(3494) <= a and b;
    outputs(3495) <= not (a and b);
    outputs(3496) <= not (a xor b);
    outputs(3497) <= b;
    outputs(3498) <= a and b;
    outputs(3499) <= not a;
    outputs(3500) <= a and not b;
    outputs(3501) <= not b or a;
    outputs(3502) <= a and b;
    outputs(3503) <= b;
    outputs(3504) <= a and b;
    outputs(3505) <= a xor b;
    outputs(3506) <= b and not a;
    outputs(3507) <= b;
    outputs(3508) <= not (a xor b);
    outputs(3509) <= a and not b;
    outputs(3510) <= not (a and b);
    outputs(3511) <= b;
    outputs(3512) <= a;
    outputs(3513) <= b;
    outputs(3514) <= a;
    outputs(3515) <= a;
    outputs(3516) <= not a;
    outputs(3517) <= a;
    outputs(3518) <= not b;
    outputs(3519) <= not (a or b);
    outputs(3520) <= a xor b;
    outputs(3521) <= a xor b;
    outputs(3522) <= b;
    outputs(3523) <= a and b;
    outputs(3524) <= not (a or b);
    outputs(3525) <= a and not b;
    outputs(3526) <= not a;
    outputs(3527) <= a xor b;
    outputs(3528) <= not b;
    outputs(3529) <= a xor b;
    outputs(3530) <= not (a xor b);
    outputs(3531) <= a and b;
    outputs(3532) <= not (a or b);
    outputs(3533) <= a and not b;
    outputs(3534) <= a xor b;
    outputs(3535) <= not (a xor b);
    outputs(3536) <= b;
    outputs(3537) <= not (a xor b);
    outputs(3538) <= b;
    outputs(3539) <= b;
    outputs(3540) <= not b;
    outputs(3541) <= b and not a;
    outputs(3542) <= not b;
    outputs(3543) <= b and not a;
    outputs(3544) <= not a;
    outputs(3545) <= not b;
    outputs(3546) <= not b;
    outputs(3547) <= b and not a;
    outputs(3548) <= b and not a;
    outputs(3549) <= b and not a;
    outputs(3550) <= a xor b;
    outputs(3551) <= not b;
    outputs(3552) <= a and not b;
    outputs(3553) <= b;
    outputs(3554) <= b and not a;
    outputs(3555) <= not a;
    outputs(3556) <= not b;
    outputs(3557) <= a;
    outputs(3558) <= not (a or b);
    outputs(3559) <= a;
    outputs(3560) <= not (a xor b);
    outputs(3561) <= not a;
    outputs(3562) <= not (a xor b);
    outputs(3563) <= a;
    outputs(3564) <= a and b;
    outputs(3565) <= not (a xor b);
    outputs(3566) <= not b;
    outputs(3567) <= not b;
    outputs(3568) <= b;
    outputs(3569) <= a;
    outputs(3570) <= b;
    outputs(3571) <= not b;
    outputs(3572) <= not b;
    outputs(3573) <= a;
    outputs(3574) <= a xor b;
    outputs(3575) <= not a;
    outputs(3576) <= a and not b;
    outputs(3577) <= not a;
    outputs(3578) <= not a;
    outputs(3579) <= not b;
    outputs(3580) <= b and not a;
    outputs(3581) <= not (a or b);
    outputs(3582) <= a;
    outputs(3583) <= not (a xor b);
    outputs(3584) <= a xor b;
    outputs(3585) <= a xor b;
    outputs(3586) <= not a or b;
    outputs(3587) <= a;
    outputs(3588) <= not (a or b);
    outputs(3589) <= not a;
    outputs(3590) <= a;
    outputs(3591) <= not b;
    outputs(3592) <= a xor b;
    outputs(3593) <= not (a xor b);
    outputs(3594) <= not (a xor b);
    outputs(3595) <= not a;
    outputs(3596) <= a xor b;
    outputs(3597) <= not (a or b);
    outputs(3598) <= not (a or b);
    outputs(3599) <= b and not a;
    outputs(3600) <= not a;
    outputs(3601) <= not a;
    outputs(3602) <= not a or b;
    outputs(3603) <= not (a and b);
    outputs(3604) <= not (a xor b);
    outputs(3605) <= not b or a;
    outputs(3606) <= a and b;
    outputs(3607) <= not b or a;
    outputs(3608) <= a and not b;
    outputs(3609) <= not (a xor b);
    outputs(3610) <= not (a xor b);
    outputs(3611) <= b;
    outputs(3612) <= not a;
    outputs(3613) <= a and not b;
    outputs(3614) <= a xor b;
    outputs(3615) <= a xor b;
    outputs(3616) <= a;
    outputs(3617) <= not (a or b);
    outputs(3618) <= a and not b;
    outputs(3619) <= a and b;
    outputs(3620) <= b and not a;
    outputs(3621) <= not a;
    outputs(3622) <= b and not a;
    outputs(3623) <= not a;
    outputs(3624) <= not (a xor b);
    outputs(3625) <= a and b;
    outputs(3626) <= b and not a;
    outputs(3627) <= not a;
    outputs(3628) <= a xor b;
    outputs(3629) <= a;
    outputs(3630) <= not b;
    outputs(3631) <= not (a xor b);
    outputs(3632) <= not a;
    outputs(3633) <= a;
    outputs(3634) <= not (a xor b);
    outputs(3635) <= b;
    outputs(3636) <= not b;
    outputs(3637) <= not b;
    outputs(3638) <= not b;
    outputs(3639) <= not b;
    outputs(3640) <= a;
    outputs(3641) <= not (a xor b);
    outputs(3642) <= a or b;
    outputs(3643) <= b;
    outputs(3644) <= a;
    outputs(3645) <= not b;
    outputs(3646) <= not b or a;
    outputs(3647) <= not (a xor b);
    outputs(3648) <= not (a or b);
    outputs(3649) <= not a;
    outputs(3650) <= a or b;
    outputs(3651) <= not a;
    outputs(3652) <= a;
    outputs(3653) <= a and b;
    outputs(3654) <= b;
    outputs(3655) <= not a;
    outputs(3656) <= a;
    outputs(3657) <= a;
    outputs(3658) <= b and not a;
    outputs(3659) <= not (a and b);
    outputs(3660) <= not b;
    outputs(3661) <= not (a xor b);
    outputs(3662) <= a xor b;
    outputs(3663) <= not a;
    outputs(3664) <= a and not b;
    outputs(3665) <= a and b;
    outputs(3666) <= a and b;
    outputs(3667) <= a;
    outputs(3668) <= a xor b;
    outputs(3669) <= not (a xor b);
    outputs(3670) <= not b;
    outputs(3671) <= not b or a;
    outputs(3672) <= a or b;
    outputs(3673) <= a xor b;
    outputs(3674) <= not a;
    outputs(3675) <= not a;
    outputs(3676) <= not (a or b);
    outputs(3677) <= not b;
    outputs(3678) <= not a;
    outputs(3679) <= b and not a;
    outputs(3680) <= a;
    outputs(3681) <= not b;
    outputs(3682) <= b and not a;
    outputs(3683) <= not a;
    outputs(3684) <= a;
    outputs(3685) <= a xor b;
    outputs(3686) <= not (a and b);
    outputs(3687) <= a and b;
    outputs(3688) <= not b;
    outputs(3689) <= not b;
    outputs(3690) <= a;
    outputs(3691) <= not a;
    outputs(3692) <= a and b;
    outputs(3693) <= a;
    outputs(3694) <= not a;
    outputs(3695) <= not a;
    outputs(3696) <= a;
    outputs(3697) <= not (a or b);
    outputs(3698) <= not (a or b);
    outputs(3699) <= a and not b;
    outputs(3700) <= not a;
    outputs(3701) <= not a;
    outputs(3702) <= not a or b;
    outputs(3703) <= not (a and b);
    outputs(3704) <= not (a or b);
    outputs(3705) <= a and b;
    outputs(3706) <= not (a or b);
    outputs(3707) <= a xor b;
    outputs(3708) <= b and not a;
    outputs(3709) <= not b;
    outputs(3710) <= not (a xor b);
    outputs(3711) <= not b;
    outputs(3712) <= b;
    outputs(3713) <= a;
    outputs(3714) <= a;
    outputs(3715) <= not (a xor b);
    outputs(3716) <= not b;
    outputs(3717) <= b and not a;
    outputs(3718) <= a and not b;
    outputs(3719) <= not a;
    outputs(3720) <= b;
    outputs(3721) <= b;
    outputs(3722) <= b;
    outputs(3723) <= not b;
    outputs(3724) <= b;
    outputs(3725) <= not b;
    outputs(3726) <= not a;
    outputs(3727) <= not a;
    outputs(3728) <= not (a or b);
    outputs(3729) <= b;
    outputs(3730) <= a;
    outputs(3731) <= not a;
    outputs(3732) <= b and not a;
    outputs(3733) <= not b;
    outputs(3734) <= not b;
    outputs(3735) <= a xor b;
    outputs(3736) <= b and not a;
    outputs(3737) <= not b or a;
    outputs(3738) <= b;
    outputs(3739) <= a xor b;
    outputs(3740) <= a;
    outputs(3741) <= b and not a;
    outputs(3742) <= not b or a;
    outputs(3743) <= not b;
    outputs(3744) <= a and b;
    outputs(3745) <= not b;
    outputs(3746) <= not b;
    outputs(3747) <= a;
    outputs(3748) <= b and not a;
    outputs(3749) <= b;
    outputs(3750) <= not a;
    outputs(3751) <= not b;
    outputs(3752) <= not (a or b);
    outputs(3753) <= not (a or b);
    outputs(3754) <= not b;
    outputs(3755) <= not a;
    outputs(3756) <= not b;
    outputs(3757) <= a;
    outputs(3758) <= not b;
    outputs(3759) <= a;
    outputs(3760) <= b;
    outputs(3761) <= a xor b;
    outputs(3762) <= not b;
    outputs(3763) <= not (a or b);
    outputs(3764) <= not (a xor b);
    outputs(3765) <= not (a xor b);
    outputs(3766) <= not (a xor b);
    outputs(3767) <= a and not b;
    outputs(3768) <= not (a or b);
    outputs(3769) <= not (a and b);
    outputs(3770) <= a;
    outputs(3771) <= a xor b;
    outputs(3772) <= not b;
    outputs(3773) <= not b;
    outputs(3774) <= a;
    outputs(3775) <= not (a or b);
    outputs(3776) <= not a;
    outputs(3777) <= a and b;
    outputs(3778) <= a and not b;
    outputs(3779) <= not (a or b);
    outputs(3780) <= not a or b;
    outputs(3781) <= b and not a;
    outputs(3782) <= not (a xor b);
    outputs(3783) <= a xor b;
    outputs(3784) <= a and not b;
    outputs(3785) <= not a;
    outputs(3786) <= a;
    outputs(3787) <= not a;
    outputs(3788) <= not b;
    outputs(3789) <= a xor b;
    outputs(3790) <= not a;
    outputs(3791) <= not a;
    outputs(3792) <= a and b;
    outputs(3793) <= b and not a;
    outputs(3794) <= not b;
    outputs(3795) <= a and b;
    outputs(3796) <= not (a xor b);
    outputs(3797) <= b and not a;
    outputs(3798) <= a or b;
    outputs(3799) <= not a or b;
    outputs(3800) <= a or b;
    outputs(3801) <= a and not b;
    outputs(3802) <= not a;
    outputs(3803) <= not b or a;
    outputs(3804) <= not (a xor b);
    outputs(3805) <= not (a or b);
    outputs(3806) <= a xor b;
    outputs(3807) <= not a;
    outputs(3808) <= not a;
    outputs(3809) <= a;
    outputs(3810) <= b;
    outputs(3811) <= a and not b;
    outputs(3812) <= b;
    outputs(3813) <= a and b;
    outputs(3814) <= not (a xor b);
    outputs(3815) <= not a;
    outputs(3816) <= a xor b;
    outputs(3817) <= not b;
    outputs(3818) <= a;
    outputs(3819) <= a and b;
    outputs(3820) <= a;
    outputs(3821) <= a xor b;
    outputs(3822) <= a and not b;
    outputs(3823) <= a and b;
    outputs(3824) <= not b;
    outputs(3825) <= a;
    outputs(3826) <= not (a xor b);
    outputs(3827) <= a xor b;
    outputs(3828) <= a and not b;
    outputs(3829) <= not (a or b);
    outputs(3830) <= b;
    outputs(3831) <= a;
    outputs(3832) <= b and not a;
    outputs(3833) <= not b;
    outputs(3834) <= b;
    outputs(3835) <= a xor b;
    outputs(3836) <= a or b;
    outputs(3837) <= a and b;
    outputs(3838) <= not a or b;
    outputs(3839) <= a and not b;
    outputs(3840) <= not b;
    outputs(3841) <= b and not a;
    outputs(3842) <= a xor b;
    outputs(3843) <= not a;
    outputs(3844) <= b;
    outputs(3845) <= b and not a;
    outputs(3846) <= not b;
    outputs(3847) <= a and b;
    outputs(3848) <= not b or a;
    outputs(3849) <= a xor b;
    outputs(3850) <= not a;
    outputs(3851) <= not (a xor b);
    outputs(3852) <= b;
    outputs(3853) <= a xor b;
    outputs(3854) <= not (a or b);
    outputs(3855) <= b;
    outputs(3856) <= a;
    outputs(3857) <= a;
    outputs(3858) <= a and not b;
    outputs(3859) <= not (a xor b);
    outputs(3860) <= a or b;
    outputs(3861) <= b;
    outputs(3862) <= not b or a;
    outputs(3863) <= not (a xor b);
    outputs(3864) <= not (a xor b);
    outputs(3865) <= not a;
    outputs(3866) <= b and not a;
    outputs(3867) <= a and b;
    outputs(3868) <= not (a or b);
    outputs(3869) <= a;
    outputs(3870) <= a or b;
    outputs(3871) <= a and b;
    outputs(3872) <= b;
    outputs(3873) <= b;
    outputs(3874) <= not b or a;
    outputs(3875) <= a xor b;
    outputs(3876) <= not (a xor b);
    outputs(3877) <= a;
    outputs(3878) <= not (a or b);
    outputs(3879) <= not a;
    outputs(3880) <= b and not a;
    outputs(3881) <= not b;
    outputs(3882) <= a;
    outputs(3883) <= not a;
    outputs(3884) <= not (a xor b);
    outputs(3885) <= a or b;
    outputs(3886) <= not (a xor b);
    outputs(3887) <= not (a xor b);
    outputs(3888) <= a and b;
    outputs(3889) <= not (a xor b);
    outputs(3890) <= not (a xor b);
    outputs(3891) <= not (a xor b);
    outputs(3892) <= not b;
    outputs(3893) <= not a;
    outputs(3894) <= b;
    outputs(3895) <= b and not a;
    outputs(3896) <= not b;
    outputs(3897) <= not a;
    outputs(3898) <= not (a or b);
    outputs(3899) <= b;
    outputs(3900) <= a xor b;
    outputs(3901) <= a;
    outputs(3902) <= not a or b;
    outputs(3903) <= not b;
    outputs(3904) <= a xor b;
    outputs(3905) <= not a or b;
    outputs(3906) <= b;
    outputs(3907) <= not b;
    outputs(3908) <= a;
    outputs(3909) <= a and b;
    outputs(3910) <= not (a or b);
    outputs(3911) <= a or b;
    outputs(3912) <= not (a xor b);
    outputs(3913) <= not (a xor b);
    outputs(3914) <= a xor b;
    outputs(3915) <= a or b;
    outputs(3916) <= a;
    outputs(3917) <= a and b;
    outputs(3918) <= a and not b;
    outputs(3919) <= b and not a;
    outputs(3920) <= not b or a;
    outputs(3921) <= a xor b;
    outputs(3922) <= a and b;
    outputs(3923) <= a;
    outputs(3924) <= a;
    outputs(3925) <= not b;
    outputs(3926) <= not a;
    outputs(3927) <= not a or b;
    outputs(3928) <= a xor b;
    outputs(3929) <= not a;
    outputs(3930) <= not (a xor b);
    outputs(3931) <= a xor b;
    outputs(3932) <= not a;
    outputs(3933) <= not a;
    outputs(3934) <= not a;
    outputs(3935) <= not b;
    outputs(3936) <= not (a xor b);
    outputs(3937) <= a;
    outputs(3938) <= not (a or b);
    outputs(3939) <= not a or b;
    outputs(3940) <= not (a xor b);
    outputs(3941) <= a xor b;
    outputs(3942) <= not (a xor b);
    outputs(3943) <= b and not a;
    outputs(3944) <= not a or b;
    outputs(3945) <= a xor b;
    outputs(3946) <= not b;
    outputs(3947) <= not a;
    outputs(3948) <= a;
    outputs(3949) <= a xor b;
    outputs(3950) <= a;
    outputs(3951) <= a and not b;
    outputs(3952) <= not b;
    outputs(3953) <= b;
    outputs(3954) <= a xor b;
    outputs(3955) <= not (a or b);
    outputs(3956) <= b;
    outputs(3957) <= not (a xor b);
    outputs(3958) <= not (a xor b);
    outputs(3959) <= a;
    outputs(3960) <= not (a xor b);
    outputs(3961) <= not (a xor b);
    outputs(3962) <= not a or b;
    outputs(3963) <= a and b;
    outputs(3964) <= not (a xor b);
    outputs(3965) <= b;
    outputs(3966) <= a or b;
    outputs(3967) <= a xor b;
    outputs(3968) <= a;
    outputs(3969) <= not (a xor b);
    outputs(3970) <= b;
    outputs(3971) <= not (a xor b);
    outputs(3972) <= a xor b;
    outputs(3973) <= a and b;
    outputs(3974) <= a and not b;
    outputs(3975) <= not (a xor b);
    outputs(3976) <= a or b;
    outputs(3977) <= b;
    outputs(3978) <= b and not a;
    outputs(3979) <= b;
    outputs(3980) <= a xor b;
    outputs(3981) <= a and b;
    outputs(3982) <= a xor b;
    outputs(3983) <= a;
    outputs(3984) <= not b or a;
    outputs(3985) <= not b;
    outputs(3986) <= a;
    outputs(3987) <= not (a xor b);
    outputs(3988) <= b;
    outputs(3989) <= a;
    outputs(3990) <= not (a xor b);
    outputs(3991) <= b;
    outputs(3992) <= not (a xor b);
    outputs(3993) <= a and not b;
    outputs(3994) <= a xor b;
    outputs(3995) <= not (a xor b);
    outputs(3996) <= not (a xor b);
    outputs(3997) <= a;
    outputs(3998) <= not b or a;
    outputs(3999) <= not (a or b);
    outputs(4000) <= not b;
    outputs(4001) <= a;
    outputs(4002) <= a xor b;
    outputs(4003) <= not (a xor b);
    outputs(4004) <= not b;
    outputs(4005) <= b;
    outputs(4006) <= not a;
    outputs(4007) <= not b;
    outputs(4008) <= b and not a;
    outputs(4009) <= not (a or b);
    outputs(4010) <= not (a xor b);
    outputs(4011) <= a xor b;
    outputs(4012) <= a;
    outputs(4013) <= not (a or b);
    outputs(4014) <= not a;
    outputs(4015) <= not (a xor b);
    outputs(4016) <= not a;
    outputs(4017) <= not b;
    outputs(4018) <= a;
    outputs(4019) <= not b;
    outputs(4020) <= b and not a;
    outputs(4021) <= not b;
    outputs(4022) <= a and not b;
    outputs(4023) <= not a;
    outputs(4024) <= not a;
    outputs(4025) <= not (a xor b);
    outputs(4026) <= not b;
    outputs(4027) <= a and b;
    outputs(4028) <= a;
    outputs(4029) <= not (a xor b);
    outputs(4030) <= not a;
    outputs(4031) <= not b or a;
    outputs(4032) <= a xor b;
    outputs(4033) <= not a or b;
    outputs(4034) <= not (a xor b);
    outputs(4035) <= not a or b;
    outputs(4036) <= a;
    outputs(4037) <= b;
    outputs(4038) <= a;
    outputs(4039) <= not (a and b);
    outputs(4040) <= not (a xor b);
    outputs(4041) <= not (a or b);
    outputs(4042) <= a xor b;
    outputs(4043) <= not (a xor b);
    outputs(4044) <= not b;
    outputs(4045) <= a xor b;
    outputs(4046) <= not b;
    outputs(4047) <= not (a xor b);
    outputs(4048) <= not a;
    outputs(4049) <= a xor b;
    outputs(4050) <= b;
    outputs(4051) <= b;
    outputs(4052) <= b;
    outputs(4053) <= not a;
    outputs(4054) <= not (a and b);
    outputs(4055) <= not a;
    outputs(4056) <= not (a and b);
    outputs(4057) <= not (a xor b);
    outputs(4058) <= a;
    outputs(4059) <= b;
    outputs(4060) <= a xor b;
    outputs(4061) <= a;
    outputs(4062) <= not b or a;
    outputs(4063) <= b;
    outputs(4064) <= b;
    outputs(4065) <= a or b;
    outputs(4066) <= not b;
    outputs(4067) <= a and b;
    outputs(4068) <= not (a xor b);
    outputs(4069) <= not (a xor b);
    outputs(4070) <= not (a or b);
    outputs(4071) <= not (a or b);
    outputs(4072) <= b;
    outputs(4073) <= a and b;
    outputs(4074) <= not a;
    outputs(4075) <= a and not b;
    outputs(4076) <= a;
    outputs(4077) <= not (a xor b);
    outputs(4078) <= not (a or b);
    outputs(4079) <= a and b;
    outputs(4080) <= a and not b;
    outputs(4081) <= a;
    outputs(4082) <= b;
    outputs(4083) <= a xor b;
    outputs(4084) <= not (a or b);
    outputs(4085) <= b and not a;
    outputs(4086) <= a;
    outputs(4087) <= a xor b;
    outputs(4088) <= not a or b;
    outputs(4089) <= b and not a;
    outputs(4090) <= not a;
    outputs(4091) <= a and b;
    outputs(4092) <= not b;
    outputs(4093) <= a or b;
    outputs(4094) <= not a;
    outputs(4095) <= a;
    outputs(4096) <= a xor b;
    outputs(4097) <= a;
    outputs(4098) <= a xor b;
    outputs(4099) <= a xor b;
    outputs(4100) <= b;
    outputs(4101) <= not b;
    outputs(4102) <= a and b;
    outputs(4103) <= not (a xor b);
    outputs(4104) <= not (a and b);
    outputs(4105) <= not a or b;
    outputs(4106) <= not a or b;
    outputs(4107) <= a and b;
    outputs(4108) <= not (a xor b);
    outputs(4109) <= not a;
    outputs(4110) <= a;
    outputs(4111) <= a;
    outputs(4112) <= a xor b;
    outputs(4113) <= not (a and b);
    outputs(4114) <= not b;
    outputs(4115) <= not (a and b);
    outputs(4116) <= not a;
    outputs(4117) <= not a;
    outputs(4118) <= a;
    outputs(4119) <= a or b;
    outputs(4120) <= a;
    outputs(4121) <= a and not b;
    outputs(4122) <= a and b;
    outputs(4123) <= a;
    outputs(4124) <= a xor b;
    outputs(4125) <= a xor b;
    outputs(4126) <= a and b;
    outputs(4127) <= not (a xor b);
    outputs(4128) <= a and not b;
    outputs(4129) <= a and not b;
    outputs(4130) <= a or b;
    outputs(4131) <= not (a or b);
    outputs(4132) <= b;
    outputs(4133) <= b;
    outputs(4134) <= a xor b;
    outputs(4135) <= a;
    outputs(4136) <= not (a or b);
    outputs(4137) <= not a;
    outputs(4138) <= not (a xor b);
    outputs(4139) <= a and not b;
    outputs(4140) <= not (a and b);
    outputs(4141) <= b;
    outputs(4142) <= not (a and b);
    outputs(4143) <= not (a xor b);
    outputs(4144) <= b;
    outputs(4145) <= not b;
    outputs(4146) <= not b or a;
    outputs(4147) <= not (a xor b);
    outputs(4148) <= not (a or b);
    outputs(4149) <= not b;
    outputs(4150) <= not (a or b);
    outputs(4151) <= a xor b;
    outputs(4152) <= not b;
    outputs(4153) <= not (a xor b);
    outputs(4154) <= not b or a;
    outputs(4155) <= not b;
    outputs(4156) <= b and not a;
    outputs(4157) <= b;
    outputs(4158) <= not a or b;
    outputs(4159) <= not (a xor b);
    outputs(4160) <= a xor b;
    outputs(4161) <= b;
    outputs(4162) <= a xor b;
    outputs(4163) <= not a;
    outputs(4164) <= a and not b;
    outputs(4165) <= not b;
    outputs(4166) <= a xor b;
    outputs(4167) <= a;
    outputs(4168) <= not (a and b);
    outputs(4169) <= not a;
    outputs(4170) <= a;
    outputs(4171) <= not b;
    outputs(4172) <= not b or a;
    outputs(4173) <= not b;
    outputs(4174) <= not b;
    outputs(4175) <= a;
    outputs(4176) <= not (a xor b);
    outputs(4177) <= a and b;
    outputs(4178) <= a;
    outputs(4179) <= a;
    outputs(4180) <= not b or a;
    outputs(4181) <= b;
    outputs(4182) <= b;
    outputs(4183) <= b;
    outputs(4184) <= not (a xor b);
    outputs(4185) <= b and not a;
    outputs(4186) <= b and not a;
    outputs(4187) <= not (a xor b);
    outputs(4188) <= a or b;
    outputs(4189) <= not (a xor b);
    outputs(4190) <= a xor b;
    outputs(4191) <= a xor b;
    outputs(4192) <= not (a and b);
    outputs(4193) <= not a;
    outputs(4194) <= not b;
    outputs(4195) <= a and not b;
    outputs(4196) <= not (a xor b);
    outputs(4197) <= b and not a;
    outputs(4198) <= b;
    outputs(4199) <= not a;
    outputs(4200) <= a xor b;
    outputs(4201) <= a;
    outputs(4202) <= not b;
    outputs(4203) <= not a;
    outputs(4204) <= not (a xor b);
    outputs(4205) <= a and b;
    outputs(4206) <= a;
    outputs(4207) <= not (a xor b);
    outputs(4208) <= a xor b;
    outputs(4209) <= b;
    outputs(4210) <= b;
    outputs(4211) <= a;
    outputs(4212) <= not b;
    outputs(4213) <= not (a xor b);
    outputs(4214) <= not a;
    outputs(4215) <= not b;
    outputs(4216) <= b;
    outputs(4217) <= a;
    outputs(4218) <= not b;
    outputs(4219) <= a;
    outputs(4220) <= not b or a;
    outputs(4221) <= a and b;
    outputs(4222) <= a;
    outputs(4223) <= not b;
    outputs(4224) <= not (a and b);
    outputs(4225) <= not a;
    outputs(4226) <= not b;
    outputs(4227) <= not (a or b);
    outputs(4228) <= not (a or b);
    outputs(4229) <= a and not b;
    outputs(4230) <= not (a or b);
    outputs(4231) <= a and not b;
    outputs(4232) <= not a;
    outputs(4233) <= not (a xor b);
    outputs(4234) <= b;
    outputs(4235) <= a and not b;
    outputs(4236) <= not (a xor b);
    outputs(4237) <= a and b;
    outputs(4238) <= not b;
    outputs(4239) <= not b or a;
    outputs(4240) <= not b;
    outputs(4241) <= not b or a;
    outputs(4242) <= a xor b;
    outputs(4243) <= a xor b;
    outputs(4244) <= not a;
    outputs(4245) <= not a;
    outputs(4246) <= not (a xor b);
    outputs(4247) <= b;
    outputs(4248) <= a and not b;
    outputs(4249) <= a and b;
    outputs(4250) <= not a or b;
    outputs(4251) <= not b;
    outputs(4252) <= not (a xor b);
    outputs(4253) <= not (a xor b);
    outputs(4254) <= not (a xor b);
    outputs(4255) <= not (a xor b);
    outputs(4256) <= not a;
    outputs(4257) <= a and b;
    outputs(4258) <= not b;
    outputs(4259) <= b;
    outputs(4260) <= not b or a;
    outputs(4261) <= not a;
    outputs(4262) <= a xor b;
    outputs(4263) <= not (a xor b);
    outputs(4264) <= a;
    outputs(4265) <= a and b;
    outputs(4266) <= a and b;
    outputs(4267) <= a xor b;
    outputs(4268) <= a;
    outputs(4269) <= b and not a;
    outputs(4270) <= not (a xor b);
    outputs(4271) <= b;
    outputs(4272) <= a;
    outputs(4273) <= not a;
    outputs(4274) <= a and b;
    outputs(4275) <= not b or a;
    outputs(4276) <= a and not b;
    outputs(4277) <= b and not a;
    outputs(4278) <= a xor b;
    outputs(4279) <= not a;
    outputs(4280) <= b and not a;
    outputs(4281) <= not a or b;
    outputs(4282) <= not (a or b);
    outputs(4283) <= a xor b;
    outputs(4284) <= not b;
    outputs(4285) <= not a;
    outputs(4286) <= not a;
    outputs(4287) <= not a;
    outputs(4288) <= not a;
    outputs(4289) <= a and b;
    outputs(4290) <= not (a and b);
    outputs(4291) <= not (a and b);
    outputs(4292) <= not a or b;
    outputs(4293) <= not a;
    outputs(4294) <= b;
    outputs(4295) <= b and not a;
    outputs(4296) <= not (a xor b);
    outputs(4297) <= not b or a;
    outputs(4298) <= not (a xor b);
    outputs(4299) <= not (a xor b);
    outputs(4300) <= a xor b;
    outputs(4301) <= not a;
    outputs(4302) <= b;
    outputs(4303) <= not (a and b);
    outputs(4304) <= b;
    outputs(4305) <= a and not b;
    outputs(4306) <= a and b;
    outputs(4307) <= not b;
    outputs(4308) <= not a;
    outputs(4309) <= a xor b;
    outputs(4310) <= not (a xor b);
    outputs(4311) <= b;
    outputs(4312) <= a;
    outputs(4313) <= a;
    outputs(4314) <= not a or b;
    outputs(4315) <= a and b;
    outputs(4316) <= b;
    outputs(4317) <= not (a xor b);
    outputs(4318) <= a and not b;
    outputs(4319) <= not b;
    outputs(4320) <= a xor b;
    outputs(4321) <= not a or b;
    outputs(4322) <= not b;
    outputs(4323) <= not a;
    outputs(4324) <= not b;
    outputs(4325) <= a xor b;
    outputs(4326) <= a xor b;
    outputs(4327) <= not a or b;
    outputs(4328) <= not (a or b);
    outputs(4329) <= not (a xor b);
    outputs(4330) <= a;
    outputs(4331) <= a;
    outputs(4332) <= not a or b;
    outputs(4333) <= not a or b;
    outputs(4334) <= not (a xor b);
    outputs(4335) <= b;
    outputs(4336) <= a and b;
    outputs(4337) <= not a;
    outputs(4338) <= a xor b;
    outputs(4339) <= not a or b;
    outputs(4340) <= not b;
    outputs(4341) <= a xor b;
    outputs(4342) <= not a;
    outputs(4343) <= not (a xor b);
    outputs(4344) <= not a;
    outputs(4345) <= not b;
    outputs(4346) <= b;
    outputs(4347) <= not (a or b);
    outputs(4348) <= a;
    outputs(4349) <= a and b;
    outputs(4350) <= a xor b;
    outputs(4351) <= b and not a;
    outputs(4352) <= a and not b;
    outputs(4353) <= not (a xor b);
    outputs(4354) <= not b;
    outputs(4355) <= a xor b;
    outputs(4356) <= not (a xor b);
    outputs(4357) <= not a;
    outputs(4358) <= not b;
    outputs(4359) <= b;
    outputs(4360) <= not (a or b);
    outputs(4361) <= not a or b;
    outputs(4362) <= b;
    outputs(4363) <= not b;
    outputs(4364) <= not (a and b);
    outputs(4365) <= not (a and b);
    outputs(4366) <= not a;
    outputs(4367) <= a and b;
    outputs(4368) <= not a;
    outputs(4369) <= not (a and b);
    outputs(4370) <= not b or a;
    outputs(4371) <= not (a xor b);
    outputs(4372) <= not (a xor b);
    outputs(4373) <= a;
    outputs(4374) <= a and not b;
    outputs(4375) <= not a or b;
    outputs(4376) <= not (a or b);
    outputs(4377) <= not b or a;
    outputs(4378) <= not b;
    outputs(4379) <= a xor b;
    outputs(4380) <= not (a xor b);
    outputs(4381) <= not b or a;
    outputs(4382) <= not (a and b);
    outputs(4383) <= not b;
    outputs(4384) <= not a;
    outputs(4385) <= b;
    outputs(4386) <= not b;
    outputs(4387) <= b and not a;
    outputs(4388) <= a;
    outputs(4389) <= a and b;
    outputs(4390) <= not a;
    outputs(4391) <= a;
    outputs(4392) <= not (a xor b);
    outputs(4393) <= b;
    outputs(4394) <= not (a and b);
    outputs(4395) <= not a;
    outputs(4396) <= not a;
    outputs(4397) <= b;
    outputs(4398) <= a xor b;
    outputs(4399) <= not b;
    outputs(4400) <= not (a xor b);
    outputs(4401) <= not (a and b);
    outputs(4402) <= not b;
    outputs(4403) <= a and not b;
    outputs(4404) <= a and b;
    outputs(4405) <= not (a xor b);
    outputs(4406) <= b;
    outputs(4407) <= not (a xor b);
    outputs(4408) <= a and b;
    outputs(4409) <= not b;
    outputs(4410) <= a and b;
    outputs(4411) <= b and not a;
    outputs(4412) <= b and not a;
    outputs(4413) <= a xor b;
    outputs(4414) <= not (a xor b);
    outputs(4415) <= a xor b;
    outputs(4416) <= not (a xor b);
    outputs(4417) <= b and not a;
    outputs(4418) <= not (a xor b);
    outputs(4419) <= a xor b;
    outputs(4420) <= not (a xor b);
    outputs(4421) <= not a;
    outputs(4422) <= not (a xor b);
    outputs(4423) <= not b;
    outputs(4424) <= not (a xor b);
    outputs(4425) <= not (a xor b);
    outputs(4426) <= not a;
    outputs(4427) <= a;
    outputs(4428) <= not (a xor b);
    outputs(4429) <= not a;
    outputs(4430) <= not (a xor b);
    outputs(4431) <= b;
    outputs(4432) <= a and not b;
    outputs(4433) <= not (a xor b);
    outputs(4434) <= not a;
    outputs(4435) <= a and b;
    outputs(4436) <= a;
    outputs(4437) <= not b or a;
    outputs(4438) <= not a;
    outputs(4439) <= not (a xor b);
    outputs(4440) <= not (a xor b);
    outputs(4441) <= not b;
    outputs(4442) <= a xor b;
    outputs(4443) <= a and not b;
    outputs(4444) <= b and not a;
    outputs(4445) <= a xor b;
    outputs(4446) <= not (a xor b);
    outputs(4447) <= a xor b;
    outputs(4448) <= a xor b;
    outputs(4449) <= a;
    outputs(4450) <= not (a xor b);
    outputs(4451) <= not a;
    outputs(4452) <= a xor b;
    outputs(4453) <= a xor b;
    outputs(4454) <= not a or b;
    outputs(4455) <= a;
    outputs(4456) <= not a;
    outputs(4457) <= a and not b;
    outputs(4458) <= not a;
    outputs(4459) <= not (a xor b);
    outputs(4460) <= a;
    outputs(4461) <= a;
    outputs(4462) <= not a;
    outputs(4463) <= not b;
    outputs(4464) <= a or b;
    outputs(4465) <= a and b;
    outputs(4466) <= not (a xor b);
    outputs(4467) <= a xor b;
    outputs(4468) <= not a;
    outputs(4469) <= not b or a;
    outputs(4470) <= a and b;
    outputs(4471) <= a;
    outputs(4472) <= a and not b;
    outputs(4473) <= not (a or b);
    outputs(4474) <= not (a and b);
    outputs(4475) <= a or b;
    outputs(4476) <= not b or a;
    outputs(4477) <= not (a xor b);
    outputs(4478) <= a xor b;
    outputs(4479) <= a;
    outputs(4480) <= a xor b;
    outputs(4481) <= not (a xor b);
    outputs(4482) <= not a or b;
    outputs(4483) <= a or b;
    outputs(4484) <= not (a or b);
    outputs(4485) <= b and not a;
    outputs(4486) <= b;
    outputs(4487) <= a;
    outputs(4488) <= a xor b;
    outputs(4489) <= b;
    outputs(4490) <= a and not b;
    outputs(4491) <= b;
    outputs(4492) <= not a;
    outputs(4493) <= a xor b;
    outputs(4494) <= not a;
    outputs(4495) <= b;
    outputs(4496) <= b;
    outputs(4497) <= a;
    outputs(4498) <= a xor b;
    outputs(4499) <= not b or a;
    outputs(4500) <= b;
    outputs(4501) <= not (a or b);
    outputs(4502) <= b and not a;
    outputs(4503) <= a;
    outputs(4504) <= not (a xor b);
    outputs(4505) <= a or b;
    outputs(4506) <= not a;
    outputs(4507) <= b and not a;
    outputs(4508) <= not b;
    outputs(4509) <= not (a xor b);
    outputs(4510) <= not (a xor b);
    outputs(4511) <= a xor b;
    outputs(4512) <= b;
    outputs(4513) <= a xor b;
    outputs(4514) <= a;
    outputs(4515) <= a;
    outputs(4516) <= not a;
    outputs(4517) <= a or b;
    outputs(4518) <= a and b;
    outputs(4519) <= a and b;
    outputs(4520) <= not (a or b);
    outputs(4521) <= a and b;
    outputs(4522) <= not b or a;
    outputs(4523) <= not b;
    outputs(4524) <= b;
    outputs(4525) <= not (a xor b);
    outputs(4526) <= a and b;
    outputs(4527) <= not (a xor b);
    outputs(4528) <= a xor b;
    outputs(4529) <= not b;
    outputs(4530) <= a xor b;
    outputs(4531) <= a and b;
    outputs(4532) <= a xor b;
    outputs(4533) <= not a;
    outputs(4534) <= a xor b;
    outputs(4535) <= not (a xor b);
    outputs(4536) <= b;
    outputs(4537) <= not (a xor b);
    outputs(4538) <= not b or a;
    outputs(4539) <= a xor b;
    outputs(4540) <= a and b;
    outputs(4541) <= a;
    outputs(4542) <= a and b;
    outputs(4543) <= a xor b;
    outputs(4544) <= a xor b;
    outputs(4545) <= b;
    outputs(4546) <= b;
    outputs(4547) <= b and not a;
    outputs(4548) <= a xor b;
    outputs(4549) <= b and not a;
    outputs(4550) <= a;
    outputs(4551) <= a xor b;
    outputs(4552) <= a xor b;
    outputs(4553) <= b;
    outputs(4554) <= a xor b;
    outputs(4555) <= not b or a;
    outputs(4556) <= not (a xor b);
    outputs(4557) <= b;
    outputs(4558) <= a;
    outputs(4559) <= not b;
    outputs(4560) <= not (a xor b);
    outputs(4561) <= not b;
    outputs(4562) <= b;
    outputs(4563) <= a xor b;
    outputs(4564) <= not b or a;
    outputs(4565) <= not b or a;
    outputs(4566) <= not (a and b);
    outputs(4567) <= a xor b;
    outputs(4568) <= a xor b;
    outputs(4569) <= not a or b;
    outputs(4570) <= a or b;
    outputs(4571) <= not b;
    outputs(4572) <= not (a xor b);
    outputs(4573) <= a or b;
    outputs(4574) <= a;
    outputs(4575) <= a xor b;
    outputs(4576) <= not (a xor b);
    outputs(4577) <= b;
    outputs(4578) <= b;
    outputs(4579) <= b;
    outputs(4580) <= b;
    outputs(4581) <= not a;
    outputs(4582) <= not (a xor b);
    outputs(4583) <= not (a xor b);
    outputs(4584) <= not a;
    outputs(4585) <= not a;
    outputs(4586) <= a xor b;
    outputs(4587) <= not a;
    outputs(4588) <= b and not a;
    outputs(4589) <= not (a and b);
    outputs(4590) <= b;
    outputs(4591) <= not b or a;
    outputs(4592) <= a and b;
    outputs(4593) <= a and b;
    outputs(4594) <= not (a xor b);
    outputs(4595) <= not (a xor b);
    outputs(4596) <= not (a xor b);
    outputs(4597) <= not b or a;
    outputs(4598) <= a xor b;
    outputs(4599) <= not a;
    outputs(4600) <= a and not b;
    outputs(4601) <= not b;
    outputs(4602) <= a xor b;
    outputs(4603) <= a;
    outputs(4604) <= b and not a;
    outputs(4605) <= a xor b;
    outputs(4606) <= not a;
    outputs(4607) <= a and b;
    outputs(4608) <= a and b;
    outputs(4609) <= b and not a;
    outputs(4610) <= not (a or b);
    outputs(4611) <= not a;
    outputs(4612) <= not b;
    outputs(4613) <= not a;
    outputs(4614) <= not (a xor b);
    outputs(4615) <= b and not a;
    outputs(4616) <= b;
    outputs(4617) <= not (a or b);
    outputs(4618) <= not a;
    outputs(4619) <= not (a xor b);
    outputs(4620) <= b;
    outputs(4621) <= a xor b;
    outputs(4622) <= not b;
    outputs(4623) <= not a;
    outputs(4624) <= a;
    outputs(4625) <= not (a xor b);
    outputs(4626) <= a and b;
    outputs(4627) <= b;
    outputs(4628) <= not a;
    outputs(4629) <= b;
    outputs(4630) <= not b;
    outputs(4631) <= b;
    outputs(4632) <= a and b;
    outputs(4633) <= not a;
    outputs(4634) <= not (a or b);
    outputs(4635) <= b;
    outputs(4636) <= b;
    outputs(4637) <= a xor b;
    outputs(4638) <= not (a and b);
    outputs(4639) <= not b;
    outputs(4640) <= not b or a;
    outputs(4641) <= not b;
    outputs(4642) <= b;
    outputs(4643) <= a xor b;
    outputs(4644) <= not a;
    outputs(4645) <= not a;
    outputs(4646) <= not a or b;
    outputs(4647) <= a;
    outputs(4648) <= not a;
    outputs(4649) <= a and not b;
    outputs(4650) <= a and not b;
    outputs(4651) <= b and not a;
    outputs(4652) <= a;
    outputs(4653) <= not (a xor b);
    outputs(4654) <= not b;
    outputs(4655) <= b and not a;
    outputs(4656) <= a xor b;
    outputs(4657) <= a;
    outputs(4658) <= b and not a;
    outputs(4659) <= a xor b;
    outputs(4660) <= a and not b;
    outputs(4661) <= b;
    outputs(4662) <= not b;
    outputs(4663) <= b;
    outputs(4664) <= not a;
    outputs(4665) <= a xor b;
    outputs(4666) <= a;
    outputs(4667) <= not (a xor b);
    outputs(4668) <= b and not a;
    outputs(4669) <= not a or b;
    outputs(4670) <= not (a xor b);
    outputs(4671) <= b;
    outputs(4672) <= b;
    outputs(4673) <= a;
    outputs(4674) <= not (a xor b);
    outputs(4675) <= b;
    outputs(4676) <= a;
    outputs(4677) <= not (a and b);
    outputs(4678) <= a;
    outputs(4679) <= not (a xor b);
    outputs(4680) <= b and not a;
    outputs(4681) <= not (a and b);
    outputs(4682) <= not (a xor b);
    outputs(4683) <= not (a or b);
    outputs(4684) <= a;
    outputs(4685) <= not a;
    outputs(4686) <= not b or a;
    outputs(4687) <= not a;
    outputs(4688) <= a;
    outputs(4689) <= a and not b;
    outputs(4690) <= not b;
    outputs(4691) <= a and b;
    outputs(4692) <= a and not b;
    outputs(4693) <= not b;
    outputs(4694) <= not (a or b);
    outputs(4695) <= not a;
    outputs(4696) <= a;
    outputs(4697) <= a and not b;
    outputs(4698) <= a and not b;
    outputs(4699) <= not a or b;
    outputs(4700) <= a;
    outputs(4701) <= a xor b;
    outputs(4702) <= a and b;
    outputs(4703) <= b and not a;
    outputs(4704) <= not (a and b);
    outputs(4705) <= a xor b;
    outputs(4706) <= b;
    outputs(4707) <= not (a or b);
    outputs(4708) <= a;
    outputs(4709) <= not b;
    outputs(4710) <= a;
    outputs(4711) <= not a;
    outputs(4712) <= a;
    outputs(4713) <= a and b;
    outputs(4714) <= b;
    outputs(4715) <= a and b;
    outputs(4716) <= not a;
    outputs(4717) <= not (a xor b);
    outputs(4718) <= a;
    outputs(4719) <= a;
    outputs(4720) <= not b;
    outputs(4721) <= b;
    outputs(4722) <= not (a or b);
    outputs(4723) <= not (a xor b);
    outputs(4724) <= b and not a;
    outputs(4725) <= a xor b;
    outputs(4726) <= a and not b;
    outputs(4727) <= b;
    outputs(4728) <= not a;
    outputs(4729) <= not b;
    outputs(4730) <= b and not a;
    outputs(4731) <= a and b;
    outputs(4732) <= a xor b;
    outputs(4733) <= a xor b;
    outputs(4734) <= not a;
    outputs(4735) <= not b;
    outputs(4736) <= b and not a;
    outputs(4737) <= not (a xor b);
    outputs(4738) <= a;
    outputs(4739) <= b;
    outputs(4740) <= b;
    outputs(4741) <= not a;
    outputs(4742) <= a xor b;
    outputs(4743) <= a and not b;
    outputs(4744) <= b and not a;
    outputs(4745) <= a and not b;
    outputs(4746) <= b;
    outputs(4747) <= not (a xor b);
    outputs(4748) <= not (a xor b);
    outputs(4749) <= a;
    outputs(4750) <= not a;
    outputs(4751) <= not a;
    outputs(4752) <= not b;
    outputs(4753) <= a xor b;
    outputs(4754) <= not a or b;
    outputs(4755) <= a;
    outputs(4756) <= b;
    outputs(4757) <= a;
    outputs(4758) <= a xor b;
    outputs(4759) <= b;
    outputs(4760) <= not (a or b);
    outputs(4761) <= not (a xor b);
    outputs(4762) <= not (a and b);
    outputs(4763) <= a xor b;
    outputs(4764) <= b;
    outputs(4765) <= a;
    outputs(4766) <= not b or a;
    outputs(4767) <= not (a or b);
    outputs(4768) <= a and b;
    outputs(4769) <= a;
    outputs(4770) <= not b;
    outputs(4771) <= not (a xor b);
    outputs(4772) <= a xor b;
    outputs(4773) <= not a;
    outputs(4774) <= not (a xor b);
    outputs(4775) <= not b or a;
    outputs(4776) <= a xor b;
    outputs(4777) <= a;
    outputs(4778) <= a and b;
    outputs(4779) <= not (a xor b);
    outputs(4780) <= not a;
    outputs(4781) <= not (a or b);
    outputs(4782) <= a;
    outputs(4783) <= not a;
    outputs(4784) <= not (a xor b);
    outputs(4785) <= not a;
    outputs(4786) <= not (a xor b);
    outputs(4787) <= b;
    outputs(4788) <= not b;
    outputs(4789) <= not a;
    outputs(4790) <= not (a xor b);
    outputs(4791) <= not a;
    outputs(4792) <= a and not b;
    outputs(4793) <= not b;
    outputs(4794) <= not (a and b);
    outputs(4795) <= b;
    outputs(4796) <= b;
    outputs(4797) <= b and not a;
    outputs(4798) <= not (a xor b);
    outputs(4799) <= a and b;
    outputs(4800) <= not b or a;
    outputs(4801) <= not (a and b);
    outputs(4802) <= not (a or b);
    outputs(4803) <= a xor b;
    outputs(4804) <= not (a xor b);
    outputs(4805) <= 1'b0;
    outputs(4806) <= not a;
    outputs(4807) <= not a;
    outputs(4808) <= a and b;
    outputs(4809) <= not (a xor b);
    outputs(4810) <= a and not b;
    outputs(4811) <= not (a xor b);
    outputs(4812) <= not b;
    outputs(4813) <= a or b;
    outputs(4814) <= a or b;
    outputs(4815) <= a and not b;
    outputs(4816) <= b;
    outputs(4817) <= b;
    outputs(4818) <= a xor b;
    outputs(4819) <= not a;
    outputs(4820) <= not b;
    outputs(4821) <= a and not b;
    outputs(4822) <= not (a xor b);
    outputs(4823) <= a and b;
    outputs(4824) <= b and not a;
    outputs(4825) <= not (a xor b);
    outputs(4826) <= b;
    outputs(4827) <= a or b;
    outputs(4828) <= not (a xor b);
    outputs(4829) <= not b or a;
    outputs(4830) <= not b;
    outputs(4831) <= not b or a;
    outputs(4832) <= a xor b;
    outputs(4833) <= not (a xor b);
    outputs(4834) <= b;
    outputs(4835) <= a and not b;
    outputs(4836) <= b;
    outputs(4837) <= a xor b;
    outputs(4838) <= not (a or b);
    outputs(4839) <= not (a or b);
    outputs(4840) <= b;
    outputs(4841) <= not (a or b);
    outputs(4842) <= b and not a;
    outputs(4843) <= a and not b;
    outputs(4844) <= b and not a;
    outputs(4845) <= b;
    outputs(4846) <= a xor b;
    outputs(4847) <= a;
    outputs(4848) <= a;
    outputs(4849) <= b;
    outputs(4850) <= b and not a;
    outputs(4851) <= not a or b;
    outputs(4852) <= b;
    outputs(4853) <= b and not a;
    outputs(4854) <= a;
    outputs(4855) <= b;
    outputs(4856) <= not (a xor b);
    outputs(4857) <= not (a xor b);
    outputs(4858) <= a;
    outputs(4859) <= not b;
    outputs(4860) <= b and not a;
    outputs(4861) <= a or b;
    outputs(4862) <= a or b;
    outputs(4863) <= not (a xor b);
    outputs(4864) <= a and not b;
    outputs(4865) <= b;
    outputs(4866) <= not (a or b);
    outputs(4867) <= b;
    outputs(4868) <= not a;
    outputs(4869) <= not a;
    outputs(4870) <= b;
    outputs(4871) <= a and b;
    outputs(4872) <= not (a xor b);
    outputs(4873) <= not (a and b);
    outputs(4874) <= not (a and b);
    outputs(4875) <= a and not b;
    outputs(4876) <= a and b;
    outputs(4877) <= not (a xor b);
    outputs(4878) <= a;
    outputs(4879) <= b;
    outputs(4880) <= not (a xor b);
    outputs(4881) <= a and not b;
    outputs(4882) <= a xor b;
    outputs(4883) <= not (a and b);
    outputs(4884) <= a and b;
    outputs(4885) <= b and not a;
    outputs(4886) <= b;
    outputs(4887) <= b;
    outputs(4888) <= not (a xor b);
    outputs(4889) <= not (a or b);
    outputs(4890) <= b;
    outputs(4891) <= a and not b;
    outputs(4892) <= b and not a;
    outputs(4893) <= not (a xor b);
    outputs(4894) <= a and not b;
    outputs(4895) <= a or b;
    outputs(4896) <= not b;
    outputs(4897) <= not b;
    outputs(4898) <= a;
    outputs(4899) <= a xor b;
    outputs(4900) <= a xor b;
    outputs(4901) <= b and not a;
    outputs(4902) <= not (a or b);
    outputs(4903) <= a xor b;
    outputs(4904) <= b;
    outputs(4905) <= not b;
    outputs(4906) <= a xor b;
    outputs(4907) <= a;
    outputs(4908) <= a and not b;
    outputs(4909) <= not b;
    outputs(4910) <= not a;
    outputs(4911) <= b and not a;
    outputs(4912) <= b;
    outputs(4913) <= b;
    outputs(4914) <= b;
    outputs(4915) <= b and not a;
    outputs(4916) <= a and not b;
    outputs(4917) <= not (a xor b);
    outputs(4918) <= not (a xor b);
    outputs(4919) <= not (a xor b);
    outputs(4920) <= not (a xor b);
    outputs(4921) <= not (a or b);
    outputs(4922) <= not a;
    outputs(4923) <= not b;
    outputs(4924) <= a and not b;
    outputs(4925) <= not a;
    outputs(4926) <= b and not a;
    outputs(4927) <= not a;
    outputs(4928) <= b;
    outputs(4929) <= a xor b;
    outputs(4930) <= a;
    outputs(4931) <= not (a xor b);
    outputs(4932) <= not b;
    outputs(4933) <= not b;
    outputs(4934) <= b;
    outputs(4935) <= not b;
    outputs(4936) <= not b;
    outputs(4937) <= not b;
    outputs(4938) <= a;
    outputs(4939) <= not a;
    outputs(4940) <= not b;
    outputs(4941) <= a and b;
    outputs(4942) <= not a or b;
    outputs(4943) <= b;
    outputs(4944) <= not (a xor b);
    outputs(4945) <= not a;
    outputs(4946) <= a xor b;
    outputs(4947) <= a;
    outputs(4948) <= not (a or b);
    outputs(4949) <= not (a or b);
    outputs(4950) <= a or b;
    outputs(4951) <= a and not b;
    outputs(4952) <= b;
    outputs(4953) <= not (a xor b);
    outputs(4954) <= not (a and b);
    outputs(4955) <= a or b;
    outputs(4956) <= not b;
    outputs(4957) <= not a;
    outputs(4958) <= not a;
    outputs(4959) <= not (a xor b);
    outputs(4960) <= not b or a;
    outputs(4961) <= not a;
    outputs(4962) <= b;
    outputs(4963) <= a xor b;
    outputs(4964) <= a and b;
    outputs(4965) <= a;
    outputs(4966) <= a xor b;
    outputs(4967) <= not a;
    outputs(4968) <= not (a and b);
    outputs(4969) <= not b or a;
    outputs(4970) <= not (a and b);
    outputs(4971) <= not a;
    outputs(4972) <= b;
    outputs(4973) <= not a;
    outputs(4974) <= not a;
    outputs(4975) <= a or b;
    outputs(4976) <= not (a xor b);
    outputs(4977) <= not b;
    outputs(4978) <= not b or a;
    outputs(4979) <= b;
    outputs(4980) <= b;
    outputs(4981) <= not b or a;
    outputs(4982) <= a and b;
    outputs(4983) <= not (a xor b);
    outputs(4984) <= a xor b;
    outputs(4985) <= a;
    outputs(4986) <= b;
    outputs(4987) <= not b;
    outputs(4988) <= a and not b;
    outputs(4989) <= not (a or b);
    outputs(4990) <= not a;
    outputs(4991) <= b;
    outputs(4992) <= b and not a;
    outputs(4993) <= not b;
    outputs(4994) <= not b;
    outputs(4995) <= not a;
    outputs(4996) <= not (a xor b);
    outputs(4997) <= a and not b;
    outputs(4998) <= not (a xor b);
    outputs(4999) <= not a;
    outputs(5000) <= not (a xor b);
    outputs(5001) <= a;
    outputs(5002) <= not b;
    outputs(5003) <= not (a xor b);
    outputs(5004) <= not a;
    outputs(5005) <= a;
    outputs(5006) <= a or b;
    outputs(5007) <= b;
    outputs(5008) <= not (a xor b);
    outputs(5009) <= not b or a;
    outputs(5010) <= not b;
    outputs(5011) <= a xor b;
    outputs(5012) <= not (a and b);
    outputs(5013) <= a;
    outputs(5014) <= not (a xor b);
    outputs(5015) <= b;
    outputs(5016) <= a;
    outputs(5017) <= not (a or b);
    outputs(5018) <= a and b;
    outputs(5019) <= b;
    outputs(5020) <= b;
    outputs(5021) <= a and b;
    outputs(5022) <= a;
    outputs(5023) <= a xor b;
    outputs(5024) <= a and not b;
    outputs(5025) <= b;
    outputs(5026) <= b and not a;
    outputs(5027) <= not (a xor b);
    outputs(5028) <= b;
    outputs(5029) <= a and not b;
    outputs(5030) <= not (a or b);
    outputs(5031) <= a and b;
    outputs(5032) <= b;
    outputs(5033) <= not a;
    outputs(5034) <= a or b;
    outputs(5035) <= not a or b;
    outputs(5036) <= not (a xor b);
    outputs(5037) <= not b;
    outputs(5038) <= a and not b;
    outputs(5039) <= not (a or b);
    outputs(5040) <= a and b;
    outputs(5041) <= b and not a;
    outputs(5042) <= not a or b;
    outputs(5043) <= not (a and b);
    outputs(5044) <= a xor b;
    outputs(5045) <= a;
    outputs(5046) <= not (a and b);
    outputs(5047) <= not (a or b);
    outputs(5048) <= not (a xor b);
    outputs(5049) <= not (a or b);
    outputs(5050) <= a;
    outputs(5051) <= a and b;
    outputs(5052) <= a and b;
    outputs(5053) <= b and not a;
    outputs(5054) <= b;
    outputs(5055) <= a and b;
    outputs(5056) <= a xor b;
    outputs(5057) <= not (a xor b);
    outputs(5058) <= b;
    outputs(5059) <= not a;
    outputs(5060) <= a xor b;
    outputs(5061) <= not (a and b);
    outputs(5062) <= a and b;
    outputs(5063) <= not b;
    outputs(5064) <= not a;
    outputs(5065) <= a xor b;
    outputs(5066) <= a xor b;
    outputs(5067) <= b;
    outputs(5068) <= a xor b;
    outputs(5069) <= not (a or b);
    outputs(5070) <= a;
    outputs(5071) <= not b;
    outputs(5072) <= a xor b;
    outputs(5073) <= not a;
    outputs(5074) <= a and not b;
    outputs(5075) <= a xor b;
    outputs(5076) <= a;
    outputs(5077) <= b;
    outputs(5078) <= a;
    outputs(5079) <= not b;
    outputs(5080) <= b and not a;
    outputs(5081) <= a;
    outputs(5082) <= not b;
    outputs(5083) <= not b or a;
    outputs(5084) <= a;
    outputs(5085) <= b;
    outputs(5086) <= not a or b;
    outputs(5087) <= not b;
    outputs(5088) <= b and not a;
    outputs(5089) <= a and b;
    outputs(5090) <= a xor b;
    outputs(5091) <= not (a xor b);
    outputs(5092) <= a and b;
    outputs(5093) <= a;
    outputs(5094) <= not (a or b);
    outputs(5095) <= b;
    outputs(5096) <= a xor b;
    outputs(5097) <= not (a xor b);
    outputs(5098) <= b;
    outputs(5099) <= b;
    outputs(5100) <= b and not a;
    outputs(5101) <= a xor b;
    outputs(5102) <= a xor b;
    outputs(5103) <= b and not a;
    outputs(5104) <= a;
    outputs(5105) <= a xor b;
    outputs(5106) <= not b;
    outputs(5107) <= a and not b;
    outputs(5108) <= not b;
    outputs(5109) <= a and not b;
    outputs(5110) <= a xor b;
    outputs(5111) <= b and not a;
    outputs(5112) <= b;
    outputs(5113) <= a or b;
    outputs(5114) <= b and not a;
    outputs(5115) <= not (a xor b);
    outputs(5116) <= not (a and b);
    outputs(5117) <= b and not a;
    outputs(5118) <= a;
    outputs(5119) <= not (a xor b);
    outputs(5120) <= a;
    outputs(5121) <= a and not b;
    outputs(5122) <= not b;
    outputs(5123) <= not (a xor b);
    outputs(5124) <= a and not b;
    outputs(5125) <= a xor b;
    outputs(5126) <= a;
    outputs(5127) <= not a;
    outputs(5128) <= not a;
    outputs(5129) <= not a;
    outputs(5130) <= not b;
    outputs(5131) <= not (a xor b);
    outputs(5132) <= not (a or b);
    outputs(5133) <= not (a and b);
    outputs(5134) <= a;
    outputs(5135) <= not a;
    outputs(5136) <= not (a or b);
    outputs(5137) <= not (a xor b);
    outputs(5138) <= a and b;
    outputs(5139) <= not b;
    outputs(5140) <= not (a or b);
    outputs(5141) <= a;
    outputs(5142) <= not (a xor b);
    outputs(5143) <= b;
    outputs(5144) <= a and not b;
    outputs(5145) <= not (a xor b);
    outputs(5146) <= not (a xor b);
    outputs(5147) <= b and not a;
    outputs(5148) <= a xor b;
    outputs(5149) <= not b;
    outputs(5150) <= not (a or b);
    outputs(5151) <= not a;
    outputs(5152) <= b and not a;
    outputs(5153) <= b;
    outputs(5154) <= a;
    outputs(5155) <= not (a xor b);
    outputs(5156) <= a xor b;
    outputs(5157) <= a;
    outputs(5158) <= not b;
    outputs(5159) <= a xor b;
    outputs(5160) <= not (a or b);
    outputs(5161) <= not a;
    outputs(5162) <= b;
    outputs(5163) <= not (a and b);
    outputs(5164) <= a and b;
    outputs(5165) <= not b or a;
    outputs(5166) <= b;
    outputs(5167) <= not a;
    outputs(5168) <= a and not b;
    outputs(5169) <= a;
    outputs(5170) <= a;
    outputs(5171) <= not a;
    outputs(5172) <= not a;
    outputs(5173) <= not b;
    outputs(5174) <= not (a or b);
    outputs(5175) <= not (a and b);
    outputs(5176) <= not (a or b);
    outputs(5177) <= not a;
    outputs(5178) <= not b or a;
    outputs(5179) <= a;
    outputs(5180) <= not a or b;
    outputs(5181) <= not b or a;
    outputs(5182) <= not (a xor b);
    outputs(5183) <= b;
    outputs(5184) <= not a;
    outputs(5185) <= a xor b;
    outputs(5186) <= not a;
    outputs(5187) <= not b;
    outputs(5188) <= not b;
    outputs(5189) <= a;
    outputs(5190) <= not a;
    outputs(5191) <= not (a xor b);
    outputs(5192) <= not (a xor b);
    outputs(5193) <= not b;
    outputs(5194) <= not a;
    outputs(5195) <= b;
    outputs(5196) <= not (a xor b);
    outputs(5197) <= not (a xor b);
    outputs(5198) <= b;
    outputs(5199) <= a;
    outputs(5200) <= not (a or b);
    outputs(5201) <= a and b;
    outputs(5202) <= b;
    outputs(5203) <= a and b;
    outputs(5204) <= a;
    outputs(5205) <= a xor b;
    outputs(5206) <= a and not b;
    outputs(5207) <= a and not b;
    outputs(5208) <= b;
    outputs(5209) <= not b or a;
    outputs(5210) <= not b;
    outputs(5211) <= a and b;
    outputs(5212) <= a;
    outputs(5213) <= not (a or b);
    outputs(5214) <= not b or a;
    outputs(5215) <= a and not b;
    outputs(5216) <= not (a xor b);
    outputs(5217) <= not a;
    outputs(5218) <= not b;
    outputs(5219) <= b and not a;
    outputs(5220) <= b;
    outputs(5221) <= not (a and b);
    outputs(5222) <= a xor b;
    outputs(5223) <= b and not a;
    outputs(5224) <= b;
    outputs(5225) <= a and b;
    outputs(5226) <= a xor b;
    outputs(5227) <= a xor b;
    outputs(5228) <= not (a xor b);
    outputs(5229) <= b;
    outputs(5230) <= a and not b;
    outputs(5231) <= a;
    outputs(5232) <= b;
    outputs(5233) <= a and b;
    outputs(5234) <= not b;
    outputs(5235) <= b;
    outputs(5236) <= b and not a;
    outputs(5237) <= not (a or b);
    outputs(5238) <= not (a xor b);
    outputs(5239) <= b;
    outputs(5240) <= a xor b;
    outputs(5241) <= not a;
    outputs(5242) <= not b;
    outputs(5243) <= not a;
    outputs(5244) <= not (a xor b);
    outputs(5245) <= not (a and b);
    outputs(5246) <= not b;
    outputs(5247) <= a;
    outputs(5248) <= not a;
    outputs(5249) <= not (a or b);
    outputs(5250) <= a;
    outputs(5251) <= a xor b;
    outputs(5252) <= b;
    outputs(5253) <= not (a xor b);
    outputs(5254) <= a xor b;
    outputs(5255) <= a;
    outputs(5256) <= not b;
    outputs(5257) <= a xor b;
    outputs(5258) <= a xor b;
    outputs(5259) <= a;
    outputs(5260) <= not b;
    outputs(5261) <= not b or a;
    outputs(5262) <= a and not b;
    outputs(5263) <= a;
    outputs(5264) <= not (a xor b);
    outputs(5265) <= a and b;
    outputs(5266) <= a xor b;
    outputs(5267) <= not b;
    outputs(5268) <= b and not a;
    outputs(5269) <= b;
    outputs(5270) <= not (a or b);
    outputs(5271) <= not (a xor b);
    outputs(5272) <= not b;
    outputs(5273) <= b and not a;
    outputs(5274) <= a xor b;
    outputs(5275) <= not a;
    outputs(5276) <= not (a or b);
    outputs(5277) <= b and not a;
    outputs(5278) <= not (a xor b);
    outputs(5279) <= a xor b;
    outputs(5280) <= b;
    outputs(5281) <= not b or a;
    outputs(5282) <= a xor b;
    outputs(5283) <= not (a or b);
    outputs(5284) <= not b;
    outputs(5285) <= a and b;
    outputs(5286) <= a xor b;
    outputs(5287) <= not a or b;
    outputs(5288) <= not (a or b);
    outputs(5289) <= not (a xor b);
    outputs(5290) <= a;
    outputs(5291) <= not b;
    outputs(5292) <= a;
    outputs(5293) <= a and not b;
    outputs(5294) <= b and not a;
    outputs(5295) <= a or b;
    outputs(5296) <= a or b;
    outputs(5297) <= not (a and b);
    outputs(5298) <= a;
    outputs(5299) <= b and not a;
    outputs(5300) <= b;
    outputs(5301) <= b and not a;
    outputs(5302) <= not (a xor b);
    outputs(5303) <= b and not a;
    outputs(5304) <= not b;
    outputs(5305) <= not b;
    outputs(5306) <= b;
    outputs(5307) <= not b;
    outputs(5308) <= a xor b;
    outputs(5309) <= a and b;
    outputs(5310) <= a xor b;
    outputs(5311) <= a and b;
    outputs(5312) <= a or b;
    outputs(5313) <= a and not b;
    outputs(5314) <= not a;
    outputs(5315) <= not (a xor b);
    outputs(5316) <= b;
    outputs(5317) <= a;
    outputs(5318) <= a and b;
    outputs(5319) <= a xor b;
    outputs(5320) <= b;
    outputs(5321) <= not (a xor b);
    outputs(5322) <= not a;
    outputs(5323) <= a and not b;
    outputs(5324) <= not b or a;
    outputs(5325) <= b and not a;
    outputs(5326) <= not a;
    outputs(5327) <= not a;
    outputs(5328) <= a and not b;
    outputs(5329) <= a xor b;
    outputs(5330) <= not b;
    outputs(5331) <= a xor b;
    outputs(5332) <= not b;
    outputs(5333) <= a and not b;
    outputs(5334) <= not (a or b);
    outputs(5335) <= a xor b;
    outputs(5336) <= not b;
    outputs(5337) <= b;
    outputs(5338) <= not (a xor b);
    outputs(5339) <= not b;
    outputs(5340) <= not a;
    outputs(5341) <= a and b;
    outputs(5342) <= not (a or b);
    outputs(5343) <= not b;
    outputs(5344) <= not a;
    outputs(5345) <= not a;
    outputs(5346) <= not b or a;
    outputs(5347) <= not a;
    outputs(5348) <= not b or a;
    outputs(5349) <= b;
    outputs(5350) <= not (a and b);
    outputs(5351) <= not a;
    outputs(5352) <= b and not a;
    outputs(5353) <= a or b;
    outputs(5354) <= a;
    outputs(5355) <= a and not b;
    outputs(5356) <= not a;
    outputs(5357) <= b;
    outputs(5358) <= a and not b;
    outputs(5359) <= a;
    outputs(5360) <= a xor b;
    outputs(5361) <= a;
    outputs(5362) <= a;
    outputs(5363) <= not a;
    outputs(5364) <= not a or b;
    outputs(5365) <= a;
    outputs(5366) <= a or b;
    outputs(5367) <= a;
    outputs(5368) <= a xor b;
    outputs(5369) <= b;
    outputs(5370) <= a xor b;
    outputs(5371) <= not a;
    outputs(5372) <= b and not a;
    outputs(5373) <= not b;
    outputs(5374) <= not (a xor b);
    outputs(5375) <= not b or a;
    outputs(5376) <= b and not a;
    outputs(5377) <= a and b;
    outputs(5378) <= not a;
    outputs(5379) <= not (a xor b);
    outputs(5380) <= not (a xor b);
    outputs(5381) <= not a or b;
    outputs(5382) <= a and not b;
    outputs(5383) <= not b or a;
    outputs(5384) <= b and not a;
    outputs(5385) <= a and b;
    outputs(5386) <= not a;
    outputs(5387) <= not a;
    outputs(5388) <= not b;
    outputs(5389) <= not (a xor b);
    outputs(5390) <= not a;
    outputs(5391) <= not (a or b);
    outputs(5392) <= a xor b;
    outputs(5393) <= b;
    outputs(5394) <= a and not b;
    outputs(5395) <= a;
    outputs(5396) <= b;
    outputs(5397) <= a;
    outputs(5398) <= not (a xor b);
    outputs(5399) <= not a;
    outputs(5400) <= a;
    outputs(5401) <= b;
    outputs(5402) <= b and not a;
    outputs(5403) <= a;
    outputs(5404) <= b;
    outputs(5405) <= not (a or b);
    outputs(5406) <= a or b;
    outputs(5407) <= not b;
    outputs(5408) <= not (a xor b);
    outputs(5409) <= a xor b;
    outputs(5410) <= a xor b;
    outputs(5411) <= not (a xor b);
    outputs(5412) <= not (a and b);
    outputs(5413) <= a;
    outputs(5414) <= not a;
    outputs(5415) <= not b;
    outputs(5416) <= a xor b;
    outputs(5417) <= not a;
    outputs(5418) <= a and b;
    outputs(5419) <= not b;
    outputs(5420) <= not b or a;
    outputs(5421) <= not (a or b);
    outputs(5422) <= b;
    outputs(5423) <= not (a or b);
    outputs(5424) <= a and b;
    outputs(5425) <= b and not a;
    outputs(5426) <= not (a xor b);
    outputs(5427) <= not b;
    outputs(5428) <= not a;
    outputs(5429) <= a xor b;
    outputs(5430) <= b;
    outputs(5431) <= not (a xor b);
    outputs(5432) <= not b or a;
    outputs(5433) <= a and not b;
    outputs(5434) <= not b or a;
    outputs(5435) <= not b;
    outputs(5436) <= a xor b;
    outputs(5437) <= a or b;
    outputs(5438) <= b;
    outputs(5439) <= not a;
    outputs(5440) <= not a;
    outputs(5441) <= a and b;
    outputs(5442) <= a and not b;
    outputs(5443) <= not a;
    outputs(5444) <= not a;
    outputs(5445) <= a;
    outputs(5446) <= a xor b;
    outputs(5447) <= a;
    outputs(5448) <= not b;
    outputs(5449) <= a;
    outputs(5450) <= b and not a;
    outputs(5451) <= a and b;
    outputs(5452) <= b;
    outputs(5453) <= b and not a;
    outputs(5454) <= b;
    outputs(5455) <= a xor b;
    outputs(5456) <= not a;
    outputs(5457) <= a xor b;
    outputs(5458) <= a and not b;
    outputs(5459) <= not a;
    outputs(5460) <= b and not a;
    outputs(5461) <= not a;
    outputs(5462) <= a xor b;
    outputs(5463) <= a xor b;
    outputs(5464) <= b;
    outputs(5465) <= a and not b;
    outputs(5466) <= a xor b;
    outputs(5467) <= not b or a;
    outputs(5468) <= not a;
    outputs(5469) <= a;
    outputs(5470) <= not a;
    outputs(5471) <= not (a xor b);
    outputs(5472) <= b;
    outputs(5473) <= not a;
    outputs(5474) <= not (a or b);
    outputs(5475) <= b;
    outputs(5476) <= a and b;
    outputs(5477) <= not (a xor b);
    outputs(5478) <= a and not b;
    outputs(5479) <= a;
    outputs(5480) <= not a;
    outputs(5481) <= not (a xor b);
    outputs(5482) <= a;
    outputs(5483) <= a and b;
    outputs(5484) <= a xor b;
    outputs(5485) <= a;
    outputs(5486) <= a and not b;
    outputs(5487) <= a and b;
    outputs(5488) <= not (a xor b);
    outputs(5489) <= a or b;
    outputs(5490) <= not a;
    outputs(5491) <= b;
    outputs(5492) <= not (a or b);
    outputs(5493) <= not a;
    outputs(5494) <= b;
    outputs(5495) <= a and not b;
    outputs(5496) <= not (a xor b);
    outputs(5497) <= not a or b;
    outputs(5498) <= b;
    outputs(5499) <= a and b;
    outputs(5500) <= a and b;
    outputs(5501) <= not (a xor b);
    outputs(5502) <= a xor b;
    outputs(5503) <= not a;
    outputs(5504) <= a and b;
    outputs(5505) <= not (a xor b);
    outputs(5506) <= a xor b;
    outputs(5507) <= not b;
    outputs(5508) <= a or b;
    outputs(5509) <= not b;
    outputs(5510) <= a and b;
    outputs(5511) <= not a;
    outputs(5512) <= not b or a;
    outputs(5513) <= b;
    outputs(5514) <= not a or b;
    outputs(5515) <= b;
    outputs(5516) <= b and not a;
    outputs(5517) <= not (a and b);
    outputs(5518) <= b and not a;
    outputs(5519) <= not a or b;
    outputs(5520) <= a xor b;
    outputs(5521) <= a;
    outputs(5522) <= a xor b;
    outputs(5523) <= not b;
    outputs(5524) <= a xor b;
    outputs(5525) <= not (a xor b);
    outputs(5526) <= b;
    outputs(5527) <= not (a xor b);
    outputs(5528) <= a xor b;
    outputs(5529) <= not (a or b);
    outputs(5530) <= a xor b;
    outputs(5531) <= b;
    outputs(5532) <= a xor b;
    outputs(5533) <= not a;
    outputs(5534) <= not a;
    outputs(5535) <= not a;
    outputs(5536) <= b;
    outputs(5537) <= b;
    outputs(5538) <= not (a or b);
    outputs(5539) <= a xor b;
    outputs(5540) <= not (a xor b);
    outputs(5541) <= a and not b;
    outputs(5542) <= not (a xor b);
    outputs(5543) <= not a;
    outputs(5544) <= b and not a;
    outputs(5545) <= not (a xor b);
    outputs(5546) <= b;
    outputs(5547) <= not a;
    outputs(5548) <= not (a or b);
    outputs(5549) <= a xor b;
    outputs(5550) <= a xor b;
    outputs(5551) <= a;
    outputs(5552) <= a xor b;
    outputs(5553) <= not (a or b);
    outputs(5554) <= not b;
    outputs(5555) <= not b;
    outputs(5556) <= a xor b;
    outputs(5557) <= a;
    outputs(5558) <= not b;
    outputs(5559) <= not (a xor b);
    outputs(5560) <= a and not b;
    outputs(5561) <= not (a xor b);
    outputs(5562) <= not a;
    outputs(5563) <= not (a xor b);
    outputs(5564) <= not a;
    outputs(5565) <= a xor b;
    outputs(5566) <= a xor b;
    outputs(5567) <= not (a or b);
    outputs(5568) <= a xor b;
    outputs(5569) <= a;
    outputs(5570) <= not b;
    outputs(5571) <= a xor b;
    outputs(5572) <= not a or b;
    outputs(5573) <= a;
    outputs(5574) <= not (a or b);
    outputs(5575) <= not b;
    outputs(5576) <= a xor b;
    outputs(5577) <= not (a or b);
    outputs(5578) <= a xor b;
    outputs(5579) <= not b;
    outputs(5580) <= b and not a;
    outputs(5581) <= b and not a;
    outputs(5582) <= a and b;
    outputs(5583) <= not a;
    outputs(5584) <= not (a xor b);
    outputs(5585) <= a xor b;
    outputs(5586) <= not a;
    outputs(5587) <= not b;
    outputs(5588) <= a;
    outputs(5589) <= not b;
    outputs(5590) <= not (a xor b);
    outputs(5591) <= not b or a;
    outputs(5592) <= not (a xor b);
    outputs(5593) <= not (a xor b);
    outputs(5594) <= a;
    outputs(5595) <= not b or a;
    outputs(5596) <= b and not a;
    outputs(5597) <= b;
    outputs(5598) <= a;
    outputs(5599) <= a;
    outputs(5600) <= a and not b;
    outputs(5601) <= b;
    outputs(5602) <= a and not b;
    outputs(5603) <= not b;
    outputs(5604) <= a;
    outputs(5605) <= not (a xor b);
    outputs(5606) <= b and not a;
    outputs(5607) <= not b;
    outputs(5608) <= a;
    outputs(5609) <= not b;
    outputs(5610) <= b;
    outputs(5611) <= a or b;
    outputs(5612) <= a;
    outputs(5613) <= not b;
    outputs(5614) <= b;
    outputs(5615) <= not (a and b);
    outputs(5616) <= a;
    outputs(5617) <= not (a or b);
    outputs(5618) <= a xor b;
    outputs(5619) <= not a;
    outputs(5620) <= not b;
    outputs(5621) <= a or b;
    outputs(5622) <= b and not a;
    outputs(5623) <= a xor b;
    outputs(5624) <= not (a or b);
    outputs(5625) <= b and not a;
    outputs(5626) <= a and not b;
    outputs(5627) <= not a;
    outputs(5628) <= a and not b;
    outputs(5629) <= b and not a;
    outputs(5630) <= b;
    outputs(5631) <= a and b;
    outputs(5632) <= a and not b;
    outputs(5633) <= a xor b;
    outputs(5634) <= b and not a;
    outputs(5635) <= a;
    outputs(5636) <= b and not a;
    outputs(5637) <= a;
    outputs(5638) <= a xor b;
    outputs(5639) <= not b;
    outputs(5640) <= not b;
    outputs(5641) <= b;
    outputs(5642) <= a and not b;
    outputs(5643) <= a and b;
    outputs(5644) <= b and not a;
    outputs(5645) <= not (a xor b);
    outputs(5646) <= a and b;
    outputs(5647) <= not b;
    outputs(5648) <= a;
    outputs(5649) <= not b or a;
    outputs(5650) <= a xor b;
    outputs(5651) <= not (a xor b);
    outputs(5652) <= not (a and b);
    outputs(5653) <= b;
    outputs(5654) <= not a;
    outputs(5655) <= b and not a;
    outputs(5656) <= a and not b;
    outputs(5657) <= not a;
    outputs(5658) <= b;
    outputs(5659) <= a xor b;
    outputs(5660) <= not b;
    outputs(5661) <= b;
    outputs(5662) <= b;
    outputs(5663) <= not b or a;
    outputs(5664) <= not a;
    outputs(5665) <= b and not a;
    outputs(5666) <= a xor b;
    outputs(5667) <= b and not a;
    outputs(5668) <= a and not b;
    outputs(5669) <= not (a xor b);
    outputs(5670) <= not b;
    outputs(5671) <= b and not a;
    outputs(5672) <= not (a or b);
    outputs(5673) <= a and b;
    outputs(5674) <= a or b;
    outputs(5675) <= not (a or b);
    outputs(5676) <= not (a xor b);
    outputs(5677) <= a and b;
    outputs(5678) <= not (a or b);
    outputs(5679) <= not (a xor b);
    outputs(5680) <= b and not a;
    outputs(5681) <= a;
    outputs(5682) <= not (a or b);
    outputs(5683) <= a and not b;
    outputs(5684) <= a or b;
    outputs(5685) <= not (a or b);
    outputs(5686) <= not b;
    outputs(5687) <= a and not b;
    outputs(5688) <= not b;
    outputs(5689) <= a;
    outputs(5690) <= not (a or b);
    outputs(5691) <= a xor b;
    outputs(5692) <= a;
    outputs(5693) <= a xor b;
    outputs(5694) <= a;
    outputs(5695) <= not b;
    outputs(5696) <= not a;
    outputs(5697) <= a xor b;
    outputs(5698) <= b and not a;
    outputs(5699) <= a xor b;
    outputs(5700) <= not b;
    outputs(5701) <= not b;
    outputs(5702) <= not b;
    outputs(5703) <= not (a xor b);
    outputs(5704) <= a;
    outputs(5705) <= not (a or b);
    outputs(5706) <= a xor b;
    outputs(5707) <= not (a or b);
    outputs(5708) <= not (a xor b);
    outputs(5709) <= b and not a;
    outputs(5710) <= b and not a;
    outputs(5711) <= a and b;
    outputs(5712) <= b and not a;
    outputs(5713) <= not b;
    outputs(5714) <= not (a xor b);
    outputs(5715) <= not (a or b);
    outputs(5716) <= not (a or b);
    outputs(5717) <= b;
    outputs(5718) <= a;
    outputs(5719) <= not b or a;
    outputs(5720) <= a and not b;
    outputs(5721) <= not (a xor b);
    outputs(5722) <= not b;
    outputs(5723) <= a and b;
    outputs(5724) <= a;
    outputs(5725) <= a xor b;
    outputs(5726) <= not b or a;
    outputs(5727) <= b and not a;
    outputs(5728) <= not a;
    outputs(5729) <= not a;
    outputs(5730) <= a xor b;
    outputs(5731) <= not a;
    outputs(5732) <= a;
    outputs(5733) <= not (a or b);
    outputs(5734) <= a xor b;
    outputs(5735) <= b;
    outputs(5736) <= not a;
    outputs(5737) <= a and not b;
    outputs(5738) <= not (a or b);
    outputs(5739) <= not b;
    outputs(5740) <= b;
    outputs(5741) <= not b;
    outputs(5742) <= not b;
    outputs(5743) <= b;
    outputs(5744) <= not a;
    outputs(5745) <= not b;
    outputs(5746) <= b;
    outputs(5747) <= b;
    outputs(5748) <= not (a or b);
    outputs(5749) <= b;
    outputs(5750) <= not b;
    outputs(5751) <= a xor b;
    outputs(5752) <= not (a xor b);
    outputs(5753) <= not (a xor b);
    outputs(5754) <= b and not a;
    outputs(5755) <= a xor b;
    outputs(5756) <= not (a xor b);
    outputs(5757) <= not b or a;
    outputs(5758) <= b and not a;
    outputs(5759) <= not b;
    outputs(5760) <= not (a xor b);
    outputs(5761) <= a;
    outputs(5762) <= b and not a;
    outputs(5763) <= a;
    outputs(5764) <= not (a xor b);
    outputs(5765) <= a and not b;
    outputs(5766) <= not b;
    outputs(5767) <= a and b;
    outputs(5768) <= not a or b;
    outputs(5769) <= not b;
    outputs(5770) <= not b;
    outputs(5771) <= not (a xor b);
    outputs(5772) <= not b;
    outputs(5773) <= b;
    outputs(5774) <= b and not a;
    outputs(5775) <= not (a xor b);
    outputs(5776) <= not a;
    outputs(5777) <= not a or b;
    outputs(5778) <= b and not a;
    outputs(5779) <= a xor b;
    outputs(5780) <= not b;
    outputs(5781) <= a and not b;
    outputs(5782) <= b and not a;
    outputs(5783) <= not (a or b);
    outputs(5784) <= not (a or b);
    outputs(5785) <= not a;
    outputs(5786) <= a xor b;
    outputs(5787) <= a and b;
    outputs(5788) <= not (a xor b);
    outputs(5789) <= not a or b;
    outputs(5790) <= b;
    outputs(5791) <= a xor b;
    outputs(5792) <= b;
    outputs(5793) <= a or b;
    outputs(5794) <= not a;
    outputs(5795) <= not a;
    outputs(5796) <= b;
    outputs(5797) <= a;
    outputs(5798) <= not b;
    outputs(5799) <= a;
    outputs(5800) <= not b;
    outputs(5801) <= not a;
    outputs(5802) <= a xor b;
    outputs(5803) <= a xor b;
    outputs(5804) <= not (a or b);
    outputs(5805) <= a or b;
    outputs(5806) <= not b;
    outputs(5807) <= not (a or b);
    outputs(5808) <= not a;
    outputs(5809) <= a and not b;
    outputs(5810) <= not b;
    outputs(5811) <= not a;
    outputs(5812) <= not a or b;
    outputs(5813) <= not a;
    outputs(5814) <= not (a xor b);
    outputs(5815) <= b and not a;
    outputs(5816) <= a;
    outputs(5817) <= not a;
    outputs(5818) <= not a;
    outputs(5819) <= a and b;
    outputs(5820) <= not (a or b);
    outputs(5821) <= a and b;
    outputs(5822) <= b and not a;
    outputs(5823) <= not a;
    outputs(5824) <= not (a or b);
    outputs(5825) <= a;
    outputs(5826) <= a xor b;
    outputs(5827) <= a xor b;
    outputs(5828) <= not a;
    outputs(5829) <= a or b;
    outputs(5830) <= a xor b;
    outputs(5831) <= a and b;
    outputs(5832) <= a and b;
    outputs(5833) <= not (a or b);
    outputs(5834) <= not b or a;
    outputs(5835) <= a;
    outputs(5836) <= not a;
    outputs(5837) <= b;
    outputs(5838) <= not a or b;
    outputs(5839) <= b;
    outputs(5840) <= b;
    outputs(5841) <= a xor b;
    outputs(5842) <= b and not a;
    outputs(5843) <= a;
    outputs(5844) <= not a;
    outputs(5845) <= a;
    outputs(5846) <= not a or b;
    outputs(5847) <= not b;
    outputs(5848) <= b and not a;
    outputs(5849) <= a and b;
    outputs(5850) <= not b or a;
    outputs(5851) <= not (a or b);
    outputs(5852) <= a;
    outputs(5853) <= not a;
    outputs(5854) <= not a;
    outputs(5855) <= not (a or b);
    outputs(5856) <= not (a xor b);
    outputs(5857) <= not a;
    outputs(5858) <= a xor b;
    outputs(5859) <= a;
    outputs(5860) <= not (a and b);
    outputs(5861) <= not (a xor b);
    outputs(5862) <= b;
    outputs(5863) <= not b or a;
    outputs(5864) <= not a;
    outputs(5865) <= not a;
    outputs(5866) <= not a or b;
    outputs(5867) <= b;
    outputs(5868) <= not b;
    outputs(5869) <= a;
    outputs(5870) <= b;
    outputs(5871) <= b;
    outputs(5872) <= not (a xor b);
    outputs(5873) <= not (a xor b);
    outputs(5874) <= b;
    outputs(5875) <= not (a xor b);
    outputs(5876) <= not (a or b);
    outputs(5877) <= not b;
    outputs(5878) <= not b or a;
    outputs(5879) <= b;
    outputs(5880) <= not b;
    outputs(5881) <= not b or a;
    outputs(5882) <= a or b;
    outputs(5883) <= a and b;
    outputs(5884) <= a;
    outputs(5885) <= b and not a;
    outputs(5886) <= b;
    outputs(5887) <= b;
    outputs(5888) <= a and not b;
    outputs(5889) <= not a;
    outputs(5890) <= b;
    outputs(5891) <= not (a xor b);
    outputs(5892) <= not b;
    outputs(5893) <= not b;
    outputs(5894) <= not a or b;
    outputs(5895) <= a;
    outputs(5896) <= not (a or b);
    outputs(5897) <= not b;
    outputs(5898) <= not a;
    outputs(5899) <= a xor b;
    outputs(5900) <= a and b;
    outputs(5901) <= a xor b;
    outputs(5902) <= not (a or b);
    outputs(5903) <= b;
    outputs(5904) <= not (a and b);
    outputs(5905) <= not b;
    outputs(5906) <= a;
    outputs(5907) <= not a;
    outputs(5908) <= a and b;
    outputs(5909) <= a and not b;
    outputs(5910) <= not (a or b);
    outputs(5911) <= not a or b;
    outputs(5912) <= not a;
    outputs(5913) <= a and not b;
    outputs(5914) <= not b;
    outputs(5915) <= a;
    outputs(5916) <= a and b;
    outputs(5917) <= b and not a;
    outputs(5918) <= a or b;
    outputs(5919) <= not b;
    outputs(5920) <= b and not a;
    outputs(5921) <= a and b;
    outputs(5922) <= not b;
    outputs(5923) <= not (a xor b);
    outputs(5924) <= a;
    outputs(5925) <= b;
    outputs(5926) <= b and not a;
    outputs(5927) <= a or b;
    outputs(5928) <= not a;
    outputs(5929) <= b;
    outputs(5930) <= a and b;
    outputs(5931) <= b and not a;
    outputs(5932) <= not b;
    outputs(5933) <= a or b;
    outputs(5934) <= not (a or b);
    outputs(5935) <= not b;
    outputs(5936) <= not (a and b);
    outputs(5937) <= not b;
    outputs(5938) <= a and not b;
    outputs(5939) <= b and not a;
    outputs(5940) <= not (a or b);
    outputs(5941) <= a and not b;
    outputs(5942) <= a and b;
    outputs(5943) <= not a;
    outputs(5944) <= not (a xor b);
    outputs(5945) <= a;
    outputs(5946) <= not a;
    outputs(5947) <= b and not a;
    outputs(5948) <= b;
    outputs(5949) <= not a;
    outputs(5950) <= not b or a;
    outputs(5951) <= not (a xor b);
    outputs(5952) <= b and not a;
    outputs(5953) <= not (a xor b);
    outputs(5954) <= not b;
    outputs(5955) <= a;
    outputs(5956) <= not b;
    outputs(5957) <= not a;
    outputs(5958) <= not (a xor b);
    outputs(5959) <= a and b;
    outputs(5960) <= not a;
    outputs(5961) <= not (a or b);
    outputs(5962) <= not (a xor b);
    outputs(5963) <= not (a xor b);
    outputs(5964) <= not (a xor b);
    outputs(5965) <= not b;
    outputs(5966) <= not a;
    outputs(5967) <= not (a or b);
    outputs(5968) <= a or b;
    outputs(5969) <= a xor b;
    outputs(5970) <= not (a or b);
    outputs(5971) <= a xor b;
    outputs(5972) <= a or b;
    outputs(5973) <= a xor b;
    outputs(5974) <= b and not a;
    outputs(5975) <= a and not b;
    outputs(5976) <= not a;
    outputs(5977) <= not (a or b);
    outputs(5978) <= not (a xor b);
    outputs(5979) <= not (a or b);
    outputs(5980) <= b;
    outputs(5981) <= b and not a;
    outputs(5982) <= not (a or b);
    outputs(5983) <= not (a xor b);
    outputs(5984) <= not a;
    outputs(5985) <= a and b;
    outputs(5986) <= a and not b;
    outputs(5987) <= b;
    outputs(5988) <= b;
    outputs(5989) <= not b;
    outputs(5990) <= not b;
    outputs(5991) <= a;
    outputs(5992) <= b;
    outputs(5993) <= a xor b;
    outputs(5994) <= b and not a;
    outputs(5995) <= a xor b;
    outputs(5996) <= not (a xor b);
    outputs(5997) <= not (a or b);
    outputs(5998) <= not (a and b);
    outputs(5999) <= a xor b;
    outputs(6000) <= a and not b;
    outputs(6001) <= a or b;
    outputs(6002) <= not (a xor b);
    outputs(6003) <= not b or a;
    outputs(6004) <= not a;
    outputs(6005) <= not a;
    outputs(6006) <= not a;
    outputs(6007) <= b and not a;
    outputs(6008) <= b;
    outputs(6009) <= b;
    outputs(6010) <= a;
    outputs(6011) <= not (a or b);
    outputs(6012) <= not b;
    outputs(6013) <= a or b;
    outputs(6014) <= b;
    outputs(6015) <= a or b;
    outputs(6016) <= not (a and b);
    outputs(6017) <= not (a xor b);
    outputs(6018) <= a and b;
    outputs(6019) <= a xor b;
    outputs(6020) <= a and b;
    outputs(6021) <= not b or a;
    outputs(6022) <= a and b;
    outputs(6023) <= not a;
    outputs(6024) <= a;
    outputs(6025) <= not (a xor b);
    outputs(6026) <= not (a or b);
    outputs(6027) <= b;
    outputs(6028) <= a xor b;
    outputs(6029) <= a;
    outputs(6030) <= a;
    outputs(6031) <= not a;
    outputs(6032) <= not (a xor b);
    outputs(6033) <= a;
    outputs(6034) <= b and not a;
    outputs(6035) <= a xor b;
    outputs(6036) <= a xor b;
    outputs(6037) <= a xor b;
    outputs(6038) <= b;
    outputs(6039) <= not a;
    outputs(6040) <= not b;
    outputs(6041) <= not a or b;
    outputs(6042) <= a xor b;
    outputs(6043) <= not a or b;
    outputs(6044) <= a xor b;
    outputs(6045) <= not b;
    outputs(6046) <= a and not b;
    outputs(6047) <= a;
    outputs(6048) <= not b;
    outputs(6049) <= b;
    outputs(6050) <= not a;
    outputs(6051) <= not (a or b);
    outputs(6052) <= a xor b;
    outputs(6053) <= not a;
    outputs(6054) <= not b;
    outputs(6055) <= not (a xor b);
    outputs(6056) <= a and not b;
    outputs(6057) <= not (a xor b);
    outputs(6058) <= a and not b;
    outputs(6059) <= not (a xor b);
    outputs(6060) <= a and b;
    outputs(6061) <= a;
    outputs(6062) <= b;
    outputs(6063) <= b and not a;
    outputs(6064) <= b;
    outputs(6065) <= not (a xor b);
    outputs(6066) <= a and not b;
    outputs(6067) <= b and not a;
    outputs(6068) <= not (a xor b);
    outputs(6069) <= a;
    outputs(6070) <= a xor b;
    outputs(6071) <= a and b;
    outputs(6072) <= not b;
    outputs(6073) <= not a;
    outputs(6074) <= not (a or b);
    outputs(6075) <= not b;
    outputs(6076) <= not a;
    outputs(6077) <= not a;
    outputs(6078) <= not (a xor b);
    outputs(6079) <= b;
    outputs(6080) <= not a;
    outputs(6081) <= b and not a;
    outputs(6082) <= not a;
    outputs(6083) <= not (a xor b);
    outputs(6084) <= b and not a;
    outputs(6085) <= a xor b;
    outputs(6086) <= a;
    outputs(6087) <= not (a xor b);
    outputs(6088) <= not (a or b);
    outputs(6089) <= b;
    outputs(6090) <= not a;
    outputs(6091) <= not a or b;
    outputs(6092) <= b;
    outputs(6093) <= a;
    outputs(6094) <= not b or a;
    outputs(6095) <= b;
    outputs(6096) <= not (a or b);
    outputs(6097) <= a and not b;
    outputs(6098) <= not (a and b);
    outputs(6099) <= not b;
    outputs(6100) <= a xor b;
    outputs(6101) <= not (a or b);
    outputs(6102) <= a and not b;
    outputs(6103) <= not b;
    outputs(6104) <= not (a or b);
    outputs(6105) <= not a;
    outputs(6106) <= not b;
    outputs(6107) <= not (a xor b);
    outputs(6108) <= a xor b;
    outputs(6109) <= b and not a;
    outputs(6110) <= a and not b;
    outputs(6111) <= not (a xor b);
    outputs(6112) <= b;
    outputs(6113) <= a and not b;
    outputs(6114) <= a;
    outputs(6115) <= not a;
    outputs(6116) <= a and b;
    outputs(6117) <= a and not b;
    outputs(6118) <= a and b;
    outputs(6119) <= a and b;
    outputs(6120) <= a and not b;
    outputs(6121) <= not (a or b);
    outputs(6122) <= not a;
    outputs(6123) <= a xor b;
    outputs(6124) <= a;
    outputs(6125) <= a xor b;
    outputs(6126) <= a;
    outputs(6127) <= a;
    outputs(6128) <= not b;
    outputs(6129) <= not (a or b);
    outputs(6130) <= a;
    outputs(6131) <= a xor b;
    outputs(6132) <= b and not a;
    outputs(6133) <= not b;
    outputs(6134) <= a and b;
    outputs(6135) <= a;
    outputs(6136) <= not b;
    outputs(6137) <= b;
    outputs(6138) <= a and not b;
    outputs(6139) <= b;
    outputs(6140) <= a and not b;
    outputs(6141) <= not (a or b);
    outputs(6142) <= b and not a;
    outputs(6143) <= a and b;
    outputs(6144) <= a xor b;
    outputs(6145) <= not b;
    outputs(6146) <= not (a xor b);
    outputs(6147) <= not b;
    outputs(6148) <= not a;
    outputs(6149) <= not b or a;
    outputs(6150) <= a xor b;
    outputs(6151) <= not a or b;
    outputs(6152) <= not b;
    outputs(6153) <= not (a and b);
    outputs(6154) <= a xor b;
    outputs(6155) <= a and b;
    outputs(6156) <= b and not a;
    outputs(6157) <= b;
    outputs(6158) <= a and not b;
    outputs(6159) <= a xor b;
    outputs(6160) <= not a;
    outputs(6161) <= not (a and b);
    outputs(6162) <= b;
    outputs(6163) <= b;
    outputs(6164) <= a;
    outputs(6165) <= not b or a;
    outputs(6166) <= b;
    outputs(6167) <= not b;
    outputs(6168) <= a;
    outputs(6169) <= b;
    outputs(6170) <= not a;
    outputs(6171) <= a;
    outputs(6172) <= not b;
    outputs(6173) <= not a;
    outputs(6174) <= not b;
    outputs(6175) <= not (a and b);
    outputs(6176) <= a;
    outputs(6177) <= a and b;
    outputs(6178) <= a;
    outputs(6179) <= not (a or b);
    outputs(6180) <= not a;
    outputs(6181) <= a;
    outputs(6182) <= b;
    outputs(6183) <= a or b;
    outputs(6184) <= a xor b;
    outputs(6185) <= a or b;
    outputs(6186) <= a;
    outputs(6187) <= not (a or b);
    outputs(6188) <= not (a xor b);
    outputs(6189) <= b and not a;
    outputs(6190) <= b and not a;
    outputs(6191) <= b;
    outputs(6192) <= not b;
    outputs(6193) <= a xor b;
    outputs(6194) <= not (a and b);
    outputs(6195) <= a and not b;
    outputs(6196) <= not b;
    outputs(6197) <= not a;
    outputs(6198) <= not b;
    outputs(6199) <= a and not b;
    outputs(6200) <= a xor b;
    outputs(6201) <= a and b;
    outputs(6202) <= not a or b;
    outputs(6203) <= not (a or b);
    outputs(6204) <= not a;
    outputs(6205) <= not (a xor b);
    outputs(6206) <= not b;
    outputs(6207) <= a and not b;
    outputs(6208) <= not b;
    outputs(6209) <= a;
    outputs(6210) <= not a;
    outputs(6211) <= not (a and b);
    outputs(6212) <= not b;
    outputs(6213) <= a or b;
    outputs(6214) <= not (a or b);
    outputs(6215) <= not b;
    outputs(6216) <= not (a and b);
    outputs(6217) <= not b;
    outputs(6218) <= a xor b;
    outputs(6219) <= not (a xor b);
    outputs(6220) <= a and not b;
    outputs(6221) <= not a;
    outputs(6222) <= a and b;
    outputs(6223) <= not (a or b);
    outputs(6224) <= a xor b;
    outputs(6225) <= b and not a;
    outputs(6226) <= a xor b;
    outputs(6227) <= a;
    outputs(6228) <= a;
    outputs(6229) <= not a;
    outputs(6230) <= not (a xor b);
    outputs(6231) <= a;
    outputs(6232) <= b;
    outputs(6233) <= b and not a;
    outputs(6234) <= not a;
    outputs(6235) <= a;
    outputs(6236) <= b;
    outputs(6237) <= not a;
    outputs(6238) <= b;
    outputs(6239) <= a xor b;
    outputs(6240) <= not (a and b);
    outputs(6241) <= a;
    outputs(6242) <= not (a xor b);
    outputs(6243) <= b;
    outputs(6244) <= not (a or b);
    outputs(6245) <= b and not a;
    outputs(6246) <= b;
    outputs(6247) <= not b or a;
    outputs(6248) <= not (a xor b);
    outputs(6249) <= not b or a;
    outputs(6250) <= a and not b;
    outputs(6251) <= a and b;
    outputs(6252) <= b;
    outputs(6253) <= a xor b;
    outputs(6254) <= not a;
    outputs(6255) <= a;
    outputs(6256) <= not (a xor b);
    outputs(6257) <= not (a and b);
    outputs(6258) <= not b;
    outputs(6259) <= a;
    outputs(6260) <= a xor b;
    outputs(6261) <= a or b;
    outputs(6262) <= a xor b;
    outputs(6263) <= a xor b;
    outputs(6264) <= not a or b;
    outputs(6265) <= a and b;
    outputs(6266) <= a and b;
    outputs(6267) <= not b or a;
    outputs(6268) <= a and b;
    outputs(6269) <= not a;
    outputs(6270) <= not (a and b);
    outputs(6271) <= a xor b;
    outputs(6272) <= not b;
    outputs(6273) <= a xor b;
    outputs(6274) <= not b or a;
    outputs(6275) <= not (a xor b);
    outputs(6276) <= a and b;
    outputs(6277) <= a xor b;
    outputs(6278) <= a xor b;
    outputs(6279) <= a and b;
    outputs(6280) <= b;
    outputs(6281) <= not b;
    outputs(6282) <= not a;
    outputs(6283) <= b;
    outputs(6284) <= not (a xor b);
    outputs(6285) <= a;
    outputs(6286) <= not a or b;
    outputs(6287) <= a xor b;
    outputs(6288) <= a xor b;
    outputs(6289) <= not (a xor b);
    outputs(6290) <= not b;
    outputs(6291) <= b;
    outputs(6292) <= not a;
    outputs(6293) <= b;
    outputs(6294) <= not (a and b);
    outputs(6295) <= not (a xor b);
    outputs(6296) <= b and not a;
    outputs(6297) <= not b;
    outputs(6298) <= not (a xor b);
    outputs(6299) <= not b or a;
    outputs(6300) <= a xor b;
    outputs(6301) <= a and not b;
    outputs(6302) <= not (a xor b);
    outputs(6303) <= not b;
    outputs(6304) <= not b;
    outputs(6305) <= not b;
    outputs(6306) <= a xor b;
    outputs(6307) <= a;
    outputs(6308) <= not (a and b);
    outputs(6309) <= not (a or b);
    outputs(6310) <= a xor b;
    outputs(6311) <= a or b;
    outputs(6312) <= a;
    outputs(6313) <= not b;
    outputs(6314) <= b;
    outputs(6315) <= not b;
    outputs(6316) <= not (a xor b);
    outputs(6317) <= not b;
    outputs(6318) <= not a;
    outputs(6319) <= b and not a;
    outputs(6320) <= a;
    outputs(6321) <= a or b;
    outputs(6322) <= not (a xor b);
    outputs(6323) <= a and b;
    outputs(6324) <= a xor b;
    outputs(6325) <= not (a and b);
    outputs(6326) <= not (a and b);
    outputs(6327) <= not (a and b);
    outputs(6328) <= not b or a;
    outputs(6329) <= b;
    outputs(6330) <= a xor b;
    outputs(6331) <= not b;
    outputs(6332) <= a xor b;
    outputs(6333) <= a;
    outputs(6334) <= a xor b;
    outputs(6335) <= not (a or b);
    outputs(6336) <= a and not b;
    outputs(6337) <= not (a xor b);
    outputs(6338) <= not (a xor b);
    outputs(6339) <= a or b;
    outputs(6340) <= a xor b;
    outputs(6341) <= a xor b;
    outputs(6342) <= b;
    outputs(6343) <= b;
    outputs(6344) <= b and not a;
    outputs(6345) <= not b or a;
    outputs(6346) <= not (a and b);
    outputs(6347) <= a;
    outputs(6348) <= a xor b;
    outputs(6349) <= not (a or b);
    outputs(6350) <= b;
    outputs(6351) <= a or b;
    outputs(6352) <= not (a xor b);
    outputs(6353) <= a xor b;
    outputs(6354) <= not (a and b);
    outputs(6355) <= not (a xor b);
    outputs(6356) <= a xor b;
    outputs(6357) <= not b or a;
    outputs(6358) <= a xor b;
    outputs(6359) <= not (a xor b);
    outputs(6360) <= a and not b;
    outputs(6361) <= a xor b;
    outputs(6362) <= not a;
    outputs(6363) <= a;
    outputs(6364) <= a xor b;
    outputs(6365) <= not b or a;
    outputs(6366) <= a xor b;
    outputs(6367) <= a or b;
    outputs(6368) <= not b;
    outputs(6369) <= not b;
    outputs(6370) <= not (a xor b);
    outputs(6371) <= a xor b;
    outputs(6372) <= not (a xor b);
    outputs(6373) <= a and not b;
    outputs(6374) <= not (a and b);
    outputs(6375) <= not a or b;
    outputs(6376) <= not (a xor b);
    outputs(6377) <= a or b;
    outputs(6378) <= not b or a;
    outputs(6379) <= not b or a;
    outputs(6380) <= not b;
    outputs(6381) <= not (a xor b);
    outputs(6382) <= not a or b;
    outputs(6383) <= not a;
    outputs(6384) <= a;
    outputs(6385) <= a xor b;
    outputs(6386) <= a;
    outputs(6387) <= a and b;
    outputs(6388) <= b;
    outputs(6389) <= a;
    outputs(6390) <= a;
    outputs(6391) <= not a or b;
    outputs(6392) <= a;
    outputs(6393) <= a and not b;
    outputs(6394) <= not b;
    outputs(6395) <= not b;
    outputs(6396) <= b;
    outputs(6397) <= a or b;
    outputs(6398) <= not b or a;
    outputs(6399) <= not a;
    outputs(6400) <= not a;
    outputs(6401) <= a and not b;
    outputs(6402) <= not a;
    outputs(6403) <= a and b;
    outputs(6404) <= a and not b;
    outputs(6405) <= not (a xor b);
    outputs(6406) <= not (a xor b);
    outputs(6407) <= not b;
    outputs(6408) <= not (a or b);
    outputs(6409) <= a or b;
    outputs(6410) <= a xor b;
    outputs(6411) <= not (a or b);
    outputs(6412) <= a;
    outputs(6413) <= a xor b;
    outputs(6414) <= not (a xor b);
    outputs(6415) <= b and not a;
    outputs(6416) <= not (a xor b);
    outputs(6417) <= not b;
    outputs(6418) <= a xor b;
    outputs(6419) <= not (a xor b);
    outputs(6420) <= b;
    outputs(6421) <= not (a and b);
    outputs(6422) <= not (a xor b);
    outputs(6423) <= a and b;
    outputs(6424) <= not b;
    outputs(6425) <= not (a xor b);
    outputs(6426) <= b and not a;
    outputs(6427) <= b;
    outputs(6428) <= not (a or b);
    outputs(6429) <= not b or a;
    outputs(6430) <= a xor b;
    outputs(6431) <= b;
    outputs(6432) <= not b or a;
    outputs(6433) <= a and b;
    outputs(6434) <= a;
    outputs(6435) <= not (a xor b);
    outputs(6436) <= a;
    outputs(6437) <= b and not a;
    outputs(6438) <= not b;
    outputs(6439) <= b;
    outputs(6440) <= a xor b;
    outputs(6441) <= b and not a;
    outputs(6442) <= not (a xor b);
    outputs(6443) <= a xor b;
    outputs(6444) <= not (a or b);
    outputs(6445) <= a;
    outputs(6446) <= b;
    outputs(6447) <= a;
    outputs(6448) <= not (a xor b);
    outputs(6449) <= not (a or b);
    outputs(6450) <= not a;
    outputs(6451) <= not b or a;
    outputs(6452) <= a xor b;
    outputs(6453) <= a and not b;
    outputs(6454) <= not b or a;
    outputs(6455) <= not (a and b);
    outputs(6456) <= not (a and b);
    outputs(6457) <= not (a xor b);
    outputs(6458) <= not a or b;
    outputs(6459) <= a and b;
    outputs(6460) <= not (a xor b);
    outputs(6461) <= a xor b;
    outputs(6462) <= not b;
    outputs(6463) <= not b or a;
    outputs(6464) <= not (a xor b);
    outputs(6465) <= a;
    outputs(6466) <= a or b;
    outputs(6467) <= a;
    outputs(6468) <= a xor b;
    outputs(6469) <= not (a and b);
    outputs(6470) <= not a;
    outputs(6471) <= not b;
    outputs(6472) <= not (a xor b);
    outputs(6473) <= not (a xor b);
    outputs(6474) <= not b;
    outputs(6475) <= a or b;
    outputs(6476) <= a;
    outputs(6477) <= b;
    outputs(6478) <= a and not b;
    outputs(6479) <= not a or b;
    outputs(6480) <= b;
    outputs(6481) <= b;
    outputs(6482) <= a;
    outputs(6483) <= not a;
    outputs(6484) <= a;
    outputs(6485) <= not (a and b);
    outputs(6486) <= not a or b;
    outputs(6487) <= not (a xor b);
    outputs(6488) <= a;
    outputs(6489) <= a and not b;
    outputs(6490) <= b;
    outputs(6491) <= not a or b;
    outputs(6492) <= not (a or b);
    outputs(6493) <= not a;
    outputs(6494) <= b;
    outputs(6495) <= b;
    outputs(6496) <= not b;
    outputs(6497) <= b;
    outputs(6498) <= a;
    outputs(6499) <= b and not a;
    outputs(6500) <= a and b;
    outputs(6501) <= not (a xor b);
    outputs(6502) <= a and b;
    outputs(6503) <= a;
    outputs(6504) <= a and b;
    outputs(6505) <= not b;
    outputs(6506) <= not (a xor b);
    outputs(6507) <= a and not b;
    outputs(6508) <= not (a xor b);
    outputs(6509) <= b;
    outputs(6510) <= a and not b;
    outputs(6511) <= b;
    outputs(6512) <= b and not a;
    outputs(6513) <= a;
    outputs(6514) <= not b or a;
    outputs(6515) <= a xor b;
    outputs(6516) <= not (a xor b);
    outputs(6517) <= not a or b;
    outputs(6518) <= not b;
    outputs(6519) <= a;
    outputs(6520) <= not a or b;
    outputs(6521) <= not b;
    outputs(6522) <= not a or b;
    outputs(6523) <= a;
    outputs(6524) <= not b;
    outputs(6525) <= a xor b;
    outputs(6526) <= not a;
    outputs(6527) <= a or b;
    outputs(6528) <= not (a xor b);
    outputs(6529) <= b;
    outputs(6530) <= not a;
    outputs(6531) <= not b;
    outputs(6532) <= not (a xor b);
    outputs(6533) <= b and not a;
    outputs(6534) <= not (a xor b);
    outputs(6535) <= not (a and b);
    outputs(6536) <= a xor b;
    outputs(6537) <= not (a xor b);
    outputs(6538) <= b;
    outputs(6539) <= a xor b;
    outputs(6540) <= b;
    outputs(6541) <= not a;
    outputs(6542) <= not b or a;
    outputs(6543) <= not a or b;
    outputs(6544) <= a or b;
    outputs(6545) <= a;
    outputs(6546) <= a or b;
    outputs(6547) <= a or b;
    outputs(6548) <= not a or b;
    outputs(6549) <= a;
    outputs(6550) <= a and b;
    outputs(6551) <= not b;
    outputs(6552) <= not (a xor b);
    outputs(6553) <= b;
    outputs(6554) <= not a or b;
    outputs(6555) <= not a;
    outputs(6556) <= not (a or b);
    outputs(6557) <= not a or b;
    outputs(6558) <= not b;
    outputs(6559) <= not (a xor b);
    outputs(6560) <= not a;
    outputs(6561) <= not a or b;
    outputs(6562) <= b;
    outputs(6563) <= not a;
    outputs(6564) <= a;
    outputs(6565) <= a or b;
    outputs(6566) <= not a;
    outputs(6567) <= not a;
    outputs(6568) <= not a;
    outputs(6569) <= b;
    outputs(6570) <= a xor b;
    outputs(6571) <= not b;
    outputs(6572) <= not a or b;
    outputs(6573) <= not a or b;
    outputs(6574) <= a or b;
    outputs(6575) <= a;
    outputs(6576) <= a xor b;
    outputs(6577) <= not (a or b);
    outputs(6578) <= not (a xor b);
    outputs(6579) <= a and b;
    outputs(6580) <= not a;
    outputs(6581) <= not (a or b);
    outputs(6582) <= not b;
    outputs(6583) <= b;
    outputs(6584) <= a and b;
    outputs(6585) <= not a;
    outputs(6586) <= not (a and b);
    outputs(6587) <= a and b;
    outputs(6588) <= a xor b;
    outputs(6589) <= not b;
    outputs(6590) <= not a;
    outputs(6591) <= not b;
    outputs(6592) <= a xor b;
    outputs(6593) <= not b;
    outputs(6594) <= not (a or b);
    outputs(6595) <= not a;
    outputs(6596) <= not a;
    outputs(6597) <= not b or a;
    outputs(6598) <= not a or b;
    outputs(6599) <= not a;
    outputs(6600) <= not a or b;
    outputs(6601) <= not (a xor b);
    outputs(6602) <= not a;
    outputs(6603) <= a and b;
    outputs(6604) <= not b;
    outputs(6605) <= a xor b;
    outputs(6606) <= not a;
    outputs(6607) <= not (a xor b);
    outputs(6608) <= not (a and b);
    outputs(6609) <= a;
    outputs(6610) <= not a;
    outputs(6611) <= a and b;
    outputs(6612) <= b;
    outputs(6613) <= a and not b;
    outputs(6614) <= not b;
    outputs(6615) <= not b;
    outputs(6616) <= not (a or b);
    outputs(6617) <= not a;
    outputs(6618) <= b;
    outputs(6619) <= not (a or b);
    outputs(6620) <= not (a xor b);
    outputs(6621) <= a or b;
    outputs(6622) <= b and not a;
    outputs(6623) <= not (a xor b);
    outputs(6624) <= not b;
    outputs(6625) <= not (a xor b);
    outputs(6626) <= not a;
    outputs(6627) <= not a or b;
    outputs(6628) <= a xor b;
    outputs(6629) <= a;
    outputs(6630) <= a;
    outputs(6631) <= a;
    outputs(6632) <= not (a or b);
    outputs(6633) <= a xor b;
    outputs(6634) <= not (a xor b);
    outputs(6635) <= a and b;
    outputs(6636) <= not (a xor b);
    outputs(6637) <= not b or a;
    outputs(6638) <= not (a and b);
    outputs(6639) <= b and not a;
    outputs(6640) <= not (a xor b);
    outputs(6641) <= not b or a;
    outputs(6642) <= b;
    outputs(6643) <= b and not a;
    outputs(6644) <= not b or a;
    outputs(6645) <= b;
    outputs(6646) <= not a;
    outputs(6647) <= b;
    outputs(6648) <= a xor b;
    outputs(6649) <= not a or b;
    outputs(6650) <= not (a and b);
    outputs(6651) <= a xor b;
    outputs(6652) <= a xor b;
    outputs(6653) <= b;
    outputs(6654) <= a and not b;
    outputs(6655) <= not a;
    outputs(6656) <= a xor b;
    outputs(6657) <= not (a xor b);
    outputs(6658) <= not b or a;
    outputs(6659) <= b;
    outputs(6660) <= a;
    outputs(6661) <= not b;
    outputs(6662) <= b and not a;
    outputs(6663) <= a or b;
    outputs(6664) <= a xor b;
    outputs(6665) <= not (a or b);
    outputs(6666) <= not (a xor b);
    outputs(6667) <= not (a xor b);
    outputs(6668) <= a and b;
    outputs(6669) <= not (a xor b);
    outputs(6670) <= a and b;
    outputs(6671) <= a or b;
    outputs(6672) <= not (a xor b);
    outputs(6673) <= not a or b;
    outputs(6674) <= b;
    outputs(6675) <= not (a xor b);
    outputs(6676) <= not (a or b);
    outputs(6677) <= not b;
    outputs(6678) <= a and b;
    outputs(6679) <= b and not a;
    outputs(6680) <= a xor b;
    outputs(6681) <= b;
    outputs(6682) <= not b or a;
    outputs(6683) <= a xor b;
    outputs(6684) <= not (a xor b);
    outputs(6685) <= a and not b;
    outputs(6686) <= a;
    outputs(6687) <= not a or b;
    outputs(6688) <= a xor b;
    outputs(6689) <= a and not b;
    outputs(6690) <= not b;
    outputs(6691) <= not (a xor b);
    outputs(6692) <= a;
    outputs(6693) <= a;
    outputs(6694) <= b;
    outputs(6695) <= not (a xor b);
    outputs(6696) <= a and not b;
    outputs(6697) <= not a;
    outputs(6698) <= not (a xor b);
    outputs(6699) <= a xor b;
    outputs(6700) <= not (a and b);
    outputs(6701) <= a xor b;
    outputs(6702) <= a xor b;
    outputs(6703) <= a xor b;
    outputs(6704) <= not b;
    outputs(6705) <= not b or a;
    outputs(6706) <= not (a xor b);
    outputs(6707) <= not a or b;
    outputs(6708) <= not a;
    outputs(6709) <= a and b;
    outputs(6710) <= not (a xor b);
    outputs(6711) <= not b or a;
    outputs(6712) <= a xor b;
    outputs(6713) <= a;
    outputs(6714) <= not b or a;
    outputs(6715) <= a;
    outputs(6716) <= a or b;
    outputs(6717) <= not a or b;
    outputs(6718) <= a and not b;
    outputs(6719) <= b;
    outputs(6720) <= b;
    outputs(6721) <= not (a xor b);
    outputs(6722) <= b and not a;
    outputs(6723) <= not b or a;
    outputs(6724) <= a and b;
    outputs(6725) <= not a;
    outputs(6726) <= not (a xor b);
    outputs(6727) <= b;
    outputs(6728) <= a;
    outputs(6729) <= not (a xor b);
    outputs(6730) <= not b;
    outputs(6731) <= b;
    outputs(6732) <= a;
    outputs(6733) <= not (a and b);
    outputs(6734) <= a and b;
    outputs(6735) <= not a or b;
    outputs(6736) <= not (a xor b);
    outputs(6737) <= a xor b;
    outputs(6738) <= a xor b;
    outputs(6739) <= a xor b;
    outputs(6740) <= a or b;
    outputs(6741) <= not (a xor b);
    outputs(6742) <= b;
    outputs(6743) <= not (a xor b);
    outputs(6744) <= a or b;
    outputs(6745) <= b and not a;
    outputs(6746) <= not b;
    outputs(6747) <= not (a and b);
    outputs(6748) <= not a or b;
    outputs(6749) <= not (a xor b);
    outputs(6750) <= a and not b;
    outputs(6751) <= not (a xor b);
    outputs(6752) <= not a;
    outputs(6753) <= not a;
    outputs(6754) <= a xor b;
    outputs(6755) <= a;
    outputs(6756) <= not a;
    outputs(6757) <= not a or b;
    outputs(6758) <= a and not b;
    outputs(6759) <= not a;
    outputs(6760) <= not (a and b);
    outputs(6761) <= b;
    outputs(6762) <= a xor b;
    outputs(6763) <= not (a and b);
    outputs(6764) <= not (a xor b);
    outputs(6765) <= not (a or b);
    outputs(6766) <= a or b;
    outputs(6767) <= b and not a;
    outputs(6768) <= a or b;
    outputs(6769) <= not b;
    outputs(6770) <= b;
    outputs(6771) <= a;
    outputs(6772) <= not (a xor b);
    outputs(6773) <= a or b;
    outputs(6774) <= not (a and b);
    outputs(6775) <= not b;
    outputs(6776) <= not a or b;
    outputs(6777) <= b;
    outputs(6778) <= a;
    outputs(6779) <= a;
    outputs(6780) <= a xor b;
    outputs(6781) <= not a;
    outputs(6782) <= not a;
    outputs(6783) <= a or b;
    outputs(6784) <= b;
    outputs(6785) <= not a or b;
    outputs(6786) <= not a;
    outputs(6787) <= a or b;
    outputs(6788) <= not b;
    outputs(6789) <= a xor b;
    outputs(6790) <= a;
    outputs(6791) <= b and not a;
    outputs(6792) <= a and not b;
    outputs(6793) <= not b;
    outputs(6794) <= not a or b;
    outputs(6795) <= not (a and b);
    outputs(6796) <= not b;
    outputs(6797) <= a xor b;
    outputs(6798) <= not (a or b);
    outputs(6799) <= a and b;
    outputs(6800) <= not a;
    outputs(6801) <= not (a xor b);
    outputs(6802) <= b and not a;
    outputs(6803) <= a xor b;
    outputs(6804) <= not a or b;
    outputs(6805) <= a xor b;
    outputs(6806) <= not (a xor b);
    outputs(6807) <= not a or b;
    outputs(6808) <= b;
    outputs(6809) <= not a or b;
    outputs(6810) <= not (a xor b);
    outputs(6811) <= not (a xor b);
    outputs(6812) <= not a or b;
    outputs(6813) <= b and not a;
    outputs(6814) <= not a or b;
    outputs(6815) <= a xor b;
    outputs(6816) <= not a;
    outputs(6817) <= not (a xor b);
    outputs(6818) <= b;
    outputs(6819) <= b;
    outputs(6820) <= not b or a;
    outputs(6821) <= a;
    outputs(6822) <= not b;
    outputs(6823) <= a xor b;
    outputs(6824) <= a;
    outputs(6825) <= a;
    outputs(6826) <= a or b;
    outputs(6827) <= not (a xor b);
    outputs(6828) <= not (a xor b);
    outputs(6829) <= b;
    outputs(6830) <= not (a and b);
    outputs(6831) <= b and not a;
    outputs(6832) <= a and b;
    outputs(6833) <= not (a xor b);
    outputs(6834) <= a xor b;
    outputs(6835) <= not b or a;
    outputs(6836) <= a;
    outputs(6837) <= not b;
    outputs(6838) <= b and not a;
    outputs(6839) <= a xor b;
    outputs(6840) <= a xor b;
    outputs(6841) <= a;
    outputs(6842) <= a xor b;
    outputs(6843) <= not a or b;
    outputs(6844) <= a or b;
    outputs(6845) <= not b;
    outputs(6846) <= not a;
    outputs(6847) <= not (a or b);
    outputs(6848) <= b and not a;
    outputs(6849) <= a and b;
    outputs(6850) <= not (a xor b);
    outputs(6851) <= a;
    outputs(6852) <= a and b;
    outputs(6853) <= b and not a;
    outputs(6854) <= a;
    outputs(6855) <= not a;
    outputs(6856) <= a;
    outputs(6857) <= a and not b;
    outputs(6858) <= not (a xor b);
    outputs(6859) <= a xor b;
    outputs(6860) <= not b;
    outputs(6861) <= not b;
    outputs(6862) <= not (a xor b);
    outputs(6863) <= a xor b;
    outputs(6864) <= b;
    outputs(6865) <= not a or b;
    outputs(6866) <= a xor b;
    outputs(6867) <= not a;
    outputs(6868) <= not a;
    outputs(6869) <= b;
    outputs(6870) <= a xor b;
    outputs(6871) <= a and b;
    outputs(6872) <= a;
    outputs(6873) <= a or b;
    outputs(6874) <= a;
    outputs(6875) <= a and not b;
    outputs(6876) <= not a;
    outputs(6877) <= a xor b;
    outputs(6878) <= not a or b;
    outputs(6879) <= a;
    outputs(6880) <= b and not a;
    outputs(6881) <= a and not b;
    outputs(6882) <= b;
    outputs(6883) <= not a;
    outputs(6884) <= b;
    outputs(6885) <= not (a or b);
    outputs(6886) <= not b or a;
    outputs(6887) <= not b;
    outputs(6888) <= not b or a;
    outputs(6889) <= a xor b;
    outputs(6890) <= b and not a;
    outputs(6891) <= not a or b;
    outputs(6892) <= not (a and b);
    outputs(6893) <= not a or b;
    outputs(6894) <= a and not b;
    outputs(6895) <= a and b;
    outputs(6896) <= not b;
    outputs(6897) <= not (a or b);
    outputs(6898) <= a xor b;
    outputs(6899) <= a and b;
    outputs(6900) <= not a;
    outputs(6901) <= a;
    outputs(6902) <= not b or a;
    outputs(6903) <= not b;
    outputs(6904) <= b;
    outputs(6905) <= b and not a;
    outputs(6906) <= not (a and b);
    outputs(6907) <= b;
    outputs(6908) <= a;
    outputs(6909) <= a or b;
    outputs(6910) <= not a;
    outputs(6911) <= b;
    outputs(6912) <= b;
    outputs(6913) <= not a;
    outputs(6914) <= a and b;
    outputs(6915) <= not b;
    outputs(6916) <= not (a xor b);
    outputs(6917) <= a and b;
    outputs(6918) <= b;
    outputs(6919) <= b;
    outputs(6920) <= b;
    outputs(6921) <= a and b;
    outputs(6922) <= not (a xor b);
    outputs(6923) <= a xor b;
    outputs(6924) <= a and not b;
    outputs(6925) <= b and not a;
    outputs(6926) <= not b;
    outputs(6927) <= a and not b;
    outputs(6928) <= not a;
    outputs(6929) <= not b;
    outputs(6930) <= a xor b;
    outputs(6931) <= a xor b;
    outputs(6932) <= not a or b;
    outputs(6933) <= b;
    outputs(6934) <= b;
    outputs(6935) <= b;
    outputs(6936) <= not a;
    outputs(6937) <= not a;
    outputs(6938) <= b and not a;
    outputs(6939) <= not b;
    outputs(6940) <= a and b;
    outputs(6941) <= b and not a;
    outputs(6942) <= not b;
    outputs(6943) <= a and not b;
    outputs(6944) <= not b;
    outputs(6945) <= not (a or b);
    outputs(6946) <= not b;
    outputs(6947) <= b;
    outputs(6948) <= not a;
    outputs(6949) <= b;
    outputs(6950) <= a and not b;
    outputs(6951) <= b and not a;
    outputs(6952) <= not a or b;
    outputs(6953) <= not b or a;
    outputs(6954) <= not a;
    outputs(6955) <= not a or b;
    outputs(6956) <= not b;
    outputs(6957) <= not (a and b);
    outputs(6958) <= a and not b;
    outputs(6959) <= not b or a;
    outputs(6960) <= not a or b;
    outputs(6961) <= not (a xor b);
    outputs(6962) <= a xor b;
    outputs(6963) <= b;
    outputs(6964) <= a;
    outputs(6965) <= b;
    outputs(6966) <= b;
    outputs(6967) <= not a or b;
    outputs(6968) <= a and not b;
    outputs(6969) <= not a;
    outputs(6970) <= b and not a;
    outputs(6971) <= b and not a;
    outputs(6972) <= a xor b;
    outputs(6973) <= not b;
    outputs(6974) <= a and not b;
    outputs(6975) <= not a or b;
    outputs(6976) <= a and b;
    outputs(6977) <= not a or b;
    outputs(6978) <= a and not b;
    outputs(6979) <= a xor b;
    outputs(6980) <= a and not b;
    outputs(6981) <= a and not b;
    outputs(6982) <= a;
    outputs(6983) <= a and b;
    outputs(6984) <= not a;
    outputs(6985) <= a and not b;
    outputs(6986) <= a xor b;
    outputs(6987) <= not a;
    outputs(6988) <= not a;
    outputs(6989) <= not a;
    outputs(6990) <= not (a xor b);
    outputs(6991) <= a xor b;
    outputs(6992) <= a and b;
    outputs(6993) <= a and not b;
    outputs(6994) <= b and not a;
    outputs(6995) <= b;
    outputs(6996) <= not b or a;
    outputs(6997) <= not (a or b);
    outputs(6998) <= a and b;
    outputs(6999) <= not b or a;
    outputs(7000) <= not (a xor b);
    outputs(7001) <= not a or b;
    outputs(7002) <= b and not a;
    outputs(7003) <= a xor b;
    outputs(7004) <= a and not b;
    outputs(7005) <= not a;
    outputs(7006) <= not (a or b);
    outputs(7007) <= not (a xor b);
    outputs(7008) <= not (a or b);
    outputs(7009) <= not b;
    outputs(7010) <= not a or b;
    outputs(7011) <= not (a xor b);
    outputs(7012) <= not (a xor b);
    outputs(7013) <= a and b;
    outputs(7014) <= not (a or b);
    outputs(7015) <= b;
    outputs(7016) <= a xor b;
    outputs(7017) <= not b;
    outputs(7018) <= not b or a;
    outputs(7019) <= not (a xor b);
    outputs(7020) <= not a or b;
    outputs(7021) <= b and not a;
    outputs(7022) <= not b;
    outputs(7023) <= a xor b;
    outputs(7024) <= a and b;
    outputs(7025) <= a xor b;
    outputs(7026) <= not (a and b);
    outputs(7027) <= b;
    outputs(7028) <= a;
    outputs(7029) <= a;
    outputs(7030) <= b;
    outputs(7031) <= a and not b;
    outputs(7032) <= a and b;
    outputs(7033) <= not b;
    outputs(7034) <= a xor b;
    outputs(7035) <= a and b;
    outputs(7036) <= not a or b;
    outputs(7037) <= a and b;
    outputs(7038) <= a and not b;
    outputs(7039) <= not (a or b);
    outputs(7040) <= not a;
    outputs(7041) <= a and b;
    outputs(7042) <= a or b;
    outputs(7043) <= a or b;
    outputs(7044) <= b;
    outputs(7045) <= not a;
    outputs(7046) <= not b;
    outputs(7047) <= not (a and b);
    outputs(7048) <= not a or b;
    outputs(7049) <= not a;
    outputs(7050) <= b and not a;
    outputs(7051) <= a xor b;
    outputs(7052) <= a xor b;
    outputs(7053) <= a and not b;
    outputs(7054) <= not a or b;
    outputs(7055) <= a xor b;
    outputs(7056) <= a and not b;
    outputs(7057) <= not (a or b);
    outputs(7058) <= b;
    outputs(7059) <= not a or b;
    outputs(7060) <= a xor b;
    outputs(7061) <= not (a xor b);
    outputs(7062) <= not (a xor b);
    outputs(7063) <= b and not a;
    outputs(7064) <= a;
    outputs(7065) <= not (a and b);
    outputs(7066) <= a;
    outputs(7067) <= not (a or b);
    outputs(7068) <= not b;
    outputs(7069) <= b;
    outputs(7070) <= not a or b;
    outputs(7071) <= not (a or b);
    outputs(7072) <= not (a and b);
    outputs(7073) <= b;
    outputs(7074) <= a xor b;
    outputs(7075) <= b and not a;
    outputs(7076) <= b and not a;
    outputs(7077) <= b and not a;
    outputs(7078) <= not (a xor b);
    outputs(7079) <= a xor b;
    outputs(7080) <= a xor b;
    outputs(7081) <= not (a xor b);
    outputs(7082) <= a and not b;
    outputs(7083) <= not (a or b);
    outputs(7084) <= a;
    outputs(7085) <= a xor b;
    outputs(7086) <= not b;
    outputs(7087) <= not (a and b);
    outputs(7088) <= not (a xor b);
    outputs(7089) <= not a;
    outputs(7090) <= not a or b;
    outputs(7091) <= not (a or b);
    outputs(7092) <= not (a xor b);
    outputs(7093) <= not a or b;
    outputs(7094) <= b and not a;
    outputs(7095) <= not b;
    outputs(7096) <= not (a xor b);
    outputs(7097) <= not a;
    outputs(7098) <= a or b;
    outputs(7099) <= a;
    outputs(7100) <= not (a or b);
    outputs(7101) <= a xor b;
    outputs(7102) <= not (a xor b);
    outputs(7103) <= a;
    outputs(7104) <= a;
    outputs(7105) <= not b;
    outputs(7106) <= a and not b;
    outputs(7107) <= a xor b;
    outputs(7108) <= a and not b;
    outputs(7109) <= not a;
    outputs(7110) <= not b or a;
    outputs(7111) <= b and not a;
    outputs(7112) <= not (a xor b);
    outputs(7113) <= a and b;
    outputs(7114) <= not a;
    outputs(7115) <= b;
    outputs(7116) <= a or b;
    outputs(7117) <= not (a xor b);
    outputs(7118) <= a xor b;
    outputs(7119) <= b and not a;
    outputs(7120) <= b;
    outputs(7121) <= a;
    outputs(7122) <= a and not b;
    outputs(7123) <= not b or a;
    outputs(7124) <= a and not b;
    outputs(7125) <= not (a or b);
    outputs(7126) <= not (a or b);
    outputs(7127) <= a and b;
    outputs(7128) <= a and b;
    outputs(7129) <= not a;
    outputs(7130) <= a and b;
    outputs(7131) <= not (a or b);
    outputs(7132) <= not b or a;
    outputs(7133) <= b;
    outputs(7134) <= a;
    outputs(7135) <= a;
    outputs(7136) <= not (a xor b);
    outputs(7137) <= not a;
    outputs(7138) <= not b;
    outputs(7139) <= a and b;
    outputs(7140) <= a and not b;
    outputs(7141) <= a;
    outputs(7142) <= a xor b;
    outputs(7143) <= not b;
    outputs(7144) <= a and not b;
    outputs(7145) <= a and not b;
    outputs(7146) <= not a or b;
    outputs(7147) <= a xor b;
    outputs(7148) <= b;
    outputs(7149) <= not (a or b);
    outputs(7150) <= a xor b;
    outputs(7151) <= not b;
    outputs(7152) <= a and not b;
    outputs(7153) <= b and not a;
    outputs(7154) <= not (a or b);
    outputs(7155) <= b;
    outputs(7156) <= a and b;
    outputs(7157) <= not (a xor b);
    outputs(7158) <= not (a xor b);
    outputs(7159) <= not b or a;
    outputs(7160) <= not b or a;
    outputs(7161) <= a and b;
    outputs(7162) <= a xor b;
    outputs(7163) <= a;
    outputs(7164) <= a or b;
    outputs(7165) <= not a;
    outputs(7166) <= a;
    outputs(7167) <= a xor b;
    outputs(7168) <= a and b;
    outputs(7169) <= a xor b;
    outputs(7170) <= b and not a;
    outputs(7171) <= not a;
    outputs(7172) <= not a;
    outputs(7173) <= not b;
    outputs(7174) <= b and not a;
    outputs(7175) <= a xor b;
    outputs(7176) <= a xor b;
    outputs(7177) <= a and not b;
    outputs(7178) <= not a;
    outputs(7179) <= a and not b;
    outputs(7180) <= a and b;
    outputs(7181) <= not (a or b);
    outputs(7182) <= a or b;
    outputs(7183) <= a xor b;
    outputs(7184) <= not b;
    outputs(7185) <= b;
    outputs(7186) <= a and not b;
    outputs(7187) <= b and not a;
    outputs(7188) <= a xor b;
    outputs(7189) <= not (a or b);
    outputs(7190) <= not b or a;
    outputs(7191) <= not a;
    outputs(7192) <= not (a xor b);
    outputs(7193) <= a and not b;
    outputs(7194) <= a and not b;
    outputs(7195) <= a or b;
    outputs(7196) <= not (a or b);
    outputs(7197) <= not (a xor b);
    outputs(7198) <= b and not a;
    outputs(7199) <= a and not b;
    outputs(7200) <= a and not b;
    outputs(7201) <= a;
    outputs(7202) <= not b;
    outputs(7203) <= a;
    outputs(7204) <= a and not b;
    outputs(7205) <= b and not a;
    outputs(7206) <= b;
    outputs(7207) <= not a;
    outputs(7208) <= b;
    outputs(7209) <= a xor b;
    outputs(7210) <= a xor b;
    outputs(7211) <= not b;
    outputs(7212) <= a and b;
    outputs(7213) <= a or b;
    outputs(7214) <= not b;
    outputs(7215) <= not (a xor b);
    outputs(7216) <= a and not b;
    outputs(7217) <= not b or a;
    outputs(7218) <= a xor b;
    outputs(7219) <= a xor b;
    outputs(7220) <= not a;
    outputs(7221) <= b;
    outputs(7222) <= b and not a;
    outputs(7223) <= a;
    outputs(7224) <= b;
    outputs(7225) <= a;
    outputs(7226) <= not b;
    outputs(7227) <= not b;
    outputs(7228) <= a;
    outputs(7229) <= not a;
    outputs(7230) <= not a;
    outputs(7231) <= a xor b;
    outputs(7232) <= not a;
    outputs(7233) <= a;
    outputs(7234) <= a xor b;
    outputs(7235) <= a xor b;
    outputs(7236) <= a xor b;
    outputs(7237) <= not a;
    outputs(7238) <= not a;
    outputs(7239) <= not a;
    outputs(7240) <= b and not a;
    outputs(7241) <= a xor b;
    outputs(7242) <= not (a xor b);
    outputs(7243) <= not a;
    outputs(7244) <= not (a xor b);
    outputs(7245) <= not b;
    outputs(7246) <= b;
    outputs(7247) <= a;
    outputs(7248) <= b and not a;
    outputs(7249) <= a;
    outputs(7250) <= b and not a;
    outputs(7251) <= not (a or b);
    outputs(7252) <= b;
    outputs(7253) <= a;
    outputs(7254) <= not b or a;
    outputs(7255) <= a and not b;
    outputs(7256) <= not (a or b);
    outputs(7257) <= not b;
    outputs(7258) <= not a or b;
    outputs(7259) <= b;
    outputs(7260) <= a and b;
    outputs(7261) <= a;
    outputs(7262) <= not (a xor b);
    outputs(7263) <= b;
    outputs(7264) <= not (a and b);
    outputs(7265) <= b;
    outputs(7266) <= not b;
    outputs(7267) <= not (a or b);
    outputs(7268) <= a and not b;
    outputs(7269) <= b and not a;
    outputs(7270) <= not a;
    outputs(7271) <= not (a xor b);
    outputs(7272) <= a or b;
    outputs(7273) <= not b;
    outputs(7274) <= not a;
    outputs(7275) <= a;
    outputs(7276) <= a and b;
    outputs(7277) <= b and not a;
    outputs(7278) <= b and not a;
    outputs(7279) <= not (a and b);
    outputs(7280) <= not (a or b);
    outputs(7281) <= a;
    outputs(7282) <= not a;
    outputs(7283) <= a;
    outputs(7284) <= b and not a;
    outputs(7285) <= not a or b;
    outputs(7286) <= b and not a;
    outputs(7287) <= a and b;
    outputs(7288) <= a;
    outputs(7289) <= not b or a;
    outputs(7290) <= a;
    outputs(7291) <= not (a or b);
    outputs(7292) <= not a;
    outputs(7293) <= a and b;
    outputs(7294) <= not (a and b);
    outputs(7295) <= a and not b;
    outputs(7296) <= not b;
    outputs(7297) <= not b;
    outputs(7298) <= not a;
    outputs(7299) <= not (a xor b);
    outputs(7300) <= not a;
    outputs(7301) <= not (a xor b);
    outputs(7302) <= not b;
    outputs(7303) <= a or b;
    outputs(7304) <= not (a or b);
    outputs(7305) <= a xor b;
    outputs(7306) <= a xor b;
    outputs(7307) <= b;
    outputs(7308) <= not a;
    outputs(7309) <= not a;
    outputs(7310) <= a and not b;
    outputs(7311) <= b;
    outputs(7312) <= not b;
    outputs(7313) <= a and b;
    outputs(7314) <= a and b;
    outputs(7315) <= a xor b;
    outputs(7316) <= b and not a;
    outputs(7317) <= a xor b;
    outputs(7318) <= not b;
    outputs(7319) <= b;
    outputs(7320) <= a and b;
    outputs(7321) <= a and not b;
    outputs(7322) <= b;
    outputs(7323) <= a xor b;
    outputs(7324) <= a xor b;
    outputs(7325) <= a xor b;
    outputs(7326) <= not (a xor b);
    outputs(7327) <= not (a or b);
    outputs(7328) <= not b;
    outputs(7329) <= a and b;
    outputs(7330) <= b and not a;
    outputs(7331) <= not a;
    outputs(7332) <= not b;
    outputs(7333) <= a and not b;
    outputs(7334) <= a;
    outputs(7335) <= not (a or b);
    outputs(7336) <= a xor b;
    outputs(7337) <= not a;
    outputs(7338) <= b;
    outputs(7339) <= a and not b;
    outputs(7340) <= b and not a;
    outputs(7341) <= not b;
    outputs(7342) <= not a;
    outputs(7343) <= b;
    outputs(7344) <= a xor b;
    outputs(7345) <= a xor b;
    outputs(7346) <= not (a xor b);
    outputs(7347) <= not (a xor b);
    outputs(7348) <= not b;
    outputs(7349) <= not a;
    outputs(7350) <= b and not a;
    outputs(7351) <= a;
    outputs(7352) <= not b;
    outputs(7353) <= not b;
    outputs(7354) <= not a;
    outputs(7355) <= not a;
    outputs(7356) <= a;
    outputs(7357) <= a;
    outputs(7358) <= not (a or b);
    outputs(7359) <= not (a or b);
    outputs(7360) <= not (a xor b);
    outputs(7361) <= not (a xor b);
    outputs(7362) <= a or b;
    outputs(7363) <= not (a xor b);
    outputs(7364) <= b;
    outputs(7365) <= not b;
    outputs(7366) <= not a;
    outputs(7367) <= b;
    outputs(7368) <= a xor b;
    outputs(7369) <= a xor b;
    outputs(7370) <= not (a and b);
    outputs(7371) <= not (a xor b);
    outputs(7372) <= not b;
    outputs(7373) <= b and not a;
    outputs(7374) <= not b;
    outputs(7375) <= a xor b;
    outputs(7376) <= not b;
    outputs(7377) <= not (a xor b);
    outputs(7378) <= a;
    outputs(7379) <= not a;
    outputs(7380) <= not (a or b);
    outputs(7381) <= not (a xor b);
    outputs(7382) <= not (a xor b);
    outputs(7383) <= not a;
    outputs(7384) <= b;
    outputs(7385) <= b;
    outputs(7386) <= a and b;
    outputs(7387) <= not b;
    outputs(7388) <= a;
    outputs(7389) <= a and not b;
    outputs(7390) <= a;
    outputs(7391) <= not (a xor b);
    outputs(7392) <= not (a xor b);
    outputs(7393) <= a xor b;
    outputs(7394) <= b;
    outputs(7395) <= a and b;
    outputs(7396) <= b;
    outputs(7397) <= a xor b;
    outputs(7398) <= not a;
    outputs(7399) <= a and not b;
    outputs(7400) <= not (a xor b);
    outputs(7401) <= not b;
    outputs(7402) <= not (a or b);
    outputs(7403) <= not (a xor b);
    outputs(7404) <= a and not b;
    outputs(7405) <= not (a xor b);
    outputs(7406) <= not (a or b);
    outputs(7407) <= not a or b;
    outputs(7408) <= a and b;
    outputs(7409) <= not a or b;
    outputs(7410) <= not b;
    outputs(7411) <= not b;
    outputs(7412) <= a and not b;
    outputs(7413) <= not (a xor b);
    outputs(7414) <= a xor b;
    outputs(7415) <= a and not b;
    outputs(7416) <= b;
    outputs(7417) <= a xor b;
    outputs(7418) <= b and not a;
    outputs(7419) <= a and not b;
    outputs(7420) <= not (a or b);
    outputs(7421) <= b;
    outputs(7422) <= not a;
    outputs(7423) <= a and b;
    outputs(7424) <= b and not a;
    outputs(7425) <= not a;
    outputs(7426) <= a and b;
    outputs(7427) <= not b;
    outputs(7428) <= b;
    outputs(7429) <= not (a xor b);
    outputs(7430) <= not (a or b);
    outputs(7431) <= not (a xor b);
    outputs(7432) <= a or b;
    outputs(7433) <= not (a or b);
    outputs(7434) <= not (a or b);
    outputs(7435) <= b;
    outputs(7436) <= a and not b;
    outputs(7437) <= b;
    outputs(7438) <= a;
    outputs(7439) <= not (a xor b);
    outputs(7440) <= a;
    outputs(7441) <= a xor b;
    outputs(7442) <= not a;
    outputs(7443) <= a and not b;
    outputs(7444) <= not (a and b);
    outputs(7445) <= not b;
    outputs(7446) <= not a;
    outputs(7447) <= not (a xor b);
    outputs(7448) <= not (a and b);
    outputs(7449) <= a xor b;
    outputs(7450) <= not (a and b);
    outputs(7451) <= not a;
    outputs(7452) <= not (a or b);
    outputs(7453) <= b;
    outputs(7454) <= not (a or b);
    outputs(7455) <= not (a or b);
    outputs(7456) <= not (a xor b);
    outputs(7457) <= not b;
    outputs(7458) <= a and not b;
    outputs(7459) <= not (a xor b);
    outputs(7460) <= a xor b;
    outputs(7461) <= a xor b;
    outputs(7462) <= not (a or b);
    outputs(7463) <= a xor b;
    outputs(7464) <= a;
    outputs(7465) <= not (a xor b);
    outputs(7466) <= b and not a;
    outputs(7467) <= not a or b;
    outputs(7468) <= a xor b;
    outputs(7469) <= not a;
    outputs(7470) <= not (a xor b);
    outputs(7471) <= not b;
    outputs(7472) <= a and b;
    outputs(7473) <= b;
    outputs(7474) <= not a;
    outputs(7475) <= a;
    outputs(7476) <= not b;
    outputs(7477) <= not b;
    outputs(7478) <= b;
    outputs(7479) <= not b;
    outputs(7480) <= a and b;
    outputs(7481) <= not a;
    outputs(7482) <= not (a xor b);
    outputs(7483) <= a and b;
    outputs(7484) <= b and not a;
    outputs(7485) <= a;
    outputs(7486) <= a or b;
    outputs(7487) <= a xor b;
    outputs(7488) <= a and not b;
    outputs(7489) <= b and not a;
    outputs(7490) <= not a;
    outputs(7491) <= a;
    outputs(7492) <= a xor b;
    outputs(7493) <= a;
    outputs(7494) <= b;
    outputs(7495) <= a xor b;
    outputs(7496) <= not (a or b);
    outputs(7497) <= a and b;
    outputs(7498) <= not (a or b);
    outputs(7499) <= not (a xor b);
    outputs(7500) <= b;
    outputs(7501) <= a xor b;
    outputs(7502) <= a;
    outputs(7503) <= a;
    outputs(7504) <= a xor b;
    outputs(7505) <= a xor b;
    outputs(7506) <= a;
    outputs(7507) <= a;
    outputs(7508) <= b and not a;
    outputs(7509) <= not (a or b);
    outputs(7510) <= not (a or b);
    outputs(7511) <= b;
    outputs(7512) <= not b;
    outputs(7513) <= not (a or b);
    outputs(7514) <= a;
    outputs(7515) <= a and not b;
    outputs(7516) <= not (a and b);
    outputs(7517) <= not a or b;
    outputs(7518) <= a and not b;
    outputs(7519) <= not (a xor b);
    outputs(7520) <= not b;
    outputs(7521) <= b;
    outputs(7522) <= b and not a;
    outputs(7523) <= a xor b;
    outputs(7524) <= a;
    outputs(7525) <= not (a xor b);
    outputs(7526) <= a and b;
    outputs(7527) <= not (a or b);
    outputs(7528) <= a;
    outputs(7529) <= not (a xor b);
    outputs(7530) <= not (a and b);
    outputs(7531) <= a xor b;
    outputs(7532) <= not b;
    outputs(7533) <= a and not b;
    outputs(7534) <= b;
    outputs(7535) <= a or b;
    outputs(7536) <= a;
    outputs(7537) <= a;
    outputs(7538) <= not (a xor b);
    outputs(7539) <= a or b;
    outputs(7540) <= a or b;
    outputs(7541) <= b;
    outputs(7542) <= not b;
    outputs(7543) <= not (a xor b);
    outputs(7544) <= a xor b;
    outputs(7545) <= not b;
    outputs(7546) <= a;
    outputs(7547) <= not (a xor b);
    outputs(7548) <= a xor b;
    outputs(7549) <= not a or b;
    outputs(7550) <= b;
    outputs(7551) <= a;
    outputs(7552) <= not b;
    outputs(7553) <= a xor b;
    outputs(7554) <= b;
    outputs(7555) <= b;
    outputs(7556) <= not (a or b);
    outputs(7557) <= a xor b;
    outputs(7558) <= a xor b;
    outputs(7559) <= a xor b;
    outputs(7560) <= b and not a;
    outputs(7561) <= a;
    outputs(7562) <= not (a xor b);
    outputs(7563) <= a;
    outputs(7564) <= a xor b;
    outputs(7565) <= not b or a;
    outputs(7566) <= a xor b;
    outputs(7567) <= not (a xor b);
    outputs(7568) <= not a;
    outputs(7569) <= not b;
    outputs(7570) <= not b;
    outputs(7571) <= b and not a;
    outputs(7572) <= not (a xor b);
    outputs(7573) <= a xor b;
    outputs(7574) <= not a;
    outputs(7575) <= not (a or b);
    outputs(7576) <= a xor b;
    outputs(7577) <= a and not b;
    outputs(7578) <= a;
    outputs(7579) <= a;
    outputs(7580) <= a xor b;
    outputs(7581) <= a and b;
    outputs(7582) <= not (a xor b);
    outputs(7583) <= not (a xor b);
    outputs(7584) <= b and not a;
    outputs(7585) <= not (a or b);
    outputs(7586) <= not (a or b);
    outputs(7587) <= not (a xor b);
    outputs(7588) <= a xor b;
    outputs(7589) <= not (a xor b);
    outputs(7590) <= not b;
    outputs(7591) <= not (a xor b);
    outputs(7592) <= a xor b;
    outputs(7593) <= not b;
    outputs(7594) <= a;
    outputs(7595) <= not a;
    outputs(7596) <= not (a xor b);
    outputs(7597) <= not b;
    outputs(7598) <= a;
    outputs(7599) <= not (a xor b);
    outputs(7600) <= not (a xor b);
    outputs(7601) <= b;
    outputs(7602) <= not (a xor b);
    outputs(7603) <= a xor b;
    outputs(7604) <= b and not a;
    outputs(7605) <= not (a or b);
    outputs(7606) <= a;
    outputs(7607) <= not a;
    outputs(7608) <= not a or b;
    outputs(7609) <= a;
    outputs(7610) <= not a;
    outputs(7611) <= b;
    outputs(7612) <= b and not a;
    outputs(7613) <= a xor b;
    outputs(7614) <= a and not b;
    outputs(7615) <= a xor b;
    outputs(7616) <= not a or b;
    outputs(7617) <= a and b;
    outputs(7618) <= not (a xor b);
    outputs(7619) <= a and b;
    outputs(7620) <= not a;
    outputs(7621) <= a or b;
    outputs(7622) <= a;
    outputs(7623) <= a;
    outputs(7624) <= a and b;
    outputs(7625) <= a xor b;
    outputs(7626) <= b;
    outputs(7627) <= a;
    outputs(7628) <= b;
    outputs(7629) <= not (a xor b);
    outputs(7630) <= not b or a;
    outputs(7631) <= a xor b;
    outputs(7632) <= not a;
    outputs(7633) <= not a;
    outputs(7634) <= not b;
    outputs(7635) <= a;
    outputs(7636) <= not (a xor b);
    outputs(7637) <= not (a xor b);
    outputs(7638) <= a and not b;
    outputs(7639) <= b;
    outputs(7640) <= not (a or b);
    outputs(7641) <= a xor b;
    outputs(7642) <= b and not a;
    outputs(7643) <= a or b;
    outputs(7644) <= a and b;
    outputs(7645) <= b and not a;
    outputs(7646) <= a and b;
    outputs(7647) <= not (a xor b);
    outputs(7648) <= not (a xor b);
    outputs(7649) <= a;
    outputs(7650) <= b and not a;
    outputs(7651) <= not a;
    outputs(7652) <= a xor b;
    outputs(7653) <= a;
    outputs(7654) <= not a;
    outputs(7655) <= a and not b;
    outputs(7656) <= a xor b;
    outputs(7657) <= a and b;
    outputs(7658) <= not (a xor b);
    outputs(7659) <= not (a and b);
    outputs(7660) <= a;
    outputs(7661) <= a and b;
    outputs(7662) <= b and not a;
    outputs(7663) <= b;
    outputs(7664) <= not b or a;
    outputs(7665) <= not (a xor b);
    outputs(7666) <= not a;
    outputs(7667) <= b and not a;
    outputs(7668) <= not b;
    outputs(7669) <= a and not b;
    outputs(7670) <= b;
    outputs(7671) <= not a;
    outputs(7672) <= b;
    outputs(7673) <= not a;
    outputs(7674) <= not b;
    outputs(7675) <= a and not b;
    outputs(7676) <= b;
    outputs(7677) <= a and b;
    outputs(7678) <= not b;
    outputs(7679) <= a or b;
end Behavioral;
