library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(12799 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(12799 downto 0);
    signal layer1_outputs : std_logic_vector(12799 downto 0);
    signal layer2_outputs : std_logic_vector(12799 downto 0);

begin

    layer0_outputs(0) <= not(inputs(220));
    layer0_outputs(1) <= not(inputs(64));
    layer0_outputs(2) <= '1';
    layer0_outputs(3) <= not(inputs(117));
    layer0_outputs(4) <= not(inputs(25));
    layer0_outputs(5) <= inputs(55);
    layer0_outputs(6) <= not(inputs(167));
    layer0_outputs(7) <= not((inputs(117)) and (inputs(121)));
    layer0_outputs(8) <= (inputs(0)) xor (inputs(107));
    layer0_outputs(9) <= not(inputs(53));
    layer0_outputs(10) <= not(inputs(61));
    layer0_outputs(11) <= (inputs(43)) or (inputs(109));
    layer0_outputs(12) <= (inputs(210)) xor (inputs(202));
    layer0_outputs(13) <= (inputs(127)) or (inputs(11));
    layer0_outputs(14) <= not(inputs(244)) or (inputs(239));
    layer0_outputs(15) <= not(inputs(65)) or (inputs(145));
    layer0_outputs(16) <= (inputs(112)) or (inputs(248));
    layer0_outputs(17) <= not(inputs(245));
    layer0_outputs(18) <= not(inputs(159));
    layer0_outputs(19) <= (inputs(145)) or (inputs(7));
    layer0_outputs(20) <= not(inputs(11)) or (inputs(97));
    layer0_outputs(21) <= inputs(231);
    layer0_outputs(22) <= (inputs(47)) or (inputs(77));
    layer0_outputs(23) <= inputs(89);
    layer0_outputs(24) <= (inputs(14)) and (inputs(14));
    layer0_outputs(25) <= not(inputs(173)) or (inputs(48));
    layer0_outputs(26) <= (inputs(44)) xor (inputs(210));
    layer0_outputs(27) <= not((inputs(143)) xor (inputs(101)));
    layer0_outputs(28) <= (inputs(245)) or (inputs(205));
    layer0_outputs(29) <= (inputs(117)) or (inputs(102));
    layer0_outputs(30) <= not(inputs(115));
    layer0_outputs(31) <= (inputs(137)) and not (inputs(87));
    layer0_outputs(32) <= not((inputs(73)) and (inputs(28)));
    layer0_outputs(33) <= '0';
    layer0_outputs(34) <= not(inputs(76));
    layer0_outputs(35) <= not(inputs(12)) or (inputs(81));
    layer0_outputs(36) <= not((inputs(125)) or (inputs(94)));
    layer0_outputs(37) <= not(inputs(219)) or (inputs(21));
    layer0_outputs(38) <= not(inputs(212)) or (inputs(61));
    layer0_outputs(39) <= (inputs(49)) xor (inputs(4));
    layer0_outputs(40) <= inputs(196);
    layer0_outputs(41) <= not((inputs(145)) xor (inputs(120)));
    layer0_outputs(42) <= not(inputs(120));
    layer0_outputs(43) <= not(inputs(56)) or (inputs(42));
    layer0_outputs(44) <= not((inputs(217)) or (inputs(190)));
    layer0_outputs(45) <= (inputs(4)) or (inputs(221));
    layer0_outputs(46) <= (inputs(200)) and not (inputs(3));
    layer0_outputs(47) <= not(inputs(120));
    layer0_outputs(48) <= (inputs(230)) and not (inputs(120));
    layer0_outputs(49) <= not(inputs(213));
    layer0_outputs(50) <= '0';
    layer0_outputs(51) <= not(inputs(213)) or (inputs(54));
    layer0_outputs(52) <= not(inputs(133)) or (inputs(166));
    layer0_outputs(53) <= not(inputs(87));
    layer0_outputs(54) <= inputs(151);
    layer0_outputs(55) <= (inputs(129)) and not (inputs(80));
    layer0_outputs(56) <= (inputs(213)) or (inputs(131));
    layer0_outputs(57) <= (inputs(139)) and not (inputs(70));
    layer0_outputs(58) <= '0';
    layer0_outputs(59) <= not((inputs(251)) xor (inputs(107)));
    layer0_outputs(60) <= (inputs(123)) and not (inputs(180));
    layer0_outputs(61) <= not((inputs(213)) and (inputs(151)));
    layer0_outputs(62) <= not((inputs(103)) or (inputs(22)));
    layer0_outputs(63) <= not(inputs(132)) or (inputs(231));
    layer0_outputs(64) <= (inputs(252)) xor (inputs(28));
    layer0_outputs(65) <= not((inputs(94)) xor (inputs(181)));
    layer0_outputs(66) <= inputs(34);
    layer0_outputs(67) <= not(inputs(94));
    layer0_outputs(68) <= '0';
    layer0_outputs(69) <= inputs(133);
    layer0_outputs(70) <= not(inputs(170)) or (inputs(66));
    layer0_outputs(71) <= (inputs(10)) and not (inputs(169));
    layer0_outputs(72) <= (inputs(66)) xor (inputs(49));
    layer0_outputs(73) <= not(inputs(35));
    layer0_outputs(74) <= not(inputs(209));
    layer0_outputs(75) <= not(inputs(100)) or (inputs(9));
    layer0_outputs(76) <= (inputs(175)) xor (inputs(126));
    layer0_outputs(77) <= (inputs(213)) or (inputs(195));
    layer0_outputs(78) <= inputs(6);
    layer0_outputs(79) <= not(inputs(161));
    layer0_outputs(80) <= not(inputs(208));
    layer0_outputs(81) <= inputs(71);
    layer0_outputs(82) <= inputs(109);
    layer0_outputs(83) <= (inputs(8)) and (inputs(9));
    layer0_outputs(84) <= (inputs(159)) xor (inputs(169));
    layer0_outputs(85) <= inputs(176);
    layer0_outputs(86) <= not((inputs(173)) xor (inputs(63)));
    layer0_outputs(87) <= not(inputs(227)) or (inputs(154));
    layer0_outputs(88) <= not((inputs(170)) or (inputs(69)));
    layer0_outputs(89) <= not(inputs(39));
    layer0_outputs(90) <= '1';
    layer0_outputs(91) <= inputs(161);
    layer0_outputs(92) <= (inputs(71)) xor (inputs(23));
    layer0_outputs(93) <= not(inputs(17)) or (inputs(151));
    layer0_outputs(94) <= not(inputs(103));
    layer0_outputs(95) <= inputs(2);
    layer0_outputs(96) <= '1';
    layer0_outputs(97) <= not(inputs(76));
    layer0_outputs(98) <= not((inputs(178)) or (inputs(118)));
    layer0_outputs(99) <= (inputs(87)) and (inputs(95));
    layer0_outputs(100) <= inputs(212);
    layer0_outputs(101) <= '1';
    layer0_outputs(102) <= not(inputs(236)) or (inputs(93));
    layer0_outputs(103) <= not(inputs(233));
    layer0_outputs(104) <= not((inputs(21)) xor (inputs(64)));
    layer0_outputs(105) <= not(inputs(90));
    layer0_outputs(106) <= (inputs(218)) or (inputs(131));
    layer0_outputs(107) <= not((inputs(48)) or (inputs(180)));
    layer0_outputs(108) <= (inputs(128)) and not (inputs(248));
    layer0_outputs(109) <= inputs(131);
    layer0_outputs(110) <= (inputs(133)) or (inputs(213));
    layer0_outputs(111) <= '0';
    layer0_outputs(112) <= not((inputs(40)) xor (inputs(255)));
    layer0_outputs(113) <= not(inputs(228));
    layer0_outputs(114) <= not(inputs(182));
    layer0_outputs(115) <= (inputs(205)) and not (inputs(249));
    layer0_outputs(116) <= (inputs(178)) and not (inputs(67));
    layer0_outputs(117) <= inputs(212);
    layer0_outputs(118) <= inputs(229);
    layer0_outputs(119) <= not(inputs(90)) or (inputs(160));
    layer0_outputs(120) <= not(inputs(35)) or (inputs(25));
    layer0_outputs(121) <= '1';
    layer0_outputs(122) <= (inputs(118)) and not (inputs(15));
    layer0_outputs(123) <= not((inputs(32)) or (inputs(167)));
    layer0_outputs(124) <= not(inputs(50)) or (inputs(202));
    layer0_outputs(125) <= '0';
    layer0_outputs(126) <= not(inputs(227)) or (inputs(108));
    layer0_outputs(127) <= (inputs(52)) and not (inputs(182));
    layer0_outputs(128) <= (inputs(125)) or (inputs(144));
    layer0_outputs(129) <= inputs(190);
    layer0_outputs(130) <= inputs(9);
    layer0_outputs(131) <= not((inputs(245)) or (inputs(10)));
    layer0_outputs(132) <= (inputs(41)) or (inputs(96));
    layer0_outputs(133) <= (inputs(56)) and not (inputs(112));
    layer0_outputs(134) <= '0';
    layer0_outputs(135) <= (inputs(245)) and not (inputs(218));
    layer0_outputs(136) <= inputs(162);
    layer0_outputs(137) <= (inputs(216)) and not (inputs(199));
    layer0_outputs(138) <= not(inputs(26));
    layer0_outputs(139) <= (inputs(83)) xor (inputs(134));
    layer0_outputs(140) <= '0';
    layer0_outputs(141) <= (inputs(51)) or (inputs(91));
    layer0_outputs(142) <= inputs(76);
    layer0_outputs(143) <= not(inputs(57));
    layer0_outputs(144) <= not(inputs(180));
    layer0_outputs(145) <= not((inputs(143)) or (inputs(142)));
    layer0_outputs(146) <= not((inputs(91)) or (inputs(171)));
    layer0_outputs(147) <= not(inputs(108));
    layer0_outputs(148) <= not(inputs(10)) or (inputs(211));
    layer0_outputs(149) <= not(inputs(85));
    layer0_outputs(150) <= not((inputs(138)) and (inputs(98)));
    layer0_outputs(151) <= inputs(109);
    layer0_outputs(152) <= not(inputs(237));
    layer0_outputs(153) <= inputs(205);
    layer0_outputs(154) <= inputs(55);
    layer0_outputs(155) <= inputs(106);
    layer0_outputs(156) <= inputs(25);
    layer0_outputs(157) <= (inputs(11)) and (inputs(217));
    layer0_outputs(158) <= inputs(179);
    layer0_outputs(159) <= inputs(73);
    layer0_outputs(160) <= (inputs(44)) and not (inputs(115));
    layer0_outputs(161) <= not((inputs(131)) and (inputs(60)));
    layer0_outputs(162) <= (inputs(1)) and (inputs(125));
    layer0_outputs(163) <= (inputs(186)) and (inputs(230));
    layer0_outputs(164) <= (inputs(239)) and not (inputs(21));
    layer0_outputs(165) <= (inputs(115)) xor (inputs(7));
    layer0_outputs(166) <= (inputs(102)) xor (inputs(64));
    layer0_outputs(167) <= inputs(25);
    layer0_outputs(168) <= not(inputs(206));
    layer0_outputs(169) <= not(inputs(84)) or (inputs(175));
    layer0_outputs(170) <= (inputs(229)) xor (inputs(159));
    layer0_outputs(171) <= inputs(146);
    layer0_outputs(172) <= not((inputs(100)) xor (inputs(98)));
    layer0_outputs(173) <= (inputs(83)) and not (inputs(254));
    layer0_outputs(174) <= not(inputs(166));
    layer0_outputs(175) <= not((inputs(166)) xor (inputs(95)));
    layer0_outputs(176) <= not((inputs(34)) xor (inputs(203)));
    layer0_outputs(177) <= (inputs(145)) or (inputs(113));
    layer0_outputs(178) <= not(inputs(152));
    layer0_outputs(179) <= not((inputs(195)) or (inputs(254)));
    layer0_outputs(180) <= not(inputs(206));
    layer0_outputs(181) <= not(inputs(148)) or (inputs(253));
    layer0_outputs(182) <= (inputs(151)) xor (inputs(110));
    layer0_outputs(183) <= (inputs(113)) or (inputs(3));
    layer0_outputs(184) <= inputs(194);
    layer0_outputs(185) <= not(inputs(20)) or (inputs(108));
    layer0_outputs(186) <= not(inputs(91));
    layer0_outputs(187) <= (inputs(90)) or (inputs(175));
    layer0_outputs(188) <= not((inputs(111)) or (inputs(26)));
    layer0_outputs(189) <= not((inputs(145)) and (inputs(43)));
    layer0_outputs(190) <= inputs(150);
    layer0_outputs(191) <= (inputs(193)) and not (inputs(209));
    layer0_outputs(192) <= inputs(142);
    layer0_outputs(193) <= inputs(112);
    layer0_outputs(194) <= not(inputs(22));
    layer0_outputs(195) <= (inputs(104)) and not (inputs(145));
    layer0_outputs(196) <= not(inputs(152));
    layer0_outputs(197) <= not((inputs(196)) or (inputs(209)));
    layer0_outputs(198) <= (inputs(238)) xor (inputs(189));
    layer0_outputs(199) <= not(inputs(183)) or (inputs(40));
    layer0_outputs(200) <= not((inputs(64)) xor (inputs(197)));
    layer0_outputs(201) <= not((inputs(178)) and (inputs(57)));
    layer0_outputs(202) <= not((inputs(20)) xor (inputs(14)));
    layer0_outputs(203) <= not(inputs(166));
    layer0_outputs(204) <= (inputs(64)) and not (inputs(253));
    layer0_outputs(205) <= not((inputs(228)) or (inputs(62)));
    layer0_outputs(206) <= (inputs(214)) xor (inputs(174));
    layer0_outputs(207) <= (inputs(15)) and not (inputs(9));
    layer0_outputs(208) <= inputs(99);
    layer0_outputs(209) <= inputs(136);
    layer0_outputs(210) <= inputs(157);
    layer0_outputs(211) <= inputs(225);
    layer0_outputs(212) <= not(inputs(199));
    layer0_outputs(213) <= not(inputs(157));
    layer0_outputs(214) <= (inputs(253)) and not (inputs(113));
    layer0_outputs(215) <= inputs(151);
    layer0_outputs(216) <= '1';
    layer0_outputs(217) <= not((inputs(84)) or (inputs(186)));
    layer0_outputs(218) <= not(inputs(235));
    layer0_outputs(219) <= not((inputs(204)) or (inputs(249)));
    layer0_outputs(220) <= not(inputs(82));
    layer0_outputs(221) <= not((inputs(86)) xor (inputs(66)));
    layer0_outputs(222) <= not((inputs(247)) or (inputs(192)));
    layer0_outputs(223) <= inputs(229);
    layer0_outputs(224) <= not(inputs(155));
    layer0_outputs(225) <= (inputs(10)) xor (inputs(4));
    layer0_outputs(226) <= not(inputs(9)) or (inputs(16));
    layer0_outputs(227) <= not(inputs(162)) or (inputs(150));
    layer0_outputs(228) <= not((inputs(35)) xor (inputs(105)));
    layer0_outputs(229) <= not((inputs(161)) xor (inputs(165)));
    layer0_outputs(230) <= not((inputs(249)) or (inputs(253)));
    layer0_outputs(231) <= (inputs(163)) or (inputs(206));
    layer0_outputs(232) <= inputs(205);
    layer0_outputs(233) <= not(inputs(115));
    layer0_outputs(234) <= (inputs(144)) xor (inputs(40));
    layer0_outputs(235) <= (inputs(13)) and not (inputs(130));
    layer0_outputs(236) <= not((inputs(224)) or (inputs(161)));
    layer0_outputs(237) <= (inputs(29)) or (inputs(213));
    layer0_outputs(238) <= not((inputs(156)) or (inputs(236)));
    layer0_outputs(239) <= (inputs(104)) and not (inputs(213));
    layer0_outputs(240) <= not(inputs(75));
    layer0_outputs(241) <= not(inputs(100));
    layer0_outputs(242) <= not(inputs(41));
    layer0_outputs(243) <= (inputs(93)) or (inputs(26));
    layer0_outputs(244) <= not((inputs(248)) and (inputs(129)));
    layer0_outputs(245) <= inputs(194);
    layer0_outputs(246) <= not(inputs(70));
    layer0_outputs(247) <= not((inputs(209)) xor (inputs(108)));
    layer0_outputs(248) <= not((inputs(117)) xor (inputs(69)));
    layer0_outputs(249) <= not(inputs(183)) or (inputs(46));
    layer0_outputs(250) <= inputs(136);
    layer0_outputs(251) <= not((inputs(158)) xor (inputs(108)));
    layer0_outputs(252) <= (inputs(17)) xor (inputs(32));
    layer0_outputs(253) <= not((inputs(25)) xor (inputs(176)));
    layer0_outputs(254) <= not(inputs(221));
    layer0_outputs(255) <= (inputs(202)) and not (inputs(163));
    layer0_outputs(256) <= (inputs(37)) or (inputs(46));
    layer0_outputs(257) <= not((inputs(114)) or (inputs(83)));
    layer0_outputs(258) <= (inputs(122)) xor (inputs(174));
    layer0_outputs(259) <= '1';
    layer0_outputs(260) <= (inputs(199)) and not (inputs(96));
    layer0_outputs(261) <= not((inputs(102)) and (inputs(193)));
    layer0_outputs(262) <= not(inputs(161)) or (inputs(192));
    layer0_outputs(263) <= (inputs(220)) or (inputs(223));
    layer0_outputs(264) <= inputs(21);
    layer0_outputs(265) <= (inputs(88)) and not (inputs(255));
    layer0_outputs(266) <= (inputs(84)) and not (inputs(72));
    layer0_outputs(267) <= (inputs(229)) xor (inputs(19));
    layer0_outputs(268) <= not((inputs(207)) or (inputs(119)));
    layer0_outputs(269) <= inputs(178);
    layer0_outputs(270) <= (inputs(22)) or (inputs(61));
    layer0_outputs(271) <= not(inputs(77));
    layer0_outputs(272) <= not((inputs(136)) xor (inputs(103)));
    layer0_outputs(273) <= inputs(230);
    layer0_outputs(274) <= (inputs(197)) and not (inputs(4));
    layer0_outputs(275) <= not(inputs(136));
    layer0_outputs(276) <= not(inputs(76));
    layer0_outputs(277) <= not((inputs(100)) and (inputs(106)));
    layer0_outputs(278) <= not(inputs(45));
    layer0_outputs(279) <= inputs(145);
    layer0_outputs(280) <= inputs(164);
    layer0_outputs(281) <= not((inputs(98)) xor (inputs(154)));
    layer0_outputs(282) <= not(inputs(79)) or (inputs(172));
    layer0_outputs(283) <= not(inputs(137));
    layer0_outputs(284) <= not((inputs(141)) xor (inputs(46)));
    layer0_outputs(285) <= inputs(22);
    layer0_outputs(286) <= not(inputs(162));
    layer0_outputs(287) <= (inputs(23)) and not (inputs(29));
    layer0_outputs(288) <= not(inputs(249)) or (inputs(64));
    layer0_outputs(289) <= (inputs(8)) or (inputs(239));
    layer0_outputs(290) <= inputs(165);
    layer0_outputs(291) <= not((inputs(98)) or (inputs(126)));
    layer0_outputs(292) <= not(inputs(42)) or (inputs(184));
    layer0_outputs(293) <= not(inputs(81));
    layer0_outputs(294) <= not(inputs(137));
    layer0_outputs(295) <= '0';
    layer0_outputs(296) <= not(inputs(72)) or (inputs(5));
    layer0_outputs(297) <= '0';
    layer0_outputs(298) <= inputs(170);
    layer0_outputs(299) <= not((inputs(63)) xor (inputs(42)));
    layer0_outputs(300) <= not(inputs(99)) or (inputs(235));
    layer0_outputs(301) <= (inputs(56)) or (inputs(13));
    layer0_outputs(302) <= inputs(29);
    layer0_outputs(303) <= (inputs(137)) xor (inputs(131));
    layer0_outputs(304) <= inputs(137);
    layer0_outputs(305) <= (inputs(174)) or (inputs(75));
    layer0_outputs(306) <= not((inputs(197)) or (inputs(128)));
    layer0_outputs(307) <= (inputs(26)) or (inputs(3));
    layer0_outputs(308) <= not((inputs(4)) and (inputs(67)));
    layer0_outputs(309) <= not(inputs(147));
    layer0_outputs(310) <= not((inputs(185)) and (inputs(141)));
    layer0_outputs(311) <= not(inputs(97));
    layer0_outputs(312) <= not((inputs(240)) and (inputs(184)));
    layer0_outputs(313) <= not(inputs(143));
    layer0_outputs(314) <= not(inputs(184));
    layer0_outputs(315) <= not((inputs(59)) or (inputs(15)));
    layer0_outputs(316) <= inputs(236);
    layer0_outputs(317) <= not(inputs(151)) or (inputs(63));
    layer0_outputs(318) <= (inputs(150)) and not (inputs(12));
    layer0_outputs(319) <= not((inputs(208)) or (inputs(31)));
    layer0_outputs(320) <= '1';
    layer0_outputs(321) <= inputs(253);
    layer0_outputs(322) <= not((inputs(145)) xor (inputs(238)));
    layer0_outputs(323) <= inputs(15);
    layer0_outputs(324) <= not((inputs(86)) and (inputs(31)));
    layer0_outputs(325) <= (inputs(90)) and not (inputs(176));
    layer0_outputs(326) <= inputs(100);
    layer0_outputs(327) <= (inputs(119)) or (inputs(174));
    layer0_outputs(328) <= (inputs(112)) or (inputs(132));
    layer0_outputs(329) <= not(inputs(173)) or (inputs(22));
    layer0_outputs(330) <= inputs(63);
    layer0_outputs(331) <= (inputs(194)) or (inputs(237));
    layer0_outputs(332) <= not(inputs(158)) or (inputs(81));
    layer0_outputs(333) <= not(inputs(38));
    layer0_outputs(334) <= (inputs(139)) or (inputs(43));
    layer0_outputs(335) <= not((inputs(45)) or (inputs(238)));
    layer0_outputs(336) <= not(inputs(215));
    layer0_outputs(337) <= (inputs(172)) and (inputs(233));
    layer0_outputs(338) <= (inputs(104)) and not (inputs(197));
    layer0_outputs(339) <= not((inputs(188)) or (inputs(16)));
    layer0_outputs(340) <= (inputs(215)) and not (inputs(131));
    layer0_outputs(341) <= not(inputs(42)) or (inputs(204));
    layer0_outputs(342) <= (inputs(161)) and not (inputs(67));
    layer0_outputs(343) <= not((inputs(60)) and (inputs(81)));
    layer0_outputs(344) <= '1';
    layer0_outputs(345) <= inputs(13);
    layer0_outputs(346) <= not(inputs(254)) or (inputs(166));
    layer0_outputs(347) <= (inputs(65)) xor (inputs(90));
    layer0_outputs(348) <= (inputs(140)) or (inputs(73));
    layer0_outputs(349) <= not(inputs(41));
    layer0_outputs(350) <= not(inputs(196)) or (inputs(34));
    layer0_outputs(351) <= not((inputs(110)) or (inputs(240)));
    layer0_outputs(352) <= not(inputs(22)) or (inputs(152));
    layer0_outputs(353) <= not((inputs(54)) xor (inputs(37)));
    layer0_outputs(354) <= not(inputs(248));
    layer0_outputs(355) <= not(inputs(109));
    layer0_outputs(356) <= not(inputs(103)) or (inputs(127));
    layer0_outputs(357) <= (inputs(30)) and not (inputs(79));
    layer0_outputs(358) <= inputs(155);
    layer0_outputs(359) <= not((inputs(75)) or (inputs(200)));
    layer0_outputs(360) <= not(inputs(102)) or (inputs(1));
    layer0_outputs(361) <= inputs(137);
    layer0_outputs(362) <= (inputs(84)) xor (inputs(81));
    layer0_outputs(363) <= inputs(98);
    layer0_outputs(364) <= (inputs(21)) xor (inputs(93));
    layer0_outputs(365) <= not((inputs(186)) and (inputs(58)));
    layer0_outputs(366) <= not(inputs(88)) or (inputs(191));
    layer0_outputs(367) <= inputs(85);
    layer0_outputs(368) <= (inputs(206)) and not (inputs(13));
    layer0_outputs(369) <= (inputs(146)) and (inputs(219));
    layer0_outputs(370) <= not(inputs(229));
    layer0_outputs(371) <= '1';
    layer0_outputs(372) <= not(inputs(104));
    layer0_outputs(373) <= inputs(90);
    layer0_outputs(374) <= not(inputs(115));
    layer0_outputs(375) <= (inputs(20)) and (inputs(206));
    layer0_outputs(376) <= (inputs(237)) xor (inputs(206));
    layer0_outputs(377) <= inputs(6);
    layer0_outputs(378) <= (inputs(51)) or (inputs(255));
    layer0_outputs(379) <= (inputs(35)) xor (inputs(72));
    layer0_outputs(380) <= not(inputs(93));
    layer0_outputs(381) <= not(inputs(11)) or (inputs(28));
    layer0_outputs(382) <= (inputs(194)) and not (inputs(0));
    layer0_outputs(383) <= not(inputs(110)) or (inputs(95));
    layer0_outputs(384) <= (inputs(236)) or (inputs(103));
    layer0_outputs(385) <= (inputs(49)) or (inputs(25));
    layer0_outputs(386) <= not(inputs(6));
    layer0_outputs(387) <= not(inputs(78));
    layer0_outputs(388) <= inputs(94);
    layer0_outputs(389) <= (inputs(197)) and (inputs(255));
    layer0_outputs(390) <= (inputs(39)) xor (inputs(120));
    layer0_outputs(391) <= not((inputs(98)) xor (inputs(68)));
    layer0_outputs(392) <= not(inputs(228)) or (inputs(254));
    layer0_outputs(393) <= not(inputs(94));
    layer0_outputs(394) <= (inputs(223)) xor (inputs(191));
    layer0_outputs(395) <= inputs(133);
    layer0_outputs(396) <= not((inputs(244)) xor (inputs(106)));
    layer0_outputs(397) <= not(inputs(230)) or (inputs(54));
    layer0_outputs(398) <= not((inputs(114)) or (inputs(30)));
    layer0_outputs(399) <= inputs(229);
    layer0_outputs(400) <= (inputs(164)) and (inputs(125));
    layer0_outputs(401) <= not(inputs(146));
    layer0_outputs(402) <= inputs(43);
    layer0_outputs(403) <= not(inputs(185));
    layer0_outputs(404) <= not((inputs(208)) or (inputs(154)));
    layer0_outputs(405) <= not((inputs(22)) or (inputs(236)));
    layer0_outputs(406) <= (inputs(92)) and not (inputs(255));
    layer0_outputs(407) <= not(inputs(74));
    layer0_outputs(408) <= not(inputs(232));
    layer0_outputs(409) <= not(inputs(234));
    layer0_outputs(410) <= not(inputs(169));
    layer0_outputs(411) <= (inputs(48)) and not (inputs(179));
    layer0_outputs(412) <= (inputs(38)) and (inputs(229));
    layer0_outputs(413) <= (inputs(108)) xor (inputs(4));
    layer0_outputs(414) <= not(inputs(172)) or (inputs(133));
    layer0_outputs(415) <= (inputs(242)) or (inputs(212));
    layer0_outputs(416) <= (inputs(3)) and not (inputs(141));
    layer0_outputs(417) <= not((inputs(123)) xor (inputs(132)));
    layer0_outputs(418) <= (inputs(88)) and not (inputs(208));
    layer0_outputs(419) <= not(inputs(160));
    layer0_outputs(420) <= '0';
    layer0_outputs(421) <= not((inputs(32)) or (inputs(231)));
    layer0_outputs(422) <= inputs(105);
    layer0_outputs(423) <= (inputs(63)) or (inputs(45));
    layer0_outputs(424) <= not(inputs(218));
    layer0_outputs(425) <= (inputs(52)) and not (inputs(4));
    layer0_outputs(426) <= (inputs(140)) xor (inputs(175));
    layer0_outputs(427) <= not((inputs(100)) xor (inputs(3)));
    layer0_outputs(428) <= (inputs(142)) or (inputs(29));
    layer0_outputs(429) <= inputs(214);
    layer0_outputs(430) <= not(inputs(83)) or (inputs(252));
    layer0_outputs(431) <= (inputs(95)) xor (inputs(57));
    layer0_outputs(432) <= (inputs(34)) xor (inputs(97));
    layer0_outputs(433) <= (inputs(88)) or (inputs(106));
    layer0_outputs(434) <= (inputs(111)) xor (inputs(45));
    layer0_outputs(435) <= (inputs(55)) or (inputs(175));
    layer0_outputs(436) <= not(inputs(57));
    layer0_outputs(437) <= (inputs(219)) and not (inputs(94));
    layer0_outputs(438) <= (inputs(63)) and not (inputs(227));
    layer0_outputs(439) <= (inputs(29)) and not (inputs(70));
    layer0_outputs(440) <= not(inputs(165));
    layer0_outputs(441) <= not(inputs(119));
    layer0_outputs(442) <= (inputs(156)) and not (inputs(126));
    layer0_outputs(443) <= not((inputs(79)) or (inputs(104)));
    layer0_outputs(444) <= (inputs(237)) and (inputs(67));
    layer0_outputs(445) <= not((inputs(253)) xor (inputs(87)));
    layer0_outputs(446) <= inputs(111);
    layer0_outputs(447) <= inputs(182);
    layer0_outputs(448) <= (inputs(151)) xor (inputs(33));
    layer0_outputs(449) <= not((inputs(237)) or (inputs(87)));
    layer0_outputs(450) <= not((inputs(144)) xor (inputs(201)));
    layer0_outputs(451) <= (inputs(121)) and not (inputs(48));
    layer0_outputs(452) <= (inputs(21)) and (inputs(102));
    layer0_outputs(453) <= '1';
    layer0_outputs(454) <= not((inputs(42)) and (inputs(240)));
    layer0_outputs(455) <= (inputs(216)) and not (inputs(56));
    layer0_outputs(456) <= not((inputs(43)) and (inputs(29)));
    layer0_outputs(457) <= (inputs(123)) or (inputs(227));
    layer0_outputs(458) <= (inputs(199)) or (inputs(60));
    layer0_outputs(459) <= not(inputs(102));
    layer0_outputs(460) <= not((inputs(122)) and (inputs(43)));
    layer0_outputs(461) <= '1';
    layer0_outputs(462) <= not(inputs(188));
    layer0_outputs(463) <= not(inputs(61));
    layer0_outputs(464) <= not(inputs(37));
    layer0_outputs(465) <= not(inputs(129));
    layer0_outputs(466) <= (inputs(71)) or (inputs(148));
    layer0_outputs(467) <= (inputs(74)) and not (inputs(254));
    layer0_outputs(468) <= (inputs(9)) and not (inputs(208));
    layer0_outputs(469) <= not(inputs(26)) or (inputs(181));
    layer0_outputs(470) <= (inputs(64)) and (inputs(77));
    layer0_outputs(471) <= (inputs(72)) xor (inputs(179));
    layer0_outputs(472) <= not((inputs(89)) xor (inputs(28)));
    layer0_outputs(473) <= not(inputs(250));
    layer0_outputs(474) <= not(inputs(171)) or (inputs(35));
    layer0_outputs(475) <= '0';
    layer0_outputs(476) <= not(inputs(27));
    layer0_outputs(477) <= not(inputs(134)) or (inputs(31));
    layer0_outputs(478) <= (inputs(3)) and (inputs(210));
    layer0_outputs(479) <= (inputs(167)) or (inputs(110));
    layer0_outputs(480) <= not(inputs(15));
    layer0_outputs(481) <= not((inputs(179)) xor (inputs(174)));
    layer0_outputs(482) <= (inputs(7)) and not (inputs(44));
    layer0_outputs(483) <= not((inputs(225)) or (inputs(201)));
    layer0_outputs(484) <= '1';
    layer0_outputs(485) <= not((inputs(52)) or (inputs(111)));
    layer0_outputs(486) <= (inputs(36)) xor (inputs(71));
    layer0_outputs(487) <= (inputs(223)) or (inputs(82));
    layer0_outputs(488) <= (inputs(38)) and not (inputs(153));
    layer0_outputs(489) <= not(inputs(94));
    layer0_outputs(490) <= (inputs(3)) xor (inputs(99));
    layer0_outputs(491) <= not((inputs(158)) or (inputs(183)));
    layer0_outputs(492) <= not((inputs(36)) or (inputs(76)));
    layer0_outputs(493) <= not((inputs(157)) or (inputs(173)));
    layer0_outputs(494) <= (inputs(160)) and not (inputs(14));
    layer0_outputs(495) <= not((inputs(174)) or (inputs(132)));
    layer0_outputs(496) <= not(inputs(229));
    layer0_outputs(497) <= inputs(251);
    layer0_outputs(498) <= (inputs(237)) or (inputs(186));
    layer0_outputs(499) <= (inputs(130)) and not (inputs(121));
    layer0_outputs(500) <= (inputs(135)) and not (inputs(231));
    layer0_outputs(501) <= not(inputs(134));
    layer0_outputs(502) <= inputs(249);
    layer0_outputs(503) <= not((inputs(192)) or (inputs(77)));
    layer0_outputs(504) <= (inputs(7)) or (inputs(219));
    layer0_outputs(505) <= (inputs(67)) xor (inputs(204));
    layer0_outputs(506) <= inputs(63);
    layer0_outputs(507) <= (inputs(119)) and not (inputs(241));
    layer0_outputs(508) <= not(inputs(83)) or (inputs(24));
    layer0_outputs(509) <= '1';
    layer0_outputs(510) <= not((inputs(190)) or (inputs(181)));
    layer0_outputs(511) <= not(inputs(40)) or (inputs(185));
    layer0_outputs(512) <= not(inputs(202));
    layer0_outputs(513) <= not((inputs(240)) xor (inputs(156)));
    layer0_outputs(514) <= not(inputs(16));
    layer0_outputs(515) <= (inputs(67)) or (inputs(82));
    layer0_outputs(516) <= not((inputs(54)) xor (inputs(105)));
    layer0_outputs(517) <= not(inputs(56)) or (inputs(241));
    layer0_outputs(518) <= '0';
    layer0_outputs(519) <= not((inputs(177)) xor (inputs(209)));
    layer0_outputs(520) <= (inputs(202)) and not (inputs(175));
    layer0_outputs(521) <= not((inputs(214)) and (inputs(222)));
    layer0_outputs(522) <= not(inputs(170));
    layer0_outputs(523) <= inputs(87);
    layer0_outputs(524) <= not((inputs(21)) xor (inputs(255)));
    layer0_outputs(525) <= not((inputs(12)) xor (inputs(171)));
    layer0_outputs(526) <= not((inputs(168)) or (inputs(210)));
    layer0_outputs(527) <= not(inputs(158));
    layer0_outputs(528) <= inputs(162);
    layer0_outputs(529) <= (inputs(153)) and not (inputs(54));
    layer0_outputs(530) <= (inputs(133)) or (inputs(84));
    layer0_outputs(531) <= not(inputs(20)) or (inputs(232));
    layer0_outputs(532) <= not(inputs(204)) or (inputs(30));
    layer0_outputs(533) <= not((inputs(169)) and (inputs(163)));
    layer0_outputs(534) <= '1';
    layer0_outputs(535) <= not(inputs(82));
    layer0_outputs(536) <= not(inputs(255)) or (inputs(59));
    layer0_outputs(537) <= '0';
    layer0_outputs(538) <= not(inputs(71)) or (inputs(16));
    layer0_outputs(539) <= not(inputs(148)) or (inputs(26));
    layer0_outputs(540) <= (inputs(247)) and not (inputs(77));
    layer0_outputs(541) <= (inputs(242)) or (inputs(210));
    layer0_outputs(542) <= inputs(107);
    layer0_outputs(543) <= not((inputs(129)) xor (inputs(138)));
    layer0_outputs(544) <= (inputs(50)) and not (inputs(45));
    layer0_outputs(545) <= (inputs(251)) or (inputs(212));
    layer0_outputs(546) <= (inputs(241)) or (inputs(135));
    layer0_outputs(547) <= not((inputs(51)) or (inputs(118)));
    layer0_outputs(548) <= inputs(166);
    layer0_outputs(549) <= not(inputs(105));
    layer0_outputs(550) <= not((inputs(171)) and (inputs(200)));
    layer0_outputs(551) <= not(inputs(78));
    layer0_outputs(552) <= (inputs(189)) xor (inputs(110));
    layer0_outputs(553) <= not(inputs(253));
    layer0_outputs(554) <= (inputs(218)) xor (inputs(124));
    layer0_outputs(555) <= not(inputs(172));
    layer0_outputs(556) <= (inputs(22)) or (inputs(213));
    layer0_outputs(557) <= not((inputs(31)) and (inputs(233)));
    layer0_outputs(558) <= not(inputs(113));
    layer0_outputs(559) <= inputs(100);
    layer0_outputs(560) <= not((inputs(0)) or (inputs(149)));
    layer0_outputs(561) <= (inputs(226)) or (inputs(65));
    layer0_outputs(562) <= not(inputs(25));
    layer0_outputs(563) <= not(inputs(100)) or (inputs(164));
    layer0_outputs(564) <= inputs(215);
    layer0_outputs(565) <= (inputs(115)) and not (inputs(58));
    layer0_outputs(566) <= (inputs(86)) xor (inputs(229));
    layer0_outputs(567) <= not(inputs(10));
    layer0_outputs(568) <= not((inputs(88)) and (inputs(54)));
    layer0_outputs(569) <= not((inputs(73)) xor (inputs(95)));
    layer0_outputs(570) <= not((inputs(212)) or (inputs(223)));
    layer0_outputs(571) <= (inputs(102)) and not (inputs(88));
    layer0_outputs(572) <= (inputs(88)) or (inputs(48));
    layer0_outputs(573) <= (inputs(223)) or (inputs(218));
    layer0_outputs(574) <= not(inputs(191));
    layer0_outputs(575) <= not(inputs(127));
    layer0_outputs(576) <= not(inputs(145));
    layer0_outputs(577) <= not((inputs(72)) xor (inputs(179)));
    layer0_outputs(578) <= (inputs(120)) or (inputs(44));
    layer0_outputs(579) <= not((inputs(67)) xor (inputs(24)));
    layer0_outputs(580) <= not((inputs(203)) xor (inputs(157)));
    layer0_outputs(581) <= inputs(114);
    layer0_outputs(582) <= not((inputs(176)) or (inputs(206)));
    layer0_outputs(583) <= (inputs(18)) xor (inputs(238));
    layer0_outputs(584) <= not((inputs(147)) or (inputs(180)));
    layer0_outputs(585) <= not((inputs(57)) or (inputs(161)));
    layer0_outputs(586) <= not(inputs(13));
    layer0_outputs(587) <= (inputs(136)) and (inputs(233));
    layer0_outputs(588) <= not(inputs(154));
    layer0_outputs(589) <= (inputs(37)) and not (inputs(143));
    layer0_outputs(590) <= not((inputs(45)) xor (inputs(251)));
    layer0_outputs(591) <= not(inputs(154));
    layer0_outputs(592) <= not((inputs(160)) or (inputs(76)));
    layer0_outputs(593) <= (inputs(223)) xor (inputs(108));
    layer0_outputs(594) <= (inputs(242)) or (inputs(225));
    layer0_outputs(595) <= inputs(221);
    layer0_outputs(596) <= (inputs(253)) and not (inputs(51));
    layer0_outputs(597) <= (inputs(51)) and not (inputs(165));
    layer0_outputs(598) <= not(inputs(90)) or (inputs(244));
    layer0_outputs(599) <= (inputs(246)) and not (inputs(17));
    layer0_outputs(600) <= inputs(60);
    layer0_outputs(601) <= not((inputs(212)) or (inputs(76)));
    layer0_outputs(602) <= not(inputs(162));
    layer0_outputs(603) <= (inputs(36)) or (inputs(12));
    layer0_outputs(604) <= not((inputs(89)) xor (inputs(91)));
    layer0_outputs(605) <= (inputs(55)) xor (inputs(99));
    layer0_outputs(606) <= (inputs(105)) and not (inputs(22));
    layer0_outputs(607) <= inputs(102);
    layer0_outputs(608) <= inputs(109);
    layer0_outputs(609) <= not(inputs(72));
    layer0_outputs(610) <= not((inputs(184)) xor (inputs(178)));
    layer0_outputs(611) <= '1';
    layer0_outputs(612) <= not(inputs(85));
    layer0_outputs(613) <= not(inputs(76));
    layer0_outputs(614) <= not(inputs(247));
    layer0_outputs(615) <= not(inputs(167)) or (inputs(150));
    layer0_outputs(616) <= (inputs(68)) xor (inputs(115));
    layer0_outputs(617) <= not(inputs(114));
    layer0_outputs(618) <= not(inputs(111)) or (inputs(169));
    layer0_outputs(619) <= not((inputs(130)) and (inputs(57)));
    layer0_outputs(620) <= (inputs(25)) and not (inputs(126));
    layer0_outputs(621) <= (inputs(188)) xor (inputs(109));
    layer0_outputs(622) <= not(inputs(84)) or (inputs(209));
    layer0_outputs(623) <= (inputs(216)) and (inputs(204));
    layer0_outputs(624) <= (inputs(99)) or (inputs(45));
    layer0_outputs(625) <= not((inputs(24)) or (inputs(5)));
    layer0_outputs(626) <= inputs(68);
    layer0_outputs(627) <= not(inputs(2));
    layer0_outputs(628) <= inputs(13);
    layer0_outputs(629) <= (inputs(56)) or (inputs(245));
    layer0_outputs(630) <= not((inputs(187)) xor (inputs(36)));
    layer0_outputs(631) <= inputs(202);
    layer0_outputs(632) <= (inputs(103)) and not (inputs(192));
    layer0_outputs(633) <= '1';
    layer0_outputs(634) <= (inputs(32)) or (inputs(220));
    layer0_outputs(635) <= (inputs(58)) xor (inputs(214));
    layer0_outputs(636) <= '1';
    layer0_outputs(637) <= inputs(5);
    layer0_outputs(638) <= not(inputs(18)) or (inputs(221));
    layer0_outputs(639) <= not(inputs(69)) or (inputs(144));
    layer0_outputs(640) <= (inputs(225)) and not (inputs(31));
    layer0_outputs(641) <= not(inputs(38));
    layer0_outputs(642) <= (inputs(208)) and not (inputs(77));
    layer0_outputs(643) <= '0';
    layer0_outputs(644) <= '1';
    layer0_outputs(645) <= not(inputs(118)) or (inputs(137));
    layer0_outputs(646) <= not(inputs(81));
    layer0_outputs(647) <= not(inputs(28));
    layer0_outputs(648) <= (inputs(1)) xor (inputs(166));
    layer0_outputs(649) <= not((inputs(173)) or (inputs(232)));
    layer0_outputs(650) <= not(inputs(102));
    layer0_outputs(651) <= '0';
    layer0_outputs(652) <= not(inputs(26));
    layer0_outputs(653) <= (inputs(100)) or (inputs(199));
    layer0_outputs(654) <= inputs(193);
    layer0_outputs(655) <= inputs(41);
    layer0_outputs(656) <= not(inputs(181));
    layer0_outputs(657) <= not((inputs(184)) and (inputs(164)));
    layer0_outputs(658) <= not((inputs(169)) or (inputs(142)));
    layer0_outputs(659) <= not(inputs(208));
    layer0_outputs(660) <= not((inputs(41)) or (inputs(75)));
    layer0_outputs(661) <= '1';
    layer0_outputs(662) <= (inputs(84)) or (inputs(80));
    layer0_outputs(663) <= not((inputs(112)) or (inputs(37)));
    layer0_outputs(664) <= (inputs(182)) and (inputs(121));
    layer0_outputs(665) <= not(inputs(196));
    layer0_outputs(666) <= not(inputs(145)) or (inputs(240));
    layer0_outputs(667) <= inputs(166);
    layer0_outputs(668) <= not((inputs(254)) or (inputs(174)));
    layer0_outputs(669) <= not(inputs(154));
    layer0_outputs(670) <= not((inputs(2)) or (inputs(18)));
    layer0_outputs(671) <= inputs(164);
    layer0_outputs(672) <= (inputs(205)) and (inputs(44));
    layer0_outputs(673) <= not(inputs(27)) or (inputs(83));
    layer0_outputs(674) <= (inputs(207)) or (inputs(110));
    layer0_outputs(675) <= (inputs(168)) or (inputs(144));
    layer0_outputs(676) <= not(inputs(53)) or (inputs(17));
    layer0_outputs(677) <= inputs(178);
    layer0_outputs(678) <= (inputs(13)) xor (inputs(44));
    layer0_outputs(679) <= inputs(9);
    layer0_outputs(680) <= (inputs(12)) and not (inputs(220));
    layer0_outputs(681) <= not(inputs(113));
    layer0_outputs(682) <= (inputs(225)) xor (inputs(195));
    layer0_outputs(683) <= not((inputs(126)) xor (inputs(143)));
    layer0_outputs(684) <= inputs(204);
    layer0_outputs(685) <= inputs(230);
    layer0_outputs(686) <= (inputs(9)) and not (inputs(137));
    layer0_outputs(687) <= not((inputs(58)) and (inputs(157)));
    layer0_outputs(688) <= '1';
    layer0_outputs(689) <= (inputs(79)) and not (inputs(105));
    layer0_outputs(690) <= inputs(90);
    layer0_outputs(691) <= (inputs(62)) and (inputs(95));
    layer0_outputs(692) <= (inputs(18)) xor (inputs(153));
    layer0_outputs(693) <= not(inputs(140)) or (inputs(72));
    layer0_outputs(694) <= (inputs(208)) and not (inputs(124));
    layer0_outputs(695) <= '0';
    layer0_outputs(696) <= (inputs(101)) xor (inputs(198));
    layer0_outputs(697) <= inputs(63);
    layer0_outputs(698) <= (inputs(212)) or (inputs(104));
    layer0_outputs(699) <= (inputs(169)) xor (inputs(118));
    layer0_outputs(700) <= '0';
    layer0_outputs(701) <= (inputs(10)) and not (inputs(217));
    layer0_outputs(702) <= inputs(127);
    layer0_outputs(703) <= not(inputs(99));
    layer0_outputs(704) <= (inputs(87)) and not (inputs(221));
    layer0_outputs(705) <= not(inputs(117));
    layer0_outputs(706) <= inputs(154);
    layer0_outputs(707) <= not(inputs(174));
    layer0_outputs(708) <= (inputs(209)) and (inputs(116));
    layer0_outputs(709) <= not((inputs(189)) or (inputs(23)));
    layer0_outputs(710) <= not(inputs(108)) or (inputs(133));
    layer0_outputs(711) <= (inputs(230)) and not (inputs(80));
    layer0_outputs(712) <= not(inputs(100)) or (inputs(94));
    layer0_outputs(713) <= not((inputs(208)) or (inputs(163)));
    layer0_outputs(714) <= not(inputs(159)) or (inputs(13));
    layer0_outputs(715) <= (inputs(243)) or (inputs(204));
    layer0_outputs(716) <= not((inputs(219)) or (inputs(215)));
    layer0_outputs(717) <= (inputs(110)) xor (inputs(14));
    layer0_outputs(718) <= not(inputs(24));
    layer0_outputs(719) <= inputs(22);
    layer0_outputs(720) <= (inputs(74)) and not (inputs(252));
    layer0_outputs(721) <= (inputs(254)) and not (inputs(40));
    layer0_outputs(722) <= not((inputs(27)) xor (inputs(153)));
    layer0_outputs(723) <= not(inputs(90));
    layer0_outputs(724) <= not(inputs(59)) or (inputs(71));
    layer0_outputs(725) <= not(inputs(85));
    layer0_outputs(726) <= (inputs(170)) or (inputs(98));
    layer0_outputs(727) <= (inputs(98)) xor (inputs(115));
    layer0_outputs(728) <= not(inputs(119)) or (inputs(178));
    layer0_outputs(729) <= not((inputs(246)) xor (inputs(215)));
    layer0_outputs(730) <= not(inputs(179)) or (inputs(94));
    layer0_outputs(731) <= not(inputs(48));
    layer0_outputs(732) <= not(inputs(244));
    layer0_outputs(733) <= (inputs(251)) xor (inputs(105));
    layer0_outputs(734) <= not(inputs(38));
    layer0_outputs(735) <= (inputs(237)) and not (inputs(128));
    layer0_outputs(736) <= (inputs(214)) xor (inputs(212));
    layer0_outputs(737) <= not((inputs(47)) and (inputs(32)));
    layer0_outputs(738) <= not(inputs(141));
    layer0_outputs(739) <= inputs(33);
    layer0_outputs(740) <= (inputs(156)) and not (inputs(153));
    layer0_outputs(741) <= (inputs(150)) and not (inputs(220));
    layer0_outputs(742) <= (inputs(147)) xor (inputs(113));
    layer0_outputs(743) <= '0';
    layer0_outputs(744) <= inputs(69);
    layer0_outputs(745) <= (inputs(150)) and not (inputs(249));
    layer0_outputs(746) <= not((inputs(143)) or (inputs(138)));
    layer0_outputs(747) <= (inputs(239)) and not (inputs(250));
    layer0_outputs(748) <= inputs(234);
    layer0_outputs(749) <= not((inputs(72)) and (inputs(72)));
    layer0_outputs(750) <= inputs(168);
    layer0_outputs(751) <= not((inputs(25)) xor (inputs(220)));
    layer0_outputs(752) <= not((inputs(251)) or (inputs(198)));
    layer0_outputs(753) <= (inputs(173)) xor (inputs(68));
    layer0_outputs(754) <= (inputs(158)) or (inputs(225));
    layer0_outputs(755) <= not((inputs(248)) or (inputs(229)));
    layer0_outputs(756) <= (inputs(196)) xor (inputs(110));
    layer0_outputs(757) <= (inputs(116)) and not (inputs(245));
    layer0_outputs(758) <= (inputs(220)) xor (inputs(192));
    layer0_outputs(759) <= (inputs(62)) xor (inputs(122));
    layer0_outputs(760) <= (inputs(182)) and not (inputs(58));
    layer0_outputs(761) <= (inputs(183)) and not (inputs(130));
    layer0_outputs(762) <= inputs(235);
    layer0_outputs(763) <= not(inputs(104));
    layer0_outputs(764) <= not((inputs(64)) xor (inputs(173)));
    layer0_outputs(765) <= (inputs(184)) or (inputs(170));
    layer0_outputs(766) <= (inputs(137)) and not (inputs(48));
    layer0_outputs(767) <= inputs(23);
    layer0_outputs(768) <= inputs(154);
    layer0_outputs(769) <= (inputs(79)) or (inputs(178));
    layer0_outputs(770) <= (inputs(213)) and (inputs(71));
    layer0_outputs(771) <= (inputs(48)) xor (inputs(137));
    layer0_outputs(772) <= not(inputs(156)) or (inputs(37));
    layer0_outputs(773) <= not((inputs(194)) or (inputs(4)));
    layer0_outputs(774) <= not((inputs(210)) and (inputs(143)));
    layer0_outputs(775) <= (inputs(191)) and not (inputs(223));
    layer0_outputs(776) <= (inputs(83)) or (inputs(69));
    layer0_outputs(777) <= inputs(187);
    layer0_outputs(778) <= inputs(234);
    layer0_outputs(779) <= not(inputs(141)) or (inputs(44));
    layer0_outputs(780) <= not(inputs(79));
    layer0_outputs(781) <= not(inputs(76)) or (inputs(197));
    layer0_outputs(782) <= not(inputs(43));
    layer0_outputs(783) <= not(inputs(181)) or (inputs(166));
    layer0_outputs(784) <= not((inputs(154)) or (inputs(163)));
    layer0_outputs(785) <= inputs(45);
    layer0_outputs(786) <= inputs(166);
    layer0_outputs(787) <= (inputs(26)) or (inputs(208));
    layer0_outputs(788) <= (inputs(149)) and (inputs(90));
    layer0_outputs(789) <= '1';
    layer0_outputs(790) <= (inputs(61)) or (inputs(101));
    layer0_outputs(791) <= not((inputs(193)) or (inputs(47)));
    layer0_outputs(792) <= not((inputs(175)) or (inputs(166)));
    layer0_outputs(793) <= (inputs(139)) and (inputs(75));
    layer0_outputs(794) <= (inputs(97)) and not (inputs(106));
    layer0_outputs(795) <= not((inputs(51)) xor (inputs(102)));
    layer0_outputs(796) <= not(inputs(152)) or (inputs(55));
    layer0_outputs(797) <= inputs(151);
    layer0_outputs(798) <= not(inputs(210));
    layer0_outputs(799) <= inputs(75);
    layer0_outputs(800) <= not(inputs(28));
    layer0_outputs(801) <= not((inputs(238)) xor (inputs(106)));
    layer0_outputs(802) <= not(inputs(162));
    layer0_outputs(803) <= not(inputs(18)) or (inputs(239));
    layer0_outputs(804) <= not(inputs(167)) or (inputs(116));
    layer0_outputs(805) <= not(inputs(88)) or (inputs(33));
    layer0_outputs(806) <= not(inputs(153));
    layer0_outputs(807) <= (inputs(56)) and (inputs(29));
    layer0_outputs(808) <= inputs(41);
    layer0_outputs(809) <= not(inputs(255)) or (inputs(247));
    layer0_outputs(810) <= inputs(167);
    layer0_outputs(811) <= (inputs(144)) xor (inputs(104));
    layer0_outputs(812) <= inputs(75);
    layer0_outputs(813) <= not((inputs(6)) and (inputs(81)));
    layer0_outputs(814) <= inputs(234);
    layer0_outputs(815) <= (inputs(198)) and not (inputs(82));
    layer0_outputs(816) <= (inputs(42)) xor (inputs(61));
    layer0_outputs(817) <= not((inputs(185)) or (inputs(65)));
    layer0_outputs(818) <= not((inputs(194)) xor (inputs(55)));
    layer0_outputs(819) <= not(inputs(67));
    layer0_outputs(820) <= (inputs(150)) and not (inputs(175));
    layer0_outputs(821) <= (inputs(186)) xor (inputs(207));
    layer0_outputs(822) <= (inputs(232)) or (inputs(249));
    layer0_outputs(823) <= not(inputs(7)) or (inputs(236));
    layer0_outputs(824) <= (inputs(40)) and not (inputs(61));
    layer0_outputs(825) <= not((inputs(111)) xor (inputs(138)));
    layer0_outputs(826) <= not(inputs(87));
    layer0_outputs(827) <= not((inputs(28)) or (inputs(66)));
    layer0_outputs(828) <= not(inputs(51)) or (inputs(165));
    layer0_outputs(829) <= inputs(4);
    layer0_outputs(830) <= not(inputs(122)) or (inputs(131));
    layer0_outputs(831) <= (inputs(2)) and (inputs(207));
    layer0_outputs(832) <= not(inputs(79)) or (inputs(48));
    layer0_outputs(833) <= not((inputs(74)) xor (inputs(0)));
    layer0_outputs(834) <= (inputs(141)) and not (inputs(253));
    layer0_outputs(835) <= (inputs(144)) and not (inputs(16));
    layer0_outputs(836) <= inputs(152);
    layer0_outputs(837) <= not(inputs(228));
    layer0_outputs(838) <= '1';
    layer0_outputs(839) <= not((inputs(98)) or (inputs(193)));
    layer0_outputs(840) <= (inputs(20)) and not (inputs(220));
    layer0_outputs(841) <= '1';
    layer0_outputs(842) <= not(inputs(80));
    layer0_outputs(843) <= not(inputs(200));
    layer0_outputs(844) <= (inputs(171)) xor (inputs(124));
    layer0_outputs(845) <= not(inputs(231));
    layer0_outputs(846) <= (inputs(89)) or (inputs(180));
    layer0_outputs(847) <= (inputs(158)) or (inputs(184));
    layer0_outputs(848) <= not((inputs(211)) and (inputs(123)));
    layer0_outputs(849) <= not((inputs(163)) xor (inputs(126)));
    layer0_outputs(850) <= not((inputs(241)) xor (inputs(191)));
    layer0_outputs(851) <= not((inputs(212)) or (inputs(189)));
    layer0_outputs(852) <= inputs(213);
    layer0_outputs(853) <= (inputs(114)) xor (inputs(252));
    layer0_outputs(854) <= inputs(181);
    layer0_outputs(855) <= inputs(54);
    layer0_outputs(856) <= not(inputs(155));
    layer0_outputs(857) <= inputs(51);
    layer0_outputs(858) <= not(inputs(204));
    layer0_outputs(859) <= inputs(181);
    layer0_outputs(860) <= not((inputs(7)) xor (inputs(26)));
    layer0_outputs(861) <= inputs(172);
    layer0_outputs(862) <= (inputs(49)) and not (inputs(178));
    layer0_outputs(863) <= not((inputs(183)) xor (inputs(45)));
    layer0_outputs(864) <= not(inputs(149)) or (inputs(18));
    layer0_outputs(865) <= (inputs(201)) xor (inputs(209));
    layer0_outputs(866) <= (inputs(158)) or (inputs(77));
    layer0_outputs(867) <= (inputs(109)) and not (inputs(98));
    layer0_outputs(868) <= (inputs(251)) or (inputs(15));
    layer0_outputs(869) <= (inputs(50)) and not (inputs(35));
    layer0_outputs(870) <= not((inputs(137)) and (inputs(19)));
    layer0_outputs(871) <= not(inputs(248));
    layer0_outputs(872) <= not((inputs(83)) xor (inputs(222)));
    layer0_outputs(873) <= not(inputs(38)) or (inputs(44));
    layer0_outputs(874) <= not(inputs(136));
    layer0_outputs(875) <= (inputs(154)) or (inputs(51));
    layer0_outputs(876) <= not(inputs(95));
    layer0_outputs(877) <= inputs(57);
    layer0_outputs(878) <= not((inputs(24)) or (inputs(107)));
    layer0_outputs(879) <= (inputs(229)) xor (inputs(190));
    layer0_outputs(880) <= (inputs(21)) and not (inputs(160));
    layer0_outputs(881) <= (inputs(115)) and not (inputs(186));
    layer0_outputs(882) <= not(inputs(23)) or (inputs(181));
    layer0_outputs(883) <= (inputs(144)) xor (inputs(15));
    layer0_outputs(884) <= not((inputs(159)) xor (inputs(195)));
    layer0_outputs(885) <= not(inputs(80));
    layer0_outputs(886) <= (inputs(87)) or (inputs(202));
    layer0_outputs(887) <= (inputs(192)) xor (inputs(244));
    layer0_outputs(888) <= (inputs(89)) and not (inputs(32));
    layer0_outputs(889) <= inputs(63);
    layer0_outputs(890) <= not(inputs(128));
    layer0_outputs(891) <= inputs(96);
    layer0_outputs(892) <= (inputs(211)) or (inputs(178));
    layer0_outputs(893) <= '0';
    layer0_outputs(894) <= inputs(178);
    layer0_outputs(895) <= not(inputs(170));
    layer0_outputs(896) <= (inputs(251)) or (inputs(98));
    layer0_outputs(897) <= inputs(162);
    layer0_outputs(898) <= not((inputs(186)) and (inputs(163)));
    layer0_outputs(899) <= (inputs(17)) xor (inputs(94));
    layer0_outputs(900) <= not((inputs(98)) or (inputs(172)));
    layer0_outputs(901) <= (inputs(177)) xor (inputs(82));
    layer0_outputs(902) <= (inputs(184)) and (inputs(141));
    layer0_outputs(903) <= not((inputs(113)) or (inputs(138)));
    layer0_outputs(904) <= (inputs(219)) or (inputs(20));
    layer0_outputs(905) <= '0';
    layer0_outputs(906) <= (inputs(243)) or (inputs(48));
    layer0_outputs(907) <= not(inputs(36)) or (inputs(206));
    layer0_outputs(908) <= not(inputs(120));
    layer0_outputs(909) <= not(inputs(227)) or (inputs(12));
    layer0_outputs(910) <= not(inputs(169)) or (inputs(68));
    layer0_outputs(911) <= not((inputs(109)) or (inputs(142)));
    layer0_outputs(912) <= not(inputs(243));
    layer0_outputs(913) <= not(inputs(218));
    layer0_outputs(914) <= (inputs(173)) and not (inputs(244));
    layer0_outputs(915) <= not(inputs(213));
    layer0_outputs(916) <= not(inputs(224));
    layer0_outputs(917) <= not(inputs(98));
    layer0_outputs(918) <= (inputs(62)) and not (inputs(134));
    layer0_outputs(919) <= (inputs(200)) and not (inputs(47));
    layer0_outputs(920) <= not(inputs(162)) or (inputs(49));
    layer0_outputs(921) <= (inputs(247)) and not (inputs(18));
    layer0_outputs(922) <= not(inputs(206));
    layer0_outputs(923) <= inputs(205);
    layer0_outputs(924) <= not(inputs(212));
    layer0_outputs(925) <= not(inputs(163)) or (inputs(36));
    layer0_outputs(926) <= (inputs(61)) and not (inputs(210));
    layer0_outputs(927) <= not(inputs(158));
    layer0_outputs(928) <= (inputs(61)) xor (inputs(75));
    layer0_outputs(929) <= not(inputs(228));
    layer0_outputs(930) <= not(inputs(6));
    layer0_outputs(931) <= (inputs(186)) and not (inputs(95));
    layer0_outputs(932) <= (inputs(174)) or (inputs(45));
    layer0_outputs(933) <= inputs(200);
    layer0_outputs(934) <= (inputs(61)) xor (inputs(28));
    layer0_outputs(935) <= inputs(64);
    layer0_outputs(936) <= not(inputs(233));
    layer0_outputs(937) <= not(inputs(143)) or (inputs(24));
    layer0_outputs(938) <= inputs(151);
    layer0_outputs(939) <= not(inputs(122)) or (inputs(95));
    layer0_outputs(940) <= (inputs(248)) xor (inputs(208));
    layer0_outputs(941) <= not(inputs(171));
    layer0_outputs(942) <= not((inputs(253)) or (inputs(233)));
    layer0_outputs(943) <= (inputs(15)) or (inputs(36));
    layer0_outputs(944) <= inputs(213);
    layer0_outputs(945) <= '0';
    layer0_outputs(946) <= (inputs(104)) xor (inputs(148));
    layer0_outputs(947) <= '0';
    layer0_outputs(948) <= (inputs(4)) xor (inputs(115));
    layer0_outputs(949) <= not(inputs(140)) or (inputs(241));
    layer0_outputs(950) <= inputs(116);
    layer0_outputs(951) <= inputs(167);
    layer0_outputs(952) <= (inputs(159)) and not (inputs(114));
    layer0_outputs(953) <= (inputs(158)) or (inputs(192));
    layer0_outputs(954) <= (inputs(35)) and not (inputs(253));
    layer0_outputs(955) <= not(inputs(218));
    layer0_outputs(956) <= not(inputs(213));
    layer0_outputs(957) <= (inputs(165)) xor (inputs(168));
    layer0_outputs(958) <= (inputs(122)) and not (inputs(65));
    layer0_outputs(959) <= inputs(56);
    layer0_outputs(960) <= not(inputs(183)) or (inputs(61));
    layer0_outputs(961) <= not(inputs(241)) or (inputs(251));
    layer0_outputs(962) <= not((inputs(255)) and (inputs(138)));
    layer0_outputs(963) <= (inputs(226)) and not (inputs(94));
    layer0_outputs(964) <= (inputs(76)) and not (inputs(254));
    layer0_outputs(965) <= not(inputs(8)) or (inputs(240));
    layer0_outputs(966) <= (inputs(202)) or (inputs(212));
    layer0_outputs(967) <= '0';
    layer0_outputs(968) <= inputs(123);
    layer0_outputs(969) <= '1';
    layer0_outputs(970) <= not((inputs(36)) xor (inputs(162)));
    layer0_outputs(971) <= not(inputs(167));
    layer0_outputs(972) <= (inputs(184)) and (inputs(48));
    layer0_outputs(973) <= not((inputs(11)) xor (inputs(224)));
    layer0_outputs(974) <= not((inputs(26)) xor (inputs(232)));
    layer0_outputs(975) <= inputs(93);
    layer0_outputs(976) <= not((inputs(20)) or (inputs(5)));
    layer0_outputs(977) <= not((inputs(45)) xor (inputs(59)));
    layer0_outputs(978) <= not(inputs(182));
    layer0_outputs(979) <= '1';
    layer0_outputs(980) <= not(inputs(132));
    layer0_outputs(981) <= inputs(168);
    layer0_outputs(982) <= not((inputs(118)) or (inputs(192)));
    layer0_outputs(983) <= not(inputs(139)) or (inputs(107));
    layer0_outputs(984) <= not((inputs(37)) or (inputs(98)));
    layer0_outputs(985) <= '0';
    layer0_outputs(986) <= not((inputs(101)) or (inputs(233)));
    layer0_outputs(987) <= not((inputs(33)) or (inputs(58)));
    layer0_outputs(988) <= not(inputs(18));
    layer0_outputs(989) <= (inputs(132)) xor (inputs(112));
    layer0_outputs(990) <= (inputs(180)) or (inputs(158));
    layer0_outputs(991) <= inputs(8);
    layer0_outputs(992) <= inputs(144);
    layer0_outputs(993) <= (inputs(213)) and not (inputs(39));
    layer0_outputs(994) <= not(inputs(25));
    layer0_outputs(995) <= '0';
    layer0_outputs(996) <= (inputs(118)) xor (inputs(166));
    layer0_outputs(997) <= inputs(232);
    layer0_outputs(998) <= (inputs(121)) xor (inputs(2));
    layer0_outputs(999) <= '1';
    layer0_outputs(1000) <= inputs(88);
    layer0_outputs(1001) <= (inputs(241)) and not (inputs(140));
    layer0_outputs(1002) <= not(inputs(62));
    layer0_outputs(1003) <= (inputs(195)) or (inputs(82));
    layer0_outputs(1004) <= (inputs(114)) or (inputs(133));
    layer0_outputs(1005) <= not((inputs(244)) or (inputs(190)));
    layer0_outputs(1006) <= '1';
    layer0_outputs(1007) <= inputs(218);
    layer0_outputs(1008) <= inputs(85);
    layer0_outputs(1009) <= not(inputs(77));
    layer0_outputs(1010) <= not(inputs(131));
    layer0_outputs(1011) <= (inputs(98)) or (inputs(132));
    layer0_outputs(1012) <= inputs(166);
    layer0_outputs(1013) <= inputs(56);
    layer0_outputs(1014) <= not(inputs(104)) or (inputs(114));
    layer0_outputs(1015) <= (inputs(117)) and (inputs(39));
    layer0_outputs(1016) <= (inputs(151)) or (inputs(2));
    layer0_outputs(1017) <= not(inputs(153));
    layer0_outputs(1018) <= (inputs(89)) xor (inputs(145));
    layer0_outputs(1019) <= not(inputs(229));
    layer0_outputs(1020) <= (inputs(229)) xor (inputs(161));
    layer0_outputs(1021) <= (inputs(152)) or (inputs(163));
    layer0_outputs(1022) <= inputs(169);
    layer0_outputs(1023) <= (inputs(255)) or (inputs(141));
    layer0_outputs(1024) <= (inputs(171)) and not (inputs(119));
    layer0_outputs(1025) <= not(inputs(149)) or (inputs(4));
    layer0_outputs(1026) <= (inputs(71)) or (inputs(157));
    layer0_outputs(1027) <= not((inputs(227)) or (inputs(233)));
    layer0_outputs(1028) <= not(inputs(244)) or (inputs(113));
    layer0_outputs(1029) <= not(inputs(89));
    layer0_outputs(1030) <= not(inputs(165));
    layer0_outputs(1031) <= not(inputs(229)) or (inputs(109));
    layer0_outputs(1032) <= inputs(69);
    layer0_outputs(1033) <= not(inputs(100)) or (inputs(225));
    layer0_outputs(1034) <= not((inputs(62)) or (inputs(223)));
    layer0_outputs(1035) <= inputs(173);
    layer0_outputs(1036) <= not(inputs(131));
    layer0_outputs(1037) <= not(inputs(39));
    layer0_outputs(1038) <= (inputs(166)) xor (inputs(163));
    layer0_outputs(1039) <= not(inputs(28));
    layer0_outputs(1040) <= (inputs(109)) xor (inputs(60));
    layer0_outputs(1041) <= (inputs(237)) and (inputs(143));
    layer0_outputs(1042) <= inputs(177);
    layer0_outputs(1043) <= not(inputs(56)) or (inputs(173));
    layer0_outputs(1044) <= not(inputs(180)) or (inputs(54));
    layer0_outputs(1045) <= not(inputs(0)) or (inputs(215));
    layer0_outputs(1046) <= (inputs(127)) xor (inputs(65));
    layer0_outputs(1047) <= (inputs(49)) xor (inputs(53));
    layer0_outputs(1048) <= not((inputs(144)) or (inputs(114)));
    layer0_outputs(1049) <= inputs(122);
    layer0_outputs(1050) <= inputs(236);
    layer0_outputs(1051) <= not((inputs(173)) and (inputs(111)));
    layer0_outputs(1052) <= inputs(122);
    layer0_outputs(1053) <= not(inputs(119));
    layer0_outputs(1054) <= (inputs(179)) and (inputs(148));
    layer0_outputs(1055) <= (inputs(13)) and (inputs(238));
    layer0_outputs(1056) <= not(inputs(181)) or (inputs(98));
    layer0_outputs(1057) <= not((inputs(166)) and (inputs(119)));
    layer0_outputs(1058) <= inputs(248);
    layer0_outputs(1059) <= (inputs(204)) and not (inputs(29));
    layer0_outputs(1060) <= (inputs(67)) and not (inputs(2));
    layer0_outputs(1061) <= (inputs(170)) or (inputs(133));
    layer0_outputs(1062) <= not(inputs(50)) or (inputs(231));
    layer0_outputs(1063) <= not((inputs(125)) xor (inputs(1)));
    layer0_outputs(1064) <= (inputs(154)) and not (inputs(169));
    layer0_outputs(1065) <= (inputs(106)) and not (inputs(227));
    layer0_outputs(1066) <= (inputs(58)) and not (inputs(227));
    layer0_outputs(1067) <= not(inputs(115));
    layer0_outputs(1068) <= not((inputs(155)) and (inputs(39)));
    layer0_outputs(1069) <= inputs(146);
    layer0_outputs(1070) <= not((inputs(31)) xor (inputs(137)));
    layer0_outputs(1071) <= not(inputs(45));
    layer0_outputs(1072) <= inputs(130);
    layer0_outputs(1073) <= not((inputs(163)) or (inputs(176)));
    layer0_outputs(1074) <= inputs(116);
    layer0_outputs(1075) <= not(inputs(66));
    layer0_outputs(1076) <= not(inputs(91)) or (inputs(123));
    layer0_outputs(1077) <= (inputs(35)) or (inputs(234));
    layer0_outputs(1078) <= not(inputs(8));
    layer0_outputs(1079) <= not(inputs(167));
    layer0_outputs(1080) <= not(inputs(126)) or (inputs(174));
    layer0_outputs(1081) <= not((inputs(57)) xor (inputs(72)));
    layer0_outputs(1082) <= not(inputs(42));
    layer0_outputs(1083) <= not((inputs(144)) and (inputs(28)));
    layer0_outputs(1084) <= not(inputs(36));
    layer0_outputs(1085) <= (inputs(62)) xor (inputs(79));
    layer0_outputs(1086) <= (inputs(70)) and not (inputs(59));
    layer0_outputs(1087) <= inputs(38);
    layer0_outputs(1088) <= inputs(56);
    layer0_outputs(1089) <= (inputs(46)) or (inputs(54));
    layer0_outputs(1090) <= not(inputs(67));
    layer0_outputs(1091) <= not(inputs(253)) or (inputs(32));
    layer0_outputs(1092) <= inputs(161);
    layer0_outputs(1093) <= inputs(217);
    layer0_outputs(1094) <= (inputs(98)) or (inputs(239));
    layer0_outputs(1095) <= inputs(250);
    layer0_outputs(1096) <= '0';
    layer0_outputs(1097) <= not(inputs(220));
    layer0_outputs(1098) <= '1';
    layer0_outputs(1099) <= not(inputs(230));
    layer0_outputs(1100) <= not(inputs(84));
    layer0_outputs(1101) <= (inputs(114)) or (inputs(167));
    layer0_outputs(1102) <= (inputs(8)) and not (inputs(3));
    layer0_outputs(1103) <= '0';
    layer0_outputs(1104) <= (inputs(120)) and not (inputs(33));
    layer0_outputs(1105) <= (inputs(200)) and not (inputs(73));
    layer0_outputs(1106) <= '1';
    layer0_outputs(1107) <= '0';
    layer0_outputs(1108) <= not(inputs(7));
    layer0_outputs(1109) <= (inputs(177)) xor (inputs(8));
    layer0_outputs(1110) <= not((inputs(237)) and (inputs(38)));
    layer0_outputs(1111) <= inputs(87);
    layer0_outputs(1112) <= not(inputs(82));
    layer0_outputs(1113) <= not(inputs(168)) or (inputs(90));
    layer0_outputs(1114) <= (inputs(118)) or (inputs(68));
    layer0_outputs(1115) <= not(inputs(34));
    layer0_outputs(1116) <= not((inputs(92)) and (inputs(108)));
    layer0_outputs(1117) <= '0';
    layer0_outputs(1118) <= not((inputs(148)) and (inputs(251)));
    layer0_outputs(1119) <= inputs(246);
    layer0_outputs(1120) <= '0';
    layer0_outputs(1121) <= not((inputs(228)) xor (inputs(62)));
    layer0_outputs(1122) <= not(inputs(57)) or (inputs(83));
    layer0_outputs(1123) <= (inputs(139)) xor (inputs(205));
    layer0_outputs(1124) <= not((inputs(201)) or (inputs(20)));
    layer0_outputs(1125) <= (inputs(192)) or (inputs(119));
    layer0_outputs(1126) <= (inputs(169)) or (inputs(120));
    layer0_outputs(1127) <= (inputs(102)) or (inputs(119));
    layer0_outputs(1128) <= (inputs(196)) and not (inputs(78));
    layer0_outputs(1129) <= (inputs(251)) xor (inputs(203));
    layer0_outputs(1130) <= not((inputs(247)) or (inputs(43)));
    layer0_outputs(1131) <= inputs(76);
    layer0_outputs(1132) <= inputs(1);
    layer0_outputs(1133) <= (inputs(83)) or (inputs(239));
    layer0_outputs(1134) <= (inputs(20)) xor (inputs(77));
    layer0_outputs(1135) <= (inputs(127)) or (inputs(213));
    layer0_outputs(1136) <= inputs(92);
    layer0_outputs(1137) <= (inputs(60)) xor (inputs(28));
    layer0_outputs(1138) <= (inputs(238)) or (inputs(210));
    layer0_outputs(1139) <= not(inputs(88)) or (inputs(239));
    layer0_outputs(1140) <= inputs(50);
    layer0_outputs(1141) <= '1';
    layer0_outputs(1142) <= (inputs(1)) or (inputs(187));
    layer0_outputs(1143) <= not((inputs(155)) or (inputs(196)));
    layer0_outputs(1144) <= not(inputs(198)) or (inputs(105));
    layer0_outputs(1145) <= not(inputs(60)) or (inputs(71));
    layer0_outputs(1146) <= not((inputs(127)) xor (inputs(203)));
    layer0_outputs(1147) <= not((inputs(62)) or (inputs(37)));
    layer0_outputs(1148) <= (inputs(239)) xor (inputs(87));
    layer0_outputs(1149) <= '0';
    layer0_outputs(1150) <= inputs(156);
    layer0_outputs(1151) <= not((inputs(73)) or (inputs(226)));
    layer0_outputs(1152) <= not(inputs(230));
    layer0_outputs(1153) <= (inputs(24)) and not (inputs(235));
    layer0_outputs(1154) <= inputs(201);
    layer0_outputs(1155) <= inputs(139);
    layer0_outputs(1156) <= not((inputs(132)) and (inputs(214)));
    layer0_outputs(1157) <= not((inputs(113)) xor (inputs(68)));
    layer0_outputs(1158) <= not((inputs(17)) xor (inputs(2)));
    layer0_outputs(1159) <= inputs(93);
    layer0_outputs(1160) <= not(inputs(152)) or (inputs(60));
    layer0_outputs(1161) <= (inputs(22)) xor (inputs(157));
    layer0_outputs(1162) <= inputs(27);
    layer0_outputs(1163) <= not((inputs(10)) and (inputs(216)));
    layer0_outputs(1164) <= (inputs(127)) or (inputs(183));
    layer0_outputs(1165) <= (inputs(86)) xor (inputs(117));
    layer0_outputs(1166) <= not((inputs(112)) xor (inputs(210)));
    layer0_outputs(1167) <= not(inputs(9));
    layer0_outputs(1168) <= not(inputs(200));
    layer0_outputs(1169) <= not((inputs(107)) and (inputs(139)));
    layer0_outputs(1170) <= not(inputs(160));
    layer0_outputs(1171) <= inputs(195);
    layer0_outputs(1172) <= not(inputs(39));
    layer0_outputs(1173) <= not((inputs(179)) xor (inputs(26)));
    layer0_outputs(1174) <= not((inputs(243)) or (inputs(210)));
    layer0_outputs(1175) <= not((inputs(222)) xor (inputs(21)));
    layer0_outputs(1176) <= (inputs(244)) xor (inputs(203));
    layer0_outputs(1177) <= (inputs(98)) xor (inputs(165));
    layer0_outputs(1178) <= not(inputs(62));
    layer0_outputs(1179) <= inputs(8);
    layer0_outputs(1180) <= inputs(52);
    layer0_outputs(1181) <= (inputs(215)) and (inputs(123));
    layer0_outputs(1182) <= not((inputs(170)) and (inputs(56)));
    layer0_outputs(1183) <= not((inputs(199)) and (inputs(202)));
    layer0_outputs(1184) <= inputs(62);
    layer0_outputs(1185) <= inputs(145);
    layer0_outputs(1186) <= (inputs(109)) or (inputs(207));
    layer0_outputs(1187) <= inputs(90);
    layer0_outputs(1188) <= (inputs(189)) and not (inputs(80));
    layer0_outputs(1189) <= not((inputs(216)) xor (inputs(11)));
    layer0_outputs(1190) <= (inputs(0)) and not (inputs(128));
    layer0_outputs(1191) <= (inputs(30)) and not (inputs(45));
    layer0_outputs(1192) <= not((inputs(57)) xor (inputs(113)));
    layer0_outputs(1193) <= not(inputs(224)) or (inputs(223));
    layer0_outputs(1194) <= inputs(214);
    layer0_outputs(1195) <= (inputs(181)) and not (inputs(39));
    layer0_outputs(1196) <= not((inputs(38)) xor (inputs(136)));
    layer0_outputs(1197) <= not((inputs(159)) and (inputs(240)));
    layer0_outputs(1198) <= (inputs(118)) and (inputs(120));
    layer0_outputs(1199) <= (inputs(140)) or (inputs(53));
    layer0_outputs(1200) <= not(inputs(38));
    layer0_outputs(1201) <= inputs(229);
    layer0_outputs(1202) <= (inputs(55)) and (inputs(205));
    layer0_outputs(1203) <= (inputs(55)) or (inputs(58));
    layer0_outputs(1204) <= (inputs(130)) and not (inputs(243));
    layer0_outputs(1205) <= not(inputs(22)) or (inputs(225));
    layer0_outputs(1206) <= inputs(230);
    layer0_outputs(1207) <= inputs(124);
    layer0_outputs(1208) <= (inputs(33)) or (inputs(166));
    layer0_outputs(1209) <= inputs(141);
    layer0_outputs(1210) <= inputs(206);
    layer0_outputs(1211) <= inputs(171);
    layer0_outputs(1212) <= not((inputs(168)) or (inputs(98)));
    layer0_outputs(1213) <= not(inputs(3));
    layer0_outputs(1214) <= not(inputs(49));
    layer0_outputs(1215) <= not(inputs(132)) or (inputs(251));
    layer0_outputs(1216) <= (inputs(161)) xor (inputs(23));
    layer0_outputs(1217) <= inputs(85);
    layer0_outputs(1218) <= inputs(69);
    layer0_outputs(1219) <= not((inputs(79)) or (inputs(162)));
    layer0_outputs(1220) <= not((inputs(27)) or (inputs(64)));
    layer0_outputs(1221) <= not((inputs(186)) or (inputs(78)));
    layer0_outputs(1222) <= (inputs(17)) xor (inputs(168));
    layer0_outputs(1223) <= not(inputs(145)) or (inputs(62));
    layer0_outputs(1224) <= (inputs(92)) and not (inputs(140));
    layer0_outputs(1225) <= not(inputs(54));
    layer0_outputs(1226) <= not((inputs(53)) or (inputs(200)));
    layer0_outputs(1227) <= not((inputs(210)) and (inputs(11)));
    layer0_outputs(1228) <= not((inputs(131)) xor (inputs(127)));
    layer0_outputs(1229) <= (inputs(77)) and not (inputs(172));
    layer0_outputs(1230) <= not(inputs(135));
    layer0_outputs(1231) <= (inputs(242)) xor (inputs(189));
    layer0_outputs(1232) <= (inputs(107)) and not (inputs(0));
    layer0_outputs(1233) <= not(inputs(133));
    layer0_outputs(1234) <= (inputs(191)) or (inputs(84));
    layer0_outputs(1235) <= inputs(246);
    layer0_outputs(1236) <= not(inputs(53)) or (inputs(93));
    layer0_outputs(1237) <= (inputs(146)) or (inputs(51));
    layer0_outputs(1238) <= not((inputs(253)) or (inputs(120)));
    layer0_outputs(1239) <= not((inputs(111)) xor (inputs(5)));
    layer0_outputs(1240) <= not((inputs(27)) or (inputs(21)));
    layer0_outputs(1241) <= inputs(180);
    layer0_outputs(1242) <= (inputs(51)) xor (inputs(71));
    layer0_outputs(1243) <= not(inputs(210));
    layer0_outputs(1244) <= (inputs(211)) or (inputs(37));
    layer0_outputs(1245) <= (inputs(12)) xor (inputs(2));
    layer0_outputs(1246) <= not((inputs(130)) or (inputs(253)));
    layer0_outputs(1247) <= not(inputs(8)) or (inputs(127));
    layer0_outputs(1248) <= (inputs(10)) and (inputs(27));
    layer0_outputs(1249) <= not((inputs(172)) or (inputs(100)));
    layer0_outputs(1250) <= not(inputs(215));
    layer0_outputs(1251) <= not(inputs(122)) or (inputs(241));
    layer0_outputs(1252) <= (inputs(164)) or (inputs(109));
    layer0_outputs(1253) <= inputs(198);
    layer0_outputs(1254) <= not((inputs(253)) and (inputs(166)));
    layer0_outputs(1255) <= not(inputs(86));
    layer0_outputs(1256) <= not((inputs(157)) or (inputs(77)));
    layer0_outputs(1257) <= not(inputs(152)) or (inputs(87));
    layer0_outputs(1258) <= inputs(72);
    layer0_outputs(1259) <= (inputs(121)) and not (inputs(194));
    layer0_outputs(1260) <= (inputs(245)) or (inputs(94));
    layer0_outputs(1261) <= (inputs(151)) xor (inputs(34));
    layer0_outputs(1262) <= (inputs(189)) and not (inputs(188));
    layer0_outputs(1263) <= (inputs(144)) and not (inputs(44));
    layer0_outputs(1264) <= not(inputs(137));
    layer0_outputs(1265) <= not(inputs(177));
    layer0_outputs(1266) <= not(inputs(180));
    layer0_outputs(1267) <= inputs(209);
    layer0_outputs(1268) <= (inputs(241)) or (inputs(202));
    layer0_outputs(1269) <= (inputs(134)) and (inputs(44));
    layer0_outputs(1270) <= not(inputs(220));
    layer0_outputs(1271) <= (inputs(90)) or (inputs(217));
    layer0_outputs(1272) <= (inputs(89)) and not (inputs(23));
    layer0_outputs(1273) <= not((inputs(209)) or (inputs(150)));
    layer0_outputs(1274) <= inputs(160);
    layer0_outputs(1275) <= not(inputs(214));
    layer0_outputs(1276) <= not(inputs(219));
    layer0_outputs(1277) <= not((inputs(19)) or (inputs(92)));
    layer0_outputs(1278) <= inputs(204);
    layer0_outputs(1279) <= not(inputs(237)) or (inputs(227));
    layer0_outputs(1280) <= not((inputs(64)) or (inputs(188)));
    layer0_outputs(1281) <= not((inputs(133)) and (inputs(122)));
    layer0_outputs(1282) <= not((inputs(176)) or (inputs(156)));
    layer0_outputs(1283) <= '0';
    layer0_outputs(1284) <= (inputs(250)) and not (inputs(0));
    layer0_outputs(1285) <= '0';
    layer0_outputs(1286) <= (inputs(80)) and not (inputs(223));
    layer0_outputs(1287) <= not(inputs(123));
    layer0_outputs(1288) <= inputs(110);
    layer0_outputs(1289) <= not(inputs(216));
    layer0_outputs(1290) <= not(inputs(152)) or (inputs(245));
    layer0_outputs(1291) <= inputs(116);
    layer0_outputs(1292) <= (inputs(220)) or (inputs(170));
    layer0_outputs(1293) <= (inputs(216)) xor (inputs(171));
    layer0_outputs(1294) <= inputs(94);
    layer0_outputs(1295) <= not(inputs(212));
    layer0_outputs(1296) <= inputs(91);
    layer0_outputs(1297) <= inputs(210);
    layer0_outputs(1298) <= (inputs(183)) xor (inputs(196));
    layer0_outputs(1299) <= not((inputs(125)) or (inputs(178)));
    layer0_outputs(1300) <= inputs(236);
    layer0_outputs(1301) <= not(inputs(233)) or (inputs(83));
    layer0_outputs(1302) <= '0';
    layer0_outputs(1303) <= (inputs(120)) and not (inputs(239));
    layer0_outputs(1304) <= not(inputs(218)) or (inputs(143));
    layer0_outputs(1305) <= (inputs(99)) or (inputs(29));
    layer0_outputs(1306) <= not(inputs(128));
    layer0_outputs(1307) <= not(inputs(191));
    layer0_outputs(1308) <= inputs(158);
    layer0_outputs(1309) <= not(inputs(99));
    layer0_outputs(1310) <= not((inputs(237)) or (inputs(199)));
    layer0_outputs(1311) <= inputs(106);
    layer0_outputs(1312) <= not((inputs(193)) and (inputs(222)));
    layer0_outputs(1313) <= not(inputs(237)) or (inputs(86));
    layer0_outputs(1314) <= not((inputs(36)) or (inputs(177)));
    layer0_outputs(1315) <= not((inputs(211)) and (inputs(38)));
    layer0_outputs(1316) <= (inputs(62)) xor (inputs(4));
    layer0_outputs(1317) <= (inputs(71)) and not (inputs(123));
    layer0_outputs(1318) <= inputs(119);
    layer0_outputs(1319) <= not(inputs(108)) or (inputs(17));
    layer0_outputs(1320) <= inputs(73);
    layer0_outputs(1321) <= not(inputs(41));
    layer0_outputs(1322) <= (inputs(244)) and not (inputs(219));
    layer0_outputs(1323) <= (inputs(183)) and not (inputs(130));
    layer0_outputs(1324) <= not(inputs(84)) or (inputs(72));
    layer0_outputs(1325) <= (inputs(176)) xor (inputs(138));
    layer0_outputs(1326) <= inputs(98);
    layer0_outputs(1327) <= inputs(37);
    layer0_outputs(1328) <= (inputs(250)) and not (inputs(49));
    layer0_outputs(1329) <= (inputs(159)) and (inputs(2));
    layer0_outputs(1330) <= (inputs(27)) or (inputs(50));
    layer0_outputs(1331) <= not(inputs(122)) or (inputs(42));
    layer0_outputs(1332) <= (inputs(206)) or (inputs(202));
    layer0_outputs(1333) <= not(inputs(105));
    layer0_outputs(1334) <= (inputs(41)) xor (inputs(67));
    layer0_outputs(1335) <= (inputs(138)) and not (inputs(166));
    layer0_outputs(1336) <= inputs(240);
    layer0_outputs(1337) <= (inputs(51)) xor (inputs(164));
    layer0_outputs(1338) <= (inputs(62)) and not (inputs(254));
    layer0_outputs(1339) <= not(inputs(79));
    layer0_outputs(1340) <= '1';
    layer0_outputs(1341) <= (inputs(17)) and not (inputs(232));
    layer0_outputs(1342) <= (inputs(165)) and not (inputs(111));
    layer0_outputs(1343) <= not(inputs(126));
    layer0_outputs(1344) <= not((inputs(253)) and (inputs(144)));
    layer0_outputs(1345) <= not(inputs(122)) or (inputs(27));
    layer0_outputs(1346) <= (inputs(107)) or (inputs(48));
    layer0_outputs(1347) <= (inputs(172)) xor (inputs(190));
    layer0_outputs(1348) <= not(inputs(132)) or (inputs(57));
    layer0_outputs(1349) <= not(inputs(84));
    layer0_outputs(1350) <= not(inputs(227));
    layer0_outputs(1351) <= not((inputs(160)) or (inputs(66)));
    layer0_outputs(1352) <= (inputs(207)) xor (inputs(250));
    layer0_outputs(1353) <= inputs(102);
    layer0_outputs(1354) <= '1';
    layer0_outputs(1355) <= (inputs(64)) and (inputs(5));
    layer0_outputs(1356) <= inputs(109);
    layer0_outputs(1357) <= not(inputs(234)) or (inputs(6));
    layer0_outputs(1358) <= (inputs(207)) and (inputs(109));
    layer0_outputs(1359) <= not(inputs(146)) or (inputs(62));
    layer0_outputs(1360) <= (inputs(124)) or (inputs(8));
    layer0_outputs(1361) <= inputs(126);
    layer0_outputs(1362) <= (inputs(213)) or (inputs(208));
    layer0_outputs(1363) <= not(inputs(22));
    layer0_outputs(1364) <= (inputs(97)) or (inputs(227));
    layer0_outputs(1365) <= not((inputs(174)) and (inputs(204)));
    layer0_outputs(1366) <= not(inputs(58)) or (inputs(117));
    layer0_outputs(1367) <= not((inputs(111)) xor (inputs(239)));
    layer0_outputs(1368) <= not(inputs(148));
    layer0_outputs(1369) <= (inputs(245)) and (inputs(202));
    layer0_outputs(1370) <= not((inputs(162)) xor (inputs(233)));
    layer0_outputs(1371) <= not(inputs(142));
    layer0_outputs(1372) <= inputs(59);
    layer0_outputs(1373) <= not((inputs(230)) and (inputs(165)));
    layer0_outputs(1374) <= not(inputs(174)) or (inputs(132));
    layer0_outputs(1375) <= not(inputs(106));
    layer0_outputs(1376) <= not((inputs(104)) or (inputs(31)));
    layer0_outputs(1377) <= inputs(126);
    layer0_outputs(1378) <= (inputs(29)) or (inputs(120));
    layer0_outputs(1379) <= (inputs(85)) and not (inputs(74));
    layer0_outputs(1380) <= not((inputs(97)) and (inputs(187)));
    layer0_outputs(1381) <= '1';
    layer0_outputs(1382) <= not(inputs(172));
    layer0_outputs(1383) <= not(inputs(6));
    layer0_outputs(1384) <= (inputs(74)) and (inputs(100));
    layer0_outputs(1385) <= (inputs(231)) and (inputs(226));
    layer0_outputs(1386) <= not(inputs(251));
    layer0_outputs(1387) <= '0';
    layer0_outputs(1388) <= not(inputs(26)) or (inputs(252));
    layer0_outputs(1389) <= not(inputs(88));
    layer0_outputs(1390) <= (inputs(130)) or (inputs(218));
    layer0_outputs(1391) <= (inputs(100)) and not (inputs(126));
    layer0_outputs(1392) <= '1';
    layer0_outputs(1393) <= inputs(43);
    layer0_outputs(1394) <= not(inputs(20)) or (inputs(114));
    layer0_outputs(1395) <= inputs(126);
    layer0_outputs(1396) <= '1';
    layer0_outputs(1397) <= not(inputs(129)) or (inputs(66));
    layer0_outputs(1398) <= not(inputs(120)) or (inputs(12));
    layer0_outputs(1399) <= inputs(209);
    layer0_outputs(1400) <= not(inputs(193));
    layer0_outputs(1401) <= not((inputs(15)) xor (inputs(147)));
    layer0_outputs(1402) <= (inputs(182)) and not (inputs(209));
    layer0_outputs(1403) <= not(inputs(70));
    layer0_outputs(1404) <= (inputs(240)) xor (inputs(139));
    layer0_outputs(1405) <= not((inputs(20)) xor (inputs(81)));
    layer0_outputs(1406) <= not((inputs(28)) or (inputs(160)));
    layer0_outputs(1407) <= (inputs(175)) and not (inputs(255));
    layer0_outputs(1408) <= (inputs(32)) and (inputs(99));
    layer0_outputs(1409) <= not((inputs(116)) or (inputs(61)));
    layer0_outputs(1410) <= inputs(120);
    layer0_outputs(1411) <= inputs(239);
    layer0_outputs(1412) <= inputs(71);
    layer0_outputs(1413) <= (inputs(184)) and (inputs(9));
    layer0_outputs(1414) <= inputs(28);
    layer0_outputs(1415) <= not((inputs(30)) xor (inputs(76)));
    layer0_outputs(1416) <= '0';
    layer0_outputs(1417) <= not((inputs(186)) or (inputs(194)));
    layer0_outputs(1418) <= (inputs(123)) xor (inputs(68));
    layer0_outputs(1419) <= (inputs(13)) or (inputs(176));
    layer0_outputs(1420) <= (inputs(121)) and not (inputs(168));
    layer0_outputs(1421) <= not(inputs(9));
    layer0_outputs(1422) <= (inputs(26)) and not (inputs(201));
    layer0_outputs(1423) <= inputs(113);
    layer0_outputs(1424) <= not((inputs(128)) xor (inputs(231)));
    layer0_outputs(1425) <= inputs(201);
    layer0_outputs(1426) <= not(inputs(94));
    layer0_outputs(1427) <= not(inputs(8)) or (inputs(241));
    layer0_outputs(1428) <= (inputs(13)) or (inputs(92));
    layer0_outputs(1429) <= (inputs(222)) or (inputs(203));
    layer0_outputs(1430) <= not(inputs(134)) or (inputs(43));
    layer0_outputs(1431) <= not((inputs(148)) xor (inputs(151)));
    layer0_outputs(1432) <= not(inputs(205)) or (inputs(198));
    layer0_outputs(1433) <= not((inputs(167)) and (inputs(110)));
    layer0_outputs(1434) <= (inputs(69)) or (inputs(130));
    layer0_outputs(1435) <= (inputs(203)) and (inputs(95));
    layer0_outputs(1436) <= not(inputs(228)) or (inputs(132));
    layer0_outputs(1437) <= not((inputs(205)) or (inputs(188)));
    layer0_outputs(1438) <= inputs(152);
    layer0_outputs(1439) <= not((inputs(18)) xor (inputs(26)));
    layer0_outputs(1440) <= (inputs(7)) or (inputs(109));
    layer0_outputs(1441) <= (inputs(231)) and (inputs(181));
    layer0_outputs(1442) <= not(inputs(124));
    layer0_outputs(1443) <= not(inputs(157));
    layer0_outputs(1444) <= inputs(134);
    layer0_outputs(1445) <= (inputs(132)) or (inputs(80));
    layer0_outputs(1446) <= inputs(144);
    layer0_outputs(1447) <= not((inputs(222)) or (inputs(201)));
    layer0_outputs(1448) <= not(inputs(157)) or (inputs(65));
    layer0_outputs(1449) <= inputs(202);
    layer0_outputs(1450) <= (inputs(45)) xor (inputs(19));
    layer0_outputs(1451) <= (inputs(64)) xor (inputs(126));
    layer0_outputs(1452) <= inputs(3);
    layer0_outputs(1453) <= (inputs(48)) or (inputs(80));
    layer0_outputs(1454) <= (inputs(47)) and not (inputs(255));
    layer0_outputs(1455) <= (inputs(101)) or (inputs(143));
    layer0_outputs(1456) <= (inputs(150)) or (inputs(164));
    layer0_outputs(1457) <= inputs(214);
    layer0_outputs(1458) <= not(inputs(199)) or (inputs(97));
    layer0_outputs(1459) <= inputs(226);
    layer0_outputs(1460) <= not(inputs(40));
    layer0_outputs(1461) <= '1';
    layer0_outputs(1462) <= not(inputs(137));
    layer0_outputs(1463) <= (inputs(183)) or (inputs(86));
    layer0_outputs(1464) <= not(inputs(99)) or (inputs(30));
    layer0_outputs(1465) <= inputs(87);
    layer0_outputs(1466) <= (inputs(226)) and not (inputs(124));
    layer0_outputs(1467) <= not((inputs(4)) xor (inputs(60)));
    layer0_outputs(1468) <= not(inputs(165));
    layer0_outputs(1469) <= (inputs(109)) and not (inputs(249));
    layer0_outputs(1470) <= not(inputs(41));
    layer0_outputs(1471) <= not(inputs(128));
    layer0_outputs(1472) <= not(inputs(213)) or (inputs(143));
    layer0_outputs(1473) <= (inputs(31)) and not (inputs(129));
    layer0_outputs(1474) <= not(inputs(120));
    layer0_outputs(1475) <= not(inputs(55));
    layer0_outputs(1476) <= (inputs(188)) or (inputs(204));
    layer0_outputs(1477) <= inputs(96);
    layer0_outputs(1478) <= (inputs(54)) and not (inputs(74));
    layer0_outputs(1479) <= not((inputs(186)) and (inputs(179)));
    layer0_outputs(1480) <= inputs(98);
    layer0_outputs(1481) <= (inputs(165)) or (inputs(161));
    layer0_outputs(1482) <= not(inputs(120));
    layer0_outputs(1483) <= not((inputs(2)) and (inputs(5)));
    layer0_outputs(1484) <= (inputs(170)) or (inputs(63));
    layer0_outputs(1485) <= (inputs(99)) xor (inputs(54));
    layer0_outputs(1486) <= not(inputs(206));
    layer0_outputs(1487) <= not((inputs(172)) or (inputs(179)));
    layer0_outputs(1488) <= not(inputs(230));
    layer0_outputs(1489) <= not(inputs(59)) or (inputs(250));
    layer0_outputs(1490) <= (inputs(106)) or (inputs(12));
    layer0_outputs(1491) <= not(inputs(26));
    layer0_outputs(1492) <= '1';
    layer0_outputs(1493) <= inputs(148);
    layer0_outputs(1494) <= not(inputs(188)) or (inputs(223));
    layer0_outputs(1495) <= not(inputs(240));
    layer0_outputs(1496) <= not(inputs(63));
    layer0_outputs(1497) <= (inputs(236)) and not (inputs(228));
    layer0_outputs(1498) <= not((inputs(182)) or (inputs(36)));
    layer0_outputs(1499) <= (inputs(155)) and not (inputs(141));
    layer0_outputs(1500) <= not((inputs(82)) or (inputs(72)));
    layer0_outputs(1501) <= not(inputs(244)) or (inputs(238));
    layer0_outputs(1502) <= (inputs(22)) or (inputs(185));
    layer0_outputs(1503) <= (inputs(228)) and not (inputs(101));
    layer0_outputs(1504) <= (inputs(180)) and not (inputs(79));
    layer0_outputs(1505) <= not((inputs(180)) or (inputs(49)));
    layer0_outputs(1506) <= not((inputs(50)) and (inputs(47)));
    layer0_outputs(1507) <= not(inputs(143)) or (inputs(171));
    layer0_outputs(1508) <= '0';
    layer0_outputs(1509) <= (inputs(249)) and (inputs(59));
    layer0_outputs(1510) <= (inputs(69)) and not (inputs(178));
    layer0_outputs(1511) <= (inputs(58)) or (inputs(118));
    layer0_outputs(1512) <= not((inputs(2)) xor (inputs(237)));
    layer0_outputs(1513) <= not((inputs(64)) and (inputs(234)));
    layer0_outputs(1514) <= not(inputs(102)) or (inputs(17));
    layer0_outputs(1515) <= not(inputs(61));
    layer0_outputs(1516) <= inputs(37);
    layer0_outputs(1517) <= inputs(135);
    layer0_outputs(1518) <= (inputs(160)) xor (inputs(180));
    layer0_outputs(1519) <= inputs(216);
    layer0_outputs(1520) <= inputs(151);
    layer0_outputs(1521) <= not((inputs(1)) xor (inputs(59)));
    layer0_outputs(1522) <= (inputs(253)) and (inputs(11));
    layer0_outputs(1523) <= (inputs(31)) and (inputs(216));
    layer0_outputs(1524) <= (inputs(87)) or (inputs(89));
    layer0_outputs(1525) <= not((inputs(147)) or (inputs(162)));
    layer0_outputs(1526) <= inputs(59);
    layer0_outputs(1527) <= (inputs(116)) xor (inputs(169));
    layer0_outputs(1528) <= not(inputs(246)) or (inputs(138));
    layer0_outputs(1529) <= inputs(99);
    layer0_outputs(1530) <= not((inputs(21)) and (inputs(155)));
    layer0_outputs(1531) <= inputs(230);
    layer0_outputs(1532) <= (inputs(54)) or (inputs(29));
    layer0_outputs(1533) <= (inputs(182)) and not (inputs(252));
    layer0_outputs(1534) <= not((inputs(55)) xor (inputs(9)));
    layer0_outputs(1535) <= not((inputs(184)) xor (inputs(239)));
    layer0_outputs(1536) <= inputs(165);
    layer0_outputs(1537) <= (inputs(210)) or (inputs(80));
    layer0_outputs(1538) <= not(inputs(38));
    layer0_outputs(1539) <= (inputs(234)) or (inputs(1));
    layer0_outputs(1540) <= (inputs(25)) or (inputs(34));
    layer0_outputs(1541) <= not((inputs(161)) or (inputs(207)));
    layer0_outputs(1542) <= inputs(9);
    layer0_outputs(1543) <= not(inputs(134)) or (inputs(133));
    layer0_outputs(1544) <= not(inputs(107)) or (inputs(25));
    layer0_outputs(1545) <= not(inputs(148)) or (inputs(93));
    layer0_outputs(1546) <= not(inputs(166));
    layer0_outputs(1547) <= '1';
    layer0_outputs(1548) <= inputs(151);
    layer0_outputs(1549) <= '1';
    layer0_outputs(1550) <= not(inputs(203));
    layer0_outputs(1551) <= (inputs(12)) or (inputs(128));
    layer0_outputs(1552) <= inputs(179);
    layer0_outputs(1553) <= not((inputs(198)) and (inputs(186)));
    layer0_outputs(1554) <= not(inputs(68));
    layer0_outputs(1555) <= inputs(43);
    layer0_outputs(1556) <= not(inputs(81));
    layer0_outputs(1557) <= inputs(213);
    layer0_outputs(1558) <= inputs(220);
    layer0_outputs(1559) <= inputs(239);
    layer0_outputs(1560) <= not((inputs(17)) or (inputs(43)));
    layer0_outputs(1561) <= not((inputs(83)) or (inputs(52)));
    layer0_outputs(1562) <= not(inputs(100));
    layer0_outputs(1563) <= not((inputs(241)) xor (inputs(119)));
    layer0_outputs(1564) <= not(inputs(32)) or (inputs(121));
    layer0_outputs(1565) <= not(inputs(157));
    layer0_outputs(1566) <= (inputs(115)) or (inputs(157));
    layer0_outputs(1567) <= not(inputs(102)) or (inputs(223));
    layer0_outputs(1568) <= not(inputs(74));
    layer0_outputs(1569) <= not(inputs(254));
    layer0_outputs(1570) <= not(inputs(233));
    layer0_outputs(1571) <= not((inputs(233)) and (inputs(26)));
    layer0_outputs(1572) <= inputs(200);
    layer0_outputs(1573) <= (inputs(238)) and not (inputs(3));
    layer0_outputs(1574) <= inputs(23);
    layer0_outputs(1575) <= (inputs(14)) and not (inputs(26));
    layer0_outputs(1576) <= not(inputs(107)) or (inputs(192));
    layer0_outputs(1577) <= inputs(26);
    layer0_outputs(1578) <= (inputs(190)) or (inputs(243));
    layer0_outputs(1579) <= not((inputs(1)) or (inputs(54)));
    layer0_outputs(1580) <= not((inputs(197)) and (inputs(90)));
    layer0_outputs(1581) <= not((inputs(219)) xor (inputs(52)));
    layer0_outputs(1582) <= inputs(25);
    layer0_outputs(1583) <= inputs(7);
    layer0_outputs(1584) <= not((inputs(86)) xor (inputs(164)));
    layer0_outputs(1585) <= inputs(92);
    layer0_outputs(1586) <= (inputs(221)) or (inputs(228));
    layer0_outputs(1587) <= not(inputs(135));
    layer0_outputs(1588) <= inputs(120);
    layer0_outputs(1589) <= (inputs(203)) or (inputs(118));
    layer0_outputs(1590) <= '0';
    layer0_outputs(1591) <= inputs(150);
    layer0_outputs(1592) <= not((inputs(228)) or (inputs(233)));
    layer0_outputs(1593) <= (inputs(7)) and not (inputs(224));
    layer0_outputs(1594) <= not(inputs(18));
    layer0_outputs(1595) <= '1';
    layer0_outputs(1596) <= inputs(252);
    layer0_outputs(1597) <= not((inputs(181)) or (inputs(180)));
    layer0_outputs(1598) <= not((inputs(165)) or (inputs(142)));
    layer0_outputs(1599) <= inputs(103);
    layer0_outputs(1600) <= '1';
    layer0_outputs(1601) <= '0';
    layer0_outputs(1602) <= inputs(200);
    layer0_outputs(1603) <= (inputs(203)) or (inputs(115));
    layer0_outputs(1604) <= not((inputs(189)) xor (inputs(143)));
    layer0_outputs(1605) <= not(inputs(165)) or (inputs(140));
    layer0_outputs(1606) <= inputs(232);
    layer0_outputs(1607) <= not((inputs(198)) xor (inputs(58)));
    layer0_outputs(1608) <= inputs(126);
    layer0_outputs(1609) <= (inputs(209)) xor (inputs(32));
    layer0_outputs(1610) <= (inputs(171)) xor (inputs(253));
    layer0_outputs(1611) <= (inputs(205)) xor (inputs(186));
    layer0_outputs(1612) <= inputs(121);
    layer0_outputs(1613) <= not(inputs(76)) or (inputs(156));
    layer0_outputs(1614) <= (inputs(225)) or (inputs(62));
    layer0_outputs(1615) <= '1';
    layer0_outputs(1616) <= inputs(70);
    layer0_outputs(1617) <= (inputs(112)) and not (inputs(218));
    layer0_outputs(1618) <= not(inputs(38));
    layer0_outputs(1619) <= (inputs(233)) or (inputs(114));
    layer0_outputs(1620) <= (inputs(211)) and not (inputs(28));
    layer0_outputs(1621) <= not(inputs(198)) or (inputs(94));
    layer0_outputs(1622) <= inputs(131);
    layer0_outputs(1623) <= not(inputs(219));
    layer0_outputs(1624) <= not((inputs(245)) or (inputs(237)));
    layer0_outputs(1625) <= not((inputs(149)) or (inputs(70)));
    layer0_outputs(1626) <= inputs(190);
    layer0_outputs(1627) <= inputs(181);
    layer0_outputs(1628) <= (inputs(227)) or (inputs(48));
    layer0_outputs(1629) <= (inputs(116)) xor (inputs(118));
    layer0_outputs(1630) <= not(inputs(93)) or (inputs(216));
    layer0_outputs(1631) <= inputs(133);
    layer0_outputs(1632) <= (inputs(44)) or (inputs(129));
    layer0_outputs(1633) <= not(inputs(118)) or (inputs(175));
    layer0_outputs(1634) <= not(inputs(102)) or (inputs(218));
    layer0_outputs(1635) <= inputs(88);
    layer0_outputs(1636) <= not(inputs(102)) or (inputs(74));
    layer0_outputs(1637) <= (inputs(6)) or (inputs(129));
    layer0_outputs(1638) <= (inputs(214)) or (inputs(230));
    layer0_outputs(1639) <= (inputs(216)) and not (inputs(138));
    layer0_outputs(1640) <= (inputs(205)) or (inputs(254));
    layer0_outputs(1641) <= (inputs(180)) and (inputs(66));
    layer0_outputs(1642) <= not(inputs(164));
    layer0_outputs(1643) <= (inputs(52)) and not (inputs(202));
    layer0_outputs(1644) <= not(inputs(137));
    layer0_outputs(1645) <= (inputs(50)) or (inputs(249));
    layer0_outputs(1646) <= (inputs(233)) and not (inputs(79));
    layer0_outputs(1647) <= (inputs(184)) xor (inputs(146));
    layer0_outputs(1648) <= inputs(24);
    layer0_outputs(1649) <= not(inputs(132));
    layer0_outputs(1650) <= (inputs(78)) and not (inputs(150));
    layer0_outputs(1651) <= not((inputs(191)) or (inputs(207)));
    layer0_outputs(1652) <= inputs(201);
    layer0_outputs(1653) <= (inputs(108)) and not (inputs(205));
    layer0_outputs(1654) <= (inputs(247)) and not (inputs(113));
    layer0_outputs(1655) <= not(inputs(164));
    layer0_outputs(1656) <= not((inputs(228)) or (inputs(93)));
    layer0_outputs(1657) <= not(inputs(69)) or (inputs(93));
    layer0_outputs(1658) <= not((inputs(169)) xor (inputs(150)));
    layer0_outputs(1659) <= inputs(18);
    layer0_outputs(1660) <= (inputs(53)) and not (inputs(15));
    layer0_outputs(1661) <= (inputs(164)) or (inputs(62));
    layer0_outputs(1662) <= inputs(91);
    layer0_outputs(1663) <= not((inputs(177)) or (inputs(139)));
    layer0_outputs(1664) <= (inputs(1)) xor (inputs(21));
    layer0_outputs(1665) <= (inputs(77)) xor (inputs(228));
    layer0_outputs(1666) <= (inputs(148)) and (inputs(197));
    layer0_outputs(1667) <= not(inputs(251));
    layer0_outputs(1668) <= not(inputs(70));
    layer0_outputs(1669) <= not((inputs(191)) or (inputs(25)));
    layer0_outputs(1670) <= '0';
    layer0_outputs(1671) <= not((inputs(76)) or (inputs(208)));
    layer0_outputs(1672) <= not(inputs(186)) or (inputs(82));
    layer0_outputs(1673) <= (inputs(157)) and not (inputs(66));
    layer0_outputs(1674) <= (inputs(200)) and not (inputs(222));
    layer0_outputs(1675) <= not(inputs(101)) or (inputs(49));
    layer0_outputs(1676) <= (inputs(133)) or (inputs(66));
    layer0_outputs(1677) <= inputs(78);
    layer0_outputs(1678) <= not(inputs(141));
    layer0_outputs(1679) <= not((inputs(58)) xor (inputs(89)));
    layer0_outputs(1680) <= (inputs(69)) xor (inputs(173));
    layer0_outputs(1681) <= inputs(246);
    layer0_outputs(1682) <= not(inputs(193)) or (inputs(1));
    layer0_outputs(1683) <= not(inputs(70));
    layer0_outputs(1684) <= (inputs(108)) or (inputs(23));
    layer0_outputs(1685) <= (inputs(96)) xor (inputs(10));
    layer0_outputs(1686) <= not(inputs(33));
    layer0_outputs(1687) <= inputs(56);
    layer0_outputs(1688) <= (inputs(80)) or (inputs(196));
    layer0_outputs(1689) <= (inputs(169)) xor (inputs(110));
    layer0_outputs(1690) <= not(inputs(248)) or (inputs(2));
    layer0_outputs(1691) <= not(inputs(134)) or (inputs(121));
    layer0_outputs(1692) <= (inputs(230)) and not (inputs(50));
    layer0_outputs(1693) <= (inputs(108)) and not (inputs(226));
    layer0_outputs(1694) <= (inputs(77)) and not (inputs(241));
    layer0_outputs(1695) <= not(inputs(16));
    layer0_outputs(1696) <= not(inputs(172));
    layer0_outputs(1697) <= inputs(154);
    layer0_outputs(1698) <= not((inputs(208)) and (inputs(234)));
    layer0_outputs(1699) <= not((inputs(97)) or (inputs(68)));
    layer0_outputs(1700) <= inputs(157);
    layer0_outputs(1701) <= (inputs(192)) or (inputs(155));
    layer0_outputs(1702) <= not((inputs(85)) xor (inputs(170)));
    layer0_outputs(1703) <= not(inputs(151)) or (inputs(132));
    layer0_outputs(1704) <= (inputs(191)) and not (inputs(31));
    layer0_outputs(1705) <= (inputs(110)) and not (inputs(223));
    layer0_outputs(1706) <= not(inputs(150)) or (inputs(112));
    layer0_outputs(1707) <= (inputs(196)) xor (inputs(104));
    layer0_outputs(1708) <= not(inputs(11)) or (inputs(223));
    layer0_outputs(1709) <= not(inputs(26)) or (inputs(182));
    layer0_outputs(1710) <= inputs(161);
    layer0_outputs(1711) <= (inputs(7)) and not (inputs(163));
    layer0_outputs(1712) <= inputs(142);
    layer0_outputs(1713) <= inputs(115);
    layer0_outputs(1714) <= not((inputs(239)) or (inputs(239)));
    layer0_outputs(1715) <= not((inputs(39)) or (inputs(29)));
    layer0_outputs(1716) <= not((inputs(251)) or (inputs(200)));
    layer0_outputs(1717) <= inputs(192);
    layer0_outputs(1718) <= not(inputs(20)) or (inputs(128));
    layer0_outputs(1719) <= inputs(41);
    layer0_outputs(1720) <= not(inputs(92));
    layer0_outputs(1721) <= inputs(237);
    layer0_outputs(1722) <= not(inputs(219));
    layer0_outputs(1723) <= '1';
    layer0_outputs(1724) <= (inputs(33)) xor (inputs(138));
    layer0_outputs(1725) <= '0';
    layer0_outputs(1726) <= (inputs(27)) and not (inputs(210));
    layer0_outputs(1727) <= not(inputs(28)) or (inputs(223));
    layer0_outputs(1728) <= inputs(152);
    layer0_outputs(1729) <= not(inputs(53)) or (inputs(85));
    layer0_outputs(1730) <= (inputs(20)) or (inputs(79));
    layer0_outputs(1731) <= not(inputs(78));
    layer0_outputs(1732) <= (inputs(14)) xor (inputs(72));
    layer0_outputs(1733) <= (inputs(70)) or (inputs(61));
    layer0_outputs(1734) <= (inputs(199)) or (inputs(65));
    layer0_outputs(1735) <= not(inputs(144));
    layer0_outputs(1736) <= not(inputs(4));
    layer0_outputs(1737) <= (inputs(108)) and not (inputs(207));
    layer0_outputs(1738) <= not((inputs(152)) and (inputs(203)));
    layer0_outputs(1739) <= not(inputs(142)) or (inputs(229));
    layer0_outputs(1740) <= not(inputs(111));
    layer0_outputs(1741) <= (inputs(40)) and not (inputs(178));
    layer0_outputs(1742) <= not((inputs(96)) xor (inputs(68)));
    layer0_outputs(1743) <= not(inputs(248)) or (inputs(73));
    layer0_outputs(1744) <= not((inputs(50)) or (inputs(9)));
    layer0_outputs(1745) <= not(inputs(61)) or (inputs(27));
    layer0_outputs(1746) <= '0';
    layer0_outputs(1747) <= not((inputs(115)) xor (inputs(178)));
    layer0_outputs(1748) <= not(inputs(191)) or (inputs(251));
    layer0_outputs(1749) <= (inputs(191)) or (inputs(31));
    layer0_outputs(1750) <= not(inputs(54)) or (inputs(13));
    layer0_outputs(1751) <= (inputs(71)) and not (inputs(220));
    layer0_outputs(1752) <= not(inputs(231)) or (inputs(53));
    layer0_outputs(1753) <= not((inputs(153)) or (inputs(248)));
    layer0_outputs(1754) <= (inputs(92)) xor (inputs(129));
    layer0_outputs(1755) <= not((inputs(152)) xor (inputs(121)));
    layer0_outputs(1756) <= inputs(147);
    layer0_outputs(1757) <= not(inputs(40));
    layer0_outputs(1758) <= (inputs(218)) and (inputs(94));
    layer0_outputs(1759) <= inputs(23);
    layer0_outputs(1760) <= inputs(203);
    layer0_outputs(1761) <= not(inputs(229));
    layer0_outputs(1762) <= not((inputs(89)) xor (inputs(38)));
    layer0_outputs(1763) <= not(inputs(231));
    layer0_outputs(1764) <= not(inputs(226)) or (inputs(220));
    layer0_outputs(1765) <= (inputs(70)) or (inputs(147));
    layer0_outputs(1766) <= not(inputs(163)) or (inputs(214));
    layer0_outputs(1767) <= not(inputs(87)) or (inputs(24));
    layer0_outputs(1768) <= (inputs(94)) or (inputs(8));
    layer0_outputs(1769) <= not(inputs(147)) or (inputs(239));
    layer0_outputs(1770) <= not(inputs(30));
    layer0_outputs(1771) <= inputs(180);
    layer0_outputs(1772) <= (inputs(149)) or (inputs(198));
    layer0_outputs(1773) <= inputs(118);
    layer0_outputs(1774) <= not((inputs(192)) or (inputs(234)));
    layer0_outputs(1775) <= (inputs(117)) and not (inputs(65));
    layer0_outputs(1776) <= not((inputs(3)) xor (inputs(33)));
    layer0_outputs(1777) <= not(inputs(113)) or (inputs(233));
    layer0_outputs(1778) <= not(inputs(16));
    layer0_outputs(1779) <= (inputs(183)) and not (inputs(130));
    layer0_outputs(1780) <= not((inputs(213)) or (inputs(127)));
    layer0_outputs(1781) <= not((inputs(151)) and (inputs(231)));
    layer0_outputs(1782) <= (inputs(8)) and (inputs(73));
    layer0_outputs(1783) <= not((inputs(187)) or (inputs(172)));
    layer0_outputs(1784) <= not(inputs(113)) or (inputs(134));
    layer0_outputs(1785) <= not((inputs(0)) or (inputs(8)));
    layer0_outputs(1786) <= not(inputs(80)) or (inputs(144));
    layer0_outputs(1787) <= not(inputs(60)) or (inputs(32));
    layer0_outputs(1788) <= not(inputs(56));
    layer0_outputs(1789) <= not(inputs(199));
    layer0_outputs(1790) <= (inputs(138)) or (inputs(91));
    layer0_outputs(1791) <= '0';
    layer0_outputs(1792) <= (inputs(94)) or (inputs(60));
    layer0_outputs(1793) <= (inputs(97)) xor (inputs(240));
    layer0_outputs(1794) <= (inputs(244)) or (inputs(190));
    layer0_outputs(1795) <= not((inputs(237)) xor (inputs(173)));
    layer0_outputs(1796) <= (inputs(75)) and not (inputs(193));
    layer0_outputs(1797) <= (inputs(118)) or (inputs(19));
    layer0_outputs(1798) <= (inputs(77)) or (inputs(30));
    layer0_outputs(1799) <= (inputs(83)) and (inputs(67));
    layer0_outputs(1800) <= not(inputs(247));
    layer0_outputs(1801) <= inputs(240);
    layer0_outputs(1802) <= not(inputs(176)) or (inputs(194));
    layer0_outputs(1803) <= inputs(236);
    layer0_outputs(1804) <= not(inputs(61));
    layer0_outputs(1805) <= inputs(42);
    layer0_outputs(1806) <= (inputs(43)) xor (inputs(58));
    layer0_outputs(1807) <= (inputs(57)) or (inputs(247));
    layer0_outputs(1808) <= not(inputs(85));
    layer0_outputs(1809) <= not(inputs(30)) or (inputs(86));
    layer0_outputs(1810) <= (inputs(183)) and not (inputs(129));
    layer0_outputs(1811) <= not((inputs(213)) and (inputs(173)));
    layer0_outputs(1812) <= not((inputs(208)) xor (inputs(4)));
    layer0_outputs(1813) <= not(inputs(19));
    layer0_outputs(1814) <= (inputs(212)) and not (inputs(90));
    layer0_outputs(1815) <= not((inputs(71)) or (inputs(17)));
    layer0_outputs(1816) <= not(inputs(168)) or (inputs(63));
    layer0_outputs(1817) <= not(inputs(172)) or (inputs(154));
    layer0_outputs(1818) <= not((inputs(120)) or (inputs(241)));
    layer0_outputs(1819) <= not(inputs(69)) or (inputs(121));
    layer0_outputs(1820) <= '1';
    layer0_outputs(1821) <= inputs(206);
    layer0_outputs(1822) <= (inputs(162)) xor (inputs(113));
    layer0_outputs(1823) <= not(inputs(210));
    layer0_outputs(1824) <= not(inputs(189)) or (inputs(10));
    layer0_outputs(1825) <= not((inputs(172)) or (inputs(112)));
    layer0_outputs(1826) <= (inputs(110)) or (inputs(181));
    layer0_outputs(1827) <= not((inputs(179)) or (inputs(111)));
    layer0_outputs(1828) <= not((inputs(131)) xor (inputs(112)));
    layer0_outputs(1829) <= not((inputs(73)) or (inputs(187)));
    layer0_outputs(1830) <= not(inputs(28));
    layer0_outputs(1831) <= inputs(94);
    layer0_outputs(1832) <= not(inputs(231)) or (inputs(252));
    layer0_outputs(1833) <= (inputs(130)) or (inputs(133));
    layer0_outputs(1834) <= not((inputs(16)) or (inputs(160)));
    layer0_outputs(1835) <= not((inputs(94)) xor (inputs(25)));
    layer0_outputs(1836) <= (inputs(134)) and not (inputs(15));
    layer0_outputs(1837) <= not((inputs(161)) xor (inputs(88)));
    layer0_outputs(1838) <= inputs(252);
    layer0_outputs(1839) <= (inputs(88)) and not (inputs(28));
    layer0_outputs(1840) <= not((inputs(156)) or (inputs(93)));
    layer0_outputs(1841) <= not(inputs(116));
    layer0_outputs(1842) <= not((inputs(103)) or (inputs(67)));
    layer0_outputs(1843) <= (inputs(48)) and not (inputs(31));
    layer0_outputs(1844) <= not(inputs(233));
    layer0_outputs(1845) <= (inputs(19)) or (inputs(218));
    layer0_outputs(1846) <= not(inputs(70)) or (inputs(50));
    layer0_outputs(1847) <= (inputs(193)) or (inputs(105));
    layer0_outputs(1848) <= not(inputs(41)) or (inputs(170));
    layer0_outputs(1849) <= inputs(177);
    layer0_outputs(1850) <= (inputs(12)) and not (inputs(208));
    layer0_outputs(1851) <= inputs(155);
    layer0_outputs(1852) <= not(inputs(209));
    layer0_outputs(1853) <= inputs(126);
    layer0_outputs(1854) <= not(inputs(249));
    layer0_outputs(1855) <= (inputs(100)) and not (inputs(142));
    layer0_outputs(1856) <= (inputs(161)) or (inputs(227));
    layer0_outputs(1857) <= not(inputs(251)) or (inputs(48));
    layer0_outputs(1858) <= not((inputs(90)) xor (inputs(119)));
    layer0_outputs(1859) <= not(inputs(16));
    layer0_outputs(1860) <= (inputs(245)) or (inputs(141));
    layer0_outputs(1861) <= not(inputs(77));
    layer0_outputs(1862) <= not(inputs(37));
    layer0_outputs(1863) <= (inputs(239)) xor (inputs(206));
    layer0_outputs(1864) <= inputs(236);
    layer0_outputs(1865) <= (inputs(237)) and not (inputs(74));
    layer0_outputs(1866) <= not(inputs(197)) or (inputs(68));
    layer0_outputs(1867) <= (inputs(131)) or (inputs(65));
    layer0_outputs(1868) <= not((inputs(187)) or (inputs(37)));
    layer0_outputs(1869) <= inputs(245);
    layer0_outputs(1870) <= (inputs(16)) or (inputs(191));
    layer0_outputs(1871) <= (inputs(43)) or (inputs(22));
    layer0_outputs(1872) <= not((inputs(149)) or (inputs(229)));
    layer0_outputs(1873) <= (inputs(228)) and not (inputs(252));
    layer0_outputs(1874) <= (inputs(212)) or (inputs(187));
    layer0_outputs(1875) <= (inputs(210)) or (inputs(216));
    layer0_outputs(1876) <= not((inputs(133)) xor (inputs(152)));
    layer0_outputs(1877) <= (inputs(193)) and (inputs(193));
    layer0_outputs(1878) <= (inputs(139)) xor (inputs(164));
    layer0_outputs(1879) <= inputs(123);
    layer0_outputs(1880) <= not((inputs(175)) xor (inputs(189)));
    layer0_outputs(1881) <= not((inputs(183)) and (inputs(252)));
    layer0_outputs(1882) <= not(inputs(74)) or (inputs(156));
    layer0_outputs(1883) <= (inputs(24)) and not (inputs(129));
    layer0_outputs(1884) <= not(inputs(67));
    layer0_outputs(1885) <= (inputs(78)) and not (inputs(173));
    layer0_outputs(1886) <= not(inputs(48));
    layer0_outputs(1887) <= (inputs(8)) and not (inputs(164));
    layer0_outputs(1888) <= (inputs(86)) xor (inputs(177));
    layer0_outputs(1889) <= (inputs(205)) and not (inputs(21));
    layer0_outputs(1890) <= (inputs(161)) and not (inputs(150));
    layer0_outputs(1891) <= (inputs(107)) and not (inputs(193));
    layer0_outputs(1892) <= not((inputs(219)) or (inputs(206)));
    layer0_outputs(1893) <= not(inputs(117)) or (inputs(92));
    layer0_outputs(1894) <= not(inputs(178)) or (inputs(17));
    layer0_outputs(1895) <= not(inputs(245));
    layer0_outputs(1896) <= inputs(97);
    layer0_outputs(1897) <= not(inputs(128));
    layer0_outputs(1898) <= (inputs(151)) or (inputs(55));
    layer0_outputs(1899) <= inputs(147);
    layer0_outputs(1900) <= (inputs(103)) or (inputs(77));
    layer0_outputs(1901) <= (inputs(157)) or (inputs(79));
    layer0_outputs(1902) <= (inputs(60)) or (inputs(77));
    layer0_outputs(1903) <= not(inputs(150));
    layer0_outputs(1904) <= not(inputs(252)) or (inputs(252));
    layer0_outputs(1905) <= (inputs(21)) or (inputs(121));
    layer0_outputs(1906) <= not(inputs(100));
    layer0_outputs(1907) <= (inputs(237)) and not (inputs(74));
    layer0_outputs(1908) <= not(inputs(8)) or (inputs(15));
    layer0_outputs(1909) <= not(inputs(165));
    layer0_outputs(1910) <= (inputs(173)) xor (inputs(215));
    layer0_outputs(1911) <= inputs(37);
    layer0_outputs(1912) <= (inputs(41)) xor (inputs(9));
    layer0_outputs(1913) <= (inputs(165)) or (inputs(148));
    layer0_outputs(1914) <= not((inputs(37)) xor (inputs(82)));
    layer0_outputs(1915) <= not(inputs(178));
    layer0_outputs(1916) <= not(inputs(193));
    layer0_outputs(1917) <= not(inputs(164));
    layer0_outputs(1918) <= not(inputs(119)) or (inputs(163));
    layer0_outputs(1919) <= not((inputs(49)) or (inputs(192)));
    layer0_outputs(1920) <= not(inputs(199)) or (inputs(217));
    layer0_outputs(1921) <= (inputs(152)) and not (inputs(26));
    layer0_outputs(1922) <= (inputs(84)) or (inputs(156));
    layer0_outputs(1923) <= not(inputs(47));
    layer0_outputs(1924) <= (inputs(208)) or (inputs(192));
    layer0_outputs(1925) <= (inputs(205)) and not (inputs(32));
    layer0_outputs(1926) <= not(inputs(25));
    layer0_outputs(1927) <= not(inputs(51)) or (inputs(168));
    layer0_outputs(1928) <= (inputs(161)) or (inputs(178));
    layer0_outputs(1929) <= (inputs(208)) or (inputs(5));
    layer0_outputs(1930) <= (inputs(128)) xor (inputs(33));
    layer0_outputs(1931) <= not(inputs(3));
    layer0_outputs(1932) <= not(inputs(115)) or (inputs(17));
    layer0_outputs(1933) <= not((inputs(120)) or (inputs(96)));
    layer0_outputs(1934) <= (inputs(147)) or (inputs(115));
    layer0_outputs(1935) <= not(inputs(45)) or (inputs(41));
    layer0_outputs(1936) <= (inputs(76)) xor (inputs(235));
    layer0_outputs(1937) <= not(inputs(163)) or (inputs(167));
    layer0_outputs(1938) <= (inputs(198)) and not (inputs(93));
    layer0_outputs(1939) <= inputs(141);
    layer0_outputs(1940) <= not(inputs(34)) or (inputs(66));
    layer0_outputs(1941) <= not(inputs(135));
    layer0_outputs(1942) <= (inputs(106)) xor (inputs(180));
    layer0_outputs(1943) <= not(inputs(88)) or (inputs(225));
    layer0_outputs(1944) <= (inputs(155)) and not (inputs(110));
    layer0_outputs(1945) <= not(inputs(71));
    layer0_outputs(1946) <= (inputs(229)) or (inputs(208));
    layer0_outputs(1947) <= not(inputs(211)) or (inputs(22));
    layer0_outputs(1948) <= (inputs(84)) xor (inputs(21));
    layer0_outputs(1949) <= not((inputs(147)) or (inputs(156)));
    layer0_outputs(1950) <= (inputs(208)) and not (inputs(0));
    layer0_outputs(1951) <= not((inputs(169)) or (inputs(150)));
    layer0_outputs(1952) <= not(inputs(228));
    layer0_outputs(1953) <= not(inputs(67));
    layer0_outputs(1954) <= '1';
    layer0_outputs(1955) <= not(inputs(67));
    layer0_outputs(1956) <= inputs(123);
    layer0_outputs(1957) <= not(inputs(41)) or (inputs(111));
    layer0_outputs(1958) <= (inputs(6)) or (inputs(227));
    layer0_outputs(1959) <= inputs(4);
    layer0_outputs(1960) <= inputs(220);
    layer0_outputs(1961) <= inputs(92);
    layer0_outputs(1962) <= inputs(171);
    layer0_outputs(1963) <= (inputs(236)) or (inputs(55));
    layer0_outputs(1964) <= inputs(255);
    layer0_outputs(1965) <= (inputs(118)) or (inputs(251));
    layer0_outputs(1966) <= inputs(148);
    layer0_outputs(1967) <= not((inputs(112)) or (inputs(247)));
    layer0_outputs(1968) <= not(inputs(27));
    layer0_outputs(1969) <= not(inputs(244)) or (inputs(203));
    layer0_outputs(1970) <= (inputs(34)) or (inputs(69));
    layer0_outputs(1971) <= not(inputs(87));
    layer0_outputs(1972) <= (inputs(130)) and not (inputs(32));
    layer0_outputs(1973) <= (inputs(192)) or (inputs(17));
    layer0_outputs(1974) <= (inputs(103)) and not (inputs(109));
    layer0_outputs(1975) <= not(inputs(106));
    layer0_outputs(1976) <= not((inputs(243)) and (inputs(16)));
    layer0_outputs(1977) <= (inputs(55)) xor (inputs(10));
    layer0_outputs(1978) <= inputs(141);
    layer0_outputs(1979) <= (inputs(242)) and not (inputs(66));
    layer0_outputs(1980) <= not((inputs(146)) or (inputs(179)));
    layer0_outputs(1981) <= not((inputs(115)) or (inputs(101)));
    layer0_outputs(1982) <= not(inputs(134)) or (inputs(144));
    layer0_outputs(1983) <= not(inputs(82));
    layer0_outputs(1984) <= not(inputs(97));
    layer0_outputs(1985) <= not(inputs(237));
    layer0_outputs(1986) <= (inputs(122)) and not (inputs(81));
    layer0_outputs(1987) <= not(inputs(149)) or (inputs(206));
    layer0_outputs(1988) <= '1';
    layer0_outputs(1989) <= not(inputs(193));
    layer0_outputs(1990) <= not(inputs(108)) or (inputs(39));
    layer0_outputs(1991) <= (inputs(179)) or (inputs(111));
    layer0_outputs(1992) <= '0';
    layer0_outputs(1993) <= not(inputs(183)) or (inputs(112));
    layer0_outputs(1994) <= (inputs(231)) or (inputs(176));
    layer0_outputs(1995) <= not(inputs(104));
    layer0_outputs(1996) <= '0';
    layer0_outputs(1997) <= (inputs(7)) or (inputs(75));
    layer0_outputs(1998) <= (inputs(171)) and (inputs(224));
    layer0_outputs(1999) <= (inputs(20)) or (inputs(70));
    layer0_outputs(2000) <= (inputs(67)) and not (inputs(65));
    layer0_outputs(2001) <= not((inputs(184)) or (inputs(127)));
    layer0_outputs(2002) <= not((inputs(183)) or (inputs(55)));
    layer0_outputs(2003) <= not((inputs(180)) xor (inputs(177)));
    layer0_outputs(2004) <= not((inputs(244)) or (inputs(95)));
    layer0_outputs(2005) <= '0';
    layer0_outputs(2006) <= '1';
    layer0_outputs(2007) <= not((inputs(118)) and (inputs(51)));
    layer0_outputs(2008) <= not(inputs(66)) or (inputs(142));
    layer0_outputs(2009) <= '0';
    layer0_outputs(2010) <= (inputs(117)) or (inputs(221));
    layer0_outputs(2011) <= not(inputs(117)) or (inputs(121));
    layer0_outputs(2012) <= (inputs(28)) or (inputs(244));
    layer0_outputs(2013) <= (inputs(146)) or (inputs(219));
    layer0_outputs(2014) <= (inputs(32)) and not (inputs(79));
    layer0_outputs(2015) <= (inputs(242)) or (inputs(194));
    layer0_outputs(2016) <= (inputs(9)) xor (inputs(57));
    layer0_outputs(2017) <= not(inputs(16));
    layer0_outputs(2018) <= (inputs(208)) and not (inputs(200));
    layer0_outputs(2019) <= not(inputs(170));
    layer0_outputs(2020) <= (inputs(17)) xor (inputs(171));
    layer0_outputs(2021) <= inputs(14);
    layer0_outputs(2022) <= not(inputs(230));
    layer0_outputs(2023) <= not(inputs(167));
    layer0_outputs(2024) <= (inputs(56)) or (inputs(228));
    layer0_outputs(2025) <= (inputs(31)) or (inputs(43));
    layer0_outputs(2026) <= not((inputs(89)) or (inputs(99)));
    layer0_outputs(2027) <= (inputs(139)) and not (inputs(224));
    layer0_outputs(2028) <= not(inputs(239));
    layer0_outputs(2029) <= not((inputs(35)) xor (inputs(220)));
    layer0_outputs(2030) <= not(inputs(35));
    layer0_outputs(2031) <= not((inputs(0)) xor (inputs(221)));
    layer0_outputs(2032) <= not(inputs(25));
    layer0_outputs(2033) <= (inputs(171)) and (inputs(245));
    layer0_outputs(2034) <= not(inputs(130));
    layer0_outputs(2035) <= not(inputs(26));
    layer0_outputs(2036) <= inputs(168);
    layer0_outputs(2037) <= (inputs(237)) or (inputs(149));
    layer0_outputs(2038) <= not(inputs(153));
    layer0_outputs(2039) <= (inputs(162)) or (inputs(176));
    layer0_outputs(2040) <= inputs(254);
    layer0_outputs(2041) <= not(inputs(67));
    layer0_outputs(2042) <= (inputs(132)) xor (inputs(149));
    layer0_outputs(2043) <= not(inputs(46));
    layer0_outputs(2044) <= not((inputs(85)) and (inputs(62)));
    layer0_outputs(2045) <= not(inputs(228)) or (inputs(53));
    layer0_outputs(2046) <= inputs(7);
    layer0_outputs(2047) <= not((inputs(146)) or (inputs(175)));
    layer0_outputs(2048) <= '0';
    layer0_outputs(2049) <= (inputs(131)) xor (inputs(21));
    layer0_outputs(2050) <= not(inputs(164));
    layer0_outputs(2051) <= not(inputs(197));
    layer0_outputs(2052) <= inputs(178);
    layer0_outputs(2053) <= (inputs(189)) and not (inputs(12));
    layer0_outputs(2054) <= not(inputs(255)) or (inputs(122));
    layer0_outputs(2055) <= not((inputs(248)) or (inputs(42)));
    layer0_outputs(2056) <= not(inputs(91));
    layer0_outputs(2057) <= inputs(93);
    layer0_outputs(2058) <= not((inputs(178)) xor (inputs(232)));
    layer0_outputs(2059) <= not(inputs(159)) or (inputs(64));
    layer0_outputs(2060) <= inputs(121);
    layer0_outputs(2061) <= not(inputs(117));
    layer0_outputs(2062) <= inputs(67);
    layer0_outputs(2063) <= not(inputs(117));
    layer0_outputs(2064) <= not((inputs(227)) and (inputs(247)));
    layer0_outputs(2065) <= not((inputs(214)) xor (inputs(199)));
    layer0_outputs(2066) <= (inputs(86)) and not (inputs(150));
    layer0_outputs(2067) <= not((inputs(65)) or (inputs(164)));
    layer0_outputs(2068) <= not(inputs(160)) or (inputs(255));
    layer0_outputs(2069) <= not((inputs(181)) xor (inputs(208)));
    layer0_outputs(2070) <= not(inputs(126));
    layer0_outputs(2071) <= not(inputs(57));
    layer0_outputs(2072) <= (inputs(204)) and not (inputs(41));
    layer0_outputs(2073) <= (inputs(128)) and (inputs(210));
    layer0_outputs(2074) <= not((inputs(130)) xor (inputs(147)));
    layer0_outputs(2075) <= not((inputs(203)) xor (inputs(97)));
    layer0_outputs(2076) <= (inputs(199)) or (inputs(184));
    layer0_outputs(2077) <= '0';
    layer0_outputs(2078) <= not((inputs(247)) or (inputs(18)));
    layer0_outputs(2079) <= not(inputs(82)) or (inputs(24));
    layer0_outputs(2080) <= (inputs(232)) xor (inputs(113));
    layer0_outputs(2081) <= not((inputs(3)) or (inputs(186)));
    layer0_outputs(2082) <= not(inputs(3)) or (inputs(112));
    layer0_outputs(2083) <= inputs(81);
    layer0_outputs(2084) <= (inputs(152)) and not (inputs(9));
    layer0_outputs(2085) <= not((inputs(254)) or (inputs(253)));
    layer0_outputs(2086) <= not(inputs(186)) or (inputs(5));
    layer0_outputs(2087) <= not(inputs(167)) or (inputs(190));
    layer0_outputs(2088) <= (inputs(208)) xor (inputs(212));
    layer0_outputs(2089) <= not(inputs(213)) or (inputs(30));
    layer0_outputs(2090) <= inputs(208);
    layer0_outputs(2091) <= not(inputs(167)) or (inputs(143));
    layer0_outputs(2092) <= inputs(114);
    layer0_outputs(2093) <= (inputs(23)) or (inputs(124));
    layer0_outputs(2094) <= not(inputs(193)) or (inputs(11));
    layer0_outputs(2095) <= '1';
    layer0_outputs(2096) <= not((inputs(77)) or (inputs(109)));
    layer0_outputs(2097) <= not((inputs(240)) xor (inputs(154)));
    layer0_outputs(2098) <= '1';
    layer0_outputs(2099) <= (inputs(205)) and not (inputs(112));
    layer0_outputs(2100) <= (inputs(28)) xor (inputs(103));
    layer0_outputs(2101) <= not(inputs(34)) or (inputs(202));
    layer0_outputs(2102) <= not(inputs(41)) or (inputs(224));
    layer0_outputs(2103) <= not((inputs(99)) and (inputs(121)));
    layer0_outputs(2104) <= inputs(65);
    layer0_outputs(2105) <= '0';
    layer0_outputs(2106) <= (inputs(45)) and not (inputs(241));
    layer0_outputs(2107) <= inputs(81);
    layer0_outputs(2108) <= (inputs(122)) and not (inputs(97));
    layer0_outputs(2109) <= not(inputs(74));
    layer0_outputs(2110) <= (inputs(172)) or (inputs(226));
    layer0_outputs(2111) <= (inputs(240)) and not (inputs(191));
    layer0_outputs(2112) <= not(inputs(222)) or (inputs(114));
    layer0_outputs(2113) <= (inputs(243)) or (inputs(208));
    layer0_outputs(2114) <= not((inputs(207)) xor (inputs(236)));
    layer0_outputs(2115) <= not((inputs(91)) or (inputs(236)));
    layer0_outputs(2116) <= not((inputs(212)) xor (inputs(234)));
    layer0_outputs(2117) <= not(inputs(7));
    layer0_outputs(2118) <= not(inputs(83)) or (inputs(96));
    layer0_outputs(2119) <= not(inputs(139));
    layer0_outputs(2120) <= not(inputs(108)) or (inputs(223));
    layer0_outputs(2121) <= (inputs(127)) and not (inputs(11));
    layer0_outputs(2122) <= not((inputs(246)) and (inputs(80)));
    layer0_outputs(2123) <= inputs(182);
    layer0_outputs(2124) <= not(inputs(227)) or (inputs(82));
    layer0_outputs(2125) <= not((inputs(225)) or (inputs(152)));
    layer0_outputs(2126) <= not((inputs(117)) or (inputs(113)));
    layer0_outputs(2127) <= not(inputs(218)) or (inputs(31));
    layer0_outputs(2128) <= not((inputs(3)) or (inputs(96)));
    layer0_outputs(2129) <= inputs(113);
    layer0_outputs(2130) <= inputs(72);
    layer0_outputs(2131) <= '1';
    layer0_outputs(2132) <= inputs(212);
    layer0_outputs(2133) <= '1';
    layer0_outputs(2134) <= not(inputs(123));
    layer0_outputs(2135) <= (inputs(196)) and not (inputs(76));
    layer0_outputs(2136) <= not((inputs(211)) or (inputs(87)));
    layer0_outputs(2137) <= inputs(212);
    layer0_outputs(2138) <= not(inputs(20));
    layer0_outputs(2139) <= not(inputs(216)) or (inputs(246));
    layer0_outputs(2140) <= (inputs(250)) or (inputs(189));
    layer0_outputs(2141) <= not((inputs(139)) xor (inputs(164)));
    layer0_outputs(2142) <= (inputs(9)) and not (inputs(63));
    layer0_outputs(2143) <= not((inputs(196)) or (inputs(112)));
    layer0_outputs(2144) <= (inputs(46)) and not (inputs(145));
    layer0_outputs(2145) <= not(inputs(23));
    layer0_outputs(2146) <= (inputs(74)) and (inputs(13));
    layer0_outputs(2147) <= not((inputs(30)) and (inputs(123)));
    layer0_outputs(2148) <= not((inputs(57)) and (inputs(3)));
    layer0_outputs(2149) <= (inputs(199)) and not (inputs(255));
    layer0_outputs(2150) <= not(inputs(198)) or (inputs(16));
    layer0_outputs(2151) <= (inputs(160)) and not (inputs(147));
    layer0_outputs(2152) <= not(inputs(73));
    layer0_outputs(2153) <= not(inputs(182));
    layer0_outputs(2154) <= (inputs(205)) xor (inputs(21));
    layer0_outputs(2155) <= (inputs(216)) or (inputs(246));
    layer0_outputs(2156) <= not(inputs(162));
    layer0_outputs(2157) <= (inputs(201)) or (inputs(227));
    layer0_outputs(2158) <= inputs(234);
    layer0_outputs(2159) <= not(inputs(21)) or (inputs(228));
    layer0_outputs(2160) <= (inputs(253)) and not (inputs(187));
    layer0_outputs(2161) <= not((inputs(74)) or (inputs(167)));
    layer0_outputs(2162) <= not(inputs(229)) or (inputs(103));
    layer0_outputs(2163) <= not((inputs(15)) or (inputs(4)));
    layer0_outputs(2164) <= not((inputs(109)) xor (inputs(41)));
    layer0_outputs(2165) <= not(inputs(48));
    layer0_outputs(2166) <= (inputs(80)) or (inputs(9));
    layer0_outputs(2167) <= (inputs(194)) or (inputs(249));
    layer0_outputs(2168) <= (inputs(104)) and not (inputs(190));
    layer0_outputs(2169) <= (inputs(159)) xor (inputs(106));
    layer0_outputs(2170) <= not((inputs(107)) and (inputs(37)));
    layer0_outputs(2171) <= (inputs(236)) or (inputs(173));
    layer0_outputs(2172) <= (inputs(166)) and not (inputs(214));
    layer0_outputs(2173) <= (inputs(36)) xor (inputs(97));
    layer0_outputs(2174) <= (inputs(236)) xor (inputs(10));
    layer0_outputs(2175) <= (inputs(89)) xor (inputs(106));
    layer0_outputs(2176) <= inputs(60);
    layer0_outputs(2177) <= not(inputs(65));
    layer0_outputs(2178) <= not((inputs(230)) or (inputs(176)));
    layer0_outputs(2179) <= inputs(232);
    layer0_outputs(2180) <= inputs(164);
    layer0_outputs(2181) <= (inputs(229)) and not (inputs(37));
    layer0_outputs(2182) <= (inputs(135)) and not (inputs(62));
    layer0_outputs(2183) <= not((inputs(69)) xor (inputs(226)));
    layer0_outputs(2184) <= inputs(151);
    layer0_outputs(2185) <= not((inputs(148)) xor (inputs(155)));
    layer0_outputs(2186) <= not(inputs(86));
    layer0_outputs(2187) <= inputs(149);
    layer0_outputs(2188) <= (inputs(12)) or (inputs(227));
    layer0_outputs(2189) <= inputs(27);
    layer0_outputs(2190) <= not((inputs(32)) or (inputs(208)));
    layer0_outputs(2191) <= (inputs(116)) and not (inputs(0));
    layer0_outputs(2192) <= not(inputs(92)) or (inputs(180));
    layer0_outputs(2193) <= (inputs(234)) and not (inputs(150));
    layer0_outputs(2194) <= not((inputs(117)) xor (inputs(239)));
    layer0_outputs(2195) <= (inputs(192)) and not (inputs(0));
    layer0_outputs(2196) <= not((inputs(175)) or (inputs(158)));
    layer0_outputs(2197) <= not((inputs(133)) xor (inputs(177)));
    layer0_outputs(2198) <= (inputs(217)) xor (inputs(163));
    layer0_outputs(2199) <= inputs(199);
    layer0_outputs(2200) <= (inputs(198)) and not (inputs(208));
    layer0_outputs(2201) <= not((inputs(60)) xor (inputs(43)));
    layer0_outputs(2202) <= (inputs(162)) or (inputs(176));
    layer0_outputs(2203) <= not((inputs(155)) or (inputs(52)));
    layer0_outputs(2204) <= inputs(159);
    layer0_outputs(2205) <= not((inputs(190)) or (inputs(150)));
    layer0_outputs(2206) <= (inputs(220)) and not (inputs(243));
    layer0_outputs(2207) <= (inputs(83)) xor (inputs(84));
    layer0_outputs(2208) <= inputs(234);
    layer0_outputs(2209) <= not(inputs(85));
    layer0_outputs(2210) <= (inputs(127)) and not (inputs(251));
    layer0_outputs(2211) <= (inputs(130)) and not (inputs(39));
    layer0_outputs(2212) <= inputs(101);
    layer0_outputs(2213) <= not((inputs(77)) or (inputs(176)));
    layer0_outputs(2214) <= not(inputs(184));
    layer0_outputs(2215) <= (inputs(185)) xor (inputs(80));
    layer0_outputs(2216) <= not(inputs(91)) or (inputs(40));
    layer0_outputs(2217) <= inputs(141);
    layer0_outputs(2218) <= not(inputs(161));
    layer0_outputs(2219) <= inputs(117);
    layer0_outputs(2220) <= (inputs(64)) xor (inputs(5));
    layer0_outputs(2221) <= not(inputs(139));
    layer0_outputs(2222) <= (inputs(177)) xor (inputs(136));
    layer0_outputs(2223) <= not((inputs(230)) xor (inputs(190)));
    layer0_outputs(2224) <= inputs(127);
    layer0_outputs(2225) <= not((inputs(81)) or (inputs(124)));
    layer0_outputs(2226) <= not((inputs(0)) or (inputs(30)));
    layer0_outputs(2227) <= '0';
    layer0_outputs(2228) <= not(inputs(19));
    layer0_outputs(2229) <= (inputs(88)) and not (inputs(85));
    layer0_outputs(2230) <= inputs(164);
    layer0_outputs(2231) <= (inputs(56)) and not (inputs(197));
    layer0_outputs(2232) <= (inputs(13)) and (inputs(243));
    layer0_outputs(2233) <= not(inputs(48));
    layer0_outputs(2234) <= not((inputs(198)) or (inputs(47)));
    layer0_outputs(2235) <= not(inputs(211)) or (inputs(108));
    layer0_outputs(2236) <= (inputs(111)) or (inputs(165));
    layer0_outputs(2237) <= inputs(16);
    layer0_outputs(2238) <= not((inputs(122)) xor (inputs(93)));
    layer0_outputs(2239) <= (inputs(42)) or (inputs(241));
    layer0_outputs(2240) <= (inputs(64)) and not (inputs(173));
    layer0_outputs(2241) <= '0';
    layer0_outputs(2242) <= inputs(220);
    layer0_outputs(2243) <= not(inputs(74));
    layer0_outputs(2244) <= not(inputs(10));
    layer0_outputs(2245) <= (inputs(213)) xor (inputs(200));
    layer0_outputs(2246) <= not(inputs(240)) or (inputs(50));
    layer0_outputs(2247) <= (inputs(116)) and not (inputs(4));
    layer0_outputs(2248) <= not(inputs(231)) or (inputs(237));
    layer0_outputs(2249) <= (inputs(31)) xor (inputs(166));
    layer0_outputs(2250) <= not(inputs(140)) or (inputs(61));
    layer0_outputs(2251) <= inputs(114);
    layer0_outputs(2252) <= (inputs(228)) or (inputs(251));
    layer0_outputs(2253) <= (inputs(214)) and not (inputs(15));
    layer0_outputs(2254) <= not(inputs(94));
    layer0_outputs(2255) <= (inputs(77)) xor (inputs(228));
    layer0_outputs(2256) <= inputs(66);
    layer0_outputs(2257) <= (inputs(86)) and not (inputs(160));
    layer0_outputs(2258) <= inputs(175);
    layer0_outputs(2259) <= (inputs(47)) or (inputs(15));
    layer0_outputs(2260) <= (inputs(179)) and not (inputs(34));
    layer0_outputs(2261) <= not(inputs(109)) or (inputs(154));
    layer0_outputs(2262) <= inputs(247);
    layer0_outputs(2263) <= (inputs(107)) and not (inputs(205));
    layer0_outputs(2264) <= not((inputs(145)) xor (inputs(143)));
    layer0_outputs(2265) <= inputs(157);
    layer0_outputs(2266) <= not(inputs(214));
    layer0_outputs(2267) <= not(inputs(163));
    layer0_outputs(2268) <= not(inputs(164));
    layer0_outputs(2269) <= not(inputs(188));
    layer0_outputs(2270) <= not((inputs(194)) or (inputs(31)));
    layer0_outputs(2271) <= not(inputs(150)) or (inputs(155));
    layer0_outputs(2272) <= not(inputs(206)) or (inputs(39));
    layer0_outputs(2273) <= '1';
    layer0_outputs(2274) <= inputs(22);
    layer0_outputs(2275) <= (inputs(145)) xor (inputs(204));
    layer0_outputs(2276) <= not((inputs(230)) and (inputs(124)));
    layer0_outputs(2277) <= not(inputs(56)) or (inputs(247));
    layer0_outputs(2278) <= (inputs(1)) xor (inputs(226));
    layer0_outputs(2279) <= (inputs(74)) or (inputs(106));
    layer0_outputs(2280) <= (inputs(195)) and not (inputs(79));
    layer0_outputs(2281) <= '0';
    layer0_outputs(2282) <= inputs(248);
    layer0_outputs(2283) <= (inputs(27)) xor (inputs(78));
    layer0_outputs(2284) <= not((inputs(41)) and (inputs(75)));
    layer0_outputs(2285) <= not((inputs(130)) xor (inputs(245)));
    layer0_outputs(2286) <= not((inputs(238)) and (inputs(59)));
    layer0_outputs(2287) <= not(inputs(129)) or (inputs(181));
    layer0_outputs(2288) <= not(inputs(194));
    layer0_outputs(2289) <= not(inputs(129));
    layer0_outputs(2290) <= (inputs(2)) or (inputs(39));
    layer0_outputs(2291) <= not((inputs(202)) and (inputs(242)));
    layer0_outputs(2292) <= not((inputs(230)) xor (inputs(230)));
    layer0_outputs(2293) <= not(inputs(84));
    layer0_outputs(2294) <= (inputs(129)) xor (inputs(252));
    layer0_outputs(2295) <= (inputs(33)) and not (inputs(6));
    layer0_outputs(2296) <= not((inputs(150)) or (inputs(82)));
    layer0_outputs(2297) <= (inputs(116)) and not (inputs(5));
    layer0_outputs(2298) <= (inputs(245)) and not (inputs(186));
    layer0_outputs(2299) <= not(inputs(180)) or (inputs(160));
    layer0_outputs(2300) <= inputs(98);
    layer0_outputs(2301) <= not(inputs(55)) or (inputs(38));
    layer0_outputs(2302) <= not((inputs(162)) xor (inputs(229)));
    layer0_outputs(2303) <= not(inputs(74));
    layer0_outputs(2304) <= (inputs(157)) and (inputs(144));
    layer0_outputs(2305) <= not(inputs(23));
    layer0_outputs(2306) <= not(inputs(250)) or (inputs(9));
    layer0_outputs(2307) <= not(inputs(91)) or (inputs(208));
    layer0_outputs(2308) <= (inputs(57)) and not (inputs(168));
    layer0_outputs(2309) <= not((inputs(156)) xor (inputs(35)));
    layer0_outputs(2310) <= inputs(121);
    layer0_outputs(2311) <= not(inputs(99));
    layer0_outputs(2312) <= not((inputs(95)) or (inputs(32)));
    layer0_outputs(2313) <= '0';
    layer0_outputs(2314) <= (inputs(96)) and not (inputs(113));
    layer0_outputs(2315) <= (inputs(126)) and (inputs(92));
    layer0_outputs(2316) <= inputs(76);
    layer0_outputs(2317) <= not(inputs(82)) or (inputs(171));
    layer0_outputs(2318) <= not(inputs(112)) or (inputs(210));
    layer0_outputs(2319) <= not(inputs(154));
    layer0_outputs(2320) <= '1';
    layer0_outputs(2321) <= (inputs(25)) and not (inputs(155));
    layer0_outputs(2322) <= (inputs(137)) or (inputs(170));
    layer0_outputs(2323) <= inputs(94);
    layer0_outputs(2324) <= not(inputs(30)) or (inputs(10));
    layer0_outputs(2325) <= not(inputs(83));
    layer0_outputs(2326) <= not((inputs(41)) or (inputs(14)));
    layer0_outputs(2327) <= not((inputs(107)) xor (inputs(142)));
    layer0_outputs(2328) <= not(inputs(166)) or (inputs(238));
    layer0_outputs(2329) <= not(inputs(1)) or (inputs(207));
    layer0_outputs(2330) <= inputs(182);
    layer0_outputs(2331) <= (inputs(201)) or (inputs(6));
    layer0_outputs(2332) <= (inputs(50)) and (inputs(152));
    layer0_outputs(2333) <= not(inputs(238)) or (inputs(87));
    layer0_outputs(2334) <= (inputs(227)) and not (inputs(252));
    layer0_outputs(2335) <= not(inputs(98)) or (inputs(17));
    layer0_outputs(2336) <= not((inputs(146)) xor (inputs(87)));
    layer0_outputs(2337) <= not(inputs(68));
    layer0_outputs(2338) <= not(inputs(213)) or (inputs(146));
    layer0_outputs(2339) <= not(inputs(135));
    layer0_outputs(2340) <= (inputs(75)) xor (inputs(47));
    layer0_outputs(2341) <= (inputs(180)) or (inputs(106));
    layer0_outputs(2342) <= (inputs(126)) and not (inputs(19));
    layer0_outputs(2343) <= (inputs(71)) or (inputs(71));
    layer0_outputs(2344) <= (inputs(64)) and not (inputs(206));
    layer0_outputs(2345) <= (inputs(23)) and not (inputs(32));
    layer0_outputs(2346) <= (inputs(230)) and not (inputs(152));
    layer0_outputs(2347) <= not(inputs(181));
    layer0_outputs(2348) <= (inputs(162)) xor (inputs(249));
    layer0_outputs(2349) <= (inputs(176)) or (inputs(1));
    layer0_outputs(2350) <= not(inputs(91)) or (inputs(158));
    layer0_outputs(2351) <= not(inputs(10));
    layer0_outputs(2352) <= not((inputs(177)) xor (inputs(20)));
    layer0_outputs(2353) <= not((inputs(81)) or (inputs(39)));
    layer0_outputs(2354) <= not((inputs(231)) or (inputs(132)));
    layer0_outputs(2355) <= '0';
    layer0_outputs(2356) <= (inputs(197)) and not (inputs(124));
    layer0_outputs(2357) <= not((inputs(137)) or (inputs(63)));
    layer0_outputs(2358) <= not(inputs(101));
    layer0_outputs(2359) <= not(inputs(72));
    layer0_outputs(2360) <= '1';
    layer0_outputs(2361) <= (inputs(199)) xor (inputs(1));
    layer0_outputs(2362) <= (inputs(147)) and not (inputs(93));
    layer0_outputs(2363) <= (inputs(83)) xor (inputs(190));
    layer0_outputs(2364) <= not((inputs(96)) or (inputs(151)));
    layer0_outputs(2365) <= (inputs(38)) and (inputs(122));
    layer0_outputs(2366) <= (inputs(77)) and (inputs(232));
    layer0_outputs(2367) <= (inputs(38)) and not (inputs(70));
    layer0_outputs(2368) <= not(inputs(182)) or (inputs(127));
    layer0_outputs(2369) <= not(inputs(42));
    layer0_outputs(2370) <= (inputs(174)) or (inputs(169));
    layer0_outputs(2371) <= not(inputs(99));
    layer0_outputs(2372) <= not(inputs(204)) or (inputs(14));
    layer0_outputs(2373) <= (inputs(91)) and (inputs(247));
    layer0_outputs(2374) <= (inputs(120)) and not (inputs(16));
    layer0_outputs(2375) <= not((inputs(97)) xor (inputs(228)));
    layer0_outputs(2376) <= (inputs(139)) xor (inputs(61));
    layer0_outputs(2377) <= not((inputs(254)) or (inputs(46)));
    layer0_outputs(2378) <= not((inputs(225)) xor (inputs(162)));
    layer0_outputs(2379) <= not(inputs(77)) or (inputs(235));
    layer0_outputs(2380) <= not((inputs(32)) or (inputs(52)));
    layer0_outputs(2381) <= not((inputs(80)) xor (inputs(84)));
    layer0_outputs(2382) <= not(inputs(146));
    layer0_outputs(2383) <= not(inputs(189));
    layer0_outputs(2384) <= not((inputs(81)) or (inputs(211)));
    layer0_outputs(2385) <= (inputs(8)) and not (inputs(42));
    layer0_outputs(2386) <= inputs(244);
    layer0_outputs(2387) <= '0';
    layer0_outputs(2388) <= '1';
    layer0_outputs(2389) <= (inputs(81)) and (inputs(158));
    layer0_outputs(2390) <= not((inputs(160)) or (inputs(147)));
    layer0_outputs(2391) <= not(inputs(41));
    layer0_outputs(2392) <= (inputs(76)) or (inputs(101));
    layer0_outputs(2393) <= inputs(106);
    layer0_outputs(2394) <= (inputs(49)) and not (inputs(15));
    layer0_outputs(2395) <= (inputs(52)) xor (inputs(80));
    layer0_outputs(2396) <= '1';
    layer0_outputs(2397) <= '1';
    layer0_outputs(2398) <= inputs(32);
    layer0_outputs(2399) <= not((inputs(171)) xor (inputs(218)));
    layer0_outputs(2400) <= not(inputs(55));
    layer0_outputs(2401) <= inputs(54);
    layer0_outputs(2402) <= (inputs(135)) or (inputs(122));
    layer0_outputs(2403) <= '1';
    layer0_outputs(2404) <= not((inputs(248)) xor (inputs(208)));
    layer0_outputs(2405) <= not(inputs(39));
    layer0_outputs(2406) <= inputs(168);
    layer0_outputs(2407) <= not(inputs(48));
    layer0_outputs(2408) <= not(inputs(84));
    layer0_outputs(2409) <= (inputs(119)) and (inputs(159));
    layer0_outputs(2410) <= not((inputs(132)) or (inputs(249)));
    layer0_outputs(2411) <= not(inputs(70)) or (inputs(60));
    layer0_outputs(2412) <= inputs(63);
    layer0_outputs(2413) <= not((inputs(128)) or (inputs(75)));
    layer0_outputs(2414) <= not((inputs(8)) and (inputs(222)));
    layer0_outputs(2415) <= not((inputs(140)) xor (inputs(142)));
    layer0_outputs(2416) <= not(inputs(106)) or (inputs(185));
    layer0_outputs(2417) <= inputs(153);
    layer0_outputs(2418) <= (inputs(194)) and not (inputs(11));
    layer0_outputs(2419) <= (inputs(110)) xor (inputs(49));
    layer0_outputs(2420) <= not(inputs(55));
    layer0_outputs(2421) <= (inputs(49)) or (inputs(216));
    layer0_outputs(2422) <= (inputs(213)) or (inputs(141));
    layer0_outputs(2423) <= not(inputs(100));
    layer0_outputs(2424) <= not(inputs(196));
    layer0_outputs(2425) <= not(inputs(101)) or (inputs(33));
    layer0_outputs(2426) <= (inputs(24)) and not (inputs(135));
    layer0_outputs(2427) <= not(inputs(94));
    layer0_outputs(2428) <= '1';
    layer0_outputs(2429) <= (inputs(40)) xor (inputs(24));
    layer0_outputs(2430) <= not(inputs(165));
    layer0_outputs(2431) <= not((inputs(59)) xor (inputs(223)));
    layer0_outputs(2432) <= not(inputs(49));
    layer0_outputs(2433) <= inputs(140);
    layer0_outputs(2434) <= (inputs(224)) and not (inputs(112));
    layer0_outputs(2435) <= not((inputs(41)) xor (inputs(215)));
    layer0_outputs(2436) <= (inputs(96)) xor (inputs(247));
    layer0_outputs(2437) <= inputs(235);
    layer0_outputs(2438) <= inputs(21);
    layer0_outputs(2439) <= inputs(76);
    layer0_outputs(2440) <= not((inputs(186)) xor (inputs(174)));
    layer0_outputs(2441) <= not(inputs(69));
    layer0_outputs(2442) <= not((inputs(78)) or (inputs(40)));
    layer0_outputs(2443) <= not((inputs(112)) or (inputs(125)));
    layer0_outputs(2444) <= not((inputs(51)) or (inputs(237)));
    layer0_outputs(2445) <= not((inputs(233)) and (inputs(77)));
    layer0_outputs(2446) <= not(inputs(234));
    layer0_outputs(2447) <= not(inputs(114)) or (inputs(243));
    layer0_outputs(2448) <= not((inputs(170)) or (inputs(8)));
    layer0_outputs(2449) <= '1';
    layer0_outputs(2450) <= (inputs(218)) and (inputs(159));
    layer0_outputs(2451) <= inputs(160);
    layer0_outputs(2452) <= (inputs(59)) or (inputs(59));
    layer0_outputs(2453) <= not(inputs(39));
    layer0_outputs(2454) <= not(inputs(114));
    layer0_outputs(2455) <= not((inputs(22)) or (inputs(38)));
    layer0_outputs(2456) <= (inputs(77)) or (inputs(146));
    layer0_outputs(2457) <= (inputs(160)) and not (inputs(202));
    layer0_outputs(2458) <= not((inputs(171)) xor (inputs(217)));
    layer0_outputs(2459) <= (inputs(121)) or (inputs(180));
    layer0_outputs(2460) <= not(inputs(110));
    layer0_outputs(2461) <= not((inputs(87)) or (inputs(237)));
    layer0_outputs(2462) <= (inputs(125)) xor (inputs(208));
    layer0_outputs(2463) <= inputs(142);
    layer0_outputs(2464) <= inputs(151);
    layer0_outputs(2465) <= inputs(17);
    layer0_outputs(2466) <= not(inputs(59));
    layer0_outputs(2467) <= not(inputs(123)) or (inputs(72));
    layer0_outputs(2468) <= not(inputs(15)) or (inputs(8));
    layer0_outputs(2469) <= (inputs(197)) and not (inputs(97));
    layer0_outputs(2470) <= not(inputs(74));
    layer0_outputs(2471) <= (inputs(30)) and not (inputs(85));
    layer0_outputs(2472) <= (inputs(96)) or (inputs(114));
    layer0_outputs(2473) <= (inputs(69)) and not (inputs(224));
    layer0_outputs(2474) <= not(inputs(116));
    layer0_outputs(2475) <= (inputs(157)) and (inputs(58));
    layer0_outputs(2476) <= not(inputs(116)) or (inputs(201));
    layer0_outputs(2477) <= '1';
    layer0_outputs(2478) <= not((inputs(12)) or (inputs(19)));
    layer0_outputs(2479) <= (inputs(62)) and not (inputs(15));
    layer0_outputs(2480) <= (inputs(114)) xor (inputs(137));
    layer0_outputs(2481) <= not((inputs(227)) or (inputs(167)));
    layer0_outputs(2482) <= not(inputs(204)) or (inputs(147));
    layer0_outputs(2483) <= not(inputs(53));
    layer0_outputs(2484) <= not(inputs(169)) or (inputs(90));
    layer0_outputs(2485) <= not(inputs(193));
    layer0_outputs(2486) <= not((inputs(224)) or (inputs(145)));
    layer0_outputs(2487) <= not((inputs(126)) or (inputs(33)));
    layer0_outputs(2488) <= not(inputs(234));
    layer0_outputs(2489) <= not(inputs(33));
    layer0_outputs(2490) <= not(inputs(40));
    layer0_outputs(2491) <= (inputs(172)) and (inputs(11));
    layer0_outputs(2492) <= not((inputs(221)) or (inputs(228)));
    layer0_outputs(2493) <= not(inputs(187)) or (inputs(253));
    layer0_outputs(2494) <= (inputs(165)) or (inputs(182));
    layer0_outputs(2495) <= '0';
    layer0_outputs(2496) <= not(inputs(196)) or (inputs(241));
    layer0_outputs(2497) <= (inputs(17)) xor (inputs(9));
    layer0_outputs(2498) <= not(inputs(213)) or (inputs(35));
    layer0_outputs(2499) <= inputs(203);
    layer0_outputs(2500) <= inputs(171);
    layer0_outputs(2501) <= not(inputs(150)) or (inputs(140));
    layer0_outputs(2502) <= not((inputs(173)) or (inputs(255)));
    layer0_outputs(2503) <= inputs(248);
    layer0_outputs(2504) <= (inputs(72)) and not (inputs(207));
    layer0_outputs(2505) <= not((inputs(209)) or (inputs(97)));
    layer0_outputs(2506) <= not(inputs(181));
    layer0_outputs(2507) <= not(inputs(105)) or (inputs(78));
    layer0_outputs(2508) <= not((inputs(184)) or (inputs(200)));
    layer0_outputs(2509) <= (inputs(105)) or (inputs(237));
    layer0_outputs(2510) <= not(inputs(248));
    layer0_outputs(2511) <= not(inputs(35)) or (inputs(221));
    layer0_outputs(2512) <= inputs(116);
    layer0_outputs(2513) <= not(inputs(149)) or (inputs(203));
    layer0_outputs(2514) <= not(inputs(230)) or (inputs(239));
    layer0_outputs(2515) <= not(inputs(107));
    layer0_outputs(2516) <= inputs(63);
    layer0_outputs(2517) <= not(inputs(74));
    layer0_outputs(2518) <= (inputs(3)) xor (inputs(219));
    layer0_outputs(2519) <= not((inputs(202)) or (inputs(246)));
    layer0_outputs(2520) <= not((inputs(178)) or (inputs(212)));
    layer0_outputs(2521) <= (inputs(60)) or (inputs(79));
    layer0_outputs(2522) <= not((inputs(73)) or (inputs(207)));
    layer0_outputs(2523) <= (inputs(67)) and not (inputs(165));
    layer0_outputs(2524) <= not(inputs(14));
    layer0_outputs(2525) <= not((inputs(171)) and (inputs(229)));
    layer0_outputs(2526) <= (inputs(4)) or (inputs(175));
    layer0_outputs(2527) <= not((inputs(187)) or (inputs(248)));
    layer0_outputs(2528) <= '0';
    layer0_outputs(2529) <= (inputs(92)) or (inputs(223));
    layer0_outputs(2530) <= inputs(100);
    layer0_outputs(2531) <= inputs(104);
    layer0_outputs(2532) <= not(inputs(137)) or (inputs(80));
    layer0_outputs(2533) <= (inputs(126)) and not (inputs(75));
    layer0_outputs(2534) <= (inputs(15)) and (inputs(4));
    layer0_outputs(2535) <= inputs(180);
    layer0_outputs(2536) <= not((inputs(144)) or (inputs(194)));
    layer0_outputs(2537) <= not(inputs(24));
    layer0_outputs(2538) <= not(inputs(185));
    layer0_outputs(2539) <= not(inputs(233));
    layer0_outputs(2540) <= (inputs(59)) or (inputs(51));
    layer0_outputs(2541) <= not((inputs(93)) or (inputs(4)));
    layer0_outputs(2542) <= not(inputs(52));
    layer0_outputs(2543) <= inputs(65);
    layer0_outputs(2544) <= not((inputs(104)) or (inputs(133)));
    layer0_outputs(2545) <= (inputs(55)) or (inputs(198));
    layer0_outputs(2546) <= inputs(23);
    layer0_outputs(2547) <= inputs(194);
    layer0_outputs(2548) <= not((inputs(52)) or (inputs(108)));
    layer0_outputs(2549) <= (inputs(88)) or (inputs(216));
    layer0_outputs(2550) <= (inputs(196)) and not (inputs(251));
    layer0_outputs(2551) <= (inputs(143)) xor (inputs(185));
    layer0_outputs(2552) <= (inputs(136)) and not (inputs(175));
    layer0_outputs(2553) <= not(inputs(35)) or (inputs(5));
    layer0_outputs(2554) <= '0';
    layer0_outputs(2555) <= inputs(209);
    layer0_outputs(2556) <= inputs(61);
    layer0_outputs(2557) <= '0';
    layer0_outputs(2558) <= (inputs(184)) and not (inputs(174));
    layer0_outputs(2559) <= not(inputs(250));
    layer0_outputs(2560) <= (inputs(183)) xor (inputs(126));
    layer0_outputs(2561) <= not((inputs(60)) or (inputs(52)));
    layer0_outputs(2562) <= not(inputs(27)) or (inputs(32));
    layer0_outputs(2563) <= not(inputs(53));
    layer0_outputs(2564) <= (inputs(9)) xor (inputs(43));
    layer0_outputs(2565) <= inputs(95);
    layer0_outputs(2566) <= (inputs(70)) xor (inputs(201));
    layer0_outputs(2567) <= (inputs(71)) and not (inputs(100));
    layer0_outputs(2568) <= (inputs(224)) and not (inputs(228));
    layer0_outputs(2569) <= '1';
    layer0_outputs(2570) <= (inputs(76)) and not (inputs(186));
    layer0_outputs(2571) <= not(inputs(54)) or (inputs(0));
    layer0_outputs(2572) <= not((inputs(231)) or (inputs(2)));
    layer0_outputs(2573) <= inputs(113);
    layer0_outputs(2574) <= '1';
    layer0_outputs(2575) <= not(inputs(250));
    layer0_outputs(2576) <= not(inputs(188));
    layer0_outputs(2577) <= not(inputs(214));
    layer0_outputs(2578) <= not((inputs(97)) or (inputs(83)));
    layer0_outputs(2579) <= '0';
    layer0_outputs(2580) <= '1';
    layer0_outputs(2581) <= (inputs(206)) and not (inputs(39));
    layer0_outputs(2582) <= (inputs(109)) or (inputs(114));
    layer0_outputs(2583) <= inputs(218);
    layer0_outputs(2584) <= not((inputs(92)) xor (inputs(111)));
    layer0_outputs(2585) <= (inputs(82)) and not (inputs(16));
    layer0_outputs(2586) <= (inputs(132)) xor (inputs(24));
    layer0_outputs(2587) <= inputs(172);
    layer0_outputs(2588) <= not(inputs(156));
    layer0_outputs(2589) <= not(inputs(164));
    layer0_outputs(2590) <= not(inputs(64));
    layer0_outputs(2591) <= not((inputs(150)) xor (inputs(89)));
    layer0_outputs(2592) <= (inputs(29)) and not (inputs(43));
    layer0_outputs(2593) <= not(inputs(5));
    layer0_outputs(2594) <= not(inputs(96)) or (inputs(249));
    layer0_outputs(2595) <= inputs(135);
    layer0_outputs(2596) <= (inputs(85)) and not (inputs(105));
    layer0_outputs(2597) <= (inputs(106)) xor (inputs(237));
    layer0_outputs(2598) <= (inputs(61)) or (inputs(22));
    layer0_outputs(2599) <= not((inputs(170)) xor (inputs(252)));
    layer0_outputs(2600) <= inputs(71);
    layer0_outputs(2601) <= not(inputs(164)) or (inputs(148));
    layer0_outputs(2602) <= '0';
    layer0_outputs(2603) <= not(inputs(222)) or (inputs(234));
    layer0_outputs(2604) <= not(inputs(102));
    layer0_outputs(2605) <= not(inputs(148));
    layer0_outputs(2606) <= not(inputs(24));
    layer0_outputs(2607) <= not((inputs(183)) or (inputs(212)));
    layer0_outputs(2608) <= (inputs(13)) and not (inputs(115));
    layer0_outputs(2609) <= inputs(188);
    layer0_outputs(2610) <= not(inputs(115));
    layer0_outputs(2611) <= '1';
    layer0_outputs(2612) <= (inputs(240)) and not (inputs(145));
    layer0_outputs(2613) <= '1';
    layer0_outputs(2614) <= not(inputs(66)) or (inputs(55));
    layer0_outputs(2615) <= (inputs(136)) and (inputs(123));
    layer0_outputs(2616) <= (inputs(226)) or (inputs(193));
    layer0_outputs(2617) <= not(inputs(117));
    layer0_outputs(2618) <= not(inputs(158));
    layer0_outputs(2619) <= not(inputs(121)) or (inputs(53));
    layer0_outputs(2620) <= (inputs(122)) xor (inputs(173));
    layer0_outputs(2621) <= '1';
    layer0_outputs(2622) <= inputs(0);
    layer0_outputs(2623) <= inputs(176);
    layer0_outputs(2624) <= not(inputs(90));
    layer0_outputs(2625) <= inputs(152);
    layer0_outputs(2626) <= not((inputs(85)) or (inputs(139)));
    layer0_outputs(2627) <= not(inputs(253));
    layer0_outputs(2628) <= (inputs(80)) or (inputs(4));
    layer0_outputs(2629) <= inputs(47);
    layer0_outputs(2630) <= (inputs(64)) xor (inputs(147));
    layer0_outputs(2631) <= (inputs(57)) xor (inputs(95));
    layer0_outputs(2632) <= (inputs(141)) and not (inputs(11));
    layer0_outputs(2633) <= '0';
    layer0_outputs(2634) <= inputs(146);
    layer0_outputs(2635) <= (inputs(12)) xor (inputs(119));
    layer0_outputs(2636) <= inputs(87);
    layer0_outputs(2637) <= (inputs(55)) and not (inputs(107));
    layer0_outputs(2638) <= not(inputs(217));
    layer0_outputs(2639) <= not((inputs(146)) xor (inputs(181)));
    layer0_outputs(2640) <= inputs(26);
    layer0_outputs(2641) <= '0';
    layer0_outputs(2642) <= '0';
    layer0_outputs(2643) <= not((inputs(89)) or (inputs(151)));
    layer0_outputs(2644) <= (inputs(125)) xor (inputs(123));
    layer0_outputs(2645) <= not((inputs(151)) xor (inputs(140)));
    layer0_outputs(2646) <= (inputs(148)) xor (inputs(102));
    layer0_outputs(2647) <= (inputs(208)) or (inputs(222));
    layer0_outputs(2648) <= (inputs(81)) or (inputs(248));
    layer0_outputs(2649) <= not((inputs(93)) and (inputs(217)));
    layer0_outputs(2650) <= (inputs(50)) and not (inputs(239));
    layer0_outputs(2651) <= (inputs(214)) or (inputs(78));
    layer0_outputs(2652) <= (inputs(171)) or (inputs(188));
    layer0_outputs(2653) <= (inputs(101)) and (inputs(76));
    layer0_outputs(2654) <= inputs(214);
    layer0_outputs(2655) <= (inputs(167)) or (inputs(80));
    layer0_outputs(2656) <= not(inputs(252)) or (inputs(84));
    layer0_outputs(2657) <= not((inputs(78)) or (inputs(208)));
    layer0_outputs(2658) <= not((inputs(202)) or (inputs(38)));
    layer0_outputs(2659) <= not(inputs(56));
    layer0_outputs(2660) <= '0';
    layer0_outputs(2661) <= inputs(71);
    layer0_outputs(2662) <= not(inputs(157));
    layer0_outputs(2663) <= not(inputs(108)) or (inputs(56));
    layer0_outputs(2664) <= not(inputs(219));
    layer0_outputs(2665) <= inputs(111);
    layer0_outputs(2666) <= not((inputs(218)) or (inputs(217)));
    layer0_outputs(2667) <= not(inputs(116));
    layer0_outputs(2668) <= (inputs(39)) and not (inputs(169));
    layer0_outputs(2669) <= not(inputs(147)) or (inputs(248));
    layer0_outputs(2670) <= (inputs(53)) and not (inputs(34));
    layer0_outputs(2671) <= not(inputs(152));
    layer0_outputs(2672) <= not(inputs(163));
    layer0_outputs(2673) <= not(inputs(104)) or (inputs(123));
    layer0_outputs(2674) <= (inputs(189)) and not (inputs(15));
    layer0_outputs(2675) <= not(inputs(123));
    layer0_outputs(2676) <= (inputs(76)) and not (inputs(81));
    layer0_outputs(2677) <= not(inputs(208));
    layer0_outputs(2678) <= inputs(64);
    layer0_outputs(2679) <= inputs(8);
    layer0_outputs(2680) <= inputs(145);
    layer0_outputs(2681) <= (inputs(84)) or (inputs(246));
    layer0_outputs(2682) <= inputs(22);
    layer0_outputs(2683) <= (inputs(250)) or (inputs(102));
    layer0_outputs(2684) <= '1';
    layer0_outputs(2685) <= not(inputs(186));
    layer0_outputs(2686) <= inputs(75);
    layer0_outputs(2687) <= not((inputs(93)) or (inputs(221)));
    layer0_outputs(2688) <= not((inputs(33)) or (inputs(34)));
    layer0_outputs(2689) <= inputs(77);
    layer0_outputs(2690) <= (inputs(188)) or (inputs(203));
    layer0_outputs(2691) <= (inputs(43)) and not (inputs(181));
    layer0_outputs(2692) <= not((inputs(120)) and (inputs(115)));
    layer0_outputs(2693) <= (inputs(195)) or (inputs(15));
    layer0_outputs(2694) <= not(inputs(247)) or (inputs(37));
    layer0_outputs(2695) <= not(inputs(229)) or (inputs(234));
    layer0_outputs(2696) <= (inputs(107)) and not (inputs(197));
    layer0_outputs(2697) <= not((inputs(60)) or (inputs(238)));
    layer0_outputs(2698) <= inputs(182);
    layer0_outputs(2699) <= not(inputs(85)) or (inputs(249));
    layer0_outputs(2700) <= inputs(124);
    layer0_outputs(2701) <= (inputs(116)) or (inputs(60));
    layer0_outputs(2702) <= (inputs(220)) and not (inputs(94));
    layer0_outputs(2703) <= '1';
    layer0_outputs(2704) <= not((inputs(130)) or (inputs(16)));
    layer0_outputs(2705) <= (inputs(170)) and not (inputs(209));
    layer0_outputs(2706) <= (inputs(149)) and not (inputs(13));
    layer0_outputs(2707) <= not(inputs(66));
    layer0_outputs(2708) <= (inputs(29)) xor (inputs(248));
    layer0_outputs(2709) <= (inputs(124)) and not (inputs(222));
    layer0_outputs(2710) <= not(inputs(222));
    layer0_outputs(2711) <= '1';
    layer0_outputs(2712) <= not(inputs(1));
    layer0_outputs(2713) <= (inputs(38)) or (inputs(240));
    layer0_outputs(2714) <= not((inputs(56)) or (inputs(71)));
    layer0_outputs(2715) <= not(inputs(22));
    layer0_outputs(2716) <= inputs(130);
    layer0_outputs(2717) <= inputs(66);
    layer0_outputs(2718) <= not(inputs(116)) or (inputs(23));
    layer0_outputs(2719) <= '0';
    layer0_outputs(2720) <= not(inputs(172)) or (inputs(94));
    layer0_outputs(2721) <= not(inputs(18));
    layer0_outputs(2722) <= not((inputs(218)) xor (inputs(240)));
    layer0_outputs(2723) <= '1';
    layer0_outputs(2724) <= (inputs(21)) and not (inputs(216));
    layer0_outputs(2725) <= inputs(193);
    layer0_outputs(2726) <= (inputs(98)) or (inputs(27));
    layer0_outputs(2727) <= inputs(22);
    layer0_outputs(2728) <= inputs(134);
    layer0_outputs(2729) <= (inputs(63)) and not (inputs(242));
    layer0_outputs(2730) <= (inputs(79)) and not (inputs(169));
    layer0_outputs(2731) <= (inputs(224)) and not (inputs(94));
    layer0_outputs(2732) <= not((inputs(36)) or (inputs(2)));
    layer0_outputs(2733) <= not((inputs(10)) or (inputs(152)));
    layer0_outputs(2734) <= inputs(253);
    layer0_outputs(2735) <= (inputs(110)) or (inputs(204));
    layer0_outputs(2736) <= '0';
    layer0_outputs(2737) <= not(inputs(57)) or (inputs(225));
    layer0_outputs(2738) <= not((inputs(211)) or (inputs(242)));
    layer0_outputs(2739) <= not(inputs(225));
    layer0_outputs(2740) <= not((inputs(28)) or (inputs(34)));
    layer0_outputs(2741) <= (inputs(113)) xor (inputs(103));
    layer0_outputs(2742) <= not(inputs(212));
    layer0_outputs(2743) <= inputs(255);
    layer0_outputs(2744) <= (inputs(55)) and not (inputs(17));
    layer0_outputs(2745) <= not(inputs(232)) or (inputs(93));
    layer0_outputs(2746) <= not(inputs(212)) or (inputs(223));
    layer0_outputs(2747) <= not(inputs(47)) or (inputs(242));
    layer0_outputs(2748) <= (inputs(221)) and not (inputs(67));
    layer0_outputs(2749) <= not((inputs(106)) or (inputs(203)));
    layer0_outputs(2750) <= (inputs(83)) and not (inputs(110));
    layer0_outputs(2751) <= '0';
    layer0_outputs(2752) <= not((inputs(131)) xor (inputs(69)));
    layer0_outputs(2753) <= not(inputs(206));
    layer0_outputs(2754) <= not(inputs(244));
    layer0_outputs(2755) <= (inputs(228)) and not (inputs(14));
    layer0_outputs(2756) <= not((inputs(232)) and (inputs(151)));
    layer0_outputs(2757) <= (inputs(71)) and not (inputs(112));
    layer0_outputs(2758) <= not(inputs(205));
    layer0_outputs(2759) <= not(inputs(12));
    layer0_outputs(2760) <= not(inputs(154));
    layer0_outputs(2761) <= (inputs(251)) and not (inputs(73));
    layer0_outputs(2762) <= (inputs(24)) and (inputs(52));
    layer0_outputs(2763) <= not((inputs(163)) xor (inputs(125)));
    layer0_outputs(2764) <= not(inputs(9));
    layer0_outputs(2765) <= inputs(99);
    layer0_outputs(2766) <= (inputs(17)) xor (inputs(2));
    layer0_outputs(2767) <= (inputs(207)) and not (inputs(14));
    layer0_outputs(2768) <= not(inputs(77));
    layer0_outputs(2769) <= inputs(15);
    layer0_outputs(2770) <= not((inputs(114)) or (inputs(54)));
    layer0_outputs(2771) <= not((inputs(26)) or (inputs(27)));
    layer0_outputs(2772) <= (inputs(83)) and (inputs(83));
    layer0_outputs(2773) <= not((inputs(192)) or (inputs(128)));
    layer0_outputs(2774) <= not(inputs(36));
    layer0_outputs(2775) <= not(inputs(114));
    layer0_outputs(2776) <= (inputs(240)) and (inputs(167));
    layer0_outputs(2777) <= (inputs(230)) or (inputs(47));
    layer0_outputs(2778) <= not((inputs(91)) or (inputs(224)));
    layer0_outputs(2779) <= (inputs(12)) and not (inputs(50));
    layer0_outputs(2780) <= (inputs(85)) xor (inputs(111));
    layer0_outputs(2781) <= inputs(24);
    layer0_outputs(2782) <= not(inputs(159)) or (inputs(215));
    layer0_outputs(2783) <= (inputs(135)) or (inputs(105));
    layer0_outputs(2784) <= not(inputs(206)) or (inputs(250));
    layer0_outputs(2785) <= not(inputs(126)) or (inputs(191));
    layer0_outputs(2786) <= not(inputs(45)) or (inputs(225));
    layer0_outputs(2787) <= not(inputs(122));
    layer0_outputs(2788) <= not(inputs(209));
    layer0_outputs(2789) <= (inputs(30)) xor (inputs(112));
    layer0_outputs(2790) <= inputs(51);
    layer0_outputs(2791) <= (inputs(159)) or (inputs(128));
    layer0_outputs(2792) <= (inputs(147)) or (inputs(236));
    layer0_outputs(2793) <= '1';
    layer0_outputs(2794) <= inputs(18);
    layer0_outputs(2795) <= not((inputs(95)) or (inputs(29)));
    layer0_outputs(2796) <= (inputs(77)) or (inputs(123));
    layer0_outputs(2797) <= '0';
    layer0_outputs(2798) <= inputs(190);
    layer0_outputs(2799) <= (inputs(161)) xor (inputs(230));
    layer0_outputs(2800) <= (inputs(58)) xor (inputs(138));
    layer0_outputs(2801) <= (inputs(99)) xor (inputs(71));
    layer0_outputs(2802) <= (inputs(14)) and not (inputs(220));
    layer0_outputs(2803) <= not((inputs(68)) xor (inputs(159)));
    layer0_outputs(2804) <= (inputs(210)) and (inputs(240));
    layer0_outputs(2805) <= (inputs(95)) xor (inputs(41));
    layer0_outputs(2806) <= inputs(164);
    layer0_outputs(2807) <= not((inputs(22)) or (inputs(95)));
    layer0_outputs(2808) <= '0';
    layer0_outputs(2809) <= inputs(57);
    layer0_outputs(2810) <= not(inputs(197)) or (inputs(47));
    layer0_outputs(2811) <= not(inputs(119)) or (inputs(216));
    layer0_outputs(2812) <= '0';
    layer0_outputs(2813) <= inputs(17);
    layer0_outputs(2814) <= '0';
    layer0_outputs(2815) <= not(inputs(133)) or (inputs(222));
    layer0_outputs(2816) <= (inputs(203)) xor (inputs(79));
    layer0_outputs(2817) <= inputs(147);
    layer0_outputs(2818) <= (inputs(90)) and not (inputs(233));
    layer0_outputs(2819) <= (inputs(189)) or (inputs(209));
    layer0_outputs(2820) <= (inputs(237)) and not (inputs(88));
    layer0_outputs(2821) <= not((inputs(216)) and (inputs(203)));
    layer0_outputs(2822) <= not((inputs(253)) and (inputs(44)));
    layer0_outputs(2823) <= not((inputs(77)) xor (inputs(29)));
    layer0_outputs(2824) <= inputs(55);
    layer0_outputs(2825) <= not(inputs(103));
    layer0_outputs(2826) <= not(inputs(84));
    layer0_outputs(2827) <= (inputs(106)) or (inputs(101));
    layer0_outputs(2828) <= inputs(209);
    layer0_outputs(2829) <= inputs(153);
    layer0_outputs(2830) <= inputs(128);
    layer0_outputs(2831) <= inputs(31);
    layer0_outputs(2832) <= not((inputs(174)) and (inputs(59)));
    layer0_outputs(2833) <= not((inputs(70)) or (inputs(147)));
    layer0_outputs(2834) <= not((inputs(72)) or (inputs(253)));
    layer0_outputs(2835) <= inputs(151);
    layer0_outputs(2836) <= not(inputs(0));
    layer0_outputs(2837) <= not(inputs(161));
    layer0_outputs(2838) <= not(inputs(104));
    layer0_outputs(2839) <= not(inputs(148));
    layer0_outputs(2840) <= not(inputs(97));
    layer0_outputs(2841) <= not(inputs(225)) or (inputs(67));
    layer0_outputs(2842) <= not(inputs(202));
    layer0_outputs(2843) <= not(inputs(207)) or (inputs(242));
    layer0_outputs(2844) <= (inputs(60)) or (inputs(123));
    layer0_outputs(2845) <= not(inputs(180));
    layer0_outputs(2846) <= not(inputs(7)) or (inputs(161));
    layer0_outputs(2847) <= not(inputs(178));
    layer0_outputs(2848) <= (inputs(143)) or (inputs(4));
    layer0_outputs(2849) <= (inputs(136)) and not (inputs(3));
    layer0_outputs(2850) <= not((inputs(1)) xor (inputs(54)));
    layer0_outputs(2851) <= inputs(166);
    layer0_outputs(2852) <= not((inputs(128)) xor (inputs(146)));
    layer0_outputs(2853) <= (inputs(40)) and not (inputs(149));
    layer0_outputs(2854) <= (inputs(29)) xor (inputs(88));
    layer0_outputs(2855) <= not((inputs(116)) or (inputs(223)));
    layer0_outputs(2856) <= not(inputs(183));
    layer0_outputs(2857) <= not(inputs(69));
    layer0_outputs(2858) <= not((inputs(84)) xor (inputs(164)));
    layer0_outputs(2859) <= not(inputs(163));
    layer0_outputs(2860) <= (inputs(130)) or (inputs(199));
    layer0_outputs(2861) <= not((inputs(62)) or (inputs(134)));
    layer0_outputs(2862) <= inputs(169);
    layer0_outputs(2863) <= (inputs(27)) or (inputs(172));
    layer0_outputs(2864) <= (inputs(54)) or (inputs(13));
    layer0_outputs(2865) <= (inputs(202)) or (inputs(176));
    layer0_outputs(2866) <= not((inputs(172)) or (inputs(203)));
    layer0_outputs(2867) <= not(inputs(99));
    layer0_outputs(2868) <= inputs(10);
    layer0_outputs(2869) <= inputs(161);
    layer0_outputs(2870) <= (inputs(34)) or (inputs(6));
    layer0_outputs(2871) <= not((inputs(63)) xor (inputs(19)));
    layer0_outputs(2872) <= not((inputs(57)) or (inputs(160)));
    layer0_outputs(2873) <= not(inputs(148));
    layer0_outputs(2874) <= not(inputs(28));
    layer0_outputs(2875) <= (inputs(147)) or (inputs(209));
    layer0_outputs(2876) <= inputs(165);
    layer0_outputs(2877) <= not(inputs(96));
    layer0_outputs(2878) <= '1';
    layer0_outputs(2879) <= (inputs(162)) or (inputs(198));
    layer0_outputs(2880) <= inputs(240);
    layer0_outputs(2881) <= (inputs(167)) xor (inputs(129));
    layer0_outputs(2882) <= inputs(128);
    layer0_outputs(2883) <= not((inputs(150)) or (inputs(198)));
    layer0_outputs(2884) <= (inputs(45)) and not (inputs(254));
    layer0_outputs(2885) <= not((inputs(42)) xor (inputs(15)));
    layer0_outputs(2886) <= (inputs(5)) and not (inputs(158));
    layer0_outputs(2887) <= (inputs(100)) xor (inputs(69));
    layer0_outputs(2888) <= inputs(5);
    layer0_outputs(2889) <= (inputs(159)) and (inputs(129));
    layer0_outputs(2890) <= not(inputs(136)) or (inputs(185));
    layer0_outputs(2891) <= not((inputs(143)) xor (inputs(152)));
    layer0_outputs(2892) <= (inputs(129)) and not (inputs(254));
    layer0_outputs(2893) <= (inputs(25)) and not (inputs(178));
    layer0_outputs(2894) <= not((inputs(2)) and (inputs(162)));
    layer0_outputs(2895) <= not(inputs(73));
    layer0_outputs(2896) <= not(inputs(114));
    layer0_outputs(2897) <= not((inputs(139)) xor (inputs(141)));
    layer0_outputs(2898) <= inputs(27);
    layer0_outputs(2899) <= (inputs(97)) xor (inputs(187));
    layer0_outputs(2900) <= (inputs(223)) and (inputs(213));
    layer0_outputs(2901) <= (inputs(9)) and not (inputs(190));
    layer0_outputs(2902) <= not(inputs(221));
    layer0_outputs(2903) <= not(inputs(13));
    layer0_outputs(2904) <= not((inputs(159)) and (inputs(179)));
    layer0_outputs(2905) <= not(inputs(178));
    layer0_outputs(2906) <= not((inputs(26)) or (inputs(226)));
    layer0_outputs(2907) <= not(inputs(14));
    layer0_outputs(2908) <= not((inputs(27)) or (inputs(132)));
    layer0_outputs(2909) <= '0';
    layer0_outputs(2910) <= not(inputs(90)) or (inputs(112));
    layer0_outputs(2911) <= not(inputs(34));
    layer0_outputs(2912) <= inputs(151);
    layer0_outputs(2913) <= inputs(191);
    layer0_outputs(2914) <= not(inputs(214)) or (inputs(173));
    layer0_outputs(2915) <= '0';
    layer0_outputs(2916) <= not((inputs(134)) xor (inputs(248)));
    layer0_outputs(2917) <= (inputs(147)) and not (inputs(63));
    layer0_outputs(2918) <= not((inputs(83)) xor (inputs(0)));
    layer0_outputs(2919) <= inputs(211);
    layer0_outputs(2920) <= (inputs(23)) and (inputs(26));
    layer0_outputs(2921) <= (inputs(194)) or (inputs(221));
    layer0_outputs(2922) <= not((inputs(96)) or (inputs(70)));
    layer0_outputs(2923) <= not(inputs(86));
    layer0_outputs(2924) <= inputs(195);
    layer0_outputs(2925) <= not((inputs(198)) xor (inputs(77)));
    layer0_outputs(2926) <= inputs(150);
    layer0_outputs(2927) <= not(inputs(201));
    layer0_outputs(2928) <= not((inputs(249)) and (inputs(244)));
    layer0_outputs(2929) <= not(inputs(183)) or (inputs(216));
    layer0_outputs(2930) <= inputs(236);
    layer0_outputs(2931) <= (inputs(230)) and not (inputs(35));
    layer0_outputs(2932) <= not(inputs(135));
    layer0_outputs(2933) <= not((inputs(159)) and (inputs(243)));
    layer0_outputs(2934) <= not((inputs(223)) or (inputs(152)));
    layer0_outputs(2935) <= (inputs(178)) xor (inputs(180));
    layer0_outputs(2936) <= not(inputs(170)) or (inputs(85));
    layer0_outputs(2937) <= not((inputs(55)) xor (inputs(55)));
    layer0_outputs(2938) <= (inputs(234)) xor (inputs(86));
    layer0_outputs(2939) <= inputs(211);
    layer0_outputs(2940) <= (inputs(27)) and not (inputs(140));
    layer0_outputs(2941) <= (inputs(173)) and not (inputs(3));
    layer0_outputs(2942) <= (inputs(22)) and (inputs(41));
    layer0_outputs(2943) <= (inputs(10)) and not (inputs(246));
    layer0_outputs(2944) <= not((inputs(49)) or (inputs(29)));
    layer0_outputs(2945) <= inputs(220);
    layer0_outputs(2946) <= (inputs(221)) and not (inputs(177));
    layer0_outputs(2947) <= (inputs(212)) or (inputs(127));
    layer0_outputs(2948) <= (inputs(206)) or (inputs(217));
    layer0_outputs(2949) <= not(inputs(72));
    layer0_outputs(2950) <= (inputs(54)) or (inputs(101));
    layer0_outputs(2951) <= inputs(75);
    layer0_outputs(2952) <= (inputs(221)) and not (inputs(41));
    layer0_outputs(2953) <= not((inputs(233)) or (inputs(200)));
    layer0_outputs(2954) <= inputs(192);
    layer0_outputs(2955) <= not((inputs(193)) or (inputs(133)));
    layer0_outputs(2956) <= inputs(207);
    layer0_outputs(2957) <= (inputs(61)) or (inputs(181));
    layer0_outputs(2958) <= not(inputs(48));
    layer0_outputs(2959) <= (inputs(245)) or (inputs(177));
    layer0_outputs(2960) <= not((inputs(251)) xor (inputs(164)));
    layer0_outputs(2961) <= (inputs(148)) xor (inputs(3));
    layer0_outputs(2962) <= inputs(4);
    layer0_outputs(2963) <= (inputs(70)) and (inputs(127));
    layer0_outputs(2964) <= inputs(169);
    layer0_outputs(2965) <= inputs(71);
    layer0_outputs(2966) <= (inputs(206)) or (inputs(238));
    layer0_outputs(2967) <= not((inputs(53)) xor (inputs(221)));
    layer0_outputs(2968) <= not((inputs(90)) xor (inputs(162)));
    layer0_outputs(2969) <= inputs(90);
    layer0_outputs(2970) <= not(inputs(137));
    layer0_outputs(2971) <= '0';
    layer0_outputs(2972) <= not(inputs(196));
    layer0_outputs(2973) <= not(inputs(106)) or (inputs(46));
    layer0_outputs(2974) <= (inputs(176)) or (inputs(233));
    layer0_outputs(2975) <= (inputs(109)) or (inputs(95));
    layer0_outputs(2976) <= not((inputs(225)) or (inputs(242)));
    layer0_outputs(2977) <= not((inputs(82)) or (inputs(215)));
    layer0_outputs(2978) <= inputs(31);
    layer0_outputs(2979) <= not(inputs(72));
    layer0_outputs(2980) <= not((inputs(19)) and (inputs(46)));
    layer0_outputs(2981) <= (inputs(235)) xor (inputs(116));
    layer0_outputs(2982) <= inputs(109);
    layer0_outputs(2983) <= (inputs(191)) or (inputs(49));
    layer0_outputs(2984) <= not((inputs(227)) or (inputs(209)));
    layer0_outputs(2985) <= not(inputs(151)) or (inputs(210));
    layer0_outputs(2986) <= not(inputs(73)) or (inputs(55));
    layer0_outputs(2987) <= not((inputs(222)) xor (inputs(60)));
    layer0_outputs(2988) <= (inputs(37)) and not (inputs(18));
    layer0_outputs(2989) <= '0';
    layer0_outputs(2990) <= not(inputs(71));
    layer0_outputs(2991) <= not(inputs(130));
    layer0_outputs(2992) <= (inputs(81)) xor (inputs(147));
    layer0_outputs(2993) <= not(inputs(211));
    layer0_outputs(2994) <= not((inputs(101)) xor (inputs(112)));
    layer0_outputs(2995) <= not((inputs(224)) or (inputs(31)));
    layer0_outputs(2996) <= '0';
    layer0_outputs(2997) <= inputs(87);
    layer0_outputs(2998) <= (inputs(104)) and (inputs(188));
    layer0_outputs(2999) <= not(inputs(0));
    layer0_outputs(3000) <= inputs(62);
    layer0_outputs(3001) <= not((inputs(62)) xor (inputs(17)));
    layer0_outputs(3002) <= not(inputs(99)) or (inputs(3));
    layer0_outputs(3003) <= (inputs(188)) and not (inputs(102));
    layer0_outputs(3004) <= (inputs(50)) and not (inputs(122));
    layer0_outputs(3005) <= (inputs(63)) and not (inputs(161));
    layer0_outputs(3006) <= inputs(197);
    layer0_outputs(3007) <= not((inputs(162)) or (inputs(52)));
    layer0_outputs(3008) <= not((inputs(3)) or (inputs(189)));
    layer0_outputs(3009) <= (inputs(81)) or (inputs(139));
    layer0_outputs(3010) <= not((inputs(230)) or (inputs(113)));
    layer0_outputs(3011) <= not(inputs(176)) or (inputs(250));
    layer0_outputs(3012) <= not((inputs(188)) and (inputs(179)));
    layer0_outputs(3013) <= '0';
    layer0_outputs(3014) <= (inputs(194)) and not (inputs(18));
    layer0_outputs(3015) <= not(inputs(105)) or (inputs(145));
    layer0_outputs(3016) <= '0';
    layer0_outputs(3017) <= inputs(223);
    layer0_outputs(3018) <= '0';
    layer0_outputs(3019) <= (inputs(195)) xor (inputs(244));
    layer0_outputs(3020) <= '0';
    layer0_outputs(3021) <= (inputs(6)) or (inputs(210));
    layer0_outputs(3022) <= inputs(158);
    layer0_outputs(3023) <= inputs(129);
    layer0_outputs(3024) <= not((inputs(95)) xor (inputs(167)));
    layer0_outputs(3025) <= inputs(78);
    layer0_outputs(3026) <= inputs(217);
    layer0_outputs(3027) <= '1';
    layer0_outputs(3028) <= not(inputs(97));
    layer0_outputs(3029) <= not(inputs(99));
    layer0_outputs(3030) <= not((inputs(177)) xor (inputs(198)));
    layer0_outputs(3031) <= (inputs(50)) or (inputs(248));
    layer0_outputs(3032) <= (inputs(28)) or (inputs(34));
    layer0_outputs(3033) <= (inputs(49)) xor (inputs(139));
    layer0_outputs(3034) <= not((inputs(59)) xor (inputs(172)));
    layer0_outputs(3035) <= (inputs(107)) and not (inputs(82));
    layer0_outputs(3036) <= '0';
    layer0_outputs(3037) <= (inputs(71)) and not (inputs(22));
    layer0_outputs(3038) <= not((inputs(31)) or (inputs(219)));
    layer0_outputs(3039) <= (inputs(53)) xor (inputs(132));
    layer0_outputs(3040) <= (inputs(238)) or (inputs(88));
    layer0_outputs(3041) <= not(inputs(34));
    layer0_outputs(3042) <= not(inputs(109));
    layer0_outputs(3043) <= '0';
    layer0_outputs(3044) <= inputs(115);
    layer0_outputs(3045) <= not(inputs(81)) or (inputs(170));
    layer0_outputs(3046) <= not(inputs(24)) or (inputs(118));
    layer0_outputs(3047) <= inputs(136);
    layer0_outputs(3048) <= (inputs(77)) xor (inputs(237));
    layer0_outputs(3049) <= inputs(157);
    layer0_outputs(3050) <= (inputs(119)) and not (inputs(31));
    layer0_outputs(3051) <= inputs(229);
    layer0_outputs(3052) <= not((inputs(236)) and (inputs(25)));
    layer0_outputs(3053) <= inputs(36);
    layer0_outputs(3054) <= not((inputs(238)) or (inputs(99)));
    layer0_outputs(3055) <= (inputs(234)) and (inputs(11));
    layer0_outputs(3056) <= (inputs(40)) and (inputs(250));
    layer0_outputs(3057) <= not(inputs(219));
    layer0_outputs(3058) <= not(inputs(168));
    layer0_outputs(3059) <= not(inputs(60)) or (inputs(164));
    layer0_outputs(3060) <= not((inputs(254)) or (inputs(179)));
    layer0_outputs(3061) <= not(inputs(123)) or (inputs(161));
    layer0_outputs(3062) <= not((inputs(184)) or (inputs(185)));
    layer0_outputs(3063) <= not(inputs(235)) or (inputs(112));
    layer0_outputs(3064) <= not((inputs(204)) or (inputs(120)));
    layer0_outputs(3065) <= not((inputs(41)) or (inputs(49)));
    layer0_outputs(3066) <= not((inputs(134)) xor (inputs(114)));
    layer0_outputs(3067) <= inputs(182);
    layer0_outputs(3068) <= not((inputs(229)) or (inputs(177)));
    layer0_outputs(3069) <= (inputs(58)) and not (inputs(178));
    layer0_outputs(3070) <= (inputs(50)) or (inputs(89));
    layer0_outputs(3071) <= not(inputs(101));
    layer0_outputs(3072) <= (inputs(248)) and not (inputs(121));
    layer0_outputs(3073) <= '0';
    layer0_outputs(3074) <= not((inputs(92)) or (inputs(60)));
    layer0_outputs(3075) <= (inputs(170)) xor (inputs(67));
    layer0_outputs(3076) <= (inputs(142)) xor (inputs(198));
    layer0_outputs(3077) <= '0';
    layer0_outputs(3078) <= not((inputs(49)) and (inputs(230)));
    layer0_outputs(3079) <= not(inputs(219));
    layer0_outputs(3080) <= inputs(58);
    layer0_outputs(3081) <= inputs(241);
    layer0_outputs(3082) <= inputs(35);
    layer0_outputs(3083) <= inputs(222);
    layer0_outputs(3084) <= inputs(75);
    layer0_outputs(3085) <= not(inputs(100)) or (inputs(109));
    layer0_outputs(3086) <= not((inputs(29)) or (inputs(131)));
    layer0_outputs(3087) <= not((inputs(201)) or (inputs(188)));
    layer0_outputs(3088) <= not((inputs(180)) or (inputs(153)));
    layer0_outputs(3089) <= inputs(185);
    layer0_outputs(3090) <= inputs(67);
    layer0_outputs(3091) <= (inputs(34)) and not (inputs(11));
    layer0_outputs(3092) <= (inputs(137)) and not (inputs(32));
    layer0_outputs(3093) <= not((inputs(227)) or (inputs(34)));
    layer0_outputs(3094) <= (inputs(12)) or (inputs(115));
    layer0_outputs(3095) <= not((inputs(139)) xor (inputs(175)));
    layer0_outputs(3096) <= (inputs(20)) xor (inputs(169));
    layer0_outputs(3097) <= not(inputs(23)) or (inputs(143));
    layer0_outputs(3098) <= inputs(87);
    layer0_outputs(3099) <= not((inputs(50)) and (inputs(184)));
    layer0_outputs(3100) <= not(inputs(172));
    layer0_outputs(3101) <= (inputs(30)) and not (inputs(155));
    layer0_outputs(3102) <= (inputs(187)) or (inputs(13));
    layer0_outputs(3103) <= not((inputs(243)) or (inputs(134)));
    layer0_outputs(3104) <= (inputs(255)) and not (inputs(251));
    layer0_outputs(3105) <= not(inputs(138));
    layer0_outputs(3106) <= (inputs(224)) and not (inputs(131));
    layer0_outputs(3107) <= inputs(46);
    layer0_outputs(3108) <= inputs(24);
    layer0_outputs(3109) <= not(inputs(104));
    layer0_outputs(3110) <= not(inputs(189)) or (inputs(228));
    layer0_outputs(3111) <= not((inputs(163)) xor (inputs(182)));
    layer0_outputs(3112) <= not(inputs(64)) or (inputs(43));
    layer0_outputs(3113) <= not(inputs(66)) or (inputs(157));
    layer0_outputs(3114) <= inputs(24);
    layer0_outputs(3115) <= not(inputs(91)) or (inputs(214));
    layer0_outputs(3116) <= (inputs(232)) and not (inputs(56));
    layer0_outputs(3117) <= inputs(94);
    layer0_outputs(3118) <= not((inputs(21)) xor (inputs(45)));
    layer0_outputs(3119) <= not((inputs(182)) or (inputs(35)));
    layer0_outputs(3120) <= (inputs(34)) or (inputs(9));
    layer0_outputs(3121) <= not(inputs(119));
    layer0_outputs(3122) <= inputs(211);
    layer0_outputs(3123) <= not(inputs(30)) or (inputs(127));
    layer0_outputs(3124) <= '0';
    layer0_outputs(3125) <= (inputs(228)) or (inputs(194));
    layer0_outputs(3126) <= (inputs(218)) and not (inputs(115));
    layer0_outputs(3127) <= inputs(62);
    layer0_outputs(3128) <= '1';
    layer0_outputs(3129) <= inputs(40);
    layer0_outputs(3130) <= inputs(119);
    layer0_outputs(3131) <= not(inputs(43));
    layer0_outputs(3132) <= (inputs(118)) or (inputs(211));
    layer0_outputs(3133) <= not((inputs(155)) or (inputs(255)));
    layer0_outputs(3134) <= inputs(73);
    layer0_outputs(3135) <= not(inputs(209));
    layer0_outputs(3136) <= not((inputs(6)) or (inputs(192)));
    layer0_outputs(3137) <= (inputs(57)) and not (inputs(50));
    layer0_outputs(3138) <= not(inputs(72));
    layer0_outputs(3139) <= not(inputs(57));
    layer0_outputs(3140) <= not((inputs(146)) or (inputs(95)));
    layer0_outputs(3141) <= (inputs(221)) and (inputs(123));
    layer0_outputs(3142) <= not((inputs(210)) or (inputs(144)));
    layer0_outputs(3143) <= inputs(69);
    layer0_outputs(3144) <= (inputs(78)) or (inputs(223));
    layer0_outputs(3145) <= not((inputs(51)) xor (inputs(46)));
    layer0_outputs(3146) <= inputs(115);
    layer0_outputs(3147) <= inputs(166);
    layer0_outputs(3148) <= not(inputs(91)) or (inputs(146));
    layer0_outputs(3149) <= (inputs(26)) and not (inputs(252));
    layer0_outputs(3150) <= not((inputs(18)) or (inputs(118)));
    layer0_outputs(3151) <= inputs(148);
    layer0_outputs(3152) <= not((inputs(23)) xor (inputs(124)));
    layer0_outputs(3153) <= not(inputs(30));
    layer0_outputs(3154) <= '0';
    layer0_outputs(3155) <= not(inputs(129)) or (inputs(220));
    layer0_outputs(3156) <= not(inputs(45)) or (inputs(173));
    layer0_outputs(3157) <= not((inputs(132)) xor (inputs(255)));
    layer0_outputs(3158) <= (inputs(220)) and not (inputs(1));
    layer0_outputs(3159) <= not(inputs(98));
    layer0_outputs(3160) <= not(inputs(12));
    layer0_outputs(3161) <= (inputs(180)) xor (inputs(25));
    layer0_outputs(3162) <= not((inputs(129)) or (inputs(99)));
    layer0_outputs(3163) <= (inputs(76)) or (inputs(141));
    layer0_outputs(3164) <= (inputs(14)) or (inputs(120));
    layer0_outputs(3165) <= not((inputs(163)) or (inputs(85)));
    layer0_outputs(3166) <= not(inputs(235)) or (inputs(47));
    layer0_outputs(3167) <= inputs(208);
    layer0_outputs(3168) <= (inputs(35)) and not (inputs(251));
    layer0_outputs(3169) <= not((inputs(142)) and (inputs(120)));
    layer0_outputs(3170) <= inputs(103);
    layer0_outputs(3171) <= not(inputs(165));
    layer0_outputs(3172) <= inputs(86);
    layer0_outputs(3173) <= (inputs(35)) or (inputs(174));
    layer0_outputs(3174) <= not((inputs(253)) and (inputs(5)));
    layer0_outputs(3175) <= inputs(216);
    layer0_outputs(3176) <= (inputs(40)) and not (inputs(108));
    layer0_outputs(3177) <= (inputs(220)) or (inputs(175));
    layer0_outputs(3178) <= (inputs(34)) and not (inputs(128));
    layer0_outputs(3179) <= not(inputs(215)) or (inputs(60));
    layer0_outputs(3180) <= (inputs(96)) or (inputs(98));
    layer0_outputs(3181) <= not(inputs(221)) or (inputs(7));
    layer0_outputs(3182) <= '0';
    layer0_outputs(3183) <= (inputs(57)) and (inputs(212));
    layer0_outputs(3184) <= inputs(88);
    layer0_outputs(3185) <= (inputs(52)) and not (inputs(134));
    layer0_outputs(3186) <= not(inputs(149));
    layer0_outputs(3187) <= (inputs(248)) or (inputs(231));
    layer0_outputs(3188) <= not((inputs(148)) and (inputs(142)));
    layer0_outputs(3189) <= not((inputs(203)) or (inputs(4)));
    layer0_outputs(3190) <= not((inputs(164)) and (inputs(140)));
    layer0_outputs(3191) <= '1';
    layer0_outputs(3192) <= not(inputs(204));
    layer0_outputs(3193) <= (inputs(8)) and not (inputs(14));
    layer0_outputs(3194) <= (inputs(102)) and not (inputs(131));
    layer0_outputs(3195) <= not(inputs(37));
    layer0_outputs(3196) <= (inputs(240)) xor (inputs(118));
    layer0_outputs(3197) <= not((inputs(50)) xor (inputs(60)));
    layer0_outputs(3198) <= not((inputs(73)) xor (inputs(171)));
    layer0_outputs(3199) <= not(inputs(172)) or (inputs(147));
    layer0_outputs(3200) <= inputs(45);
    layer0_outputs(3201) <= (inputs(81)) and not (inputs(190));
    layer0_outputs(3202) <= not((inputs(195)) or (inputs(225)));
    layer0_outputs(3203) <= not((inputs(149)) or (inputs(134)));
    layer0_outputs(3204) <= not((inputs(177)) or (inputs(83)));
    layer0_outputs(3205) <= not(inputs(98)) or (inputs(111));
    layer0_outputs(3206) <= not(inputs(102));
    layer0_outputs(3207) <= (inputs(248)) and (inputs(111));
    layer0_outputs(3208) <= not(inputs(9));
    layer0_outputs(3209) <= not((inputs(204)) or (inputs(235)));
    layer0_outputs(3210) <= not((inputs(97)) xor (inputs(145)));
    layer0_outputs(3211) <= not((inputs(236)) or (inputs(32)));
    layer0_outputs(3212) <= (inputs(22)) xor (inputs(48));
    layer0_outputs(3213) <= (inputs(32)) xor (inputs(70));
    layer0_outputs(3214) <= inputs(151);
    layer0_outputs(3215) <= not(inputs(212));
    layer0_outputs(3216) <= (inputs(42)) and not (inputs(103));
    layer0_outputs(3217) <= not((inputs(68)) xor (inputs(35)));
    layer0_outputs(3218) <= not(inputs(192));
    layer0_outputs(3219) <= (inputs(58)) and not (inputs(48));
    layer0_outputs(3220) <= not(inputs(124)) or (inputs(157));
    layer0_outputs(3221) <= not((inputs(105)) xor (inputs(171)));
    layer0_outputs(3222) <= inputs(129);
    layer0_outputs(3223) <= (inputs(151)) or (inputs(239));
    layer0_outputs(3224) <= not(inputs(117));
    layer0_outputs(3225) <= (inputs(245)) and not (inputs(14));
    layer0_outputs(3226) <= not(inputs(222)) or (inputs(36));
    layer0_outputs(3227) <= not(inputs(93));
    layer0_outputs(3228) <= (inputs(251)) xor (inputs(151));
    layer0_outputs(3229) <= (inputs(130)) or (inputs(152));
    layer0_outputs(3230) <= not((inputs(157)) xor (inputs(109)));
    layer0_outputs(3231) <= (inputs(146)) xor (inputs(229));
    layer0_outputs(3232) <= (inputs(236)) xor (inputs(17));
    layer0_outputs(3233) <= (inputs(251)) or (inputs(153));
    layer0_outputs(3234) <= not(inputs(131)) or (inputs(73));
    layer0_outputs(3235) <= (inputs(112)) and (inputs(196));
    layer0_outputs(3236) <= (inputs(130)) or (inputs(134));
    layer0_outputs(3237) <= not(inputs(249));
    layer0_outputs(3238) <= not(inputs(85));
    layer0_outputs(3239) <= (inputs(186)) and not (inputs(98));
    layer0_outputs(3240) <= '1';
    layer0_outputs(3241) <= (inputs(90)) and not (inputs(238));
    layer0_outputs(3242) <= (inputs(206)) xor (inputs(107));
    layer0_outputs(3243) <= inputs(229);
    layer0_outputs(3244) <= not(inputs(202));
    layer0_outputs(3245) <= not((inputs(26)) xor (inputs(159)));
    layer0_outputs(3246) <= not(inputs(156));
    layer0_outputs(3247) <= not((inputs(15)) or (inputs(254)));
    layer0_outputs(3248) <= (inputs(203)) xor (inputs(140));
    layer0_outputs(3249) <= not(inputs(93));
    layer0_outputs(3250) <= (inputs(146)) or (inputs(110));
    layer0_outputs(3251) <= (inputs(237)) xor (inputs(207));
    layer0_outputs(3252) <= not(inputs(224));
    layer0_outputs(3253) <= inputs(120);
    layer0_outputs(3254) <= not((inputs(229)) or (inputs(244)));
    layer0_outputs(3255) <= '1';
    layer0_outputs(3256) <= not(inputs(58));
    layer0_outputs(3257) <= (inputs(36)) xor (inputs(210));
    layer0_outputs(3258) <= (inputs(199)) and not (inputs(135));
    layer0_outputs(3259) <= not(inputs(188)) or (inputs(112));
    layer0_outputs(3260) <= (inputs(100)) or (inputs(253));
    layer0_outputs(3261) <= not((inputs(10)) or (inputs(4)));
    layer0_outputs(3262) <= (inputs(235)) and not (inputs(119));
    layer0_outputs(3263) <= (inputs(137)) and not (inputs(54));
    layer0_outputs(3264) <= not(inputs(10));
    layer0_outputs(3265) <= (inputs(39)) or (inputs(97));
    layer0_outputs(3266) <= not((inputs(109)) and (inputs(194)));
    layer0_outputs(3267) <= inputs(228);
    layer0_outputs(3268) <= not(inputs(112)) or (inputs(127));
    layer0_outputs(3269) <= not(inputs(18)) or (inputs(13));
    layer0_outputs(3270) <= inputs(73);
    layer0_outputs(3271) <= not(inputs(166));
    layer0_outputs(3272) <= not((inputs(147)) xor (inputs(97)));
    layer0_outputs(3273) <= not((inputs(114)) or (inputs(148)));
    layer0_outputs(3274) <= inputs(175);
    layer0_outputs(3275) <= (inputs(176)) or (inputs(99));
    layer0_outputs(3276) <= not(inputs(90));
    layer0_outputs(3277) <= not((inputs(182)) and (inputs(18)));
    layer0_outputs(3278) <= inputs(121);
    layer0_outputs(3279) <= (inputs(145)) and not (inputs(59));
    layer0_outputs(3280) <= '1';
    layer0_outputs(3281) <= not((inputs(4)) xor (inputs(16)));
    layer0_outputs(3282) <= not(inputs(137));
    layer0_outputs(3283) <= (inputs(40)) and not (inputs(129));
    layer0_outputs(3284) <= not(inputs(164));
    layer0_outputs(3285) <= (inputs(40)) or (inputs(20));
    layer0_outputs(3286) <= inputs(199);
    layer0_outputs(3287) <= inputs(250);
    layer0_outputs(3288) <= (inputs(110)) and (inputs(63));
    layer0_outputs(3289) <= not(inputs(8));
    layer0_outputs(3290) <= (inputs(156)) and (inputs(217));
    layer0_outputs(3291) <= (inputs(143)) or (inputs(231));
    layer0_outputs(3292) <= inputs(158);
    layer0_outputs(3293) <= not(inputs(173));
    layer0_outputs(3294) <= (inputs(226)) or (inputs(223));
    layer0_outputs(3295) <= (inputs(201)) xor (inputs(233));
    layer0_outputs(3296) <= not((inputs(172)) and (inputs(245)));
    layer0_outputs(3297) <= not(inputs(11));
    layer0_outputs(3298) <= inputs(217);
    layer0_outputs(3299) <= not(inputs(42));
    layer0_outputs(3300) <= not(inputs(76));
    layer0_outputs(3301) <= (inputs(248)) and not (inputs(106));
    layer0_outputs(3302) <= (inputs(1)) and (inputs(82));
    layer0_outputs(3303) <= not(inputs(100));
    layer0_outputs(3304) <= not(inputs(72)) or (inputs(82));
    layer0_outputs(3305) <= not((inputs(221)) and (inputs(221)));
    layer0_outputs(3306) <= not(inputs(217));
    layer0_outputs(3307) <= not((inputs(242)) or (inputs(127)));
    layer0_outputs(3308) <= (inputs(248)) and not (inputs(75));
    layer0_outputs(3309) <= inputs(232);
    layer0_outputs(3310) <= (inputs(242)) and not (inputs(98));
    layer0_outputs(3311) <= not((inputs(116)) or (inputs(254)));
    layer0_outputs(3312) <= (inputs(29)) and (inputs(145));
    layer0_outputs(3313) <= (inputs(128)) xor (inputs(164));
    layer0_outputs(3314) <= not(inputs(43)) or (inputs(239));
    layer0_outputs(3315) <= inputs(65);
    layer0_outputs(3316) <= not(inputs(166)) or (inputs(62));
    layer0_outputs(3317) <= (inputs(170)) and not (inputs(226));
    layer0_outputs(3318) <= not(inputs(20)) or (inputs(192));
    layer0_outputs(3319) <= not((inputs(1)) or (inputs(238)));
    layer0_outputs(3320) <= inputs(123);
    layer0_outputs(3321) <= (inputs(15)) and not (inputs(53));
    layer0_outputs(3322) <= (inputs(245)) xor (inputs(214));
    layer0_outputs(3323) <= not((inputs(1)) or (inputs(35)));
    layer0_outputs(3324) <= not(inputs(59)) or (inputs(16));
    layer0_outputs(3325) <= not(inputs(70)) or (inputs(145));
    layer0_outputs(3326) <= '1';
    layer0_outputs(3327) <= not((inputs(85)) xor (inputs(229)));
    layer0_outputs(3328) <= inputs(53);
    layer0_outputs(3329) <= not((inputs(191)) or (inputs(78)));
    layer0_outputs(3330) <= not(inputs(188));
    layer0_outputs(3331) <= (inputs(122)) and not (inputs(164));
    layer0_outputs(3332) <= (inputs(208)) xor (inputs(222));
    layer0_outputs(3333) <= not((inputs(48)) or (inputs(119)));
    layer0_outputs(3334) <= not((inputs(60)) xor (inputs(186)));
    layer0_outputs(3335) <= not((inputs(133)) and (inputs(136)));
    layer0_outputs(3336) <= '1';
    layer0_outputs(3337) <= not(inputs(251)) or (inputs(55));
    layer0_outputs(3338) <= not((inputs(120)) and (inputs(72)));
    layer0_outputs(3339) <= not(inputs(237));
    layer0_outputs(3340) <= (inputs(218)) xor (inputs(186));
    layer0_outputs(3341) <= not(inputs(7));
    layer0_outputs(3342) <= (inputs(64)) or (inputs(2));
    layer0_outputs(3343) <= (inputs(158)) xor (inputs(78));
    layer0_outputs(3344) <= not((inputs(20)) xor (inputs(237)));
    layer0_outputs(3345) <= (inputs(214)) or (inputs(95));
    layer0_outputs(3346) <= not(inputs(117)) or (inputs(94));
    layer0_outputs(3347) <= not(inputs(178));
    layer0_outputs(3348) <= not((inputs(236)) or (inputs(215)));
    layer0_outputs(3349) <= not((inputs(15)) xor (inputs(145)));
    layer0_outputs(3350) <= not((inputs(181)) or (inputs(194)));
    layer0_outputs(3351) <= (inputs(199)) or (inputs(234));
    layer0_outputs(3352) <= not((inputs(68)) or (inputs(198)));
    layer0_outputs(3353) <= not((inputs(222)) or (inputs(216)));
    layer0_outputs(3354) <= not((inputs(133)) xor (inputs(86)));
    layer0_outputs(3355) <= not((inputs(25)) or (inputs(143)));
    layer0_outputs(3356) <= not(inputs(19));
    layer0_outputs(3357) <= '0';
    layer0_outputs(3358) <= (inputs(222)) or (inputs(198));
    layer0_outputs(3359) <= inputs(101);
    layer0_outputs(3360) <= not((inputs(210)) xor (inputs(219)));
    layer0_outputs(3361) <= not(inputs(77));
    layer0_outputs(3362) <= not(inputs(44));
    layer0_outputs(3363) <= (inputs(183)) xor (inputs(238));
    layer0_outputs(3364) <= inputs(229);
    layer0_outputs(3365) <= not(inputs(212)) or (inputs(130));
    layer0_outputs(3366) <= not(inputs(166));
    layer0_outputs(3367) <= (inputs(40)) and (inputs(38));
    layer0_outputs(3368) <= inputs(91);
    layer0_outputs(3369) <= not(inputs(91)) or (inputs(240));
    layer0_outputs(3370) <= not(inputs(179));
    layer0_outputs(3371) <= '0';
    layer0_outputs(3372) <= (inputs(205)) and not (inputs(77));
    layer0_outputs(3373) <= not(inputs(58));
    layer0_outputs(3374) <= (inputs(173)) xor (inputs(111));
    layer0_outputs(3375) <= not(inputs(148));
    layer0_outputs(3376) <= inputs(42);
    layer0_outputs(3377) <= (inputs(81)) xor (inputs(68));
    layer0_outputs(3378) <= inputs(221);
    layer0_outputs(3379) <= not((inputs(213)) or (inputs(234)));
    layer0_outputs(3380) <= not(inputs(210));
    layer0_outputs(3381) <= (inputs(38)) and not (inputs(163));
    layer0_outputs(3382) <= not((inputs(225)) or (inputs(21)));
    layer0_outputs(3383) <= not(inputs(110));
    layer0_outputs(3384) <= not(inputs(156));
    layer0_outputs(3385) <= inputs(154);
    layer0_outputs(3386) <= not(inputs(147));
    layer0_outputs(3387) <= '1';
    layer0_outputs(3388) <= '0';
    layer0_outputs(3389) <= '1';
    layer0_outputs(3390) <= not((inputs(161)) or (inputs(162)));
    layer0_outputs(3391) <= not(inputs(129));
    layer0_outputs(3392) <= (inputs(173)) xor (inputs(237));
    layer0_outputs(3393) <= '0';
    layer0_outputs(3394) <= (inputs(69)) or (inputs(25));
    layer0_outputs(3395) <= not((inputs(100)) and (inputs(140)));
    layer0_outputs(3396) <= not((inputs(42)) xor (inputs(13)));
    layer0_outputs(3397) <= inputs(231);
    layer0_outputs(3398) <= not(inputs(183));
    layer0_outputs(3399) <= not(inputs(230)) or (inputs(59));
    layer0_outputs(3400) <= not((inputs(93)) and (inputs(79)));
    layer0_outputs(3401) <= not((inputs(8)) or (inputs(128)));
    layer0_outputs(3402) <= (inputs(57)) and not (inputs(102));
    layer0_outputs(3403) <= not((inputs(96)) xor (inputs(210)));
    layer0_outputs(3404) <= not((inputs(230)) or (inputs(82)));
    layer0_outputs(3405) <= (inputs(163)) or (inputs(181));
    layer0_outputs(3406) <= not((inputs(224)) and (inputs(217)));
    layer0_outputs(3407) <= (inputs(171)) and not (inputs(49));
    layer0_outputs(3408) <= (inputs(18)) xor (inputs(0));
    layer0_outputs(3409) <= (inputs(228)) and not (inputs(174));
    layer0_outputs(3410) <= (inputs(185)) or (inputs(181));
    layer0_outputs(3411) <= not((inputs(86)) and (inputs(230)));
    layer0_outputs(3412) <= (inputs(52)) and (inputs(23));
    layer0_outputs(3413) <= not((inputs(28)) or (inputs(248)));
    layer0_outputs(3414) <= '0';
    layer0_outputs(3415) <= (inputs(101)) or (inputs(197));
    layer0_outputs(3416) <= inputs(133);
    layer0_outputs(3417) <= (inputs(110)) xor (inputs(92));
    layer0_outputs(3418) <= (inputs(179)) or (inputs(6));
    layer0_outputs(3419) <= not((inputs(217)) or (inputs(185)));
    layer0_outputs(3420) <= (inputs(231)) and not (inputs(92));
    layer0_outputs(3421) <= (inputs(208)) or (inputs(250));
    layer0_outputs(3422) <= (inputs(207)) or (inputs(238));
    layer0_outputs(3423) <= not(inputs(85)) or (inputs(32));
    layer0_outputs(3424) <= inputs(77);
    layer0_outputs(3425) <= (inputs(197)) xor (inputs(39));
    layer0_outputs(3426) <= not(inputs(48)) or (inputs(249));
    layer0_outputs(3427) <= (inputs(182)) and not (inputs(77));
    layer0_outputs(3428) <= not((inputs(228)) xor (inputs(40)));
    layer0_outputs(3429) <= not((inputs(106)) or (inputs(180)));
    layer0_outputs(3430) <= (inputs(217)) or (inputs(201));
    layer0_outputs(3431) <= inputs(13);
    layer0_outputs(3432) <= not(inputs(20));
    layer0_outputs(3433) <= not(inputs(132));
    layer0_outputs(3434) <= not(inputs(36)) or (inputs(226));
    layer0_outputs(3435) <= (inputs(179)) and not (inputs(112));
    layer0_outputs(3436) <= (inputs(144)) xor (inputs(230));
    layer0_outputs(3437) <= inputs(136);
    layer0_outputs(3438) <= (inputs(80)) or (inputs(25));
    layer0_outputs(3439) <= inputs(19);
    layer0_outputs(3440) <= '1';
    layer0_outputs(3441) <= not(inputs(201)) or (inputs(115));
    layer0_outputs(3442) <= not(inputs(7));
    layer0_outputs(3443) <= not((inputs(64)) xor (inputs(6)));
    layer0_outputs(3444) <= not(inputs(172)) or (inputs(2));
    layer0_outputs(3445) <= '0';
    layer0_outputs(3446) <= not(inputs(7)) or (inputs(168));
    layer0_outputs(3447) <= (inputs(184)) or (inputs(97));
    layer0_outputs(3448) <= inputs(146);
    layer0_outputs(3449) <= not(inputs(167)) or (inputs(41));
    layer0_outputs(3450) <= (inputs(91)) or (inputs(77));
    layer0_outputs(3451) <= not(inputs(34));
    layer0_outputs(3452) <= '0';
    layer0_outputs(3453) <= (inputs(40)) or (inputs(55));
    layer0_outputs(3454) <= inputs(139);
    layer0_outputs(3455) <= (inputs(160)) and (inputs(82));
    layer0_outputs(3456) <= not(inputs(254));
    layer0_outputs(3457) <= (inputs(165)) xor (inputs(77));
    layer0_outputs(3458) <= (inputs(180)) and (inputs(184));
    layer0_outputs(3459) <= not((inputs(134)) or (inputs(199)));
    layer0_outputs(3460) <= (inputs(134)) and not (inputs(113));
    layer0_outputs(3461) <= not((inputs(52)) or (inputs(10)));
    layer0_outputs(3462) <= (inputs(155)) or (inputs(233));
    layer0_outputs(3463) <= (inputs(19)) xor (inputs(250));
    layer0_outputs(3464) <= (inputs(90)) and not (inputs(174));
    layer0_outputs(3465) <= not((inputs(117)) or (inputs(208)));
    layer0_outputs(3466) <= not(inputs(255));
    layer0_outputs(3467) <= (inputs(146)) and not (inputs(31));
    layer0_outputs(3468) <= (inputs(226)) xor (inputs(213));
    layer0_outputs(3469) <= (inputs(154)) and not (inputs(25));
    layer0_outputs(3470) <= not((inputs(29)) xor (inputs(76)));
    layer0_outputs(3471) <= inputs(113);
    layer0_outputs(3472) <= '1';
    layer0_outputs(3473) <= (inputs(61)) or (inputs(39));
    layer0_outputs(3474) <= not(inputs(219)) or (inputs(123));
    layer0_outputs(3475) <= not(inputs(89)) or (inputs(135));
    layer0_outputs(3476) <= (inputs(10)) or (inputs(82));
    layer0_outputs(3477) <= not((inputs(16)) or (inputs(3)));
    layer0_outputs(3478) <= '1';
    layer0_outputs(3479) <= not((inputs(84)) or (inputs(52)));
    layer0_outputs(3480) <= not((inputs(74)) xor (inputs(222)));
    layer0_outputs(3481) <= not((inputs(73)) xor (inputs(135)));
    layer0_outputs(3482) <= not(inputs(22));
    layer0_outputs(3483) <= (inputs(167)) and not (inputs(189));
    layer0_outputs(3484) <= '0';
    layer0_outputs(3485) <= not(inputs(120));
    layer0_outputs(3486) <= not(inputs(195)) or (inputs(253));
    layer0_outputs(3487) <= not(inputs(188));
    layer0_outputs(3488) <= (inputs(5)) xor (inputs(125));
    layer0_outputs(3489) <= not(inputs(228));
    layer0_outputs(3490) <= (inputs(167)) or (inputs(249));
    layer0_outputs(3491) <= not(inputs(122));
    layer0_outputs(3492) <= (inputs(85)) xor (inputs(23));
    layer0_outputs(3493) <= not(inputs(72)) or (inputs(1));
    layer0_outputs(3494) <= '0';
    layer0_outputs(3495) <= not(inputs(74));
    layer0_outputs(3496) <= (inputs(76)) or (inputs(94));
    layer0_outputs(3497) <= inputs(76);
    layer0_outputs(3498) <= (inputs(197)) and (inputs(167));
    layer0_outputs(3499) <= not((inputs(174)) or (inputs(99)));
    layer0_outputs(3500) <= '0';
    layer0_outputs(3501) <= (inputs(130)) or (inputs(192));
    layer0_outputs(3502) <= not((inputs(75)) or (inputs(9)));
    layer0_outputs(3503) <= not(inputs(189));
    layer0_outputs(3504) <= not(inputs(130)) or (inputs(208));
    layer0_outputs(3505) <= not(inputs(97));
    layer0_outputs(3506) <= not(inputs(170));
    layer0_outputs(3507) <= not((inputs(52)) and (inputs(110)));
    layer0_outputs(3508) <= (inputs(136)) xor (inputs(254));
    layer0_outputs(3509) <= not(inputs(20)) or (inputs(99));
    layer0_outputs(3510) <= not((inputs(130)) or (inputs(11)));
    layer0_outputs(3511) <= (inputs(141)) and (inputs(20));
    layer0_outputs(3512) <= (inputs(54)) and not (inputs(110));
    layer0_outputs(3513) <= not(inputs(218));
    layer0_outputs(3514) <= not(inputs(117));
    layer0_outputs(3515) <= not(inputs(74));
    layer0_outputs(3516) <= '0';
    layer0_outputs(3517) <= (inputs(31)) and (inputs(27));
    layer0_outputs(3518) <= not(inputs(40));
    layer0_outputs(3519) <= not(inputs(72)) or (inputs(50));
    layer0_outputs(3520) <= not((inputs(104)) xor (inputs(62)));
    layer0_outputs(3521) <= not(inputs(6)) or (inputs(97));
    layer0_outputs(3522) <= not(inputs(211)) or (inputs(1));
    layer0_outputs(3523) <= not((inputs(48)) and (inputs(75)));
    layer0_outputs(3524) <= inputs(98);
    layer0_outputs(3525) <= (inputs(144)) xor (inputs(204));
    layer0_outputs(3526) <= '1';
    layer0_outputs(3527) <= (inputs(117)) and not (inputs(126));
    layer0_outputs(3528) <= (inputs(72)) and not (inputs(13));
    layer0_outputs(3529) <= (inputs(16)) xor (inputs(7));
    layer0_outputs(3530) <= (inputs(168)) xor (inputs(15));
    layer0_outputs(3531) <= (inputs(245)) and (inputs(249));
    layer0_outputs(3532) <= (inputs(60)) and not (inputs(38));
    layer0_outputs(3533) <= (inputs(55)) or (inputs(131));
    layer0_outputs(3534) <= inputs(89);
    layer0_outputs(3535) <= not((inputs(208)) or (inputs(24)));
    layer0_outputs(3536) <= not((inputs(51)) xor (inputs(19)));
    layer0_outputs(3537) <= (inputs(183)) and not (inputs(186));
    layer0_outputs(3538) <= (inputs(5)) xor (inputs(215));
    layer0_outputs(3539) <= inputs(78);
    layer0_outputs(3540) <= not((inputs(24)) or (inputs(8)));
    layer0_outputs(3541) <= not((inputs(88)) or (inputs(39)));
    layer0_outputs(3542) <= not((inputs(47)) or (inputs(22)));
    layer0_outputs(3543) <= (inputs(214)) and not (inputs(50));
    layer0_outputs(3544) <= (inputs(0)) xor (inputs(145));
    layer0_outputs(3545) <= not((inputs(193)) xor (inputs(254)));
    layer0_outputs(3546) <= (inputs(201)) xor (inputs(191));
    layer0_outputs(3547) <= not((inputs(33)) or (inputs(18)));
    layer0_outputs(3548) <= not(inputs(204)) or (inputs(154));
    layer0_outputs(3549) <= not(inputs(103));
    layer0_outputs(3550) <= not((inputs(53)) xor (inputs(21)));
    layer0_outputs(3551) <= not(inputs(255)) or (inputs(59));
    layer0_outputs(3552) <= (inputs(34)) xor (inputs(3));
    layer0_outputs(3553) <= (inputs(35)) and not (inputs(59));
    layer0_outputs(3554) <= (inputs(21)) xor (inputs(108));
    layer0_outputs(3555) <= (inputs(113)) xor (inputs(5));
    layer0_outputs(3556) <= inputs(26);
    layer0_outputs(3557) <= (inputs(151)) or (inputs(118));
    layer0_outputs(3558) <= (inputs(90)) and (inputs(115));
    layer0_outputs(3559) <= not(inputs(52)) or (inputs(195));
    layer0_outputs(3560) <= (inputs(96)) or (inputs(94));
    layer0_outputs(3561) <= not(inputs(117));
    layer0_outputs(3562) <= not(inputs(93));
    layer0_outputs(3563) <= not((inputs(180)) or (inputs(197)));
    layer0_outputs(3564) <= not((inputs(206)) xor (inputs(114)));
    layer0_outputs(3565) <= (inputs(238)) and (inputs(158));
    layer0_outputs(3566) <= not((inputs(168)) or (inputs(170)));
    layer0_outputs(3567) <= not(inputs(23));
    layer0_outputs(3568) <= (inputs(29)) or (inputs(17));
    layer0_outputs(3569) <= not(inputs(147));
    layer0_outputs(3570) <= inputs(49);
    layer0_outputs(3571) <= (inputs(240)) and not (inputs(29));
    layer0_outputs(3572) <= inputs(198);
    layer0_outputs(3573) <= not((inputs(146)) xor (inputs(246)));
    layer0_outputs(3574) <= (inputs(28)) or (inputs(5));
    layer0_outputs(3575) <= not(inputs(41)) or (inputs(167));
    layer0_outputs(3576) <= '0';
    layer0_outputs(3577) <= inputs(188);
    layer0_outputs(3578) <= not(inputs(41));
    layer0_outputs(3579) <= (inputs(234)) or (inputs(168));
    layer0_outputs(3580) <= not((inputs(204)) or (inputs(177)));
    layer0_outputs(3581) <= (inputs(76)) and (inputs(9));
    layer0_outputs(3582) <= inputs(193);
    layer0_outputs(3583) <= not((inputs(52)) xor (inputs(21)));
    layer0_outputs(3584) <= not(inputs(181));
    layer0_outputs(3585) <= not(inputs(112)) or (inputs(111));
    layer0_outputs(3586) <= (inputs(70)) or (inputs(119));
    layer0_outputs(3587) <= inputs(21);
    layer0_outputs(3588) <= (inputs(92)) and not (inputs(207));
    layer0_outputs(3589) <= '1';
    layer0_outputs(3590) <= not(inputs(154));
    layer0_outputs(3591) <= not((inputs(63)) or (inputs(37)));
    layer0_outputs(3592) <= not((inputs(81)) and (inputs(138)));
    layer0_outputs(3593) <= (inputs(176)) xor (inputs(253));
    layer0_outputs(3594) <= inputs(30);
    layer0_outputs(3595) <= not((inputs(144)) or (inputs(170)));
    layer0_outputs(3596) <= not(inputs(41)) or (inputs(168));
    layer0_outputs(3597) <= not(inputs(108));
    layer0_outputs(3598) <= '0';
    layer0_outputs(3599) <= (inputs(239)) or (inputs(36));
    layer0_outputs(3600) <= (inputs(167)) and (inputs(24));
    layer0_outputs(3601) <= inputs(27);
    layer0_outputs(3602) <= inputs(63);
    layer0_outputs(3603) <= (inputs(159)) or (inputs(232));
    layer0_outputs(3604) <= not(inputs(125)) or (inputs(225));
    layer0_outputs(3605) <= (inputs(24)) or (inputs(250));
    layer0_outputs(3606) <= (inputs(104)) or (inputs(83));
    layer0_outputs(3607) <= inputs(237);
    layer0_outputs(3608) <= not(inputs(183)) or (inputs(113));
    layer0_outputs(3609) <= not(inputs(20));
    layer0_outputs(3610) <= not(inputs(11));
    layer0_outputs(3611) <= inputs(146);
    layer0_outputs(3612) <= not((inputs(146)) or (inputs(46)));
    layer0_outputs(3613) <= (inputs(128)) and not (inputs(171));
    layer0_outputs(3614) <= not(inputs(253)) or (inputs(17));
    layer0_outputs(3615) <= (inputs(157)) or (inputs(236));
    layer0_outputs(3616) <= not((inputs(142)) and (inputs(133)));
    layer0_outputs(3617) <= inputs(15);
    layer0_outputs(3618) <= not((inputs(104)) and (inputs(46)));
    layer0_outputs(3619) <= not((inputs(89)) or (inputs(104)));
    layer0_outputs(3620) <= not((inputs(133)) and (inputs(232)));
    layer0_outputs(3621) <= (inputs(139)) xor (inputs(27));
    layer0_outputs(3622) <= not((inputs(23)) and (inputs(230)));
    layer0_outputs(3623) <= not((inputs(150)) or (inputs(80)));
    layer0_outputs(3624) <= not(inputs(125));
    layer0_outputs(3625) <= inputs(144);
    layer0_outputs(3626) <= (inputs(29)) or (inputs(156));
    layer0_outputs(3627) <= '0';
    layer0_outputs(3628) <= inputs(135);
    layer0_outputs(3629) <= not(inputs(9));
    layer0_outputs(3630) <= (inputs(120)) xor (inputs(154));
    layer0_outputs(3631) <= not((inputs(163)) or (inputs(140)));
    layer0_outputs(3632) <= not((inputs(71)) xor (inputs(35)));
    layer0_outputs(3633) <= not((inputs(197)) or (inputs(213)));
    layer0_outputs(3634) <= inputs(99);
    layer0_outputs(3635) <= not(inputs(228)) or (inputs(38));
    layer0_outputs(3636) <= (inputs(130)) or (inputs(50));
    layer0_outputs(3637) <= not(inputs(80));
    layer0_outputs(3638) <= not((inputs(13)) and (inputs(16)));
    layer0_outputs(3639) <= (inputs(214)) or (inputs(158));
    layer0_outputs(3640) <= (inputs(153)) or (inputs(18));
    layer0_outputs(3641) <= (inputs(37)) and (inputs(44));
    layer0_outputs(3642) <= not(inputs(56));
    layer0_outputs(3643) <= (inputs(83)) xor (inputs(127));
    layer0_outputs(3644) <= inputs(231);
    layer0_outputs(3645) <= not(inputs(130)) or (inputs(154));
    layer0_outputs(3646) <= inputs(216);
    layer0_outputs(3647) <= (inputs(155)) or (inputs(13));
    layer0_outputs(3648) <= not((inputs(69)) or (inputs(60)));
    layer0_outputs(3649) <= not((inputs(124)) and (inputs(165)));
    layer0_outputs(3650) <= not((inputs(222)) or (inputs(182)));
    layer0_outputs(3651) <= inputs(148);
    layer0_outputs(3652) <= inputs(91);
    layer0_outputs(3653) <= (inputs(236)) or (inputs(88));
    layer0_outputs(3654) <= not(inputs(172)) or (inputs(66));
    layer0_outputs(3655) <= (inputs(51)) and not (inputs(41));
    layer0_outputs(3656) <= not(inputs(112)) or (inputs(252));
    layer0_outputs(3657) <= inputs(193);
    layer0_outputs(3658) <= (inputs(243)) or (inputs(71));
    layer0_outputs(3659) <= not(inputs(131));
    layer0_outputs(3660) <= inputs(138);
    layer0_outputs(3661) <= (inputs(211)) xor (inputs(47));
    layer0_outputs(3662) <= not((inputs(120)) or (inputs(118)));
    layer0_outputs(3663) <= (inputs(17)) or (inputs(172));
    layer0_outputs(3664) <= inputs(204);
    layer0_outputs(3665) <= not(inputs(136));
    layer0_outputs(3666) <= not(inputs(15));
    layer0_outputs(3667) <= (inputs(145)) or (inputs(222));
    layer0_outputs(3668) <= not(inputs(38)) or (inputs(130));
    layer0_outputs(3669) <= not(inputs(137)) or (inputs(10));
    layer0_outputs(3670) <= (inputs(20)) or (inputs(220));
    layer0_outputs(3671) <= not(inputs(147));
    layer0_outputs(3672) <= not(inputs(162)) or (inputs(33));
    layer0_outputs(3673) <= (inputs(49)) and (inputs(80));
    layer0_outputs(3674) <= not(inputs(227));
    layer0_outputs(3675) <= (inputs(70)) and (inputs(71));
    layer0_outputs(3676) <= '1';
    layer0_outputs(3677) <= '0';
    layer0_outputs(3678) <= not(inputs(155)) or (inputs(167));
    layer0_outputs(3679) <= inputs(103);
    layer0_outputs(3680) <= not(inputs(13)) or (inputs(233));
    layer0_outputs(3681) <= not(inputs(135));
    layer0_outputs(3682) <= not(inputs(38)) or (inputs(46));
    layer0_outputs(3683) <= inputs(74);
    layer0_outputs(3684) <= (inputs(74)) and not (inputs(53));
    layer0_outputs(3685) <= inputs(98);
    layer0_outputs(3686) <= not(inputs(240));
    layer0_outputs(3687) <= not((inputs(6)) and (inputs(73)));
    layer0_outputs(3688) <= not(inputs(43)) or (inputs(167));
    layer0_outputs(3689) <= (inputs(61)) and not (inputs(96));
    layer0_outputs(3690) <= inputs(238);
    layer0_outputs(3691) <= (inputs(226)) and not (inputs(86));
    layer0_outputs(3692) <= '1';
    layer0_outputs(3693) <= inputs(123);
    layer0_outputs(3694) <= not((inputs(193)) or (inputs(249)));
    layer0_outputs(3695) <= (inputs(82)) or (inputs(116));
    layer0_outputs(3696) <= (inputs(195)) and not (inputs(33));
    layer0_outputs(3697) <= inputs(66);
    layer0_outputs(3698) <= inputs(193);
    layer0_outputs(3699) <= not((inputs(37)) xor (inputs(28)));
    layer0_outputs(3700) <= inputs(136);
    layer0_outputs(3701) <= '1';
    layer0_outputs(3702) <= not((inputs(244)) xor (inputs(182)));
    layer0_outputs(3703) <= not((inputs(175)) or (inputs(184)));
    layer0_outputs(3704) <= (inputs(151)) or (inputs(71));
    layer0_outputs(3705) <= (inputs(33)) and not (inputs(110));
    layer0_outputs(3706) <= (inputs(49)) xor (inputs(18));
    layer0_outputs(3707) <= inputs(137);
    layer0_outputs(3708) <= (inputs(203)) and not (inputs(29));
    layer0_outputs(3709) <= not((inputs(238)) or (inputs(91)));
    layer0_outputs(3710) <= not((inputs(211)) and (inputs(211)));
    layer0_outputs(3711) <= (inputs(11)) and not (inputs(172));
    layer0_outputs(3712) <= (inputs(138)) and not (inputs(192));
    layer0_outputs(3713) <= not((inputs(142)) and (inputs(250)));
    layer0_outputs(3714) <= not(inputs(152));
    layer0_outputs(3715) <= '1';
    layer0_outputs(3716) <= (inputs(149)) and not (inputs(41));
    layer0_outputs(3717) <= (inputs(61)) and not (inputs(113));
    layer0_outputs(3718) <= '1';
    layer0_outputs(3719) <= not(inputs(40)) or (inputs(178));
    layer0_outputs(3720) <= not(inputs(250)) or (inputs(140));
    layer0_outputs(3721) <= not(inputs(154));
    layer0_outputs(3722) <= inputs(82);
    layer0_outputs(3723) <= (inputs(176)) xor (inputs(83));
    layer0_outputs(3724) <= (inputs(80)) or (inputs(165));
    layer0_outputs(3725) <= (inputs(177)) and not (inputs(51));
    layer0_outputs(3726) <= not(inputs(177));
    layer0_outputs(3727) <= not(inputs(148));
    layer0_outputs(3728) <= not((inputs(32)) xor (inputs(51)));
    layer0_outputs(3729) <= (inputs(249)) and not (inputs(20));
    layer0_outputs(3730) <= inputs(121);
    layer0_outputs(3731) <= not((inputs(20)) and (inputs(185)));
    layer0_outputs(3732) <= (inputs(28)) and (inputs(111));
    layer0_outputs(3733) <= not((inputs(202)) and (inputs(215)));
    layer0_outputs(3734) <= not((inputs(43)) xor (inputs(70)));
    layer0_outputs(3735) <= '0';
    layer0_outputs(3736) <= (inputs(163)) and (inputs(131));
    layer0_outputs(3737) <= (inputs(135)) and not (inputs(195));
    layer0_outputs(3738) <= (inputs(165)) and (inputs(6));
    layer0_outputs(3739) <= (inputs(64)) or (inputs(241));
    layer0_outputs(3740) <= not(inputs(28));
    layer0_outputs(3741) <= not(inputs(112));
    layer0_outputs(3742) <= '1';
    layer0_outputs(3743) <= not((inputs(25)) xor (inputs(73)));
    layer0_outputs(3744) <= not((inputs(171)) and (inputs(132)));
    layer0_outputs(3745) <= not(inputs(167));
    layer0_outputs(3746) <= not(inputs(26)) or (inputs(254));
    layer0_outputs(3747) <= inputs(75);
    layer0_outputs(3748) <= not(inputs(197));
    layer0_outputs(3749) <= (inputs(60)) and not (inputs(222));
    layer0_outputs(3750) <= not((inputs(161)) or (inputs(79)));
    layer0_outputs(3751) <= (inputs(25)) xor (inputs(231));
    layer0_outputs(3752) <= not((inputs(156)) or (inputs(220)));
    layer0_outputs(3753) <= not(inputs(180));
    layer0_outputs(3754) <= (inputs(113)) or (inputs(200));
    layer0_outputs(3755) <= (inputs(76)) or (inputs(147));
    layer0_outputs(3756) <= (inputs(42)) or (inputs(158));
    layer0_outputs(3757) <= (inputs(179)) and not (inputs(123));
    layer0_outputs(3758) <= (inputs(155)) and (inputs(154));
    layer0_outputs(3759) <= not(inputs(253));
    layer0_outputs(3760) <= not((inputs(238)) or (inputs(169)));
    layer0_outputs(3761) <= '1';
    layer0_outputs(3762) <= not(inputs(63)) or (inputs(180));
    layer0_outputs(3763) <= not(inputs(188)) or (inputs(223));
    layer0_outputs(3764) <= not((inputs(184)) or (inputs(2)));
    layer0_outputs(3765) <= not(inputs(22));
    layer0_outputs(3766) <= (inputs(122)) and not (inputs(227));
    layer0_outputs(3767) <= inputs(123);
    layer0_outputs(3768) <= inputs(211);
    layer0_outputs(3769) <= inputs(167);
    layer0_outputs(3770) <= not(inputs(193)) or (inputs(93));
    layer0_outputs(3771) <= inputs(104);
    layer0_outputs(3772) <= not((inputs(6)) xor (inputs(34)));
    layer0_outputs(3773) <= not(inputs(61)) or (inputs(144));
    layer0_outputs(3774) <= (inputs(18)) or (inputs(38));
    layer0_outputs(3775) <= (inputs(222)) and not (inputs(38));
    layer0_outputs(3776) <= (inputs(144)) or (inputs(87));
    layer0_outputs(3777) <= not(inputs(80));
    layer0_outputs(3778) <= inputs(124);
    layer0_outputs(3779) <= not(inputs(174));
    layer0_outputs(3780) <= (inputs(163)) xor (inputs(145));
    layer0_outputs(3781) <= inputs(118);
    layer0_outputs(3782) <= inputs(204);
    layer0_outputs(3783) <= (inputs(8)) and not (inputs(99));
    layer0_outputs(3784) <= (inputs(49)) xor (inputs(152));
    layer0_outputs(3785) <= not(inputs(39)) or (inputs(29));
    layer0_outputs(3786) <= '0';
    layer0_outputs(3787) <= not(inputs(114));
    layer0_outputs(3788) <= not((inputs(99)) xor (inputs(62)));
    layer0_outputs(3789) <= not(inputs(245)) or (inputs(167));
    layer0_outputs(3790) <= inputs(145);
    layer0_outputs(3791) <= (inputs(101)) and (inputs(49));
    layer0_outputs(3792) <= not((inputs(50)) or (inputs(87)));
    layer0_outputs(3793) <= (inputs(195)) and not (inputs(63));
    layer0_outputs(3794) <= not((inputs(150)) and (inputs(67)));
    layer0_outputs(3795) <= not((inputs(125)) or (inputs(139)));
    layer0_outputs(3796) <= (inputs(230)) or (inputs(245));
    layer0_outputs(3797) <= not((inputs(190)) xor (inputs(107)));
    layer0_outputs(3798) <= not(inputs(176));
    layer0_outputs(3799) <= (inputs(170)) and not (inputs(113));
    layer0_outputs(3800) <= not(inputs(189)) or (inputs(216));
    layer0_outputs(3801) <= not(inputs(101)) or (inputs(194));
    layer0_outputs(3802) <= not(inputs(239)) or (inputs(160));
    layer0_outputs(3803) <= not((inputs(144)) or (inputs(186)));
    layer0_outputs(3804) <= (inputs(85)) and not (inputs(1));
    layer0_outputs(3805) <= not(inputs(83));
    layer0_outputs(3806) <= not((inputs(156)) xor (inputs(29)));
    layer0_outputs(3807) <= inputs(105);
    layer0_outputs(3808) <= (inputs(161)) and not (inputs(44));
    layer0_outputs(3809) <= not(inputs(251)) or (inputs(49));
    layer0_outputs(3810) <= not(inputs(101)) or (inputs(172));
    layer0_outputs(3811) <= not((inputs(33)) or (inputs(122)));
    layer0_outputs(3812) <= not((inputs(28)) and (inputs(69)));
    layer0_outputs(3813) <= '1';
    layer0_outputs(3814) <= not((inputs(199)) xor (inputs(8)));
    layer0_outputs(3815) <= not(inputs(90));
    layer0_outputs(3816) <= (inputs(89)) or (inputs(211));
    layer0_outputs(3817) <= not((inputs(15)) or (inputs(249)));
    layer0_outputs(3818) <= not((inputs(96)) xor (inputs(86)));
    layer0_outputs(3819) <= not((inputs(29)) or (inputs(44)));
    layer0_outputs(3820) <= not(inputs(198));
    layer0_outputs(3821) <= not((inputs(181)) and (inputs(116)));
    layer0_outputs(3822) <= inputs(34);
    layer0_outputs(3823) <= (inputs(235)) xor (inputs(209));
    layer0_outputs(3824) <= (inputs(42)) and (inputs(23));
    layer0_outputs(3825) <= (inputs(150)) and not (inputs(234));
    layer0_outputs(3826) <= (inputs(214)) and not (inputs(64));
    layer0_outputs(3827) <= (inputs(231)) and not (inputs(90));
    layer0_outputs(3828) <= inputs(78);
    layer0_outputs(3829) <= not(inputs(21)) or (inputs(114));
    layer0_outputs(3830) <= not((inputs(239)) and (inputs(207)));
    layer0_outputs(3831) <= not((inputs(248)) xor (inputs(218)));
    layer0_outputs(3832) <= inputs(155);
    layer0_outputs(3833) <= (inputs(103)) and not (inputs(63));
    layer0_outputs(3834) <= not((inputs(56)) and (inputs(19)));
    layer0_outputs(3835) <= '1';
    layer0_outputs(3836) <= (inputs(52)) and not (inputs(219));
    layer0_outputs(3837) <= '1';
    layer0_outputs(3838) <= not(inputs(150)) or (inputs(55));
    layer0_outputs(3839) <= not(inputs(219)) or (inputs(29));
    layer0_outputs(3840) <= not(inputs(110));
    layer0_outputs(3841) <= (inputs(153)) and not (inputs(56));
    layer0_outputs(3842) <= not(inputs(163));
    layer0_outputs(3843) <= inputs(67);
    layer0_outputs(3844) <= inputs(131);
    layer0_outputs(3845) <= (inputs(141)) or (inputs(122));
    layer0_outputs(3846) <= not(inputs(207)) or (inputs(122));
    layer0_outputs(3847) <= (inputs(4)) or (inputs(31));
    layer0_outputs(3848) <= (inputs(228)) and not (inputs(142));
    layer0_outputs(3849) <= (inputs(165)) and not (inputs(165));
    layer0_outputs(3850) <= (inputs(203)) or (inputs(255));
    layer0_outputs(3851) <= '1';
    layer0_outputs(3852) <= not(inputs(122)) or (inputs(56));
    layer0_outputs(3853) <= not(inputs(183));
    layer0_outputs(3854) <= not(inputs(119));
    layer0_outputs(3855) <= (inputs(154)) and not (inputs(204));
    layer0_outputs(3856) <= not(inputs(92)) or (inputs(40));
    layer0_outputs(3857) <= not(inputs(164));
    layer0_outputs(3858) <= not((inputs(35)) and (inputs(38)));
    layer0_outputs(3859) <= not(inputs(219)) or (inputs(237));
    layer0_outputs(3860) <= not(inputs(164)) or (inputs(254));
    layer0_outputs(3861) <= not((inputs(151)) or (inputs(15)));
    layer0_outputs(3862) <= (inputs(130)) and not (inputs(240));
    layer0_outputs(3863) <= inputs(237);
    layer0_outputs(3864) <= (inputs(207)) and not (inputs(32));
    layer0_outputs(3865) <= not(inputs(47)) or (inputs(205));
    layer0_outputs(3866) <= not(inputs(32));
    layer0_outputs(3867) <= inputs(60);
    layer0_outputs(3868) <= inputs(194);
    layer0_outputs(3869) <= not(inputs(138)) or (inputs(31));
    layer0_outputs(3870) <= not((inputs(170)) or (inputs(88)));
    layer0_outputs(3871) <= (inputs(14)) and not (inputs(239));
    layer0_outputs(3872) <= inputs(75);
    layer0_outputs(3873) <= not((inputs(80)) xor (inputs(103)));
    layer0_outputs(3874) <= not(inputs(9));
    layer0_outputs(3875) <= inputs(25);
    layer0_outputs(3876) <= '1';
    layer0_outputs(3877) <= not(inputs(168));
    layer0_outputs(3878) <= (inputs(43)) and not (inputs(101));
    layer0_outputs(3879) <= not(inputs(45));
    layer0_outputs(3880) <= inputs(213);
    layer0_outputs(3881) <= inputs(69);
    layer0_outputs(3882) <= (inputs(151)) and not (inputs(156));
    layer0_outputs(3883) <= not(inputs(135));
    layer0_outputs(3884) <= (inputs(239)) xor (inputs(89));
    layer0_outputs(3885) <= (inputs(22)) or (inputs(37));
    layer0_outputs(3886) <= not((inputs(242)) or (inputs(2)));
    layer0_outputs(3887) <= (inputs(9)) and not (inputs(205));
    layer0_outputs(3888) <= not((inputs(52)) or (inputs(26)));
    layer0_outputs(3889) <= '0';
    layer0_outputs(3890) <= (inputs(40)) and not (inputs(129));
    layer0_outputs(3891) <= not(inputs(100));
    layer0_outputs(3892) <= not(inputs(52));
    layer0_outputs(3893) <= not((inputs(119)) xor (inputs(89)));
    layer0_outputs(3894) <= not((inputs(187)) or (inputs(122)));
    layer0_outputs(3895) <= not(inputs(44));
    layer0_outputs(3896) <= (inputs(120)) and not (inputs(19));
    layer0_outputs(3897) <= (inputs(248)) and (inputs(234));
    layer0_outputs(3898) <= not(inputs(105)) or (inputs(8));
    layer0_outputs(3899) <= (inputs(132)) or (inputs(122));
    layer0_outputs(3900) <= not(inputs(91)) or (inputs(87));
    layer0_outputs(3901) <= (inputs(240)) and (inputs(142));
    layer0_outputs(3902) <= inputs(36);
    layer0_outputs(3903) <= (inputs(163)) and not (inputs(142));
    layer0_outputs(3904) <= (inputs(196)) and (inputs(74));
    layer0_outputs(3905) <= not(inputs(147)) or (inputs(109));
    layer0_outputs(3906) <= not((inputs(118)) or (inputs(117)));
    layer0_outputs(3907) <= not(inputs(17));
    layer0_outputs(3908) <= (inputs(72)) and not (inputs(186));
    layer0_outputs(3909) <= (inputs(129)) or (inputs(75));
    layer0_outputs(3910) <= not(inputs(153)) or (inputs(40));
    layer0_outputs(3911) <= inputs(108);
    layer0_outputs(3912) <= not((inputs(175)) or (inputs(158)));
    layer0_outputs(3913) <= not((inputs(62)) or (inputs(192)));
    layer0_outputs(3914) <= inputs(154);
    layer0_outputs(3915) <= (inputs(37)) or (inputs(52));
    layer0_outputs(3916) <= (inputs(66)) or (inputs(210));
    layer0_outputs(3917) <= not((inputs(37)) or (inputs(84)));
    layer0_outputs(3918) <= not(inputs(194)) or (inputs(96));
    layer0_outputs(3919) <= not(inputs(177));
    layer0_outputs(3920) <= inputs(199);
    layer0_outputs(3921) <= not((inputs(93)) or (inputs(47)));
    layer0_outputs(3922) <= (inputs(27)) or (inputs(12));
    layer0_outputs(3923) <= (inputs(36)) xor (inputs(22));
    layer0_outputs(3924) <= '1';
    layer0_outputs(3925) <= (inputs(150)) or (inputs(250));
    layer0_outputs(3926) <= inputs(204);
    layer0_outputs(3927) <= (inputs(47)) xor (inputs(55));
    layer0_outputs(3928) <= (inputs(5)) and not (inputs(159));
    layer0_outputs(3929) <= '1';
    layer0_outputs(3930) <= not(inputs(101));
    layer0_outputs(3931) <= (inputs(204)) and not (inputs(240));
    layer0_outputs(3932) <= (inputs(224)) and not (inputs(238));
    layer0_outputs(3933) <= not((inputs(176)) xor (inputs(111)));
    layer0_outputs(3934) <= not(inputs(166));
    layer0_outputs(3935) <= inputs(43);
    layer0_outputs(3936) <= not(inputs(121));
    layer0_outputs(3937) <= (inputs(231)) xor (inputs(199));
    layer0_outputs(3938) <= inputs(220);
    layer0_outputs(3939) <= (inputs(130)) and not (inputs(162));
    layer0_outputs(3940) <= not(inputs(238)) or (inputs(15));
    layer0_outputs(3941) <= not(inputs(117));
    layer0_outputs(3942) <= not((inputs(195)) xor (inputs(227)));
    layer0_outputs(3943) <= '1';
    layer0_outputs(3944) <= inputs(69);
    layer0_outputs(3945) <= not(inputs(129));
    layer0_outputs(3946) <= not((inputs(90)) or (inputs(80)));
    layer0_outputs(3947) <= '1';
    layer0_outputs(3948) <= not(inputs(37));
    layer0_outputs(3949) <= (inputs(115)) and not (inputs(239));
    layer0_outputs(3950) <= not(inputs(82)) or (inputs(82));
    layer0_outputs(3951) <= (inputs(219)) and not (inputs(142));
    layer0_outputs(3952) <= '1';
    layer0_outputs(3953) <= not(inputs(39)) or (inputs(241));
    layer0_outputs(3954) <= (inputs(107)) and (inputs(228));
    layer0_outputs(3955) <= (inputs(152)) or (inputs(245));
    layer0_outputs(3956) <= inputs(56);
    layer0_outputs(3957) <= inputs(194);
    layer0_outputs(3958) <= (inputs(9)) and not (inputs(15));
    layer0_outputs(3959) <= (inputs(142)) and (inputs(186));
    layer0_outputs(3960) <= not((inputs(231)) xor (inputs(13)));
    layer0_outputs(3961) <= inputs(175);
    layer0_outputs(3962) <= (inputs(94)) xor (inputs(178));
    layer0_outputs(3963) <= not((inputs(176)) or (inputs(109)));
    layer0_outputs(3964) <= not((inputs(74)) and (inputs(69)));
    layer0_outputs(3965) <= (inputs(232)) or (inputs(11));
    layer0_outputs(3966) <= not(inputs(11));
    layer0_outputs(3967) <= not((inputs(101)) or (inputs(235)));
    layer0_outputs(3968) <= inputs(181);
    layer0_outputs(3969) <= (inputs(115)) and not (inputs(226));
    layer0_outputs(3970) <= not(inputs(39));
    layer0_outputs(3971) <= (inputs(50)) or (inputs(187));
    layer0_outputs(3972) <= not((inputs(252)) or (inputs(234)));
    layer0_outputs(3973) <= not(inputs(139)) or (inputs(13));
    layer0_outputs(3974) <= not((inputs(39)) or (inputs(0)));
    layer0_outputs(3975) <= not((inputs(204)) xor (inputs(241)));
    layer0_outputs(3976) <= (inputs(87)) and not (inputs(238));
    layer0_outputs(3977) <= inputs(83);
    layer0_outputs(3978) <= not((inputs(196)) or (inputs(167)));
    layer0_outputs(3979) <= not(inputs(181));
    layer0_outputs(3980) <= not(inputs(220));
    layer0_outputs(3981) <= not(inputs(69));
    layer0_outputs(3982) <= inputs(75);
    layer0_outputs(3983) <= inputs(57);
    layer0_outputs(3984) <= not((inputs(241)) or (inputs(147)));
    layer0_outputs(3985) <= inputs(79);
    layer0_outputs(3986) <= not(inputs(97));
    layer0_outputs(3987) <= (inputs(243)) or (inputs(159));
    layer0_outputs(3988) <= not(inputs(208));
    layer0_outputs(3989) <= not((inputs(201)) xor (inputs(179)));
    layer0_outputs(3990) <= not(inputs(172));
    layer0_outputs(3991) <= '1';
    layer0_outputs(3992) <= '0';
    layer0_outputs(3993) <= (inputs(185)) and not (inputs(225));
    layer0_outputs(3994) <= (inputs(128)) and not (inputs(213));
    layer0_outputs(3995) <= not((inputs(201)) and (inputs(215)));
    layer0_outputs(3996) <= inputs(59);
    layer0_outputs(3997) <= (inputs(179)) and not (inputs(97));
    layer0_outputs(3998) <= not((inputs(197)) or (inputs(249)));
    layer0_outputs(3999) <= not((inputs(208)) or (inputs(197)));
    layer0_outputs(4000) <= (inputs(128)) or (inputs(37));
    layer0_outputs(4001) <= (inputs(116)) xor (inputs(66));
    layer0_outputs(4002) <= (inputs(157)) and not (inputs(58));
    layer0_outputs(4003) <= (inputs(229)) xor (inputs(0));
    layer0_outputs(4004) <= not(inputs(156));
    layer0_outputs(4005) <= (inputs(178)) or (inputs(198));
    layer0_outputs(4006) <= (inputs(253)) and not (inputs(181));
    layer0_outputs(4007) <= (inputs(104)) and not (inputs(160));
    layer0_outputs(4008) <= not(inputs(7)) or (inputs(159));
    layer0_outputs(4009) <= not(inputs(89)) or (inputs(239));
    layer0_outputs(4010) <= not((inputs(21)) or (inputs(90)));
    layer0_outputs(4011) <= not((inputs(94)) xor (inputs(175)));
    layer0_outputs(4012) <= inputs(160);
    layer0_outputs(4013) <= (inputs(205)) and (inputs(253));
    layer0_outputs(4014) <= (inputs(249)) xor (inputs(247));
    layer0_outputs(4015) <= inputs(26);
    layer0_outputs(4016) <= not((inputs(213)) xor (inputs(241)));
    layer0_outputs(4017) <= not((inputs(128)) xor (inputs(171)));
    layer0_outputs(4018) <= not((inputs(102)) or (inputs(205)));
    layer0_outputs(4019) <= not((inputs(21)) xor (inputs(229)));
    layer0_outputs(4020) <= inputs(2);
    layer0_outputs(4021) <= (inputs(128)) and (inputs(47));
    layer0_outputs(4022) <= not(inputs(109));
    layer0_outputs(4023) <= (inputs(131)) xor (inputs(131));
    layer0_outputs(4024) <= not((inputs(229)) or (inputs(65)));
    layer0_outputs(4025) <= not((inputs(89)) or (inputs(136)));
    layer0_outputs(4026) <= not(inputs(160));
    layer0_outputs(4027) <= (inputs(6)) or (inputs(195));
    layer0_outputs(4028) <= (inputs(223)) and not (inputs(143));
    layer0_outputs(4029) <= inputs(183);
    layer0_outputs(4030) <= not((inputs(217)) and (inputs(80)));
    layer0_outputs(4031) <= not((inputs(66)) or (inputs(153)));
    layer0_outputs(4032) <= not((inputs(112)) or (inputs(210)));
    layer0_outputs(4033) <= not((inputs(248)) xor (inputs(216)));
    layer0_outputs(4034) <= inputs(22);
    layer0_outputs(4035) <= not((inputs(49)) or (inputs(90)));
    layer0_outputs(4036) <= '1';
    layer0_outputs(4037) <= inputs(51);
    layer0_outputs(4038) <= not(inputs(149));
    layer0_outputs(4039) <= not(inputs(152)) or (inputs(130));
    layer0_outputs(4040) <= not((inputs(149)) xor (inputs(87)));
    layer0_outputs(4041) <= not((inputs(125)) and (inputs(152)));
    layer0_outputs(4042) <= not(inputs(119));
    layer0_outputs(4043) <= (inputs(66)) or (inputs(141));
    layer0_outputs(4044) <= not(inputs(27)) or (inputs(221));
    layer0_outputs(4045) <= '0';
    layer0_outputs(4046) <= (inputs(208)) or (inputs(74));
    layer0_outputs(4047) <= (inputs(18)) and not (inputs(103));
    layer0_outputs(4048) <= (inputs(102)) and (inputs(145));
    layer0_outputs(4049) <= (inputs(103)) and not (inputs(68));
    layer0_outputs(4050) <= (inputs(23)) or (inputs(141));
    layer0_outputs(4051) <= (inputs(32)) and not (inputs(29));
    layer0_outputs(4052) <= not(inputs(183)) or (inputs(192));
    layer0_outputs(4053) <= not(inputs(47));
    layer0_outputs(4054) <= not(inputs(184));
    layer0_outputs(4055) <= '1';
    layer0_outputs(4056) <= inputs(195);
    layer0_outputs(4057) <= not(inputs(177));
    layer0_outputs(4058) <= not((inputs(63)) or (inputs(51)));
    layer0_outputs(4059) <= inputs(235);
    layer0_outputs(4060) <= not((inputs(195)) or (inputs(43)));
    layer0_outputs(4061) <= not(inputs(149));
    layer0_outputs(4062) <= (inputs(252)) or (inputs(148));
    layer0_outputs(4063) <= '1';
    layer0_outputs(4064) <= (inputs(33)) or (inputs(122));
    layer0_outputs(4065) <= not(inputs(100));
    layer0_outputs(4066) <= not(inputs(55)) or (inputs(73));
    layer0_outputs(4067) <= inputs(160);
    layer0_outputs(4068) <= not(inputs(178)) or (inputs(166));
    layer0_outputs(4069) <= not(inputs(167));
    layer0_outputs(4070) <= not(inputs(160));
    layer0_outputs(4071) <= '0';
    layer0_outputs(4072) <= not(inputs(109)) or (inputs(33));
    layer0_outputs(4073) <= not((inputs(137)) or (inputs(64)));
    layer0_outputs(4074) <= inputs(10);
    layer0_outputs(4075) <= not(inputs(34));
    layer0_outputs(4076) <= not(inputs(104)) or (inputs(58));
    layer0_outputs(4077) <= (inputs(246)) or (inputs(81));
    layer0_outputs(4078) <= inputs(33);
    layer0_outputs(4079) <= not(inputs(35));
    layer0_outputs(4080) <= (inputs(147)) and (inputs(163));
    layer0_outputs(4081) <= not(inputs(247));
    layer0_outputs(4082) <= not((inputs(142)) xor (inputs(86)));
    layer0_outputs(4083) <= inputs(217);
    layer0_outputs(4084) <= (inputs(40)) and not (inputs(242));
    layer0_outputs(4085) <= not(inputs(210));
    layer0_outputs(4086) <= (inputs(105)) and not (inputs(250));
    layer0_outputs(4087) <= (inputs(210)) or (inputs(217));
    layer0_outputs(4088) <= inputs(169);
    layer0_outputs(4089) <= not((inputs(74)) xor (inputs(6)));
    layer0_outputs(4090) <= not(inputs(242)) or (inputs(94));
    layer0_outputs(4091) <= not(inputs(205)) or (inputs(6));
    layer0_outputs(4092) <= (inputs(53)) and not (inputs(227));
    layer0_outputs(4093) <= not(inputs(44));
    layer0_outputs(4094) <= (inputs(194)) and not (inputs(129));
    layer0_outputs(4095) <= not((inputs(196)) or (inputs(71)));
    layer0_outputs(4096) <= not(inputs(131));
    layer0_outputs(4097) <= (inputs(154)) or (inputs(71));
    layer0_outputs(4098) <= (inputs(72)) or (inputs(204));
    layer0_outputs(4099) <= (inputs(245)) or (inputs(173));
    layer0_outputs(4100) <= not(inputs(27)) or (inputs(119));
    layer0_outputs(4101) <= inputs(245);
    layer0_outputs(4102) <= inputs(40);
    layer0_outputs(4103) <= (inputs(20)) and not (inputs(137));
    layer0_outputs(4104) <= not((inputs(237)) xor (inputs(69)));
    layer0_outputs(4105) <= (inputs(35)) and (inputs(243));
    layer0_outputs(4106) <= (inputs(254)) or (inputs(8));
    layer0_outputs(4107) <= (inputs(175)) and not (inputs(114));
    layer0_outputs(4108) <= (inputs(165)) or (inputs(17));
    layer0_outputs(4109) <= not(inputs(44));
    layer0_outputs(4110) <= (inputs(154)) xor (inputs(253));
    layer0_outputs(4111) <= not(inputs(7));
    layer0_outputs(4112) <= (inputs(105)) or (inputs(128));
    layer0_outputs(4113) <= not(inputs(59));
    layer0_outputs(4114) <= (inputs(45)) and not (inputs(132));
    layer0_outputs(4115) <= (inputs(64)) or (inputs(149));
    layer0_outputs(4116) <= '0';
    layer0_outputs(4117) <= inputs(164);
    layer0_outputs(4118) <= not((inputs(118)) or (inputs(20)));
    layer0_outputs(4119) <= (inputs(246)) and not (inputs(125));
    layer0_outputs(4120) <= not(inputs(10));
    layer0_outputs(4121) <= not(inputs(145)) or (inputs(121));
    layer0_outputs(4122) <= (inputs(209)) xor (inputs(217));
    layer0_outputs(4123) <= (inputs(204)) and (inputs(45));
    layer0_outputs(4124) <= (inputs(192)) or (inputs(179));
    layer0_outputs(4125) <= not((inputs(133)) or (inputs(80)));
    layer0_outputs(4126) <= not((inputs(39)) xor (inputs(8)));
    layer0_outputs(4127) <= not(inputs(149)) or (inputs(34));
    layer0_outputs(4128) <= '0';
    layer0_outputs(4129) <= inputs(216);
    layer0_outputs(4130) <= (inputs(127)) and not (inputs(48));
    layer0_outputs(4131) <= not(inputs(219));
    layer0_outputs(4132) <= (inputs(104)) and not (inputs(253));
    layer0_outputs(4133) <= not(inputs(158)) or (inputs(204));
    layer0_outputs(4134) <= not(inputs(42)) or (inputs(235));
    layer0_outputs(4135) <= not(inputs(189)) or (inputs(66));
    layer0_outputs(4136) <= not(inputs(104)) or (inputs(98));
    layer0_outputs(4137) <= (inputs(60)) xor (inputs(223));
    layer0_outputs(4138) <= not(inputs(102));
    layer0_outputs(4139) <= '0';
    layer0_outputs(4140) <= (inputs(218)) and (inputs(10));
    layer0_outputs(4141) <= inputs(248);
    layer0_outputs(4142) <= not(inputs(136));
    layer0_outputs(4143) <= not(inputs(75)) or (inputs(103));
    layer0_outputs(4144) <= (inputs(113)) xor (inputs(197));
    layer0_outputs(4145) <= not((inputs(180)) xor (inputs(135)));
    layer0_outputs(4146) <= not(inputs(40));
    layer0_outputs(4147) <= inputs(83);
    layer0_outputs(4148) <= not(inputs(22));
    layer0_outputs(4149) <= not((inputs(146)) or (inputs(85)));
    layer0_outputs(4150) <= (inputs(63)) and not (inputs(254));
    layer0_outputs(4151) <= not(inputs(7));
    layer0_outputs(4152) <= not(inputs(167));
    layer0_outputs(4153) <= not((inputs(136)) xor (inputs(155)));
    layer0_outputs(4154) <= (inputs(128)) or (inputs(33));
    layer0_outputs(4155) <= not(inputs(155));
    layer0_outputs(4156) <= not((inputs(6)) or (inputs(47)));
    layer0_outputs(4157) <= not((inputs(142)) or (inputs(88)));
    layer0_outputs(4158) <= not((inputs(22)) xor (inputs(190)));
    layer0_outputs(4159) <= not(inputs(188)) or (inputs(207));
    layer0_outputs(4160) <= '1';
    layer0_outputs(4161) <= (inputs(157)) or (inputs(149));
    layer0_outputs(4162) <= not(inputs(168)) or (inputs(34));
    layer0_outputs(4163) <= '0';
    layer0_outputs(4164) <= not((inputs(63)) xor (inputs(32)));
    layer0_outputs(4165) <= (inputs(189)) and not (inputs(211));
    layer0_outputs(4166) <= not(inputs(166));
    layer0_outputs(4167) <= (inputs(122)) and not (inputs(8));
    layer0_outputs(4168) <= not(inputs(86));
    layer0_outputs(4169) <= not((inputs(176)) or (inputs(138)));
    layer0_outputs(4170) <= (inputs(35)) or (inputs(225));
    layer0_outputs(4171) <= not(inputs(46)) or (inputs(139));
    layer0_outputs(4172) <= not(inputs(224)) or (inputs(13));
    layer0_outputs(4173) <= (inputs(92)) xor (inputs(19));
    layer0_outputs(4174) <= not((inputs(130)) xor (inputs(150)));
    layer0_outputs(4175) <= not((inputs(146)) or (inputs(76)));
    layer0_outputs(4176) <= '1';
    layer0_outputs(4177) <= not(inputs(163));
    layer0_outputs(4178) <= (inputs(215)) or (inputs(207));
    layer0_outputs(4179) <= inputs(124);
    layer0_outputs(4180) <= (inputs(164)) and not (inputs(112));
    layer0_outputs(4181) <= (inputs(56)) and not (inputs(53));
    layer0_outputs(4182) <= inputs(209);
    layer0_outputs(4183) <= not(inputs(254));
    layer0_outputs(4184) <= not((inputs(0)) and (inputs(223)));
    layer0_outputs(4185) <= (inputs(154)) xor (inputs(137));
    layer0_outputs(4186) <= inputs(123);
    layer0_outputs(4187) <= not(inputs(160));
    layer0_outputs(4188) <= inputs(3);
    layer0_outputs(4189) <= not((inputs(149)) or (inputs(117)));
    layer0_outputs(4190) <= not(inputs(56));
    layer0_outputs(4191) <= (inputs(55)) or (inputs(39));
    layer0_outputs(4192) <= (inputs(140)) xor (inputs(127));
    layer0_outputs(4193) <= (inputs(202)) and not (inputs(181));
    layer0_outputs(4194) <= (inputs(238)) or (inputs(20));
    layer0_outputs(4195) <= '0';
    layer0_outputs(4196) <= (inputs(40)) or (inputs(245));
    layer0_outputs(4197) <= not(inputs(232));
    layer0_outputs(4198) <= (inputs(81)) and (inputs(73));
    layer0_outputs(4199) <= inputs(58);
    layer0_outputs(4200) <= not((inputs(72)) xor (inputs(47)));
    layer0_outputs(4201) <= (inputs(204)) or (inputs(32));
    layer0_outputs(4202) <= (inputs(165)) and not (inputs(129));
    layer0_outputs(4203) <= (inputs(228)) and not (inputs(88));
    layer0_outputs(4204) <= (inputs(203)) or (inputs(163));
    layer0_outputs(4205) <= inputs(194);
    layer0_outputs(4206) <= (inputs(82)) or (inputs(196));
    layer0_outputs(4207) <= not(inputs(2));
    layer0_outputs(4208) <= (inputs(224)) or (inputs(234));
    layer0_outputs(4209) <= not(inputs(120)) or (inputs(123));
    layer0_outputs(4210) <= not(inputs(243));
    layer0_outputs(4211) <= not(inputs(52)) or (inputs(134));
    layer0_outputs(4212) <= not(inputs(125));
    layer0_outputs(4213) <= '0';
    layer0_outputs(4214) <= inputs(229);
    layer0_outputs(4215) <= '0';
    layer0_outputs(4216) <= not((inputs(84)) xor (inputs(205)));
    layer0_outputs(4217) <= not(inputs(163));
    layer0_outputs(4218) <= inputs(139);
    layer0_outputs(4219) <= not((inputs(189)) and (inputs(136)));
    layer0_outputs(4220) <= (inputs(89)) xor (inputs(223));
    layer0_outputs(4221) <= inputs(146);
    layer0_outputs(4222) <= (inputs(212)) xor (inputs(157));
    layer0_outputs(4223) <= not((inputs(150)) or (inputs(45)));
    layer0_outputs(4224) <= inputs(90);
    layer0_outputs(4225) <= inputs(110);
    layer0_outputs(4226) <= not(inputs(44));
    layer0_outputs(4227) <= inputs(85);
    layer0_outputs(4228) <= not(inputs(245)) or (inputs(16));
    layer0_outputs(4229) <= not(inputs(237)) or (inputs(157));
    layer0_outputs(4230) <= (inputs(189)) or (inputs(238));
    layer0_outputs(4231) <= not((inputs(205)) and (inputs(202)));
    layer0_outputs(4232) <= not(inputs(99));
    layer0_outputs(4233) <= inputs(8);
    layer0_outputs(4234) <= (inputs(100)) and not (inputs(95));
    layer0_outputs(4235) <= not(inputs(32)) or (inputs(219));
    layer0_outputs(4236) <= (inputs(114)) and not (inputs(232));
    layer0_outputs(4237) <= inputs(76);
    layer0_outputs(4238) <= inputs(183);
    layer0_outputs(4239) <= (inputs(195)) or (inputs(194));
    layer0_outputs(4240) <= inputs(219);
    layer0_outputs(4241) <= not((inputs(190)) xor (inputs(237)));
    layer0_outputs(4242) <= not(inputs(143));
    layer0_outputs(4243) <= not(inputs(162));
    layer0_outputs(4244) <= (inputs(10)) and (inputs(24));
    layer0_outputs(4245) <= (inputs(167)) or (inputs(164));
    layer0_outputs(4246) <= not(inputs(131)) or (inputs(220));
    layer0_outputs(4247) <= not((inputs(185)) xor (inputs(174)));
    layer0_outputs(4248) <= (inputs(215)) or (inputs(202));
    layer0_outputs(4249) <= not((inputs(217)) xor (inputs(124)));
    layer0_outputs(4250) <= inputs(120);
    layer0_outputs(4251) <= not((inputs(28)) xor (inputs(49)));
    layer0_outputs(4252) <= (inputs(55)) and not (inputs(237));
    layer0_outputs(4253) <= not(inputs(29)) or (inputs(158));
    layer0_outputs(4254) <= (inputs(83)) or (inputs(98));
    layer0_outputs(4255) <= (inputs(215)) and not (inputs(158));
    layer0_outputs(4256) <= not(inputs(183)) or (inputs(183));
    layer0_outputs(4257) <= inputs(163);
    layer0_outputs(4258) <= '1';
    layer0_outputs(4259) <= (inputs(5)) and (inputs(66));
    layer0_outputs(4260) <= inputs(23);
    layer0_outputs(4261) <= not(inputs(28));
    layer0_outputs(4262) <= (inputs(34)) and not (inputs(142));
    layer0_outputs(4263) <= not(inputs(168));
    layer0_outputs(4264) <= inputs(84);
    layer0_outputs(4265) <= (inputs(229)) xor (inputs(161));
    layer0_outputs(4266) <= not(inputs(102)) or (inputs(74));
    layer0_outputs(4267) <= inputs(139);
    layer0_outputs(4268) <= not(inputs(118));
    layer0_outputs(4269) <= not((inputs(56)) or (inputs(113)));
    layer0_outputs(4270) <= not((inputs(221)) or (inputs(166)));
    layer0_outputs(4271) <= not((inputs(197)) xor (inputs(150)));
    layer0_outputs(4272) <= not((inputs(63)) or (inputs(25)));
    layer0_outputs(4273) <= not(inputs(34));
    layer0_outputs(4274) <= inputs(253);
    layer0_outputs(4275) <= inputs(153);
    layer0_outputs(4276) <= not(inputs(110)) or (inputs(118));
    layer0_outputs(4277) <= (inputs(230)) or (inputs(158));
    layer0_outputs(4278) <= (inputs(80)) or (inputs(180));
    layer0_outputs(4279) <= inputs(60);
    layer0_outputs(4280) <= not((inputs(209)) or (inputs(206)));
    layer0_outputs(4281) <= '0';
    layer0_outputs(4282) <= (inputs(171)) and not (inputs(174));
    layer0_outputs(4283) <= not((inputs(105)) or (inputs(240)));
    layer0_outputs(4284) <= (inputs(97)) or (inputs(128));
    layer0_outputs(4285) <= not(inputs(170));
    layer0_outputs(4286) <= (inputs(69)) xor (inputs(81));
    layer0_outputs(4287) <= inputs(76);
    layer0_outputs(4288) <= inputs(149);
    layer0_outputs(4289) <= not(inputs(215)) or (inputs(107));
    layer0_outputs(4290) <= (inputs(215)) and (inputs(234));
    layer0_outputs(4291) <= (inputs(36)) xor (inputs(118));
    layer0_outputs(4292) <= inputs(188);
    layer0_outputs(4293) <= not(inputs(12)) or (inputs(240));
    layer0_outputs(4294) <= (inputs(106)) and not (inputs(126));
    layer0_outputs(4295) <= not((inputs(9)) or (inputs(243)));
    layer0_outputs(4296) <= not(inputs(233));
    layer0_outputs(4297) <= not((inputs(78)) xor (inputs(92)));
    layer0_outputs(4298) <= '1';
    layer0_outputs(4299) <= '1';
    layer0_outputs(4300) <= not(inputs(238)) or (inputs(206));
    layer0_outputs(4301) <= not((inputs(189)) or (inputs(209)));
    layer0_outputs(4302) <= (inputs(207)) or (inputs(81));
    layer0_outputs(4303) <= (inputs(207)) and not (inputs(125));
    layer0_outputs(4304) <= inputs(60);
    layer0_outputs(4305) <= inputs(254);
    layer0_outputs(4306) <= inputs(58);
    layer0_outputs(4307) <= '1';
    layer0_outputs(4308) <= (inputs(64)) xor (inputs(40));
    layer0_outputs(4309) <= (inputs(179)) or (inputs(111));
    layer0_outputs(4310) <= not(inputs(205));
    layer0_outputs(4311) <= (inputs(186)) or (inputs(165));
    layer0_outputs(4312) <= not(inputs(106));
    layer0_outputs(4313) <= (inputs(175)) or (inputs(228));
    layer0_outputs(4314) <= '0';
    layer0_outputs(4315) <= not(inputs(13)) or (inputs(184));
    layer0_outputs(4316) <= not(inputs(35));
    layer0_outputs(4317) <= inputs(21);
    layer0_outputs(4318) <= not((inputs(185)) and (inputs(166)));
    layer0_outputs(4319) <= not(inputs(194)) or (inputs(168));
    layer0_outputs(4320) <= not(inputs(51));
    layer0_outputs(4321) <= not(inputs(212));
    layer0_outputs(4322) <= not(inputs(133)) or (inputs(49));
    layer0_outputs(4323) <= (inputs(132)) and (inputs(155));
    layer0_outputs(4324) <= not(inputs(168));
    layer0_outputs(4325) <= inputs(72);
    layer0_outputs(4326) <= not(inputs(254)) or (inputs(178));
    layer0_outputs(4327) <= not((inputs(105)) xor (inputs(165)));
    layer0_outputs(4328) <= not(inputs(111));
    layer0_outputs(4329) <= not((inputs(243)) or (inputs(33)));
    layer0_outputs(4330) <= (inputs(106)) xor (inputs(16));
    layer0_outputs(4331) <= not((inputs(48)) or (inputs(235)));
    layer0_outputs(4332) <= (inputs(201)) and not (inputs(142));
    layer0_outputs(4333) <= (inputs(86)) or (inputs(3));
    layer0_outputs(4334) <= not((inputs(80)) xor (inputs(51)));
    layer0_outputs(4335) <= (inputs(38)) xor (inputs(71));
    layer0_outputs(4336) <= not((inputs(178)) or (inputs(252)));
    layer0_outputs(4337) <= not((inputs(14)) or (inputs(41)));
    layer0_outputs(4338) <= not(inputs(178));
    layer0_outputs(4339) <= not(inputs(33));
    layer0_outputs(4340) <= not(inputs(45)) or (inputs(252));
    layer0_outputs(4341) <= (inputs(173)) xor (inputs(19));
    layer0_outputs(4342) <= inputs(110);
    layer0_outputs(4343) <= not(inputs(245));
    layer0_outputs(4344) <= not(inputs(192));
    layer0_outputs(4345) <= not((inputs(162)) xor (inputs(158)));
    layer0_outputs(4346) <= not((inputs(211)) or (inputs(198)));
    layer0_outputs(4347) <= inputs(101);
    layer0_outputs(4348) <= inputs(163);
    layer0_outputs(4349) <= (inputs(49)) or (inputs(26));
    layer0_outputs(4350) <= inputs(215);
    layer0_outputs(4351) <= (inputs(129)) xor (inputs(109));
    layer0_outputs(4352) <= not(inputs(25));
    layer0_outputs(4353) <= (inputs(84)) xor (inputs(82));
    layer0_outputs(4354) <= not((inputs(237)) and (inputs(58)));
    layer0_outputs(4355) <= not(inputs(66)) or (inputs(224));
    layer0_outputs(4356) <= not((inputs(94)) xor (inputs(89)));
    layer0_outputs(4357) <= '1';
    layer0_outputs(4358) <= (inputs(121)) and not (inputs(157));
    layer0_outputs(4359) <= not(inputs(35));
    layer0_outputs(4360) <= inputs(88);
    layer0_outputs(4361) <= (inputs(83)) and not (inputs(2));
    layer0_outputs(4362) <= inputs(78);
    layer0_outputs(4363) <= inputs(162);
    layer0_outputs(4364) <= not(inputs(124)) or (inputs(144));
    layer0_outputs(4365) <= inputs(189);
    layer0_outputs(4366) <= '0';
    layer0_outputs(4367) <= '1';
    layer0_outputs(4368) <= not(inputs(10));
    layer0_outputs(4369) <= not(inputs(12)) or (inputs(80));
    layer0_outputs(4370) <= not(inputs(121));
    layer0_outputs(4371) <= (inputs(149)) and not (inputs(229));
    layer0_outputs(4372) <= (inputs(78)) or (inputs(155));
    layer0_outputs(4373) <= (inputs(66)) and not (inputs(215));
    layer0_outputs(4374) <= inputs(180);
    layer0_outputs(4375) <= not((inputs(39)) or (inputs(22)));
    layer0_outputs(4376) <= not(inputs(59));
    layer0_outputs(4377) <= not((inputs(144)) or (inputs(133)));
    layer0_outputs(4378) <= not(inputs(115));
    layer0_outputs(4379) <= (inputs(194)) and not (inputs(188));
    layer0_outputs(4380) <= (inputs(168)) or (inputs(137));
    layer0_outputs(4381) <= not(inputs(137)) or (inputs(142));
    layer0_outputs(4382) <= inputs(165);
    layer0_outputs(4383) <= (inputs(206)) xor (inputs(108));
    layer0_outputs(4384) <= (inputs(120)) or (inputs(84));
    layer0_outputs(4385) <= not((inputs(129)) and (inputs(96)));
    layer0_outputs(4386) <= (inputs(48)) or (inputs(52));
    layer0_outputs(4387) <= (inputs(255)) or (inputs(193));
    layer0_outputs(4388) <= not(inputs(77)) or (inputs(178));
    layer0_outputs(4389) <= (inputs(175)) and not (inputs(142));
    layer0_outputs(4390) <= not((inputs(83)) or (inputs(177)));
    layer0_outputs(4391) <= not(inputs(172)) or (inputs(152));
    layer0_outputs(4392) <= (inputs(98)) and (inputs(42));
    layer0_outputs(4393) <= inputs(153);
    layer0_outputs(4394) <= (inputs(117)) or (inputs(248));
    layer0_outputs(4395) <= (inputs(215)) and not (inputs(71));
    layer0_outputs(4396) <= (inputs(54)) and not (inputs(149));
    layer0_outputs(4397) <= not((inputs(144)) xor (inputs(132)));
    layer0_outputs(4398) <= not((inputs(59)) or (inputs(77)));
    layer0_outputs(4399) <= not((inputs(247)) xor (inputs(143)));
    layer0_outputs(4400) <= '0';
    layer0_outputs(4401) <= not(inputs(1));
    layer0_outputs(4402) <= not((inputs(20)) xor (inputs(68)));
    layer0_outputs(4403) <= (inputs(128)) and not (inputs(70));
    layer0_outputs(4404) <= (inputs(138)) and not (inputs(27));
    layer0_outputs(4405) <= inputs(211);
    layer0_outputs(4406) <= '1';
    layer0_outputs(4407) <= not(inputs(235));
    layer0_outputs(4408) <= (inputs(214)) and not (inputs(73));
    layer0_outputs(4409) <= not((inputs(26)) or (inputs(94)));
    layer0_outputs(4410) <= (inputs(171)) and not (inputs(14));
    layer0_outputs(4411) <= not(inputs(16));
    layer0_outputs(4412) <= inputs(19);
    layer0_outputs(4413) <= inputs(246);
    layer0_outputs(4414) <= (inputs(85)) or (inputs(55));
    layer0_outputs(4415) <= (inputs(222)) and not (inputs(108));
    layer0_outputs(4416) <= (inputs(234)) and not (inputs(45));
    layer0_outputs(4417) <= inputs(109);
    layer0_outputs(4418) <= not((inputs(166)) xor (inputs(247)));
    layer0_outputs(4419) <= (inputs(33)) or (inputs(199));
    layer0_outputs(4420) <= inputs(215);
    layer0_outputs(4421) <= (inputs(106)) or (inputs(60));
    layer0_outputs(4422) <= not(inputs(242)) or (inputs(200));
    layer0_outputs(4423) <= (inputs(128)) and not (inputs(112));
    layer0_outputs(4424) <= inputs(98);
    layer0_outputs(4425) <= not((inputs(134)) xor (inputs(161)));
    layer0_outputs(4426) <= inputs(6);
    layer0_outputs(4427) <= not((inputs(1)) or (inputs(65)));
    layer0_outputs(4428) <= not(inputs(40));
    layer0_outputs(4429) <= inputs(233);
    layer0_outputs(4430) <= (inputs(75)) and (inputs(103));
    layer0_outputs(4431) <= not((inputs(89)) xor (inputs(42)));
    layer0_outputs(4432) <= inputs(127);
    layer0_outputs(4433) <= not((inputs(217)) xor (inputs(184)));
    layer0_outputs(4434) <= not(inputs(151));
    layer0_outputs(4435) <= (inputs(143)) or (inputs(89));
    layer0_outputs(4436) <= (inputs(5)) and not (inputs(144));
    layer0_outputs(4437) <= not(inputs(246)) or (inputs(178));
    layer0_outputs(4438) <= inputs(68);
    layer0_outputs(4439) <= (inputs(221)) and (inputs(144));
    layer0_outputs(4440) <= inputs(92);
    layer0_outputs(4441) <= not((inputs(197)) xor (inputs(191)));
    layer0_outputs(4442) <= inputs(114);
    layer0_outputs(4443) <= (inputs(148)) and not (inputs(152));
    layer0_outputs(4444) <= not((inputs(28)) xor (inputs(176)));
    layer0_outputs(4445) <= not(inputs(64));
    layer0_outputs(4446) <= inputs(145);
    layer0_outputs(4447) <= inputs(123);
    layer0_outputs(4448) <= not(inputs(131));
    layer0_outputs(4449) <= not((inputs(136)) or (inputs(168)));
    layer0_outputs(4450) <= (inputs(189)) and not (inputs(33));
    layer0_outputs(4451) <= (inputs(213)) or (inputs(229));
    layer0_outputs(4452) <= not((inputs(202)) or (inputs(174)));
    layer0_outputs(4453) <= inputs(89);
    layer0_outputs(4454) <= not(inputs(176)) or (inputs(4));
    layer0_outputs(4455) <= (inputs(251)) or (inputs(198));
    layer0_outputs(4456) <= not(inputs(135)) or (inputs(128));
    layer0_outputs(4457) <= not(inputs(122)) or (inputs(253));
    layer0_outputs(4458) <= not(inputs(116));
    layer0_outputs(4459) <= (inputs(24)) or (inputs(111));
    layer0_outputs(4460) <= (inputs(58)) xor (inputs(40));
    layer0_outputs(4461) <= (inputs(158)) xor (inputs(100));
    layer0_outputs(4462) <= not((inputs(10)) or (inputs(97)));
    layer0_outputs(4463) <= (inputs(7)) and not (inputs(145));
    layer0_outputs(4464) <= (inputs(104)) xor (inputs(123));
    layer0_outputs(4465) <= (inputs(58)) and not (inputs(216));
    layer0_outputs(4466) <= inputs(122);
    layer0_outputs(4467) <= not(inputs(132)) or (inputs(48));
    layer0_outputs(4468) <= (inputs(8)) and (inputs(25));
    layer0_outputs(4469) <= not(inputs(39)) or (inputs(241));
    layer0_outputs(4470) <= (inputs(129)) and not (inputs(239));
    layer0_outputs(4471) <= (inputs(178)) xor (inputs(112));
    layer0_outputs(4472) <= not((inputs(130)) or (inputs(186)));
    layer0_outputs(4473) <= not(inputs(143)) or (inputs(171));
    layer0_outputs(4474) <= not(inputs(232)) or (inputs(242));
    layer0_outputs(4475) <= not((inputs(71)) xor (inputs(203)));
    layer0_outputs(4476) <= (inputs(132)) and not (inputs(13));
    layer0_outputs(4477) <= not(inputs(99));
    layer0_outputs(4478) <= not((inputs(130)) or (inputs(132)));
    layer0_outputs(4479) <= (inputs(232)) and not (inputs(35));
    layer0_outputs(4480) <= not(inputs(79));
    layer0_outputs(4481) <= (inputs(42)) and not (inputs(170));
    layer0_outputs(4482) <= not(inputs(167)) or (inputs(46));
    layer0_outputs(4483) <= not(inputs(232));
    layer0_outputs(4484) <= not(inputs(174));
    layer0_outputs(4485) <= not(inputs(7)) or (inputs(0));
    layer0_outputs(4486) <= (inputs(118)) xor (inputs(131));
    layer0_outputs(4487) <= inputs(10);
    layer0_outputs(4488) <= not(inputs(6)) or (inputs(221));
    layer0_outputs(4489) <= not(inputs(20)) or (inputs(153));
    layer0_outputs(4490) <= (inputs(81)) xor (inputs(79));
    layer0_outputs(4491) <= inputs(94);
    layer0_outputs(4492) <= not((inputs(162)) or (inputs(7)));
    layer0_outputs(4493) <= not((inputs(109)) or (inputs(23)));
    layer0_outputs(4494) <= not((inputs(64)) xor (inputs(61)));
    layer0_outputs(4495) <= (inputs(86)) and not (inputs(249));
    layer0_outputs(4496) <= (inputs(216)) or (inputs(164));
    layer0_outputs(4497) <= (inputs(13)) or (inputs(96));
    layer0_outputs(4498) <= not(inputs(165)) or (inputs(84));
    layer0_outputs(4499) <= not(inputs(89));
    layer0_outputs(4500) <= not(inputs(8)) or (inputs(1));
    layer0_outputs(4501) <= not(inputs(63));
    layer0_outputs(4502) <= not(inputs(88)) or (inputs(227));
    layer0_outputs(4503) <= not((inputs(24)) or (inputs(1)));
    layer0_outputs(4504) <= (inputs(181)) xor (inputs(179));
    layer0_outputs(4505) <= not((inputs(225)) and (inputs(179)));
    layer0_outputs(4506) <= inputs(114);
    layer0_outputs(4507) <= (inputs(24)) and not (inputs(178));
    layer0_outputs(4508) <= not(inputs(174));
    layer0_outputs(4509) <= '0';
    layer0_outputs(4510) <= not(inputs(13)) or (inputs(151));
    layer0_outputs(4511) <= not(inputs(132)) or (inputs(45));
    layer0_outputs(4512) <= not(inputs(230));
    layer0_outputs(4513) <= not(inputs(138)) or (inputs(140));
    layer0_outputs(4514) <= not((inputs(68)) or (inputs(188)));
    layer0_outputs(4515) <= (inputs(176)) or (inputs(14));
    layer0_outputs(4516) <= not(inputs(148));
    layer0_outputs(4517) <= inputs(17);
    layer0_outputs(4518) <= not((inputs(255)) or (inputs(177)));
    layer0_outputs(4519) <= not(inputs(152)) or (inputs(203));
    layer0_outputs(4520) <= (inputs(202)) and not (inputs(108));
    layer0_outputs(4521) <= not((inputs(237)) or (inputs(164)));
    layer0_outputs(4522) <= '0';
    layer0_outputs(4523) <= not(inputs(124));
    layer0_outputs(4524) <= not(inputs(234));
    layer0_outputs(4525) <= not((inputs(126)) xor (inputs(243)));
    layer0_outputs(4526) <= not((inputs(10)) or (inputs(91)));
    layer0_outputs(4527) <= (inputs(24)) and not (inputs(115));
    layer0_outputs(4528) <= (inputs(18)) xor (inputs(91));
    layer0_outputs(4529) <= inputs(153);
    layer0_outputs(4530) <= not((inputs(168)) and (inputs(19)));
    layer0_outputs(4531) <= inputs(20);
    layer0_outputs(4532) <= not((inputs(164)) or (inputs(201)));
    layer0_outputs(4533) <= (inputs(184)) xor (inputs(83));
    layer0_outputs(4534) <= (inputs(144)) or (inputs(142));
    layer0_outputs(4535) <= not((inputs(194)) or (inputs(196)));
    layer0_outputs(4536) <= (inputs(25)) xor (inputs(71));
    layer0_outputs(4537) <= not(inputs(60));
    layer0_outputs(4538) <= not(inputs(12)) or (inputs(95));
    layer0_outputs(4539) <= not((inputs(170)) or (inputs(206)));
    layer0_outputs(4540) <= (inputs(204)) or (inputs(249));
    layer0_outputs(4541) <= not(inputs(155)) or (inputs(109));
    layer0_outputs(4542) <= not(inputs(122));
    layer0_outputs(4543) <= not((inputs(203)) and (inputs(4)));
    layer0_outputs(4544) <= (inputs(117)) or (inputs(148));
    layer0_outputs(4545) <= not(inputs(50));
    layer0_outputs(4546) <= not(inputs(209));
    layer0_outputs(4547) <= (inputs(50)) or (inputs(29));
    layer0_outputs(4548) <= '1';
    layer0_outputs(4549) <= not(inputs(104));
    layer0_outputs(4550) <= not((inputs(41)) and (inputs(228)));
    layer0_outputs(4551) <= inputs(36);
    layer0_outputs(4552) <= (inputs(104)) and not (inputs(54));
    layer0_outputs(4553) <= '0';
    layer0_outputs(4554) <= inputs(111);
    layer0_outputs(4555) <= not((inputs(252)) xor (inputs(142)));
    layer0_outputs(4556) <= (inputs(252)) or (inputs(176));
    layer0_outputs(4557) <= (inputs(138)) or (inputs(77));
    layer0_outputs(4558) <= not(inputs(122));
    layer0_outputs(4559) <= not(inputs(86));
    layer0_outputs(4560) <= not(inputs(40));
    layer0_outputs(4561) <= (inputs(83)) and (inputs(16));
    layer0_outputs(4562) <= (inputs(24)) and (inputs(26));
    layer0_outputs(4563) <= inputs(196);
    layer0_outputs(4564) <= not(inputs(148));
    layer0_outputs(4565) <= inputs(51);
    layer0_outputs(4566) <= not(inputs(229));
    layer0_outputs(4567) <= (inputs(214)) and not (inputs(156));
    layer0_outputs(4568) <= not(inputs(53)) or (inputs(192));
    layer0_outputs(4569) <= inputs(169);
    layer0_outputs(4570) <= not(inputs(187));
    layer0_outputs(4571) <= (inputs(156)) and not (inputs(12));
    layer0_outputs(4572) <= (inputs(106)) or (inputs(205));
    layer0_outputs(4573) <= (inputs(246)) xor (inputs(214));
    layer0_outputs(4574) <= not(inputs(214));
    layer0_outputs(4575) <= not(inputs(248));
    layer0_outputs(4576) <= (inputs(190)) and not (inputs(225));
    layer0_outputs(4577) <= inputs(100);
    layer0_outputs(4578) <= inputs(237);
    layer0_outputs(4579) <= not(inputs(122));
    layer0_outputs(4580) <= inputs(39);
    layer0_outputs(4581) <= (inputs(171)) and not (inputs(37));
    layer0_outputs(4582) <= (inputs(163)) or (inputs(178));
    layer0_outputs(4583) <= (inputs(143)) or (inputs(12));
    layer0_outputs(4584) <= not(inputs(179));
    layer0_outputs(4585) <= (inputs(121)) or (inputs(91));
    layer0_outputs(4586) <= (inputs(125)) xor (inputs(204));
    layer0_outputs(4587) <= (inputs(5)) or (inputs(41));
    layer0_outputs(4588) <= not(inputs(175));
    layer0_outputs(4589) <= (inputs(127)) xor (inputs(0));
    layer0_outputs(4590) <= (inputs(64)) or (inputs(75));
    layer0_outputs(4591) <= not((inputs(236)) xor (inputs(172)));
    layer0_outputs(4592) <= not(inputs(243)) or (inputs(56));
    layer0_outputs(4593) <= (inputs(220)) or (inputs(105));
    layer0_outputs(4594) <= inputs(21);
    layer0_outputs(4595) <= inputs(75);
    layer0_outputs(4596) <= not((inputs(27)) or (inputs(208)));
    layer0_outputs(4597) <= not(inputs(59)) or (inputs(205));
    layer0_outputs(4598) <= (inputs(119)) or (inputs(71));
    layer0_outputs(4599) <= not((inputs(162)) or (inputs(144)));
    layer0_outputs(4600) <= not(inputs(44));
    layer0_outputs(4601) <= not(inputs(127));
    layer0_outputs(4602) <= not((inputs(40)) or (inputs(175)));
    layer0_outputs(4603) <= inputs(233);
    layer0_outputs(4604) <= inputs(98);
    layer0_outputs(4605) <= not(inputs(24)) or (inputs(166));
    layer0_outputs(4606) <= not(inputs(246));
    layer0_outputs(4607) <= inputs(188);
    layer0_outputs(4608) <= '1';
    layer0_outputs(4609) <= not(inputs(139)) or (inputs(243));
    layer0_outputs(4610) <= not((inputs(211)) xor (inputs(16)));
    layer0_outputs(4611) <= not((inputs(199)) or (inputs(215)));
    layer0_outputs(4612) <= not((inputs(109)) or (inputs(82)));
    layer0_outputs(4613) <= not((inputs(74)) or (inputs(33)));
    layer0_outputs(4614) <= '1';
    layer0_outputs(4615) <= (inputs(181)) xor (inputs(138));
    layer0_outputs(4616) <= (inputs(227)) xor (inputs(134));
    layer0_outputs(4617) <= not(inputs(112)) or (inputs(30));
    layer0_outputs(4618) <= (inputs(145)) or (inputs(248));
    layer0_outputs(4619) <= (inputs(177)) or (inputs(247));
    layer0_outputs(4620) <= (inputs(30)) or (inputs(56));
    layer0_outputs(4621) <= not((inputs(161)) xor (inputs(218)));
    layer0_outputs(4622) <= '1';
    layer0_outputs(4623) <= (inputs(11)) or (inputs(13));
    layer0_outputs(4624) <= inputs(179);
    layer0_outputs(4625) <= inputs(184);
    layer0_outputs(4626) <= not((inputs(3)) and (inputs(157)));
    layer0_outputs(4627) <= not(inputs(154));
    layer0_outputs(4628) <= not(inputs(160));
    layer0_outputs(4629) <= not((inputs(76)) or (inputs(97)));
    layer0_outputs(4630) <= not(inputs(247)) or (inputs(12));
    layer0_outputs(4631) <= inputs(46);
    layer0_outputs(4632) <= (inputs(186)) and (inputs(179));
    layer0_outputs(4633) <= (inputs(158)) or (inputs(4));
    layer0_outputs(4634) <= (inputs(154)) and not (inputs(248));
    layer0_outputs(4635) <= not(inputs(102));
    layer0_outputs(4636) <= not((inputs(16)) or (inputs(10)));
    layer0_outputs(4637) <= not(inputs(102)) or (inputs(17));
    layer0_outputs(4638) <= '0';
    layer0_outputs(4639) <= not(inputs(220)) or (inputs(196));
    layer0_outputs(4640) <= not(inputs(29));
    layer0_outputs(4641) <= not(inputs(128)) or (inputs(3));
    layer0_outputs(4642) <= not(inputs(115)) or (inputs(31));
    layer0_outputs(4643) <= (inputs(15)) and not (inputs(20));
    layer0_outputs(4644) <= not(inputs(54)) or (inputs(180));
    layer0_outputs(4645) <= inputs(91);
    layer0_outputs(4646) <= inputs(121);
    layer0_outputs(4647) <= not((inputs(128)) xor (inputs(82)));
    layer0_outputs(4648) <= '1';
    layer0_outputs(4649) <= not((inputs(207)) xor (inputs(250)));
    layer0_outputs(4650) <= (inputs(14)) xor (inputs(47));
    layer0_outputs(4651) <= not(inputs(82));
    layer0_outputs(4652) <= not((inputs(246)) and (inputs(251)));
    layer0_outputs(4653) <= not(inputs(229));
    layer0_outputs(4654) <= inputs(5);
    layer0_outputs(4655) <= (inputs(96)) and (inputs(166));
    layer0_outputs(4656) <= (inputs(71)) and not (inputs(177));
    layer0_outputs(4657) <= not(inputs(79));
    layer0_outputs(4658) <= inputs(162);
    layer0_outputs(4659) <= not(inputs(80));
    layer0_outputs(4660) <= not(inputs(150)) or (inputs(47));
    layer0_outputs(4661) <= not(inputs(181));
    layer0_outputs(4662) <= inputs(218);
    layer0_outputs(4663) <= (inputs(103)) and not (inputs(103));
    layer0_outputs(4664) <= not((inputs(166)) and (inputs(43)));
    layer0_outputs(4665) <= (inputs(8)) or (inputs(91));
    layer0_outputs(4666) <= '1';
    layer0_outputs(4667) <= not((inputs(255)) xor (inputs(117)));
    layer0_outputs(4668) <= (inputs(100)) xor (inputs(71));
    layer0_outputs(4669) <= not(inputs(103));
    layer0_outputs(4670) <= (inputs(48)) and not (inputs(242));
    layer0_outputs(4671) <= not((inputs(200)) and (inputs(118)));
    layer0_outputs(4672) <= not((inputs(192)) or (inputs(200)));
    layer0_outputs(4673) <= not(inputs(142)) or (inputs(79));
    layer0_outputs(4674) <= not(inputs(55)) or (inputs(130));
    layer0_outputs(4675) <= (inputs(231)) and (inputs(23));
    layer0_outputs(4676) <= (inputs(147)) or (inputs(212));
    layer0_outputs(4677) <= inputs(55);
    layer0_outputs(4678) <= '1';
    layer0_outputs(4679) <= (inputs(57)) and not (inputs(187));
    layer0_outputs(4680) <= not(inputs(136)) or (inputs(99));
    layer0_outputs(4681) <= (inputs(252)) or (inputs(237));
    layer0_outputs(4682) <= (inputs(247)) xor (inputs(67));
    layer0_outputs(4683) <= not(inputs(92));
    layer0_outputs(4684) <= not(inputs(121)) or (inputs(175));
    layer0_outputs(4685) <= not((inputs(152)) xor (inputs(49)));
    layer0_outputs(4686) <= not((inputs(126)) xor (inputs(108)));
    layer0_outputs(4687) <= inputs(93);
    layer0_outputs(4688) <= not((inputs(225)) and (inputs(16)));
    layer0_outputs(4689) <= not(inputs(163)) or (inputs(241));
    layer0_outputs(4690) <= '0';
    layer0_outputs(4691) <= (inputs(250)) or (inputs(139));
    layer0_outputs(4692) <= (inputs(121)) xor (inputs(146));
    layer0_outputs(4693) <= not(inputs(117)) or (inputs(146));
    layer0_outputs(4694) <= not(inputs(60));
    layer0_outputs(4695) <= not((inputs(226)) or (inputs(239)));
    layer0_outputs(4696) <= (inputs(230)) or (inputs(32));
    layer0_outputs(4697) <= not((inputs(25)) and (inputs(22)));
    layer0_outputs(4698) <= not(inputs(106));
    layer0_outputs(4699) <= inputs(199);
    layer0_outputs(4700) <= (inputs(90)) or (inputs(74));
    layer0_outputs(4701) <= not(inputs(246));
    layer0_outputs(4702) <= not((inputs(215)) or (inputs(170)));
    layer0_outputs(4703) <= not(inputs(23)) or (inputs(160));
    layer0_outputs(4704) <= not((inputs(192)) or (inputs(176)));
    layer0_outputs(4705) <= not(inputs(62));
    layer0_outputs(4706) <= (inputs(128)) and (inputs(40));
    layer0_outputs(4707) <= not(inputs(167));
    layer0_outputs(4708) <= not(inputs(131)) or (inputs(66));
    layer0_outputs(4709) <= not(inputs(136));
    layer0_outputs(4710) <= inputs(216);
    layer0_outputs(4711) <= inputs(231);
    layer0_outputs(4712) <= (inputs(44)) and not (inputs(91));
    layer0_outputs(4713) <= (inputs(72)) and not (inputs(117));
    layer0_outputs(4714) <= (inputs(51)) or (inputs(170));
    layer0_outputs(4715) <= inputs(37);
    layer0_outputs(4716) <= (inputs(233)) xor (inputs(61));
    layer0_outputs(4717) <= (inputs(150)) and (inputs(219));
    layer0_outputs(4718) <= not(inputs(54));
    layer0_outputs(4719) <= (inputs(186)) or (inputs(98));
    layer0_outputs(4720) <= not((inputs(64)) xor (inputs(69)));
    layer0_outputs(4721) <= not((inputs(242)) and (inputs(229)));
    layer0_outputs(4722) <= (inputs(194)) and not (inputs(94));
    layer0_outputs(4723) <= not(inputs(109)) or (inputs(30));
    layer0_outputs(4724) <= not(inputs(57)) or (inputs(102));
    layer0_outputs(4725) <= not((inputs(97)) and (inputs(210)));
    layer0_outputs(4726) <= '1';
    layer0_outputs(4727) <= not((inputs(243)) xor (inputs(243)));
    layer0_outputs(4728) <= (inputs(40)) or (inputs(226));
    layer0_outputs(4729) <= inputs(204);
    layer0_outputs(4730) <= not(inputs(73));
    layer0_outputs(4731) <= not(inputs(21));
    layer0_outputs(4732) <= (inputs(114)) xor (inputs(47));
    layer0_outputs(4733) <= '1';
    layer0_outputs(4734) <= (inputs(40)) and not (inputs(68));
    layer0_outputs(4735) <= inputs(59);
    layer0_outputs(4736) <= not(inputs(208)) or (inputs(13));
    layer0_outputs(4737) <= not(inputs(87));
    layer0_outputs(4738) <= inputs(202);
    layer0_outputs(4739) <= (inputs(252)) and not (inputs(162));
    layer0_outputs(4740) <= (inputs(64)) and (inputs(3));
    layer0_outputs(4741) <= not(inputs(220));
    layer0_outputs(4742) <= not(inputs(148));
    layer0_outputs(4743) <= (inputs(221)) and not (inputs(240));
    layer0_outputs(4744) <= not((inputs(4)) xor (inputs(125)));
    layer0_outputs(4745) <= not(inputs(247));
    layer0_outputs(4746) <= (inputs(203)) or (inputs(219));
    layer0_outputs(4747) <= not((inputs(82)) or (inputs(111)));
    layer0_outputs(4748) <= (inputs(158)) or (inputs(160));
    layer0_outputs(4749) <= not(inputs(169)) or (inputs(154));
    layer0_outputs(4750) <= (inputs(84)) or (inputs(132));
    layer0_outputs(4751) <= not(inputs(110)) or (inputs(239));
    layer0_outputs(4752) <= not(inputs(37)) or (inputs(206));
    layer0_outputs(4753) <= inputs(7);
    layer0_outputs(4754) <= not((inputs(138)) or (inputs(87)));
    layer0_outputs(4755) <= not(inputs(131));
    layer0_outputs(4756) <= '1';
    layer0_outputs(4757) <= inputs(114);
    layer0_outputs(4758) <= not(inputs(109)) or (inputs(39));
    layer0_outputs(4759) <= inputs(8);
    layer0_outputs(4760) <= not(inputs(199));
    layer0_outputs(4761) <= (inputs(167)) xor (inputs(11));
    layer0_outputs(4762) <= '0';
    layer0_outputs(4763) <= not(inputs(250)) or (inputs(126));
    layer0_outputs(4764) <= not(inputs(227)) or (inputs(77));
    layer0_outputs(4765) <= (inputs(2)) or (inputs(223));
    layer0_outputs(4766) <= inputs(3);
    layer0_outputs(4767) <= (inputs(225)) and not (inputs(239));
    layer0_outputs(4768) <= (inputs(48)) and not (inputs(49));
    layer0_outputs(4769) <= (inputs(140)) or (inputs(162));
    layer0_outputs(4770) <= not(inputs(73));
    layer0_outputs(4771) <= (inputs(116)) and not (inputs(193));
    layer0_outputs(4772) <= not(inputs(25));
    layer0_outputs(4773) <= not(inputs(240));
    layer0_outputs(4774) <= (inputs(33)) and not (inputs(161));
    layer0_outputs(4775) <= not(inputs(173));
    layer0_outputs(4776) <= not(inputs(98));
    layer0_outputs(4777) <= (inputs(26)) and not (inputs(243));
    layer0_outputs(4778) <= not((inputs(35)) or (inputs(236)));
    layer0_outputs(4779) <= (inputs(27)) and (inputs(26));
    layer0_outputs(4780) <= '0';
    layer0_outputs(4781) <= not((inputs(47)) or (inputs(104)));
    layer0_outputs(4782) <= (inputs(190)) or (inputs(88));
    layer0_outputs(4783) <= '1';
    layer0_outputs(4784) <= (inputs(3)) xor (inputs(63));
    layer0_outputs(4785) <= not(inputs(185)) or (inputs(14));
    layer0_outputs(4786) <= '0';
    layer0_outputs(4787) <= '1';
    layer0_outputs(4788) <= (inputs(197)) or (inputs(156));
    layer0_outputs(4789) <= (inputs(245)) xor (inputs(201));
    layer0_outputs(4790) <= inputs(96);
    layer0_outputs(4791) <= not(inputs(101));
    layer0_outputs(4792) <= not((inputs(21)) and (inputs(25)));
    layer0_outputs(4793) <= not(inputs(69));
    layer0_outputs(4794) <= (inputs(191)) xor (inputs(149));
    layer0_outputs(4795) <= inputs(103);
    layer0_outputs(4796) <= (inputs(236)) or (inputs(109));
    layer0_outputs(4797) <= (inputs(146)) xor (inputs(25));
    layer0_outputs(4798) <= (inputs(8)) and not (inputs(164));
    layer0_outputs(4799) <= (inputs(159)) xor (inputs(0));
    layer0_outputs(4800) <= (inputs(53)) and not (inputs(118));
    layer0_outputs(4801) <= not((inputs(104)) or (inputs(203)));
    layer0_outputs(4802) <= not(inputs(117)) or (inputs(237));
    layer0_outputs(4803) <= inputs(38);
    layer0_outputs(4804) <= (inputs(217)) or (inputs(129));
    layer0_outputs(4805) <= not(inputs(8));
    layer0_outputs(4806) <= (inputs(48)) and not (inputs(255));
    layer0_outputs(4807) <= not(inputs(147));
    layer0_outputs(4808) <= not(inputs(38));
    layer0_outputs(4809) <= (inputs(184)) and not (inputs(201));
    layer0_outputs(4810) <= not(inputs(135)) or (inputs(1));
    layer0_outputs(4811) <= not(inputs(166));
    layer0_outputs(4812) <= not(inputs(110));
    layer0_outputs(4813) <= '1';
    layer0_outputs(4814) <= (inputs(61)) or (inputs(50));
    layer0_outputs(4815) <= (inputs(42)) and not (inputs(3));
    layer0_outputs(4816) <= not(inputs(191));
    layer0_outputs(4817) <= inputs(180);
    layer0_outputs(4818) <= not((inputs(185)) and (inputs(217)));
    layer0_outputs(4819) <= (inputs(102)) and (inputs(157));
    layer0_outputs(4820) <= '1';
    layer0_outputs(4821) <= not(inputs(234));
    layer0_outputs(4822) <= inputs(239);
    layer0_outputs(4823) <= not(inputs(132)) or (inputs(157));
    layer0_outputs(4824) <= (inputs(216)) and (inputs(199));
    layer0_outputs(4825) <= inputs(132);
    layer0_outputs(4826) <= inputs(235);
    layer0_outputs(4827) <= not(inputs(237)) or (inputs(250));
    layer0_outputs(4828) <= (inputs(184)) and not (inputs(67));
    layer0_outputs(4829) <= not(inputs(206)) or (inputs(184));
    layer0_outputs(4830) <= (inputs(209)) and not (inputs(65));
    layer0_outputs(4831) <= not(inputs(105));
    layer0_outputs(4832) <= not(inputs(147)) or (inputs(57));
    layer0_outputs(4833) <= not(inputs(80));
    layer0_outputs(4834) <= (inputs(201)) or (inputs(37));
    layer0_outputs(4835) <= not((inputs(67)) xor (inputs(221)));
    layer0_outputs(4836) <= not((inputs(21)) xor (inputs(229)));
    layer0_outputs(4837) <= inputs(165);
    layer0_outputs(4838) <= '1';
    layer0_outputs(4839) <= (inputs(179)) or (inputs(17));
    layer0_outputs(4840) <= inputs(105);
    layer0_outputs(4841) <= not((inputs(85)) or (inputs(147)));
    layer0_outputs(4842) <= not(inputs(157));
    layer0_outputs(4843) <= not(inputs(47));
    layer0_outputs(4844) <= not(inputs(80));
    layer0_outputs(4845) <= (inputs(11)) and not (inputs(202));
    layer0_outputs(4846) <= '1';
    layer0_outputs(4847) <= inputs(4);
    layer0_outputs(4848) <= '1';
    layer0_outputs(4849) <= not((inputs(31)) xor (inputs(159)));
    layer0_outputs(4850) <= not(inputs(83)) or (inputs(184));
    layer0_outputs(4851) <= (inputs(239)) xor (inputs(144));
    layer0_outputs(4852) <= '1';
    layer0_outputs(4853) <= not(inputs(183)) or (inputs(177));
    layer0_outputs(4854) <= (inputs(47)) or (inputs(224));
    layer0_outputs(4855) <= (inputs(49)) and (inputs(114));
    layer0_outputs(4856) <= not((inputs(113)) or (inputs(114)));
    layer0_outputs(4857) <= not(inputs(74));
    layer0_outputs(4858) <= (inputs(7)) and not (inputs(143));
    layer0_outputs(4859) <= not((inputs(163)) or (inputs(223)));
    layer0_outputs(4860) <= '0';
    layer0_outputs(4861) <= (inputs(109)) or (inputs(185));
    layer0_outputs(4862) <= not(inputs(46));
    layer0_outputs(4863) <= not(inputs(18)) or (inputs(96));
    layer0_outputs(4864) <= not(inputs(134));
    layer0_outputs(4865) <= not((inputs(106)) xor (inputs(204)));
    layer0_outputs(4866) <= not((inputs(127)) xor (inputs(193)));
    layer0_outputs(4867) <= (inputs(179)) or (inputs(234));
    layer0_outputs(4868) <= not((inputs(154)) and (inputs(66)));
    layer0_outputs(4869) <= not((inputs(143)) or (inputs(182)));
    layer0_outputs(4870) <= not((inputs(95)) or (inputs(224)));
    layer0_outputs(4871) <= not((inputs(213)) or (inputs(125)));
    layer0_outputs(4872) <= (inputs(65)) or (inputs(82));
    layer0_outputs(4873) <= not((inputs(33)) and (inputs(82)));
    layer0_outputs(4874) <= not(inputs(186)) or (inputs(6));
    layer0_outputs(4875) <= (inputs(39)) or (inputs(147));
    layer0_outputs(4876) <= (inputs(6)) or (inputs(111));
    layer0_outputs(4877) <= (inputs(185)) and not (inputs(16));
    layer0_outputs(4878) <= inputs(234);
    layer0_outputs(4879) <= (inputs(66)) xor (inputs(168));
    layer0_outputs(4880) <= not(inputs(30)) or (inputs(79));
    layer0_outputs(4881) <= inputs(37);
    layer0_outputs(4882) <= not(inputs(8));
    layer0_outputs(4883) <= not(inputs(153)) or (inputs(34));
    layer0_outputs(4884) <= '0';
    layer0_outputs(4885) <= (inputs(44)) and not (inputs(213));
    layer0_outputs(4886) <= (inputs(132)) and not (inputs(94));
    layer0_outputs(4887) <= (inputs(129)) xor (inputs(188));
    layer0_outputs(4888) <= not((inputs(23)) and (inputs(182)));
    layer0_outputs(4889) <= not((inputs(126)) or (inputs(184)));
    layer0_outputs(4890) <= not(inputs(120));
    layer0_outputs(4891) <= not(inputs(13));
    layer0_outputs(4892) <= (inputs(124)) or (inputs(101));
    layer0_outputs(4893) <= not((inputs(219)) or (inputs(230)));
    layer0_outputs(4894) <= (inputs(117)) and not (inputs(4));
    layer0_outputs(4895) <= not((inputs(244)) or (inputs(234)));
    layer0_outputs(4896) <= not(inputs(218));
    layer0_outputs(4897) <= '0';
    layer0_outputs(4898) <= (inputs(237)) or (inputs(109));
    layer0_outputs(4899) <= (inputs(139)) and not (inputs(69));
    layer0_outputs(4900) <= not((inputs(158)) xor (inputs(84)));
    layer0_outputs(4901) <= not((inputs(167)) or (inputs(183)));
    layer0_outputs(4902) <= inputs(71);
    layer0_outputs(4903) <= inputs(124);
    layer0_outputs(4904) <= not(inputs(235));
    layer0_outputs(4905) <= not(inputs(124)) or (inputs(238));
    layer0_outputs(4906) <= (inputs(12)) xor (inputs(128));
    layer0_outputs(4907) <= not(inputs(50));
    layer0_outputs(4908) <= not((inputs(153)) or (inputs(47)));
    layer0_outputs(4909) <= '1';
    layer0_outputs(4910) <= (inputs(134)) xor (inputs(224));
    layer0_outputs(4911) <= not(inputs(144));
    layer0_outputs(4912) <= inputs(182);
    layer0_outputs(4913) <= '1';
    layer0_outputs(4914) <= (inputs(205)) or (inputs(206));
    layer0_outputs(4915) <= (inputs(200)) and not (inputs(1));
    layer0_outputs(4916) <= inputs(168);
    layer0_outputs(4917) <= inputs(139);
    layer0_outputs(4918) <= not(inputs(21));
    layer0_outputs(4919) <= (inputs(225)) or (inputs(89));
    layer0_outputs(4920) <= (inputs(162)) or (inputs(160));
    layer0_outputs(4921) <= not(inputs(246));
    layer0_outputs(4922) <= (inputs(212)) and not (inputs(233));
    layer0_outputs(4923) <= inputs(74);
    layer0_outputs(4924) <= not(inputs(8));
    layer0_outputs(4925) <= '0';
    layer0_outputs(4926) <= not((inputs(38)) xor (inputs(68)));
    layer0_outputs(4927) <= (inputs(146)) or (inputs(93));
    layer0_outputs(4928) <= inputs(112);
    layer0_outputs(4929) <= not(inputs(5)) or (inputs(27));
    layer0_outputs(4930) <= inputs(218);
    layer0_outputs(4931) <= not((inputs(195)) or (inputs(192)));
    layer0_outputs(4932) <= (inputs(142)) xor (inputs(175));
    layer0_outputs(4933) <= (inputs(189)) and not (inputs(26));
    layer0_outputs(4934) <= inputs(23);
    layer0_outputs(4935) <= not(inputs(31)) or (inputs(217));
    layer0_outputs(4936) <= not((inputs(56)) xor (inputs(43)));
    layer0_outputs(4937) <= inputs(219);
    layer0_outputs(4938) <= not((inputs(6)) xor (inputs(172)));
    layer0_outputs(4939) <= not(inputs(173));
    layer0_outputs(4940) <= inputs(183);
    layer0_outputs(4941) <= inputs(144);
    layer0_outputs(4942) <= not((inputs(58)) and (inputs(95)));
    layer0_outputs(4943) <= not((inputs(27)) xor (inputs(104)));
    layer0_outputs(4944) <= (inputs(5)) and (inputs(204));
    layer0_outputs(4945) <= (inputs(145)) and not (inputs(53));
    layer0_outputs(4946) <= inputs(38);
    layer0_outputs(4947) <= (inputs(19)) and not (inputs(255));
    layer0_outputs(4948) <= inputs(67);
    layer0_outputs(4949) <= (inputs(74)) and not (inputs(179));
    layer0_outputs(4950) <= not((inputs(1)) and (inputs(215)));
    layer0_outputs(4951) <= (inputs(153)) and not (inputs(177));
    layer0_outputs(4952) <= not((inputs(53)) xor (inputs(20)));
    layer0_outputs(4953) <= not(inputs(245));
    layer0_outputs(4954) <= not(inputs(179)) or (inputs(253));
    layer0_outputs(4955) <= not(inputs(46)) or (inputs(9));
    layer0_outputs(4956) <= '0';
    layer0_outputs(4957) <= not((inputs(2)) xor (inputs(115)));
    layer0_outputs(4958) <= not((inputs(163)) or (inputs(239)));
    layer0_outputs(4959) <= inputs(155);
    layer0_outputs(4960) <= (inputs(125)) and not (inputs(238));
    layer0_outputs(4961) <= inputs(184);
    layer0_outputs(4962) <= inputs(25);
    layer0_outputs(4963) <= not((inputs(205)) or (inputs(57)));
    layer0_outputs(4964) <= (inputs(12)) and not (inputs(222));
    layer0_outputs(4965) <= (inputs(33)) xor (inputs(189));
    layer0_outputs(4966) <= not((inputs(69)) and (inputs(33)));
    layer0_outputs(4967) <= not((inputs(176)) xor (inputs(33)));
    layer0_outputs(4968) <= (inputs(112)) or (inputs(187));
    layer0_outputs(4969) <= inputs(102);
    layer0_outputs(4970) <= not(inputs(182));
    layer0_outputs(4971) <= inputs(246);
    layer0_outputs(4972) <= not((inputs(25)) xor (inputs(3)));
    layer0_outputs(4973) <= (inputs(220)) or (inputs(208));
    layer0_outputs(4974) <= not(inputs(206));
    layer0_outputs(4975) <= inputs(100);
    layer0_outputs(4976) <= not((inputs(255)) or (inputs(123)));
    layer0_outputs(4977) <= inputs(83);
    layer0_outputs(4978) <= not((inputs(139)) and (inputs(155)));
    layer0_outputs(4979) <= not(inputs(102)) or (inputs(117));
    layer0_outputs(4980) <= (inputs(33)) or (inputs(252));
    layer0_outputs(4981) <= inputs(176);
    layer0_outputs(4982) <= not(inputs(153));
    layer0_outputs(4983) <= (inputs(233)) and (inputs(15));
    layer0_outputs(4984) <= not((inputs(158)) xor (inputs(255)));
    layer0_outputs(4985) <= inputs(0);
    layer0_outputs(4986) <= not((inputs(112)) xor (inputs(232)));
    layer0_outputs(4987) <= not((inputs(212)) and (inputs(234)));
    layer0_outputs(4988) <= inputs(50);
    layer0_outputs(4989) <= inputs(141);
    layer0_outputs(4990) <= inputs(162);
    layer0_outputs(4991) <= not(inputs(78));
    layer0_outputs(4992) <= inputs(175);
    layer0_outputs(4993) <= inputs(132);
    layer0_outputs(4994) <= not((inputs(12)) xor (inputs(22)));
    layer0_outputs(4995) <= (inputs(114)) and not (inputs(207));
    layer0_outputs(4996) <= not(inputs(113));
    layer0_outputs(4997) <= (inputs(24)) and not (inputs(142));
    layer0_outputs(4998) <= not((inputs(198)) xor (inputs(61)));
    layer0_outputs(4999) <= not((inputs(80)) or (inputs(251)));
    layer0_outputs(5000) <= not((inputs(213)) or (inputs(243)));
    layer0_outputs(5001) <= not(inputs(86)) or (inputs(70));
    layer0_outputs(5002) <= (inputs(116)) and not (inputs(34));
    layer0_outputs(5003) <= not((inputs(89)) xor (inputs(228)));
    layer0_outputs(5004) <= inputs(86);
    layer0_outputs(5005) <= '1';
    layer0_outputs(5006) <= not(inputs(52));
    layer0_outputs(5007) <= (inputs(55)) and (inputs(40));
    layer0_outputs(5008) <= (inputs(173)) xor (inputs(19));
    layer0_outputs(5009) <= (inputs(234)) or (inputs(3));
    layer0_outputs(5010) <= (inputs(198)) and (inputs(95));
    layer0_outputs(5011) <= inputs(109);
    layer0_outputs(5012) <= not((inputs(125)) xor (inputs(125)));
    layer0_outputs(5013) <= inputs(165);
    layer0_outputs(5014) <= inputs(199);
    layer0_outputs(5015) <= inputs(105);
    layer0_outputs(5016) <= not(inputs(61));
    layer0_outputs(5017) <= not((inputs(220)) and (inputs(30)));
    layer0_outputs(5018) <= not((inputs(23)) xor (inputs(85)));
    layer0_outputs(5019) <= '0';
    layer0_outputs(5020) <= (inputs(116)) or (inputs(249));
    layer0_outputs(5021) <= '0';
    layer0_outputs(5022) <= inputs(54);
    layer0_outputs(5023) <= inputs(35);
    layer0_outputs(5024) <= not(inputs(75)) or (inputs(227));
    layer0_outputs(5025) <= not((inputs(77)) xor (inputs(17)));
    layer0_outputs(5026) <= not((inputs(8)) and (inputs(132)));
    layer0_outputs(5027) <= inputs(157);
    layer0_outputs(5028) <= not(inputs(7)) or (inputs(8));
    layer0_outputs(5029) <= not(inputs(148));
    layer0_outputs(5030) <= not(inputs(90)) or (inputs(221));
    layer0_outputs(5031) <= not(inputs(161));
    layer0_outputs(5032) <= (inputs(133)) or (inputs(14));
    layer0_outputs(5033) <= not((inputs(168)) or (inputs(111)));
    layer0_outputs(5034) <= not((inputs(165)) and (inputs(245)));
    layer0_outputs(5035) <= not(inputs(124));
    layer0_outputs(5036) <= inputs(23);
    layer0_outputs(5037) <= not((inputs(189)) or (inputs(249)));
    layer0_outputs(5038) <= not((inputs(72)) or (inputs(206)));
    layer0_outputs(5039) <= (inputs(100)) or (inputs(195));
    layer0_outputs(5040) <= not(inputs(59)) or (inputs(205));
    layer0_outputs(5041) <= inputs(184);
    layer0_outputs(5042) <= not((inputs(144)) xor (inputs(65)));
    layer0_outputs(5043) <= not(inputs(202));
    layer0_outputs(5044) <= inputs(23);
    layer0_outputs(5045) <= not(inputs(138));
    layer0_outputs(5046) <= (inputs(107)) and not (inputs(133));
    layer0_outputs(5047) <= not((inputs(41)) and (inputs(45)));
    layer0_outputs(5048) <= (inputs(13)) and not (inputs(245));
    layer0_outputs(5049) <= not(inputs(87)) or (inputs(37));
    layer0_outputs(5050) <= (inputs(106)) and not (inputs(47));
    layer0_outputs(5051) <= (inputs(26)) or (inputs(9));
    layer0_outputs(5052) <= not(inputs(18)) or (inputs(141));
    layer0_outputs(5053) <= not((inputs(115)) and (inputs(131)));
    layer0_outputs(5054) <= not((inputs(90)) or (inputs(146)));
    layer0_outputs(5055) <= not(inputs(219));
    layer0_outputs(5056) <= not(inputs(88)) or (inputs(80));
    layer0_outputs(5057) <= not(inputs(148));
    layer0_outputs(5058) <= (inputs(163)) xor (inputs(95));
    layer0_outputs(5059) <= (inputs(90)) and not (inputs(162));
    layer0_outputs(5060) <= (inputs(117)) and (inputs(255));
    layer0_outputs(5061) <= (inputs(36)) or (inputs(51));
    layer0_outputs(5062) <= (inputs(208)) or (inputs(205));
    layer0_outputs(5063) <= not(inputs(23));
    layer0_outputs(5064) <= (inputs(119)) and not (inputs(170));
    layer0_outputs(5065) <= inputs(77);
    layer0_outputs(5066) <= not(inputs(180)) or (inputs(89));
    layer0_outputs(5067) <= (inputs(1)) or (inputs(151));
    layer0_outputs(5068) <= inputs(35);
    layer0_outputs(5069) <= (inputs(202)) and not (inputs(97));
    layer0_outputs(5070) <= not(inputs(232));
    layer0_outputs(5071) <= (inputs(210)) and not (inputs(80));
    layer0_outputs(5072) <= (inputs(152)) xor (inputs(255));
    layer0_outputs(5073) <= not(inputs(151));
    layer0_outputs(5074) <= not((inputs(150)) or (inputs(137)));
    layer0_outputs(5075) <= (inputs(12)) xor (inputs(21));
    layer0_outputs(5076) <= not((inputs(175)) xor (inputs(246)));
    layer0_outputs(5077) <= inputs(215);
    layer0_outputs(5078) <= not(inputs(131));
    layer0_outputs(5079) <= (inputs(148)) and not (inputs(145));
    layer0_outputs(5080) <= (inputs(167)) xor (inputs(152));
    layer0_outputs(5081) <= inputs(124);
    layer0_outputs(5082) <= not((inputs(102)) and (inputs(232)));
    layer0_outputs(5083) <= not((inputs(33)) or (inputs(211)));
    layer0_outputs(5084) <= (inputs(186)) or (inputs(31));
    layer0_outputs(5085) <= (inputs(83)) and not (inputs(117));
    layer0_outputs(5086) <= not(inputs(58)) or (inputs(32));
    layer0_outputs(5087) <= not((inputs(94)) or (inputs(44)));
    layer0_outputs(5088) <= (inputs(173)) and not (inputs(255));
    layer0_outputs(5089) <= not(inputs(224)) or (inputs(15));
    layer0_outputs(5090) <= inputs(12);
    layer0_outputs(5091) <= not((inputs(66)) xor (inputs(226)));
    layer0_outputs(5092) <= (inputs(59)) and not (inputs(175));
    layer0_outputs(5093) <= (inputs(12)) or (inputs(185));
    layer0_outputs(5094) <= not((inputs(217)) xor (inputs(238)));
    layer0_outputs(5095) <= not(inputs(105));
    layer0_outputs(5096) <= (inputs(172)) xor (inputs(36));
    layer0_outputs(5097) <= '0';
    layer0_outputs(5098) <= (inputs(81)) and (inputs(35));
    layer0_outputs(5099) <= inputs(157);
    layer0_outputs(5100) <= (inputs(146)) and not (inputs(63));
    layer0_outputs(5101) <= not(inputs(19));
    layer0_outputs(5102) <= not(inputs(129));
    layer0_outputs(5103) <= (inputs(52)) or (inputs(221));
    layer0_outputs(5104) <= not(inputs(12)) or (inputs(193));
    layer0_outputs(5105) <= inputs(93);
    layer0_outputs(5106) <= (inputs(40)) and not (inputs(134));
    layer0_outputs(5107) <= not(inputs(45));
    layer0_outputs(5108) <= not(inputs(30)) or (inputs(246));
    layer0_outputs(5109) <= (inputs(70)) and (inputs(41));
    layer0_outputs(5110) <= not((inputs(232)) or (inputs(157)));
    layer0_outputs(5111) <= not((inputs(78)) or (inputs(98)));
    layer0_outputs(5112) <= not(inputs(198));
    layer0_outputs(5113) <= not((inputs(154)) or (inputs(221)));
    layer0_outputs(5114) <= (inputs(42)) or (inputs(108));
    layer0_outputs(5115) <= inputs(195);
    layer0_outputs(5116) <= not(inputs(239));
    layer0_outputs(5117) <= not((inputs(241)) or (inputs(171)));
    layer0_outputs(5118) <= (inputs(65)) and (inputs(4));
    layer0_outputs(5119) <= inputs(239);
    layer0_outputs(5120) <= inputs(24);
    layer0_outputs(5121) <= (inputs(65)) xor (inputs(74));
    layer0_outputs(5122) <= (inputs(161)) and not (inputs(124));
    layer0_outputs(5123) <= not(inputs(231));
    layer0_outputs(5124) <= inputs(107);
    layer0_outputs(5125) <= not(inputs(166)) or (inputs(91));
    layer0_outputs(5126) <= not(inputs(118)) or (inputs(24));
    layer0_outputs(5127) <= (inputs(33)) and (inputs(105));
    layer0_outputs(5128) <= not(inputs(204)) or (inputs(168));
    layer0_outputs(5129) <= not(inputs(7));
    layer0_outputs(5130) <= not((inputs(84)) xor (inputs(132)));
    layer0_outputs(5131) <= not(inputs(105));
    layer0_outputs(5132) <= not((inputs(85)) or (inputs(144)));
    layer0_outputs(5133) <= (inputs(229)) xor (inputs(197));
    layer0_outputs(5134) <= not(inputs(63));
    layer0_outputs(5135) <= (inputs(86)) and not (inputs(2));
    layer0_outputs(5136) <= (inputs(142)) or (inputs(147));
    layer0_outputs(5137) <= (inputs(198)) and not (inputs(87));
    layer0_outputs(5138) <= not((inputs(134)) or (inputs(81)));
    layer0_outputs(5139) <= not(inputs(229));
    layer0_outputs(5140) <= not(inputs(127));
    layer0_outputs(5141) <= not((inputs(176)) xor (inputs(93)));
    layer0_outputs(5142) <= not(inputs(133)) or (inputs(224));
    layer0_outputs(5143) <= not((inputs(47)) or (inputs(169)));
    layer0_outputs(5144) <= not(inputs(45)) or (inputs(48));
    layer0_outputs(5145) <= not(inputs(48)) or (inputs(24));
    layer0_outputs(5146) <= (inputs(8)) or (inputs(204));
    layer0_outputs(5147) <= (inputs(235)) or (inputs(171));
    layer0_outputs(5148) <= inputs(243);
    layer0_outputs(5149) <= (inputs(104)) xor (inputs(18));
    layer0_outputs(5150) <= '1';
    layer0_outputs(5151) <= (inputs(54)) and not (inputs(192));
    layer0_outputs(5152) <= (inputs(135)) and not (inputs(154));
    layer0_outputs(5153) <= not(inputs(255)) or (inputs(31));
    layer0_outputs(5154) <= not(inputs(82));
    layer0_outputs(5155) <= (inputs(182)) and not (inputs(91));
    layer0_outputs(5156) <= inputs(243);
    layer0_outputs(5157) <= '0';
    layer0_outputs(5158) <= not(inputs(171));
    layer0_outputs(5159) <= inputs(75);
    layer0_outputs(5160) <= (inputs(247)) and not (inputs(68));
    layer0_outputs(5161) <= not(inputs(107));
    layer0_outputs(5162) <= not((inputs(210)) or (inputs(223)));
    layer0_outputs(5163) <= not(inputs(39));
    layer0_outputs(5164) <= inputs(202);
    layer0_outputs(5165) <= inputs(83);
    layer0_outputs(5166) <= (inputs(246)) and not (inputs(91));
    layer0_outputs(5167) <= (inputs(223)) and not (inputs(221));
    layer0_outputs(5168) <= (inputs(85)) and not (inputs(243));
    layer0_outputs(5169) <= inputs(123);
    layer0_outputs(5170) <= (inputs(200)) and not (inputs(88));
    layer0_outputs(5171) <= inputs(100);
    layer0_outputs(5172) <= '0';
    layer0_outputs(5173) <= not(inputs(227)) or (inputs(133));
    layer0_outputs(5174) <= (inputs(68)) or (inputs(75));
    layer0_outputs(5175) <= inputs(86);
    layer0_outputs(5176) <= not(inputs(170)) or (inputs(65));
    layer0_outputs(5177) <= not(inputs(45)) or (inputs(169));
    layer0_outputs(5178) <= not(inputs(227));
    layer0_outputs(5179) <= not((inputs(95)) or (inputs(11)));
    layer0_outputs(5180) <= not((inputs(33)) or (inputs(35)));
    layer0_outputs(5181) <= not(inputs(70)) or (inputs(119));
    layer0_outputs(5182) <= not(inputs(24));
    layer0_outputs(5183) <= not(inputs(180));
    layer0_outputs(5184) <= not(inputs(102));
    layer0_outputs(5185) <= inputs(152);
    layer0_outputs(5186) <= not((inputs(111)) xor (inputs(31)));
    layer0_outputs(5187) <= (inputs(254)) or (inputs(222));
    layer0_outputs(5188) <= not((inputs(121)) or (inputs(166)));
    layer0_outputs(5189) <= not(inputs(100));
    layer0_outputs(5190) <= not((inputs(17)) or (inputs(88)));
    layer0_outputs(5191) <= '0';
    layer0_outputs(5192) <= (inputs(98)) or (inputs(168));
    layer0_outputs(5193) <= (inputs(81)) xor (inputs(19));
    layer0_outputs(5194) <= (inputs(208)) xor (inputs(29));
    layer0_outputs(5195) <= inputs(134);
    layer0_outputs(5196) <= not(inputs(116));
    layer0_outputs(5197) <= (inputs(181)) or (inputs(102));
    layer0_outputs(5198) <= not((inputs(194)) or (inputs(125)));
    layer0_outputs(5199) <= not((inputs(21)) or (inputs(124)));
    layer0_outputs(5200) <= (inputs(253)) or (inputs(205));
    layer0_outputs(5201) <= not(inputs(108)) or (inputs(175));
    layer0_outputs(5202) <= not(inputs(6)) or (inputs(13));
    layer0_outputs(5203) <= not((inputs(223)) or (inputs(159)));
    layer0_outputs(5204) <= not(inputs(36));
    layer0_outputs(5205) <= inputs(78);
    layer0_outputs(5206) <= not(inputs(153));
    layer0_outputs(5207) <= (inputs(53)) or (inputs(55));
    layer0_outputs(5208) <= (inputs(63)) and not (inputs(45));
    layer0_outputs(5209) <= (inputs(66)) or (inputs(48));
    layer0_outputs(5210) <= (inputs(116)) xor (inputs(98));
    layer0_outputs(5211) <= not(inputs(200));
    layer0_outputs(5212) <= not((inputs(81)) or (inputs(103)));
    layer0_outputs(5213) <= not(inputs(169)) or (inputs(72));
    layer0_outputs(5214) <= not(inputs(186)) or (inputs(8));
    layer0_outputs(5215) <= (inputs(159)) and not (inputs(155));
    layer0_outputs(5216) <= inputs(213);
    layer0_outputs(5217) <= not(inputs(90)) or (inputs(168));
    layer0_outputs(5218) <= inputs(55);
    layer0_outputs(5219) <= not(inputs(13));
    layer0_outputs(5220) <= not(inputs(216));
    layer0_outputs(5221) <= not(inputs(50)) or (inputs(199));
    layer0_outputs(5222) <= not(inputs(224));
    layer0_outputs(5223) <= not(inputs(144));
    layer0_outputs(5224) <= (inputs(80)) or (inputs(124));
    layer0_outputs(5225) <= (inputs(92)) and not (inputs(221));
    layer0_outputs(5226) <= not(inputs(190));
    layer0_outputs(5227) <= not(inputs(93));
    layer0_outputs(5228) <= '1';
    layer0_outputs(5229) <= inputs(227);
    layer0_outputs(5230) <= not(inputs(214));
    layer0_outputs(5231) <= '1';
    layer0_outputs(5232) <= (inputs(68)) xor (inputs(51));
    layer0_outputs(5233) <= not((inputs(156)) or (inputs(116)));
    layer0_outputs(5234) <= not(inputs(243)) or (inputs(57));
    layer0_outputs(5235) <= inputs(162);
    layer0_outputs(5236) <= (inputs(24)) and not (inputs(14));
    layer0_outputs(5237) <= '1';
    layer0_outputs(5238) <= not(inputs(38)) or (inputs(210));
    layer0_outputs(5239) <= inputs(24);
    layer0_outputs(5240) <= (inputs(95)) xor (inputs(225));
    layer0_outputs(5241) <= (inputs(183)) and not (inputs(155));
    layer0_outputs(5242) <= not((inputs(145)) xor (inputs(118)));
    layer0_outputs(5243) <= '1';
    layer0_outputs(5244) <= (inputs(190)) xor (inputs(13));
    layer0_outputs(5245) <= not((inputs(102)) xor (inputs(182)));
    layer0_outputs(5246) <= (inputs(81)) or (inputs(82));
    layer0_outputs(5247) <= not((inputs(81)) and (inputs(207)));
    layer0_outputs(5248) <= not((inputs(37)) xor (inputs(64)));
    layer0_outputs(5249) <= not(inputs(206));
    layer0_outputs(5250) <= not((inputs(37)) xor (inputs(146)));
    layer0_outputs(5251) <= not(inputs(83)) or (inputs(174));
    layer0_outputs(5252) <= not(inputs(156));
    layer0_outputs(5253) <= not((inputs(86)) xor (inputs(126)));
    layer0_outputs(5254) <= inputs(56);
    layer0_outputs(5255) <= not(inputs(136)) or (inputs(202));
    layer0_outputs(5256) <= '1';
    layer0_outputs(5257) <= inputs(224);
    layer0_outputs(5258) <= not((inputs(84)) or (inputs(148)));
    layer0_outputs(5259) <= not((inputs(115)) or (inputs(131)));
    layer0_outputs(5260) <= (inputs(151)) and not (inputs(140));
    layer0_outputs(5261) <= not(inputs(80));
    layer0_outputs(5262) <= not(inputs(32)) or (inputs(32));
    layer0_outputs(5263) <= (inputs(60)) or (inputs(79));
    layer0_outputs(5264) <= (inputs(68)) and (inputs(24));
    layer0_outputs(5265) <= (inputs(232)) or (inputs(67));
    layer0_outputs(5266) <= (inputs(80)) xor (inputs(110));
    layer0_outputs(5267) <= not(inputs(174)) or (inputs(186));
    layer0_outputs(5268) <= not((inputs(106)) and (inputs(137)));
    layer0_outputs(5269) <= (inputs(238)) or (inputs(238));
    layer0_outputs(5270) <= (inputs(226)) and not (inputs(217));
    layer0_outputs(5271) <= not(inputs(201)) or (inputs(207));
    layer0_outputs(5272) <= inputs(225);
    layer0_outputs(5273) <= not((inputs(238)) or (inputs(106)));
    layer0_outputs(5274) <= (inputs(136)) or (inputs(122));
    layer0_outputs(5275) <= not(inputs(103));
    layer0_outputs(5276) <= (inputs(10)) and not (inputs(31));
    layer0_outputs(5277) <= not(inputs(221));
    layer0_outputs(5278) <= not(inputs(237));
    layer0_outputs(5279) <= inputs(121);
    layer0_outputs(5280) <= (inputs(129)) xor (inputs(127));
    layer0_outputs(5281) <= (inputs(21)) and not (inputs(205));
    layer0_outputs(5282) <= (inputs(167)) and not (inputs(128));
    layer0_outputs(5283) <= not(inputs(177));
    layer0_outputs(5284) <= not(inputs(32)) or (inputs(38));
    layer0_outputs(5285) <= inputs(51);
    layer0_outputs(5286) <= not((inputs(235)) xor (inputs(186)));
    layer0_outputs(5287) <= not(inputs(247));
    layer0_outputs(5288) <= (inputs(95)) or (inputs(102));
    layer0_outputs(5289) <= not((inputs(124)) xor (inputs(7)));
    layer0_outputs(5290) <= not(inputs(58)) or (inputs(13));
    layer0_outputs(5291) <= inputs(83);
    layer0_outputs(5292) <= not(inputs(110));
    layer0_outputs(5293) <= (inputs(168)) or (inputs(126));
    layer0_outputs(5294) <= not(inputs(56));
    layer0_outputs(5295) <= not(inputs(216)) or (inputs(145));
    layer0_outputs(5296) <= not((inputs(38)) and (inputs(198)));
    layer0_outputs(5297) <= '0';
    layer0_outputs(5298) <= inputs(60);
    layer0_outputs(5299) <= not(inputs(14)) or (inputs(127));
    layer0_outputs(5300) <= inputs(50);
    layer0_outputs(5301) <= not(inputs(123));
    layer0_outputs(5302) <= not(inputs(211)) or (inputs(205));
    layer0_outputs(5303) <= not((inputs(232)) xor (inputs(16)));
    layer0_outputs(5304) <= not((inputs(168)) or (inputs(97)));
    layer0_outputs(5305) <= not(inputs(156)) or (inputs(9));
    layer0_outputs(5306) <= (inputs(124)) and not (inputs(112));
    layer0_outputs(5307) <= (inputs(148)) xor (inputs(2));
    layer0_outputs(5308) <= (inputs(157)) and not (inputs(102));
    layer0_outputs(5309) <= not((inputs(32)) xor (inputs(76)));
    layer0_outputs(5310) <= not(inputs(83)) or (inputs(161));
    layer0_outputs(5311) <= not(inputs(122)) or (inputs(223));
    layer0_outputs(5312) <= (inputs(87)) and not (inputs(48));
    layer0_outputs(5313) <= not(inputs(41)) or (inputs(60));
    layer0_outputs(5314) <= inputs(39);
    layer0_outputs(5315) <= not((inputs(161)) or (inputs(243)));
    layer0_outputs(5316) <= (inputs(208)) and not (inputs(176));
    layer0_outputs(5317) <= (inputs(5)) and not (inputs(153));
    layer0_outputs(5318) <= inputs(40);
    layer0_outputs(5319) <= not(inputs(151));
    layer0_outputs(5320) <= (inputs(69)) and not (inputs(172));
    layer0_outputs(5321) <= (inputs(255)) and not (inputs(148));
    layer0_outputs(5322) <= not((inputs(155)) xor (inputs(190)));
    layer0_outputs(5323) <= not((inputs(223)) xor (inputs(237)));
    layer0_outputs(5324) <= inputs(166);
    layer0_outputs(5325) <= (inputs(97)) or (inputs(185));
    layer0_outputs(5326) <= not(inputs(38)) or (inputs(13));
    layer0_outputs(5327) <= inputs(123);
    layer0_outputs(5328) <= not((inputs(236)) and (inputs(241)));
    layer0_outputs(5329) <= not(inputs(176)) or (inputs(146));
    layer0_outputs(5330) <= inputs(167);
    layer0_outputs(5331) <= not(inputs(24));
    layer0_outputs(5332) <= (inputs(185)) xor (inputs(136));
    layer0_outputs(5333) <= not(inputs(183));
    layer0_outputs(5334) <= (inputs(19)) and (inputs(99));
    layer0_outputs(5335) <= not((inputs(92)) xor (inputs(33)));
    layer0_outputs(5336) <= not(inputs(193));
    layer0_outputs(5337) <= (inputs(127)) and not (inputs(228));
    layer0_outputs(5338) <= inputs(84);
    layer0_outputs(5339) <= not(inputs(9));
    layer0_outputs(5340) <= not((inputs(75)) or (inputs(28)));
    layer0_outputs(5341) <= not((inputs(224)) or (inputs(4)));
    layer0_outputs(5342) <= not((inputs(160)) xor (inputs(100)));
    layer0_outputs(5343) <= not(inputs(6)) or (inputs(96));
    layer0_outputs(5344) <= (inputs(224)) and not (inputs(210));
    layer0_outputs(5345) <= not((inputs(235)) or (inputs(97)));
    layer0_outputs(5346) <= not((inputs(60)) or (inputs(46)));
    layer0_outputs(5347) <= (inputs(161)) or (inputs(217));
    layer0_outputs(5348) <= (inputs(23)) and not (inputs(59));
    layer0_outputs(5349) <= inputs(129);
    layer0_outputs(5350) <= not((inputs(94)) xor (inputs(197)));
    layer0_outputs(5351) <= (inputs(35)) xor (inputs(131));
    layer0_outputs(5352) <= (inputs(18)) xor (inputs(70));
    layer0_outputs(5353) <= (inputs(60)) and not (inputs(238));
    layer0_outputs(5354) <= (inputs(245)) xor (inputs(161));
    layer0_outputs(5355) <= not(inputs(170)) or (inputs(69));
    layer0_outputs(5356) <= not(inputs(194));
    layer0_outputs(5357) <= (inputs(19)) or (inputs(8));
    layer0_outputs(5358) <= not((inputs(28)) or (inputs(177)));
    layer0_outputs(5359) <= (inputs(243)) and not (inputs(142));
    layer0_outputs(5360) <= not(inputs(115)) or (inputs(109));
    layer0_outputs(5361) <= not((inputs(225)) or (inputs(211)));
    layer0_outputs(5362) <= not((inputs(151)) or (inputs(207)));
    layer0_outputs(5363) <= (inputs(1)) or (inputs(197));
    layer0_outputs(5364) <= not((inputs(173)) or (inputs(53)));
    layer0_outputs(5365) <= (inputs(231)) xor (inputs(255));
    layer0_outputs(5366) <= not(inputs(125));
    layer0_outputs(5367) <= (inputs(67)) and (inputs(153));
    layer0_outputs(5368) <= not(inputs(160));
    layer0_outputs(5369) <= (inputs(144)) xor (inputs(84));
    layer0_outputs(5370) <= inputs(234);
    layer0_outputs(5371) <= (inputs(162)) and not (inputs(251));
    layer0_outputs(5372) <= '1';
    layer0_outputs(5373) <= (inputs(116)) xor (inputs(128));
    layer0_outputs(5374) <= not(inputs(245));
    layer0_outputs(5375) <= (inputs(174)) and not (inputs(117));
    layer0_outputs(5376) <= inputs(212);
    layer0_outputs(5377) <= (inputs(217)) xor (inputs(210));
    layer0_outputs(5378) <= (inputs(69)) or (inputs(62));
    layer0_outputs(5379) <= not(inputs(214)) or (inputs(13));
    layer0_outputs(5380) <= not(inputs(223)) or (inputs(195));
    layer0_outputs(5381) <= inputs(41);
    layer0_outputs(5382) <= not(inputs(69)) or (inputs(101));
    layer0_outputs(5383) <= not((inputs(219)) and (inputs(114)));
    layer0_outputs(5384) <= inputs(76);
    layer0_outputs(5385) <= not(inputs(93));
    layer0_outputs(5386) <= not(inputs(166));
    layer0_outputs(5387) <= (inputs(200)) or (inputs(99));
    layer0_outputs(5388) <= '0';
    layer0_outputs(5389) <= not((inputs(63)) xor (inputs(90)));
    layer0_outputs(5390) <= (inputs(226)) and not (inputs(45));
    layer0_outputs(5391) <= not((inputs(90)) or (inputs(136)));
    layer0_outputs(5392) <= (inputs(204)) or (inputs(66));
    layer0_outputs(5393) <= not((inputs(188)) or (inputs(228)));
    layer0_outputs(5394) <= not((inputs(96)) and (inputs(74)));
    layer0_outputs(5395) <= not(inputs(253));
    layer0_outputs(5396) <= not(inputs(246)) or (inputs(119));
    layer0_outputs(5397) <= (inputs(65)) and not (inputs(108));
    layer0_outputs(5398) <= (inputs(66)) and not (inputs(79));
    layer0_outputs(5399) <= (inputs(179)) and not (inputs(160));
    layer0_outputs(5400) <= (inputs(95)) xor (inputs(19));
    layer0_outputs(5401) <= not((inputs(50)) or (inputs(86)));
    layer0_outputs(5402) <= (inputs(77)) and not (inputs(254));
    layer0_outputs(5403) <= not(inputs(225));
    layer0_outputs(5404) <= not((inputs(80)) or (inputs(196)));
    layer0_outputs(5405) <= not(inputs(211)) or (inputs(8));
    layer0_outputs(5406) <= not(inputs(251)) or (inputs(246));
    layer0_outputs(5407) <= not((inputs(210)) and (inputs(199)));
    layer0_outputs(5408) <= (inputs(97)) and (inputs(97));
    layer0_outputs(5409) <= not((inputs(189)) or (inputs(7)));
    layer0_outputs(5410) <= (inputs(112)) xor (inputs(99));
    layer0_outputs(5411) <= '1';
    layer0_outputs(5412) <= (inputs(9)) and not (inputs(191));
    layer0_outputs(5413) <= not(inputs(234));
    layer0_outputs(5414) <= (inputs(144)) and not (inputs(223));
    layer0_outputs(5415) <= not((inputs(214)) and (inputs(148)));
    layer0_outputs(5416) <= not(inputs(17)) or (inputs(222));
    layer0_outputs(5417) <= not(inputs(184));
    layer0_outputs(5418) <= inputs(151);
    layer0_outputs(5419) <= not(inputs(196)) or (inputs(113));
    layer0_outputs(5420) <= (inputs(105)) and not (inputs(161));
    layer0_outputs(5421) <= (inputs(48)) xor (inputs(17));
    layer0_outputs(5422) <= not(inputs(13));
    layer0_outputs(5423) <= not((inputs(72)) xor (inputs(12)));
    layer0_outputs(5424) <= not(inputs(188)) or (inputs(244));
    layer0_outputs(5425) <= inputs(190);
    layer0_outputs(5426) <= not((inputs(118)) xor (inputs(150)));
    layer0_outputs(5427) <= not((inputs(105)) and (inputs(179)));
    layer0_outputs(5428) <= (inputs(202)) and not (inputs(198));
    layer0_outputs(5429) <= not((inputs(134)) or (inputs(134)));
    layer0_outputs(5430) <= not(inputs(195)) or (inputs(57));
    layer0_outputs(5431) <= (inputs(46)) and not (inputs(191));
    layer0_outputs(5432) <= '0';
    layer0_outputs(5433) <= '1';
    layer0_outputs(5434) <= not(inputs(75));
    layer0_outputs(5435) <= not((inputs(164)) or (inputs(163)));
    layer0_outputs(5436) <= inputs(69);
    layer0_outputs(5437) <= (inputs(76)) and not (inputs(121));
    layer0_outputs(5438) <= inputs(103);
    layer0_outputs(5439) <= inputs(188);
    layer0_outputs(5440) <= (inputs(158)) and (inputs(212));
    layer0_outputs(5441) <= (inputs(192)) or (inputs(6));
    layer0_outputs(5442) <= not((inputs(163)) and (inputs(100)));
    layer0_outputs(5443) <= not((inputs(227)) xor (inputs(248)));
    layer0_outputs(5444) <= inputs(136);
    layer0_outputs(5445) <= (inputs(246)) and (inputs(6));
    layer0_outputs(5446) <= not((inputs(149)) and (inputs(141)));
    layer0_outputs(5447) <= not(inputs(42)) or (inputs(143));
    layer0_outputs(5448) <= inputs(73);
    layer0_outputs(5449) <= (inputs(205)) and (inputs(154));
    layer0_outputs(5450) <= inputs(56);
    layer0_outputs(5451) <= (inputs(72)) and not (inputs(58));
    layer0_outputs(5452) <= '1';
    layer0_outputs(5453) <= not((inputs(184)) xor (inputs(246)));
    layer0_outputs(5454) <= '0';
    layer0_outputs(5455) <= (inputs(198)) and not (inputs(236));
    layer0_outputs(5456) <= not(inputs(244));
    layer0_outputs(5457) <= not(inputs(55)) or (inputs(112));
    layer0_outputs(5458) <= (inputs(76)) xor (inputs(73));
    layer0_outputs(5459) <= not(inputs(148)) or (inputs(247));
    layer0_outputs(5460) <= not((inputs(107)) xor (inputs(0)));
    layer0_outputs(5461) <= (inputs(116)) xor (inputs(145));
    layer0_outputs(5462) <= not((inputs(149)) or (inputs(188)));
    layer0_outputs(5463) <= not(inputs(247)) or (inputs(223));
    layer0_outputs(5464) <= inputs(17);
    layer0_outputs(5465) <= inputs(162);
    layer0_outputs(5466) <= not((inputs(106)) xor (inputs(142)));
    layer0_outputs(5467) <= (inputs(157)) and not (inputs(239));
    layer0_outputs(5468) <= '0';
    layer0_outputs(5469) <= not(inputs(125));
    layer0_outputs(5470) <= '1';
    layer0_outputs(5471) <= (inputs(149)) xor (inputs(194));
    layer0_outputs(5472) <= (inputs(164)) xor (inputs(250));
    layer0_outputs(5473) <= not(inputs(222));
    layer0_outputs(5474) <= (inputs(199)) and not (inputs(16));
    layer0_outputs(5475) <= (inputs(56)) xor (inputs(13));
    layer0_outputs(5476) <= '0';
    layer0_outputs(5477) <= not(inputs(97));
    layer0_outputs(5478) <= (inputs(211)) and not (inputs(93));
    layer0_outputs(5479) <= (inputs(48)) and (inputs(94));
    layer0_outputs(5480) <= not(inputs(73));
    layer0_outputs(5481) <= (inputs(49)) and (inputs(111));
    layer0_outputs(5482) <= not((inputs(213)) or (inputs(14)));
    layer0_outputs(5483) <= not(inputs(61));
    layer0_outputs(5484) <= inputs(143);
    layer0_outputs(5485) <= '0';
    layer0_outputs(5486) <= not(inputs(152)) or (inputs(111));
    layer0_outputs(5487) <= '0';
    layer0_outputs(5488) <= not(inputs(147));
    layer0_outputs(5489) <= not(inputs(225));
    layer0_outputs(5490) <= not(inputs(134));
    layer0_outputs(5491) <= not(inputs(106)) or (inputs(83));
    layer0_outputs(5492) <= (inputs(156)) and not (inputs(211));
    layer0_outputs(5493) <= not(inputs(5)) or (inputs(11));
    layer0_outputs(5494) <= (inputs(246)) or (inputs(159));
    layer0_outputs(5495) <= not((inputs(184)) and (inputs(186)));
    layer0_outputs(5496) <= inputs(134);
    layer0_outputs(5497) <= not((inputs(14)) or (inputs(119)));
    layer0_outputs(5498) <= inputs(214);
    layer0_outputs(5499) <= inputs(145);
    layer0_outputs(5500) <= not(inputs(89)) or (inputs(238));
    layer0_outputs(5501) <= not((inputs(134)) or (inputs(143)));
    layer0_outputs(5502) <= (inputs(175)) xor (inputs(35));
    layer0_outputs(5503) <= not(inputs(182)) or (inputs(215));
    layer0_outputs(5504) <= (inputs(107)) xor (inputs(35));
    layer0_outputs(5505) <= (inputs(253)) and not (inputs(237));
    layer0_outputs(5506) <= '1';
    layer0_outputs(5507) <= inputs(119);
    layer0_outputs(5508) <= not(inputs(233));
    layer0_outputs(5509) <= (inputs(165)) and not (inputs(144));
    layer0_outputs(5510) <= not((inputs(24)) and (inputs(27)));
    layer0_outputs(5511) <= (inputs(186)) or (inputs(117));
    layer0_outputs(5512) <= not(inputs(43)) or (inputs(100));
    layer0_outputs(5513) <= (inputs(14)) and not (inputs(42));
    layer0_outputs(5514) <= inputs(213);
    layer0_outputs(5515) <= not((inputs(139)) or (inputs(147)));
    layer0_outputs(5516) <= (inputs(134)) or (inputs(204));
    layer0_outputs(5517) <= not(inputs(46)) or (inputs(42));
    layer0_outputs(5518) <= inputs(118);
    layer0_outputs(5519) <= (inputs(175)) or (inputs(186));
    layer0_outputs(5520) <= not(inputs(213)) or (inputs(201));
    layer0_outputs(5521) <= inputs(162);
    layer0_outputs(5522) <= not(inputs(243)) or (inputs(161));
    layer0_outputs(5523) <= inputs(85);
    layer0_outputs(5524) <= not(inputs(185));
    layer0_outputs(5525) <= '0';
    layer0_outputs(5526) <= (inputs(226)) xor (inputs(155));
    layer0_outputs(5527) <= (inputs(30)) and (inputs(34));
    layer0_outputs(5528) <= (inputs(92)) and (inputs(68));
    layer0_outputs(5529) <= (inputs(129)) or (inputs(189));
    layer0_outputs(5530) <= (inputs(89)) and not (inputs(191));
    layer0_outputs(5531) <= (inputs(172)) or (inputs(112));
    layer0_outputs(5532) <= (inputs(48)) and not (inputs(39));
    layer0_outputs(5533) <= not((inputs(231)) xor (inputs(226)));
    layer0_outputs(5534) <= not(inputs(23)) or (inputs(162));
    layer0_outputs(5535) <= (inputs(11)) and not (inputs(157));
    layer0_outputs(5536) <= not(inputs(140)) or (inputs(218));
    layer0_outputs(5537) <= inputs(85);
    layer0_outputs(5538) <= not((inputs(79)) and (inputs(192)));
    layer0_outputs(5539) <= inputs(186);
    layer0_outputs(5540) <= (inputs(154)) and not (inputs(15));
    layer0_outputs(5541) <= inputs(29);
    layer0_outputs(5542) <= not((inputs(95)) xor (inputs(60)));
    layer0_outputs(5543) <= not(inputs(199)) or (inputs(119));
    layer0_outputs(5544) <= inputs(214);
    layer0_outputs(5545) <= '1';
    layer0_outputs(5546) <= (inputs(230)) and (inputs(104));
    layer0_outputs(5547) <= (inputs(33)) or (inputs(51));
    layer0_outputs(5548) <= inputs(77);
    layer0_outputs(5549) <= not(inputs(171));
    layer0_outputs(5550) <= not((inputs(2)) or (inputs(21)));
    layer0_outputs(5551) <= inputs(77);
    layer0_outputs(5552) <= '0';
    layer0_outputs(5553) <= not((inputs(246)) or (inputs(226)));
    layer0_outputs(5554) <= not(inputs(101));
    layer0_outputs(5555) <= not(inputs(67));
    layer0_outputs(5556) <= not(inputs(129));
    layer0_outputs(5557) <= (inputs(46)) xor (inputs(32));
    layer0_outputs(5558) <= not(inputs(80));
    layer0_outputs(5559) <= (inputs(45)) xor (inputs(241));
    layer0_outputs(5560) <= not((inputs(95)) or (inputs(185)));
    layer0_outputs(5561) <= (inputs(229)) and not (inputs(94));
    layer0_outputs(5562) <= (inputs(210)) or (inputs(238));
    layer0_outputs(5563) <= not((inputs(202)) or (inputs(189)));
    layer0_outputs(5564) <= inputs(228);
    layer0_outputs(5565) <= not(inputs(33)) or (inputs(31));
    layer0_outputs(5566) <= inputs(230);
    layer0_outputs(5567) <= (inputs(120)) and not (inputs(157));
    layer0_outputs(5568) <= not(inputs(255)) or (inputs(227));
    layer0_outputs(5569) <= not(inputs(49));
    layer0_outputs(5570) <= not((inputs(149)) or (inputs(137)));
    layer0_outputs(5571) <= (inputs(103)) or (inputs(68));
    layer0_outputs(5572) <= inputs(186);
    layer0_outputs(5573) <= (inputs(31)) or (inputs(10));
    layer0_outputs(5574) <= (inputs(142)) xor (inputs(118));
    layer0_outputs(5575) <= (inputs(219)) or (inputs(212));
    layer0_outputs(5576) <= not(inputs(240)) or (inputs(28));
    layer0_outputs(5577) <= (inputs(139)) or (inputs(187));
    layer0_outputs(5578) <= inputs(136);
    layer0_outputs(5579) <= inputs(96);
    layer0_outputs(5580) <= inputs(7);
    layer0_outputs(5581) <= (inputs(130)) and not (inputs(213));
    layer0_outputs(5582) <= inputs(61);
    layer0_outputs(5583) <= not(inputs(28)) or (inputs(255));
    layer0_outputs(5584) <= not((inputs(84)) and (inputs(83)));
    layer0_outputs(5585) <= (inputs(250)) or (inputs(14));
    layer0_outputs(5586) <= (inputs(65)) and not (inputs(244));
    layer0_outputs(5587) <= not((inputs(20)) xor (inputs(188)));
    layer0_outputs(5588) <= not(inputs(40));
    layer0_outputs(5589) <= inputs(27);
    layer0_outputs(5590) <= (inputs(28)) and (inputs(85));
    layer0_outputs(5591) <= not(inputs(78));
    layer0_outputs(5592) <= not((inputs(216)) xor (inputs(234)));
    layer0_outputs(5593) <= (inputs(207)) and not (inputs(178));
    layer0_outputs(5594) <= inputs(156);
    layer0_outputs(5595) <= inputs(57);
    layer0_outputs(5596) <= (inputs(25)) xor (inputs(231));
    layer0_outputs(5597) <= not(inputs(121)) or (inputs(144));
    layer0_outputs(5598) <= (inputs(61)) and not (inputs(170));
    layer0_outputs(5599) <= (inputs(232)) or (inputs(113));
    layer0_outputs(5600) <= (inputs(194)) xor (inputs(220));
    layer0_outputs(5601) <= not(inputs(213));
    layer0_outputs(5602) <= (inputs(160)) or (inputs(245));
    layer0_outputs(5603) <= not((inputs(132)) and (inputs(157)));
    layer0_outputs(5604) <= not((inputs(180)) xor (inputs(160)));
    layer0_outputs(5605) <= (inputs(134)) or (inputs(166));
    layer0_outputs(5606) <= (inputs(114)) and (inputs(25));
    layer0_outputs(5607) <= not((inputs(213)) and (inputs(246)));
    layer0_outputs(5608) <= not(inputs(249));
    layer0_outputs(5609) <= not((inputs(150)) or (inputs(22)));
    layer0_outputs(5610) <= inputs(14);
    layer0_outputs(5611) <= not((inputs(11)) xor (inputs(207)));
    layer0_outputs(5612) <= inputs(10);
    layer0_outputs(5613) <= inputs(97);
    layer0_outputs(5614) <= not((inputs(160)) or (inputs(32)));
    layer0_outputs(5615) <= not(inputs(190));
    layer0_outputs(5616) <= not(inputs(34)) or (inputs(191));
    layer0_outputs(5617) <= not(inputs(194));
    layer0_outputs(5618) <= (inputs(231)) and (inputs(253));
    layer0_outputs(5619) <= (inputs(19)) and not (inputs(187));
    layer0_outputs(5620) <= inputs(162);
    layer0_outputs(5621) <= not(inputs(242));
    layer0_outputs(5622) <= not((inputs(44)) or (inputs(63)));
    layer0_outputs(5623) <= not((inputs(255)) or (inputs(240)));
    layer0_outputs(5624) <= not((inputs(83)) or (inputs(221)));
    layer0_outputs(5625) <= not(inputs(40));
    layer0_outputs(5626) <= not((inputs(130)) xor (inputs(206)));
    layer0_outputs(5627) <= inputs(235);
    layer0_outputs(5628) <= not(inputs(24));
    layer0_outputs(5629) <= (inputs(250)) and (inputs(182));
    layer0_outputs(5630) <= not(inputs(27)) or (inputs(103));
    layer0_outputs(5631) <= not((inputs(230)) or (inputs(65)));
    layer0_outputs(5632) <= inputs(50);
    layer0_outputs(5633) <= '1';
    layer0_outputs(5634) <= not((inputs(197)) or (inputs(78)));
    layer0_outputs(5635) <= not((inputs(18)) and (inputs(235)));
    layer0_outputs(5636) <= (inputs(113)) or (inputs(181));
    layer0_outputs(5637) <= not(inputs(90)) or (inputs(224));
    layer0_outputs(5638) <= not((inputs(145)) xor (inputs(130)));
    layer0_outputs(5639) <= inputs(195);
    layer0_outputs(5640) <= inputs(19);
    layer0_outputs(5641) <= not(inputs(29));
    layer0_outputs(5642) <= (inputs(73)) and (inputs(5));
    layer0_outputs(5643) <= inputs(34);
    layer0_outputs(5644) <= inputs(7);
    layer0_outputs(5645) <= not(inputs(62)) or (inputs(50));
    layer0_outputs(5646) <= not(inputs(104));
    layer0_outputs(5647) <= not(inputs(124));
    layer0_outputs(5648) <= (inputs(34)) xor (inputs(212));
    layer0_outputs(5649) <= not(inputs(167)) or (inputs(82));
    layer0_outputs(5650) <= not(inputs(78));
    layer0_outputs(5651) <= '0';
    layer0_outputs(5652) <= not(inputs(124));
    layer0_outputs(5653) <= not(inputs(23));
    layer0_outputs(5654) <= not(inputs(209)) or (inputs(107));
    layer0_outputs(5655) <= (inputs(150)) or (inputs(183));
    layer0_outputs(5656) <= not(inputs(57));
    layer0_outputs(5657) <= not(inputs(119));
    layer0_outputs(5658) <= (inputs(242)) or (inputs(75));
    layer0_outputs(5659) <= (inputs(156)) or (inputs(162));
    layer0_outputs(5660) <= (inputs(244)) and not (inputs(121));
    layer0_outputs(5661) <= not((inputs(103)) or (inputs(167)));
    layer0_outputs(5662) <= '1';
    layer0_outputs(5663) <= (inputs(182)) or (inputs(160));
    layer0_outputs(5664) <= not(inputs(235));
    layer0_outputs(5665) <= '0';
    layer0_outputs(5666) <= not(inputs(60)) or (inputs(129));
    layer0_outputs(5667) <= not((inputs(224)) or (inputs(25)));
    layer0_outputs(5668) <= (inputs(128)) xor (inputs(18));
    layer0_outputs(5669) <= (inputs(229)) and not (inputs(137));
    layer0_outputs(5670) <= (inputs(238)) and (inputs(25));
    layer0_outputs(5671) <= (inputs(230)) or (inputs(247));
    layer0_outputs(5672) <= not(inputs(28)) or (inputs(176));
    layer0_outputs(5673) <= inputs(99);
    layer0_outputs(5674) <= not((inputs(187)) xor (inputs(158)));
    layer0_outputs(5675) <= not(inputs(243));
    layer0_outputs(5676) <= (inputs(13)) or (inputs(100));
    layer0_outputs(5677) <= not((inputs(37)) and (inputs(19)));
    layer0_outputs(5678) <= not(inputs(232));
    layer0_outputs(5679) <= '1';
    layer0_outputs(5680) <= (inputs(94)) or (inputs(67));
    layer0_outputs(5681) <= not((inputs(49)) xor (inputs(16)));
    layer0_outputs(5682) <= not(inputs(25));
    layer0_outputs(5683) <= (inputs(145)) or (inputs(233));
    layer0_outputs(5684) <= not(inputs(47));
    layer0_outputs(5685) <= (inputs(192)) and not (inputs(94));
    layer0_outputs(5686) <= (inputs(104)) and not (inputs(254));
    layer0_outputs(5687) <= inputs(193);
    layer0_outputs(5688) <= not(inputs(56));
    layer0_outputs(5689) <= not((inputs(205)) or (inputs(53)));
    layer0_outputs(5690) <= not((inputs(123)) or (inputs(49)));
    layer0_outputs(5691) <= (inputs(235)) xor (inputs(238));
    layer0_outputs(5692) <= (inputs(86)) or (inputs(117));
    layer0_outputs(5693) <= (inputs(50)) and not (inputs(248));
    layer0_outputs(5694) <= (inputs(62)) xor (inputs(219));
    layer0_outputs(5695) <= (inputs(185)) and (inputs(157));
    layer0_outputs(5696) <= (inputs(90)) and not (inputs(20));
    layer0_outputs(5697) <= (inputs(118)) and (inputs(140));
    layer0_outputs(5698) <= '0';
    layer0_outputs(5699) <= '0';
    layer0_outputs(5700) <= inputs(8);
    layer0_outputs(5701) <= not((inputs(88)) or (inputs(53)));
    layer0_outputs(5702) <= not(inputs(58));
    layer0_outputs(5703) <= not((inputs(35)) xor (inputs(17)));
    layer0_outputs(5704) <= not(inputs(198));
    layer0_outputs(5705) <= not(inputs(131));
    layer0_outputs(5706) <= (inputs(50)) and (inputs(88));
    layer0_outputs(5707) <= inputs(241);
    layer0_outputs(5708) <= inputs(231);
    layer0_outputs(5709) <= not(inputs(135));
    layer0_outputs(5710) <= (inputs(10)) and not (inputs(87));
    layer0_outputs(5711) <= (inputs(101)) or (inputs(227));
    layer0_outputs(5712) <= (inputs(157)) and not (inputs(254));
    layer0_outputs(5713) <= (inputs(239)) and (inputs(6));
    layer0_outputs(5714) <= not(inputs(230)) or (inputs(4));
    layer0_outputs(5715) <= (inputs(125)) or (inputs(248));
    layer0_outputs(5716) <= not(inputs(145)) or (inputs(255));
    layer0_outputs(5717) <= (inputs(56)) xor (inputs(6));
    layer0_outputs(5718) <= inputs(224);
    layer0_outputs(5719) <= (inputs(160)) and not (inputs(28));
    layer0_outputs(5720) <= (inputs(99)) xor (inputs(15));
    layer0_outputs(5721) <= not(inputs(194));
    layer0_outputs(5722) <= not(inputs(84));
    layer0_outputs(5723) <= not((inputs(117)) xor (inputs(103)));
    layer0_outputs(5724) <= (inputs(37)) and not (inputs(102));
    layer0_outputs(5725) <= not(inputs(253));
    layer0_outputs(5726) <= (inputs(154)) and not (inputs(201));
    layer0_outputs(5727) <= '1';
    layer0_outputs(5728) <= inputs(245);
    layer0_outputs(5729) <= not(inputs(90));
    layer0_outputs(5730) <= not(inputs(143));
    layer0_outputs(5731) <= not((inputs(90)) and (inputs(120)));
    layer0_outputs(5732) <= (inputs(75)) and not (inputs(190));
    layer0_outputs(5733) <= not(inputs(127));
    layer0_outputs(5734) <= not(inputs(187));
    layer0_outputs(5735) <= inputs(179);
    layer0_outputs(5736) <= not(inputs(176)) or (inputs(129));
    layer0_outputs(5737) <= not((inputs(179)) xor (inputs(220)));
    layer0_outputs(5738) <= '0';
    layer0_outputs(5739) <= not(inputs(38));
    layer0_outputs(5740) <= inputs(237);
    layer0_outputs(5741) <= (inputs(236)) xor (inputs(182));
    layer0_outputs(5742) <= not(inputs(105));
    layer0_outputs(5743) <= not((inputs(136)) and (inputs(44)));
    layer0_outputs(5744) <= (inputs(126)) and not (inputs(220));
    layer0_outputs(5745) <= (inputs(86)) and not (inputs(242));
    layer0_outputs(5746) <= inputs(222);
    layer0_outputs(5747) <= (inputs(117)) and not (inputs(33));
    layer0_outputs(5748) <= not(inputs(242));
    layer0_outputs(5749) <= inputs(232);
    layer0_outputs(5750) <= inputs(118);
    layer0_outputs(5751) <= (inputs(103)) and not (inputs(251));
    layer0_outputs(5752) <= (inputs(44)) and not (inputs(187));
    layer0_outputs(5753) <= not((inputs(93)) or (inputs(76)));
    layer0_outputs(5754) <= (inputs(165)) and not (inputs(96));
    layer0_outputs(5755) <= not((inputs(231)) xor (inputs(159)));
    layer0_outputs(5756) <= inputs(96);
    layer0_outputs(5757) <= '0';
    layer0_outputs(5758) <= (inputs(87)) and not (inputs(179));
    layer0_outputs(5759) <= (inputs(148)) or (inputs(48));
    layer0_outputs(5760) <= (inputs(214)) xor (inputs(108));
    layer0_outputs(5761) <= (inputs(187)) or (inputs(176));
    layer0_outputs(5762) <= inputs(52);
    layer0_outputs(5763) <= not((inputs(252)) xor (inputs(190)));
    layer0_outputs(5764) <= not(inputs(140));
    layer0_outputs(5765) <= inputs(232);
    layer0_outputs(5766) <= (inputs(126)) and not (inputs(14));
    layer0_outputs(5767) <= not(inputs(118));
    layer0_outputs(5768) <= (inputs(107)) xor (inputs(77));
    layer0_outputs(5769) <= (inputs(247)) and (inputs(149));
    layer0_outputs(5770) <= not(inputs(21)) or (inputs(224));
    layer0_outputs(5771) <= not(inputs(214)) or (inputs(37));
    layer0_outputs(5772) <= not((inputs(223)) or (inputs(227)));
    layer0_outputs(5773) <= (inputs(109)) and not (inputs(9));
    layer0_outputs(5774) <= inputs(145);
    layer0_outputs(5775) <= not(inputs(75)) or (inputs(124));
    layer0_outputs(5776) <= not(inputs(115));
    layer0_outputs(5777) <= (inputs(144)) xor (inputs(174));
    layer0_outputs(5778) <= (inputs(128)) or (inputs(23));
    layer0_outputs(5779) <= '1';
    layer0_outputs(5780) <= not((inputs(117)) xor (inputs(149)));
    layer0_outputs(5781) <= not(inputs(95));
    layer0_outputs(5782) <= not(inputs(193)) or (inputs(65));
    layer0_outputs(5783) <= (inputs(187)) xor (inputs(131));
    layer0_outputs(5784) <= (inputs(242)) xor (inputs(244));
    layer0_outputs(5785) <= not((inputs(158)) or (inputs(110)));
    layer0_outputs(5786) <= inputs(167);
    layer0_outputs(5787) <= not((inputs(87)) xor (inputs(42)));
    layer0_outputs(5788) <= not(inputs(150)) or (inputs(22));
    layer0_outputs(5789) <= not(inputs(125));
    layer0_outputs(5790) <= '0';
    layer0_outputs(5791) <= not(inputs(236));
    layer0_outputs(5792) <= (inputs(103)) or (inputs(241));
    layer0_outputs(5793) <= (inputs(172)) or (inputs(4));
    layer0_outputs(5794) <= '1';
    layer0_outputs(5795) <= '1';
    layer0_outputs(5796) <= not((inputs(195)) and (inputs(141)));
    layer0_outputs(5797) <= not(inputs(38)) or (inputs(179));
    layer0_outputs(5798) <= (inputs(0)) and not (inputs(28));
    layer0_outputs(5799) <= (inputs(124)) and not (inputs(197));
    layer0_outputs(5800) <= (inputs(206)) and not (inputs(43));
    layer0_outputs(5801) <= not(inputs(249));
    layer0_outputs(5802) <= (inputs(1)) or (inputs(210));
    layer0_outputs(5803) <= '1';
    layer0_outputs(5804) <= (inputs(43)) or (inputs(14));
    layer0_outputs(5805) <= not(inputs(212));
    layer0_outputs(5806) <= '0';
    layer0_outputs(5807) <= not(inputs(155));
    layer0_outputs(5808) <= inputs(105);
    layer0_outputs(5809) <= (inputs(30)) xor (inputs(86));
    layer0_outputs(5810) <= (inputs(93)) and (inputs(127));
    layer0_outputs(5811) <= inputs(182);
    layer0_outputs(5812) <= inputs(164);
    layer0_outputs(5813) <= not(inputs(239)) or (inputs(200));
    layer0_outputs(5814) <= inputs(134);
    layer0_outputs(5815) <= inputs(163);
    layer0_outputs(5816) <= (inputs(190)) or (inputs(96));
    layer0_outputs(5817) <= not((inputs(150)) or (inputs(66)));
    layer0_outputs(5818) <= not(inputs(254)) or (inputs(251));
    layer0_outputs(5819) <= not(inputs(165));
    layer0_outputs(5820) <= (inputs(236)) xor (inputs(173));
    layer0_outputs(5821) <= not(inputs(117));
    layer0_outputs(5822) <= (inputs(119)) xor (inputs(74));
    layer0_outputs(5823) <= not(inputs(158)) or (inputs(28));
    layer0_outputs(5824) <= (inputs(157)) xor (inputs(226));
    layer0_outputs(5825) <= (inputs(62)) and not (inputs(14));
    layer0_outputs(5826) <= inputs(152);
    layer0_outputs(5827) <= '1';
    layer0_outputs(5828) <= not(inputs(245)) or (inputs(79));
    layer0_outputs(5829) <= (inputs(79)) or (inputs(125));
    layer0_outputs(5830) <= not(inputs(118));
    layer0_outputs(5831) <= not(inputs(58)) or (inputs(207));
    layer0_outputs(5832) <= not(inputs(85)) or (inputs(240));
    layer0_outputs(5833) <= (inputs(6)) xor (inputs(133));
    layer0_outputs(5834) <= not((inputs(89)) or (inputs(11)));
    layer0_outputs(5835) <= (inputs(190)) and not (inputs(254));
    layer0_outputs(5836) <= not(inputs(27));
    layer0_outputs(5837) <= '0';
    layer0_outputs(5838) <= (inputs(33)) and not (inputs(184));
    layer0_outputs(5839) <= not(inputs(169));
    layer0_outputs(5840) <= (inputs(56)) and not (inputs(35));
    layer0_outputs(5841) <= not((inputs(0)) or (inputs(68)));
    layer0_outputs(5842) <= inputs(48);
    layer0_outputs(5843) <= not(inputs(220));
    layer0_outputs(5844) <= (inputs(73)) and (inputs(196));
    layer0_outputs(5845) <= not((inputs(144)) or (inputs(88)));
    layer0_outputs(5846) <= not(inputs(234));
    layer0_outputs(5847) <= (inputs(28)) and not (inputs(243));
    layer0_outputs(5848) <= not(inputs(228));
    layer0_outputs(5849) <= not((inputs(70)) or (inputs(97)));
    layer0_outputs(5850) <= not(inputs(119));
    layer0_outputs(5851) <= not(inputs(62));
    layer0_outputs(5852) <= (inputs(232)) and not (inputs(36));
    layer0_outputs(5853) <= not((inputs(119)) and (inputs(71)));
    layer0_outputs(5854) <= inputs(77);
    layer0_outputs(5855) <= inputs(164);
    layer0_outputs(5856) <= inputs(167);
    layer0_outputs(5857) <= inputs(247);
    layer0_outputs(5858) <= inputs(63);
    layer0_outputs(5859) <= (inputs(98)) xor (inputs(235));
    layer0_outputs(5860) <= not(inputs(120)) or (inputs(149));
    layer0_outputs(5861) <= not(inputs(114)) or (inputs(134));
    layer0_outputs(5862) <= not((inputs(19)) xor (inputs(38)));
    layer0_outputs(5863) <= not(inputs(44)) or (inputs(117));
    layer0_outputs(5864) <= (inputs(36)) and not (inputs(231));
    layer0_outputs(5865) <= inputs(55);
    layer0_outputs(5866) <= not(inputs(79)) or (inputs(15));
    layer0_outputs(5867) <= not(inputs(178));
    layer0_outputs(5868) <= (inputs(188)) or (inputs(247));
    layer0_outputs(5869) <= inputs(159);
    layer0_outputs(5870) <= not(inputs(54)) or (inputs(92));
    layer0_outputs(5871) <= inputs(237);
    layer0_outputs(5872) <= not(inputs(249)) or (inputs(231));
    layer0_outputs(5873) <= not(inputs(171)) or (inputs(167));
    layer0_outputs(5874) <= inputs(123);
    layer0_outputs(5875) <= (inputs(192)) and not (inputs(208));
    layer0_outputs(5876) <= '1';
    layer0_outputs(5877) <= (inputs(253)) xor (inputs(179));
    layer0_outputs(5878) <= not(inputs(210));
    layer0_outputs(5879) <= (inputs(181)) or (inputs(180));
    layer0_outputs(5880) <= not((inputs(199)) or (inputs(3)));
    layer0_outputs(5881) <= (inputs(7)) and not (inputs(30));
    layer0_outputs(5882) <= not((inputs(220)) or (inputs(180)));
    layer0_outputs(5883) <= '0';
    layer0_outputs(5884) <= not(inputs(78)) or (inputs(234));
    layer0_outputs(5885) <= not(inputs(0)) or (inputs(237));
    layer0_outputs(5886) <= not(inputs(104)) or (inputs(111));
    layer0_outputs(5887) <= (inputs(113)) or (inputs(240));
    layer0_outputs(5888) <= inputs(82);
    layer0_outputs(5889) <= not(inputs(120));
    layer0_outputs(5890) <= not(inputs(85));
    layer0_outputs(5891) <= not((inputs(232)) or (inputs(234)));
    layer0_outputs(5892) <= inputs(35);
    layer0_outputs(5893) <= inputs(54);
    layer0_outputs(5894) <= inputs(180);
    layer0_outputs(5895) <= (inputs(120)) xor (inputs(213));
    layer0_outputs(5896) <= not((inputs(101)) or (inputs(86)));
    layer0_outputs(5897) <= inputs(171);
    layer0_outputs(5898) <= (inputs(168)) and not (inputs(53));
    layer0_outputs(5899) <= not((inputs(177)) or (inputs(116)));
    layer0_outputs(5900) <= inputs(101);
    layer0_outputs(5901) <= inputs(238);
    layer0_outputs(5902) <= (inputs(98)) or (inputs(223));
    layer0_outputs(5903) <= not(inputs(129));
    layer0_outputs(5904) <= not((inputs(86)) xor (inputs(149)));
    layer0_outputs(5905) <= not((inputs(107)) xor (inputs(144)));
    layer0_outputs(5906) <= not(inputs(7)) or (inputs(249));
    layer0_outputs(5907) <= inputs(217);
    layer0_outputs(5908) <= not((inputs(163)) xor (inputs(174)));
    layer0_outputs(5909) <= not((inputs(236)) xor (inputs(255)));
    layer0_outputs(5910) <= '1';
    layer0_outputs(5911) <= inputs(162);
    layer0_outputs(5912) <= (inputs(124)) or (inputs(234));
    layer0_outputs(5913) <= inputs(2);
    layer0_outputs(5914) <= not((inputs(86)) xor (inputs(55)));
    layer0_outputs(5915) <= '0';
    layer0_outputs(5916) <= not(inputs(246));
    layer0_outputs(5917) <= (inputs(140)) or (inputs(174));
    layer0_outputs(5918) <= inputs(80);
    layer0_outputs(5919) <= inputs(148);
    layer0_outputs(5920) <= inputs(45);
    layer0_outputs(5921) <= not((inputs(35)) and (inputs(20)));
    layer0_outputs(5922) <= (inputs(201)) and (inputs(202));
    layer0_outputs(5923) <= (inputs(139)) or (inputs(77));
    layer0_outputs(5924) <= not(inputs(10)) or (inputs(15));
    layer0_outputs(5925) <= not((inputs(235)) or (inputs(2)));
    layer0_outputs(5926) <= (inputs(237)) xor (inputs(179));
    layer0_outputs(5927) <= not(inputs(165));
    layer0_outputs(5928) <= (inputs(117)) and not (inputs(3));
    layer0_outputs(5929) <= '1';
    layer0_outputs(5930) <= not((inputs(60)) or (inputs(176)));
    layer0_outputs(5931) <= (inputs(178)) and not (inputs(128));
    layer0_outputs(5932) <= (inputs(121)) and not (inputs(33));
    layer0_outputs(5933) <= inputs(117);
    layer0_outputs(5934) <= not(inputs(228)) or (inputs(0));
    layer0_outputs(5935) <= (inputs(204)) or (inputs(132));
    layer0_outputs(5936) <= inputs(82);
    layer0_outputs(5937) <= (inputs(69)) or (inputs(15));
    layer0_outputs(5938) <= not((inputs(15)) xor (inputs(168)));
    layer0_outputs(5939) <= not(inputs(60));
    layer0_outputs(5940) <= inputs(98);
    layer0_outputs(5941) <= inputs(197);
    layer0_outputs(5942) <= not(inputs(184));
    layer0_outputs(5943) <= not(inputs(181));
    layer0_outputs(5944) <= inputs(203);
    layer0_outputs(5945) <= inputs(158);
    layer0_outputs(5946) <= (inputs(14)) or (inputs(183));
    layer0_outputs(5947) <= not(inputs(92));
    layer0_outputs(5948) <= not((inputs(246)) or (inputs(66)));
    layer0_outputs(5949) <= not(inputs(211)) or (inputs(166));
    layer0_outputs(5950) <= not((inputs(84)) xor (inputs(113)));
    layer0_outputs(5951) <= not(inputs(39));
    layer0_outputs(5952) <= not(inputs(201)) or (inputs(47));
    layer0_outputs(5953) <= not((inputs(56)) and (inputs(206)));
    layer0_outputs(5954) <= (inputs(177)) or (inputs(162));
    layer0_outputs(5955) <= inputs(228);
    layer0_outputs(5956) <= not(inputs(94));
    layer0_outputs(5957) <= inputs(160);
    layer0_outputs(5958) <= inputs(135);
    layer0_outputs(5959) <= not((inputs(80)) xor (inputs(230)));
    layer0_outputs(5960) <= not(inputs(120)) or (inputs(65));
    layer0_outputs(5961) <= (inputs(91)) and (inputs(40));
    layer0_outputs(5962) <= not(inputs(121)) or (inputs(56));
    layer0_outputs(5963) <= not((inputs(159)) or (inputs(127)));
    layer0_outputs(5964) <= not((inputs(236)) xor (inputs(12)));
    layer0_outputs(5965) <= (inputs(224)) xor (inputs(251));
    layer0_outputs(5966) <= (inputs(42)) and not (inputs(203));
    layer0_outputs(5967) <= inputs(124);
    layer0_outputs(5968) <= not((inputs(177)) xor (inputs(197)));
    layer0_outputs(5969) <= inputs(75);
    layer0_outputs(5970) <= not((inputs(168)) xor (inputs(180)));
    layer0_outputs(5971) <= (inputs(164)) and not (inputs(23));
    layer0_outputs(5972) <= not(inputs(129));
    layer0_outputs(5973) <= inputs(125);
    layer0_outputs(5974) <= not(inputs(23));
    layer0_outputs(5975) <= not((inputs(116)) or (inputs(89)));
    layer0_outputs(5976) <= not(inputs(0)) or (inputs(190));
    layer0_outputs(5977) <= (inputs(115)) xor (inputs(50));
    layer0_outputs(5978) <= (inputs(61)) or (inputs(233));
    layer0_outputs(5979) <= (inputs(124)) or (inputs(44));
    layer0_outputs(5980) <= (inputs(51)) or (inputs(69));
    layer0_outputs(5981) <= not((inputs(37)) or (inputs(123)));
    layer0_outputs(5982) <= (inputs(3)) xor (inputs(134));
    layer0_outputs(5983) <= (inputs(181)) xor (inputs(95));
    layer0_outputs(5984) <= (inputs(103)) and (inputs(135));
    layer0_outputs(5985) <= inputs(212);
    layer0_outputs(5986) <= (inputs(192)) or (inputs(202));
    layer0_outputs(5987) <= inputs(239);
    layer0_outputs(5988) <= inputs(139);
    layer0_outputs(5989) <= not(inputs(232));
    layer0_outputs(5990) <= not((inputs(234)) or (inputs(61)));
    layer0_outputs(5991) <= not((inputs(18)) or (inputs(197)));
    layer0_outputs(5992) <= (inputs(122)) or (inputs(110));
    layer0_outputs(5993) <= (inputs(87)) and not (inputs(215));
    layer0_outputs(5994) <= not(inputs(240));
    layer0_outputs(5995) <= (inputs(196)) and not (inputs(222));
    layer0_outputs(5996) <= not(inputs(199)) or (inputs(152));
    layer0_outputs(5997) <= not((inputs(38)) or (inputs(55)));
    layer0_outputs(5998) <= (inputs(32)) or (inputs(125));
    layer0_outputs(5999) <= not(inputs(89)) or (inputs(121));
    layer0_outputs(6000) <= inputs(233);
    layer0_outputs(6001) <= not(inputs(183));
    layer0_outputs(6002) <= not((inputs(159)) or (inputs(113)));
    layer0_outputs(6003) <= '0';
    layer0_outputs(6004) <= not((inputs(85)) xor (inputs(19)));
    layer0_outputs(6005) <= inputs(70);
    layer0_outputs(6006) <= inputs(120);
    layer0_outputs(6007) <= (inputs(189)) or (inputs(160));
    layer0_outputs(6008) <= not(inputs(87));
    layer0_outputs(6009) <= not(inputs(215));
    layer0_outputs(6010) <= not((inputs(239)) xor (inputs(137)));
    layer0_outputs(6011) <= (inputs(128)) and not (inputs(109));
    layer0_outputs(6012) <= not(inputs(232)) or (inputs(52));
    layer0_outputs(6013) <= inputs(238);
    layer0_outputs(6014) <= (inputs(18)) or (inputs(244));
    layer0_outputs(6015) <= not(inputs(178)) or (inputs(62));
    layer0_outputs(6016) <= not((inputs(125)) or (inputs(180)));
    layer0_outputs(6017) <= not((inputs(158)) and (inputs(60)));
    layer0_outputs(6018) <= not((inputs(246)) or (inputs(130)));
    layer0_outputs(6019) <= (inputs(164)) xor (inputs(233));
    layer0_outputs(6020) <= not(inputs(84));
    layer0_outputs(6021) <= not(inputs(155)) or (inputs(250));
    layer0_outputs(6022) <= not(inputs(111)) or (inputs(46));
    layer0_outputs(6023) <= (inputs(79)) or (inputs(187));
    layer0_outputs(6024) <= inputs(197);
    layer0_outputs(6025) <= not((inputs(165)) or (inputs(48)));
    layer0_outputs(6026) <= (inputs(206)) and not (inputs(201));
    layer0_outputs(6027) <= not(inputs(148));
    layer0_outputs(6028) <= not(inputs(86)) or (inputs(33));
    layer0_outputs(6029) <= (inputs(197)) or (inputs(221));
    layer0_outputs(6030) <= (inputs(143)) and not (inputs(153));
    layer0_outputs(6031) <= inputs(131);
    layer0_outputs(6032) <= not(inputs(93));
    layer0_outputs(6033) <= not(inputs(206)) or (inputs(116));
    layer0_outputs(6034) <= inputs(114);
    layer0_outputs(6035) <= inputs(56);
    layer0_outputs(6036) <= inputs(65);
    layer0_outputs(6037) <= inputs(94);
    layer0_outputs(6038) <= inputs(251);
    layer0_outputs(6039) <= not((inputs(62)) or (inputs(0)));
    layer0_outputs(6040) <= not((inputs(108)) xor (inputs(210)));
    layer0_outputs(6041) <= (inputs(167)) xor (inputs(43));
    layer0_outputs(6042) <= not((inputs(168)) xor (inputs(209)));
    layer0_outputs(6043) <= (inputs(243)) and not (inputs(145));
    layer0_outputs(6044) <= not((inputs(180)) or (inputs(31)));
    layer0_outputs(6045) <= not(inputs(80));
    layer0_outputs(6046) <= not((inputs(153)) xor (inputs(107)));
    layer0_outputs(6047) <= not(inputs(195)) or (inputs(94));
    layer0_outputs(6048) <= not(inputs(4));
    layer0_outputs(6049) <= (inputs(125)) or (inputs(212));
    layer0_outputs(6050) <= not((inputs(196)) xor (inputs(145)));
    layer0_outputs(6051) <= not(inputs(47));
    layer0_outputs(6052) <= (inputs(6)) xor (inputs(176));
    layer0_outputs(6053) <= not((inputs(2)) xor (inputs(224)));
    layer0_outputs(6054) <= not((inputs(166)) xor (inputs(202)));
    layer0_outputs(6055) <= not(inputs(89)) or (inputs(203));
    layer0_outputs(6056) <= not(inputs(96));
    layer0_outputs(6057) <= (inputs(226)) or (inputs(56));
    layer0_outputs(6058) <= inputs(136);
    layer0_outputs(6059) <= not(inputs(57)) or (inputs(151));
    layer0_outputs(6060) <= (inputs(200)) and not (inputs(35));
    layer0_outputs(6061) <= inputs(39);
    layer0_outputs(6062) <= '0';
    layer0_outputs(6063) <= inputs(253);
    layer0_outputs(6064) <= not(inputs(231));
    layer0_outputs(6065) <= not(inputs(28));
    layer0_outputs(6066) <= (inputs(96)) or (inputs(98));
    layer0_outputs(6067) <= (inputs(179)) and not (inputs(125));
    layer0_outputs(6068) <= not((inputs(33)) xor (inputs(67)));
    layer0_outputs(6069) <= not((inputs(169)) or (inputs(161)));
    layer0_outputs(6070) <= not(inputs(79)) or (inputs(1));
    layer0_outputs(6071) <= (inputs(240)) and (inputs(51));
    layer0_outputs(6072) <= not(inputs(133));
    layer0_outputs(6073) <= not((inputs(58)) xor (inputs(23)));
    layer0_outputs(6074) <= (inputs(131)) and not (inputs(85));
    layer0_outputs(6075) <= inputs(88);
    layer0_outputs(6076) <= not((inputs(143)) or (inputs(196)));
    layer0_outputs(6077) <= (inputs(187)) xor (inputs(239));
    layer0_outputs(6078) <= not((inputs(135)) xor (inputs(72)));
    layer0_outputs(6079) <= not(inputs(167));
    layer0_outputs(6080) <= not(inputs(143));
    layer0_outputs(6081) <= inputs(57);
    layer0_outputs(6082) <= inputs(98);
    layer0_outputs(6083) <= (inputs(8)) or (inputs(205));
    layer0_outputs(6084) <= '0';
    layer0_outputs(6085) <= not(inputs(167));
    layer0_outputs(6086) <= (inputs(220)) xor (inputs(128));
    layer0_outputs(6087) <= inputs(167);
    layer0_outputs(6088) <= not(inputs(117)) or (inputs(9));
    layer0_outputs(6089) <= not(inputs(198));
    layer0_outputs(6090) <= '0';
    layer0_outputs(6091) <= inputs(98);
    layer0_outputs(6092) <= (inputs(8)) and (inputs(90));
    layer0_outputs(6093) <= not((inputs(89)) xor (inputs(8)));
    layer0_outputs(6094) <= not((inputs(60)) or (inputs(125)));
    layer0_outputs(6095) <= (inputs(165)) and not (inputs(200));
    layer0_outputs(6096) <= (inputs(107)) and not (inputs(234));
    layer0_outputs(6097) <= not(inputs(42)) or (inputs(230));
    layer0_outputs(6098) <= not(inputs(100));
    layer0_outputs(6099) <= (inputs(57)) or (inputs(134));
    layer0_outputs(6100) <= inputs(100);
    layer0_outputs(6101) <= (inputs(53)) or (inputs(86));
    layer0_outputs(6102) <= not(inputs(204)) or (inputs(49));
    layer0_outputs(6103) <= not(inputs(93)) or (inputs(217));
    layer0_outputs(6104) <= not((inputs(89)) xor (inputs(42)));
    layer0_outputs(6105) <= not(inputs(119)) or (inputs(190));
    layer0_outputs(6106) <= inputs(74);
    layer0_outputs(6107) <= (inputs(90)) and (inputs(76));
    layer0_outputs(6108) <= not(inputs(118));
    layer0_outputs(6109) <= (inputs(43)) and not (inputs(175));
    layer0_outputs(6110) <= (inputs(237)) or (inputs(102));
    layer0_outputs(6111) <= not(inputs(90));
    layer0_outputs(6112) <= (inputs(236)) or (inputs(126));
    layer0_outputs(6113) <= (inputs(178)) or (inputs(48));
    layer0_outputs(6114) <= not((inputs(153)) or (inputs(185)));
    layer0_outputs(6115) <= (inputs(231)) xor (inputs(197));
    layer0_outputs(6116) <= not(inputs(233)) or (inputs(208));
    layer0_outputs(6117) <= not((inputs(99)) or (inputs(100)));
    layer0_outputs(6118) <= not((inputs(208)) or (inputs(188)));
    layer0_outputs(6119) <= not(inputs(155));
    layer0_outputs(6120) <= inputs(46);
    layer0_outputs(6121) <= inputs(194);
    layer0_outputs(6122) <= not(inputs(107));
    layer0_outputs(6123) <= not((inputs(140)) xor (inputs(112)));
    layer0_outputs(6124) <= inputs(137);
    layer0_outputs(6125) <= (inputs(46)) or (inputs(14));
    layer0_outputs(6126) <= not((inputs(152)) and (inputs(101)));
    layer0_outputs(6127) <= not(inputs(98));
    layer0_outputs(6128) <= (inputs(90)) xor (inputs(95));
    layer0_outputs(6129) <= (inputs(88)) and not (inputs(187));
    layer0_outputs(6130) <= inputs(250);
    layer0_outputs(6131) <= inputs(49);
    layer0_outputs(6132) <= (inputs(30)) xor (inputs(157));
    layer0_outputs(6133) <= not((inputs(24)) xor (inputs(206)));
    layer0_outputs(6134) <= inputs(184);
    layer0_outputs(6135) <= not(inputs(69)) or (inputs(123));
    layer0_outputs(6136) <= inputs(32);
    layer0_outputs(6137) <= (inputs(95)) xor (inputs(92));
    layer0_outputs(6138) <= not(inputs(126));
    layer0_outputs(6139) <= not(inputs(191));
    layer0_outputs(6140) <= not(inputs(57));
    layer0_outputs(6141) <= not((inputs(214)) and (inputs(126)));
    layer0_outputs(6142) <= (inputs(142)) or (inputs(137));
    layer0_outputs(6143) <= not(inputs(91));
    layer0_outputs(6144) <= not((inputs(209)) or (inputs(46)));
    layer0_outputs(6145) <= (inputs(232)) xor (inputs(248));
    layer0_outputs(6146) <= (inputs(205)) xor (inputs(87));
    layer0_outputs(6147) <= inputs(206);
    layer0_outputs(6148) <= not((inputs(198)) and (inputs(19)));
    layer0_outputs(6149) <= not(inputs(220)) or (inputs(128));
    layer0_outputs(6150) <= not((inputs(124)) xor (inputs(225)));
    layer0_outputs(6151) <= not(inputs(31));
    layer0_outputs(6152) <= inputs(23);
    layer0_outputs(6153) <= (inputs(163)) or (inputs(93));
    layer0_outputs(6154) <= not(inputs(169));
    layer0_outputs(6155) <= not(inputs(238)) or (inputs(31));
    layer0_outputs(6156) <= not(inputs(233)) or (inputs(139));
    layer0_outputs(6157) <= (inputs(96)) or (inputs(145));
    layer0_outputs(6158) <= inputs(247);
    layer0_outputs(6159) <= not((inputs(150)) or (inputs(183)));
    layer0_outputs(6160) <= not(inputs(142));
    layer0_outputs(6161) <= (inputs(182)) xor (inputs(61));
    layer0_outputs(6162) <= not((inputs(214)) and (inputs(16)));
    layer0_outputs(6163) <= not(inputs(4)) or (inputs(94));
    layer0_outputs(6164) <= not((inputs(129)) xor (inputs(132)));
    layer0_outputs(6165) <= not(inputs(23)) or (inputs(246));
    layer0_outputs(6166) <= not(inputs(59)) or (inputs(254));
    layer0_outputs(6167) <= (inputs(123)) and (inputs(63));
    layer0_outputs(6168) <= inputs(158);
    layer0_outputs(6169) <= (inputs(222)) or (inputs(6));
    layer0_outputs(6170) <= not((inputs(126)) or (inputs(60)));
    layer0_outputs(6171) <= inputs(166);
    layer0_outputs(6172) <= (inputs(65)) or (inputs(139));
    layer0_outputs(6173) <= (inputs(35)) xor (inputs(112));
    layer0_outputs(6174) <= (inputs(54)) or (inputs(209));
    layer0_outputs(6175) <= not(inputs(116));
    layer0_outputs(6176) <= (inputs(255)) xor (inputs(121));
    layer0_outputs(6177) <= not(inputs(204));
    layer0_outputs(6178) <= '1';
    layer0_outputs(6179) <= not((inputs(138)) and (inputs(134)));
    layer0_outputs(6180) <= inputs(184);
    layer0_outputs(6181) <= not((inputs(128)) or (inputs(83)));
    layer0_outputs(6182) <= inputs(6);
    layer0_outputs(6183) <= inputs(185);
    layer0_outputs(6184) <= '0';
    layer0_outputs(6185) <= inputs(86);
    layer0_outputs(6186) <= (inputs(150)) or (inputs(167));
    layer0_outputs(6187) <= not((inputs(20)) and (inputs(10)));
    layer0_outputs(6188) <= inputs(134);
    layer0_outputs(6189) <= not(inputs(192)) or (inputs(180));
    layer0_outputs(6190) <= (inputs(100)) and not (inputs(93));
    layer0_outputs(6191) <= (inputs(112)) and not (inputs(127));
    layer0_outputs(6192) <= inputs(128);
    layer0_outputs(6193) <= not(inputs(14));
    layer0_outputs(6194) <= '0';
    layer0_outputs(6195) <= not((inputs(66)) or (inputs(38)));
    layer0_outputs(6196) <= not((inputs(74)) xor (inputs(223)));
    layer0_outputs(6197) <= not((inputs(210)) or (inputs(36)));
    layer0_outputs(6198) <= not((inputs(244)) and (inputs(199)));
    layer0_outputs(6199) <= not((inputs(192)) and (inputs(189)));
    layer0_outputs(6200) <= (inputs(137)) and not (inputs(21));
    layer0_outputs(6201) <= inputs(231);
    layer0_outputs(6202) <= (inputs(55)) or (inputs(207));
    layer0_outputs(6203) <= not((inputs(125)) or (inputs(141)));
    layer0_outputs(6204) <= inputs(65);
    layer0_outputs(6205) <= not(inputs(70)) or (inputs(239));
    layer0_outputs(6206) <= inputs(200);
    layer0_outputs(6207) <= not((inputs(131)) or (inputs(71)));
    layer0_outputs(6208) <= inputs(88);
    layer0_outputs(6209) <= inputs(83);
    layer0_outputs(6210) <= not(inputs(45));
    layer0_outputs(6211) <= not((inputs(231)) or (inputs(230)));
    layer0_outputs(6212) <= not((inputs(66)) and (inputs(126)));
    layer0_outputs(6213) <= (inputs(19)) xor (inputs(238));
    layer0_outputs(6214) <= not(inputs(95)) or (inputs(34));
    layer0_outputs(6215) <= '0';
    layer0_outputs(6216) <= (inputs(135)) and not (inputs(67));
    layer0_outputs(6217) <= (inputs(106)) or (inputs(13));
    layer0_outputs(6218) <= (inputs(202)) and not (inputs(18));
    layer0_outputs(6219) <= not(inputs(181));
    layer0_outputs(6220) <= not((inputs(208)) and (inputs(201)));
    layer0_outputs(6221) <= not((inputs(76)) and (inputs(92)));
    layer0_outputs(6222) <= (inputs(115)) xor (inputs(30));
    layer0_outputs(6223) <= (inputs(30)) or (inputs(141));
    layer0_outputs(6224) <= not(inputs(83));
    layer0_outputs(6225) <= (inputs(30)) or (inputs(19));
    layer0_outputs(6226) <= not(inputs(182)) or (inputs(50));
    layer0_outputs(6227) <= (inputs(37)) or (inputs(9));
    layer0_outputs(6228) <= not(inputs(221));
    layer0_outputs(6229) <= not(inputs(157)) or (inputs(212));
    layer0_outputs(6230) <= (inputs(72)) and not (inputs(154));
    layer0_outputs(6231) <= (inputs(222)) and not (inputs(66));
    layer0_outputs(6232) <= not((inputs(167)) or (inputs(65)));
    layer0_outputs(6233) <= not(inputs(32));
    layer0_outputs(6234) <= (inputs(22)) and not (inputs(121));
    layer0_outputs(6235) <= not((inputs(23)) and (inputs(0)));
    layer0_outputs(6236) <= not((inputs(224)) or (inputs(108)));
    layer0_outputs(6237) <= not(inputs(227));
    layer0_outputs(6238) <= inputs(88);
    layer0_outputs(6239) <= not((inputs(230)) xor (inputs(207)));
    layer0_outputs(6240) <= not(inputs(133)) or (inputs(172));
    layer0_outputs(6241) <= (inputs(190)) and not (inputs(233));
    layer0_outputs(6242) <= not((inputs(64)) or (inputs(149)));
    layer0_outputs(6243) <= not((inputs(124)) xor (inputs(205)));
    layer0_outputs(6244) <= not((inputs(24)) or (inputs(28)));
    layer0_outputs(6245) <= not(inputs(253));
    layer0_outputs(6246) <= '1';
    layer0_outputs(6247) <= (inputs(18)) or (inputs(247));
    layer0_outputs(6248) <= not(inputs(210)) or (inputs(113));
    layer0_outputs(6249) <= inputs(166);
    layer0_outputs(6250) <= inputs(77);
    layer0_outputs(6251) <= (inputs(167)) or (inputs(138));
    layer0_outputs(6252) <= not(inputs(101)) or (inputs(63));
    layer0_outputs(6253) <= inputs(104);
    layer0_outputs(6254) <= (inputs(132)) xor (inputs(129));
    layer0_outputs(6255) <= not(inputs(213));
    layer0_outputs(6256) <= inputs(232);
    layer0_outputs(6257) <= not(inputs(10)) or (inputs(174));
    layer0_outputs(6258) <= (inputs(125)) or (inputs(206));
    layer0_outputs(6259) <= not(inputs(145));
    layer0_outputs(6260) <= (inputs(159)) and (inputs(190));
    layer0_outputs(6261) <= '0';
    layer0_outputs(6262) <= inputs(225);
    layer0_outputs(6263) <= not((inputs(70)) or (inputs(205)));
    layer0_outputs(6264) <= not((inputs(123)) and (inputs(242)));
    layer0_outputs(6265) <= not((inputs(77)) and (inputs(164)));
    layer0_outputs(6266) <= not(inputs(251));
    layer0_outputs(6267) <= inputs(114);
    layer0_outputs(6268) <= '1';
    layer0_outputs(6269) <= not(inputs(52)) or (inputs(234));
    layer0_outputs(6270) <= (inputs(159)) and not (inputs(253));
    layer0_outputs(6271) <= not(inputs(104)) or (inputs(239));
    layer0_outputs(6272) <= (inputs(140)) and not (inputs(202));
    layer0_outputs(6273) <= not((inputs(173)) xor (inputs(212)));
    layer0_outputs(6274) <= (inputs(52)) and (inputs(143));
    layer0_outputs(6275) <= not(inputs(126));
    layer0_outputs(6276) <= (inputs(91)) and not (inputs(65));
    layer0_outputs(6277) <= not((inputs(151)) or (inputs(252)));
    layer0_outputs(6278) <= not(inputs(159));
    layer0_outputs(6279) <= not(inputs(169));
    layer0_outputs(6280) <= not((inputs(158)) xor (inputs(85)));
    layer0_outputs(6281) <= not((inputs(207)) xor (inputs(219)));
    layer0_outputs(6282) <= not((inputs(179)) xor (inputs(210)));
    layer0_outputs(6283) <= not(inputs(33)) or (inputs(82));
    layer0_outputs(6284) <= not(inputs(35)) or (inputs(216));
    layer0_outputs(6285) <= '0';
    layer0_outputs(6286) <= not(inputs(153)) or (inputs(91));
    layer0_outputs(6287) <= not((inputs(75)) xor (inputs(87)));
    layer0_outputs(6288) <= inputs(112);
    layer0_outputs(6289) <= (inputs(121)) xor (inputs(186));
    layer0_outputs(6290) <= inputs(36);
    layer0_outputs(6291) <= not((inputs(175)) xor (inputs(111)));
    layer0_outputs(6292) <= not((inputs(118)) xor (inputs(197)));
    layer0_outputs(6293) <= '1';
    layer0_outputs(6294) <= (inputs(105)) and not (inputs(111));
    layer0_outputs(6295) <= not(inputs(225)) or (inputs(143));
    layer0_outputs(6296) <= not((inputs(150)) or (inputs(210)));
    layer0_outputs(6297) <= inputs(134);
    layer0_outputs(6298) <= not(inputs(79));
    layer0_outputs(6299) <= not(inputs(182)) or (inputs(91));
    layer0_outputs(6300) <= not(inputs(122)) or (inputs(102));
    layer0_outputs(6301) <= '1';
    layer0_outputs(6302) <= (inputs(240)) or (inputs(125));
    layer0_outputs(6303) <= not(inputs(35));
    layer0_outputs(6304) <= (inputs(233)) xor (inputs(127));
    layer0_outputs(6305) <= inputs(150);
    layer0_outputs(6306) <= (inputs(247)) and not (inputs(224));
    layer0_outputs(6307) <= (inputs(68)) xor (inputs(147));
    layer0_outputs(6308) <= not(inputs(42)) or (inputs(234));
    layer0_outputs(6309) <= not(inputs(38)) or (inputs(147));
    layer0_outputs(6310) <= not((inputs(255)) or (inputs(127)));
    layer0_outputs(6311) <= not((inputs(121)) or (inputs(44)));
    layer0_outputs(6312) <= inputs(226);
    layer0_outputs(6313) <= (inputs(85)) xor (inputs(207));
    layer0_outputs(6314) <= not(inputs(196));
    layer0_outputs(6315) <= (inputs(199)) and (inputs(23));
    layer0_outputs(6316) <= not((inputs(245)) or (inputs(49)));
    layer0_outputs(6317) <= inputs(23);
    layer0_outputs(6318) <= not(inputs(9));
    layer0_outputs(6319) <= '1';
    layer0_outputs(6320) <= not((inputs(246)) or (inputs(143)));
    layer0_outputs(6321) <= not(inputs(67)) or (inputs(251));
    layer0_outputs(6322) <= not(inputs(231));
    layer0_outputs(6323) <= not(inputs(193));
    layer0_outputs(6324) <= not(inputs(114));
    layer0_outputs(6325) <= not((inputs(41)) xor (inputs(101)));
    layer0_outputs(6326) <= not((inputs(108)) xor (inputs(63)));
    layer0_outputs(6327) <= '1';
    layer0_outputs(6328) <= (inputs(25)) and (inputs(80));
    layer0_outputs(6329) <= (inputs(219)) or (inputs(158));
    layer0_outputs(6330) <= (inputs(169)) and not (inputs(120));
    layer0_outputs(6331) <= not((inputs(91)) or (inputs(2)));
    layer0_outputs(6332) <= not((inputs(219)) or (inputs(64)));
    layer0_outputs(6333) <= not(inputs(200)) or (inputs(131));
    layer0_outputs(6334) <= inputs(23);
    layer0_outputs(6335) <= (inputs(188)) and not (inputs(179));
    layer0_outputs(6336) <= not((inputs(128)) xor (inputs(151)));
    layer0_outputs(6337) <= not(inputs(160)) or (inputs(140));
    layer0_outputs(6338) <= (inputs(55)) xor (inputs(84));
    layer0_outputs(6339) <= not((inputs(105)) xor (inputs(124)));
    layer0_outputs(6340) <= inputs(70);
    layer0_outputs(6341) <= not(inputs(230)) or (inputs(106));
    layer0_outputs(6342) <= (inputs(13)) or (inputs(86));
    layer0_outputs(6343) <= (inputs(117)) and not (inputs(222));
    layer0_outputs(6344) <= not(inputs(107));
    layer0_outputs(6345) <= (inputs(61)) and not (inputs(48));
    layer0_outputs(6346) <= inputs(94);
    layer0_outputs(6347) <= (inputs(82)) and not (inputs(55));
    layer0_outputs(6348) <= (inputs(234)) xor (inputs(204));
    layer0_outputs(6349) <= not(inputs(176));
    layer0_outputs(6350) <= inputs(156);
    layer0_outputs(6351) <= '0';
    layer0_outputs(6352) <= not(inputs(138));
    layer0_outputs(6353) <= inputs(10);
    layer0_outputs(6354) <= (inputs(79)) or (inputs(50));
    layer0_outputs(6355) <= (inputs(74)) and not (inputs(144));
    layer0_outputs(6356) <= '1';
    layer0_outputs(6357) <= inputs(73);
    layer0_outputs(6358) <= not(inputs(172)) or (inputs(50));
    layer0_outputs(6359) <= not(inputs(134)) or (inputs(141));
    layer0_outputs(6360) <= inputs(39);
    layer0_outputs(6361) <= inputs(148);
    layer0_outputs(6362) <= not(inputs(37));
    layer0_outputs(6363) <= (inputs(81)) xor (inputs(86));
    layer0_outputs(6364) <= inputs(178);
    layer0_outputs(6365) <= inputs(116);
    layer0_outputs(6366) <= inputs(204);
    layer0_outputs(6367) <= inputs(21);
    layer0_outputs(6368) <= inputs(49);
    layer0_outputs(6369) <= not(inputs(100));
    layer0_outputs(6370) <= not(inputs(164));
    layer0_outputs(6371) <= not(inputs(109));
    layer0_outputs(6372) <= '1';
    layer0_outputs(6373) <= not(inputs(84));
    layer0_outputs(6374) <= (inputs(64)) and not (inputs(68));
    layer0_outputs(6375) <= (inputs(144)) or (inputs(84));
    layer0_outputs(6376) <= inputs(209);
    layer0_outputs(6377) <= (inputs(221)) and not (inputs(141));
    layer0_outputs(6378) <= (inputs(26)) and not (inputs(178));
    layer0_outputs(6379) <= not((inputs(5)) or (inputs(20)));
    layer0_outputs(6380) <= (inputs(140)) xor (inputs(5));
    layer0_outputs(6381) <= (inputs(54)) and not (inputs(255));
    layer0_outputs(6382) <= (inputs(43)) xor (inputs(65));
    layer0_outputs(6383) <= (inputs(134)) or (inputs(172));
    layer0_outputs(6384) <= not(inputs(152));
    layer0_outputs(6385) <= not((inputs(204)) or (inputs(205)));
    layer0_outputs(6386) <= not(inputs(56)) or (inputs(143));
    layer0_outputs(6387) <= not((inputs(5)) xor (inputs(81)));
    layer0_outputs(6388) <= inputs(62);
    layer0_outputs(6389) <= not(inputs(4)) or (inputs(80));
    layer0_outputs(6390) <= (inputs(37)) and not (inputs(113));
    layer0_outputs(6391) <= (inputs(126)) xor (inputs(27));
    layer0_outputs(6392) <= not(inputs(62)) or (inputs(173));
    layer0_outputs(6393) <= not(inputs(230));
    layer0_outputs(6394) <= (inputs(64)) or (inputs(209));
    layer0_outputs(6395) <= not((inputs(157)) xor (inputs(94)));
    layer0_outputs(6396) <= not((inputs(164)) or (inputs(83)));
    layer0_outputs(6397) <= not((inputs(0)) or (inputs(73)));
    layer0_outputs(6398) <= not(inputs(39));
    layer0_outputs(6399) <= (inputs(29)) xor (inputs(192));
    layer0_outputs(6400) <= not((inputs(238)) or (inputs(30)));
    layer0_outputs(6401) <= not((inputs(5)) or (inputs(89)));
    layer0_outputs(6402) <= (inputs(171)) and not (inputs(169));
    layer0_outputs(6403) <= not((inputs(79)) xor (inputs(92)));
    layer0_outputs(6404) <= (inputs(29)) and not (inputs(55));
    layer0_outputs(6405) <= (inputs(175)) and not (inputs(14));
    layer0_outputs(6406) <= inputs(169);
    layer0_outputs(6407) <= not(inputs(172)) or (inputs(30));
    layer0_outputs(6408) <= not((inputs(221)) or (inputs(17)));
    layer0_outputs(6409) <= inputs(25);
    layer0_outputs(6410) <= inputs(183);
    layer0_outputs(6411) <= not(inputs(184)) or (inputs(18));
    layer0_outputs(6412) <= not(inputs(11));
    layer0_outputs(6413) <= inputs(163);
    layer0_outputs(6414) <= not(inputs(68));
    layer0_outputs(6415) <= inputs(113);
    layer0_outputs(6416) <= (inputs(187)) and not (inputs(33));
    layer0_outputs(6417) <= not((inputs(85)) xor (inputs(223)));
    layer0_outputs(6418) <= (inputs(233)) or (inputs(223));
    layer0_outputs(6419) <= inputs(24);
    layer0_outputs(6420) <= inputs(117);
    layer0_outputs(6421) <= (inputs(216)) and not (inputs(98));
    layer0_outputs(6422) <= (inputs(235)) or (inputs(185));
    layer0_outputs(6423) <= (inputs(234)) and not (inputs(79));
    layer0_outputs(6424) <= (inputs(148)) or (inputs(5));
    layer0_outputs(6425) <= not(inputs(161));
    layer0_outputs(6426) <= '1';
    layer0_outputs(6427) <= inputs(64);
    layer0_outputs(6428) <= not(inputs(128));
    layer0_outputs(6429) <= (inputs(221)) or (inputs(92));
    layer0_outputs(6430) <= '1';
    layer0_outputs(6431) <= (inputs(117)) and not (inputs(47));
    layer0_outputs(6432) <= (inputs(148)) and not (inputs(91));
    layer0_outputs(6433) <= (inputs(89)) and not (inputs(219));
    layer0_outputs(6434) <= not(inputs(140)) or (inputs(36));
    layer0_outputs(6435) <= (inputs(234)) and not (inputs(114));
    layer0_outputs(6436) <= not(inputs(63));
    layer0_outputs(6437) <= (inputs(101)) and not (inputs(127));
    layer0_outputs(6438) <= inputs(26);
    layer0_outputs(6439) <= not(inputs(220)) or (inputs(66));
    layer0_outputs(6440) <= not(inputs(54)) or (inputs(126));
    layer0_outputs(6441) <= not(inputs(163)) or (inputs(81));
    layer0_outputs(6442) <= inputs(248);
    layer0_outputs(6443) <= inputs(138);
    layer0_outputs(6444) <= not(inputs(68)) or (inputs(48));
    layer0_outputs(6445) <= not(inputs(241));
    layer0_outputs(6446) <= (inputs(31)) or (inputs(164));
    layer0_outputs(6447) <= not(inputs(160));
    layer0_outputs(6448) <= not(inputs(196));
    layer0_outputs(6449) <= '0';
    layer0_outputs(6450) <= not(inputs(116)) or (inputs(237));
    layer0_outputs(6451) <= not((inputs(184)) or (inputs(131)));
    layer0_outputs(6452) <= not((inputs(251)) or (inputs(243)));
    layer0_outputs(6453) <= not(inputs(218)) or (inputs(110));
    layer0_outputs(6454) <= (inputs(63)) or (inputs(2));
    layer0_outputs(6455) <= not((inputs(80)) or (inputs(221)));
    layer0_outputs(6456) <= (inputs(138)) and not (inputs(10));
    layer0_outputs(6457) <= not(inputs(127)) or (inputs(29));
    layer0_outputs(6458) <= (inputs(253)) xor (inputs(19));
    layer0_outputs(6459) <= not(inputs(115));
    layer0_outputs(6460) <= not((inputs(188)) xor (inputs(219)));
    layer0_outputs(6461) <= inputs(80);
    layer0_outputs(6462) <= inputs(83);
    layer0_outputs(6463) <= inputs(27);
    layer0_outputs(6464) <= inputs(8);
    layer0_outputs(6465) <= not((inputs(236)) xor (inputs(178)));
    layer0_outputs(6466) <= not((inputs(88)) or (inputs(59)));
    layer0_outputs(6467) <= not(inputs(25));
    layer0_outputs(6468) <= (inputs(144)) xor (inputs(205));
    layer0_outputs(6469) <= not(inputs(142)) or (inputs(153));
    layer0_outputs(6470) <= not((inputs(28)) or (inputs(21)));
    layer0_outputs(6471) <= inputs(126);
    layer0_outputs(6472) <= not((inputs(202)) xor (inputs(220)));
    layer0_outputs(6473) <= not((inputs(228)) or (inputs(99)));
    layer0_outputs(6474) <= (inputs(138)) xor (inputs(139));
    layer0_outputs(6475) <= (inputs(243)) xor (inputs(212));
    layer0_outputs(6476) <= (inputs(224)) xor (inputs(172));
    layer0_outputs(6477) <= (inputs(172)) or (inputs(31));
    layer0_outputs(6478) <= (inputs(157)) and not (inputs(131));
    layer0_outputs(6479) <= inputs(32);
    layer0_outputs(6480) <= not(inputs(54));
    layer0_outputs(6481) <= not(inputs(165)) or (inputs(242));
    layer0_outputs(6482) <= inputs(43);
    layer0_outputs(6483) <= not((inputs(25)) xor (inputs(49)));
    layer0_outputs(6484) <= not(inputs(1)) or (inputs(169));
    layer0_outputs(6485) <= (inputs(213)) or (inputs(250));
    layer0_outputs(6486) <= not((inputs(115)) and (inputs(212)));
    layer0_outputs(6487) <= (inputs(246)) and not (inputs(107));
    layer0_outputs(6488) <= (inputs(87)) or (inputs(86));
    layer0_outputs(6489) <= (inputs(74)) xor (inputs(171));
    layer0_outputs(6490) <= (inputs(125)) or (inputs(92));
    layer0_outputs(6491) <= (inputs(231)) xor (inputs(125));
    layer0_outputs(6492) <= (inputs(11)) or (inputs(51));
    layer0_outputs(6493) <= inputs(223);
    layer0_outputs(6494) <= inputs(169);
    layer0_outputs(6495) <= (inputs(22)) xor (inputs(64));
    layer0_outputs(6496) <= inputs(174);
    layer0_outputs(6497) <= '0';
    layer0_outputs(6498) <= inputs(214);
    layer0_outputs(6499) <= (inputs(161)) xor (inputs(231));
    layer0_outputs(6500) <= not((inputs(176)) xor (inputs(227)));
    layer0_outputs(6501) <= not((inputs(53)) xor (inputs(7)));
    layer0_outputs(6502) <= not(inputs(28));
    layer0_outputs(6503) <= not(inputs(207)) or (inputs(133));
    layer0_outputs(6504) <= (inputs(236)) or (inputs(118));
    layer0_outputs(6505) <= (inputs(68)) or (inputs(13));
    layer0_outputs(6506) <= (inputs(119)) or (inputs(167));
    layer0_outputs(6507) <= not((inputs(253)) and (inputs(128)));
    layer0_outputs(6508) <= (inputs(44)) or (inputs(169));
    layer0_outputs(6509) <= not((inputs(213)) or (inputs(191)));
    layer0_outputs(6510) <= (inputs(127)) and not (inputs(191));
    layer0_outputs(6511) <= not((inputs(90)) or (inputs(16)));
    layer0_outputs(6512) <= not((inputs(207)) or (inputs(204)));
    layer0_outputs(6513) <= inputs(142);
    layer0_outputs(6514) <= inputs(42);
    layer0_outputs(6515) <= (inputs(205)) or (inputs(217));
    layer0_outputs(6516) <= not((inputs(243)) or (inputs(109)));
    layer0_outputs(6517) <= inputs(91);
    layer0_outputs(6518) <= '1';
    layer0_outputs(6519) <= (inputs(180)) xor (inputs(182));
    layer0_outputs(6520) <= (inputs(53)) xor (inputs(38));
    layer0_outputs(6521) <= not((inputs(91)) and (inputs(140)));
    layer0_outputs(6522) <= '1';
    layer0_outputs(6523) <= (inputs(36)) and not (inputs(252));
    layer0_outputs(6524) <= inputs(75);
    layer0_outputs(6525) <= inputs(94);
    layer0_outputs(6526) <= inputs(58);
    layer0_outputs(6527) <= not(inputs(165)) or (inputs(191));
    layer0_outputs(6528) <= not((inputs(185)) or (inputs(252)));
    layer0_outputs(6529) <= (inputs(126)) or (inputs(81));
    layer0_outputs(6530) <= not((inputs(99)) or (inputs(98)));
    layer0_outputs(6531) <= '0';
    layer0_outputs(6532) <= inputs(101);
    layer0_outputs(6533) <= not((inputs(18)) xor (inputs(105)));
    layer0_outputs(6534) <= not(inputs(66));
    layer0_outputs(6535) <= (inputs(189)) and not (inputs(204));
    layer0_outputs(6536) <= not(inputs(249));
    layer0_outputs(6537) <= not(inputs(72));
    layer0_outputs(6538) <= not(inputs(178));
    layer0_outputs(6539) <= inputs(20);
    layer0_outputs(6540) <= (inputs(255)) xor (inputs(102));
    layer0_outputs(6541) <= not(inputs(213)) or (inputs(31));
    layer0_outputs(6542) <= (inputs(39)) xor (inputs(116));
    layer0_outputs(6543) <= (inputs(44)) and not (inputs(11));
    layer0_outputs(6544) <= not(inputs(77));
    layer0_outputs(6545) <= not((inputs(33)) or (inputs(45)));
    layer0_outputs(6546) <= not(inputs(245)) or (inputs(53));
    layer0_outputs(6547) <= (inputs(102)) and not (inputs(254));
    layer0_outputs(6548) <= not(inputs(43));
    layer0_outputs(6549) <= not(inputs(253));
    layer0_outputs(6550) <= inputs(213);
    layer0_outputs(6551) <= not(inputs(212));
    layer0_outputs(6552) <= not((inputs(244)) or (inputs(187)));
    layer0_outputs(6553) <= not(inputs(120)) or (inputs(178));
    layer0_outputs(6554) <= (inputs(227)) and not (inputs(107));
    layer0_outputs(6555) <= '0';
    layer0_outputs(6556) <= (inputs(169)) xor (inputs(106));
    layer0_outputs(6557) <= not((inputs(201)) or (inputs(97)));
    layer0_outputs(6558) <= not((inputs(65)) or (inputs(166)));
    layer0_outputs(6559) <= inputs(72);
    layer0_outputs(6560) <= not(inputs(7)) or (inputs(239));
    layer0_outputs(6561) <= inputs(219);
    layer0_outputs(6562) <= not((inputs(17)) or (inputs(187)));
    layer0_outputs(6563) <= not(inputs(143));
    layer0_outputs(6564) <= not(inputs(23)) or (inputs(20));
    layer0_outputs(6565) <= (inputs(107)) xor (inputs(105));
    layer0_outputs(6566) <= '1';
    layer0_outputs(6567) <= (inputs(41)) or (inputs(145));
    layer0_outputs(6568) <= inputs(193);
    layer0_outputs(6569) <= (inputs(51)) or (inputs(165));
    layer0_outputs(6570) <= (inputs(226)) and (inputs(200));
    layer0_outputs(6571) <= inputs(199);
    layer0_outputs(6572) <= not(inputs(100));
    layer0_outputs(6573) <= inputs(119);
    layer0_outputs(6574) <= not(inputs(105));
    layer0_outputs(6575) <= inputs(112);
    layer0_outputs(6576) <= inputs(76);
    layer0_outputs(6577) <= not((inputs(61)) xor (inputs(254)));
    layer0_outputs(6578) <= not((inputs(57)) or (inputs(157)));
    layer0_outputs(6579) <= not(inputs(127));
    layer0_outputs(6580) <= not((inputs(83)) or (inputs(63)));
    layer0_outputs(6581) <= inputs(60);
    layer0_outputs(6582) <= (inputs(179)) or (inputs(157));
    layer0_outputs(6583) <= not(inputs(76)) or (inputs(229));
    layer0_outputs(6584) <= not((inputs(198)) xor (inputs(228)));
    layer0_outputs(6585) <= inputs(0);
    layer0_outputs(6586) <= (inputs(248)) and not (inputs(43));
    layer0_outputs(6587) <= (inputs(24)) and not (inputs(113));
    layer0_outputs(6588) <= inputs(181);
    layer0_outputs(6589) <= not(inputs(84));
    layer0_outputs(6590) <= not(inputs(130));
    layer0_outputs(6591) <= (inputs(52)) and (inputs(139));
    layer0_outputs(6592) <= not(inputs(101));
    layer0_outputs(6593) <= not(inputs(6)) or (inputs(80));
    layer0_outputs(6594) <= '1';
    layer0_outputs(6595) <= not(inputs(18)) or (inputs(95));
    layer0_outputs(6596) <= (inputs(74)) or (inputs(142));
    layer0_outputs(6597) <= (inputs(177)) xor (inputs(246));
    layer0_outputs(6598) <= (inputs(121)) and not (inputs(239));
    layer0_outputs(6599) <= inputs(195);
    layer0_outputs(6600) <= not(inputs(218));
    layer0_outputs(6601) <= not(inputs(9));
    layer0_outputs(6602) <= inputs(213);
    layer0_outputs(6603) <= not(inputs(54)) or (inputs(106));
    layer0_outputs(6604) <= not(inputs(135)) or (inputs(195));
    layer0_outputs(6605) <= (inputs(112)) and not (inputs(47));
    layer0_outputs(6606) <= not(inputs(242)) or (inputs(43));
    layer0_outputs(6607) <= (inputs(162)) and not (inputs(63));
    layer0_outputs(6608) <= not((inputs(194)) and (inputs(120)));
    layer0_outputs(6609) <= '0';
    layer0_outputs(6610) <= (inputs(71)) and (inputs(19));
    layer0_outputs(6611) <= not((inputs(147)) or (inputs(219)));
    layer0_outputs(6612) <= not((inputs(90)) or (inputs(75)));
    layer0_outputs(6613) <= (inputs(179)) or (inputs(43));
    layer0_outputs(6614) <= (inputs(111)) xor (inputs(26));
    layer0_outputs(6615) <= '1';
    layer0_outputs(6616) <= not(inputs(226)) or (inputs(139));
    layer0_outputs(6617) <= not(inputs(137)) or (inputs(93));
    layer0_outputs(6618) <= (inputs(219)) and (inputs(239));
    layer0_outputs(6619) <= not(inputs(43));
    layer0_outputs(6620) <= not((inputs(170)) or (inputs(131)));
    layer0_outputs(6621) <= not(inputs(40));
    layer0_outputs(6622) <= inputs(114);
    layer0_outputs(6623) <= (inputs(0)) xor (inputs(247));
    layer0_outputs(6624) <= not((inputs(160)) xor (inputs(92)));
    layer0_outputs(6625) <= not((inputs(171)) xor (inputs(155)));
    layer0_outputs(6626) <= (inputs(190)) and not (inputs(66));
    layer0_outputs(6627) <= not((inputs(52)) or (inputs(228)));
    layer0_outputs(6628) <= (inputs(18)) xor (inputs(202));
    layer0_outputs(6629) <= not((inputs(232)) or (inputs(51)));
    layer0_outputs(6630) <= not(inputs(178));
    layer0_outputs(6631) <= inputs(102);
    layer0_outputs(6632) <= not(inputs(173));
    layer0_outputs(6633) <= not(inputs(103));
    layer0_outputs(6634) <= not((inputs(93)) or (inputs(218)));
    layer0_outputs(6635) <= (inputs(137)) and (inputs(10));
    layer0_outputs(6636) <= inputs(122);
    layer0_outputs(6637) <= not((inputs(221)) xor (inputs(157)));
    layer0_outputs(6638) <= (inputs(86)) xor (inputs(144));
    layer0_outputs(6639) <= (inputs(106)) and not (inputs(182));
    layer0_outputs(6640) <= (inputs(162)) xor (inputs(245));
    layer0_outputs(6641) <= (inputs(227)) and not (inputs(150));
    layer0_outputs(6642) <= not((inputs(53)) or (inputs(65)));
    layer0_outputs(6643) <= inputs(168);
    layer0_outputs(6644) <= not((inputs(250)) and (inputs(189)));
    layer0_outputs(6645) <= (inputs(14)) and not (inputs(199));
    layer0_outputs(6646) <= not((inputs(72)) and (inputs(108)));
    layer0_outputs(6647) <= not((inputs(162)) or (inputs(92)));
    layer0_outputs(6648) <= not(inputs(58));
    layer0_outputs(6649) <= inputs(122);
    layer0_outputs(6650) <= (inputs(22)) xor (inputs(101));
    layer0_outputs(6651) <= inputs(129);
    layer0_outputs(6652) <= not(inputs(85));
    layer0_outputs(6653) <= not(inputs(181));
    layer0_outputs(6654) <= inputs(231);
    layer0_outputs(6655) <= not(inputs(56));
    layer0_outputs(6656) <= not(inputs(130));
    layer0_outputs(6657) <= not(inputs(127));
    layer0_outputs(6658) <= (inputs(94)) and (inputs(52));
    layer0_outputs(6659) <= not(inputs(181));
    layer0_outputs(6660) <= (inputs(254)) and not (inputs(56));
    layer0_outputs(6661) <= not(inputs(67));
    layer0_outputs(6662) <= not(inputs(124));
    layer0_outputs(6663) <= inputs(132);
    layer0_outputs(6664) <= inputs(228);
    layer0_outputs(6665) <= not(inputs(20));
    layer0_outputs(6666) <= inputs(137);
    layer0_outputs(6667) <= not(inputs(7));
    layer0_outputs(6668) <= (inputs(75)) and not (inputs(136));
    layer0_outputs(6669) <= not((inputs(202)) or (inputs(110)));
    layer0_outputs(6670) <= not((inputs(146)) or (inputs(30)));
    layer0_outputs(6671) <= inputs(108);
    layer0_outputs(6672) <= inputs(208);
    layer0_outputs(6673) <= inputs(121);
    layer0_outputs(6674) <= (inputs(105)) or (inputs(155));
    layer0_outputs(6675) <= not((inputs(74)) or (inputs(80)));
    layer0_outputs(6676) <= not(inputs(129));
    layer0_outputs(6677) <= (inputs(174)) and not (inputs(46));
    layer0_outputs(6678) <= not((inputs(211)) or (inputs(57)));
    layer0_outputs(6679) <= inputs(55);
    layer0_outputs(6680) <= '1';
    layer0_outputs(6681) <= not(inputs(64));
    layer0_outputs(6682) <= inputs(20);
    layer0_outputs(6683) <= not((inputs(3)) or (inputs(154)));
    layer0_outputs(6684) <= not(inputs(245));
    layer0_outputs(6685) <= (inputs(172)) or (inputs(238));
    layer0_outputs(6686) <= not((inputs(109)) xor (inputs(34)));
    layer0_outputs(6687) <= not((inputs(18)) xor (inputs(26)));
    layer0_outputs(6688) <= not((inputs(97)) xor (inputs(102)));
    layer0_outputs(6689) <= (inputs(188)) or (inputs(144));
    layer0_outputs(6690) <= (inputs(188)) xor (inputs(189));
    layer0_outputs(6691) <= (inputs(79)) xor (inputs(2));
    layer0_outputs(6692) <= not((inputs(150)) or (inputs(52)));
    layer0_outputs(6693) <= (inputs(206)) or (inputs(230));
    layer0_outputs(6694) <= '0';
    layer0_outputs(6695) <= inputs(218);
    layer0_outputs(6696) <= not((inputs(37)) or (inputs(77)));
    layer0_outputs(6697) <= not(inputs(24));
    layer0_outputs(6698) <= inputs(84);
    layer0_outputs(6699) <= not((inputs(90)) xor (inputs(242)));
    layer0_outputs(6700) <= (inputs(225)) or (inputs(205));
    layer0_outputs(6701) <= not(inputs(52)) or (inputs(83));
    layer0_outputs(6702) <= inputs(172);
    layer0_outputs(6703) <= not(inputs(2));
    layer0_outputs(6704) <= not(inputs(193));
    layer0_outputs(6705) <= not((inputs(188)) or (inputs(210)));
    layer0_outputs(6706) <= not(inputs(9));
    layer0_outputs(6707) <= (inputs(162)) or (inputs(152));
    layer0_outputs(6708) <= (inputs(115)) or (inputs(117));
    layer0_outputs(6709) <= not((inputs(0)) xor (inputs(118)));
    layer0_outputs(6710) <= (inputs(230)) xor (inputs(168));
    layer0_outputs(6711) <= (inputs(252)) or (inputs(116));
    layer0_outputs(6712) <= (inputs(70)) or (inputs(172));
    layer0_outputs(6713) <= (inputs(120)) or (inputs(30));
    layer0_outputs(6714) <= '0';
    layer0_outputs(6715) <= inputs(22);
    layer0_outputs(6716) <= not(inputs(62));
    layer0_outputs(6717) <= not(inputs(107)) or (inputs(127));
    layer0_outputs(6718) <= (inputs(198)) and not (inputs(63));
    layer0_outputs(6719) <= inputs(23);
    layer0_outputs(6720) <= not(inputs(109));
    layer0_outputs(6721) <= (inputs(83)) or (inputs(38));
    layer0_outputs(6722) <= (inputs(77)) xor (inputs(228));
    layer0_outputs(6723) <= (inputs(0)) and not (inputs(6));
    layer0_outputs(6724) <= inputs(194);
    layer0_outputs(6725) <= (inputs(249)) or (inputs(56));
    layer0_outputs(6726) <= inputs(83);
    layer0_outputs(6727) <= not(inputs(187));
    layer0_outputs(6728) <= inputs(173);
    layer0_outputs(6729) <= not(inputs(118)) or (inputs(6));
    layer0_outputs(6730) <= not((inputs(42)) xor (inputs(11)));
    layer0_outputs(6731) <= not((inputs(239)) or (inputs(70)));
    layer0_outputs(6732) <= inputs(140);
    layer0_outputs(6733) <= (inputs(20)) and not (inputs(224));
    layer0_outputs(6734) <= not((inputs(9)) xor (inputs(111)));
    layer0_outputs(6735) <= not((inputs(38)) xor (inputs(160)));
    layer0_outputs(6736) <= (inputs(243)) xor (inputs(169));
    layer0_outputs(6737) <= inputs(163);
    layer0_outputs(6738) <= not(inputs(187)) or (inputs(0));
    layer0_outputs(6739) <= inputs(214);
    layer0_outputs(6740) <= not((inputs(177)) xor (inputs(22)));
    layer0_outputs(6741) <= not(inputs(54));
    layer0_outputs(6742) <= not((inputs(0)) and (inputs(159)));
    layer0_outputs(6743) <= not(inputs(61));
    layer0_outputs(6744) <= (inputs(120)) and not (inputs(1));
    layer0_outputs(6745) <= not((inputs(252)) xor (inputs(89)));
    layer0_outputs(6746) <= (inputs(24)) and not (inputs(222));
    layer0_outputs(6747) <= not(inputs(200)) or (inputs(46));
    layer0_outputs(6748) <= '0';
    layer0_outputs(6749) <= (inputs(90)) or (inputs(73));
    layer0_outputs(6750) <= (inputs(171)) and (inputs(181));
    layer0_outputs(6751) <= (inputs(108)) and not (inputs(47));
    layer0_outputs(6752) <= inputs(200);
    layer0_outputs(6753) <= (inputs(97)) xor (inputs(71));
    layer0_outputs(6754) <= (inputs(44)) or (inputs(15));
    layer0_outputs(6755) <= (inputs(95)) or (inputs(193));
    layer0_outputs(6756) <= not((inputs(228)) xor (inputs(155)));
    layer0_outputs(6757) <= not((inputs(147)) or (inputs(20)));
    layer0_outputs(6758) <= inputs(94);
    layer0_outputs(6759) <= not((inputs(110)) and (inputs(139)));
    layer0_outputs(6760) <= not(inputs(151));
    layer0_outputs(6761) <= (inputs(123)) and (inputs(18));
    layer0_outputs(6762) <= (inputs(101)) and (inputs(171));
    layer0_outputs(6763) <= not(inputs(36)) or (inputs(0));
    layer0_outputs(6764) <= (inputs(23)) xor (inputs(51));
    layer0_outputs(6765) <= not(inputs(179)) or (inputs(135));
    layer0_outputs(6766) <= not(inputs(207)) or (inputs(201));
    layer0_outputs(6767) <= (inputs(36)) and not (inputs(216));
    layer0_outputs(6768) <= not(inputs(90)) or (inputs(161));
    layer0_outputs(6769) <= (inputs(88)) and (inputs(240));
    layer0_outputs(6770) <= not(inputs(211));
    layer0_outputs(6771) <= not(inputs(253));
    layer0_outputs(6772) <= (inputs(57)) and (inputs(126));
    layer0_outputs(6773) <= inputs(170);
    layer0_outputs(6774) <= not(inputs(162));
    layer0_outputs(6775) <= (inputs(6)) and (inputs(71));
    layer0_outputs(6776) <= (inputs(178)) and (inputs(139));
    layer0_outputs(6777) <= (inputs(244)) or (inputs(11));
    layer0_outputs(6778) <= inputs(51);
    layer0_outputs(6779) <= inputs(108);
    layer0_outputs(6780) <= not((inputs(5)) or (inputs(78)));
    layer0_outputs(6781) <= not(inputs(99));
    layer0_outputs(6782) <= not((inputs(247)) xor (inputs(237)));
    layer0_outputs(6783) <= (inputs(25)) or (inputs(35));
    layer0_outputs(6784) <= (inputs(156)) and not (inputs(135));
    layer0_outputs(6785) <= not((inputs(2)) or (inputs(29)));
    layer0_outputs(6786) <= not((inputs(90)) or (inputs(4)));
    layer0_outputs(6787) <= not((inputs(105)) or (inputs(153)));
    layer0_outputs(6788) <= (inputs(23)) and not (inputs(96));
    layer0_outputs(6789) <= (inputs(196)) and not (inputs(78));
    layer0_outputs(6790) <= not((inputs(95)) and (inputs(139)));
    layer0_outputs(6791) <= '1';
    layer0_outputs(6792) <= not(inputs(125));
    layer0_outputs(6793) <= (inputs(178)) and not (inputs(18));
    layer0_outputs(6794) <= not(inputs(29));
    layer0_outputs(6795) <= inputs(223);
    layer0_outputs(6796) <= (inputs(172)) and (inputs(248));
    layer0_outputs(6797) <= (inputs(104)) xor (inputs(89));
    layer0_outputs(6798) <= not(inputs(65));
    layer0_outputs(6799) <= not(inputs(169));
    layer0_outputs(6800) <= not(inputs(107));
    layer0_outputs(6801) <= (inputs(137)) and (inputs(68));
    layer0_outputs(6802) <= (inputs(61)) or (inputs(39));
    layer0_outputs(6803) <= (inputs(247)) xor (inputs(18));
    layer0_outputs(6804) <= inputs(108);
    layer0_outputs(6805) <= inputs(182);
    layer0_outputs(6806) <= not(inputs(39));
    layer0_outputs(6807) <= '1';
    layer0_outputs(6808) <= not(inputs(133)) or (inputs(70));
    layer0_outputs(6809) <= (inputs(157)) or (inputs(205));
    layer0_outputs(6810) <= (inputs(99)) or (inputs(96));
    layer0_outputs(6811) <= not(inputs(36));
    layer0_outputs(6812) <= (inputs(163)) and not (inputs(107));
    layer0_outputs(6813) <= (inputs(193)) or (inputs(194));
    layer0_outputs(6814) <= not((inputs(253)) xor (inputs(144)));
    layer0_outputs(6815) <= (inputs(193)) xor (inputs(229));
    layer0_outputs(6816) <= not((inputs(12)) or (inputs(163)));
    layer0_outputs(6817) <= not(inputs(114));
    layer0_outputs(6818) <= inputs(82);
    layer0_outputs(6819) <= (inputs(18)) or (inputs(199));
    layer0_outputs(6820) <= (inputs(186)) and not (inputs(16));
    layer0_outputs(6821) <= not((inputs(182)) or (inputs(66)));
    layer0_outputs(6822) <= not((inputs(23)) or (inputs(94)));
    layer0_outputs(6823) <= not((inputs(80)) xor (inputs(9)));
    layer0_outputs(6824) <= not(inputs(44));
    layer0_outputs(6825) <= not((inputs(203)) and (inputs(90)));
    layer0_outputs(6826) <= inputs(94);
    layer0_outputs(6827) <= not((inputs(217)) or (inputs(116)));
    layer0_outputs(6828) <= not((inputs(67)) xor (inputs(69)));
    layer0_outputs(6829) <= not(inputs(189));
    layer0_outputs(6830) <= (inputs(194)) and not (inputs(21));
    layer0_outputs(6831) <= inputs(194);
    layer0_outputs(6832) <= inputs(247);
    layer0_outputs(6833) <= (inputs(187)) xor (inputs(161));
    layer0_outputs(6834) <= (inputs(17)) or (inputs(71));
    layer0_outputs(6835) <= (inputs(167)) and (inputs(41));
    layer0_outputs(6836) <= not(inputs(191));
    layer0_outputs(6837) <= not((inputs(218)) xor (inputs(15)));
    layer0_outputs(6838) <= not((inputs(197)) xor (inputs(229)));
    layer0_outputs(6839) <= '0';
    layer0_outputs(6840) <= not((inputs(182)) xor (inputs(162)));
    layer0_outputs(6841) <= not(inputs(50)) or (inputs(217));
    layer0_outputs(6842) <= not(inputs(95));
    layer0_outputs(6843) <= (inputs(60)) xor (inputs(22));
    layer0_outputs(6844) <= not(inputs(45));
    layer0_outputs(6845) <= not(inputs(35));
    layer0_outputs(6846) <= (inputs(129)) xor (inputs(74));
    layer0_outputs(6847) <= inputs(92);
    layer0_outputs(6848) <= not(inputs(75));
    layer0_outputs(6849) <= '1';
    layer0_outputs(6850) <= not(inputs(1));
    layer0_outputs(6851) <= not((inputs(208)) xor (inputs(189)));
    layer0_outputs(6852) <= not((inputs(227)) xor (inputs(96)));
    layer0_outputs(6853) <= not(inputs(169));
    layer0_outputs(6854) <= not(inputs(248));
    layer0_outputs(6855) <= (inputs(238)) or (inputs(253));
    layer0_outputs(6856) <= not((inputs(203)) or (inputs(228)));
    layer0_outputs(6857) <= (inputs(198)) and not (inputs(116));
    layer0_outputs(6858) <= (inputs(22)) xor (inputs(83));
    layer0_outputs(6859) <= not((inputs(29)) or (inputs(228)));
    layer0_outputs(6860) <= not(inputs(67));
    layer0_outputs(6861) <= not(inputs(158)) or (inputs(157));
    layer0_outputs(6862) <= not(inputs(158));
    layer0_outputs(6863) <= not((inputs(13)) or (inputs(4)));
    layer0_outputs(6864) <= (inputs(238)) and not (inputs(157));
    layer0_outputs(6865) <= (inputs(68)) xor (inputs(195));
    layer0_outputs(6866) <= (inputs(204)) and not (inputs(200));
    layer0_outputs(6867) <= (inputs(173)) and not (inputs(199));
    layer0_outputs(6868) <= (inputs(95)) or (inputs(177));
    layer0_outputs(6869) <= inputs(1);
    layer0_outputs(6870) <= (inputs(210)) or (inputs(51));
    layer0_outputs(6871) <= not(inputs(136)) or (inputs(147));
    layer0_outputs(6872) <= not((inputs(234)) or (inputs(160)));
    layer0_outputs(6873) <= not((inputs(18)) or (inputs(36)));
    layer0_outputs(6874) <= not((inputs(19)) or (inputs(51)));
    layer0_outputs(6875) <= inputs(238);
    layer0_outputs(6876) <= not((inputs(46)) or (inputs(205)));
    layer0_outputs(6877) <= (inputs(182)) and not (inputs(40));
    layer0_outputs(6878) <= not(inputs(57));
    layer0_outputs(6879) <= not(inputs(216));
    layer0_outputs(6880) <= '1';
    layer0_outputs(6881) <= not((inputs(94)) or (inputs(41)));
    layer0_outputs(6882) <= inputs(84);
    layer0_outputs(6883) <= (inputs(134)) and not (inputs(140));
    layer0_outputs(6884) <= (inputs(209)) and not (inputs(119));
    layer0_outputs(6885) <= not((inputs(25)) xor (inputs(55)));
    layer0_outputs(6886) <= (inputs(159)) and (inputs(159));
    layer0_outputs(6887) <= '0';
    layer0_outputs(6888) <= not(inputs(123)) or (inputs(46));
    layer0_outputs(6889) <= '1';
    layer0_outputs(6890) <= not(inputs(91));
    layer0_outputs(6891) <= '1';
    layer0_outputs(6892) <= not(inputs(217));
    layer0_outputs(6893) <= not(inputs(78)) or (inputs(236));
    layer0_outputs(6894) <= inputs(215);
    layer0_outputs(6895) <= (inputs(132)) and not (inputs(172));
    layer0_outputs(6896) <= not((inputs(107)) or (inputs(60)));
    layer0_outputs(6897) <= (inputs(150)) or (inputs(70));
    layer0_outputs(6898) <= not(inputs(249));
    layer0_outputs(6899) <= not((inputs(224)) or (inputs(136)));
    layer0_outputs(6900) <= not(inputs(3)) or (inputs(233));
    layer0_outputs(6901) <= not(inputs(101)) or (inputs(191));
    layer0_outputs(6902) <= (inputs(19)) and not (inputs(254));
    layer0_outputs(6903) <= not((inputs(100)) or (inputs(56)));
    layer0_outputs(6904) <= (inputs(79)) or (inputs(211));
    layer0_outputs(6905) <= (inputs(229)) xor (inputs(167));
    layer0_outputs(6906) <= not(inputs(243));
    layer0_outputs(6907) <= (inputs(107)) and (inputs(92));
    layer0_outputs(6908) <= (inputs(23)) or (inputs(109));
    layer0_outputs(6909) <= inputs(197);
    layer0_outputs(6910) <= '0';
    layer0_outputs(6911) <= not((inputs(233)) or (inputs(226)));
    layer0_outputs(6912) <= '1';
    layer0_outputs(6913) <= not(inputs(55));
    layer0_outputs(6914) <= (inputs(179)) or (inputs(34));
    layer0_outputs(6915) <= not(inputs(114)) or (inputs(74));
    layer0_outputs(6916) <= (inputs(176)) or (inputs(103));
    layer0_outputs(6917) <= not(inputs(94));
    layer0_outputs(6918) <= not(inputs(228));
    layer0_outputs(6919) <= not((inputs(201)) xor (inputs(191)));
    layer0_outputs(6920) <= not((inputs(202)) or (inputs(178)));
    layer0_outputs(6921) <= (inputs(22)) and not (inputs(158));
    layer0_outputs(6922) <= not(inputs(79));
    layer0_outputs(6923) <= not(inputs(28));
    layer0_outputs(6924) <= '1';
    layer0_outputs(6925) <= (inputs(100)) or (inputs(187));
    layer0_outputs(6926) <= not(inputs(41)) or (inputs(93));
    layer0_outputs(6927) <= (inputs(80)) xor (inputs(193));
    layer0_outputs(6928) <= not((inputs(42)) or (inputs(27)));
    layer0_outputs(6929) <= (inputs(134)) and (inputs(104));
    layer0_outputs(6930) <= not((inputs(240)) xor (inputs(127)));
    layer0_outputs(6931) <= not(inputs(129));
    layer0_outputs(6932) <= not((inputs(23)) and (inputs(158)));
    layer0_outputs(6933) <= '0';
    layer0_outputs(6934) <= (inputs(18)) or (inputs(181));
    layer0_outputs(6935) <= inputs(125);
    layer0_outputs(6936) <= (inputs(69)) or (inputs(56));
    layer0_outputs(6937) <= not(inputs(116)) or (inputs(245));
    layer0_outputs(6938) <= inputs(255);
    layer0_outputs(6939) <= inputs(129);
    layer0_outputs(6940) <= not(inputs(145));
    layer0_outputs(6941) <= '0';
    layer0_outputs(6942) <= inputs(27);
    layer0_outputs(6943) <= (inputs(14)) and not (inputs(211));
    layer0_outputs(6944) <= not((inputs(162)) xor (inputs(215)));
    layer0_outputs(6945) <= not(inputs(54));
    layer0_outputs(6946) <= (inputs(207)) or (inputs(227));
    layer0_outputs(6947) <= not(inputs(118));
    layer0_outputs(6948) <= not(inputs(121));
    layer0_outputs(6949) <= (inputs(231)) and (inputs(224));
    layer0_outputs(6950) <= (inputs(254)) xor (inputs(93));
    layer0_outputs(6951) <= not(inputs(234));
    layer0_outputs(6952) <= not(inputs(220));
    layer0_outputs(6953) <= (inputs(47)) or (inputs(4));
    layer0_outputs(6954) <= inputs(216);
    layer0_outputs(6955) <= (inputs(34)) or (inputs(151));
    layer0_outputs(6956) <= (inputs(159)) or (inputs(197));
    layer0_outputs(6957) <= inputs(203);
    layer0_outputs(6958) <= (inputs(210)) and not (inputs(40));
    layer0_outputs(6959) <= not(inputs(239));
    layer0_outputs(6960) <= not(inputs(232)) or (inputs(6));
    layer0_outputs(6961) <= not(inputs(168));
    layer0_outputs(6962) <= '1';
    layer0_outputs(6963) <= not((inputs(56)) xor (inputs(4)));
    layer0_outputs(6964) <= not(inputs(14));
    layer0_outputs(6965) <= (inputs(111)) and (inputs(55));
    layer0_outputs(6966) <= not((inputs(139)) xor (inputs(120)));
    layer0_outputs(6967) <= not(inputs(200));
    layer0_outputs(6968) <= inputs(73);
    layer0_outputs(6969) <= not((inputs(175)) or (inputs(204)));
    layer0_outputs(6970) <= inputs(144);
    layer0_outputs(6971) <= not(inputs(196));
    layer0_outputs(6972) <= not(inputs(218));
    layer0_outputs(6973) <= not(inputs(151)) or (inputs(139));
    layer0_outputs(6974) <= not(inputs(100)) or (inputs(88));
    layer0_outputs(6975) <= not(inputs(56)) or (inputs(237));
    layer0_outputs(6976) <= (inputs(230)) and not (inputs(224));
    layer0_outputs(6977) <= not((inputs(236)) or (inputs(104)));
    layer0_outputs(6978) <= (inputs(116)) and not (inputs(169));
    layer0_outputs(6979) <= (inputs(101)) and (inputs(92));
    layer0_outputs(6980) <= not((inputs(142)) or (inputs(85)));
    layer0_outputs(6981) <= inputs(92);
    layer0_outputs(6982) <= not(inputs(39)) or (inputs(127));
    layer0_outputs(6983) <= (inputs(107)) xor (inputs(73));
    layer0_outputs(6984) <= not(inputs(11)) or (inputs(72));
    layer0_outputs(6985) <= (inputs(177)) xor (inputs(8));
    layer0_outputs(6986) <= not(inputs(213)) or (inputs(13));
    layer0_outputs(6987) <= not(inputs(153));
    layer0_outputs(6988) <= (inputs(10)) or (inputs(97));
    layer0_outputs(6989) <= inputs(21);
    layer0_outputs(6990) <= (inputs(213)) or (inputs(135));
    layer0_outputs(6991) <= inputs(143);
    layer0_outputs(6992) <= (inputs(26)) xor (inputs(32));
    layer0_outputs(6993) <= not(inputs(38));
    layer0_outputs(6994) <= (inputs(70)) or (inputs(111));
    layer0_outputs(6995) <= not((inputs(204)) or (inputs(112)));
    layer0_outputs(6996) <= not(inputs(231));
    layer0_outputs(6997) <= (inputs(211)) and not (inputs(60));
    layer0_outputs(6998) <= inputs(122);
    layer0_outputs(6999) <= (inputs(44)) xor (inputs(196));
    layer0_outputs(7000) <= not(inputs(155));
    layer0_outputs(7001) <= (inputs(177)) and not (inputs(150));
    layer0_outputs(7002) <= not(inputs(243)) or (inputs(107));
    layer0_outputs(7003) <= (inputs(208)) and not (inputs(64));
    layer0_outputs(7004) <= not((inputs(163)) xor (inputs(196)));
    layer0_outputs(7005) <= not(inputs(184));
    layer0_outputs(7006) <= not((inputs(244)) and (inputs(189)));
    layer0_outputs(7007) <= not(inputs(4)) or (inputs(65));
    layer0_outputs(7008) <= not(inputs(164));
    layer0_outputs(7009) <= not(inputs(107)) or (inputs(193));
    layer0_outputs(7010) <= not((inputs(204)) xor (inputs(65)));
    layer0_outputs(7011) <= not(inputs(47));
    layer0_outputs(7012) <= not(inputs(195)) or (inputs(121));
    layer0_outputs(7013) <= not(inputs(244)) or (inputs(158));
    layer0_outputs(7014) <= (inputs(231)) and not (inputs(119));
    layer0_outputs(7015) <= inputs(253);
    layer0_outputs(7016) <= not((inputs(64)) and (inputs(255)));
    layer0_outputs(7017) <= not((inputs(194)) or (inputs(129)));
    layer0_outputs(7018) <= not((inputs(207)) or (inputs(187)));
    layer0_outputs(7019) <= (inputs(50)) or (inputs(105));
    layer0_outputs(7020) <= not(inputs(65)) or (inputs(245));
    layer0_outputs(7021) <= inputs(101);
    layer0_outputs(7022) <= not(inputs(125)) or (inputs(231));
    layer0_outputs(7023) <= '1';
    layer0_outputs(7024) <= not(inputs(135)) or (inputs(238));
    layer0_outputs(7025) <= (inputs(253)) or (inputs(1));
    layer0_outputs(7026) <= not(inputs(241)) or (inputs(211));
    layer0_outputs(7027) <= not(inputs(106));
    layer0_outputs(7028) <= not(inputs(172));
    layer0_outputs(7029) <= not(inputs(76));
    layer0_outputs(7030) <= not(inputs(6)) or (inputs(218));
    layer0_outputs(7031) <= not(inputs(198)) or (inputs(98));
    layer0_outputs(7032) <= not(inputs(188));
    layer0_outputs(7033) <= not((inputs(48)) and (inputs(12)));
    layer0_outputs(7034) <= (inputs(25)) or (inputs(225));
    layer0_outputs(7035) <= (inputs(116)) and not (inputs(34));
    layer0_outputs(7036) <= not(inputs(152));
    layer0_outputs(7037) <= (inputs(125)) and not (inputs(110));
    layer0_outputs(7038) <= (inputs(15)) and (inputs(185));
    layer0_outputs(7039) <= inputs(93);
    layer0_outputs(7040) <= inputs(86);
    layer0_outputs(7041) <= not((inputs(251)) and (inputs(19)));
    layer0_outputs(7042) <= not((inputs(50)) or (inputs(195)));
    layer0_outputs(7043) <= not(inputs(116));
    layer0_outputs(7044) <= not((inputs(51)) xor (inputs(23)));
    layer0_outputs(7045) <= not((inputs(87)) or (inputs(101)));
    layer0_outputs(7046) <= (inputs(35)) xor (inputs(147));
    layer0_outputs(7047) <= not((inputs(212)) or (inputs(46)));
    layer0_outputs(7048) <= not(inputs(113)) or (inputs(235));
    layer0_outputs(7049) <= not(inputs(241));
    layer0_outputs(7050) <= not((inputs(68)) or (inputs(78)));
    layer0_outputs(7051) <= inputs(54);
    layer0_outputs(7052) <= (inputs(52)) or (inputs(52));
    layer0_outputs(7053) <= inputs(50);
    layer0_outputs(7054) <= not(inputs(196)) or (inputs(78));
    layer0_outputs(7055) <= inputs(208);
    layer0_outputs(7056) <= (inputs(187)) and (inputs(54));
    layer0_outputs(7057) <= (inputs(184)) and not (inputs(42));
    layer0_outputs(7058) <= (inputs(27)) xor (inputs(168));
    layer0_outputs(7059) <= (inputs(65)) and (inputs(39));
    layer0_outputs(7060) <= (inputs(28)) and (inputs(149));
    layer0_outputs(7061) <= not(inputs(148));
    layer0_outputs(7062) <= (inputs(97)) or (inputs(10));
    layer0_outputs(7063) <= (inputs(34)) and not (inputs(196));
    layer0_outputs(7064) <= (inputs(27)) and not (inputs(195));
    layer0_outputs(7065) <= not(inputs(180)) or (inputs(14));
    layer0_outputs(7066) <= not(inputs(229)) or (inputs(163));
    layer0_outputs(7067) <= not(inputs(141)) or (inputs(50));
    layer0_outputs(7068) <= (inputs(166)) or (inputs(178));
    layer0_outputs(7069) <= not(inputs(210));
    layer0_outputs(7070) <= not(inputs(190)) or (inputs(12));
    layer0_outputs(7071) <= inputs(183);
    layer0_outputs(7072) <= not(inputs(244)) or (inputs(15));
    layer0_outputs(7073) <= not(inputs(14));
    layer0_outputs(7074) <= not((inputs(48)) xor (inputs(69)));
    layer0_outputs(7075) <= not(inputs(119));
    layer0_outputs(7076) <= (inputs(140)) and not (inputs(175));
    layer0_outputs(7077) <= not(inputs(151));
    layer0_outputs(7078) <= (inputs(177)) and not (inputs(239));
    layer0_outputs(7079) <= not(inputs(83));
    layer0_outputs(7080) <= (inputs(249)) or (inputs(229));
    layer0_outputs(7081) <= not((inputs(192)) xor (inputs(206)));
    layer0_outputs(7082) <= not((inputs(43)) xor (inputs(71)));
    layer0_outputs(7083) <= (inputs(36)) or (inputs(247));
    layer0_outputs(7084) <= not(inputs(224));
    layer0_outputs(7085) <= (inputs(3)) and not (inputs(142));
    layer0_outputs(7086) <= (inputs(41)) and (inputs(60));
    layer0_outputs(7087) <= not((inputs(75)) or (inputs(7)));
    layer0_outputs(7088) <= not(inputs(169));
    layer0_outputs(7089) <= (inputs(76)) xor (inputs(159));
    layer0_outputs(7090) <= not(inputs(194));
    layer0_outputs(7091) <= not((inputs(97)) xor (inputs(129)));
    layer0_outputs(7092) <= not((inputs(73)) or (inputs(74)));
    layer0_outputs(7093) <= not((inputs(87)) xor (inputs(43)));
    layer0_outputs(7094) <= not((inputs(66)) or (inputs(67)));
    layer0_outputs(7095) <= '1';
    layer0_outputs(7096) <= (inputs(47)) xor (inputs(5));
    layer0_outputs(7097) <= (inputs(250)) or (inputs(144));
    layer0_outputs(7098) <= (inputs(43)) and not (inputs(159));
    layer0_outputs(7099) <= not(inputs(213));
    layer0_outputs(7100) <= inputs(170);
    layer0_outputs(7101) <= (inputs(139)) and (inputs(45));
    layer0_outputs(7102) <= not(inputs(12));
    layer0_outputs(7103) <= inputs(202);
    layer0_outputs(7104) <= not(inputs(89));
    layer0_outputs(7105) <= not((inputs(145)) or (inputs(191)));
    layer0_outputs(7106) <= not(inputs(47));
    layer0_outputs(7107) <= not((inputs(116)) or (inputs(77)));
    layer0_outputs(7108) <= not((inputs(70)) or (inputs(93)));
    layer0_outputs(7109) <= not((inputs(123)) and (inputs(251)));
    layer0_outputs(7110) <= not(inputs(20));
    layer0_outputs(7111) <= (inputs(130)) or (inputs(34));
    layer0_outputs(7112) <= (inputs(1)) or (inputs(116));
    layer0_outputs(7113) <= not((inputs(124)) or (inputs(130)));
    layer0_outputs(7114) <= (inputs(136)) and not (inputs(203));
    layer0_outputs(7115) <= (inputs(12)) or (inputs(79));
    layer0_outputs(7116) <= (inputs(100)) and (inputs(116));
    layer0_outputs(7117) <= not((inputs(59)) and (inputs(82)));
    layer0_outputs(7118) <= (inputs(11)) and (inputs(5));
    layer0_outputs(7119) <= not(inputs(3));
    layer0_outputs(7120) <= inputs(190);
    layer0_outputs(7121) <= not((inputs(164)) xor (inputs(222)));
    layer0_outputs(7122) <= (inputs(80)) and not (inputs(212));
    layer0_outputs(7123) <= (inputs(12)) and not (inputs(162));
    layer0_outputs(7124) <= not(inputs(18)) or (inputs(127));
    layer0_outputs(7125) <= (inputs(176)) and not (inputs(226));
    layer0_outputs(7126) <= not(inputs(61)) or (inputs(16));
    layer0_outputs(7127) <= not(inputs(130));
    layer0_outputs(7128) <= (inputs(74)) and (inputs(236));
    layer0_outputs(7129) <= inputs(221);
    layer0_outputs(7130) <= not(inputs(27)) or (inputs(200));
    layer0_outputs(7131) <= inputs(92);
    layer0_outputs(7132) <= not(inputs(145)) or (inputs(235));
    layer0_outputs(7133) <= (inputs(9)) xor (inputs(219));
    layer0_outputs(7134) <= not(inputs(226));
    layer0_outputs(7135) <= inputs(249);
    layer0_outputs(7136) <= not((inputs(22)) xor (inputs(68)));
    layer0_outputs(7137) <= (inputs(21)) or (inputs(171));
    layer0_outputs(7138) <= not(inputs(157));
    layer0_outputs(7139) <= (inputs(85)) or (inputs(35));
    layer0_outputs(7140) <= not(inputs(86));
    layer0_outputs(7141) <= not(inputs(206));
    layer0_outputs(7142) <= not(inputs(172));
    layer0_outputs(7143) <= (inputs(193)) and not (inputs(216));
    layer0_outputs(7144) <= (inputs(97)) and (inputs(5));
    layer0_outputs(7145) <= (inputs(109)) and not (inputs(151));
    layer0_outputs(7146) <= inputs(158);
    layer0_outputs(7147) <= not(inputs(199));
    layer0_outputs(7148) <= (inputs(124)) and (inputs(48));
    layer0_outputs(7149) <= (inputs(207)) or (inputs(232));
    layer0_outputs(7150) <= inputs(4);
    layer0_outputs(7151) <= not(inputs(202)) or (inputs(94));
    layer0_outputs(7152) <= not(inputs(138));
    layer0_outputs(7153) <= (inputs(219)) and (inputs(201));
    layer0_outputs(7154) <= inputs(134);
    layer0_outputs(7155) <= (inputs(254)) xor (inputs(35));
    layer0_outputs(7156) <= not(inputs(67));
    layer0_outputs(7157) <= (inputs(188)) xor (inputs(252));
    layer0_outputs(7158) <= '1';
    layer0_outputs(7159) <= not((inputs(186)) and (inputs(167)));
    layer0_outputs(7160) <= not((inputs(157)) or (inputs(156)));
    layer0_outputs(7161) <= inputs(0);
    layer0_outputs(7162) <= not(inputs(150)) or (inputs(76));
    layer0_outputs(7163) <= not(inputs(182)) or (inputs(132));
    layer0_outputs(7164) <= inputs(194);
    layer0_outputs(7165) <= inputs(85);
    layer0_outputs(7166) <= (inputs(41)) xor (inputs(165));
    layer0_outputs(7167) <= (inputs(42)) and not (inputs(24));
    layer0_outputs(7168) <= not(inputs(179));
    layer0_outputs(7169) <= not(inputs(206)) or (inputs(49));
    layer0_outputs(7170) <= (inputs(69)) and not (inputs(32));
    layer0_outputs(7171) <= not(inputs(175));
    layer0_outputs(7172) <= (inputs(71)) and not (inputs(51));
    layer0_outputs(7173) <= not(inputs(197)) or (inputs(31));
    layer0_outputs(7174) <= not(inputs(141)) or (inputs(33));
    layer0_outputs(7175) <= (inputs(244)) xor (inputs(212));
    layer0_outputs(7176) <= '0';
    layer0_outputs(7177) <= not((inputs(217)) and (inputs(39)));
    layer0_outputs(7178) <= '0';
    layer0_outputs(7179) <= inputs(54);
    layer0_outputs(7180) <= (inputs(220)) xor (inputs(174));
    layer0_outputs(7181) <= not(inputs(187)) or (inputs(10));
    layer0_outputs(7182) <= not(inputs(140)) or (inputs(108));
    layer0_outputs(7183) <= inputs(62);
    layer0_outputs(7184) <= not(inputs(123));
    layer0_outputs(7185) <= (inputs(131)) or (inputs(206));
    layer0_outputs(7186) <= (inputs(245)) xor (inputs(143));
    layer0_outputs(7187) <= not(inputs(187));
    layer0_outputs(7188) <= inputs(196);
    layer0_outputs(7189) <= not((inputs(49)) or (inputs(43)));
    layer0_outputs(7190) <= not(inputs(240)) or (inputs(166));
    layer0_outputs(7191) <= inputs(209);
    layer0_outputs(7192) <= not(inputs(86));
    layer0_outputs(7193) <= (inputs(51)) and not (inputs(240));
    layer0_outputs(7194) <= not(inputs(37)) or (inputs(194));
    layer0_outputs(7195) <= not((inputs(44)) or (inputs(92)));
    layer0_outputs(7196) <= inputs(170);
    layer0_outputs(7197) <= (inputs(126)) xor (inputs(123));
    layer0_outputs(7198) <= inputs(140);
    layer0_outputs(7199) <= inputs(184);
    layer0_outputs(7200) <= not((inputs(154)) or (inputs(103)));
    layer0_outputs(7201) <= (inputs(36)) or (inputs(79));
    layer0_outputs(7202) <= not((inputs(205)) and (inputs(170)));
    layer0_outputs(7203) <= not(inputs(185));
    layer0_outputs(7204) <= (inputs(9)) and not (inputs(197));
    layer0_outputs(7205) <= (inputs(231)) and (inputs(227));
    layer0_outputs(7206) <= (inputs(93)) or (inputs(27));
    layer0_outputs(7207) <= (inputs(251)) and not (inputs(72));
    layer0_outputs(7208) <= not(inputs(196)) or (inputs(161));
    layer0_outputs(7209) <= not(inputs(136)) or (inputs(172));
    layer0_outputs(7210) <= (inputs(55)) or (inputs(109));
    layer0_outputs(7211) <= (inputs(148)) or (inputs(15));
    layer0_outputs(7212) <= '0';
    layer0_outputs(7213) <= not(inputs(171));
    layer0_outputs(7214) <= not(inputs(53));
    layer0_outputs(7215) <= not((inputs(189)) xor (inputs(187)));
    layer0_outputs(7216) <= (inputs(4)) xor (inputs(79));
    layer0_outputs(7217) <= inputs(59);
    layer0_outputs(7218) <= not(inputs(101));
    layer0_outputs(7219) <= not(inputs(224)) or (inputs(169));
    layer0_outputs(7220) <= not((inputs(65)) xor (inputs(141)));
    layer0_outputs(7221) <= (inputs(11)) or (inputs(12));
    layer0_outputs(7222) <= (inputs(148)) or (inputs(216));
    layer0_outputs(7223) <= not(inputs(81)) or (inputs(139));
    layer0_outputs(7224) <= not((inputs(45)) and (inputs(210)));
    layer0_outputs(7225) <= not((inputs(24)) xor (inputs(147)));
    layer0_outputs(7226) <= not(inputs(54));
    layer0_outputs(7227) <= (inputs(242)) and not (inputs(215));
    layer0_outputs(7228) <= not(inputs(129)) or (inputs(140));
    layer0_outputs(7229) <= not(inputs(28)) or (inputs(184));
    layer0_outputs(7230) <= inputs(200);
    layer0_outputs(7231) <= (inputs(132)) xor (inputs(51));
    layer0_outputs(7232) <= not(inputs(250));
    layer0_outputs(7233) <= not(inputs(109)) or (inputs(83));
    layer0_outputs(7234) <= not((inputs(110)) or (inputs(33)));
    layer0_outputs(7235) <= (inputs(17)) or (inputs(100));
    layer0_outputs(7236) <= (inputs(212)) and not (inputs(221));
    layer0_outputs(7237) <= not(inputs(165));
    layer0_outputs(7238) <= not(inputs(172));
    layer0_outputs(7239) <= not(inputs(101)) or (inputs(63));
    layer0_outputs(7240) <= not((inputs(197)) xor (inputs(213)));
    layer0_outputs(7241) <= not((inputs(63)) and (inputs(3)));
    layer0_outputs(7242) <= not(inputs(109));
    layer0_outputs(7243) <= not(inputs(45));
    layer0_outputs(7244) <= not(inputs(180));
    layer0_outputs(7245) <= not(inputs(64));
    layer0_outputs(7246) <= (inputs(152)) or (inputs(175));
    layer0_outputs(7247) <= (inputs(88)) xor (inputs(119));
    layer0_outputs(7248) <= inputs(171);
    layer0_outputs(7249) <= (inputs(204)) and (inputs(219));
    layer0_outputs(7250) <= (inputs(8)) or (inputs(154));
    layer0_outputs(7251) <= not((inputs(168)) xor (inputs(62)));
    layer0_outputs(7252) <= not((inputs(48)) and (inputs(0)));
    layer0_outputs(7253) <= not(inputs(25));
    layer0_outputs(7254) <= not(inputs(26)) or (inputs(17));
    layer0_outputs(7255) <= (inputs(183)) and not (inputs(172));
    layer0_outputs(7256) <= not(inputs(135)) or (inputs(76));
    layer0_outputs(7257) <= (inputs(71)) or (inputs(223));
    layer0_outputs(7258) <= (inputs(18)) or (inputs(16));
    layer0_outputs(7259) <= not(inputs(121)) or (inputs(20));
    layer0_outputs(7260) <= (inputs(190)) xor (inputs(209));
    layer0_outputs(7261) <= inputs(106);
    layer0_outputs(7262) <= not(inputs(12)) or (inputs(176));
    layer0_outputs(7263) <= (inputs(2)) and (inputs(254));
    layer0_outputs(7264) <= (inputs(137)) and not (inputs(95));
    layer0_outputs(7265) <= inputs(0);
    layer0_outputs(7266) <= not(inputs(67));
    layer0_outputs(7267) <= (inputs(7)) and not (inputs(217));
    layer0_outputs(7268) <= inputs(118);
    layer0_outputs(7269) <= not(inputs(162));
    layer0_outputs(7270) <= not(inputs(68));
    layer0_outputs(7271) <= (inputs(81)) or (inputs(143));
    layer0_outputs(7272) <= not(inputs(102)) or (inputs(176));
    layer0_outputs(7273) <= inputs(110);
    layer0_outputs(7274) <= inputs(22);
    layer0_outputs(7275) <= (inputs(19)) and not (inputs(211));
    layer0_outputs(7276) <= (inputs(96)) xor (inputs(53));
    layer0_outputs(7277) <= (inputs(92)) or (inputs(53));
    layer0_outputs(7278) <= '1';
    layer0_outputs(7279) <= (inputs(161)) xor (inputs(8));
    layer0_outputs(7280) <= (inputs(27)) and not (inputs(61));
    layer0_outputs(7281) <= (inputs(250)) and not (inputs(238));
    layer0_outputs(7282) <= not(inputs(132));
    layer0_outputs(7283) <= not(inputs(196)) or (inputs(3));
    layer0_outputs(7284) <= not(inputs(147)) or (inputs(66));
    layer0_outputs(7285) <= not((inputs(223)) xor (inputs(123)));
    layer0_outputs(7286) <= not(inputs(184));
    layer0_outputs(7287) <= not((inputs(199)) and (inputs(201)));
    layer0_outputs(7288) <= not(inputs(91)) or (inputs(160));
    layer0_outputs(7289) <= not(inputs(11)) or (inputs(117));
    layer0_outputs(7290) <= not(inputs(193));
    layer0_outputs(7291) <= not((inputs(48)) or (inputs(14)));
    layer0_outputs(7292) <= not(inputs(18));
    layer0_outputs(7293) <= (inputs(96)) or (inputs(168));
    layer0_outputs(7294) <= not((inputs(122)) or (inputs(137)));
    layer0_outputs(7295) <= inputs(138);
    layer0_outputs(7296) <= inputs(211);
    layer0_outputs(7297) <= not(inputs(135)) or (inputs(108));
    layer0_outputs(7298) <= (inputs(254)) and not (inputs(36));
    layer0_outputs(7299) <= inputs(106);
    layer0_outputs(7300) <= not((inputs(110)) and (inputs(203)));
    layer0_outputs(7301) <= (inputs(72)) and not (inputs(93));
    layer0_outputs(7302) <= (inputs(8)) and not (inputs(3));
    layer0_outputs(7303) <= (inputs(142)) xor (inputs(19));
    layer0_outputs(7304) <= not((inputs(216)) xor (inputs(248)));
    layer0_outputs(7305) <= '0';
    layer0_outputs(7306) <= not(inputs(92));
    layer0_outputs(7307) <= (inputs(128)) or (inputs(53));
    layer0_outputs(7308) <= not((inputs(14)) and (inputs(199)));
    layer0_outputs(7309) <= not(inputs(228));
    layer0_outputs(7310) <= not(inputs(214));
    layer0_outputs(7311) <= inputs(71);
    layer0_outputs(7312) <= not((inputs(14)) or (inputs(102)));
    layer0_outputs(7313) <= not((inputs(34)) xor (inputs(19)));
    layer0_outputs(7314) <= not(inputs(91)) or (inputs(160));
    layer0_outputs(7315) <= inputs(162);
    layer0_outputs(7316) <= (inputs(182)) and not (inputs(133));
    layer0_outputs(7317) <= (inputs(79)) xor (inputs(174));
    layer0_outputs(7318) <= (inputs(39)) xor (inputs(28));
    layer0_outputs(7319) <= not(inputs(158));
    layer0_outputs(7320) <= inputs(206);
    layer0_outputs(7321) <= not(inputs(244)) or (inputs(95));
    layer0_outputs(7322) <= not((inputs(59)) or (inputs(145)));
    layer0_outputs(7323) <= not((inputs(61)) or (inputs(60)));
    layer0_outputs(7324) <= inputs(86);
    layer0_outputs(7325) <= not(inputs(70));
    layer0_outputs(7326) <= (inputs(199)) and not (inputs(46));
    layer0_outputs(7327) <= '0';
    layer0_outputs(7328) <= inputs(195);
    layer0_outputs(7329) <= (inputs(91)) or (inputs(89));
    layer0_outputs(7330) <= (inputs(66)) and not (inputs(54));
    layer0_outputs(7331) <= inputs(165);
    layer0_outputs(7332) <= not(inputs(141)) or (inputs(255));
    layer0_outputs(7333) <= not(inputs(244));
    layer0_outputs(7334) <= not(inputs(107));
    layer0_outputs(7335) <= (inputs(164)) xor (inputs(228));
    layer0_outputs(7336) <= inputs(248);
    layer0_outputs(7337) <= not(inputs(37)) or (inputs(54));
    layer0_outputs(7338) <= (inputs(172)) xor (inputs(5));
    layer0_outputs(7339) <= not(inputs(21)) or (inputs(85));
    layer0_outputs(7340) <= inputs(233);
    layer0_outputs(7341) <= not((inputs(0)) or (inputs(22)));
    layer0_outputs(7342) <= inputs(108);
    layer0_outputs(7343) <= not((inputs(245)) or (inputs(29)));
    layer0_outputs(7344) <= (inputs(153)) and not (inputs(58));
    layer0_outputs(7345) <= '0';
    layer0_outputs(7346) <= not((inputs(88)) or (inputs(152)));
    layer0_outputs(7347) <= not(inputs(12)) or (inputs(223));
    layer0_outputs(7348) <= (inputs(68)) xor (inputs(65));
    layer0_outputs(7349) <= inputs(72);
    layer0_outputs(7350) <= not(inputs(40));
    layer0_outputs(7351) <= not(inputs(188));
    layer0_outputs(7352) <= not((inputs(209)) or (inputs(149)));
    layer0_outputs(7353) <= not(inputs(5)) or (inputs(54));
    layer0_outputs(7354) <= not(inputs(179)) or (inputs(35));
    layer0_outputs(7355) <= not(inputs(162));
    layer0_outputs(7356) <= (inputs(193)) and not (inputs(112));
    layer0_outputs(7357) <= not((inputs(44)) and (inputs(39)));
    layer0_outputs(7358) <= (inputs(161)) xor (inputs(141));
    layer0_outputs(7359) <= not((inputs(8)) or (inputs(154)));
    layer0_outputs(7360) <= (inputs(14)) and not (inputs(78));
    layer0_outputs(7361) <= not((inputs(155)) xor (inputs(146)));
    layer0_outputs(7362) <= not((inputs(69)) and (inputs(5)));
    layer0_outputs(7363) <= not((inputs(17)) or (inputs(230)));
    layer0_outputs(7364) <= inputs(138);
    layer0_outputs(7365) <= (inputs(105)) or (inputs(97));
    layer0_outputs(7366) <= not((inputs(99)) and (inputs(193)));
    layer0_outputs(7367) <= not(inputs(152)) or (inputs(247));
    layer0_outputs(7368) <= (inputs(147)) and not (inputs(217));
    layer0_outputs(7369) <= (inputs(121)) and not (inputs(132));
    layer0_outputs(7370) <= not((inputs(132)) xor (inputs(98)));
    layer0_outputs(7371) <= not((inputs(214)) xor (inputs(206)));
    layer0_outputs(7372) <= not(inputs(182)) or (inputs(63));
    layer0_outputs(7373) <= not((inputs(12)) xor (inputs(17)));
    layer0_outputs(7374) <= inputs(144);
    layer0_outputs(7375) <= '1';
    layer0_outputs(7376) <= (inputs(171)) or (inputs(186));
    layer0_outputs(7377) <= not(inputs(164));
    layer0_outputs(7378) <= (inputs(236)) or (inputs(243));
    layer0_outputs(7379) <= inputs(22);
    layer0_outputs(7380) <= not((inputs(181)) or (inputs(148)));
    layer0_outputs(7381) <= not(inputs(142));
    layer0_outputs(7382) <= inputs(112);
    layer0_outputs(7383) <= not((inputs(99)) or (inputs(187)));
    layer0_outputs(7384) <= (inputs(30)) and (inputs(132));
    layer0_outputs(7385) <= inputs(179);
    layer0_outputs(7386) <= not((inputs(222)) xor (inputs(235)));
    layer0_outputs(7387) <= (inputs(76)) and (inputs(190));
    layer0_outputs(7388) <= (inputs(21)) and not (inputs(77));
    layer0_outputs(7389) <= not(inputs(152)) or (inputs(45));
    layer0_outputs(7390) <= (inputs(248)) and not (inputs(30));
    layer0_outputs(7391) <= not(inputs(121)) or (inputs(149));
    layer0_outputs(7392) <= (inputs(74)) xor (inputs(24));
    layer0_outputs(7393) <= (inputs(142)) or (inputs(249));
    layer0_outputs(7394) <= not(inputs(223));
    layer0_outputs(7395) <= not(inputs(42)) or (inputs(98));
    layer0_outputs(7396) <= '1';
    layer0_outputs(7397) <= inputs(52);
    layer0_outputs(7398) <= not((inputs(119)) xor (inputs(160)));
    layer0_outputs(7399) <= not((inputs(8)) or (inputs(66)));
    layer0_outputs(7400) <= inputs(113);
    layer0_outputs(7401) <= inputs(215);
    layer0_outputs(7402) <= (inputs(53)) and not (inputs(241));
    layer0_outputs(7403) <= not(inputs(3)) or (inputs(32));
    layer0_outputs(7404) <= not((inputs(111)) or (inputs(124)));
    layer0_outputs(7405) <= '0';
    layer0_outputs(7406) <= (inputs(230)) or (inputs(51));
    layer0_outputs(7407) <= not((inputs(115)) or (inputs(43)));
    layer0_outputs(7408) <= not(inputs(103)) or (inputs(181));
    layer0_outputs(7409) <= inputs(113);
    layer0_outputs(7410) <= not(inputs(119)) or (inputs(230));
    layer0_outputs(7411) <= inputs(54);
    layer0_outputs(7412) <= '0';
    layer0_outputs(7413) <= inputs(72);
    layer0_outputs(7414) <= inputs(21);
    layer0_outputs(7415) <= not((inputs(171)) and (inputs(255)));
    layer0_outputs(7416) <= not(inputs(115)) or (inputs(104));
    layer0_outputs(7417) <= not(inputs(228));
    layer0_outputs(7418) <= not((inputs(211)) xor (inputs(115)));
    layer0_outputs(7419) <= (inputs(99)) and not (inputs(201));
    layer0_outputs(7420) <= inputs(105);
    layer0_outputs(7421) <= not((inputs(146)) or (inputs(2)));
    layer0_outputs(7422) <= inputs(181);
    layer0_outputs(7423) <= inputs(62);
    layer0_outputs(7424) <= not(inputs(11));
    layer0_outputs(7425) <= not(inputs(24));
    layer0_outputs(7426) <= (inputs(130)) or (inputs(30));
    layer0_outputs(7427) <= not((inputs(234)) or (inputs(104)));
    layer0_outputs(7428) <= not(inputs(70)) or (inputs(240));
    layer0_outputs(7429) <= inputs(134);
    layer0_outputs(7430) <= not((inputs(208)) or (inputs(172)));
    layer0_outputs(7431) <= not(inputs(86));
    layer0_outputs(7432) <= not(inputs(249)) or (inputs(84));
    layer0_outputs(7433) <= not(inputs(253));
    layer0_outputs(7434) <= '1';
    layer0_outputs(7435) <= not(inputs(57));
    layer0_outputs(7436) <= (inputs(69)) or (inputs(181));
    layer0_outputs(7437) <= inputs(42);
    layer0_outputs(7438) <= (inputs(182)) and not (inputs(168));
    layer0_outputs(7439) <= not((inputs(105)) xor (inputs(167)));
    layer0_outputs(7440) <= not(inputs(237));
    layer0_outputs(7441) <= '1';
    layer0_outputs(7442) <= (inputs(57)) xor (inputs(252));
    layer0_outputs(7443) <= inputs(210);
    layer0_outputs(7444) <= '1';
    layer0_outputs(7445) <= not(inputs(235)) or (inputs(114));
    layer0_outputs(7446) <= not((inputs(180)) or (inputs(170)));
    layer0_outputs(7447) <= not(inputs(99));
    layer0_outputs(7448) <= (inputs(184)) or (inputs(84));
    layer0_outputs(7449) <= inputs(45);
    layer0_outputs(7450) <= (inputs(207)) or (inputs(20));
    layer0_outputs(7451) <= inputs(247);
    layer0_outputs(7452) <= inputs(171);
    layer0_outputs(7453) <= (inputs(180)) xor (inputs(182));
    layer0_outputs(7454) <= not(inputs(121));
    layer0_outputs(7455) <= '1';
    layer0_outputs(7456) <= not(inputs(247)) or (inputs(57));
    layer0_outputs(7457) <= (inputs(124)) and (inputs(92));
    layer0_outputs(7458) <= not(inputs(200)) or (inputs(26));
    layer0_outputs(7459) <= (inputs(73)) xor (inputs(45));
    layer0_outputs(7460) <= not(inputs(79)) or (inputs(202));
    layer0_outputs(7461) <= not((inputs(172)) or (inputs(217)));
    layer0_outputs(7462) <= not(inputs(152));
    layer0_outputs(7463) <= (inputs(227)) or (inputs(96));
    layer0_outputs(7464) <= not((inputs(58)) or (inputs(153)));
    layer0_outputs(7465) <= (inputs(91)) and not (inputs(195));
    layer0_outputs(7466) <= not(inputs(234)) or (inputs(112));
    layer0_outputs(7467) <= not((inputs(206)) or (inputs(251)));
    layer0_outputs(7468) <= not(inputs(122));
    layer0_outputs(7469) <= inputs(58);
    layer0_outputs(7470) <= (inputs(208)) and not (inputs(113));
    layer0_outputs(7471) <= inputs(174);
    layer0_outputs(7472) <= inputs(199);
    layer0_outputs(7473) <= '0';
    layer0_outputs(7474) <= (inputs(191)) xor (inputs(172));
    layer0_outputs(7475) <= not(inputs(195));
    layer0_outputs(7476) <= (inputs(152)) and not (inputs(234));
    layer0_outputs(7477) <= not((inputs(227)) or (inputs(19)));
    layer0_outputs(7478) <= not((inputs(72)) or (inputs(143)));
    layer0_outputs(7479) <= (inputs(124)) or (inputs(37));
    layer0_outputs(7480) <= (inputs(174)) xor (inputs(126));
    layer0_outputs(7481) <= not(inputs(35));
    layer0_outputs(7482) <= not(inputs(112)) or (inputs(232));
    layer0_outputs(7483) <= (inputs(125)) or (inputs(156));
    layer0_outputs(7484) <= not(inputs(189));
    layer0_outputs(7485) <= not(inputs(197));
    layer0_outputs(7486) <= not(inputs(27));
    layer0_outputs(7487) <= (inputs(60)) and not (inputs(236));
    layer0_outputs(7488) <= (inputs(190)) or (inputs(141));
    layer0_outputs(7489) <= not((inputs(209)) xor (inputs(173)));
    layer0_outputs(7490) <= (inputs(88)) and not (inputs(3));
    layer0_outputs(7491) <= not((inputs(225)) or (inputs(15)));
    layer0_outputs(7492) <= (inputs(11)) and not (inputs(239));
    layer0_outputs(7493) <= inputs(169);
    layer0_outputs(7494) <= (inputs(229)) xor (inputs(171));
    layer0_outputs(7495) <= '0';
    layer0_outputs(7496) <= not((inputs(17)) or (inputs(196)));
    layer0_outputs(7497) <= not(inputs(127));
    layer0_outputs(7498) <= not(inputs(126));
    layer0_outputs(7499) <= not(inputs(246));
    layer0_outputs(7500) <= (inputs(189)) or (inputs(205));
    layer0_outputs(7501) <= (inputs(193)) and not (inputs(169));
    layer0_outputs(7502) <= not(inputs(74));
    layer0_outputs(7503) <= (inputs(230)) and not (inputs(152));
    layer0_outputs(7504) <= not((inputs(80)) xor (inputs(70)));
    layer0_outputs(7505) <= not(inputs(245));
    layer0_outputs(7506) <= (inputs(171)) and (inputs(214));
    layer0_outputs(7507) <= not((inputs(95)) xor (inputs(104)));
    layer0_outputs(7508) <= inputs(92);
    layer0_outputs(7509) <= (inputs(126)) or (inputs(13));
    layer0_outputs(7510) <= not(inputs(136)) or (inputs(64));
    layer0_outputs(7511) <= '0';
    layer0_outputs(7512) <= (inputs(133)) and not (inputs(190));
    layer0_outputs(7513) <= not((inputs(51)) xor (inputs(199)));
    layer0_outputs(7514) <= (inputs(83)) or (inputs(112));
    layer0_outputs(7515) <= (inputs(126)) or (inputs(181));
    layer0_outputs(7516) <= inputs(37);
    layer0_outputs(7517) <= not(inputs(95));
    layer0_outputs(7518) <= inputs(217);
    layer0_outputs(7519) <= not((inputs(74)) or (inputs(129)));
    layer0_outputs(7520) <= not((inputs(57)) and (inputs(53)));
    layer0_outputs(7521) <= inputs(81);
    layer0_outputs(7522) <= not(inputs(183)) or (inputs(207));
    layer0_outputs(7523) <= not(inputs(38)) or (inputs(201));
    layer0_outputs(7524) <= (inputs(100)) and not (inputs(80));
    layer0_outputs(7525) <= (inputs(49)) and not (inputs(209));
    layer0_outputs(7526) <= (inputs(178)) and not (inputs(31));
    layer0_outputs(7527) <= not(inputs(138));
    layer0_outputs(7528) <= (inputs(195)) xor (inputs(0));
    layer0_outputs(7529) <= (inputs(255)) or (inputs(49));
    layer0_outputs(7530) <= not(inputs(238));
    layer0_outputs(7531) <= not((inputs(86)) xor (inputs(19)));
    layer0_outputs(7532) <= not((inputs(26)) or (inputs(92)));
    layer0_outputs(7533) <= not(inputs(89)) or (inputs(248));
    layer0_outputs(7534) <= (inputs(188)) xor (inputs(179));
    layer0_outputs(7535) <= not((inputs(192)) or (inputs(95)));
    layer0_outputs(7536) <= '0';
    layer0_outputs(7537) <= not((inputs(50)) or (inputs(79)));
    layer0_outputs(7538) <= (inputs(88)) and (inputs(61));
    layer0_outputs(7539) <= inputs(242);
    layer0_outputs(7540) <= (inputs(141)) or (inputs(97));
    layer0_outputs(7541) <= inputs(218);
    layer0_outputs(7542) <= inputs(85);
    layer0_outputs(7543) <= not((inputs(114)) or (inputs(102)));
    layer0_outputs(7544) <= not(inputs(191));
    layer0_outputs(7545) <= not((inputs(192)) and (inputs(132)));
    layer0_outputs(7546) <= (inputs(187)) and not (inputs(14));
    layer0_outputs(7547) <= '1';
    layer0_outputs(7548) <= (inputs(112)) and not (inputs(238));
    layer0_outputs(7549) <= not(inputs(73));
    layer0_outputs(7550) <= not((inputs(149)) xor (inputs(221)));
    layer0_outputs(7551) <= (inputs(139)) or (inputs(106));
    layer0_outputs(7552) <= (inputs(75)) and not (inputs(81));
    layer0_outputs(7553) <= inputs(201);
    layer0_outputs(7554) <= not(inputs(87)) or (inputs(13));
    layer0_outputs(7555) <= (inputs(17)) and not (inputs(3));
    layer0_outputs(7556) <= (inputs(158)) xor (inputs(39));
    layer0_outputs(7557) <= (inputs(207)) xor (inputs(255));
    layer0_outputs(7558) <= not(inputs(9));
    layer0_outputs(7559) <= not(inputs(107)) or (inputs(40));
    layer0_outputs(7560) <= (inputs(186)) and not (inputs(102));
    layer0_outputs(7561) <= not((inputs(214)) or (inputs(183)));
    layer0_outputs(7562) <= not(inputs(3));
    layer0_outputs(7563) <= (inputs(129)) or (inputs(156));
    layer0_outputs(7564) <= (inputs(161)) or (inputs(175));
    layer0_outputs(7565) <= not((inputs(129)) or (inputs(149)));
    layer0_outputs(7566) <= not(inputs(76));
    layer0_outputs(7567) <= '0';
    layer0_outputs(7568) <= (inputs(251)) and (inputs(139));
    layer0_outputs(7569) <= not(inputs(34));
    layer0_outputs(7570) <= (inputs(183)) xor (inputs(230));
    layer0_outputs(7571) <= inputs(213);
    layer0_outputs(7572) <= '0';
    layer0_outputs(7573) <= (inputs(19)) xor (inputs(3));
    layer0_outputs(7574) <= not((inputs(31)) or (inputs(122)));
    layer0_outputs(7575) <= not((inputs(66)) xor (inputs(91)));
    layer0_outputs(7576) <= not(inputs(82)) or (inputs(240));
    layer0_outputs(7577) <= (inputs(202)) xor (inputs(111));
    layer0_outputs(7578) <= not(inputs(138));
    layer0_outputs(7579) <= (inputs(120)) and not (inputs(155));
    layer0_outputs(7580) <= (inputs(99)) or (inputs(46));
    layer0_outputs(7581) <= not((inputs(252)) xor (inputs(129)));
    layer0_outputs(7582) <= (inputs(253)) or (inputs(61));
    layer0_outputs(7583) <= inputs(38);
    layer0_outputs(7584) <= (inputs(179)) or (inputs(111));
    layer0_outputs(7585) <= not(inputs(71)) or (inputs(224));
    layer0_outputs(7586) <= inputs(177);
    layer0_outputs(7587) <= not(inputs(51));
    layer0_outputs(7588) <= not((inputs(44)) or (inputs(84)));
    layer0_outputs(7589) <= inputs(228);
    layer0_outputs(7590) <= not((inputs(138)) xor (inputs(74)));
    layer0_outputs(7591) <= (inputs(89)) xor (inputs(112));
    layer0_outputs(7592) <= (inputs(32)) xor (inputs(128));
    layer0_outputs(7593) <= not(inputs(127));
    layer0_outputs(7594) <= (inputs(158)) and not (inputs(126));
    layer0_outputs(7595) <= not((inputs(167)) or (inputs(111)));
    layer0_outputs(7596) <= not((inputs(166)) or (inputs(33)));
    layer0_outputs(7597) <= not(inputs(132)) or (inputs(190));
    layer0_outputs(7598) <= not(inputs(146));
    layer0_outputs(7599) <= not((inputs(214)) or (inputs(19)));
    layer0_outputs(7600) <= not((inputs(128)) or (inputs(58)));
    layer0_outputs(7601) <= (inputs(226)) xor (inputs(232));
    layer0_outputs(7602) <= (inputs(233)) or (inputs(26));
    layer0_outputs(7603) <= (inputs(203)) and not (inputs(42));
    layer0_outputs(7604) <= (inputs(107)) and not (inputs(153));
    layer0_outputs(7605) <= (inputs(197)) or (inputs(76));
    layer0_outputs(7606) <= not(inputs(101)) or (inputs(160));
    layer0_outputs(7607) <= (inputs(134)) and not (inputs(7));
    layer0_outputs(7608) <= not(inputs(105));
    layer0_outputs(7609) <= (inputs(235)) xor (inputs(250));
    layer0_outputs(7610) <= not(inputs(90)) or (inputs(188));
    layer0_outputs(7611) <= not(inputs(156)) or (inputs(65));
    layer0_outputs(7612) <= not((inputs(83)) xor (inputs(82)));
    layer0_outputs(7613) <= not(inputs(29)) or (inputs(50));
    layer0_outputs(7614) <= inputs(34);
    layer0_outputs(7615) <= not(inputs(8));
    layer0_outputs(7616) <= (inputs(158)) and (inputs(218));
    layer0_outputs(7617) <= not(inputs(107));
    layer0_outputs(7618) <= (inputs(107)) or (inputs(74));
    layer0_outputs(7619) <= '1';
    layer0_outputs(7620) <= not(inputs(70));
    layer0_outputs(7621) <= not(inputs(178));
    layer0_outputs(7622) <= (inputs(43)) or (inputs(218));
    layer0_outputs(7623) <= not((inputs(242)) and (inputs(235)));
    layer0_outputs(7624) <= inputs(202);
    layer0_outputs(7625) <= not((inputs(65)) xor (inputs(104)));
    layer0_outputs(7626) <= not(inputs(19)) or (inputs(178));
    layer0_outputs(7627) <= inputs(202);
    layer0_outputs(7628) <= '0';
    layer0_outputs(7629) <= (inputs(240)) and not (inputs(177));
    layer0_outputs(7630) <= inputs(85);
    layer0_outputs(7631) <= not((inputs(118)) or (inputs(164)));
    layer0_outputs(7632) <= not(inputs(74)) or (inputs(167));
    layer0_outputs(7633) <= not(inputs(68));
    layer0_outputs(7634) <= not((inputs(156)) xor (inputs(122)));
    layer0_outputs(7635) <= not(inputs(60));
    layer0_outputs(7636) <= (inputs(236)) or (inputs(161));
    layer0_outputs(7637) <= (inputs(172)) or (inputs(217));
    layer0_outputs(7638) <= not(inputs(121));
    layer0_outputs(7639) <= (inputs(12)) and not (inputs(61));
    layer0_outputs(7640) <= '1';
    layer0_outputs(7641) <= not((inputs(43)) or (inputs(106)));
    layer0_outputs(7642) <= '1';
    layer0_outputs(7643) <= not(inputs(134));
    layer0_outputs(7644) <= (inputs(224)) or (inputs(89));
    layer0_outputs(7645) <= (inputs(21)) and not (inputs(68));
    layer0_outputs(7646) <= (inputs(124)) xor (inputs(35));
    layer0_outputs(7647) <= not((inputs(8)) xor (inputs(0)));
    layer0_outputs(7648) <= not((inputs(124)) or (inputs(101)));
    layer0_outputs(7649) <= (inputs(9)) and (inputs(75));
    layer0_outputs(7650) <= not(inputs(68)) or (inputs(231));
    layer0_outputs(7651) <= (inputs(82)) and not (inputs(233));
    layer0_outputs(7652) <= not((inputs(254)) or (inputs(190)));
    layer0_outputs(7653) <= inputs(85);
    layer0_outputs(7654) <= not(inputs(68));
    layer0_outputs(7655) <= (inputs(133)) and not (inputs(188));
    layer0_outputs(7656) <= '0';
    layer0_outputs(7657) <= not((inputs(141)) or (inputs(147)));
    layer0_outputs(7658) <= (inputs(180)) or (inputs(224));
    layer0_outputs(7659) <= inputs(63);
    layer0_outputs(7660) <= not((inputs(1)) xor (inputs(224)));
    layer0_outputs(7661) <= not((inputs(247)) or (inputs(87)));
    layer0_outputs(7662) <= not((inputs(77)) xor (inputs(28)));
    layer0_outputs(7663) <= (inputs(57)) xor (inputs(0));
    layer0_outputs(7664) <= (inputs(153)) and (inputs(135));
    layer0_outputs(7665) <= not(inputs(142));
    layer0_outputs(7666) <= not(inputs(250));
    layer0_outputs(7667) <= not(inputs(177));
    layer0_outputs(7668) <= not(inputs(120)) or (inputs(28));
    layer0_outputs(7669) <= '0';
    layer0_outputs(7670) <= (inputs(118)) and not (inputs(178));
    layer0_outputs(7671) <= (inputs(253)) or (inputs(225));
    layer0_outputs(7672) <= not((inputs(180)) xor (inputs(15)));
    layer0_outputs(7673) <= inputs(10);
    layer0_outputs(7674) <= (inputs(126)) and not (inputs(147));
    layer0_outputs(7675) <= inputs(152);
    layer0_outputs(7676) <= not(inputs(96));
    layer0_outputs(7677) <= (inputs(60)) or (inputs(129));
    layer0_outputs(7678) <= not((inputs(138)) xor (inputs(109)));
    layer0_outputs(7679) <= inputs(120);
    layer0_outputs(7680) <= not(inputs(220));
    layer0_outputs(7681) <= not((inputs(171)) and (inputs(164)));
    layer0_outputs(7682) <= (inputs(174)) or (inputs(160));
    layer0_outputs(7683) <= not(inputs(52)) or (inputs(33));
    layer0_outputs(7684) <= (inputs(36)) and not (inputs(1));
    layer0_outputs(7685) <= inputs(138);
    layer0_outputs(7686) <= inputs(23);
    layer0_outputs(7687) <= not(inputs(205)) or (inputs(250));
    layer0_outputs(7688) <= (inputs(137)) and (inputs(97));
    layer0_outputs(7689) <= (inputs(231)) and (inputs(27));
    layer0_outputs(7690) <= not(inputs(106)) or (inputs(58));
    layer0_outputs(7691) <= inputs(228);
    layer0_outputs(7692) <= not(inputs(38));
    layer0_outputs(7693) <= inputs(237);
    layer0_outputs(7694) <= (inputs(117)) or (inputs(86));
    layer0_outputs(7695) <= (inputs(245)) and not (inputs(34));
    layer0_outputs(7696) <= (inputs(48)) and not (inputs(49));
    layer0_outputs(7697) <= inputs(230);
    layer0_outputs(7698) <= not(inputs(93));
    layer0_outputs(7699) <= (inputs(146)) and not (inputs(3));
    layer0_outputs(7700) <= not(inputs(90));
    layer0_outputs(7701) <= (inputs(138)) and not (inputs(103));
    layer0_outputs(7702) <= (inputs(6)) and not (inputs(143));
    layer0_outputs(7703) <= (inputs(219)) or (inputs(226));
    layer0_outputs(7704) <= not((inputs(62)) and (inputs(62)));
    layer0_outputs(7705) <= (inputs(196)) or (inputs(253));
    layer0_outputs(7706) <= (inputs(191)) or (inputs(166));
    layer0_outputs(7707) <= not(inputs(155));
    layer0_outputs(7708) <= inputs(154);
    layer0_outputs(7709) <= not(inputs(24));
    layer0_outputs(7710) <= not(inputs(88)) or (inputs(38));
    layer0_outputs(7711) <= not(inputs(48));
    layer0_outputs(7712) <= not((inputs(52)) xor (inputs(176)));
    layer0_outputs(7713) <= (inputs(235)) or (inputs(223));
    layer0_outputs(7714) <= not((inputs(113)) xor (inputs(57)));
    layer0_outputs(7715) <= inputs(162);
    layer0_outputs(7716) <= not(inputs(112));
    layer0_outputs(7717) <= not(inputs(126));
    layer0_outputs(7718) <= inputs(169);
    layer0_outputs(7719) <= not(inputs(231));
    layer0_outputs(7720) <= '0';
    layer0_outputs(7721) <= not(inputs(64));
    layer0_outputs(7722) <= not(inputs(251));
    layer0_outputs(7723) <= not(inputs(127));
    layer0_outputs(7724) <= inputs(94);
    layer0_outputs(7725) <= (inputs(103)) xor (inputs(147));
    layer0_outputs(7726) <= not((inputs(16)) or (inputs(60)));
    layer0_outputs(7727) <= (inputs(16)) and not (inputs(155));
    layer0_outputs(7728) <= not(inputs(135)) or (inputs(160));
    layer0_outputs(7729) <= inputs(110);
    layer0_outputs(7730) <= (inputs(61)) or (inputs(84));
    layer0_outputs(7731) <= (inputs(23)) xor (inputs(232));
    layer0_outputs(7732) <= not(inputs(168));
    layer0_outputs(7733) <= not(inputs(78));
    layer0_outputs(7734) <= inputs(164);
    layer0_outputs(7735) <= not((inputs(81)) or (inputs(188)));
    layer0_outputs(7736) <= not(inputs(21));
    layer0_outputs(7737) <= not((inputs(183)) and (inputs(32)));
    layer0_outputs(7738) <= (inputs(97)) or (inputs(228));
    layer0_outputs(7739) <= not((inputs(196)) or (inputs(65)));
    layer0_outputs(7740) <= not(inputs(152));
    layer0_outputs(7741) <= not((inputs(74)) or (inputs(67)));
    layer0_outputs(7742) <= not(inputs(34));
    layer0_outputs(7743) <= (inputs(225)) or (inputs(78));
    layer0_outputs(7744) <= not((inputs(241)) or (inputs(222)));
    layer0_outputs(7745) <= not(inputs(185));
    layer0_outputs(7746) <= not((inputs(8)) or (inputs(121)));
    layer0_outputs(7747) <= not(inputs(136));
    layer0_outputs(7748) <= inputs(107);
    layer0_outputs(7749) <= (inputs(180)) or (inputs(228));
    layer0_outputs(7750) <= (inputs(150)) xor (inputs(153));
    layer0_outputs(7751) <= (inputs(29)) and (inputs(21));
    layer0_outputs(7752) <= (inputs(175)) and not (inputs(57));
    layer0_outputs(7753) <= (inputs(186)) and not (inputs(123));
    layer0_outputs(7754) <= '0';
    layer0_outputs(7755) <= (inputs(183)) and not (inputs(10));
    layer0_outputs(7756) <= '0';
    layer0_outputs(7757) <= '0';
    layer0_outputs(7758) <= not(inputs(144)) or (inputs(246));
    layer0_outputs(7759) <= '0';
    layer0_outputs(7760) <= not(inputs(1));
    layer0_outputs(7761) <= inputs(62);
    layer0_outputs(7762) <= inputs(36);
    layer0_outputs(7763) <= not(inputs(213));
    layer0_outputs(7764) <= (inputs(127)) or (inputs(38));
    layer0_outputs(7765) <= not(inputs(203)) or (inputs(109));
    layer0_outputs(7766) <= not(inputs(245)) or (inputs(77));
    layer0_outputs(7767) <= inputs(139);
    layer0_outputs(7768) <= (inputs(194)) and not (inputs(126));
    layer0_outputs(7769) <= (inputs(176)) and not (inputs(82));
    layer0_outputs(7770) <= not((inputs(125)) xor (inputs(127)));
    layer0_outputs(7771) <= not(inputs(49));
    layer0_outputs(7772) <= not(inputs(140)) or (inputs(69));
    layer0_outputs(7773) <= not(inputs(225));
    layer0_outputs(7774) <= (inputs(181)) and not (inputs(99));
    layer0_outputs(7775) <= inputs(146);
    layer0_outputs(7776) <= not(inputs(181));
    layer0_outputs(7777) <= inputs(156);
    layer0_outputs(7778) <= not(inputs(46)) or (inputs(236));
    layer0_outputs(7779) <= inputs(43);
    layer0_outputs(7780) <= not((inputs(180)) or (inputs(2)));
    layer0_outputs(7781) <= not(inputs(99)) or (inputs(11));
    layer0_outputs(7782) <= not((inputs(65)) or (inputs(51)));
    layer0_outputs(7783) <= not(inputs(150));
    layer0_outputs(7784) <= (inputs(32)) and not (inputs(220));
    layer0_outputs(7785) <= (inputs(216)) or (inputs(215));
    layer0_outputs(7786) <= not(inputs(53));
    layer0_outputs(7787) <= '1';
    layer0_outputs(7788) <= not(inputs(22)) or (inputs(174));
    layer0_outputs(7789) <= (inputs(250)) xor (inputs(209));
    layer0_outputs(7790) <= inputs(144);
    layer0_outputs(7791) <= (inputs(230)) or (inputs(219));
    layer0_outputs(7792) <= not((inputs(163)) and (inputs(112)));
    layer0_outputs(7793) <= not(inputs(231));
    layer0_outputs(7794) <= (inputs(91)) and not (inputs(190));
    layer0_outputs(7795) <= (inputs(20)) or (inputs(148));
    layer0_outputs(7796) <= (inputs(145)) or (inputs(185));
    layer0_outputs(7797) <= not((inputs(76)) or (inputs(23)));
    layer0_outputs(7798) <= inputs(154);
    layer0_outputs(7799) <= not((inputs(30)) and (inputs(108)));
    layer0_outputs(7800) <= (inputs(187)) or (inputs(108));
    layer0_outputs(7801) <= not((inputs(9)) or (inputs(62)));
    layer0_outputs(7802) <= not(inputs(116)) or (inputs(169));
    layer0_outputs(7803) <= (inputs(220)) or (inputs(239));
    layer0_outputs(7804) <= not((inputs(46)) and (inputs(236)));
    layer0_outputs(7805) <= inputs(101);
    layer0_outputs(7806) <= not(inputs(198));
    layer0_outputs(7807) <= '0';
    layer0_outputs(7808) <= (inputs(78)) and not (inputs(19));
    layer0_outputs(7809) <= not(inputs(146));
    layer0_outputs(7810) <= (inputs(23)) and not (inputs(118));
    layer0_outputs(7811) <= not((inputs(192)) and (inputs(69)));
    layer0_outputs(7812) <= not(inputs(91));
    layer0_outputs(7813) <= inputs(255);
    layer0_outputs(7814) <= inputs(7);
    layer0_outputs(7815) <= not((inputs(165)) or (inputs(143)));
    layer0_outputs(7816) <= '1';
    layer0_outputs(7817) <= inputs(93);
    layer0_outputs(7818) <= not((inputs(221)) xor (inputs(253)));
    layer0_outputs(7819) <= inputs(58);
    layer0_outputs(7820) <= (inputs(150)) and not (inputs(220));
    layer0_outputs(7821) <= not(inputs(41)) or (inputs(77));
    layer0_outputs(7822) <= '1';
    layer0_outputs(7823) <= not(inputs(87)) or (inputs(214));
    layer0_outputs(7824) <= (inputs(140)) and (inputs(222));
    layer0_outputs(7825) <= inputs(5);
    layer0_outputs(7826) <= not((inputs(37)) xor (inputs(254)));
    layer0_outputs(7827) <= not((inputs(49)) or (inputs(195)));
    layer0_outputs(7828) <= not((inputs(14)) or (inputs(54)));
    layer0_outputs(7829) <= inputs(40);
    layer0_outputs(7830) <= inputs(120);
    layer0_outputs(7831) <= not(inputs(218)) or (inputs(133));
    layer0_outputs(7832) <= (inputs(53)) or (inputs(161));
    layer0_outputs(7833) <= not(inputs(132));
    layer0_outputs(7834) <= '1';
    layer0_outputs(7835) <= (inputs(69)) xor (inputs(164));
    layer0_outputs(7836) <= not(inputs(142)) or (inputs(126));
    layer0_outputs(7837) <= (inputs(67)) and not (inputs(161));
    layer0_outputs(7838) <= not(inputs(4)) or (inputs(90));
    layer0_outputs(7839) <= (inputs(95)) and not (inputs(51));
    layer0_outputs(7840) <= (inputs(164)) and (inputs(35));
    layer0_outputs(7841) <= not(inputs(133)) or (inputs(254));
    layer0_outputs(7842) <= not((inputs(43)) or (inputs(196)));
    layer0_outputs(7843) <= not(inputs(42));
    layer0_outputs(7844) <= not(inputs(99)) or (inputs(174));
    layer0_outputs(7845) <= (inputs(99)) or (inputs(23));
    layer0_outputs(7846) <= (inputs(85)) or (inputs(147));
    layer0_outputs(7847) <= not((inputs(83)) and (inputs(80)));
    layer0_outputs(7848) <= '0';
    layer0_outputs(7849) <= (inputs(89)) or (inputs(65));
    layer0_outputs(7850) <= not(inputs(179));
    layer0_outputs(7851) <= inputs(202);
    layer0_outputs(7852) <= (inputs(135)) or (inputs(107));
    layer0_outputs(7853) <= '1';
    layer0_outputs(7854) <= not((inputs(253)) or (inputs(185)));
    layer0_outputs(7855) <= not(inputs(43));
    layer0_outputs(7856) <= not(inputs(78)) or (inputs(26));
    layer0_outputs(7857) <= (inputs(106)) or (inputs(187));
    layer0_outputs(7858) <= not((inputs(250)) or (inputs(145)));
    layer0_outputs(7859) <= not(inputs(111));
    layer0_outputs(7860) <= (inputs(222)) or (inputs(111));
    layer0_outputs(7861) <= not(inputs(130));
    layer0_outputs(7862) <= (inputs(218)) and not (inputs(109));
    layer0_outputs(7863) <= inputs(91);
    layer0_outputs(7864) <= not(inputs(133));
    layer0_outputs(7865) <= not(inputs(84));
    layer0_outputs(7866) <= not((inputs(54)) or (inputs(226)));
    layer0_outputs(7867) <= (inputs(116)) or (inputs(112));
    layer0_outputs(7868) <= inputs(119);
    layer0_outputs(7869) <= not(inputs(2));
    layer0_outputs(7870) <= not((inputs(232)) xor (inputs(242)));
    layer0_outputs(7871) <= not(inputs(184));
    layer0_outputs(7872) <= not(inputs(233)) or (inputs(211));
    layer0_outputs(7873) <= not(inputs(249)) or (inputs(18));
    layer0_outputs(7874) <= not((inputs(125)) or (inputs(94)));
    layer0_outputs(7875) <= inputs(106);
    layer0_outputs(7876) <= inputs(200);
    layer0_outputs(7877) <= inputs(133);
    layer0_outputs(7878) <= (inputs(78)) or (inputs(79));
    layer0_outputs(7879) <= inputs(48);
    layer0_outputs(7880) <= not(inputs(8));
    layer0_outputs(7881) <= inputs(223);
    layer0_outputs(7882) <= not((inputs(222)) and (inputs(7)));
    layer0_outputs(7883) <= not(inputs(154));
    layer0_outputs(7884) <= (inputs(90)) and not (inputs(219));
    layer0_outputs(7885) <= inputs(107);
    layer0_outputs(7886) <= (inputs(75)) and not (inputs(235));
    layer0_outputs(7887) <= not(inputs(115));
    layer0_outputs(7888) <= (inputs(81)) xor (inputs(42));
    layer0_outputs(7889) <= (inputs(198)) xor (inputs(75));
    layer0_outputs(7890) <= not(inputs(166)) or (inputs(222));
    layer0_outputs(7891) <= not(inputs(103));
    layer0_outputs(7892) <= not((inputs(71)) xor (inputs(74)));
    layer0_outputs(7893) <= (inputs(200)) xor (inputs(201));
    layer0_outputs(7894) <= not(inputs(159)) or (inputs(151));
    layer0_outputs(7895) <= (inputs(228)) and not (inputs(132));
    layer0_outputs(7896) <= inputs(0);
    layer0_outputs(7897) <= (inputs(92)) and not (inputs(12));
    layer0_outputs(7898) <= inputs(161);
    layer0_outputs(7899) <= inputs(180);
    layer0_outputs(7900) <= (inputs(118)) xor (inputs(103));
    layer0_outputs(7901) <= inputs(168);
    layer0_outputs(7902) <= (inputs(134)) and not (inputs(105));
    layer0_outputs(7903) <= not(inputs(103));
    layer0_outputs(7904) <= inputs(100);
    layer0_outputs(7905) <= not(inputs(103)) or (inputs(1));
    layer0_outputs(7906) <= '1';
    layer0_outputs(7907) <= (inputs(193)) or (inputs(5));
    layer0_outputs(7908) <= not(inputs(194)) or (inputs(5));
    layer0_outputs(7909) <= inputs(196);
    layer0_outputs(7910) <= not(inputs(93));
    layer0_outputs(7911) <= not((inputs(152)) or (inputs(182)));
    layer0_outputs(7912) <= not((inputs(44)) xor (inputs(74)));
    layer0_outputs(7913) <= not((inputs(148)) or (inputs(148)));
    layer0_outputs(7914) <= '1';
    layer0_outputs(7915) <= inputs(141);
    layer0_outputs(7916) <= not(inputs(8));
    layer0_outputs(7917) <= inputs(24);
    layer0_outputs(7918) <= (inputs(177)) xor (inputs(234));
    layer0_outputs(7919) <= not((inputs(246)) or (inputs(207)));
    layer0_outputs(7920) <= (inputs(221)) xor (inputs(189));
    layer0_outputs(7921) <= (inputs(234)) or (inputs(207));
    layer0_outputs(7922) <= not(inputs(122));
    layer0_outputs(7923) <= (inputs(123)) xor (inputs(170));
    layer0_outputs(7924) <= not((inputs(204)) and (inputs(139)));
    layer0_outputs(7925) <= (inputs(243)) xor (inputs(210));
    layer0_outputs(7926) <= '1';
    layer0_outputs(7927) <= not((inputs(86)) xor (inputs(80)));
    layer0_outputs(7928) <= inputs(70);
    layer0_outputs(7929) <= not((inputs(155)) xor (inputs(51)));
    layer0_outputs(7930) <= not(inputs(57)) or (inputs(20));
    layer0_outputs(7931) <= inputs(44);
    layer0_outputs(7932) <= not((inputs(33)) or (inputs(236)));
    layer0_outputs(7933) <= inputs(143);
    layer0_outputs(7934) <= (inputs(151)) and not (inputs(73));
    layer0_outputs(7935) <= not(inputs(56));
    layer0_outputs(7936) <= not(inputs(194));
    layer0_outputs(7937) <= not(inputs(118));
    layer0_outputs(7938) <= not((inputs(168)) and (inputs(77)));
    layer0_outputs(7939) <= (inputs(229)) and not (inputs(104));
    layer0_outputs(7940) <= inputs(104);
    layer0_outputs(7941) <= (inputs(212)) or (inputs(6));
    layer0_outputs(7942) <= not((inputs(91)) and (inputs(163)));
    layer0_outputs(7943) <= not((inputs(0)) and (inputs(40)));
    layer0_outputs(7944) <= inputs(36);
    layer0_outputs(7945) <= not((inputs(51)) and (inputs(169)));
    layer0_outputs(7946) <= not((inputs(4)) xor (inputs(11)));
    layer0_outputs(7947) <= not((inputs(141)) or (inputs(132)));
    layer0_outputs(7948) <= (inputs(219)) and not (inputs(142));
    layer0_outputs(7949) <= (inputs(62)) xor (inputs(218));
    layer0_outputs(7950) <= not((inputs(220)) or (inputs(109)));
    layer0_outputs(7951) <= inputs(148);
    layer0_outputs(7952) <= not(inputs(223)) or (inputs(96));
    layer0_outputs(7953) <= not(inputs(187));
    layer0_outputs(7954) <= (inputs(101)) and not (inputs(115));
    layer0_outputs(7955) <= (inputs(216)) or (inputs(9));
    layer0_outputs(7956) <= (inputs(166)) xor (inputs(108));
    layer0_outputs(7957) <= inputs(108);
    layer0_outputs(7958) <= (inputs(62)) xor (inputs(247));
    layer0_outputs(7959) <= (inputs(212)) and not (inputs(111));
    layer0_outputs(7960) <= (inputs(223)) and (inputs(128));
    layer0_outputs(7961) <= not(inputs(59));
    layer0_outputs(7962) <= not(inputs(165)) or (inputs(47));
    layer0_outputs(7963) <= (inputs(210)) and not (inputs(27));
    layer0_outputs(7964) <= not(inputs(41));
    layer0_outputs(7965) <= (inputs(143)) and not (inputs(248));
    layer0_outputs(7966) <= inputs(169);
    layer0_outputs(7967) <= (inputs(89)) and not (inputs(224));
    layer0_outputs(7968) <= inputs(136);
    layer0_outputs(7969) <= (inputs(212)) or (inputs(212));
    layer0_outputs(7970) <= not(inputs(133)) or (inputs(137));
    layer0_outputs(7971) <= '1';
    layer0_outputs(7972) <= inputs(46);
    layer0_outputs(7973) <= not(inputs(65)) or (inputs(145));
    layer0_outputs(7974) <= inputs(2);
    layer0_outputs(7975) <= inputs(20);
    layer0_outputs(7976) <= '1';
    layer0_outputs(7977) <= (inputs(217)) and not (inputs(123));
    layer0_outputs(7978) <= not(inputs(214));
    layer0_outputs(7979) <= inputs(98);
    layer0_outputs(7980) <= not(inputs(110));
    layer0_outputs(7981) <= not(inputs(87)) or (inputs(73));
    layer0_outputs(7982) <= (inputs(93)) or (inputs(93));
    layer0_outputs(7983) <= inputs(111);
    layer0_outputs(7984) <= (inputs(97)) or (inputs(99));
    layer0_outputs(7985) <= '0';
    layer0_outputs(7986) <= (inputs(209)) xor (inputs(251));
    layer0_outputs(7987) <= (inputs(153)) xor (inputs(42));
    layer0_outputs(7988) <= not((inputs(55)) xor (inputs(6)));
    layer0_outputs(7989) <= (inputs(65)) xor (inputs(35));
    layer0_outputs(7990) <= not((inputs(156)) or (inputs(163)));
    layer0_outputs(7991) <= not((inputs(208)) xor (inputs(38)));
    layer0_outputs(7992) <= not(inputs(80)) or (inputs(198));
    layer0_outputs(7993) <= (inputs(190)) xor (inputs(180));
    layer0_outputs(7994) <= not((inputs(63)) xor (inputs(204)));
    layer0_outputs(7995) <= not(inputs(99));
    layer0_outputs(7996) <= not(inputs(233));
    layer0_outputs(7997) <= not(inputs(247)) or (inputs(163));
    layer0_outputs(7998) <= not(inputs(3)) or (inputs(206));
    layer0_outputs(7999) <= inputs(36);
    layer0_outputs(8000) <= (inputs(203)) xor (inputs(135));
    layer0_outputs(8001) <= not(inputs(92)) or (inputs(235));
    layer0_outputs(8002) <= (inputs(32)) xor (inputs(63));
    layer0_outputs(8003) <= not((inputs(112)) or (inputs(160)));
    layer0_outputs(8004) <= not((inputs(238)) or (inputs(191)));
    layer0_outputs(8005) <= (inputs(213)) and not (inputs(49));
    layer0_outputs(8006) <= inputs(85);
    layer0_outputs(8007) <= (inputs(92)) and not (inputs(83));
    layer0_outputs(8008) <= not((inputs(201)) or (inputs(151)));
    layer0_outputs(8009) <= not((inputs(195)) or (inputs(233)));
    layer0_outputs(8010) <= inputs(41);
    layer0_outputs(8011) <= (inputs(23)) and not (inputs(188));
    layer0_outputs(8012) <= (inputs(93)) xor (inputs(160));
    layer0_outputs(8013) <= inputs(92);
    layer0_outputs(8014) <= (inputs(46)) and not (inputs(8));
    layer0_outputs(8015) <= (inputs(65)) or (inputs(116));
    layer0_outputs(8016) <= (inputs(31)) xor (inputs(39));
    layer0_outputs(8017) <= (inputs(199)) and not (inputs(147));
    layer0_outputs(8018) <= inputs(194);
    layer0_outputs(8019) <= (inputs(16)) and not (inputs(160));
    layer0_outputs(8020) <= not(inputs(10));
    layer0_outputs(8021) <= (inputs(187)) or (inputs(49));
    layer0_outputs(8022) <= not((inputs(178)) or (inputs(245)));
    layer0_outputs(8023) <= not(inputs(149)) or (inputs(124));
    layer0_outputs(8024) <= (inputs(13)) or (inputs(2));
    layer0_outputs(8025) <= (inputs(176)) or (inputs(181));
    layer0_outputs(8026) <= not(inputs(221));
    layer0_outputs(8027) <= not(inputs(144)) or (inputs(0));
    layer0_outputs(8028) <= not(inputs(203)) or (inputs(117));
    layer0_outputs(8029) <= (inputs(115)) and not (inputs(19));
    layer0_outputs(8030) <= not((inputs(247)) and (inputs(172)));
    layer0_outputs(8031) <= not(inputs(146));
    layer0_outputs(8032) <= not(inputs(178)) or (inputs(179));
    layer0_outputs(8033) <= (inputs(50)) or (inputs(33));
    layer0_outputs(8034) <= (inputs(119)) or (inputs(237));
    layer0_outputs(8035) <= (inputs(96)) and not (inputs(77));
    layer0_outputs(8036) <= (inputs(200)) or (inputs(124));
    layer0_outputs(8037) <= not((inputs(115)) xor (inputs(173)));
    layer0_outputs(8038) <= (inputs(102)) and not (inputs(4));
    layer0_outputs(8039) <= (inputs(189)) and not (inputs(154));
    layer0_outputs(8040) <= not((inputs(229)) or (inputs(224)));
    layer0_outputs(8041) <= (inputs(175)) or (inputs(146));
    layer0_outputs(8042) <= (inputs(36)) or (inputs(2));
    layer0_outputs(8043) <= not(inputs(192));
    layer0_outputs(8044) <= (inputs(205)) or (inputs(133));
    layer0_outputs(8045) <= (inputs(161)) and (inputs(158));
    layer0_outputs(8046) <= not(inputs(170));
    layer0_outputs(8047) <= (inputs(53)) and not (inputs(144));
    layer0_outputs(8048) <= not((inputs(67)) or (inputs(230)));
    layer0_outputs(8049) <= (inputs(210)) and not (inputs(142));
    layer0_outputs(8050) <= (inputs(97)) and not (inputs(121));
    layer0_outputs(8051) <= not(inputs(54));
    layer0_outputs(8052) <= inputs(140);
    layer0_outputs(8053) <= not((inputs(82)) xor (inputs(111)));
    layer0_outputs(8054) <= (inputs(58)) xor (inputs(43));
    layer0_outputs(8055) <= not(inputs(113)) or (inputs(72));
    layer0_outputs(8056) <= not(inputs(186)) or (inputs(106));
    layer0_outputs(8057) <= not(inputs(146));
    layer0_outputs(8058) <= (inputs(242)) or (inputs(39));
    layer0_outputs(8059) <= inputs(16);
    layer0_outputs(8060) <= (inputs(143)) xor (inputs(204));
    layer0_outputs(8061) <= not((inputs(174)) or (inputs(199)));
    layer0_outputs(8062) <= inputs(119);
    layer0_outputs(8063) <= not((inputs(100)) or (inputs(141)));
    layer0_outputs(8064) <= (inputs(201)) and not (inputs(40));
    layer0_outputs(8065) <= (inputs(230)) or (inputs(176));
    layer0_outputs(8066) <= not(inputs(157));
    layer0_outputs(8067) <= not(inputs(187));
    layer0_outputs(8068) <= (inputs(60)) and not (inputs(231));
    layer0_outputs(8069) <= not(inputs(225));
    layer0_outputs(8070) <= not((inputs(254)) and (inputs(12)));
    layer0_outputs(8071) <= not(inputs(224)) or (inputs(109));
    layer0_outputs(8072) <= (inputs(144)) or (inputs(34));
    layer0_outputs(8073) <= inputs(7);
    layer0_outputs(8074) <= (inputs(123)) and not (inputs(194));
    layer0_outputs(8075) <= not(inputs(158));
    layer0_outputs(8076) <= (inputs(240)) or (inputs(64));
    layer0_outputs(8077) <= not(inputs(58));
    layer0_outputs(8078) <= (inputs(59)) or (inputs(75));
    layer0_outputs(8079) <= (inputs(150)) and not (inputs(233));
    layer0_outputs(8080) <= not((inputs(204)) or (inputs(11)));
    layer0_outputs(8081) <= not((inputs(87)) and (inputs(143)));
    layer0_outputs(8082) <= (inputs(112)) and not (inputs(87));
    layer0_outputs(8083) <= (inputs(191)) and not (inputs(104));
    layer0_outputs(8084) <= inputs(188);
    layer0_outputs(8085) <= (inputs(212)) and not (inputs(53));
    layer0_outputs(8086) <= not((inputs(205)) or (inputs(23)));
    layer0_outputs(8087) <= not(inputs(96)) or (inputs(1));
    layer0_outputs(8088) <= not((inputs(99)) or (inputs(140)));
    layer0_outputs(8089) <= not(inputs(187)) or (inputs(184));
    layer0_outputs(8090) <= inputs(120);
    layer0_outputs(8091) <= (inputs(188)) and not (inputs(110));
    layer0_outputs(8092) <= (inputs(195)) and not (inputs(2));
    layer0_outputs(8093) <= not((inputs(2)) or (inputs(200)));
    layer0_outputs(8094) <= not((inputs(159)) and (inputs(2)));
    layer0_outputs(8095) <= not((inputs(144)) xor (inputs(163)));
    layer0_outputs(8096) <= inputs(149);
    layer0_outputs(8097) <= (inputs(241)) or (inputs(202));
    layer0_outputs(8098) <= (inputs(251)) or (inputs(163));
    layer0_outputs(8099) <= not((inputs(185)) and (inputs(224)));
    layer0_outputs(8100) <= not(inputs(178));
    layer0_outputs(8101) <= not(inputs(127));
    layer0_outputs(8102) <= (inputs(253)) or (inputs(41));
    layer0_outputs(8103) <= not((inputs(189)) or (inputs(239)));
    layer0_outputs(8104) <= not(inputs(6));
    layer0_outputs(8105) <= '1';
    layer0_outputs(8106) <= not((inputs(35)) or (inputs(206)));
    layer0_outputs(8107) <= not(inputs(151)) or (inputs(185));
    layer0_outputs(8108) <= not((inputs(239)) or (inputs(246)));
    layer0_outputs(8109) <= not(inputs(229));
    layer0_outputs(8110) <= not(inputs(152));
    layer0_outputs(8111) <= inputs(154);
    layer0_outputs(8112) <= not((inputs(107)) or (inputs(15)));
    layer0_outputs(8113) <= not((inputs(200)) or (inputs(206)));
    layer0_outputs(8114) <= not((inputs(162)) or (inputs(161)));
    layer0_outputs(8115) <= not((inputs(67)) xor (inputs(128)));
    layer0_outputs(8116) <= not(inputs(61));
    layer0_outputs(8117) <= not(inputs(240));
    layer0_outputs(8118) <= inputs(35);
    layer0_outputs(8119) <= not(inputs(122)) or (inputs(181));
    layer0_outputs(8120) <= (inputs(199)) xor (inputs(89));
    layer0_outputs(8121) <= (inputs(89)) and not (inputs(81));
    layer0_outputs(8122) <= (inputs(17)) or (inputs(155));
    layer0_outputs(8123) <= not(inputs(22));
    layer0_outputs(8124) <= (inputs(235)) or (inputs(206));
    layer0_outputs(8125) <= inputs(209);
    layer0_outputs(8126) <= (inputs(34)) or (inputs(21));
    layer0_outputs(8127) <= inputs(125);
    layer0_outputs(8128) <= not(inputs(86));
    layer0_outputs(8129) <= not((inputs(56)) and (inputs(195)));
    layer0_outputs(8130) <= not((inputs(179)) or (inputs(11)));
    layer0_outputs(8131) <= (inputs(244)) and (inputs(226));
    layer0_outputs(8132) <= not((inputs(190)) or (inputs(117)));
    layer0_outputs(8133) <= not((inputs(124)) xor (inputs(92)));
    layer0_outputs(8134) <= not(inputs(215));
    layer0_outputs(8135) <= (inputs(177)) or (inputs(117));
    layer0_outputs(8136) <= not(inputs(133)) or (inputs(177));
    layer0_outputs(8137) <= not((inputs(151)) or (inputs(221)));
    layer0_outputs(8138) <= (inputs(24)) xor (inputs(72));
    layer0_outputs(8139) <= (inputs(100)) and (inputs(22));
    layer0_outputs(8140) <= not(inputs(206));
    layer0_outputs(8141) <= not(inputs(41));
    layer0_outputs(8142) <= not((inputs(171)) xor (inputs(236)));
    layer0_outputs(8143) <= not((inputs(125)) xor (inputs(19)));
    layer0_outputs(8144) <= not(inputs(160));
    layer0_outputs(8145) <= not(inputs(57));
    layer0_outputs(8146) <= not(inputs(137));
    layer0_outputs(8147) <= inputs(250);
    layer0_outputs(8148) <= not((inputs(87)) and (inputs(244)));
    layer0_outputs(8149) <= not(inputs(18));
    layer0_outputs(8150) <= not((inputs(169)) or (inputs(63)));
    layer0_outputs(8151) <= not(inputs(91));
    layer0_outputs(8152) <= inputs(221);
    layer0_outputs(8153) <= not(inputs(188)) or (inputs(32));
    layer0_outputs(8154) <= not((inputs(143)) or (inputs(12)));
    layer0_outputs(8155) <= not((inputs(10)) xor (inputs(43)));
    layer0_outputs(8156) <= not((inputs(35)) or (inputs(17)));
    layer0_outputs(8157) <= (inputs(209)) and not (inputs(1));
    layer0_outputs(8158) <= not((inputs(255)) and (inputs(15)));
    layer0_outputs(8159) <= not(inputs(214));
    layer0_outputs(8160) <= inputs(67);
    layer0_outputs(8161) <= inputs(174);
    layer0_outputs(8162) <= not(inputs(116)) or (inputs(2));
    layer0_outputs(8163) <= (inputs(138)) or (inputs(149));
    layer0_outputs(8164) <= not(inputs(46));
    layer0_outputs(8165) <= not(inputs(68));
    layer0_outputs(8166) <= not(inputs(201)) or (inputs(203));
    layer0_outputs(8167) <= inputs(151);
    layer0_outputs(8168) <= not((inputs(242)) xor (inputs(64)));
    layer0_outputs(8169) <= not((inputs(79)) xor (inputs(141)));
    layer0_outputs(8170) <= (inputs(83)) or (inputs(88));
    layer0_outputs(8171) <= not((inputs(199)) and (inputs(210)));
    layer0_outputs(8172) <= (inputs(165)) and not (inputs(166));
    layer0_outputs(8173) <= not(inputs(98)) or (inputs(238));
    layer0_outputs(8174) <= (inputs(197)) and not (inputs(101));
    layer0_outputs(8175) <= not((inputs(206)) xor (inputs(85)));
    layer0_outputs(8176) <= inputs(100);
    layer0_outputs(8177) <= (inputs(169)) xor (inputs(171));
    layer0_outputs(8178) <= (inputs(115)) or (inputs(130));
    layer0_outputs(8179) <= (inputs(89)) xor (inputs(188));
    layer0_outputs(8180) <= inputs(189);
    layer0_outputs(8181) <= (inputs(222)) and not (inputs(200));
    layer0_outputs(8182) <= inputs(133);
    layer0_outputs(8183) <= (inputs(246)) xor (inputs(198));
    layer0_outputs(8184) <= not(inputs(237));
    layer0_outputs(8185) <= not((inputs(131)) xor (inputs(101)));
    layer0_outputs(8186) <= (inputs(57)) xor (inputs(88));
    layer0_outputs(8187) <= not((inputs(126)) or (inputs(0)));
    layer0_outputs(8188) <= (inputs(72)) and not (inputs(41));
    layer0_outputs(8189) <= not(inputs(232)) or (inputs(185));
    layer0_outputs(8190) <= (inputs(37)) or (inputs(5));
    layer0_outputs(8191) <= not(inputs(230));
    layer0_outputs(8192) <= (inputs(195)) and not (inputs(239));
    layer0_outputs(8193) <= (inputs(71)) and not (inputs(120));
    layer0_outputs(8194) <= (inputs(230)) and not (inputs(20));
    layer0_outputs(8195) <= (inputs(183)) xor (inputs(125));
    layer0_outputs(8196) <= inputs(131);
    layer0_outputs(8197) <= not((inputs(200)) and (inputs(218)));
    layer0_outputs(8198) <= not((inputs(161)) or (inputs(218)));
    layer0_outputs(8199) <= not(inputs(71));
    layer0_outputs(8200) <= '1';
    layer0_outputs(8201) <= (inputs(238)) xor (inputs(143));
    layer0_outputs(8202) <= inputs(235);
    layer0_outputs(8203) <= not(inputs(45));
    layer0_outputs(8204) <= (inputs(234)) or (inputs(224));
    layer0_outputs(8205) <= (inputs(208)) or (inputs(32));
    layer0_outputs(8206) <= inputs(167);
    layer0_outputs(8207) <= (inputs(135)) and not (inputs(133));
    layer0_outputs(8208) <= (inputs(76)) and not (inputs(253));
    layer0_outputs(8209) <= (inputs(10)) or (inputs(247));
    layer0_outputs(8210) <= (inputs(195)) and not (inputs(19));
    layer0_outputs(8211) <= not(inputs(187)) or (inputs(5));
    layer0_outputs(8212) <= not(inputs(147));
    layer0_outputs(8213) <= inputs(111);
    layer0_outputs(8214) <= (inputs(172)) and not (inputs(63));
    layer0_outputs(8215) <= (inputs(235)) and not (inputs(97));
    layer0_outputs(8216) <= '0';
    layer0_outputs(8217) <= not(inputs(167));
    layer0_outputs(8218) <= not(inputs(166)) or (inputs(198));
    layer0_outputs(8219) <= (inputs(79)) xor (inputs(226));
    layer0_outputs(8220) <= (inputs(133)) xor (inputs(152));
    layer0_outputs(8221) <= not(inputs(164));
    layer0_outputs(8222) <= (inputs(65)) or (inputs(103));
    layer0_outputs(8223) <= not(inputs(98));
    layer0_outputs(8224) <= (inputs(43)) and not (inputs(234));
    layer0_outputs(8225) <= (inputs(244)) and not (inputs(120));
    layer0_outputs(8226) <= inputs(130);
    layer0_outputs(8227) <= not((inputs(241)) or (inputs(15)));
    layer0_outputs(8228) <= not(inputs(85)) or (inputs(164));
    layer0_outputs(8229) <= (inputs(211)) and (inputs(129));
    layer0_outputs(8230) <= inputs(201);
    layer0_outputs(8231) <= not((inputs(80)) or (inputs(5)));
    layer0_outputs(8232) <= inputs(21);
    layer0_outputs(8233) <= (inputs(22)) and not (inputs(18));
    layer0_outputs(8234) <= (inputs(58)) and not (inputs(176));
    layer0_outputs(8235) <= not(inputs(40)) or (inputs(113));
    layer0_outputs(8236) <= not(inputs(104)) or (inputs(102));
    layer0_outputs(8237) <= (inputs(137)) and not (inputs(178));
    layer0_outputs(8238) <= (inputs(29)) and not (inputs(142));
    layer0_outputs(8239) <= inputs(85);
    layer0_outputs(8240) <= not(inputs(255));
    layer0_outputs(8241) <= not(inputs(68));
    layer0_outputs(8242) <= inputs(233);
    layer0_outputs(8243) <= not((inputs(107)) and (inputs(23)));
    layer0_outputs(8244) <= not((inputs(120)) and (inputs(120)));
    layer0_outputs(8245) <= not(inputs(150));
    layer0_outputs(8246) <= not(inputs(149)) or (inputs(44));
    layer0_outputs(8247) <= not(inputs(68));
    layer0_outputs(8248) <= inputs(94);
    layer0_outputs(8249) <= (inputs(37)) xor (inputs(254));
    layer0_outputs(8250) <= not(inputs(90)) or (inputs(192));
    layer0_outputs(8251) <= not(inputs(111));
    layer0_outputs(8252) <= inputs(98);
    layer0_outputs(8253) <= not(inputs(173));
    layer0_outputs(8254) <= not(inputs(224)) or (inputs(181));
    layer0_outputs(8255) <= '0';
    layer0_outputs(8256) <= not(inputs(204)) or (inputs(32));
    layer0_outputs(8257) <= (inputs(236)) and not (inputs(156));
    layer0_outputs(8258) <= inputs(144);
    layer0_outputs(8259) <= '0';
    layer0_outputs(8260) <= (inputs(133)) and not (inputs(34));
    layer0_outputs(8261) <= not((inputs(133)) and (inputs(233)));
    layer0_outputs(8262) <= not((inputs(47)) or (inputs(52)));
    layer0_outputs(8263) <= not((inputs(114)) xor (inputs(156)));
    layer0_outputs(8264) <= '1';
    layer0_outputs(8265) <= not(inputs(45));
    layer0_outputs(8266) <= not((inputs(72)) or (inputs(235)));
    layer0_outputs(8267) <= not(inputs(232));
    layer0_outputs(8268) <= (inputs(176)) or (inputs(217));
    layer0_outputs(8269) <= inputs(29);
    layer0_outputs(8270) <= inputs(64);
    layer0_outputs(8271) <= not((inputs(231)) and (inputs(101)));
    layer0_outputs(8272) <= (inputs(181)) or (inputs(254));
    layer0_outputs(8273) <= (inputs(88)) and not (inputs(233));
    layer0_outputs(8274) <= not((inputs(181)) or (inputs(125)));
    layer0_outputs(8275) <= not(inputs(135));
    layer0_outputs(8276) <= not(inputs(244)) or (inputs(86));
    layer0_outputs(8277) <= (inputs(35)) or (inputs(253));
    layer0_outputs(8278) <= not(inputs(90)) or (inputs(221));
    layer0_outputs(8279) <= not(inputs(31));
    layer0_outputs(8280) <= not(inputs(8));
    layer0_outputs(8281) <= not((inputs(11)) or (inputs(66)));
    layer0_outputs(8282) <= '0';
    layer0_outputs(8283) <= not(inputs(82)) or (inputs(189));
    layer0_outputs(8284) <= not(inputs(118));
    layer0_outputs(8285) <= not(inputs(86));
    layer0_outputs(8286) <= inputs(245);
    layer0_outputs(8287) <= not(inputs(105));
    layer0_outputs(8288) <= not((inputs(149)) or (inputs(48)));
    layer0_outputs(8289) <= not(inputs(231)) or (inputs(216));
    layer0_outputs(8290) <= not(inputs(193)) or (inputs(48));
    layer0_outputs(8291) <= not(inputs(124));
    layer0_outputs(8292) <= '0';
    layer0_outputs(8293) <= inputs(40);
    layer0_outputs(8294) <= not(inputs(71));
    layer0_outputs(8295) <= inputs(110);
    layer0_outputs(8296) <= not((inputs(67)) xor (inputs(20)));
    layer0_outputs(8297) <= (inputs(65)) or (inputs(29));
    layer0_outputs(8298) <= inputs(49);
    layer0_outputs(8299) <= not((inputs(162)) or (inputs(203)));
    layer0_outputs(8300) <= not((inputs(149)) or (inputs(116)));
    layer0_outputs(8301) <= not((inputs(151)) or (inputs(227)));
    layer0_outputs(8302) <= not(inputs(91));
    layer0_outputs(8303) <= not((inputs(200)) and (inputs(166)));
    layer0_outputs(8304) <= not((inputs(110)) or (inputs(182)));
    layer0_outputs(8305) <= not((inputs(174)) or (inputs(179)));
    layer0_outputs(8306) <= not(inputs(173));
    layer0_outputs(8307) <= not(inputs(56));
    layer0_outputs(8308) <= inputs(133);
    layer0_outputs(8309) <= (inputs(182)) and not (inputs(70));
    layer0_outputs(8310) <= not(inputs(199)) or (inputs(175));
    layer0_outputs(8311) <= not(inputs(234));
    layer0_outputs(8312) <= not((inputs(248)) or (inputs(160)));
    layer0_outputs(8313) <= (inputs(196)) and not (inputs(132));
    layer0_outputs(8314) <= inputs(126);
    layer0_outputs(8315) <= not(inputs(161));
    layer0_outputs(8316) <= not(inputs(1));
    layer0_outputs(8317) <= (inputs(43)) and not (inputs(16));
    layer0_outputs(8318) <= '0';
    layer0_outputs(8319) <= not((inputs(160)) xor (inputs(228)));
    layer0_outputs(8320) <= not((inputs(193)) and (inputs(1)));
    layer0_outputs(8321) <= (inputs(131)) xor (inputs(64));
    layer0_outputs(8322) <= not((inputs(220)) or (inputs(107)));
    layer0_outputs(8323) <= (inputs(1)) xor (inputs(151));
    layer0_outputs(8324) <= (inputs(198)) and (inputs(203));
    layer0_outputs(8325) <= (inputs(73)) or (inputs(90));
    layer0_outputs(8326) <= not(inputs(79)) or (inputs(207));
    layer0_outputs(8327) <= not(inputs(4)) or (inputs(190));
    layer0_outputs(8328) <= inputs(202);
    layer0_outputs(8329) <= not((inputs(69)) or (inputs(185)));
    layer0_outputs(8330) <= not((inputs(195)) xor (inputs(59)));
    layer0_outputs(8331) <= inputs(146);
    layer0_outputs(8332) <= inputs(172);
    layer0_outputs(8333) <= not((inputs(80)) or (inputs(167)));
    layer0_outputs(8334) <= (inputs(50)) and (inputs(243));
    layer0_outputs(8335) <= not(inputs(55));
    layer0_outputs(8336) <= not((inputs(5)) or (inputs(180)));
    layer0_outputs(8337) <= not((inputs(243)) xor (inputs(12)));
    layer0_outputs(8338) <= not(inputs(83));
    layer0_outputs(8339) <= not(inputs(155)) or (inputs(15));
    layer0_outputs(8340) <= '1';
    layer0_outputs(8341) <= inputs(59);
    layer0_outputs(8342) <= (inputs(130)) or (inputs(242));
    layer0_outputs(8343) <= inputs(130);
    layer0_outputs(8344) <= (inputs(163)) or (inputs(49));
    layer0_outputs(8345) <= not((inputs(162)) or (inputs(87)));
    layer0_outputs(8346) <= not((inputs(176)) or (inputs(48)));
    layer0_outputs(8347) <= not(inputs(183));
    layer0_outputs(8348) <= not((inputs(241)) xor (inputs(165)));
    layer0_outputs(8349) <= not(inputs(1));
    layer0_outputs(8350) <= (inputs(60)) xor (inputs(43));
    layer0_outputs(8351) <= not(inputs(127)) or (inputs(13));
    layer0_outputs(8352) <= inputs(113);
    layer0_outputs(8353) <= not((inputs(145)) or (inputs(14)));
    layer0_outputs(8354) <= (inputs(5)) or (inputs(246));
    layer0_outputs(8355) <= not((inputs(2)) xor (inputs(175)));
    layer0_outputs(8356) <= not(inputs(184)) or (inputs(7));
    layer0_outputs(8357) <= (inputs(49)) or (inputs(190));
    layer0_outputs(8358) <= (inputs(113)) and not (inputs(28));
    layer0_outputs(8359) <= (inputs(243)) xor (inputs(95));
    layer0_outputs(8360) <= inputs(162);
    layer0_outputs(8361) <= inputs(57);
    layer0_outputs(8362) <= not(inputs(232)) or (inputs(126));
    layer0_outputs(8363) <= not((inputs(56)) or (inputs(5)));
    layer0_outputs(8364) <= not(inputs(49));
    layer0_outputs(8365) <= not(inputs(144)) or (inputs(143));
    layer0_outputs(8366) <= not((inputs(111)) xor (inputs(9)));
    layer0_outputs(8367) <= '0';
    layer0_outputs(8368) <= not(inputs(135)) or (inputs(92));
    layer0_outputs(8369) <= inputs(187);
    layer0_outputs(8370) <= not(inputs(42)) or (inputs(99));
    layer0_outputs(8371) <= not(inputs(69));
    layer0_outputs(8372) <= (inputs(176)) xor (inputs(88));
    layer0_outputs(8373) <= not((inputs(190)) xor (inputs(139)));
    layer0_outputs(8374) <= not(inputs(140)) or (inputs(185));
    layer0_outputs(8375) <= not((inputs(205)) or (inputs(167)));
    layer0_outputs(8376) <= not(inputs(109));
    layer0_outputs(8377) <= '1';
    layer0_outputs(8378) <= (inputs(218)) or (inputs(77));
    layer0_outputs(8379) <= (inputs(200)) or (inputs(255));
    layer0_outputs(8380) <= (inputs(11)) or (inputs(169));
    layer0_outputs(8381) <= inputs(21);
    layer0_outputs(8382) <= '0';
    layer0_outputs(8383) <= not(inputs(88));
    layer0_outputs(8384) <= (inputs(37)) xor (inputs(247));
    layer0_outputs(8385) <= not(inputs(221));
    layer0_outputs(8386) <= (inputs(8)) and not (inputs(15));
    layer0_outputs(8387) <= inputs(198);
    layer0_outputs(8388) <= not((inputs(175)) or (inputs(209)));
    layer0_outputs(8389) <= not(inputs(136)) or (inputs(252));
    layer0_outputs(8390) <= not((inputs(204)) and (inputs(182)));
    layer0_outputs(8391) <= not((inputs(226)) or (inputs(193)));
    layer0_outputs(8392) <= inputs(47);
    layer0_outputs(8393) <= not((inputs(187)) xor (inputs(37)));
    layer0_outputs(8394) <= inputs(56);
    layer0_outputs(8395) <= inputs(92);
    layer0_outputs(8396) <= inputs(178);
    layer0_outputs(8397) <= inputs(121);
    layer0_outputs(8398) <= not(inputs(119)) or (inputs(10));
    layer0_outputs(8399) <= not((inputs(250)) xor (inputs(227)));
    layer0_outputs(8400) <= not(inputs(187)) or (inputs(126));
    layer0_outputs(8401) <= inputs(149);
    layer0_outputs(8402) <= '0';
    layer0_outputs(8403) <= not(inputs(134));
    layer0_outputs(8404) <= not((inputs(181)) xor (inputs(39)));
    layer0_outputs(8405) <= (inputs(205)) and not (inputs(145));
    layer0_outputs(8406) <= not((inputs(161)) xor (inputs(16)));
    layer0_outputs(8407) <= not((inputs(138)) xor (inputs(61)));
    layer0_outputs(8408) <= not((inputs(186)) xor (inputs(147)));
    layer0_outputs(8409) <= not(inputs(94)) or (inputs(237));
    layer0_outputs(8410) <= not((inputs(117)) or (inputs(205)));
    layer0_outputs(8411) <= not((inputs(106)) xor (inputs(48)));
    layer0_outputs(8412) <= not(inputs(36)) or (inputs(144));
    layer0_outputs(8413) <= not(inputs(213));
    layer0_outputs(8414) <= (inputs(2)) or (inputs(61));
    layer0_outputs(8415) <= inputs(99);
    layer0_outputs(8416) <= (inputs(170)) xor (inputs(162));
    layer0_outputs(8417) <= not((inputs(135)) or (inputs(7)));
    layer0_outputs(8418) <= (inputs(46)) or (inputs(16));
    layer0_outputs(8419) <= inputs(185);
    layer0_outputs(8420) <= (inputs(246)) or (inputs(95));
    layer0_outputs(8421) <= inputs(212);
    layer0_outputs(8422) <= not(inputs(212)) or (inputs(111));
    layer0_outputs(8423) <= not(inputs(102));
    layer0_outputs(8424) <= (inputs(240)) and not (inputs(42));
    layer0_outputs(8425) <= not(inputs(203)) or (inputs(15));
    layer0_outputs(8426) <= not(inputs(241)) or (inputs(100));
    layer0_outputs(8427) <= not((inputs(143)) or (inputs(2)));
    layer0_outputs(8428) <= (inputs(181)) and not (inputs(148));
    layer0_outputs(8429) <= inputs(146);
    layer0_outputs(8430) <= (inputs(101)) and not (inputs(108));
    layer0_outputs(8431) <= not(inputs(145));
    layer0_outputs(8432) <= not(inputs(166)) or (inputs(191));
    layer0_outputs(8433) <= not(inputs(86));
    layer0_outputs(8434) <= not(inputs(235));
    layer0_outputs(8435) <= not((inputs(73)) xor (inputs(62)));
    layer0_outputs(8436) <= (inputs(81)) and not (inputs(204));
    layer0_outputs(8437) <= not(inputs(212)) or (inputs(47));
    layer0_outputs(8438) <= (inputs(117)) and (inputs(75));
    layer0_outputs(8439) <= (inputs(164)) and not (inputs(58));
    layer0_outputs(8440) <= not(inputs(131));
    layer0_outputs(8441) <= not(inputs(174));
    layer0_outputs(8442) <= inputs(139);
    layer0_outputs(8443) <= '1';
    layer0_outputs(8444) <= not((inputs(90)) xor (inputs(87)));
    layer0_outputs(8445) <= inputs(17);
    layer0_outputs(8446) <= not((inputs(198)) or (inputs(182)));
    layer0_outputs(8447) <= not((inputs(205)) and (inputs(52)));
    layer0_outputs(8448) <= not(inputs(36));
    layer0_outputs(8449) <= not(inputs(203)) or (inputs(164));
    layer0_outputs(8450) <= not((inputs(232)) and (inputs(147)));
    layer0_outputs(8451) <= (inputs(245)) and not (inputs(61));
    layer0_outputs(8452) <= not(inputs(245)) or (inputs(5));
    layer0_outputs(8453) <= not((inputs(53)) xor (inputs(9)));
    layer0_outputs(8454) <= not(inputs(222));
    layer0_outputs(8455) <= (inputs(58)) and (inputs(74));
    layer0_outputs(8456) <= '1';
    layer0_outputs(8457) <= not(inputs(128));
    layer0_outputs(8458) <= not((inputs(126)) or (inputs(127)));
    layer0_outputs(8459) <= inputs(118);
    layer0_outputs(8460) <= not(inputs(157)) or (inputs(29));
    layer0_outputs(8461) <= not(inputs(57)) or (inputs(161));
    layer0_outputs(8462) <= inputs(100);
    layer0_outputs(8463) <= inputs(165);
    layer0_outputs(8464) <= not(inputs(137));
    layer0_outputs(8465) <= (inputs(251)) xor (inputs(187));
    layer0_outputs(8466) <= inputs(54);
    layer0_outputs(8467) <= inputs(214);
    layer0_outputs(8468) <= (inputs(132)) and not (inputs(251));
    layer0_outputs(8469) <= (inputs(134)) and not (inputs(123));
    layer0_outputs(8470) <= (inputs(23)) or (inputs(129));
    layer0_outputs(8471) <= not((inputs(64)) or (inputs(53)));
    layer0_outputs(8472) <= (inputs(178)) and (inputs(131));
    layer0_outputs(8473) <= (inputs(158)) xor (inputs(235));
    layer0_outputs(8474) <= not((inputs(114)) or (inputs(115)));
    layer0_outputs(8475) <= inputs(96);
    layer0_outputs(8476) <= '0';
    layer0_outputs(8477) <= not((inputs(221)) or (inputs(119)));
    layer0_outputs(8478) <= inputs(202);
    layer0_outputs(8479) <= (inputs(151)) and not (inputs(115));
    layer0_outputs(8480) <= not(inputs(147)) or (inputs(14));
    layer0_outputs(8481) <= not((inputs(3)) or (inputs(180)));
    layer0_outputs(8482) <= (inputs(107)) and not (inputs(191));
    layer0_outputs(8483) <= (inputs(166)) or (inputs(24));
    layer0_outputs(8484) <= (inputs(197)) and not (inputs(141));
    layer0_outputs(8485) <= (inputs(64)) and not (inputs(242));
    layer0_outputs(8486) <= (inputs(21)) or (inputs(25));
    layer0_outputs(8487) <= not(inputs(5)) or (inputs(172));
    layer0_outputs(8488) <= not(inputs(176));
    layer0_outputs(8489) <= not(inputs(230)) or (inputs(61));
    layer0_outputs(8490) <= not(inputs(8)) or (inputs(223));
    layer0_outputs(8491) <= (inputs(64)) or (inputs(38));
    layer0_outputs(8492) <= not(inputs(154)) or (inputs(101));
    layer0_outputs(8493) <= not((inputs(27)) xor (inputs(238)));
    layer0_outputs(8494) <= inputs(50);
    layer0_outputs(8495) <= not((inputs(166)) or (inputs(30)));
    layer0_outputs(8496) <= (inputs(252)) xor (inputs(8));
    layer0_outputs(8497) <= (inputs(44)) and (inputs(117));
    layer0_outputs(8498) <= (inputs(136)) or (inputs(117));
    layer0_outputs(8499) <= inputs(155);
    layer0_outputs(8500) <= (inputs(30)) or (inputs(27));
    layer0_outputs(8501) <= not(inputs(120));
    layer0_outputs(8502) <= (inputs(28)) or (inputs(111));
    layer0_outputs(8503) <= (inputs(171)) xor (inputs(133));
    layer0_outputs(8504) <= (inputs(187)) or (inputs(46));
    layer0_outputs(8505) <= not(inputs(111)) or (inputs(220));
    layer0_outputs(8506) <= (inputs(212)) or (inputs(194));
    layer0_outputs(8507) <= inputs(118);
    layer0_outputs(8508) <= not(inputs(248));
    layer0_outputs(8509) <= (inputs(166)) and not (inputs(160));
    layer0_outputs(8510) <= inputs(37);
    layer0_outputs(8511) <= (inputs(186)) and not (inputs(105));
    layer0_outputs(8512) <= (inputs(8)) and not (inputs(241));
    layer0_outputs(8513) <= inputs(166);
    layer0_outputs(8514) <= not((inputs(119)) xor (inputs(184)));
    layer0_outputs(8515) <= inputs(181);
    layer0_outputs(8516) <= not(inputs(207)) or (inputs(15));
    layer0_outputs(8517) <= not((inputs(38)) or (inputs(16)));
    layer0_outputs(8518) <= inputs(141);
    layer0_outputs(8519) <= (inputs(147)) and not (inputs(107));
    layer0_outputs(8520) <= inputs(4);
    layer0_outputs(8521) <= inputs(201);
    layer0_outputs(8522) <= not((inputs(169)) or (inputs(138)));
    layer0_outputs(8523) <= inputs(91);
    layer0_outputs(8524) <= '1';
    layer0_outputs(8525) <= (inputs(150)) or (inputs(238));
    layer0_outputs(8526) <= not((inputs(42)) or (inputs(79)));
    layer0_outputs(8527) <= not((inputs(241)) or (inputs(175)));
    layer0_outputs(8528) <= not((inputs(87)) and (inputs(221)));
    layer0_outputs(8529) <= (inputs(165)) and not (inputs(16));
    layer0_outputs(8530) <= not(inputs(235));
    layer0_outputs(8531) <= not(inputs(219));
    layer0_outputs(8532) <= not((inputs(83)) or (inputs(10)));
    layer0_outputs(8533) <= inputs(188);
    layer0_outputs(8534) <= inputs(54);
    layer0_outputs(8535) <= not(inputs(77)) or (inputs(220));
    layer0_outputs(8536) <= (inputs(45)) or (inputs(69));
    layer0_outputs(8537) <= not(inputs(238));
    layer0_outputs(8538) <= (inputs(24)) and (inputs(248));
    layer0_outputs(8539) <= (inputs(255)) or (inputs(230));
    layer0_outputs(8540) <= not(inputs(121)) or (inputs(163));
    layer0_outputs(8541) <= not(inputs(1));
    layer0_outputs(8542) <= not(inputs(7));
    layer0_outputs(8543) <= not(inputs(135));
    layer0_outputs(8544) <= (inputs(189)) and not (inputs(242));
    layer0_outputs(8545) <= not((inputs(120)) xor (inputs(121)));
    layer0_outputs(8546) <= inputs(41);
    layer0_outputs(8547) <= (inputs(101)) and not (inputs(244));
    layer0_outputs(8548) <= not(inputs(198));
    layer0_outputs(8549) <= not(inputs(24)) or (inputs(115));
    layer0_outputs(8550) <= not((inputs(69)) xor (inputs(20)));
    layer0_outputs(8551) <= not(inputs(42)) or (inputs(221));
    layer0_outputs(8552) <= not(inputs(22));
    layer0_outputs(8553) <= (inputs(146)) and not (inputs(235));
    layer0_outputs(8554) <= inputs(24);
    layer0_outputs(8555) <= not(inputs(106)) or (inputs(193));
    layer0_outputs(8556) <= (inputs(227)) and not (inputs(155));
    layer0_outputs(8557) <= not(inputs(108));
    layer0_outputs(8558) <= (inputs(54)) or (inputs(226));
    layer0_outputs(8559) <= inputs(36);
    layer0_outputs(8560) <= not(inputs(197));
    layer0_outputs(8561) <= not(inputs(142)) or (inputs(93));
    layer0_outputs(8562) <= inputs(234);
    layer0_outputs(8563) <= (inputs(208)) xor (inputs(98));
    layer0_outputs(8564) <= (inputs(108)) and not (inputs(248));
    layer0_outputs(8565) <= not(inputs(113)) or (inputs(64));
    layer0_outputs(8566) <= not(inputs(74));
    layer0_outputs(8567) <= inputs(148);
    layer0_outputs(8568) <= inputs(222);
    layer0_outputs(8569) <= (inputs(193)) and not (inputs(73));
    layer0_outputs(8570) <= inputs(221);
    layer0_outputs(8571) <= not((inputs(102)) xor (inputs(165)));
    layer0_outputs(8572) <= (inputs(194)) and not (inputs(100));
    layer0_outputs(8573) <= inputs(39);
    layer0_outputs(8574) <= not((inputs(204)) xor (inputs(16)));
    layer0_outputs(8575) <= not(inputs(151));
    layer0_outputs(8576) <= (inputs(103)) xor (inputs(135));
    layer0_outputs(8577) <= (inputs(215)) and (inputs(215));
    layer0_outputs(8578) <= '1';
    layer0_outputs(8579) <= not((inputs(253)) or (inputs(236)));
    layer0_outputs(8580) <= inputs(52);
    layer0_outputs(8581) <= (inputs(236)) or (inputs(244));
    layer0_outputs(8582) <= not((inputs(199)) or (inputs(183)));
    layer0_outputs(8583) <= inputs(190);
    layer0_outputs(8584) <= inputs(211);
    layer0_outputs(8585) <= (inputs(227)) and not (inputs(17));
    layer0_outputs(8586) <= (inputs(180)) and not (inputs(29));
    layer0_outputs(8587) <= inputs(114);
    layer0_outputs(8588) <= not((inputs(7)) xor (inputs(214)));
    layer0_outputs(8589) <= not(inputs(118));
    layer0_outputs(8590) <= not(inputs(121));
    layer0_outputs(8591) <= (inputs(156)) or (inputs(205));
    layer0_outputs(8592) <= (inputs(157)) or (inputs(86));
    layer0_outputs(8593) <= inputs(131);
    layer0_outputs(8594) <= not((inputs(170)) xor (inputs(94)));
    layer0_outputs(8595) <= (inputs(131)) and (inputs(196));
    layer0_outputs(8596) <= (inputs(101)) xor (inputs(71));
    layer0_outputs(8597) <= not(inputs(189));
    layer0_outputs(8598) <= not(inputs(220)) or (inputs(59));
    layer0_outputs(8599) <= '1';
    layer0_outputs(8600) <= not((inputs(174)) xor (inputs(123)));
    layer0_outputs(8601) <= not((inputs(99)) xor (inputs(71)));
    layer0_outputs(8602) <= not(inputs(111));
    layer0_outputs(8603) <= not(inputs(254));
    layer0_outputs(8604) <= (inputs(119)) and not (inputs(235));
    layer0_outputs(8605) <= not((inputs(244)) and (inputs(12)));
    layer0_outputs(8606) <= (inputs(47)) and not (inputs(16));
    layer0_outputs(8607) <= inputs(77);
    layer0_outputs(8608) <= not((inputs(184)) xor (inputs(158)));
    layer0_outputs(8609) <= not(inputs(39));
    layer0_outputs(8610) <= not(inputs(43)) or (inputs(254));
    layer0_outputs(8611) <= not(inputs(85));
    layer0_outputs(8612) <= inputs(230);
    layer0_outputs(8613) <= not((inputs(89)) or (inputs(45)));
    layer0_outputs(8614) <= not((inputs(8)) or (inputs(231)));
    layer0_outputs(8615) <= not(inputs(136));
    layer0_outputs(8616) <= (inputs(19)) and not (inputs(140));
    layer0_outputs(8617) <= (inputs(179)) and not (inputs(4));
    layer0_outputs(8618) <= (inputs(233)) and (inputs(135));
    layer0_outputs(8619) <= (inputs(11)) or (inputs(12));
    layer0_outputs(8620) <= inputs(214);
    layer0_outputs(8621) <= not(inputs(117));
    layer0_outputs(8622) <= (inputs(185)) and not (inputs(126));
    layer0_outputs(8623) <= inputs(198);
    layer0_outputs(8624) <= '0';
    layer0_outputs(8625) <= (inputs(43)) or (inputs(114));
    layer0_outputs(8626) <= inputs(132);
    layer0_outputs(8627) <= not((inputs(102)) or (inputs(244)));
    layer0_outputs(8628) <= inputs(21);
    layer0_outputs(8629) <= not(inputs(78));
    layer0_outputs(8630) <= (inputs(173)) xor (inputs(71));
    layer0_outputs(8631) <= not((inputs(11)) and (inputs(173)));
    layer0_outputs(8632) <= not(inputs(140)) or (inputs(191));
    layer0_outputs(8633) <= not((inputs(165)) or (inputs(90)));
    layer0_outputs(8634) <= (inputs(52)) or (inputs(6));
    layer0_outputs(8635) <= not(inputs(230)) or (inputs(238));
    layer0_outputs(8636) <= not((inputs(91)) and (inputs(8)));
    layer0_outputs(8637) <= not(inputs(222));
    layer0_outputs(8638) <= (inputs(88)) and (inputs(14));
    layer0_outputs(8639) <= (inputs(106)) or (inputs(123));
    layer0_outputs(8640) <= (inputs(214)) or (inputs(139));
    layer0_outputs(8641) <= not(inputs(160));
    layer0_outputs(8642) <= (inputs(66)) or (inputs(30));
    layer0_outputs(8643) <= (inputs(151)) or (inputs(206));
    layer0_outputs(8644) <= (inputs(177)) and (inputs(151));
    layer0_outputs(8645) <= (inputs(50)) xor (inputs(75));
    layer0_outputs(8646) <= (inputs(53)) or (inputs(7));
    layer0_outputs(8647) <= (inputs(178)) xor (inputs(58));
    layer0_outputs(8648) <= (inputs(189)) and (inputs(219));
    layer0_outputs(8649) <= not(inputs(59));
    layer0_outputs(8650) <= not(inputs(155));
    layer0_outputs(8651) <= not(inputs(99)) or (inputs(41));
    layer0_outputs(8652) <= (inputs(169)) and not (inputs(39));
    layer0_outputs(8653) <= inputs(213);
    layer0_outputs(8654) <= not((inputs(70)) xor (inputs(177)));
    layer0_outputs(8655) <= not(inputs(45));
    layer0_outputs(8656) <= not((inputs(193)) or (inputs(63)));
    layer0_outputs(8657) <= not(inputs(200)) or (inputs(31));
    layer0_outputs(8658) <= (inputs(23)) and (inputs(25));
    layer0_outputs(8659) <= not((inputs(5)) or (inputs(1)));
    layer0_outputs(8660) <= not(inputs(134));
    layer0_outputs(8661) <= not((inputs(107)) xor (inputs(86)));
    layer0_outputs(8662) <= (inputs(86)) xor (inputs(107));
    layer0_outputs(8663) <= inputs(172);
    layer0_outputs(8664) <= not(inputs(202)) or (inputs(32));
    layer0_outputs(8665) <= (inputs(147)) and not (inputs(46));
    layer0_outputs(8666) <= not((inputs(17)) or (inputs(227)));
    layer0_outputs(8667) <= (inputs(128)) or (inputs(99));
    layer0_outputs(8668) <= '1';
    layer0_outputs(8669) <= not(inputs(190));
    layer0_outputs(8670) <= not(inputs(245)) or (inputs(68));
    layer0_outputs(8671) <= (inputs(105)) and not (inputs(20));
    layer0_outputs(8672) <= inputs(115);
    layer0_outputs(8673) <= inputs(127);
    layer0_outputs(8674) <= not(inputs(156));
    layer0_outputs(8675) <= inputs(9);
    layer0_outputs(8676) <= (inputs(47)) and not (inputs(207));
    layer0_outputs(8677) <= (inputs(250)) and (inputs(146));
    layer0_outputs(8678) <= inputs(197);
    layer0_outputs(8679) <= inputs(182);
    layer0_outputs(8680) <= (inputs(99)) and not (inputs(54));
    layer0_outputs(8681) <= (inputs(18)) or (inputs(74));
    layer0_outputs(8682) <= inputs(102);
    layer0_outputs(8683) <= not(inputs(73)) or (inputs(156));
    layer0_outputs(8684) <= inputs(130);
    layer0_outputs(8685) <= not(inputs(71)) or (inputs(246));
    layer0_outputs(8686) <= '0';
    layer0_outputs(8687) <= (inputs(247)) or (inputs(111));
    layer0_outputs(8688) <= not(inputs(44)) or (inputs(8));
    layer0_outputs(8689) <= not(inputs(38)) or (inputs(223));
    layer0_outputs(8690) <= (inputs(135)) and not (inputs(191));
    layer0_outputs(8691) <= inputs(49);
    layer0_outputs(8692) <= (inputs(70)) and not (inputs(246));
    layer0_outputs(8693) <= (inputs(130)) and (inputs(70));
    layer0_outputs(8694) <= (inputs(211)) and not (inputs(236));
    layer0_outputs(8695) <= inputs(149);
    layer0_outputs(8696) <= inputs(131);
    layer0_outputs(8697) <= not((inputs(232)) or (inputs(2)));
    layer0_outputs(8698) <= (inputs(112)) and not (inputs(126));
    layer0_outputs(8699) <= (inputs(80)) and not (inputs(218));
    layer0_outputs(8700) <= not((inputs(167)) and (inputs(44)));
    layer0_outputs(8701) <= (inputs(221)) and not (inputs(158));
    layer0_outputs(8702) <= '0';
    layer0_outputs(8703) <= not((inputs(148)) or (inputs(22)));
    layer0_outputs(8704) <= inputs(56);
    layer0_outputs(8705) <= inputs(102);
    layer0_outputs(8706) <= not(inputs(135));
    layer0_outputs(8707) <= inputs(192);
    layer0_outputs(8708) <= (inputs(238)) and (inputs(61));
    layer0_outputs(8709) <= not(inputs(77));
    layer0_outputs(8710) <= (inputs(204)) xor (inputs(101));
    layer0_outputs(8711) <= not(inputs(249));
    layer0_outputs(8712) <= (inputs(46)) or (inputs(128));
    layer0_outputs(8713) <= (inputs(93)) and not (inputs(194));
    layer0_outputs(8714) <= inputs(109);
    layer0_outputs(8715) <= not((inputs(153)) or (inputs(148)));
    layer0_outputs(8716) <= '1';
    layer0_outputs(8717) <= not((inputs(0)) and (inputs(146)));
    layer0_outputs(8718) <= not(inputs(214));
    layer0_outputs(8719) <= inputs(141);
    layer0_outputs(8720) <= (inputs(231)) and not (inputs(237));
    layer0_outputs(8721) <= not(inputs(65)) or (inputs(184));
    layer0_outputs(8722) <= not(inputs(103));
    layer0_outputs(8723) <= not(inputs(124));
    layer0_outputs(8724) <= not((inputs(220)) xor (inputs(4)));
    layer0_outputs(8725) <= (inputs(22)) and not (inputs(146));
    layer0_outputs(8726) <= (inputs(164)) xor (inputs(147));
    layer0_outputs(8727) <= not((inputs(107)) or (inputs(61)));
    layer0_outputs(8728) <= not(inputs(236));
    layer0_outputs(8729) <= '0';
    layer0_outputs(8730) <= not(inputs(72));
    layer0_outputs(8731) <= not(inputs(93));
    layer0_outputs(8732) <= not(inputs(11));
    layer0_outputs(8733) <= (inputs(51)) xor (inputs(147));
    layer0_outputs(8734) <= inputs(245);
    layer0_outputs(8735) <= (inputs(250)) or (inputs(55));
    layer0_outputs(8736) <= not((inputs(147)) or (inputs(144)));
    layer0_outputs(8737) <= not((inputs(240)) and (inputs(18)));
    layer0_outputs(8738) <= not(inputs(173));
    layer0_outputs(8739) <= not(inputs(133)) or (inputs(34));
    layer0_outputs(8740) <= (inputs(46)) or (inputs(114));
    layer0_outputs(8741) <= not(inputs(75));
    layer0_outputs(8742) <= not(inputs(23));
    layer0_outputs(8743) <= not((inputs(251)) or (inputs(218)));
    layer0_outputs(8744) <= (inputs(80)) or (inputs(196));
    layer0_outputs(8745) <= not((inputs(106)) and (inputs(198)));
    layer0_outputs(8746) <= not(inputs(235)) or (inputs(78));
    layer0_outputs(8747) <= not(inputs(159));
    layer0_outputs(8748) <= not(inputs(251)) or (inputs(38));
    layer0_outputs(8749) <= inputs(62);
    layer0_outputs(8750) <= (inputs(204)) or (inputs(37));
    layer0_outputs(8751) <= '0';
    layer0_outputs(8752) <= not(inputs(119));
    layer0_outputs(8753) <= not(inputs(214));
    layer0_outputs(8754) <= (inputs(6)) or (inputs(242));
    layer0_outputs(8755) <= (inputs(216)) or (inputs(55));
    layer0_outputs(8756) <= not((inputs(110)) xor (inputs(21)));
    layer0_outputs(8757) <= not(inputs(67)) or (inputs(225));
    layer0_outputs(8758) <= inputs(42);
    layer0_outputs(8759) <= (inputs(197)) and not (inputs(1));
    layer0_outputs(8760) <= not(inputs(99));
    layer0_outputs(8761) <= (inputs(23)) xor (inputs(106));
    layer0_outputs(8762) <= not(inputs(26));
    layer0_outputs(8763) <= not((inputs(225)) or (inputs(18)));
    layer0_outputs(8764) <= (inputs(202)) and (inputs(78));
    layer0_outputs(8765) <= (inputs(254)) and not (inputs(52));
    layer0_outputs(8766) <= (inputs(166)) and not (inputs(188));
    layer0_outputs(8767) <= inputs(164);
    layer0_outputs(8768) <= (inputs(215)) or (inputs(119));
    layer0_outputs(8769) <= not(inputs(22));
    layer0_outputs(8770) <= not((inputs(123)) or (inputs(73)));
    layer0_outputs(8771) <= not((inputs(213)) and (inputs(190)));
    layer0_outputs(8772) <= not((inputs(235)) or (inputs(210)));
    layer0_outputs(8773) <= inputs(121);
    layer0_outputs(8774) <= not(inputs(248)) or (inputs(20));
    layer0_outputs(8775) <= (inputs(141)) and not (inputs(154));
    layer0_outputs(8776) <= (inputs(201)) and not (inputs(196));
    layer0_outputs(8777) <= inputs(231);
    layer0_outputs(8778) <= (inputs(64)) xor (inputs(114));
    layer0_outputs(8779) <= not(inputs(126));
    layer0_outputs(8780) <= not((inputs(49)) and (inputs(118)));
    layer0_outputs(8781) <= (inputs(170)) or (inputs(185));
    layer0_outputs(8782) <= not(inputs(22)) or (inputs(196));
    layer0_outputs(8783) <= not(inputs(151));
    layer0_outputs(8784) <= not(inputs(95)) or (inputs(250));
    layer0_outputs(8785) <= (inputs(18)) and not (inputs(66));
    layer0_outputs(8786) <= inputs(78);
    layer0_outputs(8787) <= (inputs(81)) or (inputs(114));
    layer0_outputs(8788) <= (inputs(100)) or (inputs(189));
    layer0_outputs(8789) <= (inputs(47)) or (inputs(27));
    layer0_outputs(8790) <= (inputs(114)) or (inputs(238));
    layer0_outputs(8791) <= not((inputs(53)) xor (inputs(22)));
    layer0_outputs(8792) <= not(inputs(162));
    layer0_outputs(8793) <= not(inputs(138)) or (inputs(93));
    layer0_outputs(8794) <= not((inputs(83)) or (inputs(219)));
    layer0_outputs(8795) <= not((inputs(210)) xor (inputs(180)));
    layer0_outputs(8796) <= not(inputs(104));
    layer0_outputs(8797) <= (inputs(238)) or (inputs(72));
    layer0_outputs(8798) <= not((inputs(161)) or (inputs(126)));
    layer0_outputs(8799) <= (inputs(146)) or (inputs(68));
    layer0_outputs(8800) <= (inputs(255)) or (inputs(18));
    layer0_outputs(8801) <= (inputs(183)) and not (inputs(173));
    layer0_outputs(8802) <= (inputs(20)) and not (inputs(176));
    layer0_outputs(8803) <= (inputs(68)) and not (inputs(3));
    layer0_outputs(8804) <= (inputs(199)) and (inputs(201));
    layer0_outputs(8805) <= (inputs(129)) or (inputs(34));
    layer0_outputs(8806) <= inputs(237);
    layer0_outputs(8807) <= not((inputs(20)) xor (inputs(81)));
    layer0_outputs(8808) <= inputs(106);
    layer0_outputs(8809) <= not((inputs(62)) xor (inputs(44)));
    layer0_outputs(8810) <= inputs(251);
    layer0_outputs(8811) <= inputs(12);
    layer0_outputs(8812) <= (inputs(194)) and not (inputs(136));
    layer0_outputs(8813) <= not(inputs(217));
    layer0_outputs(8814) <= not(inputs(82));
    layer0_outputs(8815) <= not(inputs(24));
    layer0_outputs(8816) <= not((inputs(14)) and (inputs(117)));
    layer0_outputs(8817) <= not((inputs(231)) xor (inputs(21)));
    layer0_outputs(8818) <= (inputs(30)) or (inputs(69));
    layer0_outputs(8819) <= (inputs(133)) and (inputs(65));
    layer0_outputs(8820) <= inputs(57);
    layer0_outputs(8821) <= not(inputs(11));
    layer0_outputs(8822) <= not((inputs(84)) xor (inputs(218)));
    layer0_outputs(8823) <= inputs(159);
    layer0_outputs(8824) <= '1';
    layer0_outputs(8825) <= not(inputs(133));
    layer0_outputs(8826) <= not((inputs(34)) xor (inputs(125)));
    layer0_outputs(8827) <= (inputs(78)) xor (inputs(6));
    layer0_outputs(8828) <= (inputs(3)) or (inputs(57));
    layer0_outputs(8829) <= not(inputs(164));
    layer0_outputs(8830) <= not((inputs(232)) xor (inputs(246)));
    layer0_outputs(8831) <= not(inputs(54));
    layer0_outputs(8832) <= (inputs(144)) xor (inputs(194));
    layer0_outputs(8833) <= not(inputs(132));
    layer0_outputs(8834) <= not(inputs(133)) or (inputs(29));
    layer0_outputs(8835) <= not((inputs(170)) xor (inputs(238)));
    layer0_outputs(8836) <= not(inputs(171));
    layer0_outputs(8837) <= '1';
    layer0_outputs(8838) <= not((inputs(157)) xor (inputs(119)));
    layer0_outputs(8839) <= inputs(6);
    layer0_outputs(8840) <= inputs(210);
    layer0_outputs(8841) <= inputs(93);
    layer0_outputs(8842) <= not(inputs(171)) or (inputs(31));
    layer0_outputs(8843) <= (inputs(106)) and not (inputs(153));
    layer0_outputs(8844) <= not(inputs(28)) or (inputs(125));
    layer0_outputs(8845) <= '0';
    layer0_outputs(8846) <= not((inputs(241)) xor (inputs(156)));
    layer0_outputs(8847) <= not(inputs(169));
    layer0_outputs(8848) <= not((inputs(31)) or (inputs(108)));
    layer0_outputs(8849) <= inputs(9);
    layer0_outputs(8850) <= '1';
    layer0_outputs(8851) <= not(inputs(201));
    layer0_outputs(8852) <= not(inputs(210)) or (inputs(146));
    layer0_outputs(8853) <= (inputs(17)) and (inputs(227));
    layer0_outputs(8854) <= not((inputs(174)) or (inputs(193)));
    layer0_outputs(8855) <= not(inputs(233)) or (inputs(127));
    layer0_outputs(8856) <= not(inputs(195)) or (inputs(113));
    layer0_outputs(8857) <= inputs(43);
    layer0_outputs(8858) <= (inputs(106)) and not (inputs(184));
    layer0_outputs(8859) <= inputs(122);
    layer0_outputs(8860) <= (inputs(158)) xor (inputs(185));
    layer0_outputs(8861) <= (inputs(205)) and not (inputs(243));
    layer0_outputs(8862) <= not((inputs(115)) xor (inputs(128)));
    layer0_outputs(8863) <= not((inputs(192)) or (inputs(133)));
    layer0_outputs(8864) <= (inputs(229)) and not (inputs(223));
    layer0_outputs(8865) <= inputs(249);
    layer0_outputs(8866) <= not(inputs(176)) or (inputs(36));
    layer0_outputs(8867) <= (inputs(217)) or (inputs(67));
    layer0_outputs(8868) <= (inputs(98)) and not (inputs(110));
    layer0_outputs(8869) <= inputs(242);
    layer0_outputs(8870) <= not((inputs(136)) or (inputs(225)));
    layer0_outputs(8871) <= not((inputs(9)) xor (inputs(207)));
    layer0_outputs(8872) <= (inputs(50)) and (inputs(62));
    layer0_outputs(8873) <= inputs(202);
    layer0_outputs(8874) <= (inputs(75)) and (inputs(106));
    layer0_outputs(8875) <= inputs(76);
    layer0_outputs(8876) <= (inputs(183)) and not (inputs(83));
    layer0_outputs(8877) <= not((inputs(197)) xor (inputs(10)));
    layer0_outputs(8878) <= not((inputs(214)) or (inputs(181)));
    layer0_outputs(8879) <= not(inputs(185));
    layer0_outputs(8880) <= (inputs(241)) and not (inputs(214));
    layer0_outputs(8881) <= not(inputs(193));
    layer0_outputs(8882) <= not((inputs(242)) and (inputs(55)));
    layer0_outputs(8883) <= (inputs(89)) or (inputs(4));
    layer0_outputs(8884) <= not(inputs(210));
    layer0_outputs(8885) <= not(inputs(13)) or (inputs(90));
    layer0_outputs(8886) <= not(inputs(47));
    layer0_outputs(8887) <= not((inputs(37)) xor (inputs(43)));
    layer0_outputs(8888) <= not(inputs(233));
    layer0_outputs(8889) <= not((inputs(118)) xor (inputs(116)));
    layer0_outputs(8890) <= (inputs(233)) and not (inputs(150));
    layer0_outputs(8891) <= '1';
    layer0_outputs(8892) <= '1';
    layer0_outputs(8893) <= not(inputs(222));
    layer0_outputs(8894) <= not(inputs(33)) or (inputs(65));
    layer0_outputs(8895) <= inputs(165);
    layer0_outputs(8896) <= not((inputs(139)) xor (inputs(101)));
    layer0_outputs(8897) <= (inputs(4)) or (inputs(64));
    layer0_outputs(8898) <= not(inputs(100));
    layer0_outputs(8899) <= (inputs(149)) and not (inputs(38));
    layer0_outputs(8900) <= inputs(150);
    layer0_outputs(8901) <= not(inputs(78));
    layer0_outputs(8902) <= inputs(107);
    layer0_outputs(8903) <= '0';
    layer0_outputs(8904) <= (inputs(45)) and not (inputs(137));
    layer0_outputs(8905) <= (inputs(219)) and (inputs(182));
    layer0_outputs(8906) <= not(inputs(174)) or (inputs(153));
    layer0_outputs(8907) <= not((inputs(253)) or (inputs(134)));
    layer0_outputs(8908) <= not((inputs(247)) and (inputs(227)));
    layer0_outputs(8909) <= not(inputs(24));
    layer0_outputs(8910) <= '1';
    layer0_outputs(8911) <= (inputs(159)) and not (inputs(215));
    layer0_outputs(8912) <= not((inputs(249)) or (inputs(254)));
    layer0_outputs(8913) <= not(inputs(45));
    layer0_outputs(8914) <= '0';
    layer0_outputs(8915) <= not((inputs(232)) or (inputs(190)));
    layer0_outputs(8916) <= not(inputs(181));
    layer0_outputs(8917) <= inputs(119);
    layer0_outputs(8918) <= not(inputs(197));
    layer0_outputs(8919) <= '1';
    layer0_outputs(8920) <= (inputs(146)) or (inputs(50));
    layer0_outputs(8921) <= not(inputs(37));
    layer0_outputs(8922) <= inputs(140);
    layer0_outputs(8923) <= not(inputs(193)) or (inputs(39));
    layer0_outputs(8924) <= not(inputs(28)) or (inputs(253));
    layer0_outputs(8925) <= (inputs(154)) and not (inputs(3));
    layer0_outputs(8926) <= (inputs(121)) and not (inputs(93));
    layer0_outputs(8927) <= not(inputs(229));
    layer0_outputs(8928) <= inputs(58);
    layer0_outputs(8929) <= not((inputs(39)) or (inputs(47)));
    layer0_outputs(8930) <= (inputs(254)) and not (inputs(220));
    layer0_outputs(8931) <= not(inputs(136));
    layer0_outputs(8932) <= (inputs(148)) or (inputs(87));
    layer0_outputs(8933) <= not(inputs(123)) or (inputs(59));
    layer0_outputs(8934) <= not(inputs(207));
    layer0_outputs(8935) <= inputs(25);
    layer0_outputs(8936) <= inputs(100);
    layer0_outputs(8937) <= not((inputs(159)) or (inputs(32)));
    layer0_outputs(8938) <= (inputs(109)) and not (inputs(239));
    layer0_outputs(8939) <= not((inputs(53)) and (inputs(59)));
    layer0_outputs(8940) <= (inputs(197)) and not (inputs(190));
    layer0_outputs(8941) <= not(inputs(35));
    layer0_outputs(8942) <= inputs(98);
    layer0_outputs(8943) <= inputs(219);
    layer0_outputs(8944) <= inputs(114);
    layer0_outputs(8945) <= not(inputs(252));
    layer0_outputs(8946) <= inputs(245);
    layer0_outputs(8947) <= not(inputs(88)) or (inputs(34));
    layer0_outputs(8948) <= not(inputs(24)) or (inputs(97));
    layer0_outputs(8949) <= not(inputs(129));
    layer0_outputs(8950) <= inputs(250);
    layer0_outputs(8951) <= not((inputs(145)) xor (inputs(132)));
    layer0_outputs(8952) <= inputs(247);
    layer0_outputs(8953) <= not((inputs(85)) and (inputs(85)));
    layer0_outputs(8954) <= (inputs(85)) and (inputs(84));
    layer0_outputs(8955) <= not(inputs(49));
    layer0_outputs(8956) <= (inputs(253)) or (inputs(254));
    layer0_outputs(8957) <= inputs(115);
    layer0_outputs(8958) <= (inputs(91)) and not (inputs(57));
    layer0_outputs(8959) <= (inputs(191)) xor (inputs(108));
    layer0_outputs(8960) <= '1';
    layer0_outputs(8961) <= inputs(58);
    layer0_outputs(8962) <= not(inputs(93));
    layer0_outputs(8963) <= inputs(247);
    layer0_outputs(8964) <= not((inputs(170)) and (inputs(76)));
    layer0_outputs(8965) <= not(inputs(186));
    layer0_outputs(8966) <= not((inputs(225)) or (inputs(63)));
    layer0_outputs(8967) <= inputs(90);
    layer0_outputs(8968) <= inputs(73);
    layer0_outputs(8969) <= (inputs(70)) and not (inputs(191));
    layer0_outputs(8970) <= (inputs(78)) or (inputs(45));
    layer0_outputs(8971) <= not(inputs(212));
    layer0_outputs(8972) <= '0';
    layer0_outputs(8973) <= not(inputs(171));
    layer0_outputs(8974) <= (inputs(79)) xor (inputs(222));
    layer0_outputs(8975) <= not(inputs(61));
    layer0_outputs(8976) <= not(inputs(146));
    layer0_outputs(8977) <= not(inputs(160));
    layer0_outputs(8978) <= inputs(167);
    layer0_outputs(8979) <= not(inputs(29));
    layer0_outputs(8980) <= not(inputs(120));
    layer0_outputs(8981) <= (inputs(161)) or (inputs(222));
    layer0_outputs(8982) <= not((inputs(88)) xor (inputs(93)));
    layer0_outputs(8983) <= not(inputs(147));
    layer0_outputs(8984) <= not(inputs(102));
    layer0_outputs(8985) <= (inputs(191)) and (inputs(32));
    layer0_outputs(8986) <= '1';
    layer0_outputs(8987) <= (inputs(186)) xor (inputs(177));
    layer0_outputs(8988) <= not((inputs(164)) xor (inputs(176)));
    layer0_outputs(8989) <= inputs(123);
    layer0_outputs(8990) <= (inputs(22)) and not (inputs(115));
    layer0_outputs(8991) <= not(inputs(146)) or (inputs(220));
    layer0_outputs(8992) <= inputs(28);
    layer0_outputs(8993) <= '0';
    layer0_outputs(8994) <= not(inputs(11)) or (inputs(18));
    layer0_outputs(8995) <= inputs(117);
    layer0_outputs(8996) <= not((inputs(122)) xor (inputs(110)));
    layer0_outputs(8997) <= (inputs(85)) or (inputs(100));
    layer0_outputs(8998) <= (inputs(42)) and (inputs(66));
    layer0_outputs(8999) <= (inputs(91)) xor (inputs(65));
    layer0_outputs(9000) <= (inputs(47)) xor (inputs(105));
    layer0_outputs(9001) <= inputs(231);
    layer0_outputs(9002) <= (inputs(13)) or (inputs(30));
    layer0_outputs(9003) <= (inputs(49)) xor (inputs(123));
    layer0_outputs(9004) <= inputs(121);
    layer0_outputs(9005) <= (inputs(236)) xor (inputs(207));
    layer0_outputs(9006) <= not((inputs(42)) or (inputs(79)));
    layer0_outputs(9007) <= not(inputs(243)) or (inputs(135));
    layer0_outputs(9008) <= not((inputs(78)) and (inputs(88)));
    layer0_outputs(9009) <= inputs(73);
    layer0_outputs(9010) <= (inputs(158)) or (inputs(146));
    layer0_outputs(9011) <= not((inputs(2)) or (inputs(183)));
    layer0_outputs(9012) <= (inputs(203)) and (inputs(0));
    layer0_outputs(9013) <= not(inputs(16));
    layer0_outputs(9014) <= (inputs(174)) or (inputs(160));
    layer0_outputs(9015) <= inputs(155);
    layer0_outputs(9016) <= (inputs(41)) and not (inputs(238));
    layer0_outputs(9017) <= (inputs(211)) and not (inputs(88));
    layer0_outputs(9018) <= not(inputs(121));
    layer0_outputs(9019) <= (inputs(64)) xor (inputs(5));
    layer0_outputs(9020) <= (inputs(147)) or (inputs(124));
    layer0_outputs(9021) <= (inputs(228)) and not (inputs(30));
    layer0_outputs(9022) <= not((inputs(42)) or (inputs(6)));
    layer0_outputs(9023) <= (inputs(76)) and not (inputs(195));
    layer0_outputs(9024) <= inputs(176);
    layer0_outputs(9025) <= (inputs(131)) or (inputs(53));
    layer0_outputs(9026) <= not(inputs(110));
    layer0_outputs(9027) <= inputs(184);
    layer0_outputs(9028) <= (inputs(128)) xor (inputs(31));
    layer0_outputs(9029) <= '1';
    layer0_outputs(9030) <= not(inputs(211)) or (inputs(95));
    layer0_outputs(9031) <= not(inputs(166));
    layer0_outputs(9032) <= not((inputs(48)) or (inputs(106)));
    layer0_outputs(9033) <= (inputs(159)) and not (inputs(145));
    layer0_outputs(9034) <= not((inputs(178)) or (inputs(125)));
    layer0_outputs(9035) <= not(inputs(102));
    layer0_outputs(9036) <= '1';
    layer0_outputs(9037) <= inputs(74);
    layer0_outputs(9038) <= (inputs(37)) xor (inputs(252));
    layer0_outputs(9039) <= (inputs(26)) or (inputs(3));
    layer0_outputs(9040) <= not(inputs(232));
    layer0_outputs(9041) <= not((inputs(159)) and (inputs(40)));
    layer0_outputs(9042) <= inputs(92);
    layer0_outputs(9043) <= inputs(193);
    layer0_outputs(9044) <= not(inputs(130));
    layer0_outputs(9045) <= (inputs(141)) and not (inputs(19));
    layer0_outputs(9046) <= inputs(193);
    layer0_outputs(9047) <= (inputs(178)) xor (inputs(219));
    layer0_outputs(9048) <= not(inputs(13)) or (inputs(245));
    layer0_outputs(9049) <= (inputs(21)) and not (inputs(207));
    layer0_outputs(9050) <= inputs(117);
    layer0_outputs(9051) <= not((inputs(108)) or (inputs(130)));
    layer0_outputs(9052) <= (inputs(131)) and not (inputs(241));
    layer0_outputs(9053) <= inputs(97);
    layer0_outputs(9054) <= not(inputs(146));
    layer0_outputs(9055) <= not(inputs(148));
    layer0_outputs(9056) <= (inputs(229)) and not (inputs(222));
    layer0_outputs(9057) <= not(inputs(160));
    layer0_outputs(9058) <= not((inputs(137)) or (inputs(59)));
    layer0_outputs(9059) <= (inputs(141)) and (inputs(146));
    layer0_outputs(9060) <= inputs(68);
    layer0_outputs(9061) <= not((inputs(153)) xor (inputs(94)));
    layer0_outputs(9062) <= inputs(158);
    layer0_outputs(9063) <= (inputs(176)) or (inputs(50));
    layer0_outputs(9064) <= not((inputs(125)) or (inputs(49)));
    layer0_outputs(9065) <= '0';
    layer0_outputs(9066) <= not((inputs(229)) and (inputs(232)));
    layer0_outputs(9067) <= not((inputs(170)) or (inputs(236)));
    layer0_outputs(9068) <= (inputs(88)) xor (inputs(49));
    layer0_outputs(9069) <= (inputs(46)) or (inputs(66));
    layer0_outputs(9070) <= not(inputs(23)) or (inputs(240));
    layer0_outputs(9071) <= inputs(203);
    layer0_outputs(9072) <= not(inputs(223)) or (inputs(36));
    layer0_outputs(9073) <= not(inputs(70));
    layer0_outputs(9074) <= not(inputs(177)) or (inputs(42));
    layer0_outputs(9075) <= not((inputs(82)) or (inputs(54)));
    layer0_outputs(9076) <= not((inputs(49)) xor (inputs(6)));
    layer0_outputs(9077) <= (inputs(134)) and not (inputs(237));
    layer0_outputs(9078) <= '1';
    layer0_outputs(9079) <= not(inputs(212)) or (inputs(98));
    layer0_outputs(9080) <= not(inputs(112)) or (inputs(31));
    layer0_outputs(9081) <= (inputs(59)) and (inputs(62));
    layer0_outputs(9082) <= not((inputs(41)) or (inputs(190)));
    layer0_outputs(9083) <= not((inputs(175)) or (inputs(177)));
    layer0_outputs(9084) <= not((inputs(20)) or (inputs(89)));
    layer0_outputs(9085) <= (inputs(206)) and not (inputs(131));
    layer0_outputs(9086) <= inputs(127);
    layer0_outputs(9087) <= '0';
    layer0_outputs(9088) <= not(inputs(71));
    layer0_outputs(9089) <= inputs(248);
    layer0_outputs(9090) <= not(inputs(21));
    layer0_outputs(9091) <= not(inputs(174));
    layer0_outputs(9092) <= (inputs(0)) xor (inputs(62));
    layer0_outputs(9093) <= inputs(179);
    layer0_outputs(9094) <= (inputs(188)) xor (inputs(242));
    layer0_outputs(9095) <= (inputs(11)) and not (inputs(201));
    layer0_outputs(9096) <= not((inputs(201)) or (inputs(34)));
    layer0_outputs(9097) <= inputs(169);
    layer0_outputs(9098) <= (inputs(226)) and (inputs(44));
    layer0_outputs(9099) <= not((inputs(249)) xor (inputs(99)));
    layer0_outputs(9100) <= not(inputs(163)) or (inputs(31));
    layer0_outputs(9101) <= (inputs(241)) or (inputs(66));
    layer0_outputs(9102) <= not(inputs(37)) or (inputs(153));
    layer0_outputs(9103) <= not((inputs(62)) or (inputs(32)));
    layer0_outputs(9104) <= not(inputs(19));
    layer0_outputs(9105) <= not(inputs(121));
    layer0_outputs(9106) <= (inputs(126)) and not (inputs(154));
    layer0_outputs(9107) <= inputs(42);
    layer0_outputs(9108) <= not(inputs(105));
    layer0_outputs(9109) <= not(inputs(233)) or (inputs(105));
    layer0_outputs(9110) <= not(inputs(63)) or (inputs(16));
    layer0_outputs(9111) <= (inputs(180)) and not (inputs(6));
    layer0_outputs(9112) <= inputs(128);
    layer0_outputs(9113) <= (inputs(158)) or (inputs(176));
    layer0_outputs(9114) <= (inputs(108)) and (inputs(159));
    layer0_outputs(9115) <= not(inputs(81));
    layer0_outputs(9116) <= inputs(117);
    layer0_outputs(9117) <= (inputs(217)) xor (inputs(192));
    layer0_outputs(9118) <= not(inputs(118));
    layer0_outputs(9119) <= (inputs(22)) and not (inputs(73));
    layer0_outputs(9120) <= (inputs(40)) and not (inputs(217));
    layer0_outputs(9121) <= not(inputs(73)) or (inputs(210));
    layer0_outputs(9122) <= (inputs(35)) and not (inputs(125));
    layer0_outputs(9123) <= not((inputs(145)) or (inputs(30)));
    layer0_outputs(9124) <= (inputs(247)) or (inputs(228));
    layer0_outputs(9125) <= inputs(76);
    layer0_outputs(9126) <= not(inputs(127));
    layer0_outputs(9127) <= not(inputs(190));
    layer0_outputs(9128) <= inputs(230);
    layer0_outputs(9129) <= not(inputs(13)) or (inputs(80));
    layer0_outputs(9130) <= not(inputs(171));
    layer0_outputs(9131) <= not((inputs(47)) or (inputs(32)));
    layer0_outputs(9132) <= not((inputs(211)) xor (inputs(14)));
    layer0_outputs(9133) <= not((inputs(4)) or (inputs(35)));
    layer0_outputs(9134) <= not(inputs(234));
    layer0_outputs(9135) <= (inputs(39)) and not (inputs(132));
    layer0_outputs(9136) <= (inputs(107)) or (inputs(30));
    layer0_outputs(9137) <= inputs(147);
    layer0_outputs(9138) <= not(inputs(84));
    layer0_outputs(9139) <= '1';
    layer0_outputs(9140) <= not(inputs(82));
    layer0_outputs(9141) <= not((inputs(187)) xor (inputs(251)));
    layer0_outputs(9142) <= (inputs(171)) or (inputs(97));
    layer0_outputs(9143) <= inputs(133);
    layer0_outputs(9144) <= not((inputs(132)) or (inputs(61)));
    layer0_outputs(9145) <= '0';
    layer0_outputs(9146) <= not(inputs(42)) or (inputs(135));
    layer0_outputs(9147) <= (inputs(65)) and (inputs(70));
    layer0_outputs(9148) <= inputs(247);
    layer0_outputs(9149) <= (inputs(36)) xor (inputs(254));
    layer0_outputs(9150) <= (inputs(195)) and not (inputs(85));
    layer0_outputs(9151) <= '0';
    layer0_outputs(9152) <= inputs(83);
    layer0_outputs(9153) <= not(inputs(138)) or (inputs(60));
    layer0_outputs(9154) <= not((inputs(199)) or (inputs(59)));
    layer0_outputs(9155) <= (inputs(216)) and (inputs(209));
    layer0_outputs(9156) <= not((inputs(113)) xor (inputs(138)));
    layer0_outputs(9157) <= not((inputs(155)) or (inputs(35)));
    layer0_outputs(9158) <= inputs(244);
    layer0_outputs(9159) <= inputs(153);
    layer0_outputs(9160) <= not((inputs(98)) or (inputs(37)));
    layer0_outputs(9161) <= (inputs(132)) and not (inputs(252));
    layer0_outputs(9162) <= (inputs(152)) or (inputs(255));
    layer0_outputs(9163) <= not(inputs(101));
    layer0_outputs(9164) <= inputs(47);
    layer0_outputs(9165) <= inputs(128);
    layer0_outputs(9166) <= (inputs(162)) and not (inputs(243));
    layer0_outputs(9167) <= (inputs(239)) and not (inputs(214));
    layer0_outputs(9168) <= (inputs(83)) or (inputs(201));
    layer0_outputs(9169) <= not(inputs(228));
    layer0_outputs(9170) <= inputs(57);
    layer0_outputs(9171) <= not(inputs(78));
    layer0_outputs(9172) <= '1';
    layer0_outputs(9173) <= not((inputs(145)) or (inputs(90)));
    layer0_outputs(9174) <= not(inputs(121)) or (inputs(229));
    layer0_outputs(9175) <= not(inputs(107));
    layer0_outputs(9176) <= not(inputs(104));
    layer0_outputs(9177) <= (inputs(222)) and not (inputs(210));
    layer0_outputs(9178) <= (inputs(43)) or (inputs(75));
    layer0_outputs(9179) <= not(inputs(229));
    layer0_outputs(9180) <= (inputs(82)) and not (inputs(229));
    layer0_outputs(9181) <= inputs(149);
    layer0_outputs(9182) <= not(inputs(212));
    layer0_outputs(9183) <= not((inputs(154)) xor (inputs(236)));
    layer0_outputs(9184) <= '1';
    layer0_outputs(9185) <= not(inputs(73)) or (inputs(34));
    layer0_outputs(9186) <= not((inputs(46)) or (inputs(101)));
    layer0_outputs(9187) <= not(inputs(44));
    layer0_outputs(9188) <= not(inputs(209)) or (inputs(15));
    layer0_outputs(9189) <= (inputs(157)) or (inputs(172));
    layer0_outputs(9190) <= (inputs(226)) and (inputs(200));
    layer0_outputs(9191) <= not((inputs(78)) and (inputs(63)));
    layer0_outputs(9192) <= not(inputs(85));
    layer0_outputs(9193) <= '1';
    layer0_outputs(9194) <= not((inputs(142)) or (inputs(20)));
    layer0_outputs(9195) <= not(inputs(101));
    layer0_outputs(9196) <= not(inputs(169)) or (inputs(82));
    layer0_outputs(9197) <= inputs(167);
    layer0_outputs(9198) <= not(inputs(115)) or (inputs(192));
    layer0_outputs(9199) <= not(inputs(120)) or (inputs(55));
    layer0_outputs(9200) <= not((inputs(241)) xor (inputs(44)));
    layer0_outputs(9201) <= not((inputs(116)) or (inputs(87)));
    layer0_outputs(9202) <= not((inputs(238)) or (inputs(120)));
    layer0_outputs(9203) <= '0';
    layer0_outputs(9204) <= not((inputs(206)) xor (inputs(20)));
    layer0_outputs(9205) <= inputs(89);
    layer0_outputs(9206) <= not(inputs(145)) or (inputs(66));
    layer0_outputs(9207) <= not((inputs(29)) or (inputs(53)));
    layer0_outputs(9208) <= inputs(235);
    layer0_outputs(9209) <= inputs(121);
    layer0_outputs(9210) <= not(inputs(101)) or (inputs(91));
    layer0_outputs(9211) <= not(inputs(149));
    layer0_outputs(9212) <= not(inputs(202));
    layer0_outputs(9213) <= not((inputs(222)) xor (inputs(211)));
    layer0_outputs(9214) <= not((inputs(186)) xor (inputs(187)));
    layer0_outputs(9215) <= not((inputs(79)) or (inputs(25)));
    layer0_outputs(9216) <= (inputs(99)) and not (inputs(195));
    layer0_outputs(9217) <= (inputs(210)) and not (inputs(64));
    layer0_outputs(9218) <= inputs(145);
    layer0_outputs(9219) <= (inputs(101)) xor (inputs(109));
    layer0_outputs(9220) <= (inputs(90)) or (inputs(181));
    layer0_outputs(9221) <= not(inputs(90));
    layer0_outputs(9222) <= (inputs(37)) or (inputs(250));
    layer0_outputs(9223) <= not((inputs(250)) or (inputs(223)));
    layer0_outputs(9224) <= (inputs(225)) xor (inputs(189));
    layer0_outputs(9225) <= (inputs(234)) and not (inputs(175));
    layer0_outputs(9226) <= not(inputs(31));
    layer0_outputs(9227) <= not(inputs(193));
    layer0_outputs(9228) <= not((inputs(34)) or (inputs(246)));
    layer0_outputs(9229) <= inputs(156);
    layer0_outputs(9230) <= not((inputs(6)) or (inputs(131)));
    layer0_outputs(9231) <= not(inputs(156));
    layer0_outputs(9232) <= not((inputs(144)) and (inputs(101)));
    layer0_outputs(9233) <= inputs(82);
    layer0_outputs(9234) <= '0';
    layer0_outputs(9235) <= (inputs(242)) or (inputs(246));
    layer0_outputs(9236) <= (inputs(66)) and not (inputs(249));
    layer0_outputs(9237) <= not((inputs(128)) xor (inputs(130)));
    layer0_outputs(9238) <= not((inputs(243)) or (inputs(46)));
    layer0_outputs(9239) <= '0';
    layer0_outputs(9240) <= inputs(121);
    layer0_outputs(9241) <= (inputs(196)) xor (inputs(148));
    layer0_outputs(9242) <= not(inputs(37));
    layer0_outputs(9243) <= inputs(229);
    layer0_outputs(9244) <= (inputs(167)) and not (inputs(88));
    layer0_outputs(9245) <= not((inputs(191)) and (inputs(31)));
    layer0_outputs(9246) <= inputs(171);
    layer0_outputs(9247) <= (inputs(205)) or (inputs(211));
    layer0_outputs(9248) <= inputs(18);
    layer0_outputs(9249) <= not(inputs(219)) or (inputs(29));
    layer0_outputs(9250) <= not(inputs(126));
    layer0_outputs(9251) <= inputs(115);
    layer0_outputs(9252) <= '0';
    layer0_outputs(9253) <= not(inputs(203));
    layer0_outputs(9254) <= (inputs(222)) or (inputs(233));
    layer0_outputs(9255) <= inputs(163);
    layer0_outputs(9256) <= not(inputs(249)) or (inputs(0));
    layer0_outputs(9257) <= not(inputs(196));
    layer0_outputs(9258) <= not(inputs(50));
    layer0_outputs(9259) <= (inputs(19)) or (inputs(251));
    layer0_outputs(9260) <= inputs(45);
    layer0_outputs(9261) <= (inputs(103)) and not (inputs(2));
    layer0_outputs(9262) <= not(inputs(28));
    layer0_outputs(9263) <= '0';
    layer0_outputs(9264) <= (inputs(216)) and not (inputs(169));
    layer0_outputs(9265) <= not(inputs(93));
    layer0_outputs(9266) <= not(inputs(246));
    layer0_outputs(9267) <= not(inputs(51));
    layer0_outputs(9268) <= (inputs(80)) and not (inputs(99));
    layer0_outputs(9269) <= not(inputs(50));
    layer0_outputs(9270) <= (inputs(176)) and not (inputs(140));
    layer0_outputs(9271) <= inputs(87);
    layer0_outputs(9272) <= inputs(67);
    layer0_outputs(9273) <= (inputs(16)) xor (inputs(204));
    layer0_outputs(9274) <= not((inputs(142)) or (inputs(215)));
    layer0_outputs(9275) <= '1';
    layer0_outputs(9276) <= (inputs(230)) and not (inputs(28));
    layer0_outputs(9277) <= (inputs(100)) xor (inputs(189));
    layer0_outputs(9278) <= not((inputs(75)) and (inputs(9)));
    layer0_outputs(9279) <= not((inputs(16)) xor (inputs(243)));
    layer0_outputs(9280) <= not((inputs(196)) or (inputs(155)));
    layer0_outputs(9281) <= not(inputs(151));
    layer0_outputs(9282) <= (inputs(172)) and not (inputs(49));
    layer0_outputs(9283) <= not(inputs(134));
    layer0_outputs(9284) <= (inputs(50)) or (inputs(181));
    layer0_outputs(9285) <= not((inputs(223)) or (inputs(214)));
    layer0_outputs(9286) <= not((inputs(50)) or (inputs(196)));
    layer0_outputs(9287) <= not((inputs(146)) xor (inputs(248)));
    layer0_outputs(9288) <= not((inputs(112)) xor (inputs(85)));
    layer0_outputs(9289) <= inputs(165);
    layer0_outputs(9290) <= (inputs(5)) xor (inputs(34));
    layer0_outputs(9291) <= not(inputs(150));
    layer0_outputs(9292) <= inputs(94);
    layer0_outputs(9293) <= inputs(133);
    layer0_outputs(9294) <= inputs(145);
    layer0_outputs(9295) <= not((inputs(135)) or (inputs(151)));
    layer0_outputs(9296) <= inputs(108);
    layer0_outputs(9297) <= (inputs(107)) and not (inputs(129));
    layer0_outputs(9298) <= (inputs(247)) xor (inputs(114));
    layer0_outputs(9299) <= (inputs(165)) and not (inputs(53));
    layer0_outputs(9300) <= '1';
    layer0_outputs(9301) <= (inputs(166)) or (inputs(185));
    layer0_outputs(9302) <= not(inputs(221));
    layer0_outputs(9303) <= not((inputs(174)) xor (inputs(175)));
    layer0_outputs(9304) <= inputs(108);
    layer0_outputs(9305) <= not(inputs(204));
    layer0_outputs(9306) <= (inputs(79)) xor (inputs(2));
    layer0_outputs(9307) <= not(inputs(60));
    layer0_outputs(9308) <= (inputs(34)) xor (inputs(124));
    layer0_outputs(9309) <= not(inputs(24)) or (inputs(235));
    layer0_outputs(9310) <= inputs(8);
    layer0_outputs(9311) <= inputs(244);
    layer0_outputs(9312) <= (inputs(217)) xor (inputs(101));
    layer0_outputs(9313) <= inputs(226);
    layer0_outputs(9314) <= not(inputs(171));
    layer0_outputs(9315) <= inputs(113);
    layer0_outputs(9316) <= not((inputs(231)) xor (inputs(236)));
    layer0_outputs(9317) <= not(inputs(76)) or (inputs(146));
    layer0_outputs(9318) <= not((inputs(12)) or (inputs(22)));
    layer0_outputs(9319) <= inputs(178);
    layer0_outputs(9320) <= (inputs(75)) or (inputs(162));
    layer0_outputs(9321) <= (inputs(211)) and not (inputs(164));
    layer0_outputs(9322) <= inputs(154);
    layer0_outputs(9323) <= inputs(89);
    layer0_outputs(9324) <= not(inputs(29));
    layer0_outputs(9325) <= (inputs(176)) and not (inputs(78));
    layer0_outputs(9326) <= not(inputs(66));
    layer0_outputs(9327) <= (inputs(140)) and not (inputs(197));
    layer0_outputs(9328) <= not(inputs(199));
    layer0_outputs(9329) <= (inputs(163)) and not (inputs(61));
    layer0_outputs(9330) <= '1';
    layer0_outputs(9331) <= not((inputs(90)) or (inputs(173)));
    layer0_outputs(9332) <= inputs(102);
    layer0_outputs(9333) <= not((inputs(155)) or (inputs(238)));
    layer0_outputs(9334) <= (inputs(9)) and not (inputs(240));
    layer0_outputs(9335) <= inputs(125);
    layer0_outputs(9336) <= not(inputs(173));
    layer0_outputs(9337) <= not((inputs(249)) or (inputs(171)));
    layer0_outputs(9338) <= inputs(108);
    layer0_outputs(9339) <= not(inputs(244)) or (inputs(219));
    layer0_outputs(9340) <= inputs(95);
    layer0_outputs(9341) <= not((inputs(19)) xor (inputs(222)));
    layer0_outputs(9342) <= not(inputs(208)) or (inputs(67));
    layer0_outputs(9343) <= not((inputs(101)) or (inputs(172)));
    layer0_outputs(9344) <= inputs(46);
    layer0_outputs(9345) <= not(inputs(95));
    layer0_outputs(9346) <= (inputs(17)) and not (inputs(118));
    layer0_outputs(9347) <= not(inputs(126));
    layer0_outputs(9348) <= not(inputs(153));
    layer0_outputs(9349) <= inputs(226);
    layer0_outputs(9350) <= not(inputs(252)) or (inputs(189));
    layer0_outputs(9351) <= (inputs(139)) or (inputs(144));
    layer0_outputs(9352) <= inputs(241);
    layer0_outputs(9353) <= not((inputs(108)) or (inputs(114)));
    layer0_outputs(9354) <= '0';
    layer0_outputs(9355) <= not(inputs(39)) or (inputs(63));
    layer0_outputs(9356) <= not(inputs(66));
    layer0_outputs(9357) <= not(inputs(92));
    layer0_outputs(9358) <= (inputs(231)) and not (inputs(125));
    layer0_outputs(9359) <= not((inputs(175)) or (inputs(196)));
    layer0_outputs(9360) <= (inputs(19)) and not (inputs(96));
    layer0_outputs(9361) <= '1';
    layer0_outputs(9362) <= (inputs(4)) or (inputs(103));
    layer0_outputs(9363) <= inputs(100);
    layer0_outputs(9364) <= not((inputs(40)) xor (inputs(175)));
    layer0_outputs(9365) <= not((inputs(191)) xor (inputs(236)));
    layer0_outputs(9366) <= not(inputs(106));
    layer0_outputs(9367) <= not((inputs(15)) or (inputs(201)));
    layer0_outputs(9368) <= not(inputs(136));
    layer0_outputs(9369) <= not(inputs(223));
    layer0_outputs(9370) <= (inputs(14)) and not (inputs(76));
    layer0_outputs(9371) <= inputs(176);
    layer0_outputs(9372) <= (inputs(42)) and (inputs(108));
    layer0_outputs(9373) <= (inputs(183)) and (inputs(36));
    layer0_outputs(9374) <= (inputs(73)) and not (inputs(64));
    layer0_outputs(9375) <= not((inputs(40)) xor (inputs(60)));
    layer0_outputs(9376) <= (inputs(2)) or (inputs(22));
    layer0_outputs(9377) <= (inputs(39)) and (inputs(237));
    layer0_outputs(9378) <= (inputs(30)) xor (inputs(208));
    layer0_outputs(9379) <= not((inputs(149)) xor (inputs(176)));
    layer0_outputs(9380) <= inputs(203);
    layer0_outputs(9381) <= not((inputs(177)) xor (inputs(225)));
    layer0_outputs(9382) <= (inputs(78)) xor (inputs(133));
    layer0_outputs(9383) <= (inputs(91)) and not (inputs(226));
    layer0_outputs(9384) <= (inputs(159)) and not (inputs(190));
    layer0_outputs(9385) <= not((inputs(35)) xor (inputs(62)));
    layer0_outputs(9386) <= not(inputs(134));
    layer0_outputs(9387) <= (inputs(106)) and not (inputs(89));
    layer0_outputs(9388) <= inputs(150);
    layer0_outputs(9389) <= (inputs(196)) and not (inputs(3));
    layer0_outputs(9390) <= not(inputs(70));
    layer0_outputs(9391) <= not(inputs(127));
    layer0_outputs(9392) <= inputs(148);
    layer0_outputs(9393) <= not((inputs(55)) xor (inputs(49)));
    layer0_outputs(9394) <= (inputs(248)) and not (inputs(232));
    layer0_outputs(9395) <= not(inputs(117));
    layer0_outputs(9396) <= not(inputs(188));
    layer0_outputs(9397) <= not((inputs(217)) or (inputs(187)));
    layer0_outputs(9398) <= (inputs(85)) and not (inputs(26));
    layer0_outputs(9399) <= not((inputs(31)) or (inputs(3)));
    layer0_outputs(9400) <= not(inputs(23)) or (inputs(191));
    layer0_outputs(9401) <= not(inputs(246)) or (inputs(240));
    layer0_outputs(9402) <= (inputs(61)) or (inputs(43));
    layer0_outputs(9403) <= (inputs(110)) xor (inputs(163));
    layer0_outputs(9404) <= (inputs(120)) or (inputs(142));
    layer0_outputs(9405) <= '1';
    layer0_outputs(9406) <= (inputs(173)) and not (inputs(65));
    layer0_outputs(9407) <= not(inputs(81)) or (inputs(189));
    layer0_outputs(9408) <= inputs(125);
    layer0_outputs(9409) <= not((inputs(217)) or (inputs(132)));
    layer0_outputs(9410) <= (inputs(117)) and not (inputs(224));
    layer0_outputs(9411) <= not(inputs(146));
    layer0_outputs(9412) <= not(inputs(59));
    layer0_outputs(9413) <= not(inputs(108)) or (inputs(133));
    layer0_outputs(9414) <= not((inputs(178)) and (inputs(20)));
    layer0_outputs(9415) <= inputs(162);
    layer0_outputs(9416) <= not((inputs(248)) and (inputs(138)));
    layer0_outputs(9417) <= not(inputs(125));
    layer0_outputs(9418) <= not(inputs(211));
    layer0_outputs(9419) <= not(inputs(93));
    layer0_outputs(9420) <= (inputs(75)) and not (inputs(220));
    layer0_outputs(9421) <= inputs(75);
    layer0_outputs(9422) <= not((inputs(122)) xor (inputs(92)));
    layer0_outputs(9423) <= not(inputs(23)) or (inputs(249));
    layer0_outputs(9424) <= not((inputs(47)) and (inputs(229)));
    layer0_outputs(9425) <= '1';
    layer0_outputs(9426) <= (inputs(61)) xor (inputs(199));
    layer0_outputs(9427) <= not(inputs(53)) or (inputs(207));
    layer0_outputs(9428) <= (inputs(139)) and (inputs(20));
    layer0_outputs(9429) <= not((inputs(192)) or (inputs(226)));
    layer0_outputs(9430) <= not(inputs(233)) or (inputs(95));
    layer0_outputs(9431) <= not(inputs(116));
    layer0_outputs(9432) <= (inputs(52)) xor (inputs(226));
    layer0_outputs(9433) <= not(inputs(146));
    layer0_outputs(9434) <= '1';
    layer0_outputs(9435) <= inputs(169);
    layer0_outputs(9436) <= (inputs(141)) or (inputs(178));
    layer0_outputs(9437) <= (inputs(223)) xor (inputs(130));
    layer0_outputs(9438) <= not((inputs(251)) xor (inputs(255)));
    layer0_outputs(9439) <= not(inputs(127)) or (inputs(10));
    layer0_outputs(9440) <= not((inputs(130)) xor (inputs(249)));
    layer0_outputs(9441) <= not((inputs(4)) or (inputs(209)));
    layer0_outputs(9442) <= inputs(232);
    layer0_outputs(9443) <= '0';
    layer0_outputs(9444) <= not(inputs(247));
    layer0_outputs(9445) <= not(inputs(6)) or (inputs(235));
    layer0_outputs(9446) <= '0';
    layer0_outputs(9447) <= not(inputs(126)) or (inputs(245));
    layer0_outputs(9448) <= (inputs(165)) or (inputs(206));
    layer0_outputs(9449) <= not(inputs(84)) or (inputs(24));
    layer0_outputs(9450) <= not(inputs(98));
    layer0_outputs(9451) <= not(inputs(88));
    layer0_outputs(9452) <= not((inputs(187)) and (inputs(144)));
    layer0_outputs(9453) <= not(inputs(120)) or (inputs(113));
    layer0_outputs(9454) <= not(inputs(73));
    layer0_outputs(9455) <= not(inputs(176));
    layer0_outputs(9456) <= not(inputs(136));
    layer0_outputs(9457) <= not((inputs(235)) xor (inputs(208)));
    layer0_outputs(9458) <= not(inputs(22));
    layer0_outputs(9459) <= (inputs(63)) or (inputs(243));
    layer0_outputs(9460) <= (inputs(62)) xor (inputs(108));
    layer0_outputs(9461) <= '0';
    layer0_outputs(9462) <= not(inputs(91)) or (inputs(97));
    layer0_outputs(9463) <= not((inputs(109)) or (inputs(233)));
    layer0_outputs(9464) <= (inputs(112)) and not (inputs(73));
    layer0_outputs(9465) <= not(inputs(198));
    layer0_outputs(9466) <= not((inputs(0)) and (inputs(175)));
    layer0_outputs(9467) <= not((inputs(20)) or (inputs(242)));
    layer0_outputs(9468) <= inputs(214);
    layer0_outputs(9469) <= not((inputs(77)) or (inputs(123)));
    layer0_outputs(9470) <= not(inputs(159));
    layer0_outputs(9471) <= (inputs(123)) xor (inputs(45));
    layer0_outputs(9472) <= not(inputs(199)) or (inputs(191));
    layer0_outputs(9473) <= inputs(80);
    layer0_outputs(9474) <= '1';
    layer0_outputs(9475) <= not(inputs(160)) or (inputs(253));
    layer0_outputs(9476) <= not((inputs(119)) or (inputs(195)));
    layer0_outputs(9477) <= (inputs(66)) or (inputs(244));
    layer0_outputs(9478) <= '0';
    layer0_outputs(9479) <= not((inputs(72)) xor (inputs(123)));
    layer0_outputs(9480) <= (inputs(145)) and not (inputs(168));
    layer0_outputs(9481) <= '0';
    layer0_outputs(9482) <= '0';
    layer0_outputs(9483) <= (inputs(163)) or (inputs(220));
    layer0_outputs(9484) <= inputs(2);
    layer0_outputs(9485) <= not((inputs(48)) xor (inputs(252)));
    layer0_outputs(9486) <= '1';
    layer0_outputs(9487) <= not(inputs(231));
    layer0_outputs(9488) <= not((inputs(242)) and (inputs(144)));
    layer0_outputs(9489) <= not((inputs(92)) or (inputs(237)));
    layer0_outputs(9490) <= '1';
    layer0_outputs(9491) <= (inputs(194)) and not (inputs(81));
    layer0_outputs(9492) <= not((inputs(93)) xor (inputs(91)));
    layer0_outputs(9493) <= inputs(110);
    layer0_outputs(9494) <= (inputs(141)) or (inputs(79));
    layer0_outputs(9495) <= (inputs(8)) xor (inputs(191));
    layer0_outputs(9496) <= not(inputs(182));
    layer0_outputs(9497) <= (inputs(173)) xor (inputs(5));
    layer0_outputs(9498) <= not(inputs(195));
    layer0_outputs(9499) <= (inputs(93)) or (inputs(38));
    layer0_outputs(9500) <= not(inputs(108));
    layer0_outputs(9501) <= (inputs(243)) and not (inputs(224));
    layer0_outputs(9502) <= inputs(216);
    layer0_outputs(9503) <= (inputs(34)) and not (inputs(187));
    layer0_outputs(9504) <= not((inputs(186)) or (inputs(141)));
    layer0_outputs(9505) <= not(inputs(179));
    layer0_outputs(9506) <= not((inputs(11)) or (inputs(196)));
    layer0_outputs(9507) <= inputs(150);
    layer0_outputs(9508) <= inputs(0);
    layer0_outputs(9509) <= (inputs(117)) and not (inputs(93));
    layer0_outputs(9510) <= not((inputs(15)) and (inputs(190)));
    layer0_outputs(9511) <= (inputs(213)) or (inputs(73));
    layer0_outputs(9512) <= not(inputs(182));
    layer0_outputs(9513) <= inputs(70);
    layer0_outputs(9514) <= not((inputs(91)) xor (inputs(142)));
    layer0_outputs(9515) <= inputs(76);
    layer0_outputs(9516) <= '1';
    layer0_outputs(9517) <= '1';
    layer0_outputs(9518) <= inputs(6);
    layer0_outputs(9519) <= not(inputs(244));
    layer0_outputs(9520) <= not(inputs(68)) or (inputs(222));
    layer0_outputs(9521) <= not(inputs(120));
    layer0_outputs(9522) <= not(inputs(84));
    layer0_outputs(9523) <= inputs(124);
    layer0_outputs(9524) <= (inputs(195)) and not (inputs(45));
    layer0_outputs(9525) <= (inputs(146)) xor (inputs(176));
    layer0_outputs(9526) <= (inputs(203)) or (inputs(146));
    layer0_outputs(9527) <= (inputs(53)) or (inputs(69));
    layer0_outputs(9528) <= (inputs(17)) or (inputs(240));
    layer0_outputs(9529) <= (inputs(145)) and not (inputs(10));
    layer0_outputs(9530) <= not(inputs(122)) or (inputs(129));
    layer0_outputs(9531) <= inputs(55);
    layer0_outputs(9532) <= (inputs(156)) xor (inputs(190));
    layer0_outputs(9533) <= inputs(161);
    layer0_outputs(9534) <= not((inputs(236)) xor (inputs(172)));
    layer0_outputs(9535) <= (inputs(243)) or (inputs(115));
    layer0_outputs(9536) <= not(inputs(209)) or (inputs(198));
    layer0_outputs(9537) <= not(inputs(228)) or (inputs(1));
    layer0_outputs(9538) <= not((inputs(189)) xor (inputs(249)));
    layer0_outputs(9539) <= (inputs(47)) or (inputs(151));
    layer0_outputs(9540) <= not(inputs(33));
    layer0_outputs(9541) <= '0';
    layer0_outputs(9542) <= not(inputs(180)) or (inputs(173));
    layer0_outputs(9543) <= not(inputs(220)) or (inputs(22));
    layer0_outputs(9544) <= not(inputs(148)) or (inputs(105));
    layer0_outputs(9545) <= (inputs(213)) and not (inputs(47));
    layer0_outputs(9546) <= not(inputs(179));
    layer0_outputs(9547) <= (inputs(212)) and (inputs(29));
    layer0_outputs(9548) <= not(inputs(146));
    layer0_outputs(9549) <= not(inputs(222));
    layer0_outputs(9550) <= inputs(228);
    layer0_outputs(9551) <= not(inputs(203));
    layer0_outputs(9552) <= (inputs(154)) and not (inputs(245));
    layer0_outputs(9553) <= '0';
    layer0_outputs(9554) <= not((inputs(122)) or (inputs(229)));
    layer0_outputs(9555) <= inputs(247);
    layer0_outputs(9556) <= not((inputs(20)) or (inputs(61)));
    layer0_outputs(9557) <= not((inputs(44)) or (inputs(188)));
    layer0_outputs(9558) <= (inputs(96)) or (inputs(130));
    layer0_outputs(9559) <= (inputs(18)) and not (inputs(209));
    layer0_outputs(9560) <= (inputs(232)) and (inputs(166));
    layer0_outputs(9561) <= '0';
    layer0_outputs(9562) <= not(inputs(180)) or (inputs(46));
    layer0_outputs(9563) <= not(inputs(170));
    layer0_outputs(9564) <= not((inputs(167)) xor (inputs(216)));
    layer0_outputs(9565) <= (inputs(52)) xor (inputs(255));
    layer0_outputs(9566) <= not((inputs(95)) xor (inputs(189)));
    layer0_outputs(9567) <= inputs(193);
    layer0_outputs(9568) <= not(inputs(246)) or (inputs(113));
    layer0_outputs(9569) <= not((inputs(112)) xor (inputs(50)));
    layer0_outputs(9570) <= not((inputs(32)) xor (inputs(170)));
    layer0_outputs(9571) <= (inputs(99)) xor (inputs(102));
    layer0_outputs(9572) <= not((inputs(22)) xor (inputs(85)));
    layer0_outputs(9573) <= not(inputs(209));
    layer0_outputs(9574) <= not(inputs(255));
    layer0_outputs(9575) <= not(inputs(156));
    layer0_outputs(9576) <= (inputs(134)) or (inputs(26));
    layer0_outputs(9577) <= '0';
    layer0_outputs(9578) <= (inputs(66)) or (inputs(65));
    layer0_outputs(9579) <= not(inputs(142)) or (inputs(12));
    layer0_outputs(9580) <= inputs(188);
    layer0_outputs(9581) <= inputs(24);
    layer0_outputs(9582) <= not((inputs(112)) xor (inputs(116)));
    layer0_outputs(9583) <= not(inputs(147));
    layer0_outputs(9584) <= (inputs(201)) xor (inputs(203));
    layer0_outputs(9585) <= (inputs(143)) or (inputs(47));
    layer0_outputs(9586) <= not((inputs(209)) xor (inputs(246)));
    layer0_outputs(9587) <= (inputs(217)) and not (inputs(74));
    layer0_outputs(9588) <= not((inputs(156)) xor (inputs(159)));
    layer0_outputs(9589) <= (inputs(75)) xor (inputs(1));
    layer0_outputs(9590) <= (inputs(79)) and (inputs(18));
    layer0_outputs(9591) <= (inputs(223)) xor (inputs(79));
    layer0_outputs(9592) <= not(inputs(207));
    layer0_outputs(9593) <= inputs(129);
    layer0_outputs(9594) <= (inputs(82)) xor (inputs(168));
    layer0_outputs(9595) <= not((inputs(213)) or (inputs(144)));
    layer0_outputs(9596) <= not((inputs(12)) or (inputs(98)));
    layer0_outputs(9597) <= not(inputs(115));
    layer0_outputs(9598) <= not(inputs(115)) or (inputs(13));
    layer0_outputs(9599) <= not(inputs(133));
    layer0_outputs(9600) <= not(inputs(238)) or (inputs(35));
    layer0_outputs(9601) <= not(inputs(157));
    layer0_outputs(9602) <= (inputs(196)) and not (inputs(31));
    layer0_outputs(9603) <= (inputs(118)) and not (inputs(119));
    layer0_outputs(9604) <= inputs(229);
    layer0_outputs(9605) <= not((inputs(181)) and (inputs(24)));
    layer0_outputs(9606) <= not(inputs(126));
    layer0_outputs(9607) <= inputs(59);
    layer0_outputs(9608) <= not((inputs(179)) or (inputs(195)));
    layer0_outputs(9609) <= not(inputs(97));
    layer0_outputs(9610) <= not(inputs(69));
    layer0_outputs(9611) <= '0';
    layer0_outputs(9612) <= not((inputs(106)) or (inputs(171)));
    layer0_outputs(9613) <= not(inputs(7));
    layer0_outputs(9614) <= inputs(53);
    layer0_outputs(9615) <= not(inputs(190));
    layer0_outputs(9616) <= not(inputs(44)) or (inputs(146));
    layer0_outputs(9617) <= not(inputs(186)) or (inputs(165));
    layer0_outputs(9618) <= (inputs(200)) xor (inputs(231));
    layer0_outputs(9619) <= not(inputs(232)) or (inputs(225));
    layer0_outputs(9620) <= (inputs(197)) or (inputs(130));
    layer0_outputs(9621) <= inputs(24);
    layer0_outputs(9622) <= inputs(120);
    layer0_outputs(9623) <= not((inputs(72)) or (inputs(83)));
    layer0_outputs(9624) <= (inputs(24)) and not (inputs(179));
    layer0_outputs(9625) <= not(inputs(125));
    layer0_outputs(9626) <= inputs(11);
    layer0_outputs(9627) <= (inputs(23)) and not (inputs(192));
    layer0_outputs(9628) <= not(inputs(38)) or (inputs(157));
    layer0_outputs(9629) <= not(inputs(232)) or (inputs(223));
    layer0_outputs(9630) <= (inputs(178)) and not (inputs(18));
    layer0_outputs(9631) <= inputs(175);
    layer0_outputs(9632) <= inputs(24);
    layer0_outputs(9633) <= not((inputs(66)) or (inputs(154)));
    layer0_outputs(9634) <= not((inputs(175)) or (inputs(200)));
    layer0_outputs(9635) <= (inputs(213)) and (inputs(120));
    layer0_outputs(9636) <= not((inputs(171)) or (inputs(200)));
    layer0_outputs(9637) <= not(inputs(65));
    layer0_outputs(9638) <= not((inputs(73)) and (inputs(185)));
    layer0_outputs(9639) <= inputs(100);
    layer0_outputs(9640) <= (inputs(89)) and not (inputs(207));
    layer0_outputs(9641) <= (inputs(177)) or (inputs(211));
    layer0_outputs(9642) <= not((inputs(26)) and (inputs(234)));
    layer0_outputs(9643) <= (inputs(5)) or (inputs(158));
    layer0_outputs(9644) <= (inputs(100)) xor (inputs(181));
    layer0_outputs(9645) <= (inputs(223)) and not (inputs(156));
    layer0_outputs(9646) <= not(inputs(151)) or (inputs(8));
    layer0_outputs(9647) <= inputs(114);
    layer0_outputs(9648) <= not((inputs(250)) xor (inputs(81)));
    layer0_outputs(9649) <= '1';
    layer0_outputs(9650) <= (inputs(26)) and not (inputs(148));
    layer0_outputs(9651) <= not((inputs(97)) and (inputs(222)));
    layer0_outputs(9652) <= (inputs(255)) and not (inputs(121));
    layer0_outputs(9653) <= inputs(150);
    layer0_outputs(9654) <= not((inputs(50)) xor (inputs(69)));
    layer0_outputs(9655) <= inputs(77);
    layer0_outputs(9656) <= inputs(60);
    layer0_outputs(9657) <= inputs(84);
    layer0_outputs(9658) <= not((inputs(215)) or (inputs(78)));
    layer0_outputs(9659) <= not(inputs(196));
    layer0_outputs(9660) <= inputs(53);
    layer0_outputs(9661) <= not(inputs(149));
    layer0_outputs(9662) <= not((inputs(186)) or (inputs(51)));
    layer0_outputs(9663) <= not(inputs(198));
    layer0_outputs(9664) <= '0';
    layer0_outputs(9665) <= inputs(121);
    layer0_outputs(9666) <= not(inputs(229)) or (inputs(125));
    layer0_outputs(9667) <= not((inputs(193)) or (inputs(62)));
    layer0_outputs(9668) <= not(inputs(173)) or (inputs(45));
    layer0_outputs(9669) <= not(inputs(103));
    layer0_outputs(9670) <= not((inputs(155)) or (inputs(177)));
    layer0_outputs(9671) <= not(inputs(173));
    layer0_outputs(9672) <= '0';
    layer0_outputs(9673) <= not((inputs(75)) or (inputs(20)));
    layer0_outputs(9674) <= not((inputs(249)) or (inputs(11)));
    layer0_outputs(9675) <= not((inputs(18)) xor (inputs(57)));
    layer0_outputs(9676) <= not(inputs(70)) or (inputs(173));
    layer0_outputs(9677) <= (inputs(229)) and (inputs(21));
    layer0_outputs(9678) <= not(inputs(151));
    layer0_outputs(9679) <= not((inputs(112)) xor (inputs(87)));
    layer0_outputs(9680) <= (inputs(25)) or (inputs(33));
    layer0_outputs(9681) <= '0';
    layer0_outputs(9682) <= inputs(100);
    layer0_outputs(9683) <= not(inputs(204));
    layer0_outputs(9684) <= (inputs(40)) xor (inputs(191));
    layer0_outputs(9685) <= not(inputs(59)) or (inputs(191));
    layer0_outputs(9686) <= inputs(218);
    layer0_outputs(9687) <= '0';
    layer0_outputs(9688) <= not(inputs(122));
    layer0_outputs(9689) <= inputs(123);
    layer0_outputs(9690) <= not((inputs(28)) and (inputs(138)));
    layer0_outputs(9691) <= (inputs(99)) and not (inputs(215));
    layer0_outputs(9692) <= not(inputs(84));
    layer0_outputs(9693) <= not(inputs(235));
    layer0_outputs(9694) <= '1';
    layer0_outputs(9695) <= (inputs(238)) and not (inputs(17));
    layer0_outputs(9696) <= (inputs(28)) or (inputs(250));
    layer0_outputs(9697) <= inputs(224);
    layer0_outputs(9698) <= not(inputs(26)) or (inputs(198));
    layer0_outputs(9699) <= (inputs(177)) xor (inputs(174));
    layer0_outputs(9700) <= not((inputs(207)) or (inputs(94)));
    layer0_outputs(9701) <= not(inputs(140)) or (inputs(98));
    layer0_outputs(9702) <= not((inputs(169)) and (inputs(197)));
    layer0_outputs(9703) <= (inputs(58)) xor (inputs(238));
    layer0_outputs(9704) <= not(inputs(102));
    layer0_outputs(9705) <= not(inputs(135));
    layer0_outputs(9706) <= not((inputs(131)) or (inputs(226)));
    layer0_outputs(9707) <= (inputs(118)) and not (inputs(17));
    layer0_outputs(9708) <= (inputs(39)) and (inputs(57));
    layer0_outputs(9709) <= (inputs(91)) and not (inputs(34));
    layer0_outputs(9710) <= (inputs(188)) or (inputs(13));
    layer0_outputs(9711) <= not(inputs(248));
    layer0_outputs(9712) <= not(inputs(41));
    layer0_outputs(9713) <= (inputs(100)) or (inputs(100));
    layer0_outputs(9714) <= (inputs(21)) xor (inputs(255));
    layer0_outputs(9715) <= '0';
    layer0_outputs(9716) <= (inputs(126)) and not (inputs(97));
    layer0_outputs(9717) <= (inputs(63)) or (inputs(36));
    layer0_outputs(9718) <= not(inputs(229));
    layer0_outputs(9719) <= inputs(87);
    layer0_outputs(9720) <= (inputs(207)) and not (inputs(27));
    layer0_outputs(9721) <= not(inputs(103));
    layer0_outputs(9722) <= (inputs(33)) and not (inputs(174));
    layer0_outputs(9723) <= not((inputs(187)) xor (inputs(177)));
    layer0_outputs(9724) <= (inputs(87)) xor (inputs(129));
    layer0_outputs(9725) <= inputs(107);
    layer0_outputs(9726) <= not((inputs(81)) or (inputs(157)));
    layer0_outputs(9727) <= not(inputs(101));
    layer0_outputs(9728) <= '1';
    layer0_outputs(9729) <= inputs(33);
    layer0_outputs(9730) <= (inputs(4)) or (inputs(123));
    layer0_outputs(9731) <= not(inputs(49));
    layer0_outputs(9732) <= inputs(60);
    layer0_outputs(9733) <= not(inputs(36)) or (inputs(242));
    layer0_outputs(9734) <= not(inputs(192));
    layer0_outputs(9735) <= not(inputs(26)) or (inputs(54));
    layer0_outputs(9736) <= not(inputs(183));
    layer0_outputs(9737) <= not((inputs(210)) and (inputs(215)));
    layer0_outputs(9738) <= (inputs(15)) and not (inputs(217));
    layer0_outputs(9739) <= inputs(90);
    layer0_outputs(9740) <= not((inputs(132)) xor (inputs(163)));
    layer0_outputs(9741) <= not(inputs(102)) or (inputs(126));
    layer0_outputs(9742) <= (inputs(17)) and not (inputs(145));
    layer0_outputs(9743) <= not(inputs(20));
    layer0_outputs(9744) <= (inputs(96)) xor (inputs(114));
    layer0_outputs(9745) <= not(inputs(101));
    layer0_outputs(9746) <= inputs(175);
    layer0_outputs(9747) <= inputs(213);
    layer0_outputs(9748) <= inputs(29);
    layer0_outputs(9749) <= not(inputs(98)) or (inputs(75));
    layer0_outputs(9750) <= (inputs(158)) or (inputs(219));
    layer0_outputs(9751) <= not(inputs(99)) or (inputs(7));
    layer0_outputs(9752) <= not(inputs(135)) or (inputs(217));
    layer0_outputs(9753) <= not(inputs(32));
    layer0_outputs(9754) <= (inputs(172)) xor (inputs(208));
    layer0_outputs(9755) <= (inputs(65)) xor (inputs(53));
    layer0_outputs(9756) <= not((inputs(250)) or (inputs(196)));
    layer0_outputs(9757) <= inputs(159);
    layer0_outputs(9758) <= not((inputs(200)) xor (inputs(176)));
    layer0_outputs(9759) <= inputs(136);
    layer0_outputs(9760) <= not((inputs(235)) or (inputs(110)));
    layer0_outputs(9761) <= not(inputs(114)) or (inputs(114));
    layer0_outputs(9762) <= not((inputs(200)) xor (inputs(110)));
    layer0_outputs(9763) <= (inputs(21)) and not (inputs(179));
    layer0_outputs(9764) <= not(inputs(211)) or (inputs(236));
    layer0_outputs(9765) <= not(inputs(60));
    layer0_outputs(9766) <= not(inputs(131)) or (inputs(209));
    layer0_outputs(9767) <= not((inputs(70)) and (inputs(154)));
    layer0_outputs(9768) <= not(inputs(241));
    layer0_outputs(9769) <= (inputs(233)) xor (inputs(238));
    layer0_outputs(9770) <= not(inputs(85));
    layer0_outputs(9771) <= '0';
    layer0_outputs(9772) <= not(inputs(28));
    layer0_outputs(9773) <= not(inputs(57));
    layer0_outputs(9774) <= (inputs(135)) or (inputs(235));
    layer0_outputs(9775) <= (inputs(107)) and not (inputs(104));
    layer0_outputs(9776) <= (inputs(217)) and not (inputs(60));
    layer0_outputs(9777) <= (inputs(21)) or (inputs(26));
    layer0_outputs(9778) <= (inputs(79)) and not (inputs(250));
    layer0_outputs(9779) <= not(inputs(102));
    layer0_outputs(9780) <= not(inputs(104)) or (inputs(84));
    layer0_outputs(9781) <= not((inputs(40)) or (inputs(187)));
    layer0_outputs(9782) <= not((inputs(65)) and (inputs(191)));
    layer0_outputs(9783) <= not((inputs(1)) xor (inputs(96)));
    layer0_outputs(9784) <= not((inputs(170)) xor (inputs(65)));
    layer0_outputs(9785) <= (inputs(41)) and not (inputs(83));
    layer0_outputs(9786) <= inputs(22);
    layer0_outputs(9787) <= (inputs(65)) or (inputs(91));
    layer0_outputs(9788) <= (inputs(221)) xor (inputs(119));
    layer0_outputs(9789) <= (inputs(86)) and not (inputs(34));
    layer0_outputs(9790) <= (inputs(153)) and (inputs(13));
    layer0_outputs(9791) <= not(inputs(46));
    layer0_outputs(9792) <= (inputs(50)) xor (inputs(12));
    layer0_outputs(9793) <= inputs(99);
    layer0_outputs(9794) <= (inputs(227)) or (inputs(107));
    layer0_outputs(9795) <= not(inputs(207));
    layer0_outputs(9796) <= '1';
    layer0_outputs(9797) <= not(inputs(175));
    layer0_outputs(9798) <= not(inputs(50)) or (inputs(12));
    layer0_outputs(9799) <= (inputs(162)) xor (inputs(207));
    layer0_outputs(9800) <= not(inputs(75));
    layer0_outputs(9801) <= (inputs(132)) and not (inputs(160));
    layer0_outputs(9802) <= inputs(51);
    layer0_outputs(9803) <= not(inputs(22));
    layer0_outputs(9804) <= not(inputs(42));
    layer0_outputs(9805) <= not(inputs(42)) or (inputs(224));
    layer0_outputs(9806) <= (inputs(186)) xor (inputs(80));
    layer0_outputs(9807) <= (inputs(70)) xor (inputs(75));
    layer0_outputs(9808) <= not(inputs(133)) or (inputs(41));
    layer0_outputs(9809) <= (inputs(146)) or (inputs(247));
    layer0_outputs(9810) <= not(inputs(59)) or (inputs(173));
    layer0_outputs(9811) <= inputs(44);
    layer0_outputs(9812) <= not((inputs(71)) or (inputs(5)));
    layer0_outputs(9813) <= inputs(27);
    layer0_outputs(9814) <= inputs(110);
    layer0_outputs(9815) <= (inputs(2)) and (inputs(230));
    layer0_outputs(9816) <= (inputs(37)) or (inputs(124));
    layer0_outputs(9817) <= inputs(161);
    layer0_outputs(9818) <= not(inputs(60)) or (inputs(207));
    layer0_outputs(9819) <= not((inputs(2)) or (inputs(62)));
    layer0_outputs(9820) <= (inputs(213)) or (inputs(118));
    layer0_outputs(9821) <= inputs(121);
    layer0_outputs(9822) <= '1';
    layer0_outputs(9823) <= (inputs(142)) xor (inputs(80));
    layer0_outputs(9824) <= not((inputs(15)) or (inputs(74)));
    layer0_outputs(9825) <= (inputs(62)) or (inputs(32));
    layer0_outputs(9826) <= not(inputs(166));
    layer0_outputs(9827) <= inputs(131);
    layer0_outputs(9828) <= (inputs(104)) or (inputs(29));
    layer0_outputs(9829) <= inputs(137);
    layer0_outputs(9830) <= (inputs(209)) or (inputs(248));
    layer0_outputs(9831) <= not(inputs(105));
    layer0_outputs(9832) <= not(inputs(34));
    layer0_outputs(9833) <= not(inputs(140)) or (inputs(135));
    layer0_outputs(9834) <= not((inputs(165)) and (inputs(71)));
    layer0_outputs(9835) <= not(inputs(13));
    layer0_outputs(9836) <= (inputs(76)) xor (inputs(211));
    layer0_outputs(9837) <= (inputs(93)) xor (inputs(19));
    layer0_outputs(9838) <= not(inputs(82));
    layer0_outputs(9839) <= not(inputs(56));
    layer0_outputs(9840) <= (inputs(249)) and (inputs(189));
    layer0_outputs(9841) <= (inputs(167)) and not (inputs(117));
    layer0_outputs(9842) <= not((inputs(238)) and (inputs(17)));
    layer0_outputs(9843) <= not(inputs(108));
    layer0_outputs(9844) <= (inputs(245)) and (inputs(9));
    layer0_outputs(9845) <= (inputs(106)) xor (inputs(175));
    layer0_outputs(9846) <= inputs(54);
    layer0_outputs(9847) <= (inputs(111)) and not (inputs(78));
    layer0_outputs(9848) <= (inputs(13)) and (inputs(27));
    layer0_outputs(9849) <= (inputs(25)) and not (inputs(15));
    layer0_outputs(9850) <= not(inputs(192));
    layer0_outputs(9851) <= '1';
    layer0_outputs(9852) <= not(inputs(115)) or (inputs(29));
    layer0_outputs(9853) <= inputs(96);
    layer0_outputs(9854) <= (inputs(188)) and not (inputs(106));
    layer0_outputs(9855) <= not(inputs(196));
    layer0_outputs(9856) <= not(inputs(10));
    layer0_outputs(9857) <= inputs(51);
    layer0_outputs(9858) <= (inputs(53)) and not (inputs(190));
    layer0_outputs(9859) <= (inputs(239)) and (inputs(0));
    layer0_outputs(9860) <= not((inputs(75)) or (inputs(106)));
    layer0_outputs(9861) <= not(inputs(62));
    layer0_outputs(9862) <= not(inputs(42)) or (inputs(164));
    layer0_outputs(9863) <= not(inputs(59));
    layer0_outputs(9864) <= (inputs(212)) xor (inputs(244));
    layer0_outputs(9865) <= (inputs(150)) or (inputs(30));
    layer0_outputs(9866) <= not(inputs(49));
    layer0_outputs(9867) <= (inputs(85)) and not (inputs(143));
    layer0_outputs(9868) <= not(inputs(120));
    layer0_outputs(9869) <= not((inputs(177)) or (inputs(25)));
    layer0_outputs(9870) <= inputs(130);
    layer0_outputs(9871) <= not(inputs(218)) or (inputs(253));
    layer0_outputs(9872) <= inputs(232);
    layer0_outputs(9873) <= not((inputs(16)) and (inputs(138)));
    layer0_outputs(9874) <= inputs(253);
    layer0_outputs(9875) <= inputs(34);
    layer0_outputs(9876) <= not(inputs(7)) or (inputs(220));
    layer0_outputs(9877) <= not(inputs(232)) or (inputs(54));
    layer0_outputs(9878) <= (inputs(170)) xor (inputs(83));
    layer0_outputs(9879) <= inputs(183);
    layer0_outputs(9880) <= not(inputs(23));
    layer0_outputs(9881) <= not(inputs(243));
    layer0_outputs(9882) <= (inputs(127)) and not (inputs(220));
    layer0_outputs(9883) <= (inputs(149)) and not (inputs(123));
    layer0_outputs(9884) <= (inputs(87)) and not (inputs(81));
    layer0_outputs(9885) <= not(inputs(211)) or (inputs(73));
    layer0_outputs(9886) <= not((inputs(8)) xor (inputs(55)));
    layer0_outputs(9887) <= '0';
    layer0_outputs(9888) <= not(inputs(166));
    layer0_outputs(9889) <= (inputs(191)) and (inputs(6));
    layer0_outputs(9890) <= (inputs(177)) and not (inputs(135));
    layer0_outputs(9891) <= inputs(137);
    layer0_outputs(9892) <= '0';
    layer0_outputs(9893) <= not((inputs(106)) and (inputs(46)));
    layer0_outputs(9894) <= '0';
    layer0_outputs(9895) <= inputs(215);
    layer0_outputs(9896) <= not((inputs(255)) or (inputs(122)));
    layer0_outputs(9897) <= inputs(228);
    layer0_outputs(9898) <= (inputs(240)) or (inputs(156));
    layer0_outputs(9899) <= (inputs(212)) and (inputs(109));
    layer0_outputs(9900) <= inputs(98);
    layer0_outputs(9901) <= (inputs(131)) and not (inputs(33));
    layer0_outputs(9902) <= not(inputs(58));
    layer0_outputs(9903) <= not((inputs(83)) xor (inputs(132)));
    layer0_outputs(9904) <= not(inputs(136));
    layer0_outputs(9905) <= '1';
    layer0_outputs(9906) <= not(inputs(146));
    layer0_outputs(9907) <= not(inputs(136)) or (inputs(244));
    layer0_outputs(9908) <= (inputs(172)) or (inputs(55));
    layer0_outputs(9909) <= inputs(244);
    layer0_outputs(9910) <= (inputs(50)) or (inputs(60));
    layer0_outputs(9911) <= (inputs(10)) or (inputs(0));
    layer0_outputs(9912) <= not((inputs(40)) or (inputs(25)));
    layer0_outputs(9913) <= not((inputs(127)) and (inputs(141)));
    layer0_outputs(9914) <= (inputs(190)) or (inputs(123));
    layer0_outputs(9915) <= not((inputs(228)) or (inputs(187)));
    layer0_outputs(9916) <= inputs(33);
    layer0_outputs(9917) <= not(inputs(54));
    layer0_outputs(9918) <= not((inputs(128)) and (inputs(143)));
    layer0_outputs(9919) <= inputs(181);
    layer0_outputs(9920) <= inputs(231);
    layer0_outputs(9921) <= not(inputs(22)) or (inputs(240));
    layer0_outputs(9922) <= not(inputs(100));
    layer0_outputs(9923) <= not(inputs(81));
    layer0_outputs(9924) <= (inputs(153)) or (inputs(67));
    layer0_outputs(9925) <= not(inputs(16)) or (inputs(173));
    layer0_outputs(9926) <= not(inputs(56));
    layer0_outputs(9927) <= inputs(140);
    layer0_outputs(9928) <= (inputs(38)) or (inputs(131));
    layer0_outputs(9929) <= not(inputs(132));
    layer0_outputs(9930) <= (inputs(188)) or (inputs(202));
    layer0_outputs(9931) <= (inputs(205)) or (inputs(118));
    layer0_outputs(9932) <= inputs(60);
    layer0_outputs(9933) <= not(inputs(30)) or (inputs(127));
    layer0_outputs(9934) <= (inputs(71)) xor (inputs(229));
    layer0_outputs(9935) <= inputs(194);
    layer0_outputs(9936) <= not((inputs(199)) or (inputs(23)));
    layer0_outputs(9937) <= (inputs(85)) and not (inputs(140));
    layer0_outputs(9938) <= '1';
    layer0_outputs(9939) <= (inputs(144)) or (inputs(132));
    layer0_outputs(9940) <= not((inputs(52)) xor (inputs(39)));
    layer0_outputs(9941) <= '1';
    layer0_outputs(9942) <= (inputs(81)) or (inputs(215));
    layer0_outputs(9943) <= (inputs(62)) or (inputs(250));
    layer0_outputs(9944) <= (inputs(191)) or (inputs(179));
    layer0_outputs(9945) <= not((inputs(57)) xor (inputs(12)));
    layer0_outputs(9946) <= inputs(254);
    layer0_outputs(9947) <= '1';
    layer0_outputs(9948) <= (inputs(167)) and not (inputs(26));
    layer0_outputs(9949) <= inputs(165);
    layer0_outputs(9950) <= (inputs(149)) and not (inputs(0));
    layer0_outputs(9951) <= not(inputs(100));
    layer0_outputs(9952) <= not(inputs(163)) or (inputs(97));
    layer0_outputs(9953) <= inputs(25);
    layer0_outputs(9954) <= not(inputs(238));
    layer0_outputs(9955) <= (inputs(119)) and (inputs(149));
    layer0_outputs(9956) <= (inputs(245)) or (inputs(79));
    layer0_outputs(9957) <= not(inputs(25));
    layer0_outputs(9958) <= (inputs(103)) and not (inputs(127));
    layer0_outputs(9959) <= not((inputs(105)) or (inputs(66)));
    layer0_outputs(9960) <= not((inputs(223)) or (inputs(126)));
    layer0_outputs(9961) <= (inputs(190)) and not (inputs(242));
    layer0_outputs(9962) <= not((inputs(119)) xor (inputs(113)));
    layer0_outputs(9963) <= (inputs(52)) or (inputs(89));
    layer0_outputs(9964) <= (inputs(76)) and not (inputs(178));
    layer0_outputs(9965) <= (inputs(106)) or (inputs(239));
    layer0_outputs(9966) <= (inputs(46)) or (inputs(237));
    layer0_outputs(9967) <= (inputs(34)) and not (inputs(191));
    layer0_outputs(9968) <= not(inputs(48)) or (inputs(22));
    layer0_outputs(9969) <= not((inputs(192)) xor (inputs(243)));
    layer0_outputs(9970) <= (inputs(152)) and (inputs(189));
    layer0_outputs(9971) <= not((inputs(161)) xor (inputs(114)));
    layer0_outputs(9972) <= (inputs(138)) or (inputs(251));
    layer0_outputs(9973) <= inputs(94);
    layer0_outputs(9974) <= inputs(12);
    layer0_outputs(9975) <= inputs(59);
    layer0_outputs(9976) <= not((inputs(9)) xor (inputs(5)));
    layer0_outputs(9977) <= (inputs(197)) or (inputs(53));
    layer0_outputs(9978) <= (inputs(67)) xor (inputs(61));
    layer0_outputs(9979) <= (inputs(17)) and not (inputs(63));
    layer0_outputs(9980) <= inputs(213);
    layer0_outputs(9981) <= not(inputs(111)) or (inputs(244));
    layer0_outputs(9982) <= (inputs(216)) xor (inputs(161));
    layer0_outputs(9983) <= not(inputs(84));
    layer0_outputs(9984) <= not((inputs(128)) or (inputs(61)));
    layer0_outputs(9985) <= not(inputs(214)) or (inputs(125));
    layer0_outputs(9986) <= (inputs(229)) and not (inputs(95));
    layer0_outputs(9987) <= inputs(76);
    layer0_outputs(9988) <= not(inputs(11)) or (inputs(67));
    layer0_outputs(9989) <= '1';
    layer0_outputs(9990) <= inputs(205);
    layer0_outputs(9991) <= inputs(90);
    layer0_outputs(9992) <= not(inputs(191)) or (inputs(235));
    layer0_outputs(9993) <= not(inputs(160));
    layer0_outputs(9994) <= not(inputs(38)) or (inputs(112));
    layer0_outputs(9995) <= (inputs(164)) or (inputs(140));
    layer0_outputs(9996) <= not(inputs(126)) or (inputs(244));
    layer0_outputs(9997) <= not(inputs(91)) or (inputs(128));
    layer0_outputs(9998) <= (inputs(1)) or (inputs(165));
    layer0_outputs(9999) <= not(inputs(11)) or (inputs(200));
    layer0_outputs(10000) <= (inputs(251)) and (inputs(184));
    layer0_outputs(10001) <= not(inputs(7)) or (inputs(53));
    layer0_outputs(10002) <= (inputs(222)) or (inputs(246));
    layer0_outputs(10003) <= (inputs(141)) or (inputs(122));
    layer0_outputs(10004) <= not(inputs(102));
    layer0_outputs(10005) <= '0';
    layer0_outputs(10006) <= '1';
    layer0_outputs(10007) <= (inputs(67)) and (inputs(132));
    layer0_outputs(10008) <= not((inputs(25)) or (inputs(189)));
    layer0_outputs(10009) <= not((inputs(30)) and (inputs(45)));
    layer0_outputs(10010) <= inputs(123);
    layer0_outputs(10011) <= (inputs(188)) and not (inputs(153));
    layer0_outputs(10012) <= (inputs(91)) and not (inputs(235));
    layer0_outputs(10013) <= inputs(127);
    layer0_outputs(10014) <= (inputs(17)) or (inputs(154));
    layer0_outputs(10015) <= not(inputs(101)) or (inputs(126));
    layer0_outputs(10016) <= not(inputs(119));
    layer0_outputs(10017) <= (inputs(43)) or (inputs(46));
    layer0_outputs(10018) <= not(inputs(195)) or (inputs(44));
    layer0_outputs(10019) <= (inputs(95)) or (inputs(25));
    layer0_outputs(10020) <= not((inputs(251)) or (inputs(156)));
    layer0_outputs(10021) <= (inputs(29)) or (inputs(92));
    layer0_outputs(10022) <= '1';
    layer0_outputs(10023) <= (inputs(246)) and not (inputs(236));
    layer0_outputs(10024) <= not((inputs(174)) xor (inputs(62)));
    layer0_outputs(10025) <= (inputs(228)) xor (inputs(176));
    layer0_outputs(10026) <= inputs(149);
    layer0_outputs(10027) <= (inputs(248)) and not (inputs(7));
    layer0_outputs(10028) <= not((inputs(31)) xor (inputs(177)));
    layer0_outputs(10029) <= (inputs(76)) and (inputs(236));
    layer0_outputs(10030) <= not((inputs(152)) or (inputs(221)));
    layer0_outputs(10031) <= (inputs(177)) and not (inputs(96));
    layer0_outputs(10032) <= inputs(85);
    layer0_outputs(10033) <= (inputs(107)) and not (inputs(194));
    layer0_outputs(10034) <= not(inputs(24));
    layer0_outputs(10035) <= not(inputs(76));
    layer0_outputs(10036) <= not(inputs(172)) or (inputs(61));
    layer0_outputs(10037) <= inputs(130);
    layer0_outputs(10038) <= not(inputs(252));
    layer0_outputs(10039) <= not((inputs(237)) xor (inputs(93)));
    layer0_outputs(10040) <= not(inputs(246));
    layer0_outputs(10041) <= not((inputs(235)) and (inputs(246)));
    layer0_outputs(10042) <= not(inputs(209));
    layer0_outputs(10043) <= inputs(213);
    layer0_outputs(10044) <= not((inputs(155)) xor (inputs(197)));
    layer0_outputs(10045) <= not((inputs(191)) xor (inputs(100)));
    layer0_outputs(10046) <= not((inputs(206)) or (inputs(20)));
    layer0_outputs(10047) <= not((inputs(168)) or (inputs(60)));
    layer0_outputs(10048) <= (inputs(146)) and not (inputs(120));
    layer0_outputs(10049) <= inputs(211);
    layer0_outputs(10050) <= (inputs(222)) xor (inputs(78));
    layer0_outputs(10051) <= (inputs(50)) xor (inputs(155));
    layer0_outputs(10052) <= (inputs(195)) and not (inputs(110));
    layer0_outputs(10053) <= (inputs(46)) or (inputs(44));
    layer0_outputs(10054) <= not(inputs(254)) or (inputs(71));
    layer0_outputs(10055) <= inputs(197);
    layer0_outputs(10056) <= (inputs(213)) and not (inputs(14));
    layer0_outputs(10057) <= not(inputs(112));
    layer0_outputs(10058) <= not((inputs(192)) or (inputs(123)));
    layer0_outputs(10059) <= (inputs(131)) and (inputs(146));
    layer0_outputs(10060) <= not((inputs(217)) or (inputs(130)));
    layer0_outputs(10061) <= (inputs(190)) or (inputs(149));
    layer0_outputs(10062) <= inputs(86);
    layer0_outputs(10063) <= not(inputs(143));
    layer0_outputs(10064) <= not(inputs(155));
    layer0_outputs(10065) <= (inputs(113)) or (inputs(167));
    layer0_outputs(10066) <= not(inputs(190)) or (inputs(52));
    layer0_outputs(10067) <= (inputs(62)) or (inputs(160));
    layer0_outputs(10068) <= not(inputs(56));
    layer0_outputs(10069) <= not(inputs(218)) or (inputs(93));
    layer0_outputs(10070) <= not((inputs(154)) xor (inputs(4)));
    layer0_outputs(10071) <= inputs(180);
    layer0_outputs(10072) <= not((inputs(147)) xor (inputs(223)));
    layer0_outputs(10073) <= inputs(16);
    layer0_outputs(10074) <= not((inputs(206)) or (inputs(152)));
    layer0_outputs(10075) <= not(inputs(81)) or (inputs(30));
    layer0_outputs(10076) <= '0';
    layer0_outputs(10077) <= not(inputs(95)) or (inputs(172));
    layer0_outputs(10078) <= inputs(191);
    layer0_outputs(10079) <= inputs(124);
    layer0_outputs(10080) <= not((inputs(211)) or (inputs(145)));
    layer0_outputs(10081) <= (inputs(103)) xor (inputs(81));
    layer0_outputs(10082) <= inputs(97);
    layer0_outputs(10083) <= not((inputs(21)) or (inputs(31)));
    layer0_outputs(10084) <= not((inputs(25)) and (inputs(58)));
    layer0_outputs(10085) <= (inputs(227)) or (inputs(99));
    layer0_outputs(10086) <= not(inputs(196));
    layer0_outputs(10087) <= not(inputs(144));
    layer0_outputs(10088) <= inputs(29);
    layer0_outputs(10089) <= not((inputs(109)) xor (inputs(190)));
    layer0_outputs(10090) <= inputs(82);
    layer0_outputs(10091) <= not(inputs(31)) or (inputs(240));
    layer0_outputs(10092) <= inputs(73);
    layer0_outputs(10093) <= inputs(83);
    layer0_outputs(10094) <= not((inputs(47)) or (inputs(203)));
    layer0_outputs(10095) <= inputs(228);
    layer0_outputs(10096) <= not((inputs(135)) and (inputs(69)));
    layer0_outputs(10097) <= not(inputs(95)) or (inputs(65));
    layer0_outputs(10098) <= not((inputs(165)) or (inputs(249)));
    layer0_outputs(10099) <= (inputs(220)) or (inputs(207));
    layer0_outputs(10100) <= not(inputs(210));
    layer0_outputs(10101) <= inputs(223);
    layer0_outputs(10102) <= (inputs(97)) and not (inputs(151));
    layer0_outputs(10103) <= not(inputs(37));
    layer0_outputs(10104) <= not(inputs(179)) or (inputs(62));
    layer0_outputs(10105) <= (inputs(1)) and not (inputs(119));
    layer0_outputs(10106) <= (inputs(62)) and not (inputs(155));
    layer0_outputs(10107) <= not((inputs(141)) or (inputs(37)));
    layer0_outputs(10108) <= inputs(163);
    layer0_outputs(10109) <= not(inputs(124)) or (inputs(169));
    layer0_outputs(10110) <= not((inputs(98)) xor (inputs(21)));
    layer0_outputs(10111) <= inputs(63);
    layer0_outputs(10112) <= not(inputs(71));
    layer0_outputs(10113) <= not(inputs(214)) or (inputs(57));
    layer0_outputs(10114) <= (inputs(183)) and not (inputs(175));
    layer0_outputs(10115) <= (inputs(143)) or (inputs(149));
    layer0_outputs(10116) <= (inputs(245)) and not (inputs(113));
    layer0_outputs(10117) <= inputs(76);
    layer0_outputs(10118) <= (inputs(218)) and not (inputs(239));
    layer0_outputs(10119) <= (inputs(217)) or (inputs(252));
    layer0_outputs(10120) <= not(inputs(96));
    layer0_outputs(10121) <= not(inputs(36)) or (inputs(99));
    layer0_outputs(10122) <= not((inputs(96)) and (inputs(109)));
    layer0_outputs(10123) <= not(inputs(240));
    layer0_outputs(10124) <= not((inputs(179)) xor (inputs(247)));
    layer0_outputs(10125) <= inputs(243);
    layer0_outputs(10126) <= not((inputs(253)) xor (inputs(145)));
    layer0_outputs(10127) <= (inputs(86)) and not (inputs(170));
    layer0_outputs(10128) <= (inputs(178)) xor (inputs(247));
    layer0_outputs(10129) <= (inputs(211)) xor (inputs(15));
    layer0_outputs(10130) <= not((inputs(202)) xor (inputs(234)));
    layer0_outputs(10131) <= (inputs(157)) xor (inputs(8));
    layer0_outputs(10132) <= (inputs(121)) or (inputs(91));
    layer0_outputs(10133) <= not((inputs(113)) or (inputs(122)));
    layer0_outputs(10134) <= not(inputs(76));
    layer0_outputs(10135) <= not((inputs(204)) xor (inputs(144)));
    layer0_outputs(10136) <= '1';
    layer0_outputs(10137) <= (inputs(226)) or (inputs(5));
    layer0_outputs(10138) <= '1';
    layer0_outputs(10139) <= not((inputs(71)) xor (inputs(84)));
    layer0_outputs(10140) <= (inputs(47)) and not (inputs(184));
    layer0_outputs(10141) <= (inputs(11)) and not (inputs(68));
    layer0_outputs(10142) <= inputs(31);
    layer0_outputs(10143) <= (inputs(158)) and not (inputs(47));
    layer0_outputs(10144) <= (inputs(160)) xor (inputs(39));
    layer0_outputs(10145) <= (inputs(234)) and not (inputs(0));
    layer0_outputs(10146) <= not((inputs(164)) xor (inputs(135)));
    layer0_outputs(10147) <= inputs(83);
    layer0_outputs(10148) <= not(inputs(42)) or (inputs(106));
    layer0_outputs(10149) <= not((inputs(47)) or (inputs(13)));
    layer0_outputs(10150) <= inputs(191);
    layer0_outputs(10151) <= not(inputs(122)) or (inputs(174));
    layer0_outputs(10152) <= not((inputs(242)) and (inputs(186)));
    layer0_outputs(10153) <= inputs(92);
    layer0_outputs(10154) <= not((inputs(171)) or (inputs(221)));
    layer0_outputs(10155) <= not(inputs(142));
    layer0_outputs(10156) <= not(inputs(177)) or (inputs(10));
    layer0_outputs(10157) <= (inputs(75)) xor (inputs(175));
    layer0_outputs(10158) <= (inputs(31)) xor (inputs(156));
    layer0_outputs(10159) <= not((inputs(133)) or (inputs(30)));
    layer0_outputs(10160) <= inputs(137);
    layer0_outputs(10161) <= inputs(246);
    layer0_outputs(10162) <= (inputs(116)) and not (inputs(55));
    layer0_outputs(10163) <= not(inputs(114));
    layer0_outputs(10164) <= (inputs(145)) or (inputs(89));
    layer0_outputs(10165) <= not(inputs(33)) or (inputs(253));
    layer0_outputs(10166) <= not(inputs(103));
    layer0_outputs(10167) <= inputs(161);
    layer0_outputs(10168) <= not(inputs(155));
    layer0_outputs(10169) <= (inputs(180)) or (inputs(114));
    layer0_outputs(10170) <= not(inputs(149));
    layer0_outputs(10171) <= inputs(102);
    layer0_outputs(10172) <= (inputs(74)) and not (inputs(141));
    layer0_outputs(10173) <= (inputs(219)) or (inputs(251));
    layer0_outputs(10174) <= not((inputs(203)) xor (inputs(252)));
    layer0_outputs(10175) <= not((inputs(233)) or (inputs(39)));
    layer0_outputs(10176) <= not(inputs(179));
    layer0_outputs(10177) <= (inputs(22)) and not (inputs(160));
    layer0_outputs(10178) <= not(inputs(149));
    layer0_outputs(10179) <= (inputs(186)) and not (inputs(69));
    layer0_outputs(10180) <= not((inputs(52)) xor (inputs(117)));
    layer0_outputs(10181) <= not(inputs(24));
    layer0_outputs(10182) <= inputs(113);
    layer0_outputs(10183) <= not((inputs(182)) or (inputs(146)));
    layer0_outputs(10184) <= not(inputs(58)) or (inputs(210));
    layer0_outputs(10185) <= not((inputs(164)) or (inputs(56)));
    layer0_outputs(10186) <= (inputs(215)) xor (inputs(246));
    layer0_outputs(10187) <= not((inputs(128)) or (inputs(27)));
    layer0_outputs(10188) <= (inputs(100)) and (inputs(122));
    layer0_outputs(10189) <= (inputs(209)) and not (inputs(15));
    layer0_outputs(10190) <= (inputs(33)) and (inputs(48));
    layer0_outputs(10191) <= not((inputs(67)) xor (inputs(124)));
    layer0_outputs(10192) <= not(inputs(57)) or (inputs(183));
    layer0_outputs(10193) <= not(inputs(89));
    layer0_outputs(10194) <= inputs(165);
    layer0_outputs(10195) <= '1';
    layer0_outputs(10196) <= not((inputs(232)) or (inputs(211)));
    layer0_outputs(10197) <= not((inputs(117)) and (inputs(170)));
    layer0_outputs(10198) <= not((inputs(26)) or (inputs(7)));
    layer0_outputs(10199) <= inputs(68);
    layer0_outputs(10200) <= inputs(24);
    layer0_outputs(10201) <= (inputs(165)) and not (inputs(62));
    layer0_outputs(10202) <= not((inputs(58)) or (inputs(124)));
    layer0_outputs(10203) <= (inputs(35)) or (inputs(37));
    layer0_outputs(10204) <= not(inputs(176)) or (inputs(48));
    layer0_outputs(10205) <= not(inputs(207));
    layer0_outputs(10206) <= '1';
    layer0_outputs(10207) <= not((inputs(50)) or (inputs(172)));
    layer0_outputs(10208) <= not(inputs(77)) or (inputs(15));
    layer0_outputs(10209) <= inputs(0);
    layer0_outputs(10210) <= not((inputs(185)) xor (inputs(198)));
    layer0_outputs(10211) <= not(inputs(237));
    layer0_outputs(10212) <= not((inputs(160)) or (inputs(221)));
    layer0_outputs(10213) <= (inputs(30)) or (inputs(207));
    layer0_outputs(10214) <= not((inputs(126)) xor (inputs(89)));
    layer0_outputs(10215) <= inputs(224);
    layer0_outputs(10216) <= inputs(1);
    layer0_outputs(10217) <= not((inputs(225)) xor (inputs(248)));
    layer0_outputs(10218) <= not(inputs(255));
    layer0_outputs(10219) <= not(inputs(166));
    layer0_outputs(10220) <= not(inputs(43)) or (inputs(193));
    layer0_outputs(10221) <= inputs(209);
    layer0_outputs(10222) <= not(inputs(62));
    layer0_outputs(10223) <= not(inputs(116));
    layer0_outputs(10224) <= not(inputs(222)) or (inputs(116));
    layer0_outputs(10225) <= (inputs(217)) and (inputs(207));
    layer0_outputs(10226) <= not(inputs(119));
    layer0_outputs(10227) <= not(inputs(82));
    layer0_outputs(10228) <= not((inputs(194)) and (inputs(231)));
    layer0_outputs(10229) <= (inputs(126)) and not (inputs(12));
    layer0_outputs(10230) <= '0';
    layer0_outputs(10231) <= (inputs(93)) or (inputs(171));
    layer0_outputs(10232) <= inputs(179);
    layer0_outputs(10233) <= not(inputs(10)) or (inputs(152));
    layer0_outputs(10234) <= inputs(94);
    layer0_outputs(10235) <= '1';
    layer0_outputs(10236) <= not((inputs(148)) xor (inputs(68)));
    layer0_outputs(10237) <= (inputs(215)) and not (inputs(84));
    layer0_outputs(10238) <= inputs(197);
    layer0_outputs(10239) <= not(inputs(82));
    layer0_outputs(10240) <= (inputs(117)) xor (inputs(87));
    layer0_outputs(10241) <= (inputs(247)) or (inputs(91));
    layer0_outputs(10242) <= not(inputs(93));
    layer0_outputs(10243) <= inputs(216);
    layer0_outputs(10244) <= not(inputs(217)) or (inputs(141));
    layer0_outputs(10245) <= inputs(162);
    layer0_outputs(10246) <= not(inputs(99)) or (inputs(191));
    layer0_outputs(10247) <= inputs(93);
    layer0_outputs(10248) <= not(inputs(4));
    layer0_outputs(10249) <= not(inputs(212));
    layer0_outputs(10250) <= not((inputs(161)) or (inputs(172)));
    layer0_outputs(10251) <= inputs(194);
    layer0_outputs(10252) <= (inputs(203)) or (inputs(212));
    layer0_outputs(10253) <= inputs(76);
    layer0_outputs(10254) <= '0';
    layer0_outputs(10255) <= not((inputs(121)) or (inputs(165)));
    layer0_outputs(10256) <= (inputs(146)) and not (inputs(85));
    layer0_outputs(10257) <= (inputs(175)) xor (inputs(54));
    layer0_outputs(10258) <= not(inputs(26)) or (inputs(248));
    layer0_outputs(10259) <= inputs(67);
    layer0_outputs(10260) <= (inputs(212)) and not (inputs(9));
    layer0_outputs(10261) <= not(inputs(96));
    layer0_outputs(10262) <= '0';
    layer0_outputs(10263) <= not(inputs(26)) or (inputs(237));
    layer0_outputs(10264) <= inputs(122);
    layer0_outputs(10265) <= not(inputs(115)) or (inputs(233));
    layer0_outputs(10266) <= not((inputs(65)) xor (inputs(37)));
    layer0_outputs(10267) <= (inputs(9)) and (inputs(26));
    layer0_outputs(10268) <= not(inputs(78));
    layer0_outputs(10269) <= not(inputs(195)) or (inputs(159));
    layer0_outputs(10270) <= (inputs(196)) xor (inputs(2));
    layer0_outputs(10271) <= (inputs(19)) or (inputs(207));
    layer0_outputs(10272) <= not((inputs(42)) or (inputs(63)));
    layer0_outputs(10273) <= (inputs(44)) xor (inputs(63));
    layer0_outputs(10274) <= (inputs(172)) and not (inputs(13));
    layer0_outputs(10275) <= inputs(64);
    layer0_outputs(10276) <= not((inputs(49)) or (inputs(84)));
    layer0_outputs(10277) <= (inputs(132)) and not (inputs(185));
    layer0_outputs(10278) <= '0';
    layer0_outputs(10279) <= not(inputs(162)) or (inputs(93));
    layer0_outputs(10280) <= inputs(69);
    layer0_outputs(10281) <= (inputs(198)) xor (inputs(137));
    layer0_outputs(10282) <= not(inputs(203));
    layer0_outputs(10283) <= not((inputs(130)) or (inputs(161)));
    layer0_outputs(10284) <= not(inputs(113));
    layer0_outputs(10285) <= (inputs(22)) and not (inputs(222));
    layer0_outputs(10286) <= not(inputs(246));
    layer0_outputs(10287) <= inputs(125);
    layer0_outputs(10288) <= (inputs(20)) and not (inputs(28));
    layer0_outputs(10289) <= '1';
    layer0_outputs(10290) <= not((inputs(253)) or (inputs(107)));
    layer0_outputs(10291) <= (inputs(243)) xor (inputs(212));
    layer0_outputs(10292) <= not((inputs(253)) or (inputs(32)));
    layer0_outputs(10293) <= not(inputs(159));
    layer0_outputs(10294) <= (inputs(5)) or (inputs(166));
    layer0_outputs(10295) <= not((inputs(87)) and (inputs(124)));
    layer0_outputs(10296) <= (inputs(89)) and not (inputs(53));
    layer0_outputs(10297) <= inputs(77);
    layer0_outputs(10298) <= not((inputs(135)) or (inputs(71)));
    layer0_outputs(10299) <= (inputs(96)) or (inputs(66));
    layer0_outputs(10300) <= not((inputs(94)) xor (inputs(197)));
    layer0_outputs(10301) <= not(inputs(234));
    layer0_outputs(10302) <= not((inputs(142)) or (inputs(85)));
    layer0_outputs(10303) <= '0';
    layer0_outputs(10304) <= (inputs(69)) and not (inputs(145));
    layer0_outputs(10305) <= (inputs(26)) or (inputs(16));
    layer0_outputs(10306) <= inputs(156);
    layer0_outputs(10307) <= not((inputs(170)) xor (inputs(109)));
    layer0_outputs(10308) <= (inputs(231)) and (inputs(189));
    layer0_outputs(10309) <= not((inputs(172)) xor (inputs(48)));
    layer0_outputs(10310) <= not(inputs(74));
    layer0_outputs(10311) <= not(inputs(168));
    layer0_outputs(10312) <= not((inputs(182)) or (inputs(99)));
    layer0_outputs(10313) <= not((inputs(117)) xor (inputs(217)));
    layer0_outputs(10314) <= inputs(154);
    layer0_outputs(10315) <= not((inputs(35)) or (inputs(102)));
    layer0_outputs(10316) <= (inputs(108)) and (inputs(200));
    layer0_outputs(10317) <= (inputs(228)) or (inputs(197));
    layer0_outputs(10318) <= inputs(180);
    layer0_outputs(10319) <= inputs(202);
    layer0_outputs(10320) <= not(inputs(219)) or (inputs(69));
    layer0_outputs(10321) <= not(inputs(124));
    layer0_outputs(10322) <= inputs(31);
    layer0_outputs(10323) <= (inputs(125)) or (inputs(106));
    layer0_outputs(10324) <= not((inputs(130)) or (inputs(175)));
    layer0_outputs(10325) <= not(inputs(126));
    layer0_outputs(10326) <= not(inputs(221));
    layer0_outputs(10327) <= not(inputs(133));
    layer0_outputs(10328) <= not(inputs(83)) or (inputs(169));
    layer0_outputs(10329) <= (inputs(19)) or (inputs(32));
    layer0_outputs(10330) <= (inputs(216)) and not (inputs(60));
    layer0_outputs(10331) <= (inputs(217)) or (inputs(63));
    layer0_outputs(10332) <= inputs(173);
    layer0_outputs(10333) <= not((inputs(159)) xor (inputs(161)));
    layer0_outputs(10334) <= not((inputs(170)) or (inputs(203)));
    layer0_outputs(10335) <= not(inputs(157)) or (inputs(26));
    layer0_outputs(10336) <= not((inputs(3)) xor (inputs(209)));
    layer0_outputs(10337) <= not(inputs(173));
    layer0_outputs(10338) <= not(inputs(109)) or (inputs(52));
    layer0_outputs(10339) <= not(inputs(183)) or (inputs(68));
    layer0_outputs(10340) <= not((inputs(78)) or (inputs(119)));
    layer0_outputs(10341) <= (inputs(104)) or (inputs(87));
    layer0_outputs(10342) <= not((inputs(52)) and (inputs(154)));
    layer0_outputs(10343) <= not((inputs(61)) or (inputs(142)));
    layer0_outputs(10344) <= not(inputs(132)) or (inputs(3));
    layer0_outputs(10345) <= (inputs(193)) and not (inputs(91));
    layer0_outputs(10346) <= not(inputs(45));
    layer0_outputs(10347) <= inputs(5);
    layer0_outputs(10348) <= not(inputs(138)) or (inputs(65));
    layer0_outputs(10349) <= not((inputs(204)) xor (inputs(79)));
    layer0_outputs(10350) <= inputs(135);
    layer0_outputs(10351) <= inputs(60);
    layer0_outputs(10352) <= not((inputs(107)) and (inputs(133)));
    layer0_outputs(10353) <= not(inputs(255)) or (inputs(113));
    layer0_outputs(10354) <= inputs(233);
    layer0_outputs(10355) <= (inputs(10)) and not (inputs(119));
    layer0_outputs(10356) <= (inputs(59)) and not (inputs(236));
    layer0_outputs(10357) <= not((inputs(105)) and (inputs(122)));
    layer0_outputs(10358) <= (inputs(226)) or (inputs(17));
    layer0_outputs(10359) <= not((inputs(204)) and (inputs(56)));
    layer0_outputs(10360) <= not(inputs(133)) or (inputs(4));
    layer0_outputs(10361) <= (inputs(162)) and not (inputs(76));
    layer0_outputs(10362) <= not(inputs(115));
    layer0_outputs(10363) <= inputs(92);
    layer0_outputs(10364) <= not((inputs(7)) and (inputs(228)));
    layer0_outputs(10365) <= (inputs(223)) xor (inputs(51));
    layer0_outputs(10366) <= (inputs(91)) and not (inputs(116));
    layer0_outputs(10367) <= not((inputs(229)) or (inputs(225)));
    layer0_outputs(10368) <= not(inputs(175));
    layer0_outputs(10369) <= '1';
    layer0_outputs(10370) <= (inputs(98)) and not (inputs(87));
    layer0_outputs(10371) <= (inputs(90)) or (inputs(115));
    layer0_outputs(10372) <= not(inputs(251)) or (inputs(172));
    layer0_outputs(10373) <= not(inputs(182)) or (inputs(67));
    layer0_outputs(10374) <= not(inputs(167));
    layer0_outputs(10375) <= not(inputs(202));
    layer0_outputs(10376) <= not((inputs(105)) or (inputs(160)));
    layer0_outputs(10377) <= (inputs(163)) and not (inputs(224));
    layer0_outputs(10378) <= not((inputs(17)) or (inputs(143)));
    layer0_outputs(10379) <= '1';
    layer0_outputs(10380) <= (inputs(230)) and (inputs(165));
    layer0_outputs(10381) <= inputs(226);
    layer0_outputs(10382) <= inputs(96);
    layer0_outputs(10383) <= not(inputs(63)) or (inputs(254));
    layer0_outputs(10384) <= not(inputs(3));
    layer0_outputs(10385) <= inputs(120);
    layer0_outputs(10386) <= not(inputs(215));
    layer0_outputs(10387) <= not(inputs(118)) or (inputs(85));
    layer0_outputs(10388) <= not((inputs(48)) or (inputs(174)));
    layer0_outputs(10389) <= (inputs(73)) or (inputs(3));
    layer0_outputs(10390) <= (inputs(28)) and not (inputs(241));
    layer0_outputs(10391) <= not(inputs(26));
    layer0_outputs(10392) <= (inputs(192)) or (inputs(4));
    layer0_outputs(10393) <= (inputs(246)) or (inputs(154));
    layer0_outputs(10394) <= (inputs(227)) and (inputs(180));
    layer0_outputs(10395) <= (inputs(136)) and not (inputs(63));
    layer0_outputs(10396) <= (inputs(192)) xor (inputs(250));
    layer0_outputs(10397) <= not((inputs(55)) or (inputs(95)));
    layer0_outputs(10398) <= (inputs(148)) and not (inputs(137));
    layer0_outputs(10399) <= not((inputs(13)) or (inputs(52)));
    layer0_outputs(10400) <= (inputs(131)) and not (inputs(120));
    layer0_outputs(10401) <= not((inputs(129)) xor (inputs(103)));
    layer0_outputs(10402) <= (inputs(251)) xor (inputs(107));
    layer0_outputs(10403) <= '1';
    layer0_outputs(10404) <= not(inputs(198));
    layer0_outputs(10405) <= (inputs(170)) and not (inputs(87));
    layer0_outputs(10406) <= (inputs(218)) and not (inputs(18));
    layer0_outputs(10407) <= not(inputs(251)) or (inputs(242));
    layer0_outputs(10408) <= (inputs(213)) and not (inputs(158));
    layer0_outputs(10409) <= not(inputs(88));
    layer0_outputs(10410) <= not(inputs(42)) or (inputs(190));
    layer0_outputs(10411) <= (inputs(138)) xor (inputs(135));
    layer0_outputs(10412) <= inputs(248);
    layer0_outputs(10413) <= (inputs(224)) or (inputs(2));
    layer0_outputs(10414) <= '1';
    layer0_outputs(10415) <= not((inputs(40)) or (inputs(1)));
    layer0_outputs(10416) <= inputs(163);
    layer0_outputs(10417) <= not(inputs(86));
    layer0_outputs(10418) <= '0';
    layer0_outputs(10419) <= not((inputs(23)) or (inputs(36)));
    layer0_outputs(10420) <= (inputs(94)) and (inputs(136));
    layer0_outputs(10421) <= not(inputs(195)) or (inputs(136));
    layer0_outputs(10422) <= inputs(19);
    layer0_outputs(10423) <= not((inputs(40)) and (inputs(71)));
    layer0_outputs(10424) <= not((inputs(63)) xor (inputs(29)));
    layer0_outputs(10425) <= inputs(238);
    layer0_outputs(10426) <= (inputs(122)) and not (inputs(1));
    layer0_outputs(10427) <= not(inputs(37)) or (inputs(254));
    layer0_outputs(10428) <= (inputs(45)) or (inputs(208));
    layer0_outputs(10429) <= not(inputs(183));
    layer0_outputs(10430) <= not(inputs(216));
    layer0_outputs(10431) <= (inputs(202)) xor (inputs(185));
    layer0_outputs(10432) <= not((inputs(87)) xor (inputs(162)));
    layer0_outputs(10433) <= inputs(94);
    layer0_outputs(10434) <= not((inputs(158)) xor (inputs(116)));
    layer0_outputs(10435) <= (inputs(59)) or (inputs(123));
    layer0_outputs(10436) <= (inputs(36)) and not (inputs(103));
    layer0_outputs(10437) <= not((inputs(193)) or (inputs(22)));
    layer0_outputs(10438) <= inputs(105);
    layer0_outputs(10439) <= (inputs(168)) or (inputs(72));
    layer0_outputs(10440) <= not((inputs(63)) or (inputs(70)));
    layer0_outputs(10441) <= not(inputs(44)) or (inputs(238));
    layer0_outputs(10442) <= not(inputs(240)) or (inputs(175));
    layer0_outputs(10443) <= not((inputs(221)) and (inputs(249)));
    layer0_outputs(10444) <= not((inputs(5)) xor (inputs(45)));
    layer0_outputs(10445) <= (inputs(153)) and not (inputs(24));
    layer0_outputs(10446) <= (inputs(252)) or (inputs(150));
    layer0_outputs(10447) <= not((inputs(205)) or (inputs(175)));
    layer0_outputs(10448) <= (inputs(219)) and not (inputs(120));
    layer0_outputs(10449) <= inputs(212);
    layer0_outputs(10450) <= not((inputs(1)) xor (inputs(140)));
    layer0_outputs(10451) <= inputs(163);
    layer0_outputs(10452) <= (inputs(250)) xor (inputs(162));
    layer0_outputs(10453) <= (inputs(234)) xor (inputs(74));
    layer0_outputs(10454) <= (inputs(242)) or (inputs(167));
    layer0_outputs(10455) <= not(inputs(43)) or (inputs(200));
    layer0_outputs(10456) <= inputs(173);
    layer0_outputs(10457) <= not(inputs(229)) or (inputs(106));
    layer0_outputs(10458) <= (inputs(125)) and not (inputs(200));
    layer0_outputs(10459) <= (inputs(227)) and not (inputs(81));
    layer0_outputs(10460) <= (inputs(137)) xor (inputs(101));
    layer0_outputs(10461) <= (inputs(207)) or (inputs(7));
    layer0_outputs(10462) <= '1';
    layer0_outputs(10463) <= (inputs(183)) and not (inputs(13));
    layer0_outputs(10464) <= not(inputs(52)) or (inputs(71));
    layer0_outputs(10465) <= inputs(64);
    layer0_outputs(10466) <= (inputs(70)) or (inputs(58));
    layer0_outputs(10467) <= not((inputs(239)) or (inputs(159)));
    layer0_outputs(10468) <= not((inputs(193)) and (inputs(200)));
    layer0_outputs(10469) <= '1';
    layer0_outputs(10470) <= (inputs(108)) and not (inputs(48));
    layer0_outputs(10471) <= not(inputs(104));
    layer0_outputs(10472) <= not(inputs(139)) or (inputs(8));
    layer0_outputs(10473) <= inputs(76);
    layer0_outputs(10474) <= (inputs(49)) xor (inputs(22));
    layer0_outputs(10475) <= (inputs(244)) or (inputs(164));
    layer0_outputs(10476) <= '1';
    layer0_outputs(10477) <= not((inputs(9)) or (inputs(12)));
    layer0_outputs(10478) <= not((inputs(212)) or (inputs(192)));
    layer0_outputs(10479) <= not(inputs(58));
    layer0_outputs(10480) <= (inputs(103)) and not (inputs(42));
    layer0_outputs(10481) <= not((inputs(209)) xor (inputs(254)));
    layer0_outputs(10482) <= not(inputs(113));
    layer0_outputs(10483) <= not(inputs(155)) or (inputs(31));
    layer0_outputs(10484) <= not(inputs(225));
    layer0_outputs(10485) <= not((inputs(125)) xor (inputs(189)));
    layer0_outputs(10486) <= (inputs(141)) or (inputs(218));
    layer0_outputs(10487) <= (inputs(122)) and not (inputs(32));
    layer0_outputs(10488) <= (inputs(178)) or (inputs(241));
    layer0_outputs(10489) <= (inputs(40)) and (inputs(218));
    layer0_outputs(10490) <= not((inputs(129)) xor (inputs(223)));
    layer0_outputs(10491) <= (inputs(249)) and not (inputs(111));
    layer0_outputs(10492) <= (inputs(153)) and not (inputs(72));
    layer0_outputs(10493) <= not(inputs(235)) or (inputs(7));
    layer0_outputs(10494) <= not(inputs(210));
    layer0_outputs(10495) <= not((inputs(116)) or (inputs(6)));
    layer0_outputs(10496) <= (inputs(178)) and not (inputs(46));
    layer0_outputs(10497) <= not(inputs(173)) or (inputs(42));
    layer0_outputs(10498) <= not(inputs(119));
    layer0_outputs(10499) <= not(inputs(108)) or (inputs(151));
    layer0_outputs(10500) <= not((inputs(39)) or (inputs(5)));
    layer0_outputs(10501) <= not(inputs(4));
    layer0_outputs(10502) <= (inputs(166)) and not (inputs(157));
    layer0_outputs(10503) <= inputs(77);
    layer0_outputs(10504) <= not(inputs(189));
    layer0_outputs(10505) <= '1';
    layer0_outputs(10506) <= not((inputs(17)) and (inputs(117)));
    layer0_outputs(10507) <= not(inputs(219)) or (inputs(26));
    layer0_outputs(10508) <= not((inputs(246)) or (inputs(144)));
    layer0_outputs(10509) <= (inputs(21)) xor (inputs(37));
    layer0_outputs(10510) <= (inputs(174)) xor (inputs(179));
    layer0_outputs(10511) <= inputs(105);
    layer0_outputs(10512) <= (inputs(131)) and not (inputs(153));
    layer0_outputs(10513) <= not(inputs(14));
    layer0_outputs(10514) <= not((inputs(67)) or (inputs(146)));
    layer0_outputs(10515) <= not((inputs(237)) or (inputs(50)));
    layer0_outputs(10516) <= (inputs(194)) xor (inputs(219));
    layer0_outputs(10517) <= not(inputs(153)) or (inputs(108));
    layer0_outputs(10518) <= not(inputs(61));
    layer0_outputs(10519) <= inputs(24);
    layer0_outputs(10520) <= not(inputs(109));
    layer0_outputs(10521) <= '0';
    layer0_outputs(10522) <= (inputs(229)) or (inputs(191));
    layer0_outputs(10523) <= (inputs(204)) xor (inputs(224));
    layer0_outputs(10524) <= not(inputs(144)) or (inputs(255));
    layer0_outputs(10525) <= not(inputs(16));
    layer0_outputs(10526) <= not((inputs(96)) xor (inputs(139)));
    layer0_outputs(10527) <= not((inputs(30)) or (inputs(33)));
    layer0_outputs(10528) <= inputs(106);
    layer0_outputs(10529) <= (inputs(85)) and not (inputs(77));
    layer0_outputs(10530) <= not((inputs(75)) xor (inputs(19)));
    layer0_outputs(10531) <= (inputs(83)) or (inputs(233));
    layer0_outputs(10532) <= not((inputs(91)) or (inputs(111)));
    layer0_outputs(10533) <= '1';
    layer0_outputs(10534) <= not((inputs(131)) xor (inputs(145)));
    layer0_outputs(10535) <= inputs(29);
    layer0_outputs(10536) <= not((inputs(137)) and (inputs(174)));
    layer0_outputs(10537) <= (inputs(107)) xor (inputs(75));
    layer0_outputs(10538) <= not((inputs(169)) xor (inputs(123)));
    layer0_outputs(10539) <= (inputs(159)) and not (inputs(252));
    layer0_outputs(10540) <= (inputs(178)) xor (inputs(244));
    layer0_outputs(10541) <= not(inputs(7));
    layer0_outputs(10542) <= not(inputs(114));
    layer0_outputs(10543) <= not(inputs(204));
    layer0_outputs(10544) <= not(inputs(232)) or (inputs(97));
    layer0_outputs(10545) <= not((inputs(112)) xor (inputs(119)));
    layer0_outputs(10546) <= not(inputs(18));
    layer0_outputs(10547) <= not((inputs(174)) xor (inputs(17)));
    layer0_outputs(10548) <= not(inputs(198));
    layer0_outputs(10549) <= (inputs(140)) or (inputs(73));
    layer0_outputs(10550) <= inputs(152);
    layer0_outputs(10551) <= not((inputs(221)) or (inputs(13)));
    layer0_outputs(10552) <= not(inputs(56));
    layer0_outputs(10553) <= (inputs(28)) xor (inputs(154));
    layer0_outputs(10554) <= (inputs(79)) xor (inputs(206));
    layer0_outputs(10555) <= not((inputs(27)) or (inputs(107)));
    layer0_outputs(10556) <= not(inputs(2)) or (inputs(159));
    layer0_outputs(10557) <= (inputs(21)) or (inputs(253));
    layer0_outputs(10558) <= (inputs(99)) and (inputs(152));
    layer0_outputs(10559) <= (inputs(181)) and not (inputs(36));
    layer0_outputs(10560) <= not(inputs(216));
    layer0_outputs(10561) <= not(inputs(169)) or (inputs(4));
    layer0_outputs(10562) <= not((inputs(116)) xor (inputs(160)));
    layer0_outputs(10563) <= not(inputs(56)) or (inputs(18));
    layer0_outputs(10564) <= (inputs(71)) xor (inputs(188));
    layer0_outputs(10565) <= not((inputs(175)) xor (inputs(36)));
    layer0_outputs(10566) <= not((inputs(125)) xor (inputs(153)));
    layer0_outputs(10567) <= not((inputs(76)) and (inputs(90)));
    layer0_outputs(10568) <= not(inputs(30));
    layer0_outputs(10569) <= not((inputs(92)) and (inputs(138)));
    layer0_outputs(10570) <= (inputs(15)) and not (inputs(201));
    layer0_outputs(10571) <= not(inputs(208)) or (inputs(226));
    layer0_outputs(10572) <= not((inputs(100)) xor (inputs(118)));
    layer0_outputs(10573) <= (inputs(94)) xor (inputs(66));
    layer0_outputs(10574) <= (inputs(199)) and not (inputs(113));
    layer0_outputs(10575) <= not((inputs(103)) or (inputs(36)));
    layer0_outputs(10576) <= (inputs(166)) and not (inputs(18));
    layer0_outputs(10577) <= inputs(129);
    layer0_outputs(10578) <= not(inputs(51)) or (inputs(147));
    layer0_outputs(10579) <= not(inputs(51)) or (inputs(198));
    layer0_outputs(10580) <= (inputs(104)) or (inputs(67));
    layer0_outputs(10581) <= (inputs(254)) xor (inputs(181));
    layer0_outputs(10582) <= not(inputs(136));
    layer0_outputs(10583) <= (inputs(184)) and (inputs(210));
    layer0_outputs(10584) <= not(inputs(199)) or (inputs(139));
    layer0_outputs(10585) <= not(inputs(72)) or (inputs(1));
    layer0_outputs(10586) <= (inputs(231)) and (inputs(188));
    layer0_outputs(10587) <= (inputs(251)) xor (inputs(166));
    layer0_outputs(10588) <= not(inputs(129));
    layer0_outputs(10589) <= not(inputs(133)) or (inputs(18));
    layer0_outputs(10590) <= '0';
    layer0_outputs(10591) <= (inputs(130)) and not (inputs(195));
    layer0_outputs(10592) <= '1';
    layer0_outputs(10593) <= inputs(237);
    layer0_outputs(10594) <= '0';
    layer0_outputs(10595) <= inputs(19);
    layer0_outputs(10596) <= (inputs(33)) or (inputs(208));
    layer0_outputs(10597) <= not(inputs(119));
    layer0_outputs(10598) <= not((inputs(146)) xor (inputs(165)));
    layer0_outputs(10599) <= '1';
    layer0_outputs(10600) <= not((inputs(158)) or (inputs(235)));
    layer0_outputs(10601) <= (inputs(113)) and (inputs(217));
    layer0_outputs(10602) <= inputs(136);
    layer0_outputs(10603) <= (inputs(216)) or (inputs(171));
    layer0_outputs(10604) <= '1';
    layer0_outputs(10605) <= not(inputs(78)) or (inputs(112));
    layer0_outputs(10606) <= (inputs(158)) and not (inputs(205));
    layer0_outputs(10607) <= inputs(8);
    layer0_outputs(10608) <= not(inputs(107)) or (inputs(14));
    layer0_outputs(10609) <= inputs(209);
    layer0_outputs(10610) <= inputs(133);
    layer0_outputs(10611) <= (inputs(80)) or (inputs(189));
    layer0_outputs(10612) <= not(inputs(30)) or (inputs(187));
    layer0_outputs(10613) <= not(inputs(3));
    layer0_outputs(10614) <= not((inputs(182)) xor (inputs(81)));
    layer0_outputs(10615) <= not(inputs(92)) or (inputs(252));
    layer0_outputs(10616) <= inputs(43);
    layer0_outputs(10617) <= (inputs(174)) or (inputs(206));
    layer0_outputs(10618) <= inputs(76);
    layer0_outputs(10619) <= inputs(84);
    layer0_outputs(10620) <= (inputs(241)) and (inputs(224));
    layer0_outputs(10621) <= not((inputs(206)) or (inputs(221)));
    layer0_outputs(10622) <= (inputs(34)) or (inputs(47));
    layer0_outputs(10623) <= not(inputs(108));
    layer0_outputs(10624) <= inputs(138);
    layer0_outputs(10625) <= not((inputs(214)) or (inputs(105)));
    layer0_outputs(10626) <= (inputs(106)) or (inputs(73));
    layer0_outputs(10627) <= (inputs(51)) and (inputs(59));
    layer0_outputs(10628) <= not((inputs(211)) or (inputs(237)));
    layer0_outputs(10629) <= not((inputs(68)) or (inputs(220)));
    layer0_outputs(10630) <= not((inputs(133)) and (inputs(162)));
    layer0_outputs(10631) <= (inputs(188)) or (inputs(187));
    layer0_outputs(10632) <= not(inputs(53));
    layer0_outputs(10633) <= (inputs(111)) or (inputs(41));
    layer0_outputs(10634) <= (inputs(102)) and not (inputs(0));
    layer0_outputs(10635) <= (inputs(211)) xor (inputs(181));
    layer0_outputs(10636) <= inputs(11);
    layer0_outputs(10637) <= not((inputs(89)) or (inputs(221)));
    layer0_outputs(10638) <= inputs(209);
    layer0_outputs(10639) <= '1';
    layer0_outputs(10640) <= not(inputs(91));
    layer0_outputs(10641) <= not((inputs(118)) xor (inputs(79)));
    layer0_outputs(10642) <= (inputs(188)) and not (inputs(242));
    layer0_outputs(10643) <= inputs(166);
    layer0_outputs(10644) <= (inputs(57)) and (inputs(4));
    layer0_outputs(10645) <= not(inputs(2)) or (inputs(80));
    layer0_outputs(10646) <= inputs(218);
    layer0_outputs(10647) <= not((inputs(255)) or (inputs(102)));
    layer0_outputs(10648) <= (inputs(25)) or (inputs(25));
    layer0_outputs(10649) <= inputs(38);
    layer0_outputs(10650) <= not(inputs(198)) or (inputs(239));
    layer0_outputs(10651) <= (inputs(9)) or (inputs(203));
    layer0_outputs(10652) <= not((inputs(79)) xor (inputs(28)));
    layer0_outputs(10653) <= inputs(166);
    layer0_outputs(10654) <= not((inputs(164)) or (inputs(29)));
    layer0_outputs(10655) <= not((inputs(97)) or (inputs(82)));
    layer0_outputs(10656) <= not(inputs(197)) or (inputs(201));
    layer0_outputs(10657) <= not(inputs(58));
    layer0_outputs(10658) <= (inputs(177)) or (inputs(35));
    layer0_outputs(10659) <= inputs(72);
    layer0_outputs(10660) <= '0';
    layer0_outputs(10661) <= (inputs(215)) xor (inputs(171));
    layer0_outputs(10662) <= (inputs(210)) xor (inputs(104));
    layer0_outputs(10663) <= (inputs(139)) xor (inputs(219));
    layer0_outputs(10664) <= '1';
    layer0_outputs(10665) <= (inputs(104)) and not (inputs(225));
    layer0_outputs(10666) <= not(inputs(92));
    layer0_outputs(10667) <= (inputs(152)) and (inputs(40));
    layer0_outputs(10668) <= (inputs(241)) and (inputs(189));
    layer0_outputs(10669) <= not(inputs(215)) or (inputs(241));
    layer0_outputs(10670) <= not(inputs(231));
    layer0_outputs(10671) <= not(inputs(229));
    layer0_outputs(10672) <= (inputs(163)) and not (inputs(63));
    layer0_outputs(10673) <= not(inputs(197));
    layer0_outputs(10674) <= not((inputs(50)) xor (inputs(5)));
    layer0_outputs(10675) <= not(inputs(138));
    layer0_outputs(10676) <= '0';
    layer0_outputs(10677) <= not((inputs(81)) xor (inputs(147)));
    layer0_outputs(10678) <= not((inputs(171)) or (inputs(86)));
    layer0_outputs(10679) <= (inputs(15)) and not (inputs(143));
    layer0_outputs(10680) <= not(inputs(246));
    layer0_outputs(10681) <= not(inputs(104));
    layer0_outputs(10682) <= not(inputs(156)) or (inputs(254));
    layer0_outputs(10683) <= inputs(21);
    layer0_outputs(10684) <= (inputs(133)) or (inputs(6));
    layer0_outputs(10685) <= (inputs(128)) and not (inputs(82));
    layer0_outputs(10686) <= not(inputs(196));
    layer0_outputs(10687) <= inputs(183);
    layer0_outputs(10688) <= not((inputs(194)) and (inputs(119)));
    layer0_outputs(10689) <= inputs(37);
    layer0_outputs(10690) <= (inputs(227)) or (inputs(52));
    layer0_outputs(10691) <= (inputs(99)) and not (inputs(188));
    layer0_outputs(10692) <= (inputs(72)) xor (inputs(103));
    layer0_outputs(10693) <= (inputs(136)) xor (inputs(252));
    layer0_outputs(10694) <= not(inputs(94));
    layer0_outputs(10695) <= inputs(188);
    layer0_outputs(10696) <= not((inputs(28)) or (inputs(98)));
    layer0_outputs(10697) <= (inputs(212)) or (inputs(73));
    layer0_outputs(10698) <= not(inputs(162));
    layer0_outputs(10699) <= not(inputs(82)) or (inputs(192));
    layer0_outputs(10700) <= not(inputs(149));
    layer0_outputs(10701) <= not((inputs(227)) or (inputs(251)));
    layer0_outputs(10702) <= not(inputs(56));
    layer0_outputs(10703) <= not((inputs(199)) or (inputs(97)));
    layer0_outputs(10704) <= (inputs(66)) or (inputs(35));
    layer0_outputs(10705) <= (inputs(85)) and not (inputs(191));
    layer0_outputs(10706) <= (inputs(196)) xor (inputs(222));
    layer0_outputs(10707) <= inputs(134);
    layer0_outputs(10708) <= (inputs(64)) or (inputs(173));
    layer0_outputs(10709) <= (inputs(52)) and not (inputs(130));
    layer0_outputs(10710) <= not((inputs(147)) and (inputs(86)));
    layer0_outputs(10711) <= (inputs(251)) and not (inputs(168));
    layer0_outputs(10712) <= '1';
    layer0_outputs(10713) <= (inputs(26)) and not (inputs(253));
    layer0_outputs(10714) <= inputs(188);
    layer0_outputs(10715) <= not(inputs(180));
    layer0_outputs(10716) <= not((inputs(179)) or (inputs(215)));
    layer0_outputs(10717) <= inputs(70);
    layer0_outputs(10718) <= (inputs(162)) or (inputs(130));
    layer0_outputs(10719) <= '0';
    layer0_outputs(10720) <= not(inputs(129));
    layer0_outputs(10721) <= not(inputs(54));
    layer0_outputs(10722) <= (inputs(188)) or (inputs(152));
    layer0_outputs(10723) <= (inputs(58)) and (inputs(109));
    layer0_outputs(10724) <= (inputs(42)) or (inputs(54));
    layer0_outputs(10725) <= '0';
    layer0_outputs(10726) <= (inputs(156)) and not (inputs(37));
    layer0_outputs(10727) <= (inputs(32)) xor (inputs(164));
    layer0_outputs(10728) <= inputs(155);
    layer0_outputs(10729) <= not(inputs(0));
    layer0_outputs(10730) <= (inputs(193)) or (inputs(81));
    layer0_outputs(10731) <= not(inputs(227)) or (inputs(102));
    layer0_outputs(10732) <= (inputs(207)) xor (inputs(69));
    layer0_outputs(10733) <= not(inputs(242));
    layer0_outputs(10734) <= not(inputs(56));
    layer0_outputs(10735) <= (inputs(170)) and (inputs(161));
    layer0_outputs(10736) <= (inputs(101)) or (inputs(103));
    layer0_outputs(10737) <= not((inputs(58)) xor (inputs(242)));
    layer0_outputs(10738) <= inputs(233);
    layer0_outputs(10739) <= inputs(204);
    layer0_outputs(10740) <= (inputs(148)) and not (inputs(252));
    layer0_outputs(10741) <= inputs(253);
    layer0_outputs(10742) <= not(inputs(173));
    layer0_outputs(10743) <= (inputs(27)) and not (inputs(88));
    layer0_outputs(10744) <= inputs(113);
    layer0_outputs(10745) <= inputs(103);
    layer0_outputs(10746) <= (inputs(197)) or (inputs(168));
    layer0_outputs(10747) <= inputs(92);
    layer0_outputs(10748) <= not(inputs(56));
    layer0_outputs(10749) <= not((inputs(81)) xor (inputs(74)));
    layer0_outputs(10750) <= (inputs(124)) and not (inputs(253));
    layer0_outputs(10751) <= (inputs(32)) xor (inputs(95));
    layer0_outputs(10752) <= not((inputs(84)) or (inputs(173)));
    layer0_outputs(10753) <= not(inputs(142)) or (inputs(88));
    layer0_outputs(10754) <= (inputs(42)) and not (inputs(83));
    layer0_outputs(10755) <= (inputs(24)) xor (inputs(226));
    layer0_outputs(10756) <= (inputs(192)) and (inputs(135));
    layer0_outputs(10757) <= not((inputs(194)) or (inputs(153)));
    layer0_outputs(10758) <= (inputs(195)) and (inputs(43));
    layer0_outputs(10759) <= not(inputs(151));
    layer0_outputs(10760) <= not(inputs(100));
    layer0_outputs(10761) <= not(inputs(229));
    layer0_outputs(10762) <= not((inputs(126)) xor (inputs(107)));
    layer0_outputs(10763) <= (inputs(26)) or (inputs(205));
    layer0_outputs(10764) <= '0';
    layer0_outputs(10765) <= not(inputs(204));
    layer0_outputs(10766) <= inputs(88);
    layer0_outputs(10767) <= (inputs(121)) and not (inputs(243));
    layer0_outputs(10768) <= inputs(74);
    layer0_outputs(10769) <= not(inputs(187));
    layer0_outputs(10770) <= (inputs(182)) and (inputs(106));
    layer0_outputs(10771) <= '1';
    layer0_outputs(10772) <= not(inputs(102)) or (inputs(254));
    layer0_outputs(10773) <= (inputs(48)) xor (inputs(211));
    layer0_outputs(10774) <= (inputs(180)) and not (inputs(165));
    layer0_outputs(10775) <= inputs(93);
    layer0_outputs(10776) <= (inputs(28)) or (inputs(75));
    layer0_outputs(10777) <= not(inputs(167));
    layer0_outputs(10778) <= inputs(149);
    layer0_outputs(10779) <= not(inputs(146)) or (inputs(45));
    layer0_outputs(10780) <= inputs(27);
    layer0_outputs(10781) <= not(inputs(61)) or (inputs(72));
    layer0_outputs(10782) <= inputs(233);
    layer0_outputs(10783) <= not(inputs(226)) or (inputs(47));
    layer0_outputs(10784) <= not(inputs(231));
    layer0_outputs(10785) <= not(inputs(72)) or (inputs(44));
    layer0_outputs(10786) <= not((inputs(84)) xor (inputs(71)));
    layer0_outputs(10787) <= (inputs(248)) and not (inputs(20));
    layer0_outputs(10788) <= not(inputs(89));
    layer0_outputs(10789) <= inputs(134);
    layer0_outputs(10790) <= not(inputs(178));
    layer0_outputs(10791) <= (inputs(84)) xor (inputs(134));
    layer0_outputs(10792) <= (inputs(150)) and not (inputs(209));
    layer0_outputs(10793) <= not((inputs(69)) or (inputs(113)));
    layer0_outputs(10794) <= not(inputs(199)) or (inputs(2));
    layer0_outputs(10795) <= not(inputs(188)) or (inputs(68));
    layer0_outputs(10796) <= not(inputs(45));
    layer0_outputs(10797) <= not((inputs(165)) xor (inputs(205)));
    layer0_outputs(10798) <= inputs(178);
    layer0_outputs(10799) <= (inputs(74)) or (inputs(19));
    layer0_outputs(10800) <= not((inputs(89)) and (inputs(54)));
    layer0_outputs(10801) <= not(inputs(119));
    layer0_outputs(10802) <= (inputs(177)) and (inputs(224));
    layer0_outputs(10803) <= not((inputs(1)) xor (inputs(63)));
    layer0_outputs(10804) <= inputs(165);
    layer0_outputs(10805) <= not((inputs(90)) xor (inputs(181)));
    layer0_outputs(10806) <= (inputs(112)) or (inputs(193));
    layer0_outputs(10807) <= not((inputs(124)) or (inputs(255)));
    layer0_outputs(10808) <= not((inputs(234)) or (inputs(195)));
    layer0_outputs(10809) <= (inputs(78)) and not (inputs(142));
    layer0_outputs(10810) <= not((inputs(90)) xor (inputs(72)));
    layer0_outputs(10811) <= inputs(138);
    layer0_outputs(10812) <= not((inputs(7)) or (inputs(110)));
    layer0_outputs(10813) <= not(inputs(2)) or (inputs(223));
    layer0_outputs(10814) <= not(inputs(231)) or (inputs(69));
    layer0_outputs(10815) <= not((inputs(222)) and (inputs(45)));
    layer0_outputs(10816) <= (inputs(213)) or (inputs(210));
    layer0_outputs(10817) <= inputs(219);
    layer0_outputs(10818) <= not(inputs(208)) or (inputs(36));
    layer0_outputs(10819) <= (inputs(175)) or (inputs(118));
    layer0_outputs(10820) <= inputs(214);
    layer0_outputs(10821) <= not((inputs(132)) and (inputs(124)));
    layer0_outputs(10822) <= not((inputs(32)) xor (inputs(154)));
    layer0_outputs(10823) <= '1';
    layer0_outputs(10824) <= inputs(161);
    layer0_outputs(10825) <= inputs(87);
    layer0_outputs(10826) <= not((inputs(227)) or (inputs(171)));
    layer0_outputs(10827) <= not((inputs(112)) or (inputs(113)));
    layer0_outputs(10828) <= (inputs(198)) xor (inputs(36));
    layer0_outputs(10829) <= (inputs(142)) or (inputs(1));
    layer0_outputs(10830) <= (inputs(248)) and not (inputs(45));
    layer0_outputs(10831) <= inputs(50);
    layer0_outputs(10832) <= inputs(183);
    layer0_outputs(10833) <= not(inputs(87));
    layer0_outputs(10834) <= (inputs(222)) or (inputs(250));
    layer0_outputs(10835) <= not(inputs(150)) or (inputs(141));
    layer0_outputs(10836) <= inputs(205);
    layer0_outputs(10837) <= not(inputs(222)) or (inputs(133));
    layer0_outputs(10838) <= (inputs(29)) or (inputs(170));
    layer0_outputs(10839) <= (inputs(98)) or (inputs(80));
    layer0_outputs(10840) <= not(inputs(223));
    layer0_outputs(10841) <= not(inputs(176)) or (inputs(143));
    layer0_outputs(10842) <= not(inputs(25)) or (inputs(193));
    layer0_outputs(10843) <= (inputs(54)) or (inputs(109));
    layer0_outputs(10844) <= (inputs(191)) or (inputs(4));
    layer0_outputs(10845) <= (inputs(128)) xor (inputs(112));
    layer0_outputs(10846) <= not(inputs(83));
    layer0_outputs(10847) <= not(inputs(118)) or (inputs(217));
    layer0_outputs(10848) <= not(inputs(78));
    layer0_outputs(10849) <= not(inputs(145)) or (inputs(14));
    layer0_outputs(10850) <= inputs(229);
    layer0_outputs(10851) <= not(inputs(73)) or (inputs(226));
    layer0_outputs(10852) <= '0';
    layer0_outputs(10853) <= not((inputs(34)) or (inputs(116)));
    layer0_outputs(10854) <= (inputs(87)) and (inputs(203));
    layer0_outputs(10855) <= (inputs(19)) or (inputs(111));
    layer0_outputs(10856) <= inputs(105);
    layer0_outputs(10857) <= (inputs(224)) and (inputs(203));
    layer0_outputs(10858) <= not((inputs(24)) xor (inputs(81)));
    layer0_outputs(10859) <= (inputs(201)) and not (inputs(106));
    layer0_outputs(10860) <= not(inputs(91)) or (inputs(193));
    layer0_outputs(10861) <= inputs(234);
    layer0_outputs(10862) <= inputs(105);
    layer0_outputs(10863) <= (inputs(23)) and not (inputs(72));
    layer0_outputs(10864) <= (inputs(185)) or (inputs(19));
    layer0_outputs(10865) <= '0';
    layer0_outputs(10866) <= inputs(117);
    layer0_outputs(10867) <= not((inputs(104)) or (inputs(119)));
    layer0_outputs(10868) <= not((inputs(73)) and (inputs(145)));
    layer0_outputs(10869) <= not((inputs(43)) xor (inputs(197)));
    layer0_outputs(10870) <= not(inputs(203));
    layer0_outputs(10871) <= (inputs(228)) and not (inputs(119));
    layer0_outputs(10872) <= (inputs(57)) and (inputs(155));
    layer0_outputs(10873) <= inputs(182);
    layer0_outputs(10874) <= not(inputs(162));
    layer0_outputs(10875) <= not((inputs(14)) xor (inputs(124)));
    layer0_outputs(10876) <= inputs(23);
    layer0_outputs(10877) <= not(inputs(59));
    layer0_outputs(10878) <= not(inputs(89)) or (inputs(92));
    layer0_outputs(10879) <= not((inputs(105)) and (inputs(217)));
    layer0_outputs(10880) <= not(inputs(242));
    layer0_outputs(10881) <= not(inputs(127)) or (inputs(21));
    layer0_outputs(10882) <= (inputs(42)) and not (inputs(210));
    layer0_outputs(10883) <= not(inputs(164)) or (inputs(48));
    layer0_outputs(10884) <= inputs(54);
    layer0_outputs(10885) <= '0';
    layer0_outputs(10886) <= inputs(245);
    layer0_outputs(10887) <= not((inputs(212)) or (inputs(250)));
    layer0_outputs(10888) <= inputs(23);
    layer0_outputs(10889) <= (inputs(141)) xor (inputs(90));
    layer0_outputs(10890) <= not(inputs(152)) or (inputs(120));
    layer0_outputs(10891) <= (inputs(148)) and (inputs(97));
    layer0_outputs(10892) <= not(inputs(116));
    layer0_outputs(10893) <= not(inputs(103)) or (inputs(20));
    layer0_outputs(10894) <= inputs(89);
    layer0_outputs(10895) <= '1';
    layer0_outputs(10896) <= not(inputs(11)) or (inputs(2));
    layer0_outputs(10897) <= not(inputs(235)) or (inputs(199));
    layer0_outputs(10898) <= not(inputs(164));
    layer0_outputs(10899) <= not(inputs(141)) or (inputs(167));
    layer0_outputs(10900) <= (inputs(61)) and not (inputs(201));
    layer0_outputs(10901) <= (inputs(121)) or (inputs(137));
    layer0_outputs(10902) <= (inputs(27)) and not (inputs(150));
    layer0_outputs(10903) <= (inputs(126)) and not (inputs(50));
    layer0_outputs(10904) <= '0';
    layer0_outputs(10905) <= inputs(180);
    layer0_outputs(10906) <= inputs(194);
    layer0_outputs(10907) <= not(inputs(139));
    layer0_outputs(10908) <= not(inputs(171)) or (inputs(104));
    layer0_outputs(10909) <= inputs(223);
    layer0_outputs(10910) <= inputs(48);
    layer0_outputs(10911) <= '1';
    layer0_outputs(10912) <= (inputs(170)) xor (inputs(135));
    layer0_outputs(10913) <= not(inputs(89)) or (inputs(62));
    layer0_outputs(10914) <= not((inputs(138)) or (inputs(123)));
    layer0_outputs(10915) <= (inputs(89)) or (inputs(31));
    layer0_outputs(10916) <= not(inputs(86));
    layer0_outputs(10917) <= (inputs(254)) or (inputs(155));
    layer0_outputs(10918) <= not(inputs(240)) or (inputs(100));
    layer0_outputs(10919) <= not((inputs(189)) or (inputs(192)));
    layer0_outputs(10920) <= not((inputs(233)) or (inputs(245)));
    layer0_outputs(10921) <= (inputs(230)) xor (inputs(199));
    layer0_outputs(10922) <= not((inputs(138)) or (inputs(252)));
    layer0_outputs(10923) <= (inputs(239)) or (inputs(69));
    layer0_outputs(10924) <= (inputs(199)) or (inputs(213));
    layer0_outputs(10925) <= not((inputs(127)) or (inputs(166)));
    layer0_outputs(10926) <= not(inputs(236));
    layer0_outputs(10927) <= (inputs(104)) xor (inputs(174));
    layer0_outputs(10928) <= (inputs(105)) and not (inputs(69));
    layer0_outputs(10929) <= (inputs(64)) and not (inputs(107));
    layer0_outputs(10930) <= inputs(81);
    layer0_outputs(10931) <= (inputs(127)) or (inputs(46));
    layer0_outputs(10932) <= (inputs(32)) and not (inputs(79));
    layer0_outputs(10933) <= not(inputs(34)) or (inputs(6));
    layer0_outputs(10934) <= (inputs(39)) and not (inputs(120));
    layer0_outputs(10935) <= (inputs(205)) xor (inputs(126));
    layer0_outputs(10936) <= (inputs(208)) or (inputs(170));
    layer0_outputs(10937) <= not(inputs(127)) or (inputs(223));
    layer0_outputs(10938) <= not((inputs(222)) xor (inputs(22)));
    layer0_outputs(10939) <= inputs(125);
    layer0_outputs(10940) <= inputs(200);
    layer0_outputs(10941) <= '1';
    layer0_outputs(10942) <= not(inputs(255));
    layer0_outputs(10943) <= (inputs(8)) xor (inputs(144));
    layer0_outputs(10944) <= not((inputs(224)) or (inputs(40)));
    layer0_outputs(10945) <= (inputs(156)) xor (inputs(65));
    layer0_outputs(10946) <= (inputs(48)) xor (inputs(204));
    layer0_outputs(10947) <= not((inputs(34)) xor (inputs(196)));
    layer0_outputs(10948) <= (inputs(184)) and not (inputs(195));
    layer0_outputs(10949) <= not((inputs(252)) or (inputs(160)));
    layer0_outputs(10950) <= inputs(247);
    layer0_outputs(10951) <= inputs(231);
    layer0_outputs(10952) <= not(inputs(183)) or (inputs(228));
    layer0_outputs(10953) <= '1';
    layer0_outputs(10954) <= not((inputs(67)) xor (inputs(102)));
    layer0_outputs(10955) <= (inputs(83)) or (inputs(182));
    layer0_outputs(10956) <= (inputs(223)) xor (inputs(17));
    layer0_outputs(10957) <= '1';
    layer0_outputs(10958) <= not((inputs(1)) or (inputs(109)));
    layer0_outputs(10959) <= inputs(129);
    layer0_outputs(10960) <= not(inputs(148)) or (inputs(89));
    layer0_outputs(10961) <= (inputs(162)) or (inputs(113));
    layer0_outputs(10962) <= not((inputs(94)) or (inputs(117)));
    layer0_outputs(10963) <= inputs(246);
    layer0_outputs(10964) <= inputs(60);
    layer0_outputs(10965) <= (inputs(68)) and not (inputs(39));
    layer0_outputs(10966) <= not(inputs(161));
    layer0_outputs(10967) <= not((inputs(181)) or (inputs(75)));
    layer0_outputs(10968) <= not(inputs(135)) or (inputs(47));
    layer0_outputs(10969) <= (inputs(184)) or (inputs(178));
    layer0_outputs(10970) <= not(inputs(62)) or (inputs(76));
    layer0_outputs(10971) <= not((inputs(15)) or (inputs(199)));
    layer0_outputs(10972) <= (inputs(20)) xor (inputs(140));
    layer0_outputs(10973) <= not((inputs(7)) or (inputs(224)));
    layer0_outputs(10974) <= not(inputs(167)) or (inputs(154));
    layer0_outputs(10975) <= not(inputs(80)) or (inputs(2));
    layer0_outputs(10976) <= (inputs(165)) xor (inputs(148));
    layer0_outputs(10977) <= inputs(137);
    layer0_outputs(10978) <= not(inputs(176));
    layer0_outputs(10979) <= not(inputs(168));
    layer0_outputs(10980) <= inputs(164);
    layer0_outputs(10981) <= (inputs(15)) or (inputs(141));
    layer0_outputs(10982) <= inputs(190);
    layer0_outputs(10983) <= not(inputs(179));
    layer0_outputs(10984) <= not((inputs(157)) xor (inputs(25)));
    layer0_outputs(10985) <= not((inputs(80)) or (inputs(192)));
    layer0_outputs(10986) <= not(inputs(56)) or (inputs(26));
    layer0_outputs(10987) <= not(inputs(128));
    layer0_outputs(10988) <= not(inputs(168)) or (inputs(108));
    layer0_outputs(10989) <= not((inputs(233)) xor (inputs(14)));
    layer0_outputs(10990) <= (inputs(208)) xor (inputs(188));
    layer0_outputs(10991) <= not(inputs(254)) or (inputs(40));
    layer0_outputs(10992) <= inputs(37);
    layer0_outputs(10993) <= not((inputs(122)) xor (inputs(153)));
    layer0_outputs(10994) <= inputs(182);
    layer0_outputs(10995) <= (inputs(166)) and (inputs(115));
    layer0_outputs(10996) <= not(inputs(149)) or (inputs(224));
    layer0_outputs(10997) <= (inputs(203)) and not (inputs(158));
    layer0_outputs(10998) <= inputs(26);
    layer0_outputs(10999) <= not(inputs(8)) or (inputs(213));
    layer0_outputs(11000) <= not(inputs(43)) or (inputs(105));
    layer0_outputs(11001) <= (inputs(46)) and (inputs(159));
    layer0_outputs(11002) <= (inputs(111)) and not (inputs(2));
    layer0_outputs(11003) <= (inputs(6)) xor (inputs(53));
    layer0_outputs(11004) <= not(inputs(52));
    layer0_outputs(11005) <= not((inputs(134)) or (inputs(151)));
    layer0_outputs(11006) <= not(inputs(77)) or (inputs(255));
    layer0_outputs(11007) <= not(inputs(71));
    layer0_outputs(11008) <= not(inputs(17)) or (inputs(83));
    layer0_outputs(11009) <= not(inputs(59));
    layer0_outputs(11010) <= not(inputs(10)) or (inputs(237));
    layer0_outputs(11011) <= (inputs(136)) and not (inputs(30));
    layer0_outputs(11012) <= not(inputs(145));
    layer0_outputs(11013) <= inputs(232);
    layer0_outputs(11014) <= not(inputs(227));
    layer0_outputs(11015) <= (inputs(195)) and not (inputs(137));
    layer0_outputs(11016) <= not(inputs(129));
    layer0_outputs(11017) <= not(inputs(214));
    layer0_outputs(11018) <= not(inputs(232));
    layer0_outputs(11019) <= not((inputs(141)) xor (inputs(250)));
    layer0_outputs(11020) <= inputs(74);
    layer0_outputs(11021) <= not((inputs(158)) or (inputs(156)));
    layer0_outputs(11022) <= not((inputs(66)) or (inputs(79)));
    layer0_outputs(11023) <= (inputs(236)) xor (inputs(181));
    layer0_outputs(11024) <= (inputs(12)) or (inputs(6));
    layer0_outputs(11025) <= not(inputs(190));
    layer0_outputs(11026) <= not(inputs(67));
    layer0_outputs(11027) <= not(inputs(218)) or (inputs(110));
    layer0_outputs(11028) <= (inputs(45)) and not (inputs(251));
    layer0_outputs(11029) <= not((inputs(182)) and (inputs(29)));
    layer0_outputs(11030) <= not((inputs(163)) xor (inputs(117)));
    layer0_outputs(11031) <= (inputs(219)) xor (inputs(211));
    layer0_outputs(11032) <= inputs(24);
    layer0_outputs(11033) <= (inputs(104)) and not (inputs(124));
    layer0_outputs(11034) <= (inputs(208)) xor (inputs(176));
    layer0_outputs(11035) <= not((inputs(47)) or (inputs(250)));
    layer0_outputs(11036) <= '1';
    layer0_outputs(11037) <= inputs(82);
    layer0_outputs(11038) <= not((inputs(124)) xor (inputs(52)));
    layer0_outputs(11039) <= not(inputs(151)) or (inputs(115));
    layer0_outputs(11040) <= not((inputs(81)) xor (inputs(26)));
    layer0_outputs(11041) <= not(inputs(44));
    layer0_outputs(11042) <= (inputs(151)) and not (inputs(44));
    layer0_outputs(11043) <= inputs(246);
    layer0_outputs(11044) <= (inputs(223)) or (inputs(15));
    layer0_outputs(11045) <= (inputs(4)) xor (inputs(222));
    layer0_outputs(11046) <= inputs(87);
    layer0_outputs(11047) <= not(inputs(103));
    layer0_outputs(11048) <= not(inputs(218)) or (inputs(58));
    layer0_outputs(11049) <= (inputs(85)) or (inputs(15));
    layer0_outputs(11050) <= (inputs(26)) and (inputs(31));
    layer0_outputs(11051) <= not(inputs(104));
    layer0_outputs(11052) <= not((inputs(143)) xor (inputs(73)));
    layer0_outputs(11053) <= not((inputs(84)) xor (inputs(30)));
    layer0_outputs(11054) <= (inputs(197)) and not (inputs(82));
    layer0_outputs(11055) <= (inputs(202)) xor (inputs(218));
    layer0_outputs(11056) <= (inputs(98)) and (inputs(107));
    layer0_outputs(11057) <= not((inputs(70)) and (inputs(117)));
    layer0_outputs(11058) <= not((inputs(94)) xor (inputs(27)));
    layer0_outputs(11059) <= (inputs(212)) or (inputs(97));
    layer0_outputs(11060) <= (inputs(230)) xor (inputs(52));
    layer0_outputs(11061) <= not(inputs(209)) or (inputs(100));
    layer0_outputs(11062) <= not(inputs(198)) or (inputs(164));
    layer0_outputs(11063) <= '0';
    layer0_outputs(11064) <= inputs(18);
    layer0_outputs(11065) <= not(inputs(169)) or (inputs(244));
    layer0_outputs(11066) <= not(inputs(90));
    layer0_outputs(11067) <= not((inputs(153)) and (inputs(231)));
    layer0_outputs(11068) <= not(inputs(228));
    layer0_outputs(11069) <= (inputs(44)) or (inputs(52));
    layer0_outputs(11070) <= not(inputs(136)) or (inputs(60));
    layer0_outputs(11071) <= not(inputs(25));
    layer0_outputs(11072) <= inputs(42);
    layer0_outputs(11073) <= (inputs(120)) and not (inputs(129));
    layer0_outputs(11074) <= (inputs(63)) and not (inputs(241));
    layer0_outputs(11075) <= (inputs(40)) and not (inputs(160));
    layer0_outputs(11076) <= (inputs(127)) or (inputs(97));
    layer0_outputs(11077) <= (inputs(143)) xor (inputs(247));
    layer0_outputs(11078) <= inputs(53);
    layer0_outputs(11079) <= (inputs(164)) and not (inputs(170));
    layer0_outputs(11080) <= (inputs(249)) and not (inputs(40));
    layer0_outputs(11081) <= inputs(241);
    layer0_outputs(11082) <= inputs(108);
    layer0_outputs(11083) <= (inputs(153)) and not (inputs(27));
    layer0_outputs(11084) <= not(inputs(231));
    layer0_outputs(11085) <= not(inputs(142));
    layer0_outputs(11086) <= not(inputs(87));
    layer0_outputs(11087) <= not(inputs(173)) or (inputs(32));
    layer0_outputs(11088) <= inputs(176);
    layer0_outputs(11089) <= not((inputs(50)) or (inputs(148)));
    layer0_outputs(11090) <= not(inputs(151));
    layer0_outputs(11091) <= (inputs(38)) and not (inputs(241));
    layer0_outputs(11092) <= not((inputs(102)) and (inputs(79)));
    layer0_outputs(11093) <= (inputs(65)) and (inputs(10));
    layer0_outputs(11094) <= not(inputs(207));
    layer0_outputs(11095) <= not((inputs(163)) or (inputs(218)));
    layer0_outputs(11096) <= not(inputs(37));
    layer0_outputs(11097) <= not(inputs(35));
    layer0_outputs(11098) <= not(inputs(147));
    layer0_outputs(11099) <= inputs(170);
    layer0_outputs(11100) <= not((inputs(5)) xor (inputs(236)));
    layer0_outputs(11101) <= not((inputs(171)) xor (inputs(132)));
    layer0_outputs(11102) <= not(inputs(115)) or (inputs(109));
    layer0_outputs(11103) <= inputs(59);
    layer0_outputs(11104) <= not((inputs(209)) and (inputs(34)));
    layer0_outputs(11105) <= (inputs(16)) xor (inputs(143));
    layer0_outputs(11106) <= (inputs(17)) and not (inputs(119));
    layer0_outputs(11107) <= not((inputs(185)) xor (inputs(101)));
    layer0_outputs(11108) <= not(inputs(100)) or (inputs(191));
    layer0_outputs(11109) <= inputs(198);
    layer0_outputs(11110) <= (inputs(110)) and not (inputs(106));
    layer0_outputs(11111) <= (inputs(181)) and not (inputs(226));
    layer0_outputs(11112) <= inputs(151);
    layer0_outputs(11113) <= inputs(120);
    layer0_outputs(11114) <= not(inputs(152));
    layer0_outputs(11115) <= not(inputs(1)) or (inputs(242));
    layer0_outputs(11116) <= inputs(36);
    layer0_outputs(11117) <= '0';
    layer0_outputs(11118) <= '1';
    layer0_outputs(11119) <= not(inputs(2)) or (inputs(239));
    layer0_outputs(11120) <= not((inputs(221)) and (inputs(197)));
    layer0_outputs(11121) <= not(inputs(88));
    layer0_outputs(11122) <= not(inputs(153));
    layer0_outputs(11123) <= not(inputs(35)) or (inputs(104));
    layer0_outputs(11124) <= (inputs(103)) and not (inputs(34));
    layer0_outputs(11125) <= inputs(51);
    layer0_outputs(11126) <= '1';
    layer0_outputs(11127) <= not(inputs(90));
    layer0_outputs(11128) <= (inputs(178)) or (inputs(136));
    layer0_outputs(11129) <= '0';
    layer0_outputs(11130) <= not(inputs(33));
    layer0_outputs(11131) <= not((inputs(107)) xor (inputs(177)));
    layer0_outputs(11132) <= (inputs(96)) and not (inputs(178));
    layer0_outputs(11133) <= not(inputs(190)) or (inputs(111));
    layer0_outputs(11134) <= not((inputs(111)) or (inputs(157)));
    layer0_outputs(11135) <= not(inputs(60)) or (inputs(210));
    layer0_outputs(11136) <= not(inputs(229));
    layer0_outputs(11137) <= not((inputs(221)) xor (inputs(106)));
    layer0_outputs(11138) <= inputs(203);
    layer0_outputs(11139) <= not(inputs(25));
    layer0_outputs(11140) <= inputs(105);
    layer0_outputs(11141) <= inputs(0);
    layer0_outputs(11142) <= not((inputs(66)) or (inputs(201)));
    layer0_outputs(11143) <= not((inputs(135)) xor (inputs(134)));
    layer0_outputs(11144) <= inputs(114);
    layer0_outputs(11145) <= not(inputs(25)) or (inputs(181));
    layer0_outputs(11146) <= not(inputs(154)) or (inputs(195));
    layer0_outputs(11147) <= (inputs(120)) and not (inputs(30));
    layer0_outputs(11148) <= not((inputs(135)) xor (inputs(138)));
    layer0_outputs(11149) <= not((inputs(67)) or (inputs(18)));
    layer0_outputs(11150) <= not(inputs(183)) or (inputs(96));
    layer0_outputs(11151) <= not((inputs(128)) xor (inputs(160)));
    layer0_outputs(11152) <= (inputs(10)) xor (inputs(55));
    layer0_outputs(11153) <= (inputs(29)) and not (inputs(193));
    layer0_outputs(11154) <= (inputs(51)) or (inputs(220));
    layer0_outputs(11155) <= not(inputs(173)) or (inputs(207));
    layer0_outputs(11156) <= (inputs(83)) or (inputs(9));
    layer0_outputs(11157) <= (inputs(186)) and not (inputs(18));
    layer0_outputs(11158) <= inputs(46);
    layer0_outputs(11159) <= not(inputs(118));
    layer0_outputs(11160) <= not(inputs(105)) or (inputs(108));
    layer0_outputs(11161) <= (inputs(30)) and not (inputs(153));
    layer0_outputs(11162) <= (inputs(126)) and not (inputs(156));
    layer0_outputs(11163) <= not(inputs(245));
    layer0_outputs(11164) <= (inputs(13)) xor (inputs(12));
    layer0_outputs(11165) <= not((inputs(111)) or (inputs(176)));
    layer0_outputs(11166) <= not(inputs(198)) or (inputs(113));
    layer0_outputs(11167) <= not(inputs(29));
    layer0_outputs(11168) <= not((inputs(148)) or (inputs(38)));
    layer0_outputs(11169) <= not((inputs(170)) or (inputs(138)));
    layer0_outputs(11170) <= (inputs(85)) and not (inputs(191));
    layer0_outputs(11171) <= (inputs(130)) or (inputs(195));
    layer0_outputs(11172) <= inputs(56);
    layer0_outputs(11173) <= not((inputs(132)) or (inputs(94)));
    layer0_outputs(11174) <= inputs(149);
    layer0_outputs(11175) <= '1';
    layer0_outputs(11176) <= (inputs(183)) or (inputs(176));
    layer0_outputs(11177) <= (inputs(165)) or (inputs(116));
    layer0_outputs(11178) <= not((inputs(163)) xor (inputs(242)));
    layer0_outputs(11179) <= not((inputs(68)) or (inputs(174)));
    layer0_outputs(11180) <= inputs(104);
    layer0_outputs(11181) <= not(inputs(196)) or (inputs(55));
    layer0_outputs(11182) <= not(inputs(115)) or (inputs(79));
    layer0_outputs(11183) <= (inputs(184)) or (inputs(255));
    layer0_outputs(11184) <= (inputs(88)) xor (inputs(161));
    layer0_outputs(11185) <= inputs(115);
    layer0_outputs(11186) <= not(inputs(198)) or (inputs(1));
    layer0_outputs(11187) <= not((inputs(219)) xor (inputs(143)));
    layer0_outputs(11188) <= (inputs(119)) xor (inputs(212));
    layer0_outputs(11189) <= '0';
    layer0_outputs(11190) <= (inputs(87)) and not (inputs(183));
    layer0_outputs(11191) <= not((inputs(178)) xor (inputs(82)));
    layer0_outputs(11192) <= inputs(110);
    layer0_outputs(11193) <= not((inputs(195)) xor (inputs(234)));
    layer0_outputs(11194) <= not(inputs(22)) or (inputs(147));
    layer0_outputs(11195) <= not(inputs(43)) or (inputs(48));
    layer0_outputs(11196) <= (inputs(170)) or (inputs(201));
    layer0_outputs(11197) <= inputs(89);
    layer0_outputs(11198) <= not(inputs(27)) or (inputs(195));
    layer0_outputs(11199) <= not((inputs(232)) and (inputs(235)));
    layer0_outputs(11200) <= not(inputs(186));
    layer0_outputs(11201) <= not(inputs(118));
    layer0_outputs(11202) <= not((inputs(219)) or (inputs(252)));
    layer0_outputs(11203) <= not(inputs(132));
    layer0_outputs(11204) <= '0';
    layer0_outputs(11205) <= not(inputs(53));
    layer0_outputs(11206) <= inputs(199);
    layer0_outputs(11207) <= not((inputs(96)) or (inputs(192)));
    layer0_outputs(11208) <= inputs(147);
    layer0_outputs(11209) <= '0';
    layer0_outputs(11210) <= not(inputs(181)) or (inputs(28));
    layer0_outputs(11211) <= not(inputs(173)) or (inputs(41));
    layer0_outputs(11212) <= (inputs(230)) xor (inputs(208));
    layer0_outputs(11213) <= not((inputs(234)) and (inputs(252)));
    layer0_outputs(11214) <= (inputs(85)) xor (inputs(236));
    layer0_outputs(11215) <= inputs(173);
    layer0_outputs(11216) <= not((inputs(20)) or (inputs(63)));
    layer0_outputs(11217) <= (inputs(152)) xor (inputs(185));
    layer0_outputs(11218) <= inputs(221);
    layer0_outputs(11219) <= not(inputs(59));
    layer0_outputs(11220) <= inputs(139);
    layer0_outputs(11221) <= (inputs(135)) and not (inputs(161));
    layer0_outputs(11222) <= not(inputs(151)) or (inputs(65));
    layer0_outputs(11223) <= not(inputs(76)) or (inputs(0));
    layer0_outputs(11224) <= not(inputs(193));
    layer0_outputs(11225) <= inputs(82);
    layer0_outputs(11226) <= (inputs(245)) and (inputs(20));
    layer0_outputs(11227) <= not(inputs(180));
    layer0_outputs(11228) <= not(inputs(61));
    layer0_outputs(11229) <= inputs(150);
    layer0_outputs(11230) <= '1';
    layer0_outputs(11231) <= not(inputs(182));
    layer0_outputs(11232) <= not(inputs(205)) or (inputs(200));
    layer0_outputs(11233) <= (inputs(139)) and not (inputs(242));
    layer0_outputs(11234) <= not((inputs(208)) xor (inputs(43)));
    layer0_outputs(11235) <= inputs(86);
    layer0_outputs(11236) <= not(inputs(39)) or (inputs(72));
    layer0_outputs(11237) <= (inputs(129)) and not (inputs(13));
    layer0_outputs(11238) <= '1';
    layer0_outputs(11239) <= inputs(177);
    layer0_outputs(11240) <= inputs(21);
    layer0_outputs(11241) <= '0';
    layer0_outputs(11242) <= '0';
    layer0_outputs(11243) <= inputs(84);
    layer0_outputs(11244) <= inputs(36);
    layer0_outputs(11245) <= not((inputs(115)) or (inputs(78)));
    layer0_outputs(11246) <= not((inputs(62)) or (inputs(146)));
    layer0_outputs(11247) <= (inputs(158)) xor (inputs(155));
    layer0_outputs(11248) <= (inputs(72)) and not (inputs(110));
    layer0_outputs(11249) <= '1';
    layer0_outputs(11250) <= inputs(239);
    layer0_outputs(11251) <= inputs(92);
    layer0_outputs(11252) <= not(inputs(97));
    layer0_outputs(11253) <= not(inputs(71)) or (inputs(0));
    layer0_outputs(11254) <= not(inputs(163)) or (inputs(45));
    layer0_outputs(11255) <= not(inputs(79)) or (inputs(236));
    layer0_outputs(11256) <= (inputs(234)) and not (inputs(128));
    layer0_outputs(11257) <= (inputs(100)) or (inputs(35));
    layer0_outputs(11258) <= (inputs(93)) or (inputs(27));
    layer0_outputs(11259) <= not((inputs(236)) or (inputs(49)));
    layer0_outputs(11260) <= inputs(185);
    layer0_outputs(11261) <= not(inputs(59)) or (inputs(209));
    layer0_outputs(11262) <= not(inputs(216)) or (inputs(141));
    layer0_outputs(11263) <= (inputs(168)) and not (inputs(88));
    layer0_outputs(11264) <= not(inputs(231)) or (inputs(73));
    layer0_outputs(11265) <= inputs(115);
    layer0_outputs(11266) <= not((inputs(140)) xor (inputs(156)));
    layer0_outputs(11267) <= not((inputs(134)) or (inputs(131)));
    layer0_outputs(11268) <= not((inputs(115)) and (inputs(0)));
    layer0_outputs(11269) <= not(inputs(58));
    layer0_outputs(11270) <= (inputs(11)) xor (inputs(202));
    layer0_outputs(11271) <= (inputs(122)) and not (inputs(54));
    layer0_outputs(11272) <= (inputs(172)) and not (inputs(153));
    layer0_outputs(11273) <= not(inputs(85));
    layer0_outputs(11274) <= (inputs(230)) or (inputs(65));
    layer0_outputs(11275) <= not(inputs(255));
    layer0_outputs(11276) <= not((inputs(221)) or (inputs(207)));
    layer0_outputs(11277) <= not((inputs(29)) or (inputs(69)));
    layer0_outputs(11278) <= (inputs(232)) and not (inputs(103));
    layer0_outputs(11279) <= (inputs(156)) and (inputs(185));
    layer0_outputs(11280) <= not(inputs(48));
    layer0_outputs(11281) <= (inputs(204)) xor (inputs(69));
    layer0_outputs(11282) <= not((inputs(228)) and (inputs(210)));
    layer0_outputs(11283) <= not(inputs(87));
    layer0_outputs(11284) <= (inputs(218)) xor (inputs(82));
    layer0_outputs(11285) <= inputs(216);
    layer0_outputs(11286) <= not(inputs(81));
    layer0_outputs(11287) <= not(inputs(208)) or (inputs(1));
    layer0_outputs(11288) <= not(inputs(111));
    layer0_outputs(11289) <= not(inputs(181));
    layer0_outputs(11290) <= (inputs(123)) and not (inputs(9));
    layer0_outputs(11291) <= not(inputs(58));
    layer0_outputs(11292) <= '1';
    layer0_outputs(11293) <= (inputs(74)) and not (inputs(251));
    layer0_outputs(11294) <= inputs(88);
    layer0_outputs(11295) <= (inputs(179)) xor (inputs(177));
    layer0_outputs(11296) <= inputs(25);
    layer0_outputs(11297) <= not(inputs(222));
    layer0_outputs(11298) <= not((inputs(160)) or (inputs(140)));
    layer0_outputs(11299) <= (inputs(219)) xor (inputs(156));
    layer0_outputs(11300) <= not(inputs(218)) or (inputs(27));
    layer0_outputs(11301) <= not(inputs(158)) or (inputs(97));
    layer0_outputs(11302) <= (inputs(116)) and not (inputs(221));
    layer0_outputs(11303) <= not(inputs(28)) or (inputs(235));
    layer0_outputs(11304) <= not((inputs(146)) or (inputs(127)));
    layer0_outputs(11305) <= inputs(110);
    layer0_outputs(11306) <= not((inputs(69)) or (inputs(56)));
    layer0_outputs(11307) <= (inputs(121)) xor (inputs(11));
    layer0_outputs(11308) <= not(inputs(134));
    layer0_outputs(11309) <= inputs(105);
    layer0_outputs(11310) <= inputs(137);
    layer0_outputs(11311) <= not(inputs(94)) or (inputs(134));
    layer0_outputs(11312) <= (inputs(178)) xor (inputs(22));
    layer0_outputs(11313) <= (inputs(157)) or (inputs(100));
    layer0_outputs(11314) <= not(inputs(207));
    layer0_outputs(11315) <= (inputs(146)) or (inputs(145));
    layer0_outputs(11316) <= not((inputs(248)) or (inputs(247)));
    layer0_outputs(11317) <= inputs(120);
    layer0_outputs(11318) <= (inputs(10)) xor (inputs(100));
    layer0_outputs(11319) <= not((inputs(65)) xor (inputs(54)));
    layer0_outputs(11320) <= not(inputs(198)) or (inputs(214));
    layer0_outputs(11321) <= (inputs(105)) and not (inputs(69));
    layer0_outputs(11322) <= not(inputs(48));
    layer0_outputs(11323) <= not(inputs(136)) or (inputs(190));
    layer0_outputs(11324) <= (inputs(42)) and not (inputs(209));
    layer0_outputs(11325) <= (inputs(244)) and (inputs(155));
    layer0_outputs(11326) <= (inputs(132)) or (inputs(157));
    layer0_outputs(11327) <= inputs(71);
    layer0_outputs(11328) <= inputs(182);
    layer0_outputs(11329) <= (inputs(120)) and (inputs(188));
    layer0_outputs(11330) <= not(inputs(127)) or (inputs(200));
    layer0_outputs(11331) <= not((inputs(156)) and (inputs(11)));
    layer0_outputs(11332) <= not(inputs(158)) or (inputs(213));
    layer0_outputs(11333) <= (inputs(13)) xor (inputs(90));
    layer0_outputs(11334) <= not(inputs(64));
    layer0_outputs(11335) <= not((inputs(107)) xor (inputs(189)));
    layer0_outputs(11336) <= '1';
    layer0_outputs(11337) <= (inputs(236)) or (inputs(103));
    layer0_outputs(11338) <= (inputs(144)) and not (inputs(238));
    layer0_outputs(11339) <= (inputs(136)) or (inputs(42));
    layer0_outputs(11340) <= not(inputs(155)) or (inputs(77));
    layer0_outputs(11341) <= (inputs(185)) xor (inputs(142));
    layer0_outputs(11342) <= not(inputs(99));
    layer0_outputs(11343) <= (inputs(174)) xor (inputs(179));
    layer0_outputs(11344) <= not(inputs(151));
    layer0_outputs(11345) <= not((inputs(87)) xor (inputs(101)));
    layer0_outputs(11346) <= not((inputs(185)) xor (inputs(102)));
    layer0_outputs(11347) <= not(inputs(88));
    layer0_outputs(11348) <= inputs(189);
    layer0_outputs(11349) <= (inputs(29)) and not (inputs(0));
    layer0_outputs(11350) <= not(inputs(82));
    layer0_outputs(11351) <= inputs(232);
    layer0_outputs(11352) <= (inputs(233)) or (inputs(216));
    layer0_outputs(11353) <= '0';
    layer0_outputs(11354) <= not((inputs(26)) xor (inputs(57)));
    layer0_outputs(11355) <= (inputs(222)) and not (inputs(81));
    layer0_outputs(11356) <= (inputs(72)) xor (inputs(22));
    layer0_outputs(11357) <= (inputs(89)) and not (inputs(191));
    layer0_outputs(11358) <= inputs(50);
    layer0_outputs(11359) <= (inputs(236)) and not (inputs(87));
    layer0_outputs(11360) <= '1';
    layer0_outputs(11361) <= not((inputs(236)) or (inputs(13)));
    layer0_outputs(11362) <= (inputs(21)) and not (inputs(153));
    layer0_outputs(11363) <= not(inputs(247));
    layer0_outputs(11364) <= not((inputs(214)) or (inputs(27)));
    layer0_outputs(11365) <= not((inputs(155)) or (inputs(101)));
    layer0_outputs(11366) <= (inputs(97)) or (inputs(98));
    layer0_outputs(11367) <= (inputs(46)) and not (inputs(149));
    layer0_outputs(11368) <= not((inputs(81)) or (inputs(116)));
    layer0_outputs(11369) <= inputs(178);
    layer0_outputs(11370) <= (inputs(110)) xor (inputs(90));
    layer0_outputs(11371) <= (inputs(243)) and not (inputs(144));
    layer0_outputs(11372) <= inputs(214);
    layer0_outputs(11373) <= '0';
    layer0_outputs(11374) <= (inputs(89)) and not (inputs(67));
    layer0_outputs(11375) <= not(inputs(69));
    layer0_outputs(11376) <= inputs(76);
    layer0_outputs(11377) <= not(inputs(110));
    layer0_outputs(11378) <= (inputs(207)) and not (inputs(158));
    layer0_outputs(11379) <= inputs(18);
    layer0_outputs(11380) <= (inputs(136)) xor (inputs(137));
    layer0_outputs(11381) <= (inputs(86)) and not (inputs(142));
    layer0_outputs(11382) <= inputs(130);
    layer0_outputs(11383) <= not(inputs(59)) or (inputs(254));
    layer0_outputs(11384) <= (inputs(80)) or (inputs(94));
    layer0_outputs(11385) <= (inputs(77)) or (inputs(139));
    layer0_outputs(11386) <= inputs(168);
    layer0_outputs(11387) <= (inputs(157)) and not (inputs(122));
    layer0_outputs(11388) <= (inputs(39)) or (inputs(94));
    layer0_outputs(11389) <= (inputs(38)) or (inputs(140));
    layer0_outputs(11390) <= not((inputs(210)) or (inputs(69)));
    layer0_outputs(11391) <= not((inputs(43)) xor (inputs(92)));
    layer0_outputs(11392) <= not(inputs(232)) or (inputs(6));
    layer0_outputs(11393) <= not(inputs(138));
    layer0_outputs(11394) <= not((inputs(72)) or (inputs(58)));
    layer0_outputs(11395) <= not(inputs(135));
    layer0_outputs(11396) <= not(inputs(166)) or (inputs(223));
    layer0_outputs(11397) <= (inputs(133)) and (inputs(98));
    layer0_outputs(11398) <= (inputs(25)) or (inputs(24));
    layer0_outputs(11399) <= (inputs(143)) and (inputs(149));
    layer0_outputs(11400) <= (inputs(238)) xor (inputs(169));
    layer0_outputs(11401) <= not(inputs(15));
    layer0_outputs(11402) <= (inputs(29)) xor (inputs(61));
    layer0_outputs(11403) <= not(inputs(112)) or (inputs(224));
    layer0_outputs(11404) <= not((inputs(119)) or (inputs(89)));
    layer0_outputs(11405) <= (inputs(33)) and not (inputs(255));
    layer0_outputs(11406) <= not((inputs(30)) or (inputs(4)));
    layer0_outputs(11407) <= (inputs(151)) and (inputs(197));
    layer0_outputs(11408) <= (inputs(181)) and not (inputs(112));
    layer0_outputs(11409) <= not((inputs(127)) xor (inputs(110)));
    layer0_outputs(11410) <= not((inputs(121)) xor (inputs(189)));
    layer0_outputs(11411) <= (inputs(77)) and not (inputs(253));
    layer0_outputs(11412) <= not(inputs(33));
    layer0_outputs(11413) <= not((inputs(109)) or (inputs(253)));
    layer0_outputs(11414) <= not(inputs(239)) or (inputs(14));
    layer0_outputs(11415) <= not((inputs(237)) xor (inputs(224)));
    layer0_outputs(11416) <= '0';
    layer0_outputs(11417) <= inputs(167);
    layer0_outputs(11418) <= not(inputs(108));
    layer0_outputs(11419) <= (inputs(190)) and (inputs(153));
    layer0_outputs(11420) <= not((inputs(206)) or (inputs(36)));
    layer0_outputs(11421) <= not(inputs(79)) or (inputs(65));
    layer0_outputs(11422) <= not(inputs(79));
    layer0_outputs(11423) <= inputs(172);
    layer0_outputs(11424) <= (inputs(58)) and not (inputs(231));
    layer0_outputs(11425) <= not(inputs(141));
    layer0_outputs(11426) <= not(inputs(49)) or (inputs(207));
    layer0_outputs(11427) <= inputs(147);
    layer0_outputs(11428) <= (inputs(177)) and not (inputs(26));
    layer0_outputs(11429) <= (inputs(196)) and not (inputs(77));
    layer0_outputs(11430) <= not((inputs(222)) or (inputs(77)));
    layer0_outputs(11431) <= not(inputs(193)) or (inputs(157));
    layer0_outputs(11432) <= not(inputs(11));
    layer0_outputs(11433) <= not(inputs(64)) or (inputs(5));
    layer0_outputs(11434) <= (inputs(112)) and not (inputs(65));
    layer0_outputs(11435) <= inputs(186);
    layer0_outputs(11436) <= not(inputs(238));
    layer0_outputs(11437) <= (inputs(31)) or (inputs(141));
    layer0_outputs(11438) <= (inputs(211)) xor (inputs(226));
    layer0_outputs(11439) <= inputs(72);
    layer0_outputs(11440) <= (inputs(125)) and not (inputs(173));
    layer0_outputs(11441) <= (inputs(75)) xor (inputs(159));
    layer0_outputs(11442) <= not(inputs(41));
    layer0_outputs(11443) <= (inputs(29)) and not (inputs(185));
    layer0_outputs(11444) <= not(inputs(128)) or (inputs(64));
    layer0_outputs(11445) <= (inputs(147)) or (inputs(235));
    layer0_outputs(11446) <= (inputs(6)) and (inputs(227));
    layer0_outputs(11447) <= inputs(231);
    layer0_outputs(11448) <= not(inputs(201));
    layer0_outputs(11449) <= not((inputs(134)) xor (inputs(208)));
    layer0_outputs(11450) <= not(inputs(168));
    layer0_outputs(11451) <= (inputs(173)) and (inputs(198));
    layer0_outputs(11452) <= not(inputs(184));
    layer0_outputs(11453) <= '0';
    layer0_outputs(11454) <= not((inputs(176)) or (inputs(54)));
    layer0_outputs(11455) <= (inputs(216)) or (inputs(1));
    layer0_outputs(11456) <= (inputs(90)) and not (inputs(242));
    layer0_outputs(11457) <= inputs(97);
    layer0_outputs(11458) <= not((inputs(119)) xor (inputs(73)));
    layer0_outputs(11459) <= (inputs(227)) and not (inputs(95));
    layer0_outputs(11460) <= (inputs(228)) and (inputs(84));
    layer0_outputs(11461) <= inputs(165);
    layer0_outputs(11462) <= not(inputs(254));
    layer0_outputs(11463) <= not(inputs(14));
    layer0_outputs(11464) <= not((inputs(216)) and (inputs(40)));
    layer0_outputs(11465) <= inputs(227);
    layer0_outputs(11466) <= (inputs(154)) or (inputs(29));
    layer0_outputs(11467) <= (inputs(212)) and not (inputs(251));
    layer0_outputs(11468) <= not(inputs(113)) or (inputs(244));
    layer0_outputs(11469) <= not(inputs(166));
    layer0_outputs(11470) <= (inputs(111)) and not (inputs(1));
    layer0_outputs(11471) <= '0';
    layer0_outputs(11472) <= not((inputs(176)) or (inputs(249)));
    layer0_outputs(11473) <= not((inputs(114)) or (inputs(131)));
    layer0_outputs(11474) <= not(inputs(245));
    layer0_outputs(11475) <= not((inputs(162)) or (inputs(114)));
    layer0_outputs(11476) <= not(inputs(10));
    layer0_outputs(11477) <= not(inputs(220));
    layer0_outputs(11478) <= inputs(82);
    layer0_outputs(11479) <= (inputs(70)) and not (inputs(32));
    layer0_outputs(11480) <= (inputs(130)) or (inputs(31));
    layer0_outputs(11481) <= not((inputs(153)) xor (inputs(0)));
    layer0_outputs(11482) <= not(inputs(234));
    layer0_outputs(11483) <= (inputs(146)) xor (inputs(192));
    layer0_outputs(11484) <= (inputs(227)) and not (inputs(95));
    layer0_outputs(11485) <= inputs(42);
    layer0_outputs(11486) <= not((inputs(125)) or (inputs(93)));
    layer0_outputs(11487) <= not((inputs(136)) or (inputs(240)));
    layer0_outputs(11488) <= (inputs(97)) or (inputs(4));
    layer0_outputs(11489) <= '0';
    layer0_outputs(11490) <= (inputs(130)) and not (inputs(237));
    layer0_outputs(11491) <= (inputs(195)) and not (inputs(44));
    layer0_outputs(11492) <= inputs(57);
    layer0_outputs(11493) <= (inputs(106)) and (inputs(110));
    layer0_outputs(11494) <= '1';
    layer0_outputs(11495) <= not(inputs(146));
    layer0_outputs(11496) <= not((inputs(169)) or (inputs(239)));
    layer0_outputs(11497) <= not(inputs(122)) or (inputs(3));
    layer0_outputs(11498) <= inputs(139);
    layer0_outputs(11499) <= not(inputs(15));
    layer0_outputs(11500) <= (inputs(129)) or (inputs(122));
    layer0_outputs(11501) <= (inputs(60)) and not (inputs(1));
    layer0_outputs(11502) <= not(inputs(125)) or (inputs(64));
    layer0_outputs(11503) <= inputs(122);
    layer0_outputs(11504) <= '0';
    layer0_outputs(11505) <= not((inputs(99)) xor (inputs(25)));
    layer0_outputs(11506) <= not((inputs(247)) xor (inputs(249)));
    layer0_outputs(11507) <= (inputs(150)) or (inputs(78));
    layer0_outputs(11508) <= not(inputs(223)) or (inputs(229));
    layer0_outputs(11509) <= not((inputs(51)) and (inputs(150)));
    layer0_outputs(11510) <= not(inputs(43));
    layer0_outputs(11511) <= inputs(70);
    layer0_outputs(11512) <= (inputs(111)) or (inputs(176));
    layer0_outputs(11513) <= inputs(130);
    layer0_outputs(11514) <= not((inputs(235)) xor (inputs(161)));
    layer0_outputs(11515) <= not(inputs(68));
    layer0_outputs(11516) <= '1';
    layer0_outputs(11517) <= (inputs(84)) and not (inputs(172));
    layer0_outputs(11518) <= not(inputs(177)) or (inputs(112));
    layer0_outputs(11519) <= '1';
    layer0_outputs(11520) <= not((inputs(113)) xor (inputs(70)));
    layer0_outputs(11521) <= inputs(32);
    layer0_outputs(11522) <= not((inputs(19)) or (inputs(105)));
    layer0_outputs(11523) <= not(inputs(152)) or (inputs(23));
    layer0_outputs(11524) <= (inputs(243)) and (inputs(251));
    layer0_outputs(11525) <= (inputs(81)) or (inputs(175));
    layer0_outputs(11526) <= (inputs(39)) and not (inputs(103));
    layer0_outputs(11527) <= inputs(140);
    layer0_outputs(11528) <= not(inputs(148));
    layer0_outputs(11529) <= not(inputs(75));
    layer0_outputs(11530) <= not(inputs(195));
    layer0_outputs(11531) <= not((inputs(7)) or (inputs(22)));
    layer0_outputs(11532) <= (inputs(207)) and (inputs(202));
    layer0_outputs(11533) <= inputs(39);
    layer0_outputs(11534) <= not(inputs(173)) or (inputs(185));
    layer0_outputs(11535) <= inputs(9);
    layer0_outputs(11536) <= not(inputs(23));
    layer0_outputs(11537) <= not((inputs(202)) and (inputs(92)));
    layer0_outputs(11538) <= (inputs(16)) or (inputs(166));
    layer0_outputs(11539) <= (inputs(160)) or (inputs(239));
    layer0_outputs(11540) <= not(inputs(173));
    layer0_outputs(11541) <= (inputs(211)) xor (inputs(197));
    layer0_outputs(11542) <= not(inputs(199)) or (inputs(94));
    layer0_outputs(11543) <= '1';
    layer0_outputs(11544) <= (inputs(103)) xor (inputs(26));
    layer0_outputs(11545) <= inputs(223);
    layer0_outputs(11546) <= not((inputs(252)) and (inputs(140)));
    layer0_outputs(11547) <= inputs(33);
    layer0_outputs(11548) <= not(inputs(73));
    layer0_outputs(11549) <= not((inputs(132)) and (inputs(100)));
    layer0_outputs(11550) <= (inputs(181)) and not (inputs(95));
    layer0_outputs(11551) <= not((inputs(254)) or (inputs(119)));
    layer0_outputs(11552) <= (inputs(220)) and not (inputs(46));
    layer0_outputs(11553) <= not(inputs(136));
    layer0_outputs(11554) <= (inputs(7)) xor (inputs(31));
    layer0_outputs(11555) <= inputs(232);
    layer0_outputs(11556) <= not((inputs(168)) or (inputs(126)));
    layer0_outputs(11557) <= not(inputs(174));
    layer0_outputs(11558) <= inputs(83);
    layer0_outputs(11559) <= inputs(61);
    layer0_outputs(11560) <= not((inputs(176)) xor (inputs(25)));
    layer0_outputs(11561) <= inputs(37);
    layer0_outputs(11562) <= (inputs(73)) and (inputs(239));
    layer0_outputs(11563) <= (inputs(193)) and not (inputs(139));
    layer0_outputs(11564) <= (inputs(194)) or (inputs(185));
    layer0_outputs(11565) <= '0';
    layer0_outputs(11566) <= '0';
    layer0_outputs(11567) <= not((inputs(107)) or (inputs(74)));
    layer0_outputs(11568) <= '1';
    layer0_outputs(11569) <= not((inputs(119)) or (inputs(206)));
    layer0_outputs(11570) <= not((inputs(206)) or (inputs(204)));
    layer0_outputs(11571) <= not(inputs(53)) or (inputs(76));
    layer0_outputs(11572) <= not((inputs(168)) or (inputs(225)));
    layer0_outputs(11573) <= inputs(169);
    layer0_outputs(11574) <= not(inputs(78));
    layer0_outputs(11575) <= not(inputs(202)) or (inputs(31));
    layer0_outputs(11576) <= not(inputs(232)) or (inputs(60));
    layer0_outputs(11577) <= (inputs(69)) and not (inputs(216));
    layer0_outputs(11578) <= not((inputs(136)) xor (inputs(134)));
    layer0_outputs(11579) <= inputs(25);
    layer0_outputs(11580) <= (inputs(21)) or (inputs(14));
    layer0_outputs(11581) <= inputs(138);
    layer0_outputs(11582) <= (inputs(135)) or (inputs(150));
    layer0_outputs(11583) <= not(inputs(9));
    layer0_outputs(11584) <= inputs(201);
    layer0_outputs(11585) <= (inputs(86)) or (inputs(156));
    layer0_outputs(11586) <= not(inputs(61)) or (inputs(38));
    layer0_outputs(11587) <= not((inputs(35)) xor (inputs(165)));
    layer0_outputs(11588) <= (inputs(45)) and not (inputs(51));
    layer0_outputs(11589) <= not(inputs(122));
    layer0_outputs(11590) <= not((inputs(179)) and (inputs(232)));
    layer0_outputs(11591) <= not(inputs(104));
    layer0_outputs(11592) <= not(inputs(1));
    layer0_outputs(11593) <= (inputs(166)) xor (inputs(148));
    layer0_outputs(11594) <= (inputs(206)) xor (inputs(192));
    layer0_outputs(11595) <= not((inputs(141)) xor (inputs(206)));
    layer0_outputs(11596) <= not(inputs(103));
    layer0_outputs(11597) <= not(inputs(51)) or (inputs(88));
    layer0_outputs(11598) <= inputs(113);
    layer0_outputs(11599) <= not(inputs(16));
    layer0_outputs(11600) <= (inputs(178)) xor (inputs(16));
    layer0_outputs(11601) <= not(inputs(245));
    layer0_outputs(11602) <= not(inputs(153)) or (inputs(233));
    layer0_outputs(11603) <= not(inputs(182));
    layer0_outputs(11604) <= (inputs(75)) and not (inputs(243));
    layer0_outputs(11605) <= not(inputs(126));
    layer0_outputs(11606) <= (inputs(30)) and not (inputs(114));
    layer0_outputs(11607) <= inputs(228);
    layer0_outputs(11608) <= not((inputs(176)) or (inputs(47)));
    layer0_outputs(11609) <= (inputs(130)) xor (inputs(133));
    layer0_outputs(11610) <= (inputs(46)) xor (inputs(72));
    layer0_outputs(11611) <= not(inputs(157));
    layer0_outputs(11612) <= not(inputs(34)) or (inputs(200));
    layer0_outputs(11613) <= not(inputs(247));
    layer0_outputs(11614) <= (inputs(145)) xor (inputs(32));
    layer0_outputs(11615) <= (inputs(212)) and not (inputs(31));
    layer0_outputs(11616) <= inputs(92);
    layer0_outputs(11617) <= (inputs(109)) xor (inputs(52));
    layer0_outputs(11618) <= not((inputs(6)) or (inputs(211)));
    layer0_outputs(11619) <= not(inputs(105));
    layer0_outputs(11620) <= (inputs(162)) or (inputs(68));
    layer0_outputs(11621) <= not((inputs(134)) or (inputs(185)));
    layer0_outputs(11622) <= not(inputs(80));
    layer0_outputs(11623) <= (inputs(45)) and (inputs(87));
    layer0_outputs(11624) <= not((inputs(104)) or (inputs(31)));
    layer0_outputs(11625) <= not((inputs(255)) or (inputs(168)));
    layer0_outputs(11626) <= inputs(230);
    layer0_outputs(11627) <= (inputs(212)) and not (inputs(131));
    layer0_outputs(11628) <= '0';
    layer0_outputs(11629) <= inputs(88);
    layer0_outputs(11630) <= not((inputs(193)) or (inputs(216)));
    layer0_outputs(11631) <= not(inputs(39));
    layer0_outputs(11632) <= '0';
    layer0_outputs(11633) <= inputs(170);
    layer0_outputs(11634) <= inputs(44);
    layer0_outputs(11635) <= (inputs(156)) or (inputs(23));
    layer0_outputs(11636) <= not(inputs(161));
    layer0_outputs(11637) <= (inputs(4)) and not (inputs(239));
    layer0_outputs(11638) <= (inputs(235)) or (inputs(217));
    layer0_outputs(11639) <= not(inputs(233)) or (inputs(209));
    layer0_outputs(11640) <= not(inputs(147));
    layer0_outputs(11641) <= (inputs(202)) or (inputs(188));
    layer0_outputs(11642) <= not(inputs(95));
    layer0_outputs(11643) <= (inputs(70)) and not (inputs(71));
    layer0_outputs(11644) <= (inputs(217)) xor (inputs(148));
    layer0_outputs(11645) <= (inputs(42)) and not (inputs(17));
    layer0_outputs(11646) <= (inputs(25)) and not (inputs(225));
    layer0_outputs(11647) <= not((inputs(34)) or (inputs(184)));
    layer0_outputs(11648) <= not(inputs(193)) or (inputs(239));
    layer0_outputs(11649) <= (inputs(72)) or (inputs(211));
    layer0_outputs(11650) <= not((inputs(141)) or (inputs(155)));
    layer0_outputs(11651) <= not((inputs(6)) or (inputs(91)));
    layer0_outputs(11652) <= inputs(52);
    layer0_outputs(11653) <= inputs(193);
    layer0_outputs(11654) <= (inputs(29)) xor (inputs(101));
    layer0_outputs(11655) <= not(inputs(140));
    layer0_outputs(11656) <= not(inputs(228)) or (inputs(27));
    layer0_outputs(11657) <= (inputs(26)) xor (inputs(93));
    layer0_outputs(11658) <= not(inputs(104));
    layer0_outputs(11659) <= '1';
    layer0_outputs(11660) <= not((inputs(156)) and (inputs(121)));
    layer0_outputs(11661) <= not((inputs(131)) xor (inputs(119)));
    layer0_outputs(11662) <= not(inputs(213)) or (inputs(56));
    layer0_outputs(11663) <= not(inputs(18));
    layer0_outputs(11664) <= inputs(2);
    layer0_outputs(11665) <= (inputs(38)) xor (inputs(11));
    layer0_outputs(11666) <= inputs(196);
    layer0_outputs(11667) <= (inputs(69)) xor (inputs(100));
    layer0_outputs(11668) <= inputs(53);
    layer0_outputs(11669) <= (inputs(68)) or (inputs(61));
    layer0_outputs(11670) <= not(inputs(218));
    layer0_outputs(11671) <= not(inputs(193));
    layer0_outputs(11672) <= not(inputs(238));
    layer0_outputs(11673) <= (inputs(131)) and not (inputs(32));
    layer0_outputs(11674) <= (inputs(6)) and not (inputs(180));
    layer0_outputs(11675) <= inputs(102);
    layer0_outputs(11676) <= (inputs(202)) or (inputs(112));
    layer0_outputs(11677) <= (inputs(237)) xor (inputs(136));
    layer0_outputs(11678) <= not(inputs(195));
    layer0_outputs(11679) <= not(inputs(142)) or (inputs(183));
    layer0_outputs(11680) <= not(inputs(41));
    layer0_outputs(11681) <= not(inputs(92));
    layer0_outputs(11682) <= (inputs(34)) and not (inputs(51));
    layer0_outputs(11683) <= (inputs(245)) or (inputs(89));
    layer0_outputs(11684) <= inputs(241);
    layer0_outputs(11685) <= (inputs(192)) and not (inputs(70));
    layer0_outputs(11686) <= (inputs(134)) and not (inputs(186));
    layer0_outputs(11687) <= (inputs(225)) or (inputs(225));
    layer0_outputs(11688) <= not(inputs(191)) or (inputs(113));
    layer0_outputs(11689) <= not((inputs(88)) or (inputs(106)));
    layer0_outputs(11690) <= '0';
    layer0_outputs(11691) <= not(inputs(82));
    layer0_outputs(11692) <= (inputs(220)) or (inputs(216));
    layer0_outputs(11693) <= not((inputs(246)) or (inputs(162)));
    layer0_outputs(11694) <= not((inputs(145)) or (inputs(55)));
    layer0_outputs(11695) <= inputs(24);
    layer0_outputs(11696) <= not(inputs(232));
    layer0_outputs(11697) <= not((inputs(47)) or (inputs(106)));
    layer0_outputs(11698) <= (inputs(166)) and not (inputs(21));
    layer0_outputs(11699) <= inputs(115);
    layer0_outputs(11700) <= (inputs(209)) and not (inputs(247));
    layer0_outputs(11701) <= inputs(51);
    layer0_outputs(11702) <= '1';
    layer0_outputs(11703) <= inputs(118);
    layer0_outputs(11704) <= inputs(66);
    layer0_outputs(11705) <= not(inputs(148));
    layer0_outputs(11706) <= (inputs(82)) or (inputs(108));
    layer0_outputs(11707) <= not(inputs(167));
    layer0_outputs(11708) <= not((inputs(48)) or (inputs(10)));
    layer0_outputs(11709) <= not(inputs(210));
    layer0_outputs(11710) <= (inputs(54)) and (inputs(207));
    layer0_outputs(11711) <= not(inputs(233)) or (inputs(208));
    layer0_outputs(11712) <= inputs(105);
    layer0_outputs(11713) <= not(inputs(214)) or (inputs(36));
    layer0_outputs(11714) <= not(inputs(228));
    layer0_outputs(11715) <= inputs(46);
    layer0_outputs(11716) <= not(inputs(97));
    layer0_outputs(11717) <= inputs(138);
    layer0_outputs(11718) <= not(inputs(246));
    layer0_outputs(11719) <= not((inputs(135)) or (inputs(91)));
    layer0_outputs(11720) <= inputs(31);
    layer0_outputs(11721) <= inputs(129);
    layer0_outputs(11722) <= not(inputs(182)) or (inputs(174));
    layer0_outputs(11723) <= (inputs(127)) xor (inputs(92));
    layer0_outputs(11724) <= inputs(86);
    layer0_outputs(11725) <= not((inputs(66)) xor (inputs(156)));
    layer0_outputs(11726) <= (inputs(195)) xor (inputs(28));
    layer0_outputs(11727) <= not(inputs(62));
    layer0_outputs(11728) <= inputs(63);
    layer0_outputs(11729) <= not(inputs(243)) or (inputs(3));
    layer0_outputs(11730) <= not(inputs(6)) or (inputs(85));
    layer0_outputs(11731) <= (inputs(180)) and not (inputs(142));
    layer0_outputs(11732) <= not((inputs(131)) or (inputs(152)));
    layer0_outputs(11733) <= inputs(100);
    layer0_outputs(11734) <= not(inputs(206)) or (inputs(142));
    layer0_outputs(11735) <= inputs(225);
    layer0_outputs(11736) <= not((inputs(182)) and (inputs(200)));
    layer0_outputs(11737) <= not((inputs(22)) xor (inputs(27)));
    layer0_outputs(11738) <= '1';
    layer0_outputs(11739) <= (inputs(99)) and not (inputs(163));
    layer0_outputs(11740) <= inputs(38);
    layer0_outputs(11741) <= not(inputs(90));
    layer0_outputs(11742) <= '0';
    layer0_outputs(11743) <= (inputs(135)) and not (inputs(187));
    layer0_outputs(11744) <= inputs(244);
    layer0_outputs(11745) <= (inputs(210)) and (inputs(245));
    layer0_outputs(11746) <= (inputs(205)) or (inputs(18));
    layer0_outputs(11747) <= (inputs(192)) and not (inputs(253));
    layer0_outputs(11748) <= (inputs(32)) and not (inputs(241));
    layer0_outputs(11749) <= (inputs(113)) and not (inputs(95));
    layer0_outputs(11750) <= not(inputs(200)) or (inputs(244));
    layer0_outputs(11751) <= not(inputs(218));
    layer0_outputs(11752) <= (inputs(181)) and not (inputs(124));
    layer0_outputs(11753) <= not((inputs(220)) and (inputs(218)));
    layer0_outputs(11754) <= inputs(40);
    layer0_outputs(11755) <= not((inputs(203)) or (inputs(247)));
    layer0_outputs(11756) <= inputs(27);
    layer0_outputs(11757) <= not(inputs(54));
    layer0_outputs(11758) <= not((inputs(197)) or (inputs(113)));
    layer0_outputs(11759) <= not((inputs(126)) or (inputs(228)));
    layer0_outputs(11760) <= (inputs(44)) and (inputs(39));
    layer0_outputs(11761) <= (inputs(54)) or (inputs(167));
    layer0_outputs(11762) <= (inputs(109)) or (inputs(237));
    layer0_outputs(11763) <= '1';
    layer0_outputs(11764) <= (inputs(84)) and not (inputs(58));
    layer0_outputs(11765) <= not(inputs(230)) or (inputs(14));
    layer0_outputs(11766) <= (inputs(148)) and not (inputs(52));
    layer0_outputs(11767) <= '1';
    layer0_outputs(11768) <= (inputs(44)) or (inputs(22));
    layer0_outputs(11769) <= inputs(248);
    layer0_outputs(11770) <= '1';
    layer0_outputs(11771) <= inputs(86);
    layer0_outputs(11772) <= not((inputs(163)) xor (inputs(76)));
    layer0_outputs(11773) <= (inputs(41)) xor (inputs(86));
    layer0_outputs(11774) <= (inputs(26)) and (inputs(227));
    layer0_outputs(11775) <= (inputs(135)) xor (inputs(95));
    layer0_outputs(11776) <= (inputs(203)) and (inputs(200));
    layer0_outputs(11777) <= inputs(165);
    layer0_outputs(11778) <= inputs(231);
    layer0_outputs(11779) <= inputs(198);
    layer0_outputs(11780) <= not((inputs(39)) or (inputs(64)));
    layer0_outputs(11781) <= not(inputs(194));
    layer0_outputs(11782) <= not(inputs(29));
    layer0_outputs(11783) <= not(inputs(69));
    layer0_outputs(11784) <= not(inputs(77)) or (inputs(255));
    layer0_outputs(11785) <= not((inputs(236)) or (inputs(176)));
    layer0_outputs(11786) <= '0';
    layer0_outputs(11787) <= not(inputs(26));
    layer0_outputs(11788) <= not(inputs(134));
    layer0_outputs(11789) <= (inputs(213)) xor (inputs(250));
    layer0_outputs(11790) <= inputs(203);
    layer0_outputs(11791) <= inputs(103);
    layer0_outputs(11792) <= (inputs(129)) xor (inputs(92));
    layer0_outputs(11793) <= not(inputs(227)) or (inputs(226));
    layer0_outputs(11794) <= inputs(231);
    layer0_outputs(11795) <= not(inputs(91)) or (inputs(192));
    layer0_outputs(11796) <= (inputs(30)) xor (inputs(6));
    layer0_outputs(11797) <= (inputs(29)) and (inputs(200));
    layer0_outputs(11798) <= not((inputs(240)) xor (inputs(172)));
    layer0_outputs(11799) <= inputs(113);
    layer0_outputs(11800) <= inputs(103);
    layer0_outputs(11801) <= '0';
    layer0_outputs(11802) <= not(inputs(22)) or (inputs(146));
    layer0_outputs(11803) <= (inputs(33)) and not (inputs(29));
    layer0_outputs(11804) <= (inputs(72)) xor (inputs(239));
    layer0_outputs(11805) <= inputs(230);
    layer0_outputs(11806) <= not(inputs(96)) or (inputs(122));
    layer0_outputs(11807) <= not(inputs(26)) or (inputs(205));
    layer0_outputs(11808) <= not(inputs(88));
    layer0_outputs(11809) <= not((inputs(97)) or (inputs(236)));
    layer0_outputs(11810) <= not(inputs(206));
    layer0_outputs(11811) <= (inputs(63)) or (inputs(176));
    layer0_outputs(11812) <= not(inputs(31));
    layer0_outputs(11813) <= (inputs(83)) or (inputs(221));
    layer0_outputs(11814) <= (inputs(204)) xor (inputs(207));
    layer0_outputs(11815) <= not(inputs(62));
    layer0_outputs(11816) <= (inputs(54)) or (inputs(101));
    layer0_outputs(11817) <= (inputs(39)) and (inputs(152));
    layer0_outputs(11818) <= not(inputs(219)) or (inputs(109));
    layer0_outputs(11819) <= (inputs(47)) xor (inputs(203));
    layer0_outputs(11820) <= inputs(139);
    layer0_outputs(11821) <= (inputs(218)) or (inputs(245));
    layer0_outputs(11822) <= inputs(212);
    layer0_outputs(11823) <= inputs(83);
    layer0_outputs(11824) <= '1';
    layer0_outputs(11825) <= not((inputs(124)) or (inputs(19)));
    layer0_outputs(11826) <= not(inputs(116));
    layer0_outputs(11827) <= inputs(173);
    layer0_outputs(11828) <= not(inputs(184));
    layer0_outputs(11829) <= (inputs(149)) or (inputs(52));
    layer0_outputs(11830) <= not(inputs(217)) or (inputs(5));
    layer0_outputs(11831) <= not((inputs(173)) xor (inputs(105)));
    layer0_outputs(11832) <= (inputs(170)) or (inputs(171));
    layer0_outputs(11833) <= not((inputs(105)) or (inputs(67)));
    layer0_outputs(11834) <= inputs(30);
    layer0_outputs(11835) <= inputs(216);
    layer0_outputs(11836) <= (inputs(169)) and not (inputs(62));
    layer0_outputs(11837) <= not(inputs(183));
    layer0_outputs(11838) <= not((inputs(43)) or (inputs(141)));
    layer0_outputs(11839) <= (inputs(54)) xor (inputs(41));
    layer0_outputs(11840) <= (inputs(184)) and not (inputs(88));
    layer0_outputs(11841) <= '0';
    layer0_outputs(11842) <= (inputs(233)) and not (inputs(146));
    layer0_outputs(11843) <= inputs(140);
    layer0_outputs(11844) <= not(inputs(211)) or (inputs(15));
    layer0_outputs(11845) <= not(inputs(8));
    layer0_outputs(11846) <= (inputs(185)) and not (inputs(252));
    layer0_outputs(11847) <= not(inputs(219));
    layer0_outputs(11848) <= not((inputs(16)) or (inputs(245)));
    layer0_outputs(11849) <= not(inputs(192));
    layer0_outputs(11850) <= inputs(115);
    layer0_outputs(11851) <= not((inputs(249)) or (inputs(105)));
    layer0_outputs(11852) <= not((inputs(44)) or (inputs(49)));
    layer0_outputs(11853) <= not(inputs(139)) or (inputs(98));
    layer0_outputs(11854) <= not(inputs(223));
    layer0_outputs(11855) <= '1';
    layer0_outputs(11856) <= (inputs(44)) and not (inputs(182));
    layer0_outputs(11857) <= not(inputs(32)) or (inputs(10));
    layer0_outputs(11858) <= not(inputs(78));
    layer0_outputs(11859) <= inputs(73);
    layer0_outputs(11860) <= not((inputs(144)) or (inputs(171)));
    layer0_outputs(11861) <= not(inputs(27));
    layer0_outputs(11862) <= (inputs(228)) and not (inputs(58));
    layer0_outputs(11863) <= not((inputs(191)) or (inputs(203)));
    layer0_outputs(11864) <= not(inputs(45)) or (inputs(37));
    layer0_outputs(11865) <= inputs(108);
    layer0_outputs(11866) <= inputs(122);
    layer0_outputs(11867) <= inputs(83);
    layer0_outputs(11868) <= (inputs(25)) and not (inputs(111));
    layer0_outputs(11869) <= not((inputs(197)) or (inputs(68)));
    layer0_outputs(11870) <= inputs(199);
    layer0_outputs(11871) <= not(inputs(104));
    layer0_outputs(11872) <= not((inputs(64)) or (inputs(179)));
    layer0_outputs(11873) <= not((inputs(57)) and (inputs(117)));
    layer0_outputs(11874) <= (inputs(9)) or (inputs(134));
    layer0_outputs(11875) <= inputs(83);
    layer0_outputs(11876) <= inputs(23);
    layer0_outputs(11877) <= (inputs(131)) and not (inputs(224));
    layer0_outputs(11878) <= not(inputs(101));
    layer0_outputs(11879) <= (inputs(31)) and (inputs(144));
    layer0_outputs(11880) <= not(inputs(55)) or (inputs(185));
    layer0_outputs(11881) <= (inputs(235)) or (inputs(48));
    layer0_outputs(11882) <= not(inputs(252)) or (inputs(19));
    layer0_outputs(11883) <= (inputs(135)) and not (inputs(97));
    layer0_outputs(11884) <= '0';
    layer0_outputs(11885) <= not(inputs(24));
    layer0_outputs(11886) <= not((inputs(87)) or (inputs(102)));
    layer0_outputs(11887) <= (inputs(63)) xor (inputs(27));
    layer0_outputs(11888) <= not(inputs(68)) or (inputs(170));
    layer0_outputs(11889) <= not(inputs(110));
    layer0_outputs(11890) <= not((inputs(117)) or (inputs(147)));
    layer0_outputs(11891) <= inputs(246);
    layer0_outputs(11892) <= (inputs(223)) xor (inputs(193));
    layer0_outputs(11893) <= not(inputs(105)) or (inputs(217));
    layer0_outputs(11894) <= not(inputs(3));
    layer0_outputs(11895) <= (inputs(226)) and not (inputs(238));
    layer0_outputs(11896) <= not((inputs(17)) or (inputs(121)));
    layer0_outputs(11897) <= '1';
    layer0_outputs(11898) <= inputs(17);
    layer0_outputs(11899) <= (inputs(193)) xor (inputs(255));
    layer0_outputs(11900) <= (inputs(68)) and (inputs(116));
    layer0_outputs(11901) <= not(inputs(19));
    layer0_outputs(11902) <= '1';
    layer0_outputs(11903) <= inputs(131);
    layer0_outputs(11904) <= (inputs(77)) and not (inputs(154));
    layer0_outputs(11905) <= inputs(245);
    layer0_outputs(11906) <= not(inputs(36));
    layer0_outputs(11907) <= not(inputs(164));
    layer0_outputs(11908) <= not((inputs(86)) or (inputs(240)));
    layer0_outputs(11909) <= inputs(242);
    layer0_outputs(11910) <= inputs(200);
    layer0_outputs(11911) <= not(inputs(136));
    layer0_outputs(11912) <= not((inputs(191)) xor (inputs(1)));
    layer0_outputs(11913) <= (inputs(161)) and not (inputs(197));
    layer0_outputs(11914) <= (inputs(248)) and not (inputs(231));
    layer0_outputs(11915) <= inputs(163);
    layer0_outputs(11916) <= not((inputs(95)) xor (inputs(5)));
    layer0_outputs(11917) <= (inputs(169)) or (inputs(233));
    layer0_outputs(11918) <= not((inputs(175)) xor (inputs(242)));
    layer0_outputs(11919) <= (inputs(51)) and not (inputs(177));
    layer0_outputs(11920) <= not((inputs(246)) or (inputs(159)));
    layer0_outputs(11921) <= not(inputs(28));
    layer0_outputs(11922) <= not(inputs(110));
    layer0_outputs(11923) <= inputs(214);
    layer0_outputs(11924) <= (inputs(182)) xor (inputs(46));
    layer0_outputs(11925) <= (inputs(86)) or (inputs(97));
    layer0_outputs(11926) <= not(inputs(224));
    layer0_outputs(11927) <= not(inputs(102)) or (inputs(159));
    layer0_outputs(11928) <= inputs(11);
    layer0_outputs(11929) <= inputs(155);
    layer0_outputs(11930) <= not(inputs(92)) or (inputs(226));
    layer0_outputs(11931) <= inputs(228);
    layer0_outputs(11932) <= not(inputs(44)) or (inputs(198));
    layer0_outputs(11933) <= inputs(181);
    layer0_outputs(11934) <= inputs(81);
    layer0_outputs(11935) <= not((inputs(73)) or (inputs(41)));
    layer0_outputs(11936) <= not(inputs(167));
    layer0_outputs(11937) <= not(inputs(37));
    layer0_outputs(11938) <= (inputs(248)) or (inputs(213));
    layer0_outputs(11939) <= not(inputs(7)) or (inputs(184));
    layer0_outputs(11940) <= not(inputs(121));
    layer0_outputs(11941) <= inputs(216);
    layer0_outputs(11942) <= (inputs(165)) or (inputs(222));
    layer0_outputs(11943) <= not(inputs(85));
    layer0_outputs(11944) <= not((inputs(138)) or (inputs(23)));
    layer0_outputs(11945) <= inputs(180);
    layer0_outputs(11946) <= inputs(245);
    layer0_outputs(11947) <= not((inputs(141)) and (inputs(54)));
    layer0_outputs(11948) <= not(inputs(202));
    layer0_outputs(11949) <= not(inputs(128));
    layer0_outputs(11950) <= (inputs(199)) xor (inputs(46));
    layer0_outputs(11951) <= (inputs(213)) or (inputs(167));
    layer0_outputs(11952) <= inputs(104);
    layer0_outputs(11953) <= not(inputs(145));
    layer0_outputs(11954) <= not((inputs(45)) or (inputs(156)));
    layer0_outputs(11955) <= not(inputs(190));
    layer0_outputs(11956) <= not((inputs(130)) or (inputs(155)));
    layer0_outputs(11957) <= not(inputs(129));
    layer0_outputs(11958) <= inputs(201);
    layer0_outputs(11959) <= not(inputs(181));
    layer0_outputs(11960) <= not(inputs(74));
    layer0_outputs(11961) <= inputs(121);
    layer0_outputs(11962) <= not((inputs(116)) or (inputs(22)));
    layer0_outputs(11963) <= '0';
    layer0_outputs(11964) <= not((inputs(213)) or (inputs(192)));
    layer0_outputs(11965) <= inputs(2);
    layer0_outputs(11966) <= '0';
    layer0_outputs(11967) <= (inputs(113)) or (inputs(27));
    layer0_outputs(11968) <= not((inputs(87)) xor (inputs(99)));
    layer0_outputs(11969) <= not(inputs(212)) or (inputs(43));
    layer0_outputs(11970) <= not(inputs(134));
    layer0_outputs(11971) <= (inputs(115)) and not (inputs(192));
    layer0_outputs(11972) <= not(inputs(194));
    layer0_outputs(11973) <= not(inputs(58)) or (inputs(192));
    layer0_outputs(11974) <= (inputs(83)) and not (inputs(144));
    layer0_outputs(11975) <= inputs(87);
    layer0_outputs(11976) <= inputs(159);
    layer0_outputs(11977) <= not(inputs(132));
    layer0_outputs(11978) <= inputs(152);
    layer0_outputs(11979) <= not(inputs(166)) or (inputs(179));
    layer0_outputs(11980) <= (inputs(148)) or (inputs(182));
    layer0_outputs(11981) <= not((inputs(80)) or (inputs(248)));
    layer0_outputs(11982) <= not((inputs(190)) or (inputs(190)));
    layer0_outputs(11983) <= not((inputs(2)) xor (inputs(168)));
    layer0_outputs(11984) <= not(inputs(62)) or (inputs(19));
    layer0_outputs(11985) <= inputs(87);
    layer0_outputs(11986) <= inputs(57);
    layer0_outputs(11987) <= not(inputs(108)) or (inputs(68));
    layer0_outputs(11988) <= not((inputs(187)) xor (inputs(236)));
    layer0_outputs(11989) <= not((inputs(58)) xor (inputs(26)));
    layer0_outputs(11990) <= (inputs(44)) and (inputs(50));
    layer0_outputs(11991) <= not((inputs(172)) or (inputs(243)));
    layer0_outputs(11992) <= not((inputs(3)) or (inputs(10)));
    layer0_outputs(11993) <= inputs(3);
    layer0_outputs(11994) <= not(inputs(113));
    layer0_outputs(11995) <= '0';
    layer0_outputs(11996) <= not((inputs(105)) or (inputs(184)));
    layer0_outputs(11997) <= inputs(187);
    layer0_outputs(11998) <= not(inputs(100));
    layer0_outputs(11999) <= (inputs(70)) and not (inputs(225));
    layer0_outputs(12000) <= (inputs(198)) xor (inputs(168));
    layer0_outputs(12001) <= (inputs(97)) and not (inputs(51));
    layer0_outputs(12002) <= inputs(130);
    layer0_outputs(12003) <= inputs(29);
    layer0_outputs(12004) <= (inputs(193)) and not (inputs(176));
    layer0_outputs(12005) <= (inputs(32)) or (inputs(42));
    layer0_outputs(12006) <= not((inputs(67)) or (inputs(7)));
    layer0_outputs(12007) <= not((inputs(144)) or (inputs(247)));
    layer0_outputs(12008) <= not((inputs(94)) or (inputs(84)));
    layer0_outputs(12009) <= inputs(54);
    layer0_outputs(12010) <= not(inputs(196));
    layer0_outputs(12011) <= not((inputs(89)) xor (inputs(103)));
    layer0_outputs(12012) <= not(inputs(84));
    layer0_outputs(12013) <= (inputs(85)) and not (inputs(112));
    layer0_outputs(12014) <= inputs(41);
    layer0_outputs(12015) <= not((inputs(195)) or (inputs(62)));
    layer0_outputs(12016) <= not(inputs(194));
    layer0_outputs(12017) <= (inputs(113)) and not (inputs(237));
    layer0_outputs(12018) <= not(inputs(63));
    layer0_outputs(12019) <= inputs(32);
    layer0_outputs(12020) <= not((inputs(79)) and (inputs(168)));
    layer0_outputs(12021) <= (inputs(5)) xor (inputs(143));
    layer0_outputs(12022) <= (inputs(235)) and (inputs(13));
    layer0_outputs(12023) <= not((inputs(193)) and (inputs(145)));
    layer0_outputs(12024) <= (inputs(165)) or (inputs(70));
    layer0_outputs(12025) <= inputs(86);
    layer0_outputs(12026) <= not(inputs(55));
    layer0_outputs(12027) <= (inputs(159)) xor (inputs(88));
    layer0_outputs(12028) <= inputs(194);
    layer0_outputs(12029) <= not(inputs(202)) or (inputs(0));
    layer0_outputs(12030) <= not((inputs(219)) and (inputs(82)));
    layer0_outputs(12031) <= inputs(151);
    layer0_outputs(12032) <= inputs(152);
    layer0_outputs(12033) <= not(inputs(70)) or (inputs(252));
    layer0_outputs(12034) <= (inputs(202)) and not (inputs(110));
    layer0_outputs(12035) <= inputs(237);
    layer0_outputs(12036) <= not(inputs(129));
    layer0_outputs(12037) <= (inputs(204)) or (inputs(201));
    layer0_outputs(12038) <= not(inputs(133)) or (inputs(49));
    layer0_outputs(12039) <= (inputs(57)) xor (inputs(45));
    layer0_outputs(12040) <= (inputs(132)) and not (inputs(87));
    layer0_outputs(12041) <= (inputs(244)) and not (inputs(191));
    layer0_outputs(12042) <= not((inputs(100)) or (inputs(14)));
    layer0_outputs(12043) <= (inputs(195)) xor (inputs(152));
    layer0_outputs(12044) <= '1';
    layer0_outputs(12045) <= not(inputs(59));
    layer0_outputs(12046) <= not((inputs(222)) or (inputs(168)));
    layer0_outputs(12047) <= (inputs(208)) and (inputs(50));
    layer0_outputs(12048) <= not(inputs(210)) or (inputs(20));
    layer0_outputs(12049) <= not(inputs(101));
    layer0_outputs(12050) <= inputs(92);
    layer0_outputs(12051) <= '0';
    layer0_outputs(12052) <= (inputs(18)) and (inputs(81));
    layer0_outputs(12053) <= inputs(174);
    layer0_outputs(12054) <= '0';
    layer0_outputs(12055) <= not(inputs(121));
    layer0_outputs(12056) <= not(inputs(135));
    layer0_outputs(12057) <= (inputs(201)) and not (inputs(125));
    layer0_outputs(12058) <= (inputs(37)) and not (inputs(95));
    layer0_outputs(12059) <= not(inputs(97)) or (inputs(35));
    layer0_outputs(12060) <= not((inputs(245)) or (inputs(64)));
    layer0_outputs(12061) <= (inputs(213)) and not (inputs(84));
    layer0_outputs(12062) <= not(inputs(145));
    layer0_outputs(12063) <= (inputs(219)) and (inputs(238));
    layer0_outputs(12064) <= (inputs(101)) or (inputs(159));
    layer0_outputs(12065) <= not(inputs(6));
    layer0_outputs(12066) <= inputs(105);
    layer0_outputs(12067) <= not(inputs(4));
    layer0_outputs(12068) <= inputs(231);
    layer0_outputs(12069) <= '0';
    layer0_outputs(12070) <= inputs(217);
    layer0_outputs(12071) <= not(inputs(138));
    layer0_outputs(12072) <= not(inputs(75)) or (inputs(54));
    layer0_outputs(12073) <= inputs(235);
    layer0_outputs(12074) <= (inputs(97)) xor (inputs(222));
    layer0_outputs(12075) <= not(inputs(182));
    layer0_outputs(12076) <= (inputs(183)) and not (inputs(93));
    layer0_outputs(12077) <= not(inputs(213));
    layer0_outputs(12078) <= (inputs(52)) or (inputs(185));
    layer0_outputs(12079) <= not(inputs(84));
    layer0_outputs(12080) <= not(inputs(96)) or (inputs(119));
    layer0_outputs(12081) <= not((inputs(111)) or (inputs(51)));
    layer0_outputs(12082) <= not(inputs(227)) or (inputs(142));
    layer0_outputs(12083) <= (inputs(78)) and (inputs(88));
    layer0_outputs(12084) <= not(inputs(22));
    layer0_outputs(12085) <= inputs(78);
    layer0_outputs(12086) <= inputs(98);
    layer0_outputs(12087) <= (inputs(111)) xor (inputs(222));
    layer0_outputs(12088) <= (inputs(71)) and (inputs(130));
    layer0_outputs(12089) <= not(inputs(113));
    layer0_outputs(12090) <= not((inputs(189)) xor (inputs(214)));
    layer0_outputs(12091) <= not(inputs(51)) or (inputs(248));
    layer0_outputs(12092) <= not(inputs(91)) or (inputs(132));
    layer0_outputs(12093) <= not(inputs(149));
    layer0_outputs(12094) <= (inputs(206)) or (inputs(220));
    layer0_outputs(12095) <= not(inputs(224));
    layer0_outputs(12096) <= not((inputs(192)) xor (inputs(147)));
    layer0_outputs(12097) <= inputs(195);
    layer0_outputs(12098) <= (inputs(193)) and (inputs(32));
    layer0_outputs(12099) <= not(inputs(106)) or (inputs(206));
    layer0_outputs(12100) <= (inputs(244)) and not (inputs(28));
    layer0_outputs(12101) <= not(inputs(229)) or (inputs(105));
    layer0_outputs(12102) <= (inputs(180)) or (inputs(237));
    layer0_outputs(12103) <= (inputs(70)) and not (inputs(194));
    layer0_outputs(12104) <= (inputs(57)) and not (inputs(248));
    layer0_outputs(12105) <= (inputs(248)) and (inputs(10));
    layer0_outputs(12106) <= (inputs(86)) and not (inputs(230));
    layer0_outputs(12107) <= not((inputs(159)) xor (inputs(11)));
    layer0_outputs(12108) <= not((inputs(208)) or (inputs(24)));
    layer0_outputs(12109) <= '1';
    layer0_outputs(12110) <= not(inputs(116));
    layer0_outputs(12111) <= inputs(130);
    layer0_outputs(12112) <= not(inputs(163)) or (inputs(67));
    layer0_outputs(12113) <= not(inputs(230)) or (inputs(195));
    layer0_outputs(12114) <= not((inputs(0)) or (inputs(61)));
    layer0_outputs(12115) <= inputs(180);
    layer0_outputs(12116) <= not(inputs(131));
    layer0_outputs(12117) <= not(inputs(108)) or (inputs(65));
    layer0_outputs(12118) <= not((inputs(169)) xor (inputs(137)));
    layer0_outputs(12119) <= not((inputs(100)) or (inputs(96)));
    layer0_outputs(12120) <= (inputs(7)) and not (inputs(118));
    layer0_outputs(12121) <= not(inputs(146));
    layer0_outputs(12122) <= not(inputs(122)) or (inputs(248));
    layer0_outputs(12123) <= not((inputs(124)) or (inputs(249)));
    layer0_outputs(12124) <= not(inputs(204)) or (inputs(180));
    layer0_outputs(12125) <= not(inputs(132)) or (inputs(224));
    layer0_outputs(12126) <= not(inputs(179));
    layer0_outputs(12127) <= (inputs(99)) and not (inputs(32));
    layer0_outputs(12128) <= not(inputs(141)) or (inputs(222));
    layer0_outputs(12129) <= (inputs(139)) and not (inputs(246));
    layer0_outputs(12130) <= not(inputs(132)) or (inputs(104));
    layer0_outputs(12131) <= (inputs(46)) or (inputs(32));
    layer0_outputs(12132) <= not(inputs(6));
    layer0_outputs(12133) <= not(inputs(26));
    layer0_outputs(12134) <= (inputs(117)) xor (inputs(234));
    layer0_outputs(12135) <= (inputs(252)) and (inputs(217));
    layer0_outputs(12136) <= (inputs(229)) or (inputs(5));
    layer0_outputs(12137) <= not((inputs(187)) or (inputs(113)));
    layer0_outputs(12138) <= (inputs(50)) or (inputs(221));
    layer0_outputs(12139) <= inputs(149);
    layer0_outputs(12140) <= (inputs(140)) or (inputs(3));
    layer0_outputs(12141) <= inputs(85);
    layer0_outputs(12142) <= '1';
    layer0_outputs(12143) <= not((inputs(145)) or (inputs(108)));
    layer0_outputs(12144) <= not((inputs(216)) xor (inputs(248)));
    layer0_outputs(12145) <= not(inputs(141));
    layer0_outputs(12146) <= not(inputs(163)) or (inputs(253));
    layer0_outputs(12147) <= (inputs(113)) or (inputs(246));
    layer0_outputs(12148) <= not((inputs(198)) xor (inputs(242)));
    layer0_outputs(12149) <= not(inputs(53)) or (inputs(5));
    layer0_outputs(12150) <= inputs(162);
    layer0_outputs(12151) <= (inputs(60)) and not (inputs(119));
    layer0_outputs(12152) <= (inputs(156)) or (inputs(61));
    layer0_outputs(12153) <= not(inputs(72));
    layer0_outputs(12154) <= (inputs(114)) or (inputs(78));
    layer0_outputs(12155) <= not(inputs(65));
    layer0_outputs(12156) <= not(inputs(49));
    layer0_outputs(12157) <= not((inputs(246)) or (inputs(112)));
    layer0_outputs(12158) <= '1';
    layer0_outputs(12159) <= not(inputs(167));
    layer0_outputs(12160) <= (inputs(211)) or (inputs(205));
    layer0_outputs(12161) <= not(inputs(23));
    layer0_outputs(12162) <= (inputs(45)) or (inputs(8));
    layer0_outputs(12163) <= inputs(246);
    layer0_outputs(12164) <= (inputs(2)) and (inputs(216));
    layer0_outputs(12165) <= inputs(8);
    layer0_outputs(12166) <= (inputs(227)) or (inputs(254));
    layer0_outputs(12167) <= not(inputs(59));
    layer0_outputs(12168) <= not(inputs(247));
    layer0_outputs(12169) <= not(inputs(99)) or (inputs(18));
    layer0_outputs(12170) <= not(inputs(40));
    layer0_outputs(12171) <= inputs(14);
    layer0_outputs(12172) <= not(inputs(232));
    layer0_outputs(12173) <= '0';
    layer0_outputs(12174) <= not(inputs(255));
    layer0_outputs(12175) <= not((inputs(173)) or (inputs(206)));
    layer0_outputs(12176) <= (inputs(127)) or (inputs(76));
    layer0_outputs(12177) <= not(inputs(203)) or (inputs(146));
    layer0_outputs(12178) <= (inputs(43)) and not (inputs(251));
    layer0_outputs(12179) <= inputs(25);
    layer0_outputs(12180) <= inputs(136);
    layer0_outputs(12181) <= inputs(135);
    layer0_outputs(12182) <= (inputs(127)) or (inputs(194));
    layer0_outputs(12183) <= not(inputs(158));
    layer0_outputs(12184) <= not(inputs(59)) or (inputs(19));
    layer0_outputs(12185) <= (inputs(51)) or (inputs(50));
    layer0_outputs(12186) <= (inputs(230)) and not (inputs(43));
    layer0_outputs(12187) <= not((inputs(79)) xor (inputs(88)));
    layer0_outputs(12188) <= not(inputs(52)) or (inputs(145));
    layer0_outputs(12189) <= '0';
    layer0_outputs(12190) <= (inputs(184)) or (inputs(2));
    layer0_outputs(12191) <= (inputs(211)) and not (inputs(99));
    layer0_outputs(12192) <= not(inputs(169));
    layer0_outputs(12193) <= not(inputs(200));
    layer0_outputs(12194) <= inputs(37);
    layer0_outputs(12195) <= not((inputs(145)) or (inputs(96)));
    layer0_outputs(12196) <= inputs(209);
    layer0_outputs(12197) <= not(inputs(49));
    layer0_outputs(12198) <= (inputs(9)) and not (inputs(238));
    layer0_outputs(12199) <= not(inputs(76));
    layer0_outputs(12200) <= not(inputs(46));
    layer0_outputs(12201) <= (inputs(118)) or (inputs(29));
    layer0_outputs(12202) <= '0';
    layer0_outputs(12203) <= not((inputs(203)) and (inputs(115)));
    layer0_outputs(12204) <= not(inputs(128));
    layer0_outputs(12205) <= not(inputs(118));
    layer0_outputs(12206) <= (inputs(192)) and not (inputs(60));
    layer0_outputs(12207) <= not(inputs(140)) or (inputs(50));
    layer0_outputs(12208) <= not((inputs(78)) or (inputs(61)));
    layer0_outputs(12209) <= inputs(81);
    layer0_outputs(12210) <= (inputs(213)) and not (inputs(14));
    layer0_outputs(12211) <= (inputs(151)) and not (inputs(63));
    layer0_outputs(12212) <= (inputs(182)) or (inputs(3));
    layer0_outputs(12213) <= inputs(159);
    layer0_outputs(12214) <= inputs(86);
    layer0_outputs(12215) <= inputs(9);
    layer0_outputs(12216) <= (inputs(102)) xor (inputs(20));
    layer0_outputs(12217) <= not(inputs(157)) or (inputs(238));
    layer0_outputs(12218) <= inputs(205);
    layer0_outputs(12219) <= not(inputs(166)) or (inputs(110));
    layer0_outputs(12220) <= not((inputs(29)) and (inputs(42)));
    layer0_outputs(12221) <= inputs(242);
    layer0_outputs(12222) <= (inputs(90)) and not (inputs(142));
    layer0_outputs(12223) <= (inputs(192)) and not (inputs(251));
    layer0_outputs(12224) <= not((inputs(252)) xor (inputs(161)));
    layer0_outputs(12225) <= (inputs(218)) or (inputs(205));
    layer0_outputs(12226) <= not(inputs(122));
    layer0_outputs(12227) <= not(inputs(7));
    layer0_outputs(12228) <= not(inputs(136));
    layer0_outputs(12229) <= not((inputs(242)) or (inputs(110)));
    layer0_outputs(12230) <= not((inputs(191)) and (inputs(57)));
    layer0_outputs(12231) <= (inputs(188)) or (inputs(175));
    layer0_outputs(12232) <= not((inputs(56)) or (inputs(223)));
    layer0_outputs(12233) <= not(inputs(116));
    layer0_outputs(12234) <= (inputs(119)) and not (inputs(221));
    layer0_outputs(12235) <= (inputs(55)) or (inputs(0));
    layer0_outputs(12236) <= not(inputs(47)) or (inputs(16));
    layer0_outputs(12237) <= not(inputs(21));
    layer0_outputs(12238) <= not(inputs(137));
    layer0_outputs(12239) <= not((inputs(10)) or (inputs(153)));
    layer0_outputs(12240) <= inputs(230);
    layer0_outputs(12241) <= not((inputs(16)) or (inputs(45)));
    layer0_outputs(12242) <= (inputs(100)) and not (inputs(143));
    layer0_outputs(12243) <= not(inputs(229));
    layer0_outputs(12244) <= '0';
    layer0_outputs(12245) <= inputs(93);
    layer0_outputs(12246) <= not(inputs(229)) or (inputs(109));
    layer0_outputs(12247) <= not(inputs(127));
    layer0_outputs(12248) <= not(inputs(221));
    layer0_outputs(12249) <= inputs(166);
    layer0_outputs(12250) <= (inputs(40)) and not (inputs(142));
    layer0_outputs(12251) <= not((inputs(41)) xor (inputs(59)));
    layer0_outputs(12252) <= not(inputs(153)) or (inputs(197));
    layer0_outputs(12253) <= '0';
    layer0_outputs(12254) <= not((inputs(211)) or (inputs(179)));
    layer0_outputs(12255) <= not(inputs(203));
    layer0_outputs(12256) <= (inputs(149)) xor (inputs(114));
    layer0_outputs(12257) <= inputs(90);
    layer0_outputs(12258) <= not(inputs(170));
    layer0_outputs(12259) <= (inputs(172)) and not (inputs(255));
    layer0_outputs(12260) <= (inputs(214)) or (inputs(67));
    layer0_outputs(12261) <= not(inputs(194)) or (inputs(0));
    layer0_outputs(12262) <= inputs(152);
    layer0_outputs(12263) <= (inputs(92)) and (inputs(148));
    layer0_outputs(12264) <= not(inputs(138)) or (inputs(84));
    layer0_outputs(12265) <= not((inputs(140)) or (inputs(206)));
    layer0_outputs(12266) <= not(inputs(167));
    layer0_outputs(12267) <= not(inputs(57));
    layer0_outputs(12268) <= not((inputs(24)) xor (inputs(144)));
    layer0_outputs(12269) <= inputs(134);
    layer0_outputs(12270) <= not((inputs(248)) xor (inputs(235)));
    layer0_outputs(12271) <= not((inputs(57)) and (inputs(56)));
    layer0_outputs(12272) <= (inputs(11)) xor (inputs(111));
    layer0_outputs(12273) <= (inputs(76)) or (inputs(144));
    layer0_outputs(12274) <= not((inputs(76)) xor (inputs(3)));
    layer0_outputs(12275) <= not((inputs(95)) and (inputs(43)));
    layer0_outputs(12276) <= not((inputs(184)) or (inputs(82)));
    layer0_outputs(12277) <= inputs(100);
    layer0_outputs(12278) <= not(inputs(75));
    layer0_outputs(12279) <= not(inputs(70)) or (inputs(177));
    layer0_outputs(12280) <= not((inputs(105)) or (inputs(104)));
    layer0_outputs(12281) <= (inputs(153)) or (inputs(57));
    layer0_outputs(12282) <= not((inputs(207)) or (inputs(25)));
    layer0_outputs(12283) <= not(inputs(100));
    layer0_outputs(12284) <= (inputs(44)) and not (inputs(130));
    layer0_outputs(12285) <= not((inputs(193)) or (inputs(207)));
    layer0_outputs(12286) <= '1';
    layer0_outputs(12287) <= not(inputs(78)) or (inputs(206));
    layer0_outputs(12288) <= '1';
    layer0_outputs(12289) <= (inputs(183)) xor (inputs(218));
    layer0_outputs(12290) <= not(inputs(14));
    layer0_outputs(12291) <= not(inputs(231));
    layer0_outputs(12292) <= not((inputs(148)) or (inputs(101)));
    layer0_outputs(12293) <= (inputs(60)) or (inputs(9));
    layer0_outputs(12294) <= not((inputs(66)) xor (inputs(20)));
    layer0_outputs(12295) <= not(inputs(26));
    layer0_outputs(12296) <= (inputs(184)) xor (inputs(216));
    layer0_outputs(12297) <= not(inputs(234));
    layer0_outputs(12298) <= '1';
    layer0_outputs(12299) <= '1';
    layer0_outputs(12300) <= not(inputs(122));
    layer0_outputs(12301) <= not(inputs(43)) or (inputs(186));
    layer0_outputs(12302) <= inputs(214);
    layer0_outputs(12303) <= not((inputs(74)) xor (inputs(94)));
    layer0_outputs(12304) <= (inputs(224)) or (inputs(103));
    layer0_outputs(12305) <= not(inputs(37));
    layer0_outputs(12306) <= inputs(218);
    layer0_outputs(12307) <= not((inputs(245)) or (inputs(212)));
    layer0_outputs(12308) <= inputs(135);
    layer0_outputs(12309) <= (inputs(210)) or (inputs(215));
    layer0_outputs(12310) <= not((inputs(64)) or (inputs(233)));
    layer0_outputs(12311) <= not((inputs(102)) or (inputs(77)));
    layer0_outputs(12312) <= not(inputs(241)) or (inputs(195));
    layer0_outputs(12313) <= (inputs(211)) xor (inputs(8));
    layer0_outputs(12314) <= (inputs(141)) or (inputs(232));
    layer0_outputs(12315) <= '0';
    layer0_outputs(12316) <= inputs(231);
    layer0_outputs(12317) <= not(inputs(194));
    layer0_outputs(12318) <= inputs(115);
    layer0_outputs(12319) <= '1';
    layer0_outputs(12320) <= not((inputs(168)) xor (inputs(0)));
    layer0_outputs(12321) <= (inputs(96)) and (inputs(118));
    layer0_outputs(12322) <= not((inputs(216)) xor (inputs(168)));
    layer0_outputs(12323) <= not(inputs(76));
    layer0_outputs(12324) <= (inputs(135)) and not (inputs(178));
    layer0_outputs(12325) <= (inputs(211)) or (inputs(227));
    layer0_outputs(12326) <= inputs(94);
    layer0_outputs(12327) <= not(inputs(249));
    layer0_outputs(12328) <= (inputs(148)) or (inputs(177));
    layer0_outputs(12329) <= (inputs(65)) or (inputs(247));
    layer0_outputs(12330) <= inputs(180);
    layer0_outputs(12331) <= not(inputs(108));
    layer0_outputs(12332) <= not((inputs(147)) or (inputs(85)));
    layer0_outputs(12333) <= inputs(56);
    layer0_outputs(12334) <= (inputs(155)) and (inputs(2));
    layer0_outputs(12335) <= not(inputs(128));
    layer0_outputs(12336) <= not((inputs(153)) and (inputs(140)));
    layer0_outputs(12337) <= not((inputs(202)) and (inputs(158)));
    layer0_outputs(12338) <= not(inputs(187));
    layer0_outputs(12339) <= not(inputs(78));
    layer0_outputs(12340) <= not((inputs(136)) or (inputs(66)));
    layer0_outputs(12341) <= (inputs(35)) xor (inputs(91));
    layer0_outputs(12342) <= inputs(96);
    layer0_outputs(12343) <= (inputs(143)) or (inputs(127));
    layer0_outputs(12344) <= '1';
    layer0_outputs(12345) <= not(inputs(145));
    layer0_outputs(12346) <= not((inputs(94)) xor (inputs(76)));
    layer0_outputs(12347) <= (inputs(221)) and not (inputs(143));
    layer0_outputs(12348) <= not((inputs(190)) or (inputs(74)));
    layer0_outputs(12349) <= not(inputs(211));
    layer0_outputs(12350) <= not((inputs(163)) or (inputs(188)));
    layer0_outputs(12351) <= (inputs(24)) or (inputs(252));
    layer0_outputs(12352) <= inputs(169);
    layer0_outputs(12353) <= not(inputs(69)) or (inputs(214));
    layer0_outputs(12354) <= not(inputs(215));
    layer0_outputs(12355) <= inputs(30);
    layer0_outputs(12356) <= inputs(200);
    layer0_outputs(12357) <= not((inputs(201)) or (inputs(252)));
    layer0_outputs(12358) <= not((inputs(205)) or (inputs(188)));
    layer0_outputs(12359) <= not(inputs(104));
    layer0_outputs(12360) <= '1';
    layer0_outputs(12361) <= not((inputs(125)) or (inputs(133)));
    layer0_outputs(12362) <= not((inputs(254)) or (inputs(82)));
    layer0_outputs(12363) <= (inputs(222)) and not (inputs(132));
    layer0_outputs(12364) <= not((inputs(173)) or (inputs(106)));
    layer0_outputs(12365) <= (inputs(70)) or (inputs(45));
    layer0_outputs(12366) <= not(inputs(199)) or (inputs(14));
    layer0_outputs(12367) <= (inputs(48)) or (inputs(75));
    layer0_outputs(12368) <= not((inputs(19)) xor (inputs(156)));
    layer0_outputs(12369) <= (inputs(195)) xor (inputs(222));
    layer0_outputs(12370) <= not((inputs(71)) or (inputs(28)));
    layer0_outputs(12371) <= not(inputs(233));
    layer0_outputs(12372) <= not(inputs(100)) or (inputs(59));
    layer0_outputs(12373) <= (inputs(124)) and not (inputs(62));
    layer0_outputs(12374) <= not(inputs(60));
    layer0_outputs(12375) <= not((inputs(97)) or (inputs(23)));
    layer0_outputs(12376) <= not(inputs(34)) or (inputs(17));
    layer0_outputs(12377) <= (inputs(15)) xor (inputs(205));
    layer0_outputs(12378) <= not(inputs(234)) or (inputs(82));
    layer0_outputs(12379) <= not((inputs(111)) or (inputs(138)));
    layer0_outputs(12380) <= inputs(24);
    layer0_outputs(12381) <= not(inputs(49));
    layer0_outputs(12382) <= not((inputs(106)) xor (inputs(109)));
    layer0_outputs(12383) <= inputs(174);
    layer0_outputs(12384) <= not(inputs(211));
    layer0_outputs(12385) <= not(inputs(57)) or (inputs(90));
    layer0_outputs(12386) <= not((inputs(111)) or (inputs(182)));
    layer0_outputs(12387) <= not((inputs(51)) or (inputs(177)));
    layer0_outputs(12388) <= not(inputs(19));
    layer0_outputs(12389) <= not(inputs(176)) or (inputs(212));
    layer0_outputs(12390) <= not(inputs(214));
    layer0_outputs(12391) <= (inputs(160)) and not (inputs(121));
    layer0_outputs(12392) <= (inputs(0)) and (inputs(249));
    layer0_outputs(12393) <= (inputs(179)) and not (inputs(240));
    layer0_outputs(12394) <= (inputs(54)) and not (inputs(205));
    layer0_outputs(12395) <= not((inputs(66)) xor (inputs(24)));
    layer0_outputs(12396) <= (inputs(129)) or (inputs(2));
    layer0_outputs(12397) <= inputs(118);
    layer0_outputs(12398) <= not((inputs(189)) or (inputs(247)));
    layer0_outputs(12399) <= not(inputs(116));
    layer0_outputs(12400) <= (inputs(82)) xor (inputs(163));
    layer0_outputs(12401) <= not(inputs(225));
    layer0_outputs(12402) <= not(inputs(69)) or (inputs(194));
    layer0_outputs(12403) <= (inputs(103)) and not (inputs(48));
    layer0_outputs(12404) <= not(inputs(251));
    layer0_outputs(12405) <= not((inputs(23)) and (inputs(111)));
    layer0_outputs(12406) <= inputs(70);
    layer0_outputs(12407) <= (inputs(233)) xor (inputs(112));
    layer0_outputs(12408) <= not((inputs(184)) xor (inputs(16)));
    layer0_outputs(12409) <= not(inputs(7));
    layer0_outputs(12410) <= (inputs(147)) or (inputs(168));
    layer0_outputs(12411) <= (inputs(177)) xor (inputs(155));
    layer0_outputs(12412) <= not((inputs(76)) or (inputs(95)));
    layer0_outputs(12413) <= not(inputs(72));
    layer0_outputs(12414) <= (inputs(47)) and not (inputs(192));
    layer0_outputs(12415) <= not((inputs(78)) or (inputs(35)));
    layer0_outputs(12416) <= (inputs(232)) and not (inputs(127));
    layer0_outputs(12417) <= not((inputs(255)) xor (inputs(227)));
    layer0_outputs(12418) <= not(inputs(187)) or (inputs(10));
    layer0_outputs(12419) <= inputs(39);
    layer0_outputs(12420) <= not(inputs(25)) or (inputs(155));
    layer0_outputs(12421) <= inputs(250);
    layer0_outputs(12422) <= not(inputs(133));
    layer0_outputs(12423) <= not((inputs(9)) or (inputs(77)));
    layer0_outputs(12424) <= not((inputs(110)) or (inputs(121)));
    layer0_outputs(12425) <= (inputs(163)) xor (inputs(230));
    layer0_outputs(12426) <= not((inputs(26)) xor (inputs(98)));
    layer0_outputs(12427) <= '1';
    layer0_outputs(12428) <= (inputs(69)) and not (inputs(177));
    layer0_outputs(12429) <= not((inputs(173)) and (inputs(187)));
    layer0_outputs(12430) <= not(inputs(167));
    layer0_outputs(12431) <= not(inputs(162));
    layer0_outputs(12432) <= inputs(179);
    layer0_outputs(12433) <= not((inputs(63)) xor (inputs(25)));
    layer0_outputs(12434) <= (inputs(221)) and not (inputs(142));
    layer0_outputs(12435) <= (inputs(210)) and (inputs(235));
    layer0_outputs(12436) <= inputs(25);
    layer0_outputs(12437) <= not((inputs(134)) and (inputs(129)));
    layer0_outputs(12438) <= (inputs(237)) or (inputs(235));
    layer0_outputs(12439) <= not((inputs(79)) xor (inputs(29)));
    layer0_outputs(12440) <= not(inputs(183)) or (inputs(91));
    layer0_outputs(12441) <= not(inputs(183));
    layer0_outputs(12442) <= not((inputs(54)) or (inputs(204)));
    layer0_outputs(12443) <= (inputs(4)) and not (inputs(225));
    layer0_outputs(12444) <= not((inputs(102)) xor (inputs(54)));
    layer0_outputs(12445) <= inputs(130);
    layer0_outputs(12446) <= not(inputs(163)) or (inputs(208));
    layer0_outputs(12447) <= not((inputs(15)) or (inputs(159)));
    layer0_outputs(12448) <= inputs(165);
    layer0_outputs(12449) <= (inputs(249)) or (inputs(149));
    layer0_outputs(12450) <= not((inputs(132)) xor (inputs(191)));
    layer0_outputs(12451) <= not(inputs(108)) or (inputs(154));
    layer0_outputs(12452) <= not(inputs(1)) or (inputs(38));
    layer0_outputs(12453) <= not(inputs(107)) or (inputs(220));
    layer0_outputs(12454) <= not((inputs(34)) and (inputs(205)));
    layer0_outputs(12455) <= not(inputs(144));
    layer0_outputs(12456) <= not(inputs(52));
    layer0_outputs(12457) <= not((inputs(133)) or (inputs(80)));
    layer0_outputs(12458) <= not((inputs(17)) and (inputs(171)));
    layer0_outputs(12459) <= not((inputs(88)) and (inputs(26)));
    layer0_outputs(12460) <= not((inputs(10)) or (inputs(52)));
    layer0_outputs(12461) <= not(inputs(115));
    layer0_outputs(12462) <= not(inputs(234)) or (inputs(78));
    layer0_outputs(12463) <= not((inputs(55)) xor (inputs(5)));
    layer0_outputs(12464) <= not(inputs(177));
    layer0_outputs(12465) <= inputs(110);
    layer0_outputs(12466) <= (inputs(125)) and not (inputs(194));
    layer0_outputs(12467) <= not(inputs(145));
    layer0_outputs(12468) <= (inputs(87)) xor (inputs(100));
    layer0_outputs(12469) <= not(inputs(68));
    layer0_outputs(12470) <= (inputs(179)) or (inputs(45));
    layer0_outputs(12471) <= (inputs(107)) or (inputs(54));
    layer0_outputs(12472) <= inputs(10);
    layer0_outputs(12473) <= (inputs(165)) and (inputs(177));
    layer0_outputs(12474) <= not((inputs(19)) or (inputs(62)));
    layer0_outputs(12475) <= not((inputs(209)) or (inputs(194)));
    layer0_outputs(12476) <= not((inputs(66)) xor (inputs(234)));
    layer0_outputs(12477) <= (inputs(253)) or (inputs(117));
    layer0_outputs(12478) <= not((inputs(65)) xor (inputs(6)));
    layer0_outputs(12479) <= not((inputs(105)) xor (inputs(102)));
    layer0_outputs(12480) <= '1';
    layer0_outputs(12481) <= (inputs(25)) and not (inputs(208));
    layer0_outputs(12482) <= not(inputs(216));
    layer0_outputs(12483) <= not((inputs(127)) xor (inputs(4)));
    layer0_outputs(12484) <= '1';
    layer0_outputs(12485) <= not(inputs(5)) or (inputs(175));
    layer0_outputs(12486) <= (inputs(90)) and not (inputs(128));
    layer0_outputs(12487) <= not((inputs(18)) xor (inputs(118)));
    layer0_outputs(12488) <= '1';
    layer0_outputs(12489) <= (inputs(36)) and not (inputs(229));
    layer0_outputs(12490) <= not((inputs(39)) or (inputs(111)));
    layer0_outputs(12491) <= not((inputs(228)) or (inputs(163)));
    layer0_outputs(12492) <= not(inputs(254));
    layer0_outputs(12493) <= (inputs(152)) xor (inputs(149));
    layer0_outputs(12494) <= not((inputs(235)) or (inputs(181)));
    layer0_outputs(12495) <= not(inputs(63));
    layer0_outputs(12496) <= not(inputs(164));
    layer0_outputs(12497) <= (inputs(98)) xor (inputs(149));
    layer0_outputs(12498) <= (inputs(21)) xor (inputs(194));
    layer0_outputs(12499) <= inputs(79);
    layer0_outputs(12500) <= not(inputs(76));
    layer0_outputs(12501) <= not((inputs(38)) and (inputs(81)));
    layer0_outputs(12502) <= (inputs(122)) or (inputs(35));
    layer0_outputs(12503) <= (inputs(19)) or (inputs(251));
    layer0_outputs(12504) <= (inputs(87)) and (inputs(177));
    layer0_outputs(12505) <= not(inputs(220));
    layer0_outputs(12506) <= (inputs(255)) and not (inputs(149));
    layer0_outputs(12507) <= '0';
    layer0_outputs(12508) <= not((inputs(194)) xor (inputs(225)));
    layer0_outputs(12509) <= not((inputs(67)) or (inputs(174)));
    layer0_outputs(12510) <= not(inputs(92)) or (inputs(139));
    layer0_outputs(12511) <= inputs(255);
    layer0_outputs(12512) <= not(inputs(6)) or (inputs(28));
    layer0_outputs(12513) <= (inputs(189)) or (inputs(215));
    layer0_outputs(12514) <= not((inputs(135)) or (inputs(252)));
    layer0_outputs(12515) <= not(inputs(167)) or (inputs(94));
    layer0_outputs(12516) <= (inputs(49)) and not (inputs(36));
    layer0_outputs(12517) <= (inputs(150)) and (inputs(95));
    layer0_outputs(12518) <= inputs(195);
    layer0_outputs(12519) <= not((inputs(50)) xor (inputs(141)));
    layer0_outputs(12520) <= '1';
    layer0_outputs(12521) <= (inputs(117)) xor (inputs(219));
    layer0_outputs(12522) <= inputs(211);
    layer0_outputs(12523) <= not((inputs(143)) xor (inputs(75)));
    layer0_outputs(12524) <= not(inputs(23)) or (inputs(27));
    layer0_outputs(12525) <= not(inputs(225));
    layer0_outputs(12526) <= '0';
    layer0_outputs(12527) <= not(inputs(214));
    layer0_outputs(12528) <= (inputs(3)) or (inputs(30));
    layer0_outputs(12529) <= not((inputs(196)) xor (inputs(103)));
    layer0_outputs(12530) <= inputs(21);
    layer0_outputs(12531) <= inputs(121);
    layer0_outputs(12532) <= not((inputs(246)) or (inputs(210)));
    layer0_outputs(12533) <= not((inputs(28)) or (inputs(141)));
    layer0_outputs(12534) <= '1';
    layer0_outputs(12535) <= (inputs(204)) or (inputs(235));
    layer0_outputs(12536) <= (inputs(129)) or (inputs(140));
    layer0_outputs(12537) <= '1';
    layer0_outputs(12538) <= not((inputs(236)) or (inputs(230)));
    layer0_outputs(12539) <= not((inputs(29)) xor (inputs(56)));
    layer0_outputs(12540) <= (inputs(28)) xor (inputs(176));
    layer0_outputs(12541) <= (inputs(3)) xor (inputs(213));
    layer0_outputs(12542) <= inputs(36);
    layer0_outputs(12543) <= (inputs(32)) xor (inputs(93));
    layer0_outputs(12544) <= not(inputs(88)) or (inputs(98));
    layer0_outputs(12545) <= inputs(227);
    layer0_outputs(12546) <= not(inputs(45));
    layer0_outputs(12547) <= (inputs(123)) and not (inputs(149));
    layer0_outputs(12548) <= (inputs(236)) or (inputs(219));
    layer0_outputs(12549) <= (inputs(11)) and not (inputs(51));
    layer0_outputs(12550) <= not((inputs(246)) and (inputs(247)));
    layer0_outputs(12551) <= not(inputs(104));
    layer0_outputs(12552) <= inputs(28);
    layer0_outputs(12553) <= (inputs(211)) xor (inputs(165));
    layer0_outputs(12554) <= (inputs(175)) or (inputs(128));
    layer0_outputs(12555) <= (inputs(247)) and not (inputs(3));
    layer0_outputs(12556) <= (inputs(108)) or (inputs(39));
    layer0_outputs(12557) <= (inputs(234)) and not (inputs(20));
    layer0_outputs(12558) <= not(inputs(68));
    layer0_outputs(12559) <= (inputs(206)) and not (inputs(144));
    layer0_outputs(12560) <= (inputs(49)) or (inputs(41));
    layer0_outputs(12561) <= inputs(147);
    layer0_outputs(12562) <= not(inputs(67)) or (inputs(227));
    layer0_outputs(12563) <= (inputs(106)) and not (inputs(13));
    layer0_outputs(12564) <= (inputs(110)) or (inputs(131));
    layer0_outputs(12565) <= (inputs(62)) xor (inputs(71));
    layer0_outputs(12566) <= not(inputs(68));
    layer0_outputs(12567) <= not(inputs(93));
    layer0_outputs(12568) <= not((inputs(189)) xor (inputs(185)));
    layer0_outputs(12569) <= (inputs(174)) and (inputs(129));
    layer0_outputs(12570) <= (inputs(206)) or (inputs(192));
    layer0_outputs(12571) <= (inputs(67)) and not (inputs(139));
    layer0_outputs(12572) <= (inputs(137)) and not (inputs(57));
    layer0_outputs(12573) <= not((inputs(17)) or (inputs(237)));
    layer0_outputs(12574) <= '0';
    layer0_outputs(12575) <= '1';
    layer0_outputs(12576) <= (inputs(198)) and (inputs(186));
    layer0_outputs(12577) <= not((inputs(162)) xor (inputs(235)));
    layer0_outputs(12578) <= not(inputs(44));
    layer0_outputs(12579) <= not((inputs(233)) xor (inputs(176)));
    layer0_outputs(12580) <= inputs(114);
    layer0_outputs(12581) <= (inputs(49)) or (inputs(85));
    layer0_outputs(12582) <= not(inputs(161)) or (inputs(141));
    layer0_outputs(12583) <= not(inputs(20));
    layer0_outputs(12584) <= not((inputs(112)) xor (inputs(220)));
    layer0_outputs(12585) <= not(inputs(84)) or (inputs(72));
    layer0_outputs(12586) <= not((inputs(184)) and (inputs(210)));
    layer0_outputs(12587) <= inputs(93);
    layer0_outputs(12588) <= not(inputs(219)) or (inputs(135));
    layer0_outputs(12589) <= (inputs(106)) and not (inputs(179));
    layer0_outputs(12590) <= not(inputs(103)) or (inputs(195));
    layer0_outputs(12591) <= (inputs(110)) and not (inputs(78));
    layer0_outputs(12592) <= (inputs(208)) and not (inputs(187));
    layer0_outputs(12593) <= not((inputs(32)) xor (inputs(126)));
    layer0_outputs(12594) <= not(inputs(73)) or (inputs(106));
    layer0_outputs(12595) <= inputs(88);
    layer0_outputs(12596) <= not((inputs(73)) xor (inputs(78)));
    layer0_outputs(12597) <= not(inputs(124));
    layer0_outputs(12598) <= (inputs(205)) or (inputs(246));
    layer0_outputs(12599) <= (inputs(226)) and not (inputs(91));
    layer0_outputs(12600) <= not((inputs(166)) or (inputs(110)));
    layer0_outputs(12601) <= not(inputs(179)) or (inputs(61));
    layer0_outputs(12602) <= inputs(129);
    layer0_outputs(12603) <= (inputs(165)) xor (inputs(129));
    layer0_outputs(12604) <= not((inputs(186)) or (inputs(252)));
    layer0_outputs(12605) <= not((inputs(128)) xor (inputs(78)));
    layer0_outputs(12606) <= not(inputs(121)) or (inputs(65));
    layer0_outputs(12607) <= inputs(243);
    layer0_outputs(12608) <= not(inputs(176));
    layer0_outputs(12609) <= '0';
    layer0_outputs(12610) <= (inputs(47)) xor (inputs(27));
    layer0_outputs(12611) <= inputs(32);
    layer0_outputs(12612) <= not((inputs(142)) xor (inputs(108)));
    layer0_outputs(12613) <= not((inputs(58)) or (inputs(241)));
    layer0_outputs(12614) <= not(inputs(193)) or (inputs(192));
    layer0_outputs(12615) <= not((inputs(184)) xor (inputs(28)));
    layer0_outputs(12616) <= (inputs(136)) and (inputs(139));
    layer0_outputs(12617) <= (inputs(49)) or (inputs(18));
    layer0_outputs(12618) <= (inputs(196)) or (inputs(217));
    layer0_outputs(12619) <= inputs(153);
    layer0_outputs(12620) <= not((inputs(29)) xor (inputs(107)));
    layer0_outputs(12621) <= inputs(183);
    layer0_outputs(12622) <= inputs(130);
    layer0_outputs(12623) <= inputs(141);
    layer0_outputs(12624) <= not(inputs(174));
    layer0_outputs(12625) <= not(inputs(217)) or (inputs(121));
    layer0_outputs(12626) <= (inputs(81)) or (inputs(190));
    layer0_outputs(12627) <= inputs(21);
    layer0_outputs(12628) <= not(inputs(61)) or (inputs(238));
    layer0_outputs(12629) <= inputs(40);
    layer0_outputs(12630) <= not((inputs(40)) xor (inputs(24)));
    layer0_outputs(12631) <= (inputs(196)) or (inputs(155));
    layer0_outputs(12632) <= (inputs(197)) and not (inputs(124));
    layer0_outputs(12633) <= (inputs(130)) and (inputs(188));
    layer0_outputs(12634) <= not(inputs(33)) or (inputs(241));
    layer0_outputs(12635) <= not(inputs(133));
    layer0_outputs(12636) <= not(inputs(21)) or (inputs(241));
    layer0_outputs(12637) <= not(inputs(215));
    layer0_outputs(12638) <= not((inputs(211)) or (inputs(244)));
    layer0_outputs(12639) <= (inputs(142)) and not (inputs(107));
    layer0_outputs(12640) <= not(inputs(161));
    layer0_outputs(12641) <= '1';
    layer0_outputs(12642) <= not((inputs(91)) xor (inputs(95)));
    layer0_outputs(12643) <= (inputs(99)) and not (inputs(209));
    layer0_outputs(12644) <= not(inputs(15)) or (inputs(138));
    layer0_outputs(12645) <= (inputs(42)) and (inputs(86));
    layer0_outputs(12646) <= not((inputs(0)) and (inputs(87)));
    layer0_outputs(12647) <= (inputs(73)) or (inputs(30));
    layer0_outputs(12648) <= not(inputs(146));
    layer0_outputs(12649) <= (inputs(247)) and not (inputs(177));
    layer0_outputs(12650) <= (inputs(224)) and not (inputs(74));
    layer0_outputs(12651) <= not(inputs(99));
    layer0_outputs(12652) <= not(inputs(161));
    layer0_outputs(12653) <= (inputs(119)) and not (inputs(203));
    layer0_outputs(12654) <= not(inputs(82));
    layer0_outputs(12655) <= (inputs(48)) or (inputs(217));
    layer0_outputs(12656) <= inputs(27);
    layer0_outputs(12657) <= not((inputs(161)) or (inputs(18)));
    layer0_outputs(12658) <= not(inputs(75)) or (inputs(206));
    layer0_outputs(12659) <= (inputs(47)) or (inputs(142));
    layer0_outputs(12660) <= inputs(76);
    layer0_outputs(12661) <= not(inputs(116));
    layer0_outputs(12662) <= inputs(147);
    layer0_outputs(12663) <= inputs(125);
    layer0_outputs(12664) <= inputs(128);
    layer0_outputs(12665) <= not(inputs(179));
    layer0_outputs(12666) <= inputs(244);
    layer0_outputs(12667) <= not(inputs(115));
    layer0_outputs(12668) <= not(inputs(3)) or (inputs(20));
    layer0_outputs(12669) <= (inputs(61)) or (inputs(127));
    layer0_outputs(12670) <= not(inputs(120));
    layer0_outputs(12671) <= not((inputs(52)) xor (inputs(118)));
    layer0_outputs(12672) <= not((inputs(84)) xor (inputs(122)));
    layer0_outputs(12673) <= not((inputs(140)) xor (inputs(204)));
    layer0_outputs(12674) <= (inputs(137)) and not (inputs(174));
    layer0_outputs(12675) <= not(inputs(250));
    layer0_outputs(12676) <= not((inputs(73)) or (inputs(199)));
    layer0_outputs(12677) <= not(inputs(152)) or (inputs(110));
    layer0_outputs(12678) <= not((inputs(152)) xor (inputs(250)));
    layer0_outputs(12679) <= not(inputs(89));
    layer0_outputs(12680) <= not(inputs(3)) or (inputs(76));
    layer0_outputs(12681) <= inputs(84);
    layer0_outputs(12682) <= not(inputs(85)) or (inputs(173));
    layer0_outputs(12683) <= not((inputs(191)) or (inputs(244)));
    layer0_outputs(12684) <= inputs(251);
    layer0_outputs(12685) <= (inputs(102)) or (inputs(191));
    layer0_outputs(12686) <= inputs(149);
    layer0_outputs(12687) <= not((inputs(54)) and (inputs(67)));
    layer0_outputs(12688) <= not((inputs(34)) xor (inputs(136)));
    layer0_outputs(12689) <= not(inputs(133));
    layer0_outputs(12690) <= not((inputs(68)) or (inputs(227)));
    layer0_outputs(12691) <= inputs(120);
    layer0_outputs(12692) <= not(inputs(74));
    layer0_outputs(12693) <= not((inputs(240)) and (inputs(14)));
    layer0_outputs(12694) <= '0';
    layer0_outputs(12695) <= (inputs(252)) and (inputs(145));
    layer0_outputs(12696) <= '1';
    layer0_outputs(12697) <= not((inputs(179)) or (inputs(75)));
    layer0_outputs(12698) <= not(inputs(74));
    layer0_outputs(12699) <= (inputs(194)) xor (inputs(192));
    layer0_outputs(12700) <= not((inputs(76)) xor (inputs(247)));
    layer0_outputs(12701) <= inputs(77);
    layer0_outputs(12702) <= not(inputs(56));
    layer0_outputs(12703) <= inputs(228);
    layer0_outputs(12704) <= (inputs(0)) or (inputs(138));
    layer0_outputs(12705) <= not(inputs(120)) or (inputs(69));
    layer0_outputs(12706) <= inputs(154);
    layer0_outputs(12707) <= (inputs(30)) or (inputs(134));
    layer0_outputs(12708) <= (inputs(95)) or (inputs(59));
    layer0_outputs(12709) <= not((inputs(241)) and (inputs(221)));
    layer0_outputs(12710) <= '1';
    layer0_outputs(12711) <= inputs(163);
    layer0_outputs(12712) <= not((inputs(210)) xor (inputs(206)));
    layer0_outputs(12713) <= (inputs(231)) and not (inputs(82));
    layer0_outputs(12714) <= (inputs(74)) and not (inputs(27));
    layer0_outputs(12715) <= (inputs(118)) and not (inputs(108));
    layer0_outputs(12716) <= not(inputs(6));
    layer0_outputs(12717) <= not((inputs(56)) or (inputs(105)));
    layer0_outputs(12718) <= (inputs(30)) xor (inputs(46));
    layer0_outputs(12719) <= not(inputs(232)) or (inputs(222));
    layer0_outputs(12720) <= not(inputs(248)) or (inputs(5));
    layer0_outputs(12721) <= (inputs(136)) or (inputs(4));
    layer0_outputs(12722) <= not(inputs(97)) or (inputs(107));
    layer0_outputs(12723) <= '1';
    layer0_outputs(12724) <= (inputs(251)) and not (inputs(249));
    layer0_outputs(12725) <= not(inputs(244));
    layer0_outputs(12726) <= (inputs(149)) and (inputs(188));
    layer0_outputs(12727) <= (inputs(85)) or (inputs(72));
    layer0_outputs(12728) <= not(inputs(76)) or (inputs(177));
    layer0_outputs(12729) <= not(inputs(101));
    layer0_outputs(12730) <= (inputs(31)) xor (inputs(92));
    layer0_outputs(12731) <= (inputs(196)) or (inputs(141));
    layer0_outputs(12732) <= not((inputs(199)) and (inputs(253)));
    layer0_outputs(12733) <= not((inputs(86)) xor (inputs(19)));
    layer0_outputs(12734) <= not(inputs(84)) or (inputs(18));
    layer0_outputs(12735) <= (inputs(43)) and not (inputs(225));
    layer0_outputs(12736) <= not((inputs(214)) xor (inputs(2)));
    layer0_outputs(12737) <= (inputs(154)) or (inputs(174));
    layer0_outputs(12738) <= not((inputs(91)) xor (inputs(78)));
    layer0_outputs(12739) <= not((inputs(165)) xor (inputs(189)));
    layer0_outputs(12740) <= (inputs(137)) and (inputs(0));
    layer0_outputs(12741) <= (inputs(53)) and not (inputs(150));
    layer0_outputs(12742) <= inputs(186);
    layer0_outputs(12743) <= '1';
    layer0_outputs(12744) <= not(inputs(17)) or (inputs(143));
    layer0_outputs(12745) <= (inputs(64)) and (inputs(220));
    layer0_outputs(12746) <= not(inputs(178));
    layer0_outputs(12747) <= (inputs(18)) xor (inputs(223));
    layer0_outputs(12748) <= inputs(194);
    layer0_outputs(12749) <= not((inputs(61)) or (inputs(244)));
    layer0_outputs(12750) <= inputs(113);
    layer0_outputs(12751) <= (inputs(56)) and not (inputs(206));
    layer0_outputs(12752) <= not((inputs(3)) or (inputs(248)));
    layer0_outputs(12753) <= not((inputs(236)) xor (inputs(230)));
    layer0_outputs(12754) <= inputs(130);
    layer0_outputs(12755) <= not(inputs(84));
    layer0_outputs(12756) <= (inputs(142)) xor (inputs(253));
    layer0_outputs(12757) <= inputs(73);
    layer0_outputs(12758) <= (inputs(183)) and not (inputs(81));
    layer0_outputs(12759) <= inputs(64);
    layer0_outputs(12760) <= not(inputs(167)) or (inputs(194));
    layer0_outputs(12761) <= not((inputs(176)) or (inputs(254)));
    layer0_outputs(12762) <= not(inputs(252));
    layer0_outputs(12763) <= not(inputs(182)) or (inputs(63));
    layer0_outputs(12764) <= not(inputs(9)) or (inputs(131));
    layer0_outputs(12765) <= not(inputs(207));
    layer0_outputs(12766) <= inputs(154);
    layer0_outputs(12767) <= (inputs(140)) xor (inputs(143));
    layer0_outputs(12768) <= not(inputs(123));
    layer0_outputs(12769) <= (inputs(156)) or (inputs(194));
    layer0_outputs(12770) <= inputs(227);
    layer0_outputs(12771) <= not(inputs(141));
    layer0_outputs(12772) <= not(inputs(188));
    layer0_outputs(12773) <= (inputs(38)) and not (inputs(47));
    layer0_outputs(12774) <= inputs(193);
    layer0_outputs(12775) <= inputs(59);
    layer0_outputs(12776) <= not(inputs(46));
    layer0_outputs(12777) <= (inputs(59)) and not (inputs(142));
    layer0_outputs(12778) <= (inputs(186)) and not (inputs(90));
    layer0_outputs(12779) <= inputs(68);
    layer0_outputs(12780) <= not((inputs(118)) xor (inputs(72)));
    layer0_outputs(12781) <= (inputs(89)) and not (inputs(33));
    layer0_outputs(12782) <= (inputs(216)) and not (inputs(246));
    layer0_outputs(12783) <= (inputs(145)) or (inputs(148));
    layer0_outputs(12784) <= not(inputs(139)) or (inputs(94));
    layer0_outputs(12785) <= not(inputs(8));
    layer0_outputs(12786) <= (inputs(78)) and not (inputs(239));
    layer0_outputs(12787) <= inputs(178);
    layer0_outputs(12788) <= not(inputs(244));
    layer0_outputs(12789) <= not(inputs(150));
    layer0_outputs(12790) <= not((inputs(61)) or (inputs(75)));
    layer0_outputs(12791) <= not(inputs(91));
    layer0_outputs(12792) <= not(inputs(116)) or (inputs(163));
    layer0_outputs(12793) <= inputs(1);
    layer0_outputs(12794) <= '0';
    layer0_outputs(12795) <= inputs(208);
    layer0_outputs(12796) <= not(inputs(208));
    layer0_outputs(12797) <= (inputs(60)) xor (inputs(14));
    layer0_outputs(12798) <= not(inputs(64)) or (inputs(30));
    layer0_outputs(12799) <= not((inputs(46)) or (inputs(123)));
    layer1_outputs(0) <= (layer0_outputs(2066)) or (layer0_outputs(9142));
    layer1_outputs(1) <= not(layer0_outputs(705));
    layer1_outputs(2) <= not((layer0_outputs(1387)) or (layer0_outputs(10225)));
    layer1_outputs(3) <= (layer0_outputs(5591)) xor (layer0_outputs(9562));
    layer1_outputs(4) <= not(layer0_outputs(8688));
    layer1_outputs(5) <= not(layer0_outputs(3270));
    layer1_outputs(6) <= not((layer0_outputs(2997)) and (layer0_outputs(1994)));
    layer1_outputs(7) <= layer0_outputs(8907);
    layer1_outputs(8) <= (layer0_outputs(5499)) xor (layer0_outputs(10882));
    layer1_outputs(9) <= layer0_outputs(2817);
    layer1_outputs(10) <= not(layer0_outputs(1194));
    layer1_outputs(11) <= layer0_outputs(8832);
    layer1_outputs(12) <= not((layer0_outputs(8879)) xor (layer0_outputs(3779)));
    layer1_outputs(13) <= not(layer0_outputs(2526));
    layer1_outputs(14) <= (layer0_outputs(9254)) and not (layer0_outputs(5661));
    layer1_outputs(15) <= not((layer0_outputs(7713)) and (layer0_outputs(2707)));
    layer1_outputs(16) <= (layer0_outputs(1237)) or (layer0_outputs(12022));
    layer1_outputs(17) <= not(layer0_outputs(2840)) or (layer0_outputs(1304));
    layer1_outputs(18) <= not(layer0_outputs(12066));
    layer1_outputs(19) <= layer0_outputs(12780);
    layer1_outputs(20) <= not(layer0_outputs(2087));
    layer1_outputs(21) <= layer0_outputs(8733);
    layer1_outputs(22) <= not((layer0_outputs(890)) xor (layer0_outputs(10289)));
    layer1_outputs(23) <= not((layer0_outputs(12769)) or (layer0_outputs(8946)));
    layer1_outputs(24) <= layer0_outputs(12407);
    layer1_outputs(25) <= layer0_outputs(1013);
    layer1_outputs(26) <= (layer0_outputs(11276)) and (layer0_outputs(3567));
    layer1_outputs(27) <= not(layer0_outputs(4802)) or (layer0_outputs(955));
    layer1_outputs(28) <= layer0_outputs(423);
    layer1_outputs(29) <= not(layer0_outputs(7466)) or (layer0_outputs(9592));
    layer1_outputs(30) <= not((layer0_outputs(475)) and (layer0_outputs(945)));
    layer1_outputs(31) <= not(layer0_outputs(4034));
    layer1_outputs(32) <= (layer0_outputs(11518)) and not (layer0_outputs(2425));
    layer1_outputs(33) <= layer0_outputs(6689);
    layer1_outputs(34) <= not((layer0_outputs(8750)) xor (layer0_outputs(189)));
    layer1_outputs(35) <= not(layer0_outputs(998)) or (layer0_outputs(5567));
    layer1_outputs(36) <= not((layer0_outputs(8689)) and (layer0_outputs(2292)));
    layer1_outputs(37) <= layer0_outputs(1014);
    layer1_outputs(38) <= not((layer0_outputs(6853)) xor (layer0_outputs(9665)));
    layer1_outputs(39) <= not((layer0_outputs(212)) and (layer0_outputs(5953)));
    layer1_outputs(40) <= (layer0_outputs(1191)) and (layer0_outputs(4800));
    layer1_outputs(41) <= (layer0_outputs(3065)) or (layer0_outputs(12400));
    layer1_outputs(42) <= not(layer0_outputs(11806));
    layer1_outputs(43) <= (layer0_outputs(3684)) or (layer0_outputs(1723));
    layer1_outputs(44) <= not(layer0_outputs(8183));
    layer1_outputs(45) <= (layer0_outputs(10209)) and (layer0_outputs(2592));
    layer1_outputs(46) <= not(layer0_outputs(10775));
    layer1_outputs(47) <= not(layer0_outputs(6701)) or (layer0_outputs(4550));
    layer1_outputs(48) <= not(layer0_outputs(11842));
    layer1_outputs(49) <= (layer0_outputs(2326)) and (layer0_outputs(1371));
    layer1_outputs(50) <= layer0_outputs(456);
    layer1_outputs(51) <= not(layer0_outputs(10358));
    layer1_outputs(52) <= not(layer0_outputs(4381));
    layer1_outputs(53) <= not(layer0_outputs(2252));
    layer1_outputs(54) <= (layer0_outputs(5988)) or (layer0_outputs(4610));
    layer1_outputs(55) <= not((layer0_outputs(5960)) and (layer0_outputs(10623)));
    layer1_outputs(56) <= not(layer0_outputs(1042)) or (layer0_outputs(10528));
    layer1_outputs(57) <= layer0_outputs(6841);
    layer1_outputs(58) <= not((layer0_outputs(10878)) xor (layer0_outputs(11074)));
    layer1_outputs(59) <= '0';
    layer1_outputs(60) <= not((layer0_outputs(7915)) or (layer0_outputs(10817)));
    layer1_outputs(61) <= not(layer0_outputs(7775));
    layer1_outputs(62) <= not(layer0_outputs(11324));
    layer1_outputs(63) <= layer0_outputs(1489);
    layer1_outputs(64) <= layer0_outputs(1845);
    layer1_outputs(65) <= not(layer0_outputs(2430)) or (layer0_outputs(2633));
    layer1_outputs(66) <= layer0_outputs(10127);
    layer1_outputs(67) <= (layer0_outputs(8715)) and not (layer0_outputs(6801));
    layer1_outputs(68) <= layer0_outputs(5514);
    layer1_outputs(69) <= not(layer0_outputs(7739));
    layer1_outputs(70) <= (layer0_outputs(12275)) xor (layer0_outputs(3938));
    layer1_outputs(71) <= not(layer0_outputs(5218));
    layer1_outputs(72) <= layer0_outputs(9787);
    layer1_outputs(73) <= layer0_outputs(2995);
    layer1_outputs(74) <= not(layer0_outputs(9017));
    layer1_outputs(75) <= '1';
    layer1_outputs(76) <= (layer0_outputs(4841)) or (layer0_outputs(6755));
    layer1_outputs(77) <= not((layer0_outputs(9333)) xor (layer0_outputs(2163)));
    layer1_outputs(78) <= layer0_outputs(7021);
    layer1_outputs(79) <= not(layer0_outputs(6674));
    layer1_outputs(80) <= layer0_outputs(4931);
    layer1_outputs(81) <= layer0_outputs(10540);
    layer1_outputs(82) <= not(layer0_outputs(8770));
    layer1_outputs(83) <= layer0_outputs(9503);
    layer1_outputs(84) <= not(layer0_outputs(10436)) or (layer0_outputs(8280));
    layer1_outputs(85) <= (layer0_outputs(7944)) and (layer0_outputs(5314));
    layer1_outputs(86) <= (layer0_outputs(8094)) and not (layer0_outputs(2361));
    layer1_outputs(87) <= not(layer0_outputs(11629)) or (layer0_outputs(4983));
    layer1_outputs(88) <= not(layer0_outputs(7799));
    layer1_outputs(89) <= not(layer0_outputs(4778)) or (layer0_outputs(10708));
    layer1_outputs(90) <= (layer0_outputs(6645)) and not (layer0_outputs(11251));
    layer1_outputs(91) <= (layer0_outputs(4653)) and not (layer0_outputs(6602));
    layer1_outputs(92) <= (layer0_outputs(12388)) and not (layer0_outputs(7776));
    layer1_outputs(93) <= not((layer0_outputs(2784)) and (layer0_outputs(8239)));
    layer1_outputs(94) <= not((layer0_outputs(10645)) and (layer0_outputs(2180)));
    layer1_outputs(95) <= '1';
    layer1_outputs(96) <= (layer0_outputs(7947)) xor (layer0_outputs(3206));
    layer1_outputs(97) <= (layer0_outputs(3662)) and (layer0_outputs(10494));
    layer1_outputs(98) <= not(layer0_outputs(6927));
    layer1_outputs(99) <= not(layer0_outputs(12624)) or (layer0_outputs(12657));
    layer1_outputs(100) <= (layer0_outputs(6217)) and not (layer0_outputs(5122));
    layer1_outputs(101) <= layer0_outputs(5948);
    layer1_outputs(102) <= not(layer0_outputs(2157));
    layer1_outputs(103) <= not(layer0_outputs(4142));
    layer1_outputs(104) <= (layer0_outputs(7220)) and (layer0_outputs(3244));
    layer1_outputs(105) <= not(layer0_outputs(8780)) or (layer0_outputs(4581));
    layer1_outputs(106) <= (layer0_outputs(11746)) and (layer0_outputs(12422));
    layer1_outputs(107) <= not((layer0_outputs(5231)) and (layer0_outputs(4068)));
    layer1_outputs(108) <= (layer0_outputs(9329)) and not (layer0_outputs(8484));
    layer1_outputs(109) <= (layer0_outputs(7952)) and not (layer0_outputs(9678));
    layer1_outputs(110) <= layer0_outputs(8199);
    layer1_outputs(111) <= not(layer0_outputs(12019));
    layer1_outputs(112) <= layer0_outputs(675);
    layer1_outputs(113) <= (layer0_outputs(8926)) and (layer0_outputs(12146));
    layer1_outputs(114) <= (layer0_outputs(10112)) xor (layer0_outputs(7155));
    layer1_outputs(115) <= (layer0_outputs(6344)) and not (layer0_outputs(7240));
    layer1_outputs(116) <= not((layer0_outputs(1083)) or (layer0_outputs(5652)));
    layer1_outputs(117) <= not(layer0_outputs(4734)) or (layer0_outputs(12227));
    layer1_outputs(118) <= not(layer0_outputs(9647));
    layer1_outputs(119) <= not(layer0_outputs(7997));
    layer1_outputs(120) <= not(layer0_outputs(1719)) or (layer0_outputs(2083));
    layer1_outputs(121) <= not((layer0_outputs(10020)) and (layer0_outputs(32)));
    layer1_outputs(122) <= not((layer0_outputs(9058)) or (layer0_outputs(4099)));
    layer1_outputs(123) <= not((layer0_outputs(9187)) and (layer0_outputs(8732)));
    layer1_outputs(124) <= (layer0_outputs(1166)) and (layer0_outputs(4036));
    layer1_outputs(125) <= not(layer0_outputs(3944)) or (layer0_outputs(7026));
    layer1_outputs(126) <= not(layer0_outputs(6788)) or (layer0_outputs(5777));
    layer1_outputs(127) <= layer0_outputs(4253);
    layer1_outputs(128) <= not(layer0_outputs(5497));
    layer1_outputs(129) <= not((layer0_outputs(6690)) or (layer0_outputs(1125)));
    layer1_outputs(130) <= (layer0_outputs(1706)) xor (layer0_outputs(9827));
    layer1_outputs(131) <= not((layer0_outputs(5241)) xor (layer0_outputs(5659)));
    layer1_outputs(132) <= layer0_outputs(1769);
    layer1_outputs(133) <= '1';
    layer1_outputs(134) <= not((layer0_outputs(9457)) and (layer0_outputs(10544)));
    layer1_outputs(135) <= (layer0_outputs(1578)) and not (layer0_outputs(363));
    layer1_outputs(136) <= not(layer0_outputs(5662));
    layer1_outputs(137) <= not(layer0_outputs(9668)) or (layer0_outputs(4490));
    layer1_outputs(138) <= not(layer0_outputs(4217)) or (layer0_outputs(9046));
    layer1_outputs(139) <= layer0_outputs(10472);
    layer1_outputs(140) <= not(layer0_outputs(1881)) or (layer0_outputs(3124));
    layer1_outputs(141) <= not((layer0_outputs(7577)) xor (layer0_outputs(6927)));
    layer1_outputs(142) <= not(layer0_outputs(2867));
    layer1_outputs(143) <= (layer0_outputs(63)) and not (layer0_outputs(1828));
    layer1_outputs(144) <= not((layer0_outputs(1230)) and (layer0_outputs(9646)));
    layer1_outputs(145) <= layer0_outputs(2216);
    layer1_outputs(146) <= not(layer0_outputs(1433)) or (layer0_outputs(1428));
    layer1_outputs(147) <= not(layer0_outputs(142));
    layer1_outputs(148) <= '0';
    layer1_outputs(149) <= not((layer0_outputs(7066)) xor (layer0_outputs(1458)));
    layer1_outputs(150) <= (layer0_outputs(12200)) and not (layer0_outputs(7999));
    layer1_outputs(151) <= layer0_outputs(4078);
    layer1_outputs(152) <= (layer0_outputs(3620)) and not (layer0_outputs(7933));
    layer1_outputs(153) <= not((layer0_outputs(2142)) and (layer0_outputs(1594)));
    layer1_outputs(154) <= '0';
    layer1_outputs(155) <= layer0_outputs(9949);
    layer1_outputs(156) <= (layer0_outputs(6658)) or (layer0_outputs(4776));
    layer1_outputs(157) <= not((layer0_outputs(9802)) or (layer0_outputs(3045)));
    layer1_outputs(158) <= (layer0_outputs(6095)) and not (layer0_outputs(2450));
    layer1_outputs(159) <= not((layer0_outputs(727)) and (layer0_outputs(9499)));
    layer1_outputs(160) <= (layer0_outputs(11583)) xor (layer0_outputs(11423));
    layer1_outputs(161) <= (layer0_outputs(12155)) and (layer0_outputs(2583));
    layer1_outputs(162) <= not(layer0_outputs(12350)) or (layer0_outputs(1233));
    layer1_outputs(163) <= not(layer0_outputs(1375));
    layer1_outputs(164) <= not((layer0_outputs(7764)) or (layer0_outputs(8777)));
    layer1_outputs(165) <= (layer0_outputs(10011)) or (layer0_outputs(4675));
    layer1_outputs(166) <= (layer0_outputs(12082)) and not (layer0_outputs(556));
    layer1_outputs(167) <= not(layer0_outputs(4097));
    layer1_outputs(168) <= not(layer0_outputs(7367));
    layer1_outputs(169) <= layer0_outputs(5948);
    layer1_outputs(170) <= not(layer0_outputs(5224));
    layer1_outputs(171) <= not(layer0_outputs(1794));
    layer1_outputs(172) <= not(layer0_outputs(6860));
    layer1_outputs(173) <= (layer0_outputs(5758)) and (layer0_outputs(2171));
    layer1_outputs(174) <= (layer0_outputs(857)) and (layer0_outputs(6814));
    layer1_outputs(175) <= not(layer0_outputs(6515));
    layer1_outputs(176) <= (layer0_outputs(19)) xor (layer0_outputs(1162));
    layer1_outputs(177) <= layer0_outputs(5621);
    layer1_outputs(178) <= layer0_outputs(795);
    layer1_outputs(179) <= not(layer0_outputs(11137)) or (layer0_outputs(8809));
    layer1_outputs(180) <= (layer0_outputs(3016)) and not (layer0_outputs(12180));
    layer1_outputs(181) <= not((layer0_outputs(12472)) and (layer0_outputs(585)));
    layer1_outputs(182) <= not(layer0_outputs(10652));
    layer1_outputs(183) <= not(layer0_outputs(3350)) or (layer0_outputs(6695));
    layer1_outputs(184) <= not(layer0_outputs(949)) or (layer0_outputs(11490));
    layer1_outputs(185) <= not(layer0_outputs(1914));
    layer1_outputs(186) <= '1';
    layer1_outputs(187) <= not(layer0_outputs(12521));
    layer1_outputs(188) <= not(layer0_outputs(5212));
    layer1_outputs(189) <= not(layer0_outputs(8569));
    layer1_outputs(190) <= (layer0_outputs(12203)) or (layer0_outputs(2277));
    layer1_outputs(191) <= layer0_outputs(4136);
    layer1_outputs(192) <= layer0_outputs(5582);
    layer1_outputs(193) <= (layer0_outputs(389)) and (layer0_outputs(5807));
    layer1_outputs(194) <= (layer0_outputs(8132)) or (layer0_outputs(6600));
    layer1_outputs(195) <= (layer0_outputs(2561)) and not (layer0_outputs(4950));
    layer1_outputs(196) <= not((layer0_outputs(9697)) or (layer0_outputs(4271)));
    layer1_outputs(197) <= not(layer0_outputs(3386)) or (layer0_outputs(6581));
    layer1_outputs(198) <= (layer0_outputs(10606)) xor (layer0_outputs(240));
    layer1_outputs(199) <= not((layer0_outputs(144)) xor (layer0_outputs(4869)));
    layer1_outputs(200) <= not(layer0_outputs(1246));
    layer1_outputs(201) <= not(layer0_outputs(12113));
    layer1_outputs(202) <= not(layer0_outputs(9521));
    layer1_outputs(203) <= not(layer0_outputs(12352));
    layer1_outputs(204) <= not((layer0_outputs(10318)) and (layer0_outputs(9007)));
    layer1_outputs(205) <= not(layer0_outputs(8817)) or (layer0_outputs(7965));
    layer1_outputs(206) <= (layer0_outputs(5153)) and not (layer0_outputs(9432));
    layer1_outputs(207) <= layer0_outputs(12328);
    layer1_outputs(208) <= not((layer0_outputs(11745)) xor (layer0_outputs(1715)));
    layer1_outputs(209) <= (layer0_outputs(11131)) and not (layer0_outputs(7898));
    layer1_outputs(210) <= not((layer0_outputs(12506)) xor (layer0_outputs(8214)));
    layer1_outputs(211) <= layer0_outputs(7057);
    layer1_outputs(212) <= (layer0_outputs(2107)) xor (layer0_outputs(11208));
    layer1_outputs(213) <= not((layer0_outputs(6294)) and (layer0_outputs(4999)));
    layer1_outputs(214) <= (layer0_outputs(3444)) and (layer0_outputs(12653));
    layer1_outputs(215) <= not(layer0_outputs(9690));
    layer1_outputs(216) <= not((layer0_outputs(2614)) or (layer0_outputs(5573)));
    layer1_outputs(217) <= (layer0_outputs(1657)) xor (layer0_outputs(4166));
    layer1_outputs(218) <= not((layer0_outputs(8325)) xor (layer0_outputs(972)));
    layer1_outputs(219) <= not(layer0_outputs(12393));
    layer1_outputs(220) <= layer0_outputs(6117);
    layer1_outputs(221) <= (layer0_outputs(8905)) and (layer0_outputs(9876));
    layer1_outputs(222) <= (layer0_outputs(2842)) or (layer0_outputs(7084));
    layer1_outputs(223) <= (layer0_outputs(11099)) or (layer0_outputs(6660));
    layer1_outputs(224) <= layer0_outputs(949);
    layer1_outputs(225) <= not(layer0_outputs(11783));
    layer1_outputs(226) <= (layer0_outputs(2858)) and (layer0_outputs(8535));
    layer1_outputs(227) <= layer0_outputs(3212);
    layer1_outputs(228) <= (layer0_outputs(9614)) and not (layer0_outputs(2540));
    layer1_outputs(229) <= not((layer0_outputs(6032)) and (layer0_outputs(8250)));
    layer1_outputs(230) <= layer0_outputs(151);
    layer1_outputs(231) <= layer0_outputs(3905);
    layer1_outputs(232) <= not((layer0_outputs(4125)) and (layer0_outputs(12236)));
    layer1_outputs(233) <= layer0_outputs(437);
    layer1_outputs(234) <= (layer0_outputs(9969)) and (layer0_outputs(3841));
    layer1_outputs(235) <= layer0_outputs(12255);
    layer1_outputs(236) <= (layer0_outputs(6563)) and not (layer0_outputs(1463));
    layer1_outputs(237) <= not(layer0_outputs(2968));
    layer1_outputs(238) <= layer0_outputs(6975);
    layer1_outputs(239) <= layer0_outputs(6205);
    layer1_outputs(240) <= (layer0_outputs(3589)) or (layer0_outputs(8845));
    layer1_outputs(241) <= (layer0_outputs(1720)) xor (layer0_outputs(11090));
    layer1_outputs(242) <= (layer0_outputs(8873)) xor (layer0_outputs(1328));
    layer1_outputs(243) <= (layer0_outputs(1677)) xor (layer0_outputs(7462));
    layer1_outputs(244) <= (layer0_outputs(7007)) and (layer0_outputs(5034));
    layer1_outputs(245) <= (layer0_outputs(3529)) and not (layer0_outputs(6034));
    layer1_outputs(246) <= not((layer0_outputs(6858)) xor (layer0_outputs(6681)));
    layer1_outputs(247) <= not(layer0_outputs(10846)) or (layer0_outputs(1054));
    layer1_outputs(248) <= not((layer0_outputs(5050)) xor (layer0_outputs(11680)));
    layer1_outputs(249) <= not(layer0_outputs(11097));
    layer1_outputs(250) <= not(layer0_outputs(8803));
    layer1_outputs(251) <= not(layer0_outputs(7642));
    layer1_outputs(252) <= layer0_outputs(8100);
    layer1_outputs(253) <= not((layer0_outputs(11749)) or (layer0_outputs(12536)));
    layer1_outputs(254) <= not(layer0_outputs(641)) or (layer0_outputs(786));
    layer1_outputs(255) <= not(layer0_outputs(9222));
    layer1_outputs(256) <= not((layer0_outputs(3944)) or (layer0_outputs(81)));
    layer1_outputs(257) <= layer0_outputs(10876);
    layer1_outputs(258) <= not(layer0_outputs(10228)) or (layer0_outputs(2169));
    layer1_outputs(259) <= not(layer0_outputs(4502));
    layer1_outputs(260) <= (layer0_outputs(242)) and (layer0_outputs(7126));
    layer1_outputs(261) <= not((layer0_outputs(1446)) or (layer0_outputs(904)));
    layer1_outputs(262) <= not(layer0_outputs(9450));
    layer1_outputs(263) <= (layer0_outputs(1044)) and not (layer0_outputs(4662));
    layer1_outputs(264) <= not(layer0_outputs(7389));
    layer1_outputs(265) <= not(layer0_outputs(12557));
    layer1_outputs(266) <= layer0_outputs(5792);
    layer1_outputs(267) <= layer0_outputs(6538);
    layer1_outputs(268) <= (layer0_outputs(4442)) and not (layer0_outputs(8865));
    layer1_outputs(269) <= not((layer0_outputs(6232)) xor (layer0_outputs(5482)));
    layer1_outputs(270) <= layer0_outputs(264);
    layer1_outputs(271) <= (layer0_outputs(11)) xor (layer0_outputs(6511));
    layer1_outputs(272) <= not(layer0_outputs(9050));
    layer1_outputs(273) <= not((layer0_outputs(11901)) or (layer0_outputs(3333)));
    layer1_outputs(274) <= layer0_outputs(9441);
    layer1_outputs(275) <= not((layer0_outputs(10416)) or (layer0_outputs(7281)));
    layer1_outputs(276) <= not((layer0_outputs(1935)) and (layer0_outputs(9282)));
    layer1_outputs(277) <= not(layer0_outputs(7215));
    layer1_outputs(278) <= not(layer0_outputs(2740));
    layer1_outputs(279) <= not(layer0_outputs(1493));
    layer1_outputs(280) <= (layer0_outputs(9793)) xor (layer0_outputs(7994));
    layer1_outputs(281) <= (layer0_outputs(3091)) xor (layer0_outputs(10569));
    layer1_outputs(282) <= not(layer0_outputs(1298));
    layer1_outputs(283) <= not(layer0_outputs(9757));
    layer1_outputs(284) <= not(layer0_outputs(8849)) or (layer0_outputs(11879));
    layer1_outputs(285) <= layer0_outputs(12223);
    layer1_outputs(286) <= (layer0_outputs(8603)) and not (layer0_outputs(7472));
    layer1_outputs(287) <= not(layer0_outputs(10158));
    layer1_outputs(288) <= not(layer0_outputs(4996));
    layer1_outputs(289) <= not(layer0_outputs(10650));
    layer1_outputs(290) <= layer0_outputs(6913);
    layer1_outputs(291) <= not(layer0_outputs(7178));
    layer1_outputs(292) <= not((layer0_outputs(6846)) or (layer0_outputs(12759)));
    layer1_outputs(293) <= (layer0_outputs(2124)) or (layer0_outputs(1405));
    layer1_outputs(294) <= layer0_outputs(10394);
    layer1_outputs(295) <= (layer0_outputs(11555)) and not (layer0_outputs(4822));
    layer1_outputs(296) <= not((layer0_outputs(10727)) and (layer0_outputs(473)));
    layer1_outputs(297) <= not(layer0_outputs(2902));
    layer1_outputs(298) <= (layer0_outputs(8700)) or (layer0_outputs(12791));
    layer1_outputs(299) <= layer0_outputs(12411);
    layer1_outputs(300) <= not(layer0_outputs(4350)) or (layer0_outputs(2040));
    layer1_outputs(301) <= layer0_outputs(6561);
    layer1_outputs(302) <= layer0_outputs(3566);
    layer1_outputs(303) <= not(layer0_outputs(12387)) or (layer0_outputs(7237));
    layer1_outputs(304) <= layer0_outputs(398);
    layer1_outputs(305) <= not(layer0_outputs(6756));
    layer1_outputs(306) <= layer0_outputs(2807);
    layer1_outputs(307) <= (layer0_outputs(7804)) and (layer0_outputs(2138));
    layer1_outputs(308) <= not(layer0_outputs(55)) or (layer0_outputs(9987));
    layer1_outputs(309) <= (layer0_outputs(1636)) or (layer0_outputs(5931));
    layer1_outputs(310) <= '0';
    layer1_outputs(311) <= not(layer0_outputs(12364));
    layer1_outputs(312) <= not((layer0_outputs(1087)) and (layer0_outputs(5429)));
    layer1_outputs(313) <= not((layer0_outputs(4774)) or (layer0_outputs(1144)));
    layer1_outputs(314) <= not((layer0_outputs(11510)) xor (layer0_outputs(1715)));
    layer1_outputs(315) <= not(layer0_outputs(4745)) or (layer0_outputs(7320));
    layer1_outputs(316) <= not(layer0_outputs(11404));
    layer1_outputs(317) <= not((layer0_outputs(6666)) or (layer0_outputs(11875)));
    layer1_outputs(318) <= not(layer0_outputs(10784));
    layer1_outputs(319) <= '1';
    layer1_outputs(320) <= not(layer0_outputs(1045));
    layer1_outputs(321) <= not(layer0_outputs(4605)) or (layer0_outputs(11366));
    layer1_outputs(322) <= layer0_outputs(921);
    layer1_outputs(323) <= (layer0_outputs(10583)) or (layer0_outputs(12692));
    layer1_outputs(324) <= not(layer0_outputs(12645));
    layer1_outputs(325) <= (layer0_outputs(10512)) or (layer0_outputs(5163));
    layer1_outputs(326) <= not((layer0_outputs(1953)) xor (layer0_outputs(3143)));
    layer1_outputs(327) <= not(layer0_outputs(4650));
    layer1_outputs(328) <= not((layer0_outputs(2794)) or (layer0_outputs(7908)));
    layer1_outputs(329) <= not(layer0_outputs(6902));
    layer1_outputs(330) <= not(layer0_outputs(5551)) or (layer0_outputs(8274));
    layer1_outputs(331) <= (layer0_outputs(3581)) and (layer0_outputs(1043));
    layer1_outputs(332) <= not((layer0_outputs(8459)) xor (layer0_outputs(8166)));
    layer1_outputs(333) <= layer0_outputs(8016);
    layer1_outputs(334) <= not(layer0_outputs(5254));
    layer1_outputs(335) <= not((layer0_outputs(12036)) or (layer0_outputs(134)));
    layer1_outputs(336) <= layer0_outputs(1631);
    layer1_outputs(337) <= layer0_outputs(1048);
    layer1_outputs(338) <= layer0_outputs(7335);
    layer1_outputs(339) <= (layer0_outputs(9416)) or (layer0_outputs(4641));
    layer1_outputs(340) <= not(layer0_outputs(5679)) or (layer0_outputs(5503));
    layer1_outputs(341) <= (layer0_outputs(11730)) and (layer0_outputs(8668));
    layer1_outputs(342) <= not((layer0_outputs(11257)) xor (layer0_outputs(4446)));
    layer1_outputs(343) <= (layer0_outputs(3798)) and not (layer0_outputs(10909));
    layer1_outputs(344) <= layer0_outputs(581);
    layer1_outputs(345) <= not((layer0_outputs(10128)) xor (layer0_outputs(8861)));
    layer1_outputs(346) <= not(layer0_outputs(3033));
    layer1_outputs(347) <= not((layer0_outputs(7357)) and (layer0_outputs(2786)));
    layer1_outputs(348) <= layer0_outputs(11839);
    layer1_outputs(349) <= '1';
    layer1_outputs(350) <= not(layer0_outputs(8577));
    layer1_outputs(351) <= (layer0_outputs(11867)) and not (layer0_outputs(1594));
    layer1_outputs(352) <= not(layer0_outputs(8238));
    layer1_outputs(353) <= not(layer0_outputs(2163)) or (layer0_outputs(8871));
    layer1_outputs(354) <= (layer0_outputs(11289)) xor (layer0_outputs(5570));
    layer1_outputs(355) <= (layer0_outputs(10685)) and (layer0_outputs(724));
    layer1_outputs(356) <= not(layer0_outputs(660));
    layer1_outputs(357) <= (layer0_outputs(8800)) or (layer0_outputs(5112));
    layer1_outputs(358) <= not(layer0_outputs(10459)) or (layer0_outputs(405));
    layer1_outputs(359) <= not(layer0_outputs(11389));
    layer1_outputs(360) <= (layer0_outputs(4593)) or (layer0_outputs(642));
    layer1_outputs(361) <= not(layer0_outputs(3375));
    layer1_outputs(362) <= not((layer0_outputs(12568)) and (layer0_outputs(8151)));
    layer1_outputs(363) <= not((layer0_outputs(9330)) or (layer0_outputs(9407)));
    layer1_outputs(364) <= not(layer0_outputs(6419)) or (layer0_outputs(8527));
    layer1_outputs(365) <= not(layer0_outputs(640)) or (layer0_outputs(1972));
    layer1_outputs(366) <= not(layer0_outputs(6650));
    layer1_outputs(367) <= not((layer0_outputs(2469)) xor (layer0_outputs(10243)));
    layer1_outputs(368) <= layer0_outputs(10129);
    layer1_outputs(369) <= layer0_outputs(6401);
    layer1_outputs(370) <= not((layer0_outputs(7401)) and (layer0_outputs(11902)));
    layer1_outputs(371) <= (layer0_outputs(1826)) and (layer0_outputs(2769));
    layer1_outputs(372) <= not(layer0_outputs(4649)) or (layer0_outputs(6417));
    layer1_outputs(373) <= (layer0_outputs(8207)) and not (layer0_outputs(9836));
    layer1_outputs(374) <= not((layer0_outputs(1630)) xor (layer0_outputs(6482)));
    layer1_outputs(375) <= (layer0_outputs(2849)) and (layer0_outputs(10568));
    layer1_outputs(376) <= '1';
    layer1_outputs(377) <= not((layer0_outputs(8827)) xor (layer0_outputs(5398)));
    layer1_outputs(378) <= not(layer0_outputs(10101)) or (layer0_outputs(6297));
    layer1_outputs(379) <= not(layer0_outputs(9931));
    layer1_outputs(380) <= not((layer0_outputs(12432)) or (layer0_outputs(3622)));
    layer1_outputs(381) <= not(layer0_outputs(6252)) or (layer0_outputs(11712));
    layer1_outputs(382) <= layer0_outputs(6146);
    layer1_outputs(383) <= '1';
    layer1_outputs(384) <= not(layer0_outputs(7334)) or (layer0_outputs(8290));
    layer1_outputs(385) <= layer0_outputs(5783);
    layer1_outputs(386) <= not(layer0_outputs(7506));
    layer1_outputs(387) <= not(layer0_outputs(5461));
    layer1_outputs(388) <= (layer0_outputs(9350)) and not (layer0_outputs(1951));
    layer1_outputs(389) <= layer0_outputs(9468);
    layer1_outputs(390) <= not(layer0_outputs(12737)) or (layer0_outputs(7391));
    layer1_outputs(391) <= layer0_outputs(3776);
    layer1_outputs(392) <= not(layer0_outputs(3439));
    layer1_outputs(393) <= not(layer0_outputs(175)) or (layer0_outputs(1346));
    layer1_outputs(394) <= (layer0_outputs(7227)) and not (layer0_outputs(2358));
    layer1_outputs(395) <= (layer0_outputs(3035)) or (layer0_outputs(1948));
    layer1_outputs(396) <= not((layer0_outputs(11049)) xor (layer0_outputs(1075)));
    layer1_outputs(397) <= (layer0_outputs(6907)) or (layer0_outputs(6974));
    layer1_outputs(398) <= not(layer0_outputs(12370));
    layer1_outputs(399) <= layer0_outputs(294);
    layer1_outputs(400) <= '0';
    layer1_outputs(401) <= not(layer0_outputs(11084));
    layer1_outputs(402) <= layer0_outputs(4353);
    layer1_outputs(403) <= (layer0_outputs(3732)) or (layer0_outputs(1124));
    layer1_outputs(404) <= not(layer0_outputs(8968));
    layer1_outputs(405) <= not((layer0_outputs(5006)) xor (layer0_outputs(58)));
    layer1_outputs(406) <= layer0_outputs(10201);
    layer1_outputs(407) <= not(layer0_outputs(1802)) or (layer0_outputs(2316));
    layer1_outputs(408) <= (layer0_outputs(11879)) and not (layer0_outputs(10384));
    layer1_outputs(409) <= not(layer0_outputs(10422));
    layer1_outputs(410) <= not(layer0_outputs(5716));
    layer1_outputs(411) <= not(layer0_outputs(825));
    layer1_outputs(412) <= layer0_outputs(5183);
    layer1_outputs(413) <= layer0_outputs(11030);
    layer1_outputs(414) <= not(layer0_outputs(6686)) or (layer0_outputs(10253));
    layer1_outputs(415) <= not((layer0_outputs(1438)) and (layer0_outputs(9762)));
    layer1_outputs(416) <= not(layer0_outputs(1058));
    layer1_outputs(417) <= not(layer0_outputs(2949));
    layer1_outputs(418) <= not((layer0_outputs(2299)) xor (layer0_outputs(5475)));
    layer1_outputs(419) <= layer0_outputs(10410);
    layer1_outputs(420) <= not(layer0_outputs(10347));
    layer1_outputs(421) <= layer0_outputs(3960);
    layer1_outputs(422) <= layer0_outputs(8252);
    layer1_outputs(423) <= not(layer0_outputs(7476)) or (layer0_outputs(11668));
    layer1_outputs(424) <= layer0_outputs(2531);
    layer1_outputs(425) <= not(layer0_outputs(10743)) or (layer0_outputs(11146));
    layer1_outputs(426) <= layer0_outputs(2349);
    layer1_outputs(427) <= layer0_outputs(11544);
    layer1_outputs(428) <= not(layer0_outputs(11720));
    layer1_outputs(429) <= not(layer0_outputs(11176));
    layer1_outputs(430) <= not((layer0_outputs(2879)) xor (layer0_outputs(874)));
    layer1_outputs(431) <= not((layer0_outputs(9444)) xor (layer0_outputs(2862)));
    layer1_outputs(432) <= layer0_outputs(3719);
    layer1_outputs(433) <= not(layer0_outputs(12706));
    layer1_outputs(434) <= (layer0_outputs(6938)) xor (layer0_outputs(7064));
    layer1_outputs(435) <= (layer0_outputs(1397)) and (layer0_outputs(10603));
    layer1_outputs(436) <= (layer0_outputs(10970)) and not (layer0_outputs(5341));
    layer1_outputs(437) <= layer0_outputs(12372);
    layer1_outputs(438) <= layer0_outputs(331);
    layer1_outputs(439) <= layer0_outputs(8085);
    layer1_outputs(440) <= layer0_outputs(8192);
    layer1_outputs(441) <= layer0_outputs(1196);
    layer1_outputs(442) <= not(layer0_outputs(12621));
    layer1_outputs(443) <= not((layer0_outputs(8283)) xor (layer0_outputs(9911)));
    layer1_outputs(444) <= not((layer0_outputs(526)) xor (layer0_outputs(11427)));
    layer1_outputs(445) <= layer0_outputs(10490);
    layer1_outputs(446) <= layer0_outputs(12587);
    layer1_outputs(447) <= not(layer0_outputs(2103)) or (layer0_outputs(10946));
    layer1_outputs(448) <= not((layer0_outputs(4522)) or (layer0_outputs(1062)));
    layer1_outputs(449) <= (layer0_outputs(11001)) or (layer0_outputs(9088));
    layer1_outputs(450) <= not((layer0_outputs(4905)) and (layer0_outputs(12015)));
    layer1_outputs(451) <= layer0_outputs(12560);
    layer1_outputs(452) <= not(layer0_outputs(11002));
    layer1_outputs(453) <= (layer0_outputs(1973)) xor (layer0_outputs(8308));
    layer1_outputs(454) <= not(layer0_outputs(5541)) or (layer0_outputs(214));
    layer1_outputs(455) <= layer0_outputs(12566);
    layer1_outputs(456) <= not(layer0_outputs(10277));
    layer1_outputs(457) <= not((layer0_outputs(11497)) or (layer0_outputs(9593)));
    layer1_outputs(458) <= layer0_outputs(3356);
    layer1_outputs(459) <= (layer0_outputs(4424)) and (layer0_outputs(11120));
    layer1_outputs(460) <= (layer0_outputs(6243)) and (layer0_outputs(1343));
    layer1_outputs(461) <= (layer0_outputs(11969)) and not (layer0_outputs(10147));
    layer1_outputs(462) <= not(layer0_outputs(7259)) or (layer0_outputs(9973));
    layer1_outputs(463) <= (layer0_outputs(8412)) xor (layer0_outputs(11193));
    layer1_outputs(464) <= not(layer0_outputs(8626));
    layer1_outputs(465) <= (layer0_outputs(5578)) and not (layer0_outputs(8146));
    layer1_outputs(466) <= layer0_outputs(3480);
    layer1_outputs(467) <= not(layer0_outputs(1479));
    layer1_outputs(468) <= layer0_outputs(85);
    layer1_outputs(469) <= not(layer0_outputs(8614)) or (layer0_outputs(9621));
    layer1_outputs(470) <= not(layer0_outputs(4671));
    layer1_outputs(471) <= not(layer0_outputs(429));
    layer1_outputs(472) <= (layer0_outputs(1038)) or (layer0_outputs(7271));
    layer1_outputs(473) <= (layer0_outputs(9705)) and not (layer0_outputs(4854));
    layer1_outputs(474) <= not(layer0_outputs(11058));
    layer1_outputs(475) <= (layer0_outputs(6314)) and not (layer0_outputs(9656));
    layer1_outputs(476) <= (layer0_outputs(11385)) and (layer0_outputs(8999));
    layer1_outputs(477) <= not(layer0_outputs(10108));
    layer1_outputs(478) <= (layer0_outputs(6769)) or (layer0_outputs(795));
    layer1_outputs(479) <= (layer0_outputs(5159)) xor (layer0_outputs(1220));
    layer1_outputs(480) <= (layer0_outputs(11882)) and not (layer0_outputs(3178));
    layer1_outputs(481) <= layer0_outputs(5914);
    layer1_outputs(482) <= not(layer0_outputs(9926));
    layer1_outputs(483) <= not(layer0_outputs(5675));
    layer1_outputs(484) <= not(layer0_outputs(7175));
    layer1_outputs(485) <= (layer0_outputs(8386)) xor (layer0_outputs(12607));
    layer1_outputs(486) <= not((layer0_outputs(6125)) xor (layer0_outputs(7085)));
    layer1_outputs(487) <= (layer0_outputs(2388)) or (layer0_outputs(281));
    layer1_outputs(488) <= not(layer0_outputs(2288));
    layer1_outputs(489) <= not(layer0_outputs(7225));
    layer1_outputs(490) <= (layer0_outputs(533)) and not (layer0_outputs(4622));
    layer1_outputs(491) <= not((layer0_outputs(3977)) xor (layer0_outputs(3451)));
    layer1_outputs(492) <= (layer0_outputs(10907)) and (layer0_outputs(6496));
    layer1_outputs(493) <= not(layer0_outputs(10925));
    layer1_outputs(494) <= not(layer0_outputs(217));
    layer1_outputs(495) <= (layer0_outputs(11361)) and not (layer0_outputs(3217));
    layer1_outputs(496) <= not(layer0_outputs(12153));
    layer1_outputs(497) <= not(layer0_outputs(11106));
    layer1_outputs(498) <= not(layer0_outputs(2364));
    layer1_outputs(499) <= not(layer0_outputs(1296));
    layer1_outputs(500) <= '1';
    layer1_outputs(501) <= not(layer0_outputs(2930));
    layer1_outputs(502) <= not(layer0_outputs(7308)) or (layer0_outputs(615));
    layer1_outputs(503) <= layer0_outputs(3725);
    layer1_outputs(504) <= not(layer0_outputs(4444));
    layer1_outputs(505) <= (layer0_outputs(7498)) and not (layer0_outputs(4120));
    layer1_outputs(506) <= layer0_outputs(2174);
    layer1_outputs(507) <= layer0_outputs(10562);
    layer1_outputs(508) <= not((layer0_outputs(132)) and (layer0_outputs(2902)));
    layer1_outputs(509) <= not(layer0_outputs(9207));
    layer1_outputs(510) <= (layer0_outputs(9102)) xor (layer0_outputs(5056));
    layer1_outputs(511) <= not(layer0_outputs(7670)) or (layer0_outputs(3448));
    layer1_outputs(512) <= not((layer0_outputs(10103)) or (layer0_outputs(4658)));
    layer1_outputs(513) <= not(layer0_outputs(12746)) or (layer0_outputs(8956));
    layer1_outputs(514) <= not(layer0_outputs(2768)) or (layer0_outputs(203));
    layer1_outputs(515) <= layer0_outputs(10338);
    layer1_outputs(516) <= (layer0_outputs(4427)) and not (layer0_outputs(3994));
    layer1_outputs(517) <= layer0_outputs(1728);
    layer1_outputs(518) <= not(layer0_outputs(11686));
    layer1_outputs(519) <= not((layer0_outputs(1445)) xor (layer0_outputs(5168)));
    layer1_outputs(520) <= (layer0_outputs(412)) and (layer0_outputs(10843));
    layer1_outputs(521) <= (layer0_outputs(1940)) xor (layer0_outputs(3560));
    layer1_outputs(522) <= not(layer0_outputs(9314)) or (layer0_outputs(6306));
    layer1_outputs(523) <= (layer0_outputs(7480)) xor (layer0_outputs(11944));
    layer1_outputs(524) <= (layer0_outputs(6691)) xor (layer0_outputs(9140));
    layer1_outputs(525) <= not(layer0_outputs(7534));
    layer1_outputs(526) <= not(layer0_outputs(6));
    layer1_outputs(527) <= not((layer0_outputs(7526)) or (layer0_outputs(7104)));
    layer1_outputs(528) <= '1';
    layer1_outputs(529) <= layer0_outputs(2459);
    layer1_outputs(530) <= not(layer0_outputs(5622)) or (layer0_outputs(5732));
    layer1_outputs(531) <= layer0_outputs(8311);
    layer1_outputs(532) <= layer0_outputs(2882);
    layer1_outputs(533) <= not(layer0_outputs(8223));
    layer1_outputs(534) <= not(layer0_outputs(1281));
    layer1_outputs(535) <= layer0_outputs(5389);
    layer1_outputs(536) <= (layer0_outputs(8656)) xor (layer0_outputs(3974));
    layer1_outputs(537) <= '0';
    layer1_outputs(538) <= not(layer0_outputs(4319));
    layer1_outputs(539) <= not((layer0_outputs(1821)) or (layer0_outputs(7378)));
    layer1_outputs(540) <= layer0_outputs(3567);
    layer1_outputs(541) <= not((layer0_outputs(2626)) xor (layer0_outputs(2272)));
    layer1_outputs(542) <= (layer0_outputs(2688)) and not (layer0_outputs(3096));
    layer1_outputs(543) <= layer0_outputs(9628);
    layer1_outputs(544) <= not(layer0_outputs(11967));
    layer1_outputs(545) <= not(layer0_outputs(8929));
    layer1_outputs(546) <= '1';
    layer1_outputs(547) <= (layer0_outputs(943)) xor (layer0_outputs(10067));
    layer1_outputs(548) <= (layer0_outputs(1502)) and not (layer0_outputs(4964));
    layer1_outputs(549) <= not(layer0_outputs(8170)) or (layer0_outputs(9752));
    layer1_outputs(550) <= (layer0_outputs(329)) xor (layer0_outputs(12120));
    layer1_outputs(551) <= (layer0_outputs(1680)) and not (layer0_outputs(1284));
    layer1_outputs(552) <= layer0_outputs(2578);
    layer1_outputs(553) <= not((layer0_outputs(3269)) xor (layer0_outputs(5825)));
    layer1_outputs(554) <= not(layer0_outputs(2100));
    layer1_outputs(555) <= (layer0_outputs(1569)) and not (layer0_outputs(6046));
    layer1_outputs(556) <= (layer0_outputs(5084)) xor (layer0_outputs(5798));
    layer1_outputs(557) <= '0';
    layer1_outputs(558) <= not(layer0_outputs(6333)) or (layer0_outputs(2985));
    layer1_outputs(559) <= not(layer0_outputs(4998));
    layer1_outputs(560) <= (layer0_outputs(5725)) and (layer0_outputs(7874));
    layer1_outputs(561) <= layer0_outputs(7643);
    layer1_outputs(562) <= not(layer0_outputs(10621)) or (layer0_outputs(7867));
    layer1_outputs(563) <= (layer0_outputs(6628)) and (layer0_outputs(683));
    layer1_outputs(564) <= not(layer0_outputs(9531));
    layer1_outputs(565) <= (layer0_outputs(1143)) and not (layer0_outputs(6333));
    layer1_outputs(566) <= not(layer0_outputs(11224)) or (layer0_outputs(4035));
    layer1_outputs(567) <= not((layer0_outputs(4164)) xor (layer0_outputs(5906)));
    layer1_outputs(568) <= not(layer0_outputs(1347));
    layer1_outputs(569) <= not(layer0_outputs(10025));
    layer1_outputs(570) <= not(layer0_outputs(10832));
    layer1_outputs(571) <= not(layer0_outputs(9898));
    layer1_outputs(572) <= (layer0_outputs(3828)) xor (layer0_outputs(12660));
    layer1_outputs(573) <= layer0_outputs(1278);
    layer1_outputs(574) <= not((layer0_outputs(6079)) xor (layer0_outputs(10707)));
    layer1_outputs(575) <= not((layer0_outputs(12329)) xor (layer0_outputs(7055)));
    layer1_outputs(576) <= not((layer0_outputs(7945)) or (layer0_outputs(10235)));
    layer1_outputs(577) <= not((layer0_outputs(11090)) or (layer0_outputs(11685)));
    layer1_outputs(578) <= not(layer0_outputs(682)) or (layer0_outputs(5144));
    layer1_outputs(579) <= (layer0_outputs(3099)) and not (layer0_outputs(4330));
    layer1_outputs(580) <= not((layer0_outputs(6560)) and (layer0_outputs(9228)));
    layer1_outputs(581) <= (layer0_outputs(5891)) xor (layer0_outputs(10144));
    layer1_outputs(582) <= not(layer0_outputs(6349));
    layer1_outputs(583) <= (layer0_outputs(9916)) and not (layer0_outputs(3602));
    layer1_outputs(584) <= (layer0_outputs(12687)) and not (layer0_outputs(10246));
    layer1_outputs(585) <= not((layer0_outputs(3616)) xor (layer0_outputs(10806)));
    layer1_outputs(586) <= not(layer0_outputs(12418)) or (layer0_outputs(1211));
    layer1_outputs(587) <= layer0_outputs(7198);
    layer1_outputs(588) <= not(layer0_outputs(4505));
    layer1_outputs(589) <= (layer0_outputs(9054)) or (layer0_outputs(8699));
    layer1_outputs(590) <= layer0_outputs(6885);
    layer1_outputs(591) <= not(layer0_outputs(1139));
    layer1_outputs(592) <= (layer0_outputs(513)) and not (layer0_outputs(9735));
    layer1_outputs(593) <= not(layer0_outputs(10200));
    layer1_outputs(594) <= not((layer0_outputs(9065)) xor (layer0_outputs(2802)));
    layer1_outputs(595) <= not((layer0_outputs(1236)) xor (layer0_outputs(11409)));
    layer1_outputs(596) <= (layer0_outputs(7221)) and not (layer0_outputs(2903));
    layer1_outputs(597) <= not(layer0_outputs(3037));
    layer1_outputs(598) <= (layer0_outputs(5359)) and (layer0_outputs(3251));
    layer1_outputs(599) <= layer0_outputs(7928);
    layer1_outputs(600) <= not(layer0_outputs(599));
    layer1_outputs(601) <= (layer0_outputs(884)) and (layer0_outputs(6705));
    layer1_outputs(602) <= layer0_outputs(5715);
    layer1_outputs(603) <= not(layer0_outputs(2982));
    layer1_outputs(604) <= layer0_outputs(6049);
    layer1_outputs(605) <= (layer0_outputs(8495)) and not (layer0_outputs(3168));
    layer1_outputs(606) <= (layer0_outputs(10550)) and not (layer0_outputs(3904));
    layer1_outputs(607) <= not(layer0_outputs(424));
    layer1_outputs(608) <= not(layer0_outputs(1242)) or (layer0_outputs(4951));
    layer1_outputs(609) <= not((layer0_outputs(5409)) xor (layer0_outputs(8821)));
    layer1_outputs(610) <= not((layer0_outputs(12464)) and (layer0_outputs(12144)));
    layer1_outputs(611) <= not(layer0_outputs(7570));
    layer1_outputs(612) <= not(layer0_outputs(9593)) or (layer0_outputs(5097));
    layer1_outputs(613) <= not(layer0_outputs(3207));
    layer1_outputs(614) <= not(layer0_outputs(5911));
    layer1_outputs(615) <= layer0_outputs(9551);
    layer1_outputs(616) <= '0';
    layer1_outputs(617) <= layer0_outputs(9518);
    layer1_outputs(618) <= not(layer0_outputs(1036));
    layer1_outputs(619) <= '0';
    layer1_outputs(620) <= layer0_outputs(6132);
    layer1_outputs(621) <= (layer0_outputs(9922)) and (layer0_outputs(9737));
    layer1_outputs(622) <= layer0_outputs(10638);
    layer1_outputs(623) <= not((layer0_outputs(11398)) or (layer0_outputs(10424)));
    layer1_outputs(624) <= layer0_outputs(12339);
    layer1_outputs(625) <= not(layer0_outputs(6109)) or (layer0_outputs(11898));
    layer1_outputs(626) <= layer0_outputs(6354);
    layer1_outputs(627) <= not(layer0_outputs(5503));
    layer1_outputs(628) <= not((layer0_outputs(11731)) xor (layer0_outputs(3154)));
    layer1_outputs(629) <= not(layer0_outputs(11673)) or (layer0_outputs(10511));
    layer1_outputs(630) <= not(layer0_outputs(12529));
    layer1_outputs(631) <= (layer0_outputs(6483)) and (layer0_outputs(9712));
    layer1_outputs(632) <= layer0_outputs(9369);
    layer1_outputs(633) <= (layer0_outputs(2613)) or (layer0_outputs(6871));
    layer1_outputs(634) <= (layer0_outputs(1752)) and (layer0_outputs(3958));
    layer1_outputs(635) <= not(layer0_outputs(6345));
    layer1_outputs(636) <= (layer0_outputs(2140)) xor (layer0_outputs(631));
    layer1_outputs(637) <= not((layer0_outputs(6705)) and (layer0_outputs(1742)));
    layer1_outputs(638) <= layer0_outputs(4182);
    layer1_outputs(639) <= (layer0_outputs(8195)) and not (layer0_outputs(4969));
    layer1_outputs(640) <= layer0_outputs(9871);
    layer1_outputs(641) <= (layer0_outputs(4765)) and not (layer0_outputs(5088));
    layer1_outputs(642) <= (layer0_outputs(6279)) xor (layer0_outputs(12456));
    layer1_outputs(643) <= (layer0_outputs(2448)) or (layer0_outputs(1582));
    layer1_outputs(644) <= not((layer0_outputs(6439)) and (layer0_outputs(9382)));
    layer1_outputs(645) <= not(layer0_outputs(11714));
    layer1_outputs(646) <= (layer0_outputs(12311)) and not (layer0_outputs(4304));
    layer1_outputs(647) <= (layer0_outputs(11294)) xor (layer0_outputs(11722));
    layer1_outputs(648) <= layer0_outputs(6189);
    layer1_outputs(649) <= not(layer0_outputs(5114)) or (layer0_outputs(11179));
    layer1_outputs(650) <= not(layer0_outputs(10096));
    layer1_outputs(651) <= layer0_outputs(6488);
    layer1_outputs(652) <= not(layer0_outputs(5274));
    layer1_outputs(653) <= not(layer0_outputs(3935)) or (layer0_outputs(11087));
    layer1_outputs(654) <= not(layer0_outputs(8860)) or (layer0_outputs(9410));
    layer1_outputs(655) <= (layer0_outputs(2290)) and not (layer0_outputs(7640));
    layer1_outputs(656) <= not(layer0_outputs(10191));
    layer1_outputs(657) <= (layer0_outputs(3179)) xor (layer0_outputs(6859));
    layer1_outputs(658) <= (layer0_outputs(7878)) xor (layer0_outputs(9491));
    layer1_outputs(659) <= (layer0_outputs(1315)) and not (layer0_outputs(9420));
    layer1_outputs(660) <= (layer0_outputs(3300)) xor (layer0_outputs(758));
    layer1_outputs(661) <= (layer0_outputs(2523)) xor (layer0_outputs(885));
    layer1_outputs(662) <= not((layer0_outputs(12444)) or (layer0_outputs(5683)));
    layer1_outputs(663) <= not(layer0_outputs(9624)) or (layer0_outputs(3667));
    layer1_outputs(664) <= layer0_outputs(9765);
    layer1_outputs(665) <= not((layer0_outputs(8842)) or (layer0_outputs(6864)));
    layer1_outputs(666) <= '1';
    layer1_outputs(667) <= not(layer0_outputs(10349));
    layer1_outputs(668) <= (layer0_outputs(7671)) and (layer0_outputs(6252));
    layer1_outputs(669) <= not((layer0_outputs(3868)) or (layer0_outputs(6789)));
    layer1_outputs(670) <= (layer0_outputs(8020)) and not (layer0_outputs(3853));
    layer1_outputs(671) <= not((layer0_outputs(7504)) and (layer0_outputs(10588)));
    layer1_outputs(672) <= layer0_outputs(416);
    layer1_outputs(673) <= not(layer0_outputs(5219));
    layer1_outputs(674) <= layer0_outputs(10760);
    layer1_outputs(675) <= not((layer0_outputs(9004)) or (layer0_outputs(7675)));
    layer1_outputs(676) <= not(layer0_outputs(1694));
    layer1_outputs(677) <= layer0_outputs(11053);
    layer1_outputs(678) <= not((layer0_outputs(7549)) xor (layer0_outputs(7608)));
    layer1_outputs(679) <= layer0_outputs(8302);
    layer1_outputs(680) <= not(layer0_outputs(12383)) or (layer0_outputs(4928));
    layer1_outputs(681) <= not((layer0_outputs(9131)) and (layer0_outputs(9235)));
    layer1_outputs(682) <= (layer0_outputs(7744)) and not (layer0_outputs(10427));
    layer1_outputs(683) <= not(layer0_outputs(9463));
    layer1_outputs(684) <= not((layer0_outputs(12754)) or (layer0_outputs(2953)));
    layer1_outputs(685) <= layer0_outputs(2145);
    layer1_outputs(686) <= (layer0_outputs(813)) and (layer0_outputs(2231));
    layer1_outputs(687) <= '1';
    layer1_outputs(688) <= not(layer0_outputs(6089));
    layer1_outputs(689) <= (layer0_outputs(10218)) and (layer0_outputs(3861));
    layer1_outputs(690) <= not(layer0_outputs(9850));
    layer1_outputs(691) <= layer0_outputs(6771);
    layer1_outputs(692) <= layer0_outputs(9949);
    layer1_outputs(693) <= not(layer0_outputs(12775)) or (layer0_outputs(6877));
    layer1_outputs(694) <= (layer0_outputs(12589)) xor (layer0_outputs(513));
    layer1_outputs(695) <= not(layer0_outputs(10933));
    layer1_outputs(696) <= (layer0_outputs(5137)) xor (layer0_outputs(868));
    layer1_outputs(697) <= not(layer0_outputs(12756)) or (layer0_outputs(8197));
    layer1_outputs(698) <= (layer0_outputs(3968)) xor (layer0_outputs(8739));
    layer1_outputs(699) <= (layer0_outputs(11713)) and not (layer0_outputs(8088));
    layer1_outputs(700) <= layer0_outputs(7566);
    layer1_outputs(701) <= not(layer0_outputs(2488));
    layer1_outputs(702) <= layer0_outputs(3054);
    layer1_outputs(703) <= not(layer0_outputs(6661)) or (layer0_outputs(7538));
    layer1_outputs(704) <= (layer0_outputs(322)) and not (layer0_outputs(7135));
    layer1_outputs(705) <= not(layer0_outputs(1986));
    layer1_outputs(706) <= not(layer0_outputs(11318));
    layer1_outputs(707) <= layer0_outputs(3311);
    layer1_outputs(708) <= (layer0_outputs(3614)) and not (layer0_outputs(8616));
    layer1_outputs(709) <= not(layer0_outputs(1913)) or (layer0_outputs(9590));
    layer1_outputs(710) <= not(layer0_outputs(5628));
    layer1_outputs(711) <= layer0_outputs(6750);
    layer1_outputs(712) <= not(layer0_outputs(9523));
    layer1_outputs(713) <= not(layer0_outputs(11131));
    layer1_outputs(714) <= not(layer0_outputs(5053));
    layer1_outputs(715) <= (layer0_outputs(7203)) or (layer0_outputs(11905));
    layer1_outputs(716) <= not((layer0_outputs(716)) and (layer0_outputs(7801)));
    layer1_outputs(717) <= (layer0_outputs(3809)) and not (layer0_outputs(12302));
    layer1_outputs(718) <= (layer0_outputs(10432)) and (layer0_outputs(925));
    layer1_outputs(719) <= (layer0_outputs(652)) and (layer0_outputs(5845));
    layer1_outputs(720) <= (layer0_outputs(7017)) and not (layer0_outputs(6492));
    layer1_outputs(721) <= not(layer0_outputs(2311));
    layer1_outputs(722) <= layer0_outputs(5557);
    layer1_outputs(723) <= not(layer0_outputs(4777));
    layer1_outputs(724) <= layer0_outputs(2856);
    layer1_outputs(725) <= not((layer0_outputs(5191)) and (layer0_outputs(2219)));
    layer1_outputs(726) <= not(layer0_outputs(12625));
    layer1_outputs(727) <= layer0_outputs(3176);
    layer1_outputs(728) <= (layer0_outputs(2883)) and not (layer0_outputs(9907));
    layer1_outputs(729) <= not((layer0_outputs(998)) and (layer0_outputs(2986)));
    layer1_outputs(730) <= not((layer0_outputs(10028)) and (layer0_outputs(7798)));
    layer1_outputs(731) <= layer0_outputs(4563);
    layer1_outputs(732) <= not((layer0_outputs(4651)) and (layer0_outputs(3935)));
    layer1_outputs(733) <= not(layer0_outputs(5501));
    layer1_outputs(734) <= '0';
    layer1_outputs(735) <= (layer0_outputs(5495)) and not (layer0_outputs(5303));
    layer1_outputs(736) <= layer0_outputs(7386);
    layer1_outputs(737) <= (layer0_outputs(5049)) or (layer0_outputs(6677));
    layer1_outputs(738) <= (layer0_outputs(4829)) and not (layer0_outputs(12041));
    layer1_outputs(739) <= layer0_outputs(4824);
    layer1_outputs(740) <= not(layer0_outputs(7168)) or (layer0_outputs(698));
    layer1_outputs(741) <= '1';
    layer1_outputs(742) <= not(layer0_outputs(2445)) or (layer0_outputs(74));
    layer1_outputs(743) <= (layer0_outputs(6334)) and not (layer0_outputs(9533));
    layer1_outputs(744) <= not(layer0_outputs(7292)) or (layer0_outputs(12619));
    layer1_outputs(745) <= layer0_outputs(287);
    layer1_outputs(746) <= not(layer0_outputs(2468)) or (layer0_outputs(9219));
    layer1_outputs(747) <= (layer0_outputs(3890)) xor (layer0_outputs(8502));
    layer1_outputs(748) <= not(layer0_outputs(6574));
    layer1_outputs(749) <= (layer0_outputs(1377)) xor (layer0_outputs(2876));
    layer1_outputs(750) <= not((layer0_outputs(8485)) or (layer0_outputs(8710)));
    layer1_outputs(751) <= not(layer0_outputs(635));
    layer1_outputs(752) <= not(layer0_outputs(6881)) or (layer0_outputs(8812));
    layer1_outputs(753) <= (layer0_outputs(5060)) or (layer0_outputs(10485));
    layer1_outputs(754) <= not(layer0_outputs(3660)) or (layer0_outputs(6129));
    layer1_outputs(755) <= not(layer0_outputs(4888));
    layer1_outputs(756) <= not(layer0_outputs(1702));
    layer1_outputs(757) <= not(layer0_outputs(3318));
    layer1_outputs(758) <= not((layer0_outputs(1713)) and (layer0_outputs(98)));
    layer1_outputs(759) <= layer0_outputs(1971);
    layer1_outputs(760) <= (layer0_outputs(12010)) and (layer0_outputs(10977));
    layer1_outputs(761) <= (layer0_outputs(8377)) and not (layer0_outputs(8760));
    layer1_outputs(762) <= (layer0_outputs(4262)) and not (layer0_outputs(5921));
    layer1_outputs(763) <= not(layer0_outputs(10065)) or (layer0_outputs(3555));
    layer1_outputs(764) <= (layer0_outputs(6119)) xor (layer0_outputs(8590));
    layer1_outputs(765) <= not(layer0_outputs(2186)) or (layer0_outputs(10121));
    layer1_outputs(766) <= (layer0_outputs(10818)) xor (layer0_outputs(4311));
    layer1_outputs(767) <= not((layer0_outputs(10185)) or (layer0_outputs(11919)));
    layer1_outputs(768) <= (layer0_outputs(360)) and not (layer0_outputs(4533));
    layer1_outputs(769) <= layer0_outputs(6058);
    layer1_outputs(770) <= not((layer0_outputs(5629)) xor (layer0_outputs(10617)));
    layer1_outputs(771) <= not(layer0_outputs(3385));
    layer1_outputs(772) <= not(layer0_outputs(2629)) or (layer0_outputs(3257));
    layer1_outputs(773) <= not(layer0_outputs(2726));
    layer1_outputs(774) <= layer0_outputs(1637);
    layer1_outputs(775) <= (layer0_outputs(5515)) and (layer0_outputs(6245));
    layer1_outputs(776) <= not((layer0_outputs(6527)) or (layer0_outputs(8334)));
    layer1_outputs(777) <= layer0_outputs(7848);
    layer1_outputs(778) <= layer0_outputs(12615);
    layer1_outputs(779) <= (layer0_outputs(5664)) and not (layer0_outputs(10523));
    layer1_outputs(780) <= (layer0_outputs(1045)) or (layer0_outputs(10277));
    layer1_outputs(781) <= not((layer0_outputs(6228)) xor (layer0_outputs(8597)));
    layer1_outputs(782) <= layer0_outputs(2803);
    layer1_outputs(783) <= not(layer0_outputs(5366)) or (layer0_outputs(8985));
    layer1_outputs(784) <= layer0_outputs(2563);
    layer1_outputs(785) <= layer0_outputs(3443);
    layer1_outputs(786) <= (layer0_outputs(4971)) xor (layer0_outputs(2651));
    layer1_outputs(787) <= not(layer0_outputs(1153));
    layer1_outputs(788) <= layer0_outputs(12211);
    layer1_outputs(789) <= not(layer0_outputs(12008));
    layer1_outputs(790) <= (layer0_outputs(3293)) xor (layer0_outputs(3631));
    layer1_outputs(791) <= not(layer0_outputs(7266));
    layer1_outputs(792) <= (layer0_outputs(3165)) xor (layer0_outputs(3047));
    layer1_outputs(793) <= (layer0_outputs(7740)) and not (layer0_outputs(2172));
    layer1_outputs(794) <= not((layer0_outputs(10182)) or (layer0_outputs(6793)));
    layer1_outputs(795) <= not((layer0_outputs(7682)) or (layer0_outputs(2497)));
    layer1_outputs(796) <= layer0_outputs(10227);
    layer1_outputs(797) <= layer0_outputs(11057);
    layer1_outputs(798) <= layer0_outputs(5269);
    layer1_outputs(799) <= not(layer0_outputs(12656)) or (layer0_outputs(10315));
    layer1_outputs(800) <= (layer0_outputs(10119)) and not (layer0_outputs(8384));
    layer1_outputs(801) <= layer0_outputs(6054);
    layer1_outputs(802) <= layer0_outputs(12601);
    layer1_outputs(803) <= not(layer0_outputs(2369)) or (layer0_outputs(6160));
    layer1_outputs(804) <= not((layer0_outputs(7529)) or (layer0_outputs(6964)));
    layer1_outputs(805) <= (layer0_outputs(1030)) and not (layer0_outputs(1628));
    layer1_outputs(806) <= (layer0_outputs(9175)) and (layer0_outputs(8220));
    layer1_outputs(807) <= not(layer0_outputs(12637));
    layer1_outputs(808) <= layer0_outputs(9105);
    layer1_outputs(809) <= not((layer0_outputs(2848)) or (layer0_outputs(364)));
    layer1_outputs(810) <= layer0_outputs(1761);
    layer1_outputs(811) <= layer0_outputs(10958);
    layer1_outputs(812) <= not(layer0_outputs(6710));
    layer1_outputs(813) <= not(layer0_outputs(5595)) or (layer0_outputs(3775));
    layer1_outputs(814) <= (layer0_outputs(6404)) and not (layer0_outputs(1605));
    layer1_outputs(815) <= not(layer0_outputs(390));
    layer1_outputs(816) <= layer0_outputs(9243);
    layer1_outputs(817) <= (layer0_outputs(2096)) and (layer0_outputs(3513));
    layer1_outputs(818) <= '0';
    layer1_outputs(819) <= not(layer0_outputs(1054));
    layer1_outputs(820) <= (layer0_outputs(1701)) xor (layer0_outputs(8966));
    layer1_outputs(821) <= not((layer0_outputs(218)) xor (layer0_outputs(5607)));
    layer1_outputs(822) <= not((layer0_outputs(8825)) xor (layer0_outputs(5272)));
    layer1_outputs(823) <= layer0_outputs(7617);
    layer1_outputs(824) <= not(layer0_outputs(6580));
    layer1_outputs(825) <= not((layer0_outputs(5199)) and (layer0_outputs(10555)));
    layer1_outputs(826) <= layer0_outputs(8088);
    layer1_outputs(827) <= not(layer0_outputs(4994));
    layer1_outputs(828) <= not((layer0_outputs(10559)) or (layer0_outputs(1856)));
    layer1_outputs(829) <= (layer0_outputs(9114)) and (layer0_outputs(1454));
    layer1_outputs(830) <= (layer0_outputs(4176)) and not (layer0_outputs(4328));
    layer1_outputs(831) <= layer0_outputs(123);
    layer1_outputs(832) <= not(layer0_outputs(7815)) or (layer0_outputs(2416));
    layer1_outputs(833) <= layer0_outputs(10377);
    layer1_outputs(834) <= (layer0_outputs(1158)) xor (layer0_outputs(10868));
    layer1_outputs(835) <= layer0_outputs(12410);
    layer1_outputs(836) <= not(layer0_outputs(7517));
    layer1_outputs(837) <= not(layer0_outputs(2827));
    layer1_outputs(838) <= not(layer0_outputs(10026)) or (layer0_outputs(5720));
    layer1_outputs(839) <= not(layer0_outputs(6788)) or (layer0_outputs(9394));
    layer1_outputs(840) <= not((layer0_outputs(6495)) or (layer0_outputs(5646)));
    layer1_outputs(841) <= layer0_outputs(5904);
    layer1_outputs(842) <= not(layer0_outputs(12433));
    layer1_outputs(843) <= not(layer0_outputs(7284)) or (layer0_outputs(1427));
    layer1_outputs(844) <= layer0_outputs(10173);
    layer1_outputs(845) <= (layer0_outputs(11421)) and (layer0_outputs(10753));
    layer1_outputs(846) <= not((layer0_outputs(2114)) xor (layer0_outputs(5342)));
    layer1_outputs(847) <= layer0_outputs(3489);
    layer1_outputs(848) <= not(layer0_outputs(3724));
    layer1_outputs(849) <= (layer0_outputs(3362)) and not (layer0_outputs(5893));
    layer1_outputs(850) <= '1';
    layer1_outputs(851) <= not(layer0_outputs(7900));
    layer1_outputs(852) <= not(layer0_outputs(8957));
    layer1_outputs(853) <= not(layer0_outputs(8520)) or (layer0_outputs(4894));
    layer1_outputs(854) <= (layer0_outputs(8304)) and not (layer0_outputs(1890));
    layer1_outputs(855) <= not(layer0_outputs(1800));
    layer1_outputs(856) <= not(layer0_outputs(7092));
    layer1_outputs(857) <= (layer0_outputs(5863)) xor (layer0_outputs(8516));
    layer1_outputs(858) <= layer0_outputs(11737);
    layer1_outputs(859) <= not(layer0_outputs(10653));
    layer1_outputs(860) <= not((layer0_outputs(7213)) or (layer0_outputs(1068)));
    layer1_outputs(861) <= not(layer0_outputs(8344));
    layer1_outputs(862) <= (layer0_outputs(8647)) or (layer0_outputs(8493));
    layer1_outputs(863) <= not(layer0_outputs(487));
    layer1_outputs(864) <= layer0_outputs(4685);
    layer1_outputs(865) <= not(layer0_outputs(12355));
    layer1_outputs(866) <= layer0_outputs(11495);
    layer1_outputs(867) <= layer0_outputs(12218);
    layer1_outputs(868) <= not(layer0_outputs(185)) or (layer0_outputs(2025));
    layer1_outputs(869) <= not(layer0_outputs(2066));
    layer1_outputs(870) <= layer0_outputs(3082);
    layer1_outputs(871) <= not((layer0_outputs(1009)) and (layer0_outputs(2608)));
    layer1_outputs(872) <= not(layer0_outputs(6680)) or (layer0_outputs(5981));
    layer1_outputs(873) <= layer0_outputs(10245);
    layer1_outputs(874) <= layer0_outputs(11781);
    layer1_outputs(875) <= not((layer0_outputs(62)) or (layer0_outputs(6307)));
    layer1_outputs(876) <= layer0_outputs(11587);
    layer1_outputs(877) <= (layer0_outputs(4090)) or (layer0_outputs(3637));
    layer1_outputs(878) <= (layer0_outputs(5345)) xor (layer0_outputs(2704));
    layer1_outputs(879) <= layer0_outputs(8649);
    layer1_outputs(880) <= not(layer0_outputs(1412));
    layer1_outputs(881) <= layer0_outputs(3105);
    layer1_outputs(882) <= layer0_outputs(12727);
    layer1_outputs(883) <= not((layer0_outputs(8675)) and (layer0_outputs(5173)));
    layer1_outputs(884) <= layer0_outputs(6791);
    layer1_outputs(885) <= layer0_outputs(6225);
    layer1_outputs(886) <= not(layer0_outputs(6622));
    layer1_outputs(887) <= not(layer0_outputs(11522));
    layer1_outputs(888) <= not((layer0_outputs(993)) or (layer0_outputs(1361)));
    layer1_outputs(889) <= not((layer0_outputs(10207)) xor (layer0_outputs(4688)));
    layer1_outputs(890) <= (layer0_outputs(7105)) and (layer0_outputs(17));
    layer1_outputs(891) <= not(layer0_outputs(3634));
    layer1_outputs(892) <= not(layer0_outputs(7978));
    layer1_outputs(893) <= (layer0_outputs(10882)) and not (layer0_outputs(6966));
    layer1_outputs(894) <= not(layer0_outputs(11409));
    layer1_outputs(895) <= layer0_outputs(5025);
    layer1_outputs(896) <= not((layer0_outputs(10862)) xor (layer0_outputs(12306)));
    layer1_outputs(897) <= (layer0_outputs(7420)) or (layer0_outputs(2116));
    layer1_outputs(898) <= layer0_outputs(887);
    layer1_outputs(899) <= not((layer0_outputs(12254)) or (layer0_outputs(9291)));
    layer1_outputs(900) <= not((layer0_outputs(11471)) xor (layer0_outputs(5836)));
    layer1_outputs(901) <= (layer0_outputs(10901)) xor (layer0_outputs(790));
    layer1_outputs(902) <= not((layer0_outputs(12264)) or (layer0_outputs(1810)));
    layer1_outputs(903) <= not(layer0_outputs(4948));
    layer1_outputs(904) <= (layer0_outputs(7340)) or (layer0_outputs(5148));
    layer1_outputs(905) <= (layer0_outputs(1520)) and not (layer0_outputs(4933));
    layer1_outputs(906) <= not(layer0_outputs(5626));
    layer1_outputs(907) <= (layer0_outputs(612)) and (layer0_outputs(2291));
    layer1_outputs(908) <= (layer0_outputs(398)) xor (layer0_outputs(7761));
    layer1_outputs(909) <= (layer0_outputs(1666)) or (layer0_outputs(5196));
    layer1_outputs(910) <= layer0_outputs(3316);
    layer1_outputs(911) <= (layer0_outputs(4157)) or (layer0_outputs(9789));
    layer1_outputs(912) <= not((layer0_outputs(3954)) xor (layer0_outputs(9451)));
    layer1_outputs(913) <= not(layer0_outputs(8472));
    layer1_outputs(914) <= layer0_outputs(8831);
    layer1_outputs(915) <= (layer0_outputs(12564)) and not (layer0_outputs(8114));
    layer1_outputs(916) <= (layer0_outputs(8900)) and not (layer0_outputs(12446));
    layer1_outputs(917) <= not((layer0_outputs(9549)) and (layer0_outputs(5301)));
    layer1_outputs(918) <= (layer0_outputs(4660)) and not (layer0_outputs(6364));
    layer1_outputs(919) <= (layer0_outputs(5638)) and not (layer0_outputs(12335));
    layer1_outputs(920) <= not(layer0_outputs(10130)) or (layer0_outputs(9789));
    layer1_outputs(921) <= (layer0_outputs(5759)) or (layer0_outputs(9748));
    layer1_outputs(922) <= layer0_outputs(5333);
    layer1_outputs(923) <= not(layer0_outputs(8204)) or (layer0_outputs(9129));
    layer1_outputs(924) <= layer0_outputs(5814);
    layer1_outputs(925) <= (layer0_outputs(8312)) and not (layer0_outputs(3012));
    layer1_outputs(926) <= (layer0_outputs(6041)) and not (layer0_outputs(7637));
    layer1_outputs(927) <= layer0_outputs(4900);
    layer1_outputs(928) <= not((layer0_outputs(6212)) and (layer0_outputs(6654)));
    layer1_outputs(929) <= (layer0_outputs(8202)) and not (layer0_outputs(5686));
    layer1_outputs(930) <= layer0_outputs(11229);
    layer1_outputs(931) <= layer0_outputs(10613);
    layer1_outputs(932) <= (layer0_outputs(6449)) and not (layer0_outputs(1819));
    layer1_outputs(933) <= not((layer0_outputs(11185)) or (layer0_outputs(11395)));
    layer1_outputs(934) <= not(layer0_outputs(12492)) or (layer0_outputs(6549));
    layer1_outputs(935) <= layer0_outputs(8667);
    layer1_outputs(936) <= not((layer0_outputs(2809)) and (layer0_outputs(4718)));
    layer1_outputs(937) <= not(layer0_outputs(4076));
    layer1_outputs(938) <= not((layer0_outputs(11410)) xor (layer0_outputs(11633)));
    layer1_outputs(939) <= layer0_outputs(1583);
    layer1_outputs(940) <= (layer0_outputs(882)) or (layer0_outputs(897));
    layer1_outputs(941) <= not(layer0_outputs(7278)) or (layer0_outputs(8203));
    layer1_outputs(942) <= not((layer0_outputs(6887)) xor (layer0_outputs(11376)));
    layer1_outputs(943) <= not(layer0_outputs(2188));
    layer1_outputs(944) <= not((layer0_outputs(5687)) or (layer0_outputs(7893)));
    layer1_outputs(945) <= not(layer0_outputs(9128));
    layer1_outputs(946) <= layer0_outputs(5804);
    layer1_outputs(947) <= layer0_outputs(2365);
    layer1_outputs(948) <= not(layer0_outputs(9841));
    layer1_outputs(949) <= not(layer0_outputs(12679));
    layer1_outputs(950) <= (layer0_outputs(4836)) or (layer0_outputs(7817));
    layer1_outputs(951) <= not((layer0_outputs(8581)) and (layer0_outputs(1364)));
    layer1_outputs(952) <= layer0_outputs(3254);
    layer1_outputs(953) <= (layer0_outputs(8270)) or (layer0_outputs(12685));
    layer1_outputs(954) <= not(layer0_outputs(929));
    layer1_outputs(955) <= layer0_outputs(5932);
    layer1_outputs(956) <= (layer0_outputs(1172)) and not (layer0_outputs(11912));
    layer1_outputs(957) <= (layer0_outputs(3792)) or (layer0_outputs(4861));
    layer1_outputs(958) <= (layer0_outputs(7419)) and not (layer0_outputs(7776));
    layer1_outputs(959) <= '0';
    layer1_outputs(960) <= (layer0_outputs(7209)) and not (layer0_outputs(11394));
    layer1_outputs(961) <= (layer0_outputs(5289)) and not (layer0_outputs(12678));
    layer1_outputs(962) <= not(layer0_outputs(5480)) or (layer0_outputs(11611));
    layer1_outputs(963) <= (layer0_outputs(7783)) or (layer0_outputs(7655));
    layer1_outputs(964) <= not(layer0_outputs(9630));
    layer1_outputs(965) <= (layer0_outputs(6703)) or (layer0_outputs(7155));
    layer1_outputs(966) <= layer0_outputs(8163);
    layer1_outputs(967) <= (layer0_outputs(9578)) or (layer0_outputs(879));
    layer1_outputs(968) <= (layer0_outputs(7417)) or (layer0_outputs(12598));
    layer1_outputs(969) <= not(layer0_outputs(9870));
    layer1_outputs(970) <= (layer0_outputs(11256)) and not (layer0_outputs(6899));
    layer1_outputs(971) <= '1';
    layer1_outputs(972) <= not(layer0_outputs(12412));
    layer1_outputs(973) <= (layer0_outputs(8330)) and not (layer0_outputs(11183));
    layer1_outputs(974) <= not(layer0_outputs(1987)) or (layer0_outputs(8679));
    layer1_outputs(975) <= (layer0_outputs(1611)) or (layer0_outputs(11996));
    layer1_outputs(976) <= (layer0_outputs(1163)) and not (layer0_outputs(9799));
    layer1_outputs(977) <= layer0_outputs(10701);
    layer1_outputs(978) <= (layer0_outputs(3696)) and not (layer0_outputs(9304));
    layer1_outputs(979) <= not((layer0_outputs(11132)) xor (layer0_outputs(2508)));
    layer1_outputs(980) <= not(layer0_outputs(11259)) or (layer0_outputs(3417));
    layer1_outputs(981) <= layer0_outputs(1902);
    layer1_outputs(982) <= (layer0_outputs(2836)) and not (layer0_outputs(4457));
    layer1_outputs(983) <= not(layer0_outputs(6857));
    layer1_outputs(984) <= not(layer0_outputs(6869));
    layer1_outputs(985) <= layer0_outputs(5011);
    layer1_outputs(986) <= (layer0_outputs(6844)) xor (layer0_outputs(12222));
    layer1_outputs(987) <= not(layer0_outputs(2414)) or (layer0_outputs(5250));
    layer1_outputs(988) <= (layer0_outputs(8251)) and not (layer0_outputs(1946));
    layer1_outputs(989) <= (layer0_outputs(2957)) and (layer0_outputs(12366));
    layer1_outputs(990) <= (layer0_outputs(4919)) and (layer0_outputs(3349));
    layer1_outputs(991) <= (layer0_outputs(8026)) xor (layer0_outputs(4801));
    layer1_outputs(992) <= not(layer0_outputs(5614)) or (layer0_outputs(6619));
    layer1_outputs(993) <= '1';
    layer1_outputs(994) <= (layer0_outputs(11743)) and not (layer0_outputs(1582));
    layer1_outputs(995) <= not(layer0_outputs(1499)) or (layer0_outputs(6182));
    layer1_outputs(996) <= not((layer0_outputs(2514)) or (layer0_outputs(5110)));
    layer1_outputs(997) <= not(layer0_outputs(7811));
    layer1_outputs(998) <= layer0_outputs(2274);
    layer1_outputs(999) <= layer0_outputs(1504);
    layer1_outputs(1000) <= '0';
    layer1_outputs(1001) <= not(layer0_outputs(793)) or (layer0_outputs(6888));
    layer1_outputs(1002) <= (layer0_outputs(11444)) xor (layer0_outputs(3141));
    layer1_outputs(1003) <= (layer0_outputs(2352)) and not (layer0_outputs(11148));
    layer1_outputs(1004) <= not((layer0_outputs(2622)) xor (layer0_outputs(4122)));
    layer1_outputs(1005) <= (layer0_outputs(3942)) and (layer0_outputs(12252));
    layer1_outputs(1006) <= not(layer0_outputs(8621)) or (layer0_outputs(4795));
    layer1_outputs(1007) <= (layer0_outputs(7647)) and (layer0_outputs(3999));
    layer1_outputs(1008) <= (layer0_outputs(7461)) and not (layer0_outputs(4385));
    layer1_outputs(1009) <= layer0_outputs(6634);
    layer1_outputs(1010) <= not(layer0_outputs(11017));
    layer1_outputs(1011) <= layer0_outputs(2837);
    layer1_outputs(1012) <= not(layer0_outputs(7550)) or (layer0_outputs(9890));
    layer1_outputs(1013) <= layer0_outputs(12499);
    layer1_outputs(1014) <= (layer0_outputs(5456)) and not (layer0_outputs(7654));
    layer1_outputs(1015) <= not(layer0_outputs(8744)) or (layer0_outputs(8623));
    layer1_outputs(1016) <= not((layer0_outputs(10488)) or (layer0_outputs(6231)));
    layer1_outputs(1017) <= (layer0_outputs(7991)) and (layer0_outputs(878));
    layer1_outputs(1018) <= not(layer0_outputs(1320));
    layer1_outputs(1019) <= (layer0_outputs(9619)) or (layer0_outputs(5734));
    layer1_outputs(1020) <= (layer0_outputs(4371)) or (layer0_outputs(7512));
    layer1_outputs(1021) <= (layer0_outputs(5315)) and not (layer0_outputs(2935));
    layer1_outputs(1022) <= not(layer0_outputs(2452));
    layer1_outputs(1023) <= not(layer0_outputs(11545)) or (layer0_outputs(6438));
    layer1_outputs(1024) <= not((layer0_outputs(1362)) xor (layer0_outputs(6027)));
    layer1_outputs(1025) <= layer0_outputs(10810);
    layer1_outputs(1026) <= layer0_outputs(1781);
    layer1_outputs(1027) <= layer0_outputs(11974);
    layer1_outputs(1028) <= not(layer0_outputs(12375));
    layer1_outputs(1029) <= (layer0_outputs(3011)) and (layer0_outputs(12237));
    layer1_outputs(1030) <= not(layer0_outputs(952));
    layer1_outputs(1031) <= not(layer0_outputs(1363)) or (layer0_outputs(9067));
    layer1_outputs(1032) <= (layer0_outputs(1774)) xor (layer0_outputs(2167));
    layer1_outputs(1033) <= not((layer0_outputs(9161)) or (layer0_outputs(9123)));
    layer1_outputs(1034) <= not(layer0_outputs(12289));
    layer1_outputs(1035) <= (layer0_outputs(12532)) xor (layer0_outputs(7660));
    layer1_outputs(1036) <= (layer0_outputs(1209)) and (layer0_outputs(445));
    layer1_outputs(1037) <= layer0_outputs(10948);
    layer1_outputs(1038) <= not(layer0_outputs(6696));
    layer1_outputs(1039) <= (layer0_outputs(4043)) or (layer0_outputs(2909));
    layer1_outputs(1040) <= layer0_outputs(2423);
    layer1_outputs(1041) <= not((layer0_outputs(4236)) xor (layer0_outputs(6005)));
    layer1_outputs(1042) <= not(layer0_outputs(4830)) or (layer0_outputs(7660));
    layer1_outputs(1043) <= not(layer0_outputs(11742)) or (layer0_outputs(1445));
    layer1_outputs(1044) <= not(layer0_outputs(11029));
    layer1_outputs(1045) <= not(layer0_outputs(5054));
    layer1_outputs(1046) <= layer0_outputs(226);
    layer1_outputs(1047) <= not((layer0_outputs(3230)) and (layer0_outputs(12141)));
    layer1_outputs(1048) <= not(layer0_outputs(11019)) or (layer0_outputs(9389));
    layer1_outputs(1049) <= layer0_outputs(11067);
    layer1_outputs(1050) <= not((layer0_outputs(2990)) and (layer0_outputs(4729)));
    layer1_outputs(1051) <= (layer0_outputs(532)) xor (layer0_outputs(7636));
    layer1_outputs(1052) <= layer0_outputs(3781);
    layer1_outputs(1053) <= layer0_outputs(4994);
    layer1_outputs(1054) <= not((layer0_outputs(7682)) or (layer0_outputs(11381)));
    layer1_outputs(1055) <= '1';
    layer1_outputs(1056) <= layer0_outputs(7326);
    layer1_outputs(1057) <= (layer0_outputs(5708)) and not (layer0_outputs(9320));
    layer1_outputs(1058) <= not(layer0_outputs(10103)) or (layer0_outputs(853));
    layer1_outputs(1059) <= not(layer0_outputs(11140));
    layer1_outputs(1060) <= (layer0_outputs(2577)) and not (layer0_outputs(8019));
    layer1_outputs(1061) <= layer0_outputs(12070);
    layer1_outputs(1062) <= (layer0_outputs(6400)) and not (layer0_outputs(9556));
    layer1_outputs(1063) <= layer0_outputs(9919);
    layer1_outputs(1064) <= layer0_outputs(1088);
    layer1_outputs(1065) <= (layer0_outputs(3428)) and not (layer0_outputs(4690));
    layer1_outputs(1066) <= not(layer0_outputs(10382)) or (layer0_outputs(10881));
    layer1_outputs(1067) <= not(layer0_outputs(5933)) or (layer0_outputs(4864));
    layer1_outputs(1068) <= layer0_outputs(2605);
    layer1_outputs(1069) <= layer0_outputs(7255);
    layer1_outputs(1070) <= (layer0_outputs(8684)) and not (layer0_outputs(1610));
    layer1_outputs(1071) <= not(layer0_outputs(8032)) or (layer0_outputs(1113));
    layer1_outputs(1072) <= not(layer0_outputs(12616)) or (layer0_outputs(3238));
    layer1_outputs(1073) <= layer0_outputs(9489);
    layer1_outputs(1074) <= layer0_outputs(9348);
    layer1_outputs(1075) <= layer0_outputs(395);
    layer1_outputs(1076) <= layer0_outputs(3383);
    layer1_outputs(1077) <= layer0_outputs(11315);
    layer1_outputs(1078) <= (layer0_outputs(505)) xor (layer0_outputs(12691));
    layer1_outputs(1079) <= not(layer0_outputs(4310));
    layer1_outputs(1080) <= not((layer0_outputs(9109)) xor (layer0_outputs(6461)));
    layer1_outputs(1081) <= (layer0_outputs(5263)) and not (layer0_outputs(9412));
    layer1_outputs(1082) <= not((layer0_outputs(8111)) xor (layer0_outputs(6666)));
    layer1_outputs(1083) <= not(layer0_outputs(4458)) or (layer0_outputs(8916));
    layer1_outputs(1084) <= not((layer0_outputs(2330)) or (layer0_outputs(3679)));
    layer1_outputs(1085) <= (layer0_outputs(4849)) and (layer0_outputs(12670));
    layer1_outputs(1086) <= (layer0_outputs(3231)) xor (layer0_outputs(11768));
    layer1_outputs(1087) <= not(layer0_outputs(5553));
    layer1_outputs(1088) <= not((layer0_outputs(941)) or (layer0_outputs(6106)));
    layer1_outputs(1089) <= (layer0_outputs(4001)) xor (layer0_outputs(11512));
    layer1_outputs(1090) <= not(layer0_outputs(1298));
    layer1_outputs(1091) <= not((layer0_outputs(4667)) or (layer0_outputs(9221)));
    layer1_outputs(1092) <= not((layer0_outputs(10305)) and (layer0_outputs(2686)));
    layer1_outputs(1093) <= not(layer0_outputs(10767));
    layer1_outputs(1094) <= not(layer0_outputs(3460));
    layer1_outputs(1095) <= (layer0_outputs(6142)) and not (layer0_outputs(2194));
    layer1_outputs(1096) <= not((layer0_outputs(6867)) xor (layer0_outputs(10516)));
    layer1_outputs(1097) <= not(layer0_outputs(3142));
    layer1_outputs(1098) <= (layer0_outputs(948)) and not (layer0_outputs(12159));
    layer1_outputs(1099) <= layer0_outputs(5236);
    layer1_outputs(1100) <= not(layer0_outputs(11480));
    layer1_outputs(1101) <= (layer0_outputs(6260)) or (layer0_outputs(8008));
    layer1_outputs(1102) <= (layer0_outputs(6428)) and not (layer0_outputs(5804));
    layer1_outputs(1103) <= layer0_outputs(3113);
    layer1_outputs(1104) <= (layer0_outputs(353)) and not (layer0_outputs(6548));
    layer1_outputs(1105) <= not(layer0_outputs(2382));
    layer1_outputs(1106) <= not(layer0_outputs(10841)) or (layer0_outputs(4252));
    layer1_outputs(1107) <= (layer0_outputs(6826)) xor (layer0_outputs(7083));
    layer1_outputs(1108) <= (layer0_outputs(6133)) and (layer0_outputs(7184));
    layer1_outputs(1109) <= not(layer0_outputs(3496));
    layer1_outputs(1110) <= (layer0_outputs(7853)) and not (layer0_outputs(10196));
    layer1_outputs(1111) <= not((layer0_outputs(12330)) xor (layer0_outputs(8046)));
    layer1_outputs(1112) <= not(layer0_outputs(5371));
    layer1_outputs(1113) <= layer0_outputs(7762);
    layer1_outputs(1114) <= (layer0_outputs(2923)) or (layer0_outputs(12184));
    layer1_outputs(1115) <= (layer0_outputs(12376)) xor (layer0_outputs(1752));
    layer1_outputs(1116) <= not((layer0_outputs(8477)) and (layer0_outputs(1386)));
    layer1_outputs(1117) <= (layer0_outputs(5527)) xor (layer0_outputs(9866));
    layer1_outputs(1118) <= layer0_outputs(3339);
    layer1_outputs(1119) <= (layer0_outputs(1240)) xor (layer0_outputs(3031));
    layer1_outputs(1120) <= not(layer0_outputs(11014));
    layer1_outputs(1121) <= not((layer0_outputs(4136)) and (layer0_outputs(4791)));
    layer1_outputs(1122) <= layer0_outputs(4356);
    layer1_outputs(1123) <= (layer0_outputs(11568)) and not (layer0_outputs(10962));
    layer1_outputs(1124) <= (layer0_outputs(11012)) xor (layer0_outputs(11245));
    layer1_outputs(1125) <= not((layer0_outputs(7866)) and (layer0_outputs(7230)));
    layer1_outputs(1126) <= layer0_outputs(2605);
    layer1_outputs(1127) <= layer0_outputs(5091);
    layer1_outputs(1128) <= not(layer0_outputs(2247));
    layer1_outputs(1129) <= not(layer0_outputs(5990));
    layer1_outputs(1130) <= (layer0_outputs(666)) and not (layer0_outputs(8338));
    layer1_outputs(1131) <= layer0_outputs(8984);
    layer1_outputs(1132) <= not(layer0_outputs(12739)) or (layer0_outputs(6570));
    layer1_outputs(1133) <= not(layer0_outputs(12363));
    layer1_outputs(1134) <= layer0_outputs(4194);
    layer1_outputs(1135) <= not(layer0_outputs(9955)) or (layer0_outputs(9682));
    layer1_outputs(1136) <= (layer0_outputs(8018)) and not (layer0_outputs(8053));
    layer1_outputs(1137) <= (layer0_outputs(11057)) and (layer0_outputs(9524));
    layer1_outputs(1138) <= not((layer0_outputs(2979)) xor (layer0_outputs(954)));
    layer1_outputs(1139) <= not(layer0_outputs(4703));
    layer1_outputs(1140) <= (layer0_outputs(7225)) and not (layer0_outputs(7046));
    layer1_outputs(1141) <= not(layer0_outputs(12394));
    layer1_outputs(1142) <= (layer0_outputs(92)) xor (layer0_outputs(10482));
    layer1_outputs(1143) <= layer0_outputs(6710);
    layer1_outputs(1144) <= (layer0_outputs(11178)) xor (layer0_outputs(2587));
    layer1_outputs(1145) <= not(layer0_outputs(650));
    layer1_outputs(1146) <= not(layer0_outputs(8425));
    layer1_outputs(1147) <= not(layer0_outputs(5340)) or (layer0_outputs(3379));
    layer1_outputs(1148) <= not((layer0_outputs(8592)) or (layer0_outputs(1563)));
    layer1_outputs(1149) <= not(layer0_outputs(3888)) or (layer0_outputs(2353));
    layer1_outputs(1150) <= not((layer0_outputs(5893)) and (layer0_outputs(5564)));
    layer1_outputs(1151) <= not(layer0_outputs(4908)) or (layer0_outputs(11044));
    layer1_outputs(1152) <= not(layer0_outputs(11483));
    layer1_outputs(1153) <= not(layer0_outputs(1632));
    layer1_outputs(1154) <= not((layer0_outputs(8320)) or (layer0_outputs(12286)));
    layer1_outputs(1155) <= not((layer0_outputs(4770)) xor (layer0_outputs(8434)));
    layer1_outputs(1156) <= (layer0_outputs(7108)) and (layer0_outputs(3704));
    layer1_outputs(1157) <= not(layer0_outputs(341));
    layer1_outputs(1158) <= not(layer0_outputs(12758));
    layer1_outputs(1159) <= layer0_outputs(6753);
    layer1_outputs(1160) <= (layer0_outputs(6594)) and not (layer0_outputs(7437));
    layer1_outputs(1161) <= layer0_outputs(232);
    layer1_outputs(1162) <= not((layer0_outputs(2366)) or (layer0_outputs(1297)));
    layer1_outputs(1163) <= not(layer0_outputs(3826));
    layer1_outputs(1164) <= not(layer0_outputs(1371)) or (layer0_outputs(3997));
    layer1_outputs(1165) <= not(layer0_outputs(12504)) or (layer0_outputs(6528));
    layer1_outputs(1166) <= not(layer0_outputs(11955));
    layer1_outputs(1167) <= not((layer0_outputs(9020)) and (layer0_outputs(3591)));
    layer1_outputs(1168) <= not((layer0_outputs(1877)) xor (layer0_outputs(10763)));
    layer1_outputs(1169) <= not(layer0_outputs(10892)) or (layer0_outputs(3607));
    layer1_outputs(1170) <= (layer0_outputs(11250)) or (layer0_outputs(1847));
    layer1_outputs(1171) <= not(layer0_outputs(8864));
    layer1_outputs(1172) <= not((layer0_outputs(10625)) or (layer0_outputs(1574)));
    layer1_outputs(1173) <= not(layer0_outputs(5647)) or (layer0_outputs(6778));
    layer1_outputs(1174) <= layer0_outputs(5694);
    layer1_outputs(1175) <= not(layer0_outputs(9801));
    layer1_outputs(1176) <= (layer0_outputs(10360)) and (layer0_outputs(5580));
    layer1_outputs(1177) <= '1';
    layer1_outputs(1178) <= layer0_outputs(669);
    layer1_outputs(1179) <= (layer0_outputs(8093)) and not (layer0_outputs(10090));
    layer1_outputs(1180) <= (layer0_outputs(11994)) and (layer0_outputs(584));
    layer1_outputs(1181) <= not((layer0_outputs(6300)) and (layer0_outputs(1669)));
    layer1_outputs(1182) <= (layer0_outputs(12382)) and not (layer0_outputs(6581));
    layer1_outputs(1183) <= not(layer0_outputs(9194)) or (layer0_outputs(9708));
    layer1_outputs(1184) <= not(layer0_outputs(5491)) or (layer0_outputs(5901));
    layer1_outputs(1185) <= not((layer0_outputs(1063)) and (layer0_outputs(3804)));
    layer1_outputs(1186) <= (layer0_outputs(4652)) and not (layer0_outputs(5142));
    layer1_outputs(1187) <= layer0_outputs(11068);
    layer1_outputs(1188) <= (layer0_outputs(7843)) xor (layer0_outputs(7243));
    layer1_outputs(1189) <= not((layer0_outputs(12592)) or (layer0_outputs(3796)));
    layer1_outputs(1190) <= (layer0_outputs(3113)) and not (layer0_outputs(4246));
    layer1_outputs(1191) <= not(layer0_outputs(3585)) or (layer0_outputs(5192));
    layer1_outputs(1192) <= layer0_outputs(6944);
    layer1_outputs(1193) <= (layer0_outputs(8528)) or (layer0_outputs(7419));
    layer1_outputs(1194) <= not(layer0_outputs(10411));
    layer1_outputs(1195) <= (layer0_outputs(1868)) and not (layer0_outputs(5402));
    layer1_outputs(1196) <= layer0_outputs(7498);
    layer1_outputs(1197) <= not((layer0_outputs(8798)) xor (layer0_outputs(10928)));
    layer1_outputs(1198) <= (layer0_outputs(9821)) and not (layer0_outputs(5539));
    layer1_outputs(1199) <= (layer0_outputs(69)) and not (layer0_outputs(5610));
    layer1_outputs(1200) <= not((layer0_outputs(4370)) and (layer0_outputs(8415)));
    layer1_outputs(1201) <= layer0_outputs(11155);
    layer1_outputs(1202) <= (layer0_outputs(1382)) and (layer0_outputs(11808));
    layer1_outputs(1203) <= layer0_outputs(1146);
    layer1_outputs(1204) <= layer0_outputs(12238);
    layer1_outputs(1205) <= layer0_outputs(6762);
    layer1_outputs(1206) <= layer0_outputs(4817);
    layer1_outputs(1207) <= not((layer0_outputs(2300)) or (layer0_outputs(721)));
    layer1_outputs(1208) <= (layer0_outputs(2920)) or (layer0_outputs(9460));
    layer1_outputs(1209) <= not((layer0_outputs(3218)) and (layer0_outputs(5611)));
    layer1_outputs(1210) <= not(layer0_outputs(12538));
    layer1_outputs(1211) <= layer0_outputs(5294);
    layer1_outputs(1212) <= not((layer0_outputs(7104)) or (layer0_outputs(5936)));
    layer1_outputs(1213) <= layer0_outputs(7124);
    layer1_outputs(1214) <= layer0_outputs(2748);
    layer1_outputs(1215) <= (layer0_outputs(10729)) and not (layer0_outputs(5457));
    layer1_outputs(1216) <= layer0_outputs(8653);
    layer1_outputs(1217) <= layer0_outputs(5419);
    layer1_outputs(1218) <= (layer0_outputs(10300)) and not (layer0_outputs(2921));
    layer1_outputs(1219) <= (layer0_outputs(2585)) or (layer0_outputs(6131));
    layer1_outputs(1220) <= layer0_outputs(7465);
    layer1_outputs(1221) <= layer0_outputs(725);
    layer1_outputs(1222) <= (layer0_outputs(6105)) xor (layer0_outputs(9289));
    layer1_outputs(1223) <= not(layer0_outputs(5737));
    layer1_outputs(1224) <= '0';
    layer1_outputs(1225) <= not(layer0_outputs(3145)) or (layer0_outputs(8272));
    layer1_outputs(1226) <= not(layer0_outputs(1477));
    layer1_outputs(1227) <= not(layer0_outputs(2644));
    layer1_outputs(1228) <= layer0_outputs(1845);
    layer1_outputs(1229) <= layer0_outputs(5293);
    layer1_outputs(1230) <= not((layer0_outputs(11439)) and (layer0_outputs(3343)));
    layer1_outputs(1231) <= not(layer0_outputs(1689));
    layer1_outputs(1232) <= (layer0_outputs(5493)) and not (layer0_outputs(3967));
    layer1_outputs(1233) <= (layer0_outputs(1513)) and not (layer0_outputs(1777));
    layer1_outputs(1234) <= not((layer0_outputs(2991)) xor (layer0_outputs(2894)));
    layer1_outputs(1235) <= layer0_outputs(11839);
    layer1_outputs(1236) <= not(layer0_outputs(10123)) or (layer0_outputs(5740));
    layer1_outputs(1237) <= not(layer0_outputs(1439));
    layer1_outputs(1238) <= layer0_outputs(9);
    layer1_outputs(1239) <= (layer0_outputs(5274)) xor (layer0_outputs(11488));
    layer1_outputs(1240) <= not(layer0_outputs(1394));
    layer1_outputs(1241) <= not((layer0_outputs(10451)) xor (layer0_outputs(11374)));
    layer1_outputs(1242) <= not((layer0_outputs(6466)) or (layer0_outputs(4009)));
    layer1_outputs(1243) <= not((layer0_outputs(708)) and (layer0_outputs(12593)));
    layer1_outputs(1244) <= not(layer0_outputs(5490)) or (layer0_outputs(5802));
    layer1_outputs(1245) <= not(layer0_outputs(2993));
    layer1_outputs(1246) <= not((layer0_outputs(5586)) or (layer0_outputs(7363)));
    layer1_outputs(1247) <= not((layer0_outputs(6746)) and (layer0_outputs(6219)));
    layer1_outputs(1248) <= not((layer0_outputs(9578)) or (layer0_outputs(11991)));
    layer1_outputs(1249) <= (layer0_outputs(1665)) and not (layer0_outputs(1255));
    layer1_outputs(1250) <= (layer0_outputs(10372)) and not (layer0_outputs(1973));
    layer1_outputs(1251) <= not((layer0_outputs(505)) xor (layer0_outputs(1077)));
    layer1_outputs(1252) <= not((layer0_outputs(7876)) or (layer0_outputs(8355)));
    layer1_outputs(1253) <= not(layer0_outputs(5930)) or (layer0_outputs(9791));
    layer1_outputs(1254) <= layer0_outputs(11133);
    layer1_outputs(1255) <= not(layer0_outputs(3111));
    layer1_outputs(1256) <= layer0_outputs(3848);
    layer1_outputs(1257) <= not((layer0_outputs(2378)) xor (layer0_outputs(11998)));
    layer1_outputs(1258) <= not((layer0_outputs(4874)) and (layer0_outputs(2051)));
    layer1_outputs(1259) <= not(layer0_outputs(8322));
    layer1_outputs(1260) <= not(layer0_outputs(4805)) or (layer0_outputs(2615));
    layer1_outputs(1261) <= not((layer0_outputs(5361)) and (layer0_outputs(9341)));
    layer1_outputs(1262) <= layer0_outputs(10275);
    layer1_outputs(1263) <= not((layer0_outputs(4206)) or (layer0_outputs(5697)));
    layer1_outputs(1264) <= layer0_outputs(12738);
    layer1_outputs(1265) <= (layer0_outputs(3990)) and (layer0_outputs(10720));
    layer1_outputs(1266) <= not(layer0_outputs(5283)) or (layer0_outputs(5593));
    layer1_outputs(1267) <= (layer0_outputs(4118)) and (layer0_outputs(9412));
    layer1_outputs(1268) <= (layer0_outputs(4267)) or (layer0_outputs(12035));
    layer1_outputs(1269) <= not(layer0_outputs(11646)) or (layer0_outputs(9205));
    layer1_outputs(1270) <= (layer0_outputs(3558)) or (layer0_outputs(10062));
    layer1_outputs(1271) <= not((layer0_outputs(12441)) and (layer0_outputs(4187)));
    layer1_outputs(1272) <= (layer0_outputs(6806)) and not (layer0_outputs(7324));
    layer1_outputs(1273) <= not((layer0_outputs(5742)) and (layer0_outputs(764)));
    layer1_outputs(1274) <= not((layer0_outputs(621)) or (layer0_outputs(3976)));
    layer1_outputs(1275) <= (layer0_outputs(8002)) xor (layer0_outputs(4617));
    layer1_outputs(1276) <= layer0_outputs(10149);
    layer1_outputs(1277) <= not(layer0_outputs(9965));
    layer1_outputs(1278) <= (layer0_outputs(5937)) or (layer0_outputs(9209));
    layer1_outputs(1279) <= layer0_outputs(12726);
    layer1_outputs(1280) <= (layer0_outputs(8269)) or (layer0_outputs(8640));
    layer1_outputs(1281) <= layer0_outputs(699);
    layer1_outputs(1282) <= not((layer0_outputs(366)) or (layer0_outputs(1640)));
    layer1_outputs(1283) <= not(layer0_outputs(5542));
    layer1_outputs(1284) <= not(layer0_outputs(251)) or (layer0_outputs(3712));
    layer1_outputs(1285) <= (layer0_outputs(12595)) and (layer0_outputs(11978));
    layer1_outputs(1286) <= layer0_outputs(4335);
    layer1_outputs(1287) <= not((layer0_outputs(12631)) or (layer0_outputs(5445)));
    layer1_outputs(1288) <= (layer0_outputs(10877)) or (layer0_outputs(3920));
    layer1_outputs(1289) <= layer0_outputs(10862);
    layer1_outputs(1290) <= (layer0_outputs(8805)) or (layer0_outputs(9295));
    layer1_outputs(1291) <= not(layer0_outputs(996));
    layer1_outputs(1292) <= layer0_outputs(11322);
    layer1_outputs(1293) <= not(layer0_outputs(4308));
    layer1_outputs(1294) <= (layer0_outputs(4437)) and (layer0_outputs(7778));
    layer1_outputs(1295) <= (layer0_outputs(5838)) and not (layer0_outputs(10022));
    layer1_outputs(1296) <= not(layer0_outputs(5815));
    layer1_outputs(1297) <= (layer0_outputs(4599)) and not (layer0_outputs(12295));
    layer1_outputs(1298) <= '1';
    layer1_outputs(1299) <= layer0_outputs(11564);
    layer1_outputs(1300) <= layer0_outputs(9534);
    layer1_outputs(1301) <= not(layer0_outputs(7018)) or (layer0_outputs(3455));
    layer1_outputs(1302) <= not(layer0_outputs(12158)) or (layer0_outputs(6749));
    layer1_outputs(1303) <= not(layer0_outputs(2039)) or (layer0_outputs(2852));
    layer1_outputs(1304) <= not((layer0_outputs(1259)) or (layer0_outputs(4751)));
    layer1_outputs(1305) <= layer0_outputs(678);
    layer1_outputs(1306) <= not((layer0_outputs(5685)) and (layer0_outputs(4746)));
    layer1_outputs(1307) <= (layer0_outputs(7953)) and not (layer0_outputs(7676));
    layer1_outputs(1308) <= not(layer0_outputs(6812)) or (layer0_outputs(1409));
    layer1_outputs(1309) <= layer0_outputs(2945);
    layer1_outputs(1310) <= not(layer0_outputs(5941));
    layer1_outputs(1311) <= (layer0_outputs(7927)) xor (layer0_outputs(6462));
    layer1_outputs(1312) <= not((layer0_outputs(1688)) or (layer0_outputs(470)));
    layer1_outputs(1313) <= not(layer0_outputs(6529));
    layer1_outputs(1314) <= (layer0_outputs(10014)) and not (layer0_outputs(2777));
    layer1_outputs(1315) <= not(layer0_outputs(1704));
    layer1_outputs(1316) <= layer0_outputs(4453);
    layer1_outputs(1317) <= (layer0_outputs(263)) and (layer0_outputs(9447));
    layer1_outputs(1318) <= (layer0_outputs(12772)) and not (layer0_outputs(665));
    layer1_outputs(1319) <= not(layer0_outputs(5088));
    layer1_outputs(1320) <= (layer0_outputs(12297)) xor (layer0_outputs(7621));
    layer1_outputs(1321) <= not(layer0_outputs(11844));
    layer1_outputs(1322) <= not(layer0_outputs(3391)) or (layer0_outputs(10713));
    layer1_outputs(1323) <= not((layer0_outputs(2697)) and (layer0_outputs(3243)));
    layer1_outputs(1324) <= not(layer0_outputs(8320)) or (layer0_outputs(725));
    layer1_outputs(1325) <= layer0_outputs(11787);
    layer1_outputs(1326) <= not(layer0_outputs(1653));
    layer1_outputs(1327) <= not((layer0_outputs(5725)) or (layer0_outputs(2805)));
    layer1_outputs(1328) <= not((layer0_outputs(1475)) xor (layer0_outputs(4093)));
    layer1_outputs(1329) <= not((layer0_outputs(3528)) xor (layer0_outputs(9515)));
    layer1_outputs(1330) <= not(layer0_outputs(2220));
    layer1_outputs(1331) <= not((layer0_outputs(3003)) or (layer0_outputs(2340)));
    layer1_outputs(1332) <= (layer0_outputs(4369)) and not (layer0_outputs(12606));
    layer1_outputs(1333) <= not((layer0_outputs(10260)) or (layer0_outputs(1539)));
    layer1_outputs(1334) <= (layer0_outputs(6926)) or (layer0_outputs(11735));
    layer1_outputs(1335) <= layer0_outputs(664);
    layer1_outputs(1336) <= not(layer0_outputs(861));
    layer1_outputs(1337) <= (layer0_outputs(8559)) or (layer0_outputs(9833));
    layer1_outputs(1338) <= not(layer0_outputs(3150)) or (layer0_outputs(5027));
    layer1_outputs(1339) <= not(layer0_outputs(7654)) or (layer0_outputs(11114));
    layer1_outputs(1340) <= not((layer0_outputs(7645)) and (layer0_outputs(890)));
    layer1_outputs(1341) <= layer0_outputs(8563);
    layer1_outputs(1342) <= not((layer0_outputs(3989)) or (layer0_outputs(11418)));
    layer1_outputs(1343) <= not((layer0_outputs(8616)) or (layer0_outputs(7829)));
    layer1_outputs(1344) <= (layer0_outputs(1969)) xor (layer0_outputs(5474));
    layer1_outputs(1345) <= not(layer0_outputs(11761)) or (layer0_outputs(2461));
    layer1_outputs(1346) <= not((layer0_outputs(9777)) and (layer0_outputs(6088)));
    layer1_outputs(1347) <= layer0_outputs(12461);
    layer1_outputs(1348) <= not(layer0_outputs(6433));
    layer1_outputs(1349) <= not(layer0_outputs(1460));
    layer1_outputs(1350) <= not(layer0_outputs(6882));
    layer1_outputs(1351) <= not(layer0_outputs(3040));
    layer1_outputs(1352) <= '0';
    layer1_outputs(1353) <= (layer0_outputs(12276)) xor (layer0_outputs(8166));
    layer1_outputs(1354) <= not((layer0_outputs(10985)) and (layer0_outputs(2871)));
    layer1_outputs(1355) <= not(layer0_outputs(8217));
    layer1_outputs(1356) <= not(layer0_outputs(265));
    layer1_outputs(1357) <= not(layer0_outputs(2114));
    layer1_outputs(1358) <= not((layer0_outputs(10189)) or (layer0_outputs(11692)));
    layer1_outputs(1359) <= not((layer0_outputs(11006)) and (layer0_outputs(7576)));
    layer1_outputs(1360) <= not(layer0_outputs(5928));
    layer1_outputs(1361) <= '0';
    layer1_outputs(1362) <= layer0_outputs(4662);
    layer1_outputs(1363) <= layer0_outputs(347);
    layer1_outputs(1364) <= (layer0_outputs(6195)) or (layer0_outputs(8949));
    layer1_outputs(1365) <= (layer0_outputs(1956)) and not (layer0_outputs(4028));
    layer1_outputs(1366) <= not((layer0_outputs(3017)) and (layer0_outputs(8668)));
    layer1_outputs(1367) <= not(layer0_outputs(8346));
    layer1_outputs(1368) <= (layer0_outputs(8907)) xor (layer0_outputs(12040));
    layer1_outputs(1369) <= (layer0_outputs(191)) or (layer0_outputs(5003));
    layer1_outputs(1370) <= layer0_outputs(6693);
    layer1_outputs(1371) <= layer0_outputs(8772);
    layer1_outputs(1372) <= (layer0_outputs(11621)) or (layer0_outputs(10910));
    layer1_outputs(1373) <= layer0_outputs(6734);
    layer1_outputs(1374) <= (layer0_outputs(7837)) and not (layer0_outputs(9395));
    layer1_outputs(1375) <= '0';
    layer1_outputs(1376) <= (layer0_outputs(10818)) and (layer0_outputs(12337));
    layer1_outputs(1377) <= layer0_outputs(5217);
    layer1_outputs(1378) <= not(layer0_outputs(4821));
    layer1_outputs(1379) <= layer0_outputs(10171);
    layer1_outputs(1380) <= not(layer0_outputs(8725));
    layer1_outputs(1381) <= (layer0_outputs(8124)) xor (layer0_outputs(8092));
    layer1_outputs(1382) <= (layer0_outputs(9557)) and not (layer0_outputs(4098));
    layer1_outputs(1383) <= layer0_outputs(2967);
    layer1_outputs(1384) <= layer0_outputs(8795);
    layer1_outputs(1385) <= layer0_outputs(12733);
    layer1_outputs(1386) <= (layer0_outputs(6479)) and (layer0_outputs(2400));
    layer1_outputs(1387) <= layer0_outputs(11556);
    layer1_outputs(1388) <= layer0_outputs(7575);
    layer1_outputs(1389) <= not(layer0_outputs(6363));
    layer1_outputs(1390) <= (layer0_outputs(11578)) and not (layer0_outputs(8874));
    layer1_outputs(1391) <= not(layer0_outputs(1269)) or (layer0_outputs(11749));
    layer1_outputs(1392) <= not(layer0_outputs(8413)) or (layer0_outputs(1527));
    layer1_outputs(1393) <= layer0_outputs(12556);
    layer1_outputs(1394) <= not(layer0_outputs(10034));
    layer1_outputs(1395) <= not(layer0_outputs(4102));
    layer1_outputs(1396) <= not((layer0_outputs(10501)) and (layer0_outputs(11917)));
    layer1_outputs(1397) <= not((layer0_outputs(1768)) and (layer0_outputs(8725)));
    layer1_outputs(1398) <= layer0_outputs(12032);
    layer1_outputs(1399) <= (layer0_outputs(4567)) xor (layer0_outputs(7965));
    layer1_outputs(1400) <= (layer0_outputs(2094)) and not (layer0_outputs(1404));
    layer1_outputs(1401) <= (layer0_outputs(2569)) and not (layer0_outputs(5569));
    layer1_outputs(1402) <= not(layer0_outputs(12671));
    layer1_outputs(1403) <= layer0_outputs(8993);
    layer1_outputs(1404) <= not(layer0_outputs(7877));
    layer1_outputs(1405) <= layer0_outputs(11776);
    layer1_outputs(1406) <= not(layer0_outputs(1732)) or (layer0_outputs(12735));
    layer1_outputs(1407) <= (layer0_outputs(2341)) and not (layer0_outputs(2056));
    layer1_outputs(1408) <= not((layer0_outputs(1359)) and (layer0_outputs(7361)));
    layer1_outputs(1409) <= not((layer0_outputs(6848)) and (layer0_outputs(6538)));
    layer1_outputs(1410) <= '1';
    layer1_outputs(1411) <= (layer0_outputs(2285)) xor (layer0_outputs(927));
    layer1_outputs(1412) <= not(layer0_outputs(2576)) or (layer0_outputs(7209));
    layer1_outputs(1413) <= not(layer0_outputs(7477));
    layer1_outputs(1414) <= (layer0_outputs(1700)) xor (layer0_outputs(11396));
    layer1_outputs(1415) <= '1';
    layer1_outputs(1416) <= layer0_outputs(1944);
    layer1_outputs(1417) <= not(layer0_outputs(11025)) or (layer0_outputs(8090));
    layer1_outputs(1418) <= not(layer0_outputs(12428));
    layer1_outputs(1419) <= not(layer0_outputs(6000)) or (layer0_outputs(10134));
    layer1_outputs(1420) <= not(layer0_outputs(9217));
    layer1_outputs(1421) <= not((layer0_outputs(4464)) or (layer0_outputs(4944)));
    layer1_outputs(1422) <= (layer0_outputs(11597)) and (layer0_outputs(10729));
    layer1_outputs(1423) <= not(layer0_outputs(9003));
    layer1_outputs(1424) <= not(layer0_outputs(6490));
    layer1_outputs(1425) <= (layer0_outputs(3162)) and not (layer0_outputs(5187));
    layer1_outputs(1426) <= not(layer0_outputs(10607));
    layer1_outputs(1427) <= (layer0_outputs(6807)) and not (layer0_outputs(7392));
    layer1_outputs(1428) <= layer0_outputs(1646);
    layer1_outputs(1429) <= layer0_outputs(4143);
    layer1_outputs(1430) <= not(layer0_outputs(1846));
    layer1_outputs(1431) <= not(layer0_outputs(8727));
    layer1_outputs(1432) <= layer0_outputs(5069);
    layer1_outputs(1433) <= layer0_outputs(338);
    layer1_outputs(1434) <= not(layer0_outputs(11264));
    layer1_outputs(1435) <= layer0_outputs(1984);
    layer1_outputs(1436) <= not(layer0_outputs(6606));
    layer1_outputs(1437) <= layer0_outputs(457);
    layer1_outputs(1438) <= not(layer0_outputs(5822));
    layer1_outputs(1439) <= (layer0_outputs(676)) xor (layer0_outputs(4037));
    layer1_outputs(1440) <= (layer0_outputs(12320)) and (layer0_outputs(4501));
    layer1_outputs(1441) <= layer0_outputs(385);
    layer1_outputs(1442) <= (layer0_outputs(2477)) and (layer0_outputs(10281));
    layer1_outputs(1443) <= not((layer0_outputs(4458)) and (layer0_outputs(2714)));
    layer1_outputs(1444) <= layer0_outputs(12424);
    layer1_outputs(1445) <= not(layer0_outputs(8138));
    layer1_outputs(1446) <= '0';
    layer1_outputs(1447) <= layer0_outputs(1832);
    layer1_outputs(1448) <= not(layer0_outputs(1056));
    layer1_outputs(1449) <= (layer0_outputs(11638)) and (layer0_outputs(10441));
    layer1_outputs(1450) <= not(layer0_outputs(7666));
    layer1_outputs(1451) <= not((layer0_outputs(6397)) xor (layer0_outputs(1136)));
    layer1_outputs(1452) <= not(layer0_outputs(10979)) or (layer0_outputs(6315));
    layer1_outputs(1453) <= (layer0_outputs(8362)) and not (layer0_outputs(2889));
    layer1_outputs(1454) <= not(layer0_outputs(6063));
    layer1_outputs(1455) <= (layer0_outputs(12224)) xor (layer0_outputs(9533));
    layer1_outputs(1456) <= (layer0_outputs(9037)) and not (layer0_outputs(4025));
    layer1_outputs(1457) <= not((layer0_outputs(8138)) and (layer0_outputs(2811)));
    layer1_outputs(1458) <= not((layer0_outputs(5448)) or (layer0_outputs(7727)));
    layer1_outputs(1459) <= not(layer0_outputs(2001)) or (layer0_outputs(5509));
    layer1_outputs(1460) <= not((layer0_outputs(12699)) xor (layer0_outputs(12750)));
    layer1_outputs(1461) <= layer0_outputs(6732);
    layer1_outputs(1462) <= layer0_outputs(7181);
    layer1_outputs(1463) <= not(layer0_outputs(1611)) or (layer0_outputs(2942));
    layer1_outputs(1464) <= not(layer0_outputs(6110));
    layer1_outputs(1465) <= layer0_outputs(9181);
    layer1_outputs(1466) <= (layer0_outputs(5609)) and (layer0_outputs(6892));
    layer1_outputs(1467) <= not((layer0_outputs(4347)) xor (layer0_outputs(4856)));
    layer1_outputs(1468) <= (layer0_outputs(12692)) and (layer0_outputs(3973));
    layer1_outputs(1469) <= layer0_outputs(4042);
    layer1_outputs(1470) <= not((layer0_outputs(2835)) xor (layer0_outputs(455)));
    layer1_outputs(1471) <= not(layer0_outputs(6017)) or (layer0_outputs(2062));
    layer1_outputs(1472) <= not(layer0_outputs(5989));
    layer1_outputs(1473) <= not(layer0_outputs(6490));
    layer1_outputs(1474) <= layer0_outputs(5749);
    layer1_outputs(1475) <= not(layer0_outputs(1197)) or (layer0_outputs(11230));
    layer1_outputs(1476) <= not(layer0_outputs(11831));
    layer1_outputs(1477) <= not(layer0_outputs(10117));
    layer1_outputs(1478) <= (layer0_outputs(7677)) and (layer0_outputs(4057));
    layer1_outputs(1479) <= not(layer0_outputs(12276));
    layer1_outputs(1480) <= not(layer0_outputs(3549));
    layer1_outputs(1481) <= (layer0_outputs(752)) and (layer0_outputs(2754));
    layer1_outputs(1482) <= layer0_outputs(692);
    layer1_outputs(1483) <= '0';
    layer1_outputs(1484) <= not((layer0_outputs(12097)) xor (layer0_outputs(9706)));
    layer1_outputs(1485) <= not(layer0_outputs(6417));
    layer1_outputs(1486) <= not(layer0_outputs(1251));
    layer1_outputs(1487) <= (layer0_outputs(3958)) xor (layer0_outputs(5831));
    layer1_outputs(1488) <= (layer0_outputs(10804)) and (layer0_outputs(9819));
    layer1_outputs(1489) <= not((layer0_outputs(1889)) or (layer0_outputs(5604)));
    layer1_outputs(1490) <= layer0_outputs(995);
    layer1_outputs(1491) <= not(layer0_outputs(3163)) or (layer0_outputs(1950));
    layer1_outputs(1492) <= (layer0_outputs(11016)) xor (layer0_outputs(8767));
    layer1_outputs(1493) <= (layer0_outputs(10810)) and not (layer0_outputs(7425));
    layer1_outputs(1494) <= not((layer0_outputs(10242)) or (layer0_outputs(2357)));
    layer1_outputs(1495) <= not(layer0_outputs(5057));
    layer1_outputs(1496) <= not(layer0_outputs(6895));
    layer1_outputs(1497) <= not((layer0_outputs(6158)) and (layer0_outputs(9173)));
    layer1_outputs(1498) <= (layer0_outputs(7912)) and (layer0_outputs(3547));
    layer1_outputs(1499) <= layer0_outputs(4549);
    layer1_outputs(1500) <= not(layer0_outputs(12613)) or (layer0_outputs(10237));
    layer1_outputs(1501) <= (layer0_outputs(769)) or (layer0_outputs(3090));
    layer1_outputs(1502) <= (layer0_outputs(11478)) and not (layer0_outputs(10132));
    layer1_outputs(1503) <= (layer0_outputs(11858)) and not (layer0_outputs(1462));
    layer1_outputs(1504) <= not((layer0_outputs(5055)) and (layer0_outputs(9107)));
    layer1_outputs(1505) <= layer0_outputs(8552);
    layer1_outputs(1506) <= (layer0_outputs(11474)) or (layer0_outputs(33));
    layer1_outputs(1507) <= not(layer0_outputs(6920));
    layer1_outputs(1508) <= not(layer0_outputs(7118));
    layer1_outputs(1509) <= not(layer0_outputs(9513));
    layer1_outputs(1510) <= (layer0_outputs(5510)) and not (layer0_outputs(3965));
    layer1_outputs(1511) <= (layer0_outputs(8761)) or (layer0_outputs(7423));
    layer1_outputs(1512) <= layer0_outputs(2345);
    layer1_outputs(1513) <= not((layer0_outputs(7584)) and (layer0_outputs(6305)));
    layer1_outputs(1514) <= not((layer0_outputs(6998)) and (layer0_outputs(6048)));
    layer1_outputs(1515) <= not(layer0_outputs(10212));
    layer1_outputs(1516) <= (layer0_outputs(9541)) and not (layer0_outputs(4783));
    layer1_outputs(1517) <= not((layer0_outputs(5180)) xor (layer0_outputs(7110)));
    layer1_outputs(1518) <= (layer0_outputs(9609)) and (layer0_outputs(5242));
    layer1_outputs(1519) <= (layer0_outputs(9180)) and not (layer0_outputs(2061));
    layer1_outputs(1520) <= not(layer0_outputs(1805));
    layer1_outputs(1521) <= (layer0_outputs(3884)) and (layer0_outputs(3903));
    layer1_outputs(1522) <= layer0_outputs(10358);
    layer1_outputs(1523) <= (layer0_outputs(10294)) and (layer0_outputs(839));
    layer1_outputs(1524) <= not(layer0_outputs(2690));
    layer1_outputs(1525) <= (layer0_outputs(4543)) xor (layer0_outputs(6457));
    layer1_outputs(1526) <= (layer0_outputs(5412)) and not (layer0_outputs(5762));
    layer1_outputs(1527) <= not(layer0_outputs(9855));
    layer1_outputs(1528) <= (layer0_outputs(4985)) xor (layer0_outputs(7748));
    layer1_outputs(1529) <= layer0_outputs(8371);
    layer1_outputs(1530) <= layer0_outputs(10611);
    layer1_outputs(1531) <= (layer0_outputs(1922)) or (layer0_outputs(10382));
    layer1_outputs(1532) <= (layer0_outputs(7102)) or (layer0_outputs(6711));
    layer1_outputs(1533) <= not(layer0_outputs(9652));
    layer1_outputs(1534) <= not(layer0_outputs(7838));
    layer1_outputs(1535) <= (layer0_outputs(10924)) or (layer0_outputs(1262));
    layer1_outputs(1536) <= not(layer0_outputs(11513));
    layer1_outputs(1537) <= (layer0_outputs(2863)) xor (layer0_outputs(1098));
    layer1_outputs(1538) <= (layer0_outputs(9408)) and not (layer0_outputs(83));
    layer1_outputs(1539) <= layer0_outputs(11563);
    layer1_outputs(1540) <= (layer0_outputs(201)) and not (layer0_outputs(6697));
    layer1_outputs(1541) <= (layer0_outputs(10180)) or (layer0_outputs(10509));
    layer1_outputs(1542) <= (layer0_outputs(4709)) or (layer0_outputs(9118));
    layer1_outputs(1543) <= layer0_outputs(2532);
    layer1_outputs(1544) <= not((layer0_outputs(5760)) and (layer0_outputs(4798)));
    layer1_outputs(1545) <= (layer0_outputs(489)) and not (layer0_outputs(5069));
    layer1_outputs(1546) <= not(layer0_outputs(3799));
    layer1_outputs(1547) <= (layer0_outputs(6733)) and not (layer0_outputs(1734));
    layer1_outputs(1548) <= not(layer0_outputs(6946));
    layer1_outputs(1549) <= not(layer0_outputs(820));
    layer1_outputs(1550) <= (layer0_outputs(311)) and not (layer0_outputs(2375));
    layer1_outputs(1551) <= (layer0_outputs(8263)) and (layer0_outputs(447));
    layer1_outputs(1552) <= not(layer0_outputs(9986)) or (layer0_outputs(9645));
    layer1_outputs(1553) <= not(layer0_outputs(9630));
    layer1_outputs(1554) <= not(layer0_outputs(8288));
    layer1_outputs(1555) <= layer0_outputs(4881);
    layer1_outputs(1556) <= not(layer0_outputs(9828));
    layer1_outputs(1557) <= not(layer0_outputs(8434));
    layer1_outputs(1558) <= not((layer0_outputs(12632)) or (layer0_outputs(3987)));
    layer1_outputs(1559) <= not(layer0_outputs(3815));
    layer1_outputs(1560) <= layer0_outputs(8697);
    layer1_outputs(1561) <= layer0_outputs(1033);
    layer1_outputs(1562) <= layer0_outputs(10331);
    layer1_outputs(1563) <= layer0_outputs(4830);
    layer1_outputs(1564) <= (layer0_outputs(9658)) and (layer0_outputs(10922));
    layer1_outputs(1565) <= (layer0_outputs(404)) and not (layer0_outputs(9028));
    layer1_outputs(1566) <= not((layer0_outputs(11584)) and (layer0_outputs(8557)));
    layer1_outputs(1567) <= layer0_outputs(12708);
    layer1_outputs(1568) <= (layer0_outputs(8294)) and not (layer0_outputs(8888));
    layer1_outputs(1569) <= not(layer0_outputs(5794)) or (layer0_outputs(8838));
    layer1_outputs(1570) <= not((layer0_outputs(9969)) and (layer0_outputs(4926)));
    layer1_outputs(1571) <= not(layer0_outputs(2698));
    layer1_outputs(1572) <= layer0_outputs(15);
    layer1_outputs(1573) <= not((layer0_outputs(4289)) or (layer0_outputs(2690)));
    layer1_outputs(1574) <= layer0_outputs(4895);
    layer1_outputs(1575) <= not((layer0_outputs(4984)) xor (layer0_outputs(3149)));
    layer1_outputs(1576) <= not(layer0_outputs(5667));
    layer1_outputs(1577) <= not(layer0_outputs(6539)) or (layer0_outputs(7860));
    layer1_outputs(1578) <= not(layer0_outputs(221));
    layer1_outputs(1579) <= layer0_outputs(10960);
    layer1_outputs(1580) <= (layer0_outputs(4377)) xor (layer0_outputs(10072));
    layer1_outputs(1581) <= not((layer0_outputs(3031)) or (layer0_outputs(1856)));
    layer1_outputs(1582) <= not(layer0_outputs(8068));
    layer1_outputs(1583) <= not((layer0_outputs(749)) or (layer0_outputs(7256)));
    layer1_outputs(1584) <= not(layer0_outputs(10834));
    layer1_outputs(1585) <= layer0_outputs(4862);
    layer1_outputs(1586) <= layer0_outputs(6943);
    layer1_outputs(1587) <= not(layer0_outputs(2125));
    layer1_outputs(1588) <= (layer0_outputs(4399)) and (layer0_outputs(8923));
    layer1_outputs(1589) <= not(layer0_outputs(4216));
    layer1_outputs(1590) <= not((layer0_outputs(145)) and (layer0_outputs(11956)));
    layer1_outputs(1591) <= not(layer0_outputs(7470));
    layer1_outputs(1592) <= (layer0_outputs(5113)) xor (layer0_outputs(1667));
    layer1_outputs(1593) <= layer0_outputs(4761);
    layer1_outputs(1594) <= not((layer0_outputs(9073)) xor (layer0_outputs(5288)));
    layer1_outputs(1595) <= not(layer0_outputs(6127)) or (layer0_outputs(1528));
    layer1_outputs(1596) <= not(layer0_outputs(229));
    layer1_outputs(1597) <= layer0_outputs(8051);
    layer1_outputs(1598) <= (layer0_outputs(12371)) and not (layer0_outputs(1332));
    layer1_outputs(1599) <= layer0_outputs(10586);
    layer1_outputs(1600) <= not((layer0_outputs(12077)) and (layer0_outputs(10303)));
    layer1_outputs(1601) <= (layer0_outputs(10659)) and not (layer0_outputs(10780));
    layer1_outputs(1602) <= not(layer0_outputs(7428)) or (layer0_outputs(9036));
    layer1_outputs(1603) <= not(layer0_outputs(8264)) or (layer0_outputs(7532));
    layer1_outputs(1604) <= not(layer0_outputs(1807));
    layer1_outputs(1605) <= not(layer0_outputs(4927));
    layer1_outputs(1606) <= not((layer0_outputs(11710)) xor (layer0_outputs(1756)));
    layer1_outputs(1607) <= not(layer0_outputs(6556));
    layer1_outputs(1608) <= (layer0_outputs(10452)) and not (layer0_outputs(759));
    layer1_outputs(1609) <= (layer0_outputs(6907)) and not (layer0_outputs(11374));
    layer1_outputs(1610) <= (layer0_outputs(8289)) or (layer0_outputs(6507));
    layer1_outputs(1611) <= layer0_outputs(12425);
    layer1_outputs(1612) <= not(layer0_outputs(12096));
    layer1_outputs(1613) <= not((layer0_outputs(12762)) or (layer0_outputs(1586)));
    layer1_outputs(1614) <= not((layer0_outputs(10942)) xor (layer0_outputs(12542)));
    layer1_outputs(1615) <= layer0_outputs(9013);
    layer1_outputs(1616) <= not(layer0_outputs(9266));
    layer1_outputs(1617) <= not(layer0_outputs(4398));
    layer1_outputs(1618) <= not(layer0_outputs(12508)) or (layer0_outputs(6696));
    layer1_outputs(1619) <= (layer0_outputs(703)) or (layer0_outputs(8123));
    layer1_outputs(1620) <= layer0_outputs(1211);
    layer1_outputs(1621) <= not((layer0_outputs(5154)) and (layer0_outputs(401)));
    layer1_outputs(1622) <= not(layer0_outputs(579));
    layer1_outputs(1623) <= not(layer0_outputs(9601)) or (layer0_outputs(5332));
    layer1_outputs(1624) <= (layer0_outputs(3704)) or (layer0_outputs(8125));
    layer1_outputs(1625) <= not(layer0_outputs(11449));
    layer1_outputs(1626) <= (layer0_outputs(2010)) or (layer0_outputs(12739));
    layer1_outputs(1627) <= layer0_outputs(6151);
    layer1_outputs(1628) <= not(layer0_outputs(12328));
    layer1_outputs(1629) <= not(layer0_outputs(11441));
    layer1_outputs(1630) <= not(layer0_outputs(10183));
    layer1_outputs(1631) <= not(layer0_outputs(584)) or (layer0_outputs(8618));
    layer1_outputs(1632) <= (layer0_outputs(947)) xor (layer0_outputs(1030));
    layer1_outputs(1633) <= not(layer0_outputs(10393));
    layer1_outputs(1634) <= not(layer0_outputs(12746));
    layer1_outputs(1635) <= layer0_outputs(4837);
    layer1_outputs(1636) <= layer0_outputs(8507);
    layer1_outputs(1637) <= not((layer0_outputs(11390)) xor (layer0_outputs(11007)));
    layer1_outputs(1638) <= not(layer0_outputs(6451)) or (layer0_outputs(6157));
    layer1_outputs(1639) <= (layer0_outputs(10402)) xor (layer0_outputs(11078));
    layer1_outputs(1640) <= not((layer0_outputs(3072)) and (layer0_outputs(11882)));
    layer1_outputs(1641) <= (layer0_outputs(4427)) xor (layer0_outputs(10241));
    layer1_outputs(1642) <= (layer0_outputs(3673)) and not (layer0_outputs(667));
    layer1_outputs(1643) <= not(layer0_outputs(10657)) or (layer0_outputs(4108));
    layer1_outputs(1644) <= (layer0_outputs(11332)) and not (layer0_outputs(6903));
    layer1_outputs(1645) <= layer0_outputs(1674);
    layer1_outputs(1646) <= not(layer0_outputs(4665));
    layer1_outputs(1647) <= not((layer0_outputs(9008)) or (layer0_outputs(831)));
    layer1_outputs(1648) <= not(layer0_outputs(1324));
    layer1_outputs(1649) <= (layer0_outputs(648)) and (layer0_outputs(2513));
    layer1_outputs(1650) <= layer0_outputs(8155);
    layer1_outputs(1651) <= not(layer0_outputs(7730));
    layer1_outputs(1652) <= layer0_outputs(8302);
    layer1_outputs(1653) <= layer0_outputs(9296);
    layer1_outputs(1654) <= (layer0_outputs(3449)) and (layer0_outputs(1321));
    layer1_outputs(1655) <= layer0_outputs(10945);
    layer1_outputs(1656) <= not(layer0_outputs(5617)) or (layer0_outputs(10263));
    layer1_outputs(1657) <= not((layer0_outputs(5782)) xor (layer0_outputs(12312)));
    layer1_outputs(1658) <= layer0_outputs(10598);
    layer1_outputs(1659) <= not(layer0_outputs(2007));
    layer1_outputs(1660) <= not(layer0_outputs(3818));
    layer1_outputs(1661) <= layer0_outputs(2964);
    layer1_outputs(1662) <= not((layer0_outputs(2992)) and (layer0_outputs(7015)));
    layer1_outputs(1663) <= not(layer0_outputs(6413));
    layer1_outputs(1664) <= not(layer0_outputs(11520));
    layer1_outputs(1665) <= not((layer0_outputs(560)) xor (layer0_outputs(12338)));
    layer1_outputs(1666) <= (layer0_outputs(983)) and not (layer0_outputs(6435));
    layer1_outputs(1667) <= not(layer0_outputs(11674));
    layer1_outputs(1668) <= not(layer0_outputs(3411)) or (layer0_outputs(12707));
    layer1_outputs(1669) <= (layer0_outputs(11872)) and not (layer0_outputs(6946));
    layer1_outputs(1670) <= '0';
    layer1_outputs(1671) <= (layer0_outputs(1299)) and (layer0_outputs(1041));
    layer1_outputs(1672) <= layer0_outputs(2726);
    layer1_outputs(1673) <= layer0_outputs(3257);
    layer1_outputs(1674) <= not(layer0_outputs(9163)) or (layer0_outputs(470));
    layer1_outputs(1675) <= not((layer0_outputs(4197)) xor (layer0_outputs(7127)));
    layer1_outputs(1676) <= (layer0_outputs(9479)) and not (layer0_outputs(9157));
    layer1_outputs(1677) <= layer0_outputs(4244);
    layer1_outputs(1678) <= not(layer0_outputs(235));
    layer1_outputs(1679) <= (layer0_outputs(2717)) and not (layer0_outputs(8215));
    layer1_outputs(1680) <= layer0_outputs(9704);
    layer1_outputs(1681) <= (layer0_outputs(5269)) and not (layer0_outputs(2606));
    layer1_outputs(1682) <= (layer0_outputs(3203)) xor (layer0_outputs(8041));
    layer1_outputs(1683) <= layer0_outputs(12225);
    layer1_outputs(1684) <= not(layer0_outputs(2342)) or (layer0_outputs(4285));
    layer1_outputs(1685) <= layer0_outputs(10334);
    layer1_outputs(1686) <= not((layer0_outputs(12364)) or (layer0_outputs(5806)));
    layer1_outputs(1687) <= not(layer0_outputs(1082));
    layer1_outputs(1688) <= not(layer0_outputs(3390));
    layer1_outputs(1689) <= not(layer0_outputs(2256));
    layer1_outputs(1690) <= (layer0_outputs(11205)) and not (layer0_outputs(6994));
    layer1_outputs(1691) <= not(layer0_outputs(2225));
    layer1_outputs(1692) <= (layer0_outputs(4353)) xor (layer0_outputs(102));
    layer1_outputs(1693) <= (layer0_outputs(7986)) or (layer0_outputs(8885));
    layer1_outputs(1694) <= not((layer0_outputs(6508)) xor (layer0_outputs(8071)));
    layer1_outputs(1695) <= layer0_outputs(6558);
    layer1_outputs(1696) <= (layer0_outputs(6624)) and not (layer0_outputs(2374));
    layer1_outputs(1697) <= not(layer0_outputs(4463)) or (layer0_outputs(12272));
    layer1_outputs(1698) <= not(layer0_outputs(2517));
    layer1_outputs(1699) <= (layer0_outputs(12052)) or (layer0_outputs(6257));
    layer1_outputs(1700) <= not(layer0_outputs(8052)) or (layer0_outputs(11663));
    layer1_outputs(1701) <= (layer0_outputs(1279)) and not (layer0_outputs(9204));
    layer1_outputs(1702) <= not(layer0_outputs(11145)) or (layer0_outputs(2631));
    layer1_outputs(1703) <= not((layer0_outputs(11940)) and (layer0_outputs(6827)));
    layer1_outputs(1704) <= not(layer0_outputs(3026)) or (layer0_outputs(3028));
    layer1_outputs(1705) <= not(layer0_outputs(9953));
    layer1_outputs(1706) <= not((layer0_outputs(5985)) or (layer0_outputs(12125)));
    layer1_outputs(1707) <= '1';
    layer1_outputs(1708) <= not(layer0_outputs(9849)) or (layer0_outputs(12064));
    layer1_outputs(1709) <= not(layer0_outputs(12085));
    layer1_outputs(1710) <= layer0_outputs(1912);
    layer1_outputs(1711) <= not(layer0_outputs(4230));
    layer1_outputs(1712) <= not(layer0_outputs(11447));
    layer1_outputs(1713) <= not(layer0_outputs(11570)) or (layer0_outputs(12540));
    layer1_outputs(1714) <= not(layer0_outputs(540));
    layer1_outputs(1715) <= (layer0_outputs(10967)) xor (layer0_outputs(10310));
    layer1_outputs(1716) <= '0';
    layer1_outputs(1717) <= not((layer0_outputs(1872)) or (layer0_outputs(436)));
    layer1_outputs(1718) <= not(layer0_outputs(1921));
    layer1_outputs(1719) <= not(layer0_outputs(8609));
    layer1_outputs(1720) <= layer0_outputs(9868);
    layer1_outputs(1721) <= not(layer0_outputs(10542));
    layer1_outputs(1722) <= layer0_outputs(12677);
    layer1_outputs(1723) <= (layer0_outputs(11175)) and not (layer0_outputs(2741));
    layer1_outputs(1724) <= layer0_outputs(71);
    layer1_outputs(1725) <= not(layer0_outputs(3)) or (layer0_outputs(4512));
    layer1_outputs(1726) <= (layer0_outputs(5138)) and (layer0_outputs(6771));
    layer1_outputs(1727) <= layer0_outputs(9399);
    layer1_outputs(1728) <= not(layer0_outputs(11964));
    layer1_outputs(1729) <= not((layer0_outputs(628)) xor (layer0_outputs(11158)));
    layer1_outputs(1730) <= (layer0_outputs(1202)) xor (layer0_outputs(7331));
    layer1_outputs(1731) <= not(layer0_outputs(4029));
    layer1_outputs(1732) <= (layer0_outputs(10937)) and (layer0_outputs(7354));
    layer1_outputs(1733) <= (layer0_outputs(12719)) and (layer0_outputs(7107));
    layer1_outputs(1734) <= not(layer0_outputs(4496));
    layer1_outputs(1735) <= not(layer0_outputs(10632)) or (layer0_outputs(2367));
    layer1_outputs(1736) <= not(layer0_outputs(2152));
    layer1_outputs(1737) <= layer0_outputs(7923);
    layer1_outputs(1738) <= not(layer0_outputs(10796));
    layer1_outputs(1739) <= not((layer0_outputs(7883)) or (layer0_outputs(972)));
    layer1_outputs(1740) <= not((layer0_outputs(11378)) or (layer0_outputs(9935)));
    layer1_outputs(1741) <= not((layer0_outputs(8523)) or (layer0_outputs(2200)));
    layer1_outputs(1742) <= not(layer0_outputs(3662));
    layer1_outputs(1743) <= not(layer0_outputs(1026));
    layer1_outputs(1744) <= layer0_outputs(11927);
    layer1_outputs(1745) <= not(layer0_outputs(2778)) or (layer0_outputs(12470));
    layer1_outputs(1746) <= layer0_outputs(7499);
    layer1_outputs(1747) <= not(layer0_outputs(11709));
    layer1_outputs(1748) <= not((layer0_outputs(9683)) xor (layer0_outputs(2000)));
    layer1_outputs(1749) <= not((layer0_outputs(762)) xor (layer0_outputs(5511)));
    layer1_outputs(1750) <= (layer0_outputs(4674)) and (layer0_outputs(2795));
    layer1_outputs(1751) <= (layer0_outputs(9582)) and not (layer0_outputs(6));
    layer1_outputs(1752) <= not(layer0_outputs(5108)) or (layer0_outputs(9042));
    layer1_outputs(1753) <= not(layer0_outputs(2499)) or (layer0_outputs(8897));
    layer1_outputs(1754) <= layer0_outputs(1302);
    layer1_outputs(1755) <= not(layer0_outputs(6203));
    layer1_outputs(1756) <= not(layer0_outputs(1795));
    layer1_outputs(1757) <= not((layer0_outputs(11584)) xor (layer0_outputs(574)));
    layer1_outputs(1758) <= (layer0_outputs(4412)) and not (layer0_outputs(4714));
    layer1_outputs(1759) <= (layer0_outputs(3181)) and not (layer0_outputs(10981));
    layer1_outputs(1760) <= not((layer0_outputs(12634)) xor (layer0_outputs(989)));
    layer1_outputs(1761) <= not((layer0_outputs(8950)) and (layer0_outputs(9832)));
    layer1_outputs(1762) <= not((layer0_outputs(7549)) xor (layer0_outputs(9703)));
    layer1_outputs(1763) <= (layer0_outputs(9535)) and not (layer0_outputs(8213));
    layer1_outputs(1764) <= not(layer0_outputs(6530)) or (layer0_outputs(7010));
    layer1_outputs(1765) <= layer0_outputs(599);
    layer1_outputs(1766) <= not(layer0_outputs(8967)) or (layer0_outputs(5044));
    layer1_outputs(1767) <= not(layer0_outputs(3135)) or (layer0_outputs(8562));
    layer1_outputs(1768) <= layer0_outputs(9066);
    layer1_outputs(1769) <= not(layer0_outputs(5638)) or (layer0_outputs(107));
    layer1_outputs(1770) <= not(layer0_outputs(4152));
    layer1_outputs(1771) <= not(layer0_outputs(6030)) or (layer0_outputs(3741));
    layer1_outputs(1772) <= (layer0_outputs(4428)) and (layer0_outputs(11961));
    layer1_outputs(1773) <= not((layer0_outputs(11710)) or (layer0_outputs(8883)));
    layer1_outputs(1774) <= (layer0_outputs(2229)) or (layer0_outputs(3785));
    layer1_outputs(1775) <= not(layer0_outputs(1060));
    layer1_outputs(1776) <= not((layer0_outputs(12273)) xor (layer0_outputs(1851)));
    layer1_outputs(1777) <= layer0_outputs(8840);
    layer1_outputs(1778) <= not(layer0_outputs(5512));
    layer1_outputs(1779) <= not((layer0_outputs(880)) or (layer0_outputs(7525)));
    layer1_outputs(1780) <= '1';
    layer1_outputs(1781) <= layer0_outputs(4137);
    layer1_outputs(1782) <= (layer0_outputs(1844)) and not (layer0_outputs(11127));
    layer1_outputs(1783) <= (layer0_outputs(2672)) or (layer0_outputs(331));
    layer1_outputs(1784) <= (layer0_outputs(510)) or (layer0_outputs(1099));
    layer1_outputs(1785) <= (layer0_outputs(1755)) and not (layer0_outputs(11774));
    layer1_outputs(1786) <= not((layer0_outputs(8326)) xor (layer0_outputs(10257)));
    layer1_outputs(1787) <= (layer0_outputs(5270)) or (layer0_outputs(5095));
    layer1_outputs(1788) <= not(layer0_outputs(3883)) or (layer0_outputs(8119));
    layer1_outputs(1789) <= not(layer0_outputs(12118));
    layer1_outputs(1790) <= not(layer0_outputs(173));
    layer1_outputs(1791) <= not((layer0_outputs(2980)) xor (layer0_outputs(12321)));
    layer1_outputs(1792) <= layer0_outputs(7215);
    layer1_outputs(1793) <= not((layer0_outputs(9012)) or (layer0_outputs(5934)));
    layer1_outputs(1794) <= layer0_outputs(981);
    layer1_outputs(1795) <= (layer0_outputs(5689)) xor (layer0_outputs(4878));
    layer1_outputs(1796) <= not(layer0_outputs(10625));
    layer1_outputs(1797) <= not((layer0_outputs(8394)) and (layer0_outputs(7114)));
    layer1_outputs(1798) <= not(layer0_outputs(6018));
    layer1_outputs(1799) <= not(layer0_outputs(6013));
    layer1_outputs(1800) <= not(layer0_outputs(6723));
    layer1_outputs(1801) <= not((layer0_outputs(11834)) xor (layer0_outputs(4137)));
    layer1_outputs(1802) <= (layer0_outputs(5413)) and (layer0_outputs(11856));
    layer1_outputs(1803) <= not((layer0_outputs(4692)) and (layer0_outputs(10077)));
    layer1_outputs(1804) <= not(layer0_outputs(3014));
    layer1_outputs(1805) <= (layer0_outputs(10073)) and not (layer0_outputs(6655));
    layer1_outputs(1806) <= (layer0_outputs(10009)) and not (layer0_outputs(8953));
    layer1_outputs(1807) <= not(layer0_outputs(10921));
    layer1_outputs(1808) <= (layer0_outputs(11187)) and (layer0_outputs(10224));
    layer1_outputs(1809) <= (layer0_outputs(6877)) and not (layer0_outputs(2017));
    layer1_outputs(1810) <= layer0_outputs(2271);
    layer1_outputs(1811) <= not(layer0_outputs(3726));
    layer1_outputs(1812) <= (layer0_outputs(6884)) xor (layer0_outputs(951));
    layer1_outputs(1813) <= not(layer0_outputs(2115));
    layer1_outputs(1814) <= (layer0_outputs(8752)) and (layer0_outputs(8505));
    layer1_outputs(1815) <= not((layer0_outputs(9885)) and (layer0_outputs(11797)));
    layer1_outputs(1816) <= not(layer0_outputs(620));
    layer1_outputs(1817) <= not((layer0_outputs(672)) xor (layer0_outputs(198)));
    layer1_outputs(1818) <= (layer0_outputs(7998)) and (layer0_outputs(9363));
    layer1_outputs(1819) <= layer0_outputs(2955);
    layer1_outputs(1820) <= (layer0_outputs(2473)) or (layer0_outputs(6870));
    layer1_outputs(1821) <= (layer0_outputs(4775)) and (layer0_outputs(2213));
    layer1_outputs(1822) <= layer0_outputs(12303);
    layer1_outputs(1823) <= not((layer0_outputs(11899)) xor (layer0_outputs(7355)));
    layer1_outputs(1824) <= layer0_outputs(2176);
    layer1_outputs(1825) <= not((layer0_outputs(7486)) xor (layer0_outputs(2117)));
    layer1_outputs(1826) <= (layer0_outputs(5348)) or (layer0_outputs(8408));
    layer1_outputs(1827) <= not(layer0_outputs(10544));
    layer1_outputs(1828) <= (layer0_outputs(2289)) or (layer0_outputs(8290));
    layer1_outputs(1829) <= (layer0_outputs(7534)) or (layer0_outputs(7414));
    layer1_outputs(1830) <= layer0_outputs(12372);
    layer1_outputs(1831) <= layer0_outputs(1199);
    layer1_outputs(1832) <= layer0_outputs(25);
    layer1_outputs(1833) <= (layer0_outputs(2594)) and not (layer0_outputs(506));
    layer1_outputs(1834) <= (layer0_outputs(5684)) and not (layer0_outputs(707));
    layer1_outputs(1835) <= not((layer0_outputs(11033)) xor (layer0_outputs(2027)));
    layer1_outputs(1836) <= not(layer0_outputs(6085)) or (layer0_outputs(9422));
    layer1_outputs(1837) <= (layer0_outputs(4449)) and not (layer0_outputs(5170));
    layer1_outputs(1838) <= not(layer0_outputs(7610));
    layer1_outputs(1839) <= (layer0_outputs(9655)) and not (layer0_outputs(3841));
    layer1_outputs(1840) <= layer0_outputs(1622);
    layer1_outputs(1841) <= not((layer0_outputs(11816)) xor (layer0_outputs(10324)));
    layer1_outputs(1842) <= layer0_outputs(3996);
    layer1_outputs(1843) <= not(layer0_outputs(2381));
    layer1_outputs(1844) <= not(layer0_outputs(6708));
    layer1_outputs(1845) <= (layer0_outputs(12715)) xor (layer0_outputs(6251));
    layer1_outputs(1846) <= layer0_outputs(2738);
    layer1_outputs(1847) <= (layer0_outputs(6874)) xor (layer0_outputs(10458));
    layer1_outputs(1848) <= layer0_outputs(5700);
    layer1_outputs(1849) <= layer0_outputs(6596);
    layer1_outputs(1850) <= (layer0_outputs(2521)) or (layer0_outputs(7372));
    layer1_outputs(1851) <= (layer0_outputs(2295)) and not (layer0_outputs(12627));
    layer1_outputs(1852) <= (layer0_outputs(4623)) or (layer0_outputs(1651));
    layer1_outputs(1853) <= not(layer0_outputs(3154));
    layer1_outputs(1854) <= (layer0_outputs(5862)) and not (layer0_outputs(1131));
    layer1_outputs(1855) <= '1';
    layer1_outputs(1856) <= not(layer0_outputs(2888));
    layer1_outputs(1857) <= not(layer0_outputs(8932)) or (layer0_outputs(9077));
    layer1_outputs(1858) <= not(layer0_outputs(1094));
    layer1_outputs(1859) <= layer0_outputs(540);
    layer1_outputs(1860) <= not(layer0_outputs(2268)) or (layer0_outputs(5840));
    layer1_outputs(1861) <= not((layer0_outputs(7024)) and (layer0_outputs(10178)));
    layer1_outputs(1862) <= not(layer0_outputs(10187)) or (layer0_outputs(1101));
    layer1_outputs(1863) <= (layer0_outputs(11407)) and (layer0_outputs(11549));
    layer1_outputs(1864) <= '0';
    layer1_outputs(1865) <= (layer0_outputs(11339)) and (layer0_outputs(8536));
    layer1_outputs(1866) <= not((layer0_outputs(11317)) or (layer0_outputs(6883)));
    layer1_outputs(1867) <= layer0_outputs(3248);
    layer1_outputs(1868) <= (layer0_outputs(11699)) and not (layer0_outputs(2009));
    layer1_outputs(1869) <= not((layer0_outputs(5012)) xor (layer0_outputs(8551)));
    layer1_outputs(1870) <= (layer0_outputs(2260)) or (layer0_outputs(11237));
    layer1_outputs(1871) <= not(layer0_outputs(3094));
    layer1_outputs(1872) <= not(layer0_outputs(3273));
    layer1_outputs(1873) <= (layer0_outputs(1081)) and not (layer0_outputs(7779));
    layer1_outputs(1874) <= not(layer0_outputs(12712));
    layer1_outputs(1875) <= not((layer0_outputs(2306)) xor (layer0_outputs(10859)));
    layer1_outputs(1876) <= (layer0_outputs(9089)) or (layer0_outputs(5765));
    layer1_outputs(1877) <= not(layer0_outputs(2224));
    layer1_outputs(1878) <= layer0_outputs(5587);
    layer1_outputs(1879) <= not(layer0_outputs(3965)) or (layer0_outputs(9997));
    layer1_outputs(1880) <= (layer0_outputs(5711)) and not (layer0_outputs(356));
    layer1_outputs(1881) <= not((layer0_outputs(9870)) and (layer0_outputs(6039)));
    layer1_outputs(1882) <= (layer0_outputs(180)) and not (layer0_outputs(8568));
    layer1_outputs(1883) <= layer0_outputs(6765);
    layer1_outputs(1884) <= '0';
    layer1_outputs(1885) <= not(layer0_outputs(1682));
    layer1_outputs(1886) <= not(layer0_outputs(2944)) or (layer0_outputs(11648));
    layer1_outputs(1887) <= not(layer0_outputs(2960));
    layer1_outputs(1888) <= not((layer0_outputs(9951)) xor (layer0_outputs(2780)));
    layer1_outputs(1889) <= not(layer0_outputs(11836));
    layer1_outputs(1890) <= not(layer0_outputs(11384));
    layer1_outputs(1891) <= (layer0_outputs(1327)) xor (layer0_outputs(4214));
    layer1_outputs(1892) <= not((layer0_outputs(688)) xor (layer0_outputs(5062)));
    layer1_outputs(1893) <= layer0_outputs(9706);
    layer1_outputs(1894) <= not((layer0_outputs(9805)) or (layer0_outputs(3645)));
    layer1_outputs(1895) <= not(layer0_outputs(9166));
    layer1_outputs(1896) <= not((layer0_outputs(11943)) xor (layer0_outputs(7411)));
    layer1_outputs(1897) <= not(layer0_outputs(8325));
    layer1_outputs(1898) <= layer0_outputs(4952);
    layer1_outputs(1899) <= not(layer0_outputs(4619));
    layer1_outputs(1900) <= not(layer0_outputs(6406));
    layer1_outputs(1901) <= (layer0_outputs(9114)) and not (layer0_outputs(111));
    layer1_outputs(1902) <= layer0_outputs(11507);
    layer1_outputs(1903) <= layer0_outputs(439);
    layer1_outputs(1904) <= (layer0_outputs(3265)) and (layer0_outputs(6098));
    layer1_outputs(1905) <= layer0_outputs(110);
    layer1_outputs(1906) <= not((layer0_outputs(10604)) and (layer0_outputs(10940)));
    layer1_outputs(1907) <= (layer0_outputs(1838)) and not (layer0_outputs(7830));
    layer1_outputs(1908) <= not(layer0_outputs(10328));
    layer1_outputs(1909) <= not(layer0_outputs(2004));
    layer1_outputs(1910) <= (layer0_outputs(3603)) and (layer0_outputs(6140));
    layer1_outputs(1911) <= layer0_outputs(7235);
    layer1_outputs(1912) <= not(layer0_outputs(2041));
    layer1_outputs(1913) <= not(layer0_outputs(9873)) or (layer0_outputs(4893));
    layer1_outputs(1914) <= layer0_outputs(10628);
    layer1_outputs(1915) <= layer0_outputs(8142);
    layer1_outputs(1916) <= not(layer0_outputs(11578));
    layer1_outputs(1917) <= not(layer0_outputs(10964));
    layer1_outputs(1918) <= (layer0_outputs(9560)) and not (layer0_outputs(12569));
    layer1_outputs(1919) <= not(layer0_outputs(9271));
    layer1_outputs(1920) <= not((layer0_outputs(7907)) xor (layer0_outputs(8494)));
    layer1_outputs(1921) <= not(layer0_outputs(11881));
    layer1_outputs(1922) <= not(layer0_outputs(165));
    layer1_outputs(1923) <= not((layer0_outputs(5421)) or (layer0_outputs(4212)));
    layer1_outputs(1924) <= (layer0_outputs(6727)) xor (layer0_outputs(12781));
    layer1_outputs(1925) <= layer0_outputs(4412);
    layer1_outputs(1926) <= (layer0_outputs(7859)) or (layer0_outputs(11252));
    layer1_outputs(1927) <= (layer0_outputs(307)) and not (layer0_outputs(4992));
    layer1_outputs(1928) <= not(layer0_outputs(9950));
    layer1_outputs(1929) <= not(layer0_outputs(10105)) or (layer0_outputs(2377));
    layer1_outputs(1930) <= not(layer0_outputs(7561));
    layer1_outputs(1931) <= '1';
    layer1_outputs(1932) <= (layer0_outputs(7262)) and (layer0_outputs(6999));
    layer1_outputs(1933) <= not(layer0_outputs(7376));
    layer1_outputs(1934) <= '0';
    layer1_outputs(1935) <= not(layer0_outputs(10597)) or (layer0_outputs(6026));
    layer1_outputs(1936) <= layer0_outputs(7981);
    layer1_outputs(1937) <= layer0_outputs(2595);
    layer1_outputs(1938) <= layer0_outputs(8893);
    layer1_outputs(1939) <= not(layer0_outputs(9248));
    layer1_outputs(1940) <= not(layer0_outputs(1601)) or (layer0_outputs(12247));
    layer1_outputs(1941) <= layer0_outputs(6878);
    layer1_outputs(1942) <= not(layer0_outputs(1422));
    layer1_outputs(1943) <= not(layer0_outputs(3978)) or (layer0_outputs(7806));
    layer1_outputs(1944) <= not(layer0_outputs(9778));
    layer1_outputs(1945) <= layer0_outputs(10695);
    layer1_outputs(1946) <= layer0_outputs(3180);
    layer1_outputs(1947) <= not(layer0_outputs(1900));
    layer1_outputs(1948) <= (layer0_outputs(7351)) xor (layer0_outputs(6820));
    layer1_outputs(1949) <= layer0_outputs(12285);
    layer1_outputs(1950) <= (layer0_outputs(3852)) or (layer0_outputs(171));
    layer1_outputs(1951) <= (layer0_outputs(1899)) or (layer0_outputs(8085));
    layer1_outputs(1952) <= layer0_outputs(3511);
    layer1_outputs(1953) <= not(layer0_outputs(7593)) or (layer0_outputs(10607));
    layer1_outputs(1954) <= (layer0_outputs(2619)) and (layer0_outputs(10145));
    layer1_outputs(1955) <= (layer0_outputs(9828)) xor (layer0_outputs(12615));
    layer1_outputs(1956) <= (layer0_outputs(12126)) and not (layer0_outputs(6921));
    layer1_outputs(1957) <= not(layer0_outputs(8694));
    layer1_outputs(1958) <= not(layer0_outputs(4377)) or (layer0_outputs(2160));
    layer1_outputs(1959) <= (layer0_outputs(9879)) xor (layer0_outputs(7056));
    layer1_outputs(1960) <= not((layer0_outputs(11743)) or (layer0_outputs(7360)));
    layer1_outputs(1961) <= not(layer0_outputs(11603));
    layer1_outputs(1962) <= not(layer0_outputs(5253)) or (layer0_outputs(8710));
    layer1_outputs(1963) <= not(layer0_outputs(12689));
    layer1_outputs(1964) <= (layer0_outputs(7345)) and (layer0_outputs(209));
    layer1_outputs(1965) <= not(layer0_outputs(1670));
    layer1_outputs(1966) <= not(layer0_outputs(9978)) or (layer0_outputs(5741));
    layer1_outputs(1967) <= not((layer0_outputs(2083)) and (layer0_outputs(3228)));
    layer1_outputs(1968) <= not(layer0_outputs(2102));
    layer1_outputs(1969) <= not(layer0_outputs(1848));
    layer1_outputs(1970) <= not(layer0_outputs(12248));
    layer1_outputs(1971) <= layer0_outputs(12651);
    layer1_outputs(1972) <= not(layer0_outputs(3398));
    layer1_outputs(1973) <= not((layer0_outputs(3927)) xor (layer0_outputs(6372)));
    layer1_outputs(1974) <= layer0_outputs(6471);
    layer1_outputs(1975) <= not((layer0_outputs(1065)) and (layer0_outputs(3320)));
    layer1_outputs(1976) <= not(layer0_outputs(12467));
    layer1_outputs(1977) <= (layer0_outputs(1088)) and not (layer0_outputs(116));
    layer1_outputs(1978) <= not(layer0_outputs(413));
    layer1_outputs(1979) <= (layer0_outputs(6515)) and not (layer0_outputs(11447));
    layer1_outputs(1980) <= not(layer0_outputs(5811)) or (layer0_outputs(921));
    layer1_outputs(1981) <= layer0_outputs(4477);
    layer1_outputs(1982) <= (layer0_outputs(3175)) or (layer0_outputs(10930));
    layer1_outputs(1983) <= layer0_outputs(4549);
    layer1_outputs(1984) <= not(layer0_outputs(9745));
    layer1_outputs(1985) <= not(layer0_outputs(2720)) or (layer0_outputs(4743));
    layer1_outputs(1986) <= not((layer0_outputs(10426)) or (layer0_outputs(10988)));
    layer1_outputs(1987) <= layer0_outputs(5292);
    layer1_outputs(1988) <= layer0_outputs(7988);
    layer1_outputs(1989) <= not((layer0_outputs(8346)) and (layer0_outputs(2448)));
    layer1_outputs(1990) <= (layer0_outputs(277)) and not (layer0_outputs(5781));
    layer1_outputs(1991) <= (layer0_outputs(458)) xor (layer0_outputs(6081));
    layer1_outputs(1992) <= layer0_outputs(11080);
    layer1_outputs(1993) <= not((layer0_outputs(11318)) and (layer0_outputs(993)));
    layer1_outputs(1994) <= not((layer0_outputs(5182)) xor (layer0_outputs(7618)));
    layer1_outputs(1995) <= not(layer0_outputs(10233)) or (layer0_outputs(12752));
    layer1_outputs(1996) <= (layer0_outputs(11193)) and not (layer0_outputs(9306));
    layer1_outputs(1997) <= (layer0_outputs(7294)) xor (layer0_outputs(7703));
    layer1_outputs(1998) <= not(layer0_outputs(5319));
    layer1_outputs(1999) <= not((layer0_outputs(6158)) or (layer0_outputs(9196)));
    layer1_outputs(2000) <= not(layer0_outputs(12431));
    layer1_outputs(2001) <= layer0_outputs(9130);
    layer1_outputs(2002) <= not(layer0_outputs(7160));
    layer1_outputs(2003) <= (layer0_outputs(3839)) and (layer0_outputs(6600));
    layer1_outputs(2004) <= (layer0_outputs(2271)) or (layer0_outputs(8028));
    layer1_outputs(2005) <= layer0_outputs(6858);
    layer1_outputs(2006) <= not((layer0_outputs(12539)) and (layer0_outputs(4724)));
    layer1_outputs(2007) <= not(layer0_outputs(7113));
    layer1_outputs(2008) <= (layer0_outputs(6663)) xor (layer0_outputs(2441));
    layer1_outputs(2009) <= not((layer0_outputs(12270)) and (layer0_outputs(4007)));
    layer1_outputs(2010) <= not(layer0_outputs(8128)) or (layer0_outputs(9525));
    layer1_outputs(2011) <= layer0_outputs(4100);
    layer1_outputs(2012) <= (layer0_outputs(6537)) xor (layer0_outputs(9305));
    layer1_outputs(2013) <= not(layer0_outputs(3407));
    layer1_outputs(2014) <= (layer0_outputs(2368)) or (layer0_outputs(4813));
    layer1_outputs(2015) <= (layer0_outputs(6887)) or (layer0_outputs(1991));
    layer1_outputs(2016) <= not((layer0_outputs(12138)) xor (layer0_outputs(9550)));
    layer1_outputs(2017) <= not(layer0_outputs(5508));
    layer1_outputs(2018) <= not(layer0_outputs(6648)) or (layer0_outputs(10350));
    layer1_outputs(2019) <= layer0_outputs(5056);
    layer1_outputs(2020) <= not(layer0_outputs(9933));
    layer1_outputs(2021) <= not((layer0_outputs(3816)) xor (layer0_outputs(2184)));
    layer1_outputs(2022) <= not((layer0_outputs(8993)) xor (layer0_outputs(3291)));
    layer1_outputs(2023) <= layer0_outputs(11958);
    layer1_outputs(2024) <= layer0_outputs(12747);
    layer1_outputs(2025) <= (layer0_outputs(11993)) or (layer0_outputs(7063));
    layer1_outputs(2026) <= not(layer0_outputs(7094));
    layer1_outputs(2027) <= layer0_outputs(10093);
    layer1_outputs(2028) <= not((layer0_outputs(10196)) and (layer0_outputs(774)));
    layer1_outputs(2029) <= (layer0_outputs(689)) or (layer0_outputs(11876));
    layer1_outputs(2030) <= (layer0_outputs(5828)) and (layer0_outputs(5631));
    layer1_outputs(2031) <= not(layer0_outputs(188));
    layer1_outputs(2032) <= (layer0_outputs(9047)) or (layer0_outputs(3491));
    layer1_outputs(2033) <= not(layer0_outputs(3399));
    layer1_outputs(2034) <= not(layer0_outputs(11211)) or (layer0_outputs(2546));
    layer1_outputs(2035) <= not(layer0_outputs(571)) or (layer0_outputs(3682));
    layer1_outputs(2036) <= (layer0_outputs(8866)) and not (layer0_outputs(9406));
    layer1_outputs(2037) <= (layer0_outputs(3820)) and not (layer0_outputs(1708));
    layer1_outputs(2038) <= '0';
    layer1_outputs(2039) <= layer0_outputs(4850);
    layer1_outputs(2040) <= not(layer0_outputs(5872)) or (layer0_outputs(12201));
    layer1_outputs(2041) <= (layer0_outputs(5966)) and not (layer0_outputs(12094));
    layer1_outputs(2042) <= not((layer0_outputs(6388)) or (layer0_outputs(7217)));
    layer1_outputs(2043) <= (layer0_outputs(3380)) and (layer0_outputs(5368));
    layer1_outputs(2044) <= layer0_outputs(1776);
    layer1_outputs(2045) <= not(layer0_outputs(9709));
    layer1_outputs(2046) <= not(layer0_outputs(12046)) or (layer0_outputs(5553));
    layer1_outputs(2047) <= not(layer0_outputs(5703));
    layer1_outputs(2048) <= layer0_outputs(9456);
    layer1_outputs(2049) <= layer0_outputs(5771);
    layer1_outputs(2050) <= not((layer0_outputs(6945)) or (layer0_outputs(11031)));
    layer1_outputs(2051) <= not(layer0_outputs(3900)) or (layer0_outputs(9854));
    layer1_outputs(2052) <= (layer0_outputs(4826)) and not (layer0_outputs(506));
    layer1_outputs(2053) <= not(layer0_outputs(28));
    layer1_outputs(2054) <= (layer0_outputs(535)) and (layer0_outputs(5907));
    layer1_outputs(2055) <= not((layer0_outputs(2616)) or (layer0_outputs(8812)));
    layer1_outputs(2056) <= not(layer0_outputs(10034));
    layer1_outputs(2057) <= not(layer0_outputs(10968));
    layer1_outputs(2058) <= '1';
    layer1_outputs(2059) <= layer0_outputs(6706);
    layer1_outputs(2060) <= (layer0_outputs(2911)) and not (layer0_outputs(9903));
    layer1_outputs(2061) <= not(layer0_outputs(609)) or (layer0_outputs(4577));
    layer1_outputs(2062) <= (layer0_outputs(3443)) and not (layer0_outputs(10997));
    layer1_outputs(2063) <= not(layer0_outputs(11833)) or (layer0_outputs(1280));
    layer1_outputs(2064) <= (layer0_outputs(8965)) and (layer0_outputs(3275));
    layer1_outputs(2065) <= (layer0_outputs(5696)) or (layer0_outputs(8595));
    layer1_outputs(2066) <= (layer0_outputs(2891)) and not (layer0_outputs(10579));
    layer1_outputs(2067) <= layer0_outputs(11110);
    layer1_outputs(2068) <= (layer0_outputs(5303)) and not (layer0_outputs(1036));
    layer1_outputs(2069) <= '1';
    layer1_outputs(2070) <= '0';
    layer1_outputs(2071) <= not((layer0_outputs(5984)) xor (layer0_outputs(12695)));
    layer1_outputs(2072) <= not(layer0_outputs(12086));
    layer1_outputs(2073) <= not(layer0_outputs(11979));
    layer1_outputs(2074) <= (layer0_outputs(7148)) and not (layer0_outputs(5700));
    layer1_outputs(2075) <= not((layer0_outputs(10144)) or (layer0_outputs(5032)));
    layer1_outputs(2076) <= '0';
    layer1_outputs(2077) <= not((layer0_outputs(12733)) or (layer0_outputs(5885)));
    layer1_outputs(2078) <= not(layer0_outputs(573)) or (layer0_outputs(9691));
    layer1_outputs(2079) <= not(layer0_outputs(12722)) or (layer0_outputs(5471));
    layer1_outputs(2080) <= not(layer0_outputs(11561)) or (layer0_outputs(6729));
    layer1_outputs(2081) <= (layer0_outputs(8293)) xor (layer0_outputs(8730));
    layer1_outputs(2082) <= not(layer0_outputs(5772)) or (layer0_outputs(12473));
    layer1_outputs(2083) <= layer0_outputs(11323);
    layer1_outputs(2084) <= layer0_outputs(11853);
    layer1_outputs(2085) <= not(layer0_outputs(447));
    layer1_outputs(2086) <= layer0_outputs(3847);
    layer1_outputs(2087) <= not((layer0_outputs(9170)) or (layer0_outputs(5427)));
    layer1_outputs(2088) <= (layer0_outputs(9914)) and not (layer0_outputs(1131));
    layer1_outputs(2089) <= (layer0_outputs(7707)) xor (layer0_outputs(4450));
    layer1_outputs(2090) <= (layer0_outputs(553)) and (layer0_outputs(12310));
    layer1_outputs(2091) <= not((layer0_outputs(4745)) or (layer0_outputs(8534)));
    layer1_outputs(2092) <= not(layer0_outputs(2421)) or (layer0_outputs(3574));
    layer1_outputs(2093) <= not(layer0_outputs(5780)) or (layer0_outputs(378));
    layer1_outputs(2094) <= not((layer0_outputs(12717)) and (layer0_outputs(1757)));
    layer1_outputs(2095) <= not(layer0_outputs(9235)) or (layer0_outputs(6943));
    layer1_outputs(2096) <= not(layer0_outputs(8532));
    layer1_outputs(2097) <= (layer0_outputs(4661)) xor (layer0_outputs(2896));
    layer1_outputs(2098) <= not(layer0_outputs(12688)) or (layer0_outputs(1347));
    layer1_outputs(2099) <= not(layer0_outputs(2456)) or (layer0_outputs(1444));
    layer1_outputs(2100) <= not(layer0_outputs(3126));
    layer1_outputs(2101) <= layer0_outputs(1147);
    layer1_outputs(2102) <= not(layer0_outputs(2460)) or (layer0_outputs(8516));
    layer1_outputs(2103) <= layer0_outputs(5026);
    layer1_outputs(2104) <= not(layer0_outputs(5352));
    layer1_outputs(2105) <= not(layer0_outputs(3418));
    layer1_outputs(2106) <= '0';
    layer1_outputs(2107) <= layer0_outputs(6919);
    layer1_outputs(2108) <= not(layer0_outputs(492)) or (layer0_outputs(5165));
    layer1_outputs(2109) <= layer0_outputs(7925);
    layer1_outputs(2110) <= layer0_outputs(5637);
    layer1_outputs(2111) <= (layer0_outputs(12436)) and not (layer0_outputs(5455));
    layer1_outputs(2112) <= layer0_outputs(10133);
    layer1_outputs(2113) <= not(layer0_outputs(8482));
    layer1_outputs(2114) <= '1';
    layer1_outputs(2115) <= not((layer0_outputs(1273)) or (layer0_outputs(1428)));
    layer1_outputs(2116) <= not(layer0_outputs(11673));
    layer1_outputs(2117) <= not(layer0_outputs(9389));
    layer1_outputs(2118) <= layer0_outputs(4793);
    layer1_outputs(2119) <= not(layer0_outputs(10068)) or (layer0_outputs(3349));
    layer1_outputs(2120) <= (layer0_outputs(11569)) and not (layer0_outputs(12268));
    layer1_outputs(2121) <= layer0_outputs(10285);
    layer1_outputs(2122) <= (layer0_outputs(1596)) or (layer0_outputs(3936));
    layer1_outputs(2123) <= not(layer0_outputs(8783)) or (layer0_outputs(6342));
    layer1_outputs(2124) <= (layer0_outputs(5263)) and not (layer0_outputs(4743));
    layer1_outputs(2125) <= (layer0_outputs(6843)) and (layer0_outputs(3583));
    layer1_outputs(2126) <= not(layer0_outputs(720)) or (layer0_outputs(10512));
    layer1_outputs(2127) <= layer0_outputs(9487);
    layer1_outputs(2128) <= not(layer0_outputs(2016));
    layer1_outputs(2129) <= not((layer0_outputs(733)) xor (layer0_outputs(746)));
    layer1_outputs(2130) <= (layer0_outputs(12738)) and not (layer0_outputs(8841));
    layer1_outputs(2131) <= layer0_outputs(250);
    layer1_outputs(2132) <= (layer0_outputs(6265)) xor (layer0_outputs(9597));
    layer1_outputs(2133) <= layer0_outputs(39);
    layer1_outputs(2134) <= not(layer0_outputs(6866));
    layer1_outputs(2135) <= not(layer0_outputs(11516));
    layer1_outputs(2136) <= not(layer0_outputs(10964)) or (layer0_outputs(4369));
    layer1_outputs(2137) <= (layer0_outputs(6576)) and not (layer0_outputs(8557));
    layer1_outputs(2138) <= layer0_outputs(558);
    layer1_outputs(2139) <= (layer0_outputs(289)) or (layer0_outputs(2204));
    layer1_outputs(2140) <= layer0_outputs(6118);
    layer1_outputs(2141) <= layer0_outputs(1047);
    layer1_outputs(2142) <= (layer0_outputs(2289)) and (layer0_outputs(45));
    layer1_outputs(2143) <= not(layer0_outputs(454));
    layer1_outputs(2144) <= layer0_outputs(4915);
    layer1_outputs(2145) <= layer0_outputs(2692);
    layer1_outputs(2146) <= not(layer0_outputs(2064));
    layer1_outputs(2147) <= not(layer0_outputs(1212)) or (layer0_outputs(5423));
    layer1_outputs(2148) <= not((layer0_outputs(6502)) xor (layer0_outputs(5373)));
    layer1_outputs(2149) <= (layer0_outputs(4758)) and not (layer0_outputs(10008));
    layer1_outputs(2150) <= not(layer0_outputs(9959)) or (layer0_outputs(1964));
    layer1_outputs(2151) <= not(layer0_outputs(9544));
    layer1_outputs(2152) <= (layer0_outputs(1465)) or (layer0_outputs(10223));
    layer1_outputs(2153) <= (layer0_outputs(1572)) or (layer0_outputs(8790));
    layer1_outputs(2154) <= (layer0_outputs(5963)) and not (layer0_outputs(2446));
    layer1_outputs(2155) <= (layer0_outputs(5449)) and not (layer0_outputs(3723));
    layer1_outputs(2156) <= not(layer0_outputs(6238));
    layer1_outputs(2157) <= not((layer0_outputs(11348)) and (layer0_outputs(1193)));
    layer1_outputs(2158) <= not((layer0_outputs(6664)) or (layer0_outputs(3739)));
    layer1_outputs(2159) <= not((layer0_outputs(11530)) xor (layer0_outputs(5306)));
    layer1_outputs(2160) <= not(layer0_outputs(9313));
    layer1_outputs(2161) <= (layer0_outputs(3352)) and not (layer0_outputs(2230));
    layer1_outputs(2162) <= not(layer0_outputs(5240));
    layer1_outputs(2163) <= not(layer0_outputs(12241));
    layer1_outputs(2164) <= (layer0_outputs(2312)) and not (layer0_outputs(11210));
    layer1_outputs(2165) <= layer0_outputs(10995);
    layer1_outputs(2166) <= (layer0_outputs(7768)) and not (layer0_outputs(1874));
    layer1_outputs(2167) <= not(layer0_outputs(10401));
    layer1_outputs(2168) <= not(layer0_outputs(1756));
    layer1_outputs(2169) <= not(layer0_outputs(10386));
    layer1_outputs(2170) <= (layer0_outputs(3344)) and not (layer0_outputs(7179));
    layer1_outputs(2171) <= not(layer0_outputs(2190)) or (layer0_outputs(4717));
    layer1_outputs(2172) <= (layer0_outputs(6198)) xor (layer0_outputs(7154));
    layer1_outputs(2173) <= layer0_outputs(12727);
    layer1_outputs(2174) <= (layer0_outputs(12465)) or (layer0_outputs(10687));
    layer1_outputs(2175) <= layer0_outputs(1025);
    layer1_outputs(2176) <= not(layer0_outputs(1830));
    layer1_outputs(2177) <= not(layer0_outputs(8121));
    layer1_outputs(2178) <= not((layer0_outputs(3083)) xor (layer0_outputs(1140)));
    layer1_outputs(2179) <= not(layer0_outputs(10285));
    layer1_outputs(2180) <= layer0_outputs(9579);
    layer1_outputs(2181) <= layer0_outputs(43);
    layer1_outputs(2182) <= (layer0_outputs(2838)) and not (layer0_outputs(7679));
    layer1_outputs(2183) <= not((layer0_outputs(2165)) or (layer0_outputs(3180)));
    layer1_outputs(2184) <= layer0_outputs(10992);
    layer1_outputs(2185) <= not((layer0_outputs(1804)) xor (layer0_outputs(663)));
    layer1_outputs(2186) <= not(layer0_outputs(7913)) or (layer0_outputs(3199));
    layer1_outputs(2187) <= not((layer0_outputs(228)) or (layer0_outputs(1901)));
    layer1_outputs(2188) <= not(layer0_outputs(9426));
    layer1_outputs(2189) <= not(layer0_outputs(3163));
    layer1_outputs(2190) <= layer0_outputs(1236);
    layer1_outputs(2191) <= layer0_outputs(10487);
    layer1_outputs(2192) <= layer0_outputs(12562);
    layer1_outputs(2193) <= not((layer0_outputs(9501)) and (layer0_outputs(41)));
    layer1_outputs(2194) <= not(layer0_outputs(7697));
    layer1_outputs(2195) <= (layer0_outputs(4397)) and not (layer0_outputs(6493));
    layer1_outputs(2196) <= not(layer0_outputs(12006));
    layer1_outputs(2197) <= not(layer0_outputs(6268));
    layer1_outputs(2198) <= layer0_outputs(2655);
    layer1_outputs(2199) <= not(layer0_outputs(6523));
    layer1_outputs(2200) <= not((layer0_outputs(4613)) xor (layer0_outputs(7609)));
    layer1_outputs(2201) <= not(layer0_outputs(7917));
    layer1_outputs(2202) <= not(layer0_outputs(8244)) or (layer0_outputs(9895));
    layer1_outputs(2203) <= (layer0_outputs(5466)) and not (layer0_outputs(1869));
    layer1_outputs(2204) <= layer0_outputs(12110);
    layer1_outputs(2205) <= (layer0_outputs(2823)) and not (layer0_outputs(5810));
    layer1_outputs(2206) <= not(layer0_outputs(11265));
    layer1_outputs(2207) <= not((layer0_outputs(9448)) or (layer0_outputs(5152)));
    layer1_outputs(2208) <= not(layer0_outputs(12744)) or (layer0_outputs(4586));
    layer1_outputs(2209) <= layer0_outputs(11285);
    layer1_outputs(2210) <= '1';
    layer1_outputs(2211) <= (layer0_outputs(2029)) and not (layer0_outputs(6746));
    layer1_outputs(2212) <= layer0_outputs(1985);
    layer1_outputs(2213) <= not(layer0_outputs(5016)) or (layer0_outputs(4715));
    layer1_outputs(2214) <= (layer0_outputs(11413)) or (layer0_outputs(3008));
    layer1_outputs(2215) <= not((layer0_outputs(7193)) xor (layer0_outputs(4516)));
    layer1_outputs(2216) <= layer0_outputs(11239);
    layer1_outputs(2217) <= not(layer0_outputs(5043));
    layer1_outputs(2218) <= not(layer0_outputs(12205));
    layer1_outputs(2219) <= (layer0_outputs(5510)) and not (layer0_outputs(2617));
    layer1_outputs(2220) <= layer0_outputs(3978);
    layer1_outputs(2221) <= not(layer0_outputs(8896)) or (layer0_outputs(3024));
    layer1_outputs(2222) <= (layer0_outputs(3261)) xor (layer0_outputs(12690));
    layer1_outputs(2223) <= not(layer0_outputs(11149)) or (layer0_outputs(9542));
    layer1_outputs(2224) <= not((layer0_outputs(3540)) or (layer0_outputs(2240)));
    layer1_outputs(2225) <= not(layer0_outputs(8829));
    layer1_outputs(2226) <= not(layer0_outputs(12725));
    layer1_outputs(2227) <= (layer0_outputs(10472)) and not (layer0_outputs(996));
    layer1_outputs(2228) <= (layer0_outputs(5350)) and not (layer0_outputs(11359));
    layer1_outputs(2229) <= layer0_outputs(9650);
    layer1_outputs(2230) <= (layer0_outputs(12660)) and not (layer0_outputs(3170));
    layer1_outputs(2231) <= (layer0_outputs(8917)) and (layer0_outputs(3301));
    layer1_outputs(2232) <= not(layer0_outputs(9719)) or (layer0_outputs(3101));
    layer1_outputs(2233) <= not(layer0_outputs(7711)) or (layer0_outputs(11970));
    layer1_outputs(2234) <= layer0_outputs(4491);
    layer1_outputs(2235) <= not(layer0_outputs(2668)) or (layer0_outputs(10238));
    layer1_outputs(2236) <= not((layer0_outputs(12504)) and (layer0_outputs(3886)));
    layer1_outputs(2237) <= not((layer0_outputs(6601)) and (layer0_outputs(9934)));
    layer1_outputs(2238) <= (layer0_outputs(10307)) and not (layer0_outputs(3621));
    layer1_outputs(2239) <= (layer0_outputs(10526)) xor (layer0_outputs(5719));
    layer1_outputs(2240) <= not((layer0_outputs(10260)) xor (layer0_outputs(9027)));
    layer1_outputs(2241) <= layer0_outputs(6653);
    layer1_outputs(2242) <= layer0_outputs(1336);
    layer1_outputs(2243) <= (layer0_outputs(5543)) and not (layer0_outputs(10735));
    layer1_outputs(2244) <= not((layer0_outputs(5856)) and (layer0_outputs(8738)));
    layer1_outputs(2245) <= not((layer0_outputs(766)) or (layer0_outputs(1028)));
    layer1_outputs(2246) <= not(layer0_outputs(7725));
    layer1_outputs(2247) <= (layer0_outputs(9929)) and not (layer0_outputs(7694));
    layer1_outputs(2248) <= layer0_outputs(991);
    layer1_outputs(2249) <= (layer0_outputs(11060)) and (layer0_outputs(3585));
    layer1_outputs(2250) <= not(layer0_outputs(10639));
    layer1_outputs(2251) <= (layer0_outputs(4972)) and not (layer0_outputs(3517));
    layer1_outputs(2252) <= layer0_outputs(8030);
    layer1_outputs(2253) <= (layer0_outputs(8784)) and (layer0_outputs(315));
    layer1_outputs(2254) <= layer0_outputs(8295);
    layer1_outputs(2255) <= layer0_outputs(2589);
    layer1_outputs(2256) <= not(layer0_outputs(1203));
    layer1_outputs(2257) <= layer0_outputs(12767);
    layer1_outputs(2258) <= not(layer0_outputs(3434));
    layer1_outputs(2259) <= '1';
    layer1_outputs(2260) <= (layer0_outputs(10240)) and not (layer0_outputs(164));
    layer1_outputs(2261) <= not((layer0_outputs(4646)) and (layer0_outputs(11024)));
    layer1_outputs(2262) <= not(layer0_outputs(5469));
    layer1_outputs(2263) <= layer0_outputs(9846);
    layer1_outputs(2264) <= not(layer0_outputs(3151)) or (layer0_outputs(12402));
    layer1_outputs(2265) <= layer0_outputs(1867);
    layer1_outputs(2266) <= layer0_outputs(12208);
    layer1_outputs(2267) <= (layer0_outputs(854)) or (layer0_outputs(6190));
    layer1_outputs(2268) <= layer0_outputs(2950);
    layer1_outputs(2269) <= (layer0_outputs(10431)) and not (layer0_outputs(2724));
    layer1_outputs(2270) <= (layer0_outputs(8662)) and not (layer0_outputs(1676));
    layer1_outputs(2271) <= (layer0_outputs(9659)) or (layer0_outputs(6575));
    layer1_outputs(2272) <= (layer0_outputs(1864)) and not (layer0_outputs(12391));
    layer1_outputs(2273) <= (layer0_outputs(8981)) xor (layer0_outputs(3972));
    layer1_outputs(2274) <= not(layer0_outputs(5493));
    layer1_outputs(2275) <= (layer0_outputs(10755)) or (layer0_outputs(11537));
    layer1_outputs(2276) <= layer0_outputs(4482);
    layer1_outputs(2277) <= layer0_outputs(815);
    layer1_outputs(2278) <= not(layer0_outputs(11197));
    layer1_outputs(2279) <= (layer0_outputs(10562)) and not (layer0_outputs(5208));
    layer1_outputs(2280) <= (layer0_outputs(5705)) and not (layer0_outputs(1833));
    layer1_outputs(2281) <= not((layer0_outputs(12757)) and (layer0_outputs(9343)));
    layer1_outputs(2282) <= layer0_outputs(9183);
    layer1_outputs(2283) <= (layer0_outputs(2602)) and (layer0_outputs(7896));
    layer1_outputs(2284) <= not(layer0_outputs(10658)) or (layer0_outputs(2265));
    layer1_outputs(2285) <= (layer0_outputs(5537)) or (layer0_outputs(10509));
    layer1_outputs(2286) <= (layer0_outputs(65)) and not (layer0_outputs(9294));
    layer1_outputs(2287) <= (layer0_outputs(1730)) and not (layer0_outputs(11934));
    layer1_outputs(2288) <= not((layer0_outputs(11088)) or (layer0_outputs(7338)));
    layer1_outputs(2289) <= layer0_outputs(6830);
    layer1_outputs(2290) <= not((layer0_outputs(12015)) xor (layer0_outputs(5847)));
    layer1_outputs(2291) <= not((layer0_outputs(2607)) xor (layer0_outputs(11792)));
    layer1_outputs(2292) <= (layer0_outputs(4146)) xor (layer0_outputs(9125));
    layer1_outputs(2293) <= not(layer0_outputs(942));
    layer1_outputs(2294) <= not(layer0_outputs(12251));
    layer1_outputs(2295) <= (layer0_outputs(354)) and (layer0_outputs(8089));
    layer1_outputs(2296) <= not(layer0_outputs(11998));
    layer1_outputs(2297) <= (layer0_outputs(2756)) and not (layer0_outputs(3611));
    layer1_outputs(2298) <= not((layer0_outputs(11151)) xor (layer0_outputs(9768)));
    layer1_outputs(2299) <= (layer0_outputs(6558)) xor (layer0_outputs(4274));
    layer1_outputs(2300) <= (layer0_outputs(10864)) or (layer0_outputs(8473));
    layer1_outputs(2301) <= (layer0_outputs(5809)) or (layer0_outputs(8736));
    layer1_outputs(2302) <= not((layer0_outputs(3866)) and (layer0_outputs(3253)));
    layer1_outputs(2303) <= not(layer0_outputs(8294)) or (layer0_outputs(11890));
    layer1_outputs(2304) <= layer0_outputs(7631);
    layer1_outputs(2305) <= (layer0_outputs(2562)) xor (layer0_outputs(10029));
    layer1_outputs(2306) <= not(layer0_outputs(12775));
    layer1_outputs(2307) <= (layer0_outputs(7176)) and (layer0_outputs(12371));
    layer1_outputs(2308) <= not(layer0_outputs(5253)) or (layer0_outputs(7077));
    layer1_outputs(2309) <= not(layer0_outputs(7844));
    layer1_outputs(2310) <= not(layer0_outputs(11840)) or (layer0_outputs(695));
    layer1_outputs(2311) <= not(layer0_outputs(6050));
    layer1_outputs(2312) <= not((layer0_outputs(8921)) xor (layer0_outputs(8361)));
    layer1_outputs(2313) <= (layer0_outputs(9119)) and not (layer0_outputs(1989));
    layer1_outputs(2314) <= layer0_outputs(713);
    layer1_outputs(2315) <= layer0_outputs(2049);
    layer1_outputs(2316) <= not(layer0_outputs(5694));
    layer1_outputs(2317) <= (layer0_outputs(11581)) and not (layer0_outputs(4205));
    layer1_outputs(2318) <= layer0_outputs(6075);
    layer1_outputs(2319) <= (layer0_outputs(12396)) and not (layer0_outputs(3196));
    layer1_outputs(2320) <= not(layer0_outputs(8431)) or (layer0_outputs(9402));
    layer1_outputs(2321) <= not(layer0_outputs(8162));
    layer1_outputs(2322) <= not(layer0_outputs(6563)) or (layer0_outputs(1812));
    layer1_outputs(2323) <= (layer0_outputs(1064)) and not (layer0_outputs(7467));
    layer1_outputs(2324) <= (layer0_outputs(11411)) or (layer0_outputs(8878));
    layer1_outputs(2325) <= (layer0_outputs(6269)) or (layer0_outputs(4850));
    layer1_outputs(2326) <= layer0_outputs(7746);
    layer1_outputs(2327) <= not((layer0_outputs(1652)) and (layer0_outputs(4746)));
    layer1_outputs(2328) <= not(layer0_outputs(12611)) or (layer0_outputs(10605));
    layer1_outputs(2329) <= not((layer0_outputs(4829)) and (layer0_outputs(5417)));
    layer1_outputs(2330) <= not(layer0_outputs(1928));
    layer1_outputs(2331) <= layer0_outputs(3519);
    layer1_outputs(2332) <= not(layer0_outputs(9647));
    layer1_outputs(2333) <= not(layer0_outputs(12753)) or (layer0_outputs(12040));
    layer1_outputs(2334) <= not(layer0_outputs(11700));
    layer1_outputs(2335) <= layer0_outputs(11295);
    layer1_outputs(2336) <= (layer0_outputs(6248)) xor (layer0_outputs(3007));
    layer1_outputs(2337) <= (layer0_outputs(573)) or (layer0_outputs(5562));
    layer1_outputs(2338) <= not(layer0_outputs(2766));
    layer1_outputs(2339) <= not(layer0_outputs(10385));
    layer1_outputs(2340) <= not((layer0_outputs(7142)) xor (layer0_outputs(3079)));
    layer1_outputs(2341) <= not(layer0_outputs(7088));
    layer1_outputs(2342) <= not(layer0_outputs(1226));
    layer1_outputs(2343) <= (layer0_outputs(5916)) and not (layer0_outputs(1378));
    layer1_outputs(2344) <= not((layer0_outputs(6855)) or (layer0_outputs(1647)));
    layer1_outputs(2345) <= (layer0_outputs(6429)) and not (layer0_outputs(2357));
    layer1_outputs(2346) <= (layer0_outputs(8081)) and not (layer0_outputs(12409));
    layer1_outputs(2347) <= not(layer0_outputs(2634)) or (layer0_outputs(8334));
    layer1_outputs(2348) <= not((layer0_outputs(5184)) or (layer0_outputs(2394)));
    layer1_outputs(2349) <= not((layer0_outputs(4248)) or (layer0_outputs(11360)));
    layer1_outputs(2350) <= not(layer0_outputs(10662));
    layer1_outputs(2351) <= (layer0_outputs(550)) and not (layer0_outputs(12346));
    layer1_outputs(2352) <= layer0_outputs(223);
    layer1_outputs(2353) <= layer0_outputs(1599);
    layer1_outputs(2354) <= not(layer0_outputs(2110));
    layer1_outputs(2355) <= not(layer0_outputs(6009));
    layer1_outputs(2356) <= not(layer0_outputs(2405));
    layer1_outputs(2357) <= (layer0_outputs(7685)) xor (layer0_outputs(11522));
    layer1_outputs(2358) <= not((layer0_outputs(2460)) xor (layer0_outputs(7542)));
    layer1_outputs(2359) <= not(layer0_outputs(9385));
    layer1_outputs(2360) <= (layer0_outputs(4668)) xor (layer0_outputs(289));
    layer1_outputs(2361) <= not(layer0_outputs(6699));
    layer1_outputs(2362) <= not((layer0_outputs(8142)) xor (layer0_outputs(4273)));
    layer1_outputs(2363) <= not((layer0_outputs(10079)) and (layer0_outputs(6757)));
    layer1_outputs(2364) <= not(layer0_outputs(4117));
    layer1_outputs(2365) <= (layer0_outputs(5952)) or (layer0_outputs(10622));
    layer1_outputs(2366) <= '1';
    layer1_outputs(2367) <= not(layer0_outputs(5566)) or (layer0_outputs(678));
    layer1_outputs(2368) <= (layer0_outputs(3279)) or (layer0_outputs(12247));
    layer1_outputs(2369) <= layer0_outputs(9178);
    layer1_outputs(2370) <= layer0_outputs(2675);
    layer1_outputs(2371) <= not(layer0_outputs(4044));
    layer1_outputs(2372) <= not(layer0_outputs(1432)) or (layer0_outputs(1699));
    layer1_outputs(2373) <= not(layer0_outputs(7600));
    layer1_outputs(2374) <= layer0_outputs(1404);
    layer1_outputs(2375) <= not((layer0_outputs(8420)) or (layer0_outputs(10366)));
    layer1_outputs(2376) <= not(layer0_outputs(7326));
    layer1_outputs(2377) <= (layer0_outputs(5119)) or (layer0_outputs(11236));
    layer1_outputs(2378) <= not(layer0_outputs(3051));
    layer1_outputs(2379) <= (layer0_outputs(10825)) and (layer0_outputs(562));
    layer1_outputs(2380) <= not(layer0_outputs(2336));
    layer1_outputs(2381) <= not(layer0_outputs(7772)) or (layer0_outputs(9807));
    layer1_outputs(2382) <= '0';
    layer1_outputs(2383) <= layer0_outputs(4146);
    layer1_outputs(2384) <= (layer0_outputs(7314)) xor (layer0_outputs(10435));
    layer1_outputs(2385) <= (layer0_outputs(6912)) and not (layer0_outputs(3229));
    layer1_outputs(2386) <= layer0_outputs(12018);
    layer1_outputs(2387) <= (layer0_outputs(5717)) or (layer0_outputs(11064));
    layer1_outputs(2388) <= layer0_outputs(5605);
    layer1_outputs(2389) <= layer0_outputs(11143);
    layer1_outputs(2390) <= not(layer0_outputs(8682));
    layer1_outputs(2391) <= layer0_outputs(5669);
    layer1_outputs(2392) <= (layer0_outputs(9194)) or (layer0_outputs(4189));
    layer1_outputs(2393) <= layer0_outputs(5642);
    layer1_outputs(2394) <= (layer0_outputs(7627)) and (layer0_outputs(3664));
    layer1_outputs(2395) <= not(layer0_outputs(174));
    layer1_outputs(2396) <= (layer0_outputs(3226)) xor (layer0_outputs(12755));
    layer1_outputs(2397) <= layer0_outputs(11069);
    layer1_outputs(2398) <= (layer0_outputs(11826)) xor (layer0_outputs(9112));
    layer1_outputs(2399) <= (layer0_outputs(12636)) and not (layer0_outputs(8999));
    layer1_outputs(2400) <= (layer0_outputs(191)) and (layer0_outputs(9753));
    layer1_outputs(2401) <= not(layer0_outputs(12488)) or (layer0_outputs(5484));
    layer1_outputs(2402) <= (layer0_outputs(8144)) and not (layer0_outputs(280));
    layer1_outputs(2403) <= layer0_outputs(9390);
    layer1_outputs(2404) <= (layer0_outputs(10156)) and (layer0_outputs(858));
    layer1_outputs(2405) <= not((layer0_outputs(2380)) xor (layer0_outputs(926)));
    layer1_outputs(2406) <= not(layer0_outputs(7061));
    layer1_outputs(2407) <= not(layer0_outputs(3068));
    layer1_outputs(2408) <= (layer0_outputs(12474)) and not (layer0_outputs(9082));
    layer1_outputs(2409) <= (layer0_outputs(4975)) and (layer0_outputs(10087));
    layer1_outputs(2410) <= (layer0_outputs(6932)) and (layer0_outputs(6838));
    layer1_outputs(2411) <= (layer0_outputs(10775)) and not (layer0_outputs(352));
    layer1_outputs(2412) <= layer0_outputs(8773);
    layer1_outputs(2413) <= not(layer0_outputs(4119));
    layer1_outputs(2414) <= layer0_outputs(10696);
    layer1_outputs(2415) <= layer0_outputs(12630);
    layer1_outputs(2416) <= (layer0_outputs(12030)) and not (layer0_outputs(8344));
    layer1_outputs(2417) <= not(layer0_outputs(6172));
    layer1_outputs(2418) <= not((layer0_outputs(3423)) and (layer0_outputs(9798)));
    layer1_outputs(2419) <= '0';
    layer1_outputs(2420) <= not(layer0_outputs(1754)) or (layer0_outputs(10666));
    layer1_outputs(2421) <= layer0_outputs(6448);
    layer1_outputs(2422) <= not(layer0_outputs(11330)) or (layer0_outputs(2866));
    layer1_outputs(2423) <= (layer0_outputs(10209)) xor (layer0_outputs(6320));
    layer1_outputs(2424) <= not(layer0_outputs(964));
    layer1_outputs(2425) <= not(layer0_outputs(8332));
    layer1_outputs(2426) <= not((layer0_outputs(10731)) or (layer0_outputs(9359)));
    layer1_outputs(2427) <= layer0_outputs(431);
    layer1_outputs(2428) <= not(layer0_outputs(4420));
    layer1_outputs(2429) <= (layer0_outputs(8052)) and (layer0_outputs(6311));
    layer1_outputs(2430) <= layer0_outputs(6994);
    layer1_outputs(2431) <= '1';
    layer1_outputs(2432) <= (layer0_outputs(7888)) and not (layer0_outputs(5149));
    layer1_outputs(2433) <= not(layer0_outputs(7416));
    layer1_outputs(2434) <= not(layer0_outputs(4949));
    layer1_outputs(2435) <= not((layer0_outputs(11301)) and (layer0_outputs(42)));
    layer1_outputs(2436) <= layer0_outputs(8389);
    layer1_outputs(2437) <= not((layer0_outputs(1812)) xor (layer0_outputs(6716)));
    layer1_outputs(2438) <= not((layer0_outputs(4586)) and (layer0_outputs(10213)));
    layer1_outputs(2439) <= (layer0_outputs(12271)) xor (layer0_outputs(4845));
    layer1_outputs(2440) <= layer0_outputs(288);
    layer1_outputs(2441) <= layer0_outputs(4229);
    layer1_outputs(2442) <= (layer0_outputs(7831)) or (layer0_outputs(328));
    layer1_outputs(2443) <= not(layer0_outputs(3468));
    layer1_outputs(2444) <= (layer0_outputs(4667)) and not (layer0_outputs(10140));
    layer1_outputs(2445) <= (layer0_outputs(7138)) and not (layer0_outputs(8436));
    layer1_outputs(2446) <= not((layer0_outputs(10980)) and (layer0_outputs(2810)));
    layer1_outputs(2447) <= not((layer0_outputs(12417)) xor (layer0_outputs(6083)));
    layer1_outputs(2448) <= layer0_outputs(6093);
    layer1_outputs(2449) <= (layer0_outputs(701)) or (layer0_outputs(9277));
    layer1_outputs(2450) <= layer0_outputs(6533);
    layer1_outputs(2451) <= not(layer0_outputs(3052)) or (layer0_outputs(10448));
    layer1_outputs(2452) <= not(layer0_outputs(11184));
    layer1_outputs(2453) <= (layer0_outputs(2692)) and not (layer0_outputs(8697));
    layer1_outputs(2454) <= not(layer0_outputs(4816));
    layer1_outputs(2455) <= (layer0_outputs(12156)) and (layer0_outputs(9564));
    layer1_outputs(2456) <= not((layer0_outputs(12633)) xor (layer0_outputs(11323)));
    layer1_outputs(2457) <= not(layer0_outputs(4831)) or (layer0_outputs(10314));
    layer1_outputs(2458) <= layer0_outputs(1920);
    layer1_outputs(2459) <= layer0_outputs(3782);
    layer1_outputs(2460) <= (layer0_outputs(9707)) xor (layer0_outputs(6228));
    layer1_outputs(2461) <= layer0_outputs(10179);
    layer1_outputs(2462) <= layer0_outputs(6126);
    layer1_outputs(2463) <= not(layer0_outputs(10137));
    layer1_outputs(2464) <= not((layer0_outputs(4012)) xor (layer0_outputs(1614)));
    layer1_outputs(2465) <= not(layer0_outputs(8758));
    layer1_outputs(2466) <= (layer0_outputs(12068)) xor (layer0_outputs(3345));
    layer1_outputs(2467) <= '1';
    layer1_outputs(2468) <= (layer0_outputs(3432)) and (layer0_outputs(983));
    layer1_outputs(2469) <= (layer0_outputs(5797)) and not (layer0_outputs(6330));
    layer1_outputs(2470) <= (layer0_outputs(5007)) or (layer0_outputs(8321));
    layer1_outputs(2471) <= not(layer0_outputs(8154)) or (layer0_outputs(10887));
    layer1_outputs(2472) <= (layer0_outputs(988)) and not (layer0_outputs(10421));
    layer1_outputs(2473) <= layer0_outputs(5050);
    layer1_outputs(2474) <= (layer0_outputs(6554)) and (layer0_outputs(6210));
    layer1_outputs(2475) <= not(layer0_outputs(4949));
    layer1_outputs(2476) <= not(layer0_outputs(10900));
    layer1_outputs(2477) <= not(layer0_outputs(9292));
    layer1_outputs(2478) <= not(layer0_outputs(12291)) or (layer0_outputs(8071));
    layer1_outputs(2479) <= not(layer0_outputs(4003));
    layer1_outputs(2480) <= layer0_outputs(3641);
    layer1_outputs(2481) <= not(layer0_outputs(7588));
    layer1_outputs(2482) <= not(layer0_outputs(3743));
    layer1_outputs(2483) <= not((layer0_outputs(8985)) and (layer0_outputs(9491)));
    layer1_outputs(2484) <= layer0_outputs(11083);
    layer1_outputs(2485) <= not((layer0_outputs(11041)) and (layer0_outputs(2944)));
    layer1_outputs(2486) <= layer0_outputs(7851);
    layer1_outputs(2487) <= layer0_outputs(8521);
    layer1_outputs(2488) <= not((layer0_outputs(11843)) and (layer0_outputs(3887)));
    layer1_outputs(2489) <= layer0_outputs(10153);
    layer1_outputs(2490) <= layer0_outputs(11110);
    layer1_outputs(2491) <= '0';
    layer1_outputs(2492) <= (layer0_outputs(10776)) and not (layer0_outputs(888));
    layer1_outputs(2493) <= layer0_outputs(2375);
    layer1_outputs(2494) <= not((layer0_outputs(7724)) or (layer0_outputs(846)));
    layer1_outputs(2495) <= not(layer0_outputs(6172)) or (layer0_outputs(6933));
    layer1_outputs(2496) <= (layer0_outputs(379)) or (layer0_outputs(9540));
    layer1_outputs(2497) <= (layer0_outputs(1818)) and (layer0_outputs(6871));
    layer1_outputs(2498) <= (layer0_outputs(8349)) and not (layer0_outputs(1831));
    layer1_outputs(2499) <= layer0_outputs(12638);
    layer1_outputs(2500) <= not((layer0_outputs(4529)) or (layer0_outputs(7113)));
    layer1_outputs(2501) <= layer0_outputs(3525);
    layer1_outputs(2502) <= not((layer0_outputs(2373)) xor (layer0_outputs(5449)));
    layer1_outputs(2503) <= not(layer0_outputs(9659)) or (layer0_outputs(5354));
    layer1_outputs(2504) <= not(layer0_outputs(2505)) or (layer0_outputs(561));
    layer1_outputs(2505) <= not(layer0_outputs(4409)) or (layer0_outputs(8470));
    layer1_outputs(2506) <= (layer0_outputs(6588)) and not (layer0_outputs(9401));
    layer1_outputs(2507) <= (layer0_outputs(399)) and (layer0_outputs(4059));
    layer1_outputs(2508) <= (layer0_outputs(3358)) or (layer0_outputs(9086));
    layer1_outputs(2509) <= not(layer0_outputs(3115)) or (layer0_outputs(7162));
    layer1_outputs(2510) <= not(layer0_outputs(7088));
    layer1_outputs(2511) <= not(layer0_outputs(9642));
    layer1_outputs(2512) <= not((layer0_outputs(9092)) xor (layer0_outputs(6577)));
    layer1_outputs(2513) <= not((layer0_outputs(11745)) or (layer0_outputs(4290)));
    layer1_outputs(2514) <= not(layer0_outputs(6688));
    layer1_outputs(2515) <= layer0_outputs(6911);
    layer1_outputs(2516) <= layer0_outputs(6483);
    layer1_outputs(2517) <= not(layer0_outputs(1883));
    layer1_outputs(2518) <= layer0_outputs(11514);
    layer1_outputs(2519) <= not(layer0_outputs(1968));
    layer1_outputs(2520) <= '0';
    layer1_outputs(2521) <= not(layer0_outputs(8178));
    layer1_outputs(2522) <= (layer0_outputs(5684)) and (layer0_outputs(10635));
    layer1_outputs(2523) <= not((layer0_outputs(6196)) and (layer0_outputs(5307)));
    layer1_outputs(2524) <= layer0_outputs(9991);
    layer1_outputs(2525) <= not(layer0_outputs(4135));
    layer1_outputs(2526) <= not(layer0_outputs(4957));
    layer1_outputs(2527) <= (layer0_outputs(5892)) and not (layer0_outputs(4844));
    layer1_outputs(2528) <= layer0_outputs(6961);
    layer1_outputs(2529) <= (layer0_outputs(8184)) xor (layer0_outputs(11043));
    layer1_outputs(2530) <= (layer0_outputs(8378)) or (layer0_outputs(5970));
    layer1_outputs(2531) <= layer0_outputs(7809);
    layer1_outputs(2532) <= not(layer0_outputs(12627));
    layer1_outputs(2533) <= not(layer0_outputs(12435));
    layer1_outputs(2534) <= not((layer0_outputs(1809)) xor (layer0_outputs(6368)));
    layer1_outputs(2535) <= not(layer0_outputs(2284));
    layer1_outputs(2536) <= not(layer0_outputs(6589));
    layer1_outputs(2537) <= not(layer0_outputs(3720));
    layer1_outputs(2538) <= layer0_outputs(10010);
    layer1_outputs(2539) <= (layer0_outputs(10346)) and not (layer0_outputs(3745));
    layer1_outputs(2540) <= layer0_outputs(1753);
    layer1_outputs(2541) <= not((layer0_outputs(249)) and (layer0_outputs(3368)));
    layer1_outputs(2542) <= not((layer0_outputs(9823)) xor (layer0_outputs(5328)));
    layer1_outputs(2543) <= not(layer0_outputs(8692));
    layer1_outputs(2544) <= not((layer0_outputs(10145)) or (layer0_outputs(10825)));
    layer1_outputs(2545) <= not((layer0_outputs(2499)) and (layer0_outputs(11000)));
    layer1_outputs(2546) <= (layer0_outputs(11262)) and (layer0_outputs(288));
    layer1_outputs(2547) <= not((layer0_outputs(10115)) xor (layer0_outputs(12111)));
    layer1_outputs(2548) <= (layer0_outputs(11467)) and not (layer0_outputs(3799));
    layer1_outputs(2549) <= layer0_outputs(11039);
    layer1_outputs(2550) <= not(layer0_outputs(7632));
    layer1_outputs(2551) <= not(layer0_outputs(11290)) or (layer0_outputs(12306));
    layer1_outputs(2552) <= (layer0_outputs(278)) xor (layer0_outputs(3055));
    layer1_outputs(2553) <= layer0_outputs(11335);
    layer1_outputs(2554) <= not(layer0_outputs(11388)) or (layer0_outputs(8439));
    layer1_outputs(2555) <= not((layer0_outputs(11030)) or (layer0_outputs(1826)));
    layer1_outputs(2556) <= (layer0_outputs(1311)) and not (layer0_outputs(7095));
    layer1_outputs(2557) <= (layer0_outputs(842)) and not (layer0_outputs(11548));
    layer1_outputs(2558) <= not(layer0_outputs(11051)) or (layer0_outputs(11558));
    layer1_outputs(2559) <= (layer0_outputs(2913)) xor (layer0_outputs(6332));
    layer1_outputs(2560) <= layer0_outputs(4906);
    layer1_outputs(2561) <= layer0_outputs(10736);
    layer1_outputs(2562) <= not(layer0_outputs(12452)) or (layer0_outputs(5478));
    layer1_outputs(2563) <= not(layer0_outputs(1496)) or (layer0_outputs(2702));
    layer1_outputs(2564) <= layer0_outputs(4181);
    layer1_outputs(2565) <= not(layer0_outputs(11840));
    layer1_outputs(2566) <= not(layer0_outputs(11663)) or (layer0_outputs(12581));
    layer1_outputs(2567) <= not(layer0_outputs(3281));
    layer1_outputs(2568) <= layer0_outputs(10102);
    layer1_outputs(2569) <= not((layer0_outputs(6774)) xor (layer0_outputs(6393)));
    layer1_outputs(2570) <= (layer0_outputs(2402)) and not (layer0_outputs(1010));
    layer1_outputs(2571) <= not((layer0_outputs(4929)) xor (layer0_outputs(11042)));
    layer1_outputs(2572) <= layer0_outputs(3307);
    layer1_outputs(2573) <= layer0_outputs(5198);
    layer1_outputs(2574) <= not(layer0_outputs(10764));
    layer1_outputs(2575) <= not(layer0_outputs(5305)) or (layer0_outputs(11889));
    layer1_outputs(2576) <= not(layer0_outputs(8894)) or (layer0_outputs(620));
    layer1_outputs(2577) <= (layer0_outputs(9088)) or (layer0_outputs(6741));
    layer1_outputs(2578) <= not((layer0_outputs(10934)) xor (layer0_outputs(1534)));
    layer1_outputs(2579) <= not(layer0_outputs(198)) or (layer0_outputs(4636));
    layer1_outputs(2580) <= not(layer0_outputs(5946)) or (layer0_outputs(12182));
    layer1_outputs(2581) <= not(layer0_outputs(6060));
    layer1_outputs(2582) <= not(layer0_outputs(3630));
    layer1_outputs(2583) <= not((layer0_outputs(8962)) or (layer0_outputs(382)));
    layer1_outputs(2584) <= layer0_outputs(11595);
    layer1_outputs(2585) <= not((layer0_outputs(6343)) and (layer0_outputs(7171)));
    layer1_outputs(2586) <= (layer0_outputs(1580)) and (layer0_outputs(6230));
    layer1_outputs(2587) <= not(layer0_outputs(11999));
    layer1_outputs(2588) <= not(layer0_outputs(9509)) or (layer0_outputs(239));
    layer1_outputs(2589) <= layer0_outputs(434);
    layer1_outputs(2590) <= not(layer0_outputs(4266));
    layer1_outputs(2591) <= (layer0_outputs(7141)) and not (layer0_outputs(4150));
    layer1_outputs(2592) <= '0';
    layer1_outputs(2593) <= not(layer0_outputs(12702));
    layer1_outputs(2594) <= layer0_outputs(12556);
    layer1_outputs(2595) <= (layer0_outputs(5259)) or (layer0_outputs(5061));
    layer1_outputs(2596) <= (layer0_outputs(12260)) xor (layer0_outputs(9204));
    layer1_outputs(2597) <= not((layer0_outputs(1276)) and (layer0_outputs(3543)));
    layer1_outputs(2598) <= not(layer0_outputs(9104));
    layer1_outputs(2599) <= (layer0_outputs(7818)) and (layer0_outputs(12137));
    layer1_outputs(2600) <= not(layer0_outputs(200)) or (layer0_outputs(11560));
    layer1_outputs(2601) <= layer0_outputs(3758);
    layer1_outputs(2602) <= not(layer0_outputs(11347));
    layer1_outputs(2603) <= not(layer0_outputs(1417));
    layer1_outputs(2604) <= not(layer0_outputs(12544));
    layer1_outputs(2605) <= (layer0_outputs(4982)) and not (layer0_outputs(1650));
    layer1_outputs(2606) <= (layer0_outputs(9694)) and not (layer0_outputs(1798));
    layer1_outputs(2607) <= not((layer0_outputs(6985)) xor (layer0_outputs(7139)));
    layer1_outputs(2608) <= (layer0_outputs(11097)) and (layer0_outputs(5461));
    layer1_outputs(2609) <= layer0_outputs(1831);
    layer1_outputs(2610) <= (layer0_outputs(9681)) or (layer0_outputs(9982));
    layer1_outputs(2611) <= '0';
    layer1_outputs(2612) <= '0';
    layer1_outputs(2613) <= layer0_outputs(5131);
    layer1_outputs(2614) <= not(layer0_outputs(6347));
    layer1_outputs(2615) <= (layer0_outputs(12617)) xor (layer0_outputs(2126));
    layer1_outputs(2616) <= '0';
    layer1_outputs(2617) <= not((layer0_outputs(10951)) and (layer0_outputs(4339)));
    layer1_outputs(2618) <= '1';
    layer1_outputs(2619) <= (layer0_outputs(11816)) and (layer0_outputs(8266));
    layer1_outputs(2620) <= not(layer0_outputs(2267));
    layer1_outputs(2621) <= not(layer0_outputs(9475));
    layer1_outputs(2622) <= not((layer0_outputs(11911)) and (layer0_outputs(196)));
    layer1_outputs(2623) <= (layer0_outputs(9948)) xor (layer0_outputs(10621));
    layer1_outputs(2624) <= layer0_outputs(6355);
    layer1_outputs(2625) <= (layer0_outputs(3995)) and not (layer0_outputs(7643));
    layer1_outputs(2626) <= not(layer0_outputs(3351)) or (layer0_outputs(2496));
    layer1_outputs(2627) <= not((layer0_outputs(8632)) or (layer0_outputs(5850)));
    layer1_outputs(2628) <= not(layer0_outputs(5552));
    layer1_outputs(2629) <= (layer0_outputs(12267)) and (layer0_outputs(472));
    layer1_outputs(2630) <= not(layer0_outputs(3330)) or (layer0_outputs(5115));
    layer1_outputs(2631) <= layer0_outputs(5656);
    layer1_outputs(2632) <= '1';
    layer1_outputs(2633) <= layer0_outputs(12766);
    layer1_outputs(2634) <= not(layer0_outputs(2789)) or (layer0_outputs(9006));
    layer1_outputs(2635) <= not((layer0_outputs(52)) and (layer0_outputs(5854)));
    layer1_outputs(2636) <= (layer0_outputs(5817)) xor (layer0_outputs(10601));
    layer1_outputs(2637) <= not((layer0_outputs(6369)) and (layer0_outputs(907)));
    layer1_outputs(2638) <= not(layer0_outputs(4912));
    layer1_outputs(2639) <= layer0_outputs(6134);
    layer1_outputs(2640) <= not((layer0_outputs(1579)) and (layer0_outputs(7678)));
    layer1_outputs(2641) <= (layer0_outputs(9933)) and not (layer0_outputs(1840));
    layer1_outputs(2642) <= (layer0_outputs(821)) and not (layer0_outputs(3302));
    layer1_outputs(2643) <= not(layer0_outputs(7091)) or (layer0_outputs(9824));
    layer1_outputs(2644) <= layer0_outputs(6016);
    layer1_outputs(2645) <= not(layer0_outputs(2998));
    layer1_outputs(2646) <= not(layer0_outputs(5001));
    layer1_outputs(2647) <= layer0_outputs(12210);
    layer1_outputs(2648) <= layer0_outputs(4265);
    layer1_outputs(2649) <= not(layer0_outputs(1341)) or (layer0_outputs(9045));
    layer1_outputs(2650) <= not((layer0_outputs(7082)) and (layer0_outputs(657)));
    layer1_outputs(2651) <= not(layer0_outputs(11429));
    layer1_outputs(2652) <= layer0_outputs(2516);
    layer1_outputs(2653) <= layer0_outputs(6849);
    layer1_outputs(2654) <= layer0_outputs(593);
    layer1_outputs(2655) <= not(layer0_outputs(1037));
    layer1_outputs(2656) <= not(layer0_outputs(12196));
    layer1_outputs(2657) <= (layer0_outputs(10417)) xor (layer0_outputs(3159));
    layer1_outputs(2658) <= (layer0_outputs(8380)) and not (layer0_outputs(1937));
    layer1_outputs(2659) <= '1';
    layer1_outputs(2660) <= not(layer0_outputs(12256));
    layer1_outputs(2661) <= not(layer0_outputs(9798)) or (layer0_outputs(10569));
    layer1_outputs(2662) <= not(layer0_outputs(504));
    layer1_outputs(2663) <= (layer0_outputs(4967)) and not (layer0_outputs(5025));
    layer1_outputs(2664) <= layer0_outputs(3613);
    layer1_outputs(2665) <= not((layer0_outputs(6045)) xor (layer0_outputs(7263)));
    layer1_outputs(2666) <= not(layer0_outputs(8383)) or (layer0_outputs(12272));
    layer1_outputs(2667) <= (layer0_outputs(8729)) and not (layer0_outputs(11590));
    layer1_outputs(2668) <= not(layer0_outputs(10291));
    layer1_outputs(2669) <= (layer0_outputs(9345)) and not (layer0_outputs(2746));
    layer1_outputs(2670) <= not(layer0_outputs(11959));
    layer1_outputs(2671) <= not(layer0_outputs(7006));
    layer1_outputs(2672) <= not(layer0_outputs(7283));
    layer1_outputs(2673) <= not((layer0_outputs(7605)) or (layer0_outputs(8213)));
    layer1_outputs(2674) <= not(layer0_outputs(742));
    layer1_outputs(2675) <= (layer0_outputs(2318)) or (layer0_outputs(2793));
    layer1_outputs(2676) <= (layer0_outputs(10030)) or (layer0_outputs(5613));
    layer1_outputs(2677) <= not(layer0_outputs(1457)) or (layer0_outputs(10207));
    layer1_outputs(2678) <= not(layer0_outputs(471));
    layer1_outputs(2679) <= (layer0_outputs(10519)) or (layer0_outputs(1948));
    layer1_outputs(2680) <= not((layer0_outputs(7702)) and (layer0_outputs(7177)));
    layer1_outputs(2681) <= not(layer0_outputs(3297));
    layer1_outputs(2682) <= (layer0_outputs(8250)) and not (layer0_outputs(11218));
    layer1_outputs(2683) <= not(layer0_outputs(9841));
    layer1_outputs(2684) <= layer0_outputs(9864);
    layer1_outputs(2685) <= layer0_outputs(6440);
    layer1_outputs(2686) <= not(layer0_outputs(2069)) or (layer0_outputs(4336));
    layer1_outputs(2687) <= not((layer0_outputs(22)) xor (layer0_outputs(1970)));
    layer1_outputs(2688) <= (layer0_outputs(3289)) xor (layer0_outputs(36));
    layer1_outputs(2689) <= not((layer0_outputs(12259)) xor (layer0_outputs(6133)));
    layer1_outputs(2690) <= not(layer0_outputs(9608));
    layer1_outputs(2691) <= not((layer0_outputs(511)) xor (layer0_outputs(11371)));
    layer1_outputs(2692) <= not(layer0_outputs(6287));
    layer1_outputs(2693) <= not((layer0_outputs(7301)) and (layer0_outputs(11809)));
    layer1_outputs(2694) <= (layer0_outputs(10016)) or (layer0_outputs(7433));
    layer1_outputs(2695) <= (layer0_outputs(3000)) xor (layer0_outputs(3979));
    layer1_outputs(2696) <= (layer0_outputs(7736)) and not (layer0_outputs(4699));
    layer1_outputs(2697) <= not(layer0_outputs(6000));
    layer1_outputs(2698) <= (layer0_outputs(6767)) and not (layer0_outputs(6856));
    layer1_outputs(2699) <= not(layer0_outputs(4107));
    layer1_outputs(2700) <= layer0_outputs(4182);
    layer1_outputs(2701) <= (layer0_outputs(11267)) and not (layer0_outputs(6007));
    layer1_outputs(2702) <= not(layer0_outputs(4104));
    layer1_outputs(2703) <= (layer0_outputs(5791)) and (layer0_outputs(98));
    layer1_outputs(2704) <= not(layer0_outputs(11926));
    layer1_outputs(2705) <= not(layer0_outputs(7843));
    layer1_outputs(2706) <= not((layer0_outputs(1382)) xor (layer0_outputs(9324)));
    layer1_outputs(2707) <= layer0_outputs(4866);
    layer1_outputs(2708) <= (layer0_outputs(1933)) and not (layer0_outputs(12697));
    layer1_outputs(2709) <= not(layer0_outputs(10079));
    layer1_outputs(2710) <= (layer0_outputs(8274)) or (layer0_outputs(12214));
    layer1_outputs(2711) <= not(layer0_outputs(9731));
    layer1_outputs(2712) <= (layer0_outputs(11999)) and (layer0_outputs(9620));
    layer1_outputs(2713) <= not(layer0_outputs(9700));
    layer1_outputs(2714) <= layer0_outputs(6587);
    layer1_outputs(2715) <= not(layer0_outputs(6043));
    layer1_outputs(2716) <= not(layer0_outputs(7321)) or (layer0_outputs(8867));
    layer1_outputs(2717) <= (layer0_outputs(5660)) or (layer0_outputs(5255));
    layer1_outputs(2718) <= layer0_outputs(6519);
    layer1_outputs(2719) <= '1';
    layer1_outputs(2720) <= not(layer0_outputs(9568)) or (layer0_outputs(7716));
    layer1_outputs(2721) <= (layer0_outputs(306)) xor (layer0_outputs(9598));
    layer1_outputs(2722) <= not((layer0_outputs(3238)) xor (layer0_outputs(9793)));
    layer1_outputs(2723) <= layer0_outputs(9390);
    layer1_outputs(2724) <= (layer0_outputs(10739)) xor (layer0_outputs(1596));
    layer1_outputs(2725) <= not(layer0_outputs(276));
    layer1_outputs(2726) <= layer0_outputs(796);
    layer1_outputs(2727) <= not(layer0_outputs(8718));
    layer1_outputs(2728) <= not((layer0_outputs(6652)) or (layer0_outputs(4)));
    layer1_outputs(2729) <= not(layer0_outputs(12279));
    layer1_outputs(2730) <= (layer0_outputs(10852)) xor (layer0_outputs(7911));
    layer1_outputs(2731) <= not(layer0_outputs(8927));
    layer1_outputs(2732) <= not(layer0_outputs(2873));
    layer1_outputs(2733) <= (layer0_outputs(3123)) and not (layer0_outputs(8587));
    layer1_outputs(2734) <= not((layer0_outputs(12080)) xor (layer0_outputs(4188)));
    layer1_outputs(2735) <= not(layer0_outputs(5633)) or (layer0_outputs(4395));
    layer1_outputs(2736) <= (layer0_outputs(10959)) xor (layer0_outputs(2082));
    layer1_outputs(2737) <= not(layer0_outputs(495));
    layer1_outputs(2738) <= not(layer0_outputs(1871));
    layer1_outputs(2739) <= not(layer0_outputs(10244)) or (layer0_outputs(9159));
    layer1_outputs(2740) <= (layer0_outputs(89)) and not (layer0_outputs(11362));
    layer1_outputs(2741) <= (layer0_outputs(1553)) and (layer0_outputs(486));
    layer1_outputs(2742) <= layer0_outputs(11583);
    layer1_outputs(2743) <= '1';
    layer1_outputs(2744) <= not((layer0_outputs(6237)) xor (layer0_outputs(12494)));
    layer1_outputs(2745) <= not(layer0_outputs(5161));
    layer1_outputs(2746) <= layer0_outputs(2338);
    layer1_outputs(2747) <= '0';
    layer1_outputs(2748) <= (layer0_outputs(2287)) and not (layer0_outputs(2701));
    layer1_outputs(2749) <= not((layer0_outputs(2904)) xor (layer0_outputs(9251)));
    layer1_outputs(2750) <= not(layer0_outputs(5746));
    layer1_outputs(2751) <= not(layer0_outputs(4654));
    layer1_outputs(2752) <= not((layer0_outputs(9914)) or (layer0_outputs(10053)));
    layer1_outputs(2753) <= layer0_outputs(4096);
    layer1_outputs(2754) <= layer0_outputs(3053);
    layer1_outputs(2755) <= '1';
    layer1_outputs(2756) <= layer0_outputs(3395);
    layer1_outputs(2757) <= (layer0_outputs(2939)) or (layer0_outputs(12438));
    layer1_outputs(2758) <= layer0_outputs(11810);
    layer1_outputs(2759) <= (layer0_outputs(8247)) and not (layer0_outputs(4635));
    layer1_outputs(2760) <= layer0_outputs(4856);
    layer1_outputs(2761) <= layer0_outputs(3397);
    layer1_outputs(2762) <= not((layer0_outputs(10637)) or (layer0_outputs(9453)));
    layer1_outputs(2763) <= layer0_outputs(4973);
    layer1_outputs(2764) <= (layer0_outputs(9662)) xor (layer0_outputs(11654));
    layer1_outputs(2765) <= not(layer0_outputs(1546));
    layer1_outputs(2766) <= layer0_outputs(10634);
    layer1_outputs(2767) <= not(layer0_outputs(3554));
    layer1_outputs(2768) <= (layer0_outputs(5762)) or (layer0_outputs(10405));
    layer1_outputs(2769) <= (layer0_outputs(1921)) xor (layer0_outputs(3549));
    layer1_outputs(2770) <= layer0_outputs(2090);
    layer1_outputs(2771) <= not((layer0_outputs(8529)) and (layer0_outputs(11692)));
    layer1_outputs(2772) <= '1';
    layer1_outputs(2773) <= not(layer0_outputs(3789));
    layer1_outputs(2774) <= layer0_outputs(11948);
    layer1_outputs(2775) <= (layer0_outputs(8268)) or (layer0_outputs(5977));
    layer1_outputs(2776) <= not(layer0_outputs(9650));
    layer1_outputs(2777) <= not(layer0_outputs(4591));
    layer1_outputs(2778) <= not(layer0_outputs(9660));
    layer1_outputs(2779) <= (layer0_outputs(7118)) xor (layer0_outputs(3668));
    layer1_outputs(2780) <= not(layer0_outputs(5534));
    layer1_outputs(2781) <= (layer0_outputs(4336)) xor (layer0_outputs(11038));
    layer1_outputs(2782) <= not((layer0_outputs(9620)) or (layer0_outputs(2298)));
    layer1_outputs(2783) <= (layer0_outputs(10312)) or (layer0_outputs(7920));
    layer1_outputs(2784) <= '0';
    layer1_outputs(2785) <= (layer0_outputs(409)) and not (layer0_outputs(7610));
    layer1_outputs(2786) <= layer0_outputs(5524);
    layer1_outputs(2787) <= not(layer0_outputs(11800));
    layer1_outputs(2788) <= (layer0_outputs(4034)) or (layer0_outputs(4343));
    layer1_outputs(2789) <= not(layer0_outputs(687)) or (layer0_outputs(757));
    layer1_outputs(2790) <= layer0_outputs(4004);
    layer1_outputs(2791) <= not((layer0_outputs(5419)) xor (layer0_outputs(4255)));
    layer1_outputs(2792) <= layer0_outputs(2363);
    layer1_outputs(2793) <= not((layer0_outputs(10849)) and (layer0_outputs(3140)));
    layer1_outputs(2794) <= layer0_outputs(12207);
    layer1_outputs(2795) <= layer0_outputs(9679);
    layer1_outputs(2796) <= not(layer0_outputs(7001));
    layer1_outputs(2797) <= (layer0_outputs(12096)) or (layer0_outputs(9690));
    layer1_outputs(2798) <= (layer0_outputs(11592)) and (layer0_outputs(8526));
    layer1_outputs(2799) <= not((layer0_outputs(1063)) or (layer0_outputs(6718)));
    layer1_outputs(2800) <= not(layer0_outputs(2234));
    layer1_outputs(2801) <= not(layer0_outputs(9671));
    layer1_outputs(2802) <= not(layer0_outputs(7045));
    layer1_outputs(2803) <= (layer0_outputs(1229)) and (layer0_outputs(2647));
    layer1_outputs(2804) <= not((layer0_outputs(6203)) and (layer0_outputs(3139)));
    layer1_outputs(2805) <= layer0_outputs(12598);
    layer1_outputs(2806) <= not(layer0_outputs(1528)) or (layer0_outputs(2817));
    layer1_outputs(2807) <= layer0_outputs(4261);
    layer1_outputs(2808) <= (layer0_outputs(12110)) xor (layer0_outputs(7606));
    layer1_outputs(2809) <= (layer0_outputs(789)) xor (layer0_outputs(11487));
    layer1_outputs(2810) <= layer0_outputs(4737);
    layer1_outputs(2811) <= (layer0_outputs(253)) xor (layer0_outputs(6035));
    layer1_outputs(2812) <= (layer0_outputs(5818)) and not (layer0_outputs(10432));
    layer1_outputs(2813) <= not((layer0_outputs(9195)) xor (layer0_outputs(7447)));
    layer1_outputs(2814) <= layer0_outputs(10176);
    layer1_outputs(2815) <= not(layer0_outputs(2861));
    layer1_outputs(2816) <= layer0_outputs(2715);
    layer1_outputs(2817) <= not((layer0_outputs(8034)) and (layer0_outputs(5831)));
    layer1_outputs(2818) <= not(layer0_outputs(9576));
    layer1_outputs(2819) <= not((layer0_outputs(12795)) xor (layer0_outputs(9641)));
    layer1_outputs(2820) <= not((layer0_outputs(11683)) or (layer0_outputs(2910)));
    layer1_outputs(2821) <= not(layer0_outputs(7296)) or (layer0_outputs(6293));
    layer1_outputs(2822) <= (layer0_outputs(12320)) and (layer0_outputs(3479));
    layer1_outputs(2823) <= not(layer0_outputs(2052));
    layer1_outputs(2824) <= layer0_outputs(3050);
    layer1_outputs(2825) <= (layer0_outputs(10938)) and (layer0_outputs(8116));
    layer1_outputs(2826) <= not(layer0_outputs(1717));
    layer1_outputs(2827) <= '1';
    layer1_outputs(2828) <= (layer0_outputs(12478)) and not (layer0_outputs(6636));
    layer1_outputs(2829) <= layer0_outputs(2829);
    layer1_outputs(2830) <= not(layer0_outputs(9856)) or (layer0_outputs(3471));
    layer1_outputs(2831) <= not(layer0_outputs(6108));
    layer1_outputs(2832) <= not(layer0_outputs(4946));
    layer1_outputs(2833) <= not(layer0_outputs(8735));
    layer1_outputs(2834) <= not((layer0_outputs(8869)) xor (layer0_outputs(2368)));
    layer1_outputs(2835) <= layer0_outputs(8843);
    layer1_outputs(2836) <= not((layer0_outputs(8846)) and (layer0_outputs(7164)));
    layer1_outputs(2837) <= not(layer0_outputs(2625));
    layer1_outputs(2838) <= not(layer0_outputs(12186));
    layer1_outputs(2839) <= not(layer0_outputs(7093)) or (layer0_outputs(2730));
    layer1_outputs(2840) <= not(layer0_outputs(12378));
    layer1_outputs(2841) <= (layer0_outputs(8234)) xor (layer0_outputs(4237));
    layer1_outputs(2842) <= layer0_outputs(11634);
    layer1_outputs(2843) <= not((layer0_outputs(4338)) xor (layer0_outputs(1253)));
    layer1_outputs(2844) <= (layer0_outputs(12339)) and not (layer0_outputs(3084));
    layer1_outputs(2845) <= not(layer0_outputs(7260));
    layer1_outputs(2846) <= not(layer0_outputs(2650));
    layer1_outputs(2847) <= (layer0_outputs(8908)) and (layer0_outputs(3989));
    layer1_outputs(2848) <= layer0_outputs(8683);
    layer1_outputs(2849) <= (layer0_outputs(4061)) and not (layer0_outputs(1910));
    layer1_outputs(2850) <= (layer0_outputs(5744)) or (layer0_outputs(7690));
    layer1_outputs(2851) <= not((layer0_outputs(6780)) or (layer0_outputs(5773)));
    layer1_outputs(2852) <= not(layer0_outputs(6656)) or (layer0_outputs(326));
    layer1_outputs(2853) <= not(layer0_outputs(12559));
    layer1_outputs(2854) <= (layer0_outputs(6317)) and not (layer0_outputs(10788));
    layer1_outputs(2855) <= layer0_outputs(348);
    layer1_outputs(2856) <= not((layer0_outputs(11657)) and (layer0_outputs(530)));
    layer1_outputs(2857) <= layer0_outputs(12571);
    layer1_outputs(2858) <= not(layer0_outputs(8944));
    layer1_outputs(2859) <= layer0_outputs(11870);
    layer1_outputs(2860) <= (layer0_outputs(2073)) and not (layer0_outputs(11905));
    layer1_outputs(2861) <= not(layer0_outputs(1161));
    layer1_outputs(2862) <= not(layer0_outputs(10100));
    layer1_outputs(2863) <= (layer0_outputs(87)) xor (layer0_outputs(5433));
    layer1_outputs(2864) <= layer0_outputs(3633);
    layer1_outputs(2865) <= not(layer0_outputs(8666)) or (layer0_outputs(12134));
    layer1_outputs(2866) <= layer0_outputs(11038);
    layer1_outputs(2867) <= not(layer0_outputs(9811));
    layer1_outputs(2868) <= not(layer0_outputs(9364)) or (layer0_outputs(1733));
    layer1_outputs(2869) <= not(layer0_outputs(3039));
    layer1_outputs(2870) <= not(layer0_outputs(10888));
    layer1_outputs(2871) <= layer0_outputs(2727);
    layer1_outputs(2872) <= not(layer0_outputs(4268)) or (layer0_outputs(1472));
    layer1_outputs(2873) <= not(layer0_outputs(6695)) or (layer0_outputs(2550));
    layer1_outputs(2874) <= '1';
    layer1_outputs(2875) <= (layer0_outputs(4496)) xor (layer0_outputs(5670));
    layer1_outputs(2876) <= (layer0_outputs(7410)) and not (layer0_outputs(2963));
    layer1_outputs(2877) <= not(layer0_outputs(9332));
    layer1_outputs(2878) <= not((layer0_outputs(5133)) or (layer0_outputs(4430)));
    layer1_outputs(2879) <= (layer0_outputs(7515)) and (layer0_outputs(7718));
    layer1_outputs(2880) <= layer0_outputs(9532);
    layer1_outputs(2881) <= (layer0_outputs(529)) or (layer0_outputs(249));
    layer1_outputs(2882) <= not(layer0_outputs(11654));
    layer1_outputs(2883) <= (layer0_outputs(1963)) and not (layer0_outputs(235));
    layer1_outputs(2884) <= (layer0_outputs(11721)) or (layer0_outputs(9955));
    layer1_outputs(2885) <= (layer0_outputs(4583)) xor (layer0_outputs(4070));
    layer1_outputs(2886) <= not((layer0_outputs(4572)) and (layer0_outputs(7531)));
    layer1_outputs(2887) <= layer0_outputs(323);
    layer1_outputs(2888) <= not((layer0_outputs(3242)) or (layer0_outputs(10912)));
    layer1_outputs(2889) <= not(layer0_outputs(4416)) or (layer0_outputs(1535));
    layer1_outputs(2890) <= '1';
    layer1_outputs(2891) <= not((layer0_outputs(515)) or (layer0_outputs(9565)));
    layer1_outputs(2892) <= layer0_outputs(3895);
    layer1_outputs(2893) <= (layer0_outputs(12659)) and not (layer0_outputs(651));
    layer1_outputs(2894) <= not(layer0_outputs(6104));
    layer1_outputs(2895) <= layer0_outputs(5896);
    layer1_outputs(2896) <= (layer0_outputs(415)) or (layer0_outputs(5656));
    layer1_outputs(2897) <= (layer0_outputs(11876)) and not (layer0_outputs(11910));
    layer1_outputs(2898) <= not(layer0_outputs(8450));
    layer1_outputs(2899) <= not(layer0_outputs(4562)) or (layer0_outputs(5653));
    layer1_outputs(2900) <= (layer0_outputs(9723)) and not (layer0_outputs(6614));
    layer1_outputs(2901) <= not((layer0_outputs(6738)) xor (layer0_outputs(8814)));
    layer1_outputs(2902) <= layer0_outputs(9963);
    layer1_outputs(2903) <= not((layer0_outputs(2419)) and (layer0_outputs(4540)));
    layer1_outputs(2904) <= (layer0_outputs(5117)) and not (layer0_outputs(8618));
    layer1_outputs(2905) <= not(layer0_outputs(3812)) or (layer0_outputs(7962));
    layer1_outputs(2906) <= layer0_outputs(11356);
    layer1_outputs(2907) <= not((layer0_outputs(3284)) or (layer0_outputs(12794)));
    layer1_outputs(2908) <= not(layer0_outputs(6645)) or (layer0_outputs(1061));
    layer1_outputs(2909) <= (layer0_outputs(152)) and (layer0_outputs(5998));
    layer1_outputs(2910) <= not(layer0_outputs(8474));
    layer1_outputs(2911) <= (layer0_outputs(12290)) and (layer0_outputs(5766));
    layer1_outputs(2912) <= layer0_outputs(5731);
    layer1_outputs(2913) <= (layer0_outputs(6950)) or (layer0_outputs(11525));
    layer1_outputs(2914) <= not(layer0_outputs(859)) or (layer0_outputs(12718));
    layer1_outputs(2915) <= layer0_outputs(6544);
    layer1_outputs(2916) <= not(layer0_outputs(822));
    layer1_outputs(2917) <= not(layer0_outputs(520)) or (layer0_outputs(2560));
    layer1_outputs(2918) <= not(layer0_outputs(1));
    layer1_outputs(2919) <= not((layer0_outputs(830)) and (layer0_outputs(1581)));
    layer1_outputs(2920) <= (layer0_outputs(8977)) or (layer0_outputs(1232));
    layer1_outputs(2921) <= not(layer0_outputs(7803));
    layer1_outputs(2922) <= (layer0_outputs(6098)) or (layer0_outputs(309));
    layer1_outputs(2923) <= not(layer0_outputs(2395)) or (layer0_outputs(11414));
    layer1_outputs(2924) <= not(layer0_outputs(9836));
    layer1_outputs(2925) <= not((layer0_outputs(11465)) or (layer0_outputs(12650)));
    layer1_outputs(2926) <= (layer0_outputs(4728)) or (layer0_outputs(5205));
    layer1_outputs(2927) <= not(layer0_outputs(1011));
    layer1_outputs(2928) <= (layer0_outputs(10711)) and (layer0_outputs(3779));
    layer1_outputs(2929) <= not(layer0_outputs(12149));
    layer1_outputs(2930) <= '0';
    layer1_outputs(2931) <= (layer0_outputs(3324)) and not (layer0_outputs(1701));
    layer1_outputs(2932) <= (layer0_outputs(9047)) and not (layer0_outputs(2250));
    layer1_outputs(2933) <= not(layer0_outputs(9383)) or (layer0_outputs(8532));
    layer1_outputs(2934) <= not((layer0_outputs(6270)) xor (layer0_outputs(1938)));
    layer1_outputs(2935) <= '0';
    layer1_outputs(2936) <= not((layer0_outputs(7232)) xor (layer0_outputs(11553)));
    layer1_outputs(2937) <= layer0_outputs(9181);
    layer1_outputs(2938) <= not(layer0_outputs(11732));
    layer1_outputs(2939) <= not(layer0_outputs(1770));
    layer1_outputs(2940) <= (layer0_outputs(11291)) and (layer0_outputs(9500));
    layer1_outputs(2941) <= not(layer0_outputs(5008));
    layer1_outputs(2942) <= layer0_outputs(11805);
    layer1_outputs(2943) <= not((layer0_outputs(9116)) xor (layer0_outputs(9780)));
    layer1_outputs(2944) <= (layer0_outputs(2693)) and not (layer0_outputs(11443));
    layer1_outputs(2945) <= not(layer0_outputs(1517)) or (layer0_outputs(11624));
    layer1_outputs(2946) <= not(layer0_outputs(508)) or (layer0_outputs(6197));
    layer1_outputs(2947) <= not(layer0_outputs(1986));
    layer1_outputs(2948) <= layer0_outputs(12154);
    layer1_outputs(2949) <= not(layer0_outputs(12150)) or (layer0_outputs(1454));
    layer1_outputs(2950) <= layer0_outputs(12579);
    layer1_outputs(2951) <= not(layer0_outputs(5229));
    layer1_outputs(2952) <= not(layer0_outputs(9305)) or (layer0_outputs(4955));
    layer1_outputs(2953) <= (layer0_outputs(4241)) and not (layer0_outputs(5120));
    layer1_outputs(2954) <= (layer0_outputs(7790)) xor (layer0_outputs(4702));
    layer1_outputs(2955) <= layer0_outputs(4537);
    layer1_outputs(2956) <= layer0_outputs(9900);
    layer1_outputs(2957) <= not(layer0_outputs(5558));
    layer1_outputs(2958) <= (layer0_outputs(1413)) and (layer0_outputs(5964));
    layer1_outputs(2959) <= (layer0_outputs(10677)) and not (layer0_outputs(3322));
    layer1_outputs(2960) <= not(layer0_outputs(11217));
    layer1_outputs(2961) <= layer0_outputs(11295);
    layer1_outputs(2962) <= not((layer0_outputs(8510)) and (layer0_outputs(12529)));
    layer1_outputs(2963) <= not(layer0_outputs(2037));
    layer1_outputs(2964) <= not(layer0_outputs(4472));
    layer1_outputs(2965) <= layer0_outputs(9864);
    layer1_outputs(2966) <= not((layer0_outputs(8909)) or (layer0_outputs(1898)));
    layer1_outputs(2967) <= not(layer0_outputs(7378));
    layer1_outputs(2968) <= not((layer0_outputs(11046)) and (layer0_outputs(2303)));
    layer1_outputs(2969) <= (layer0_outputs(12294)) and not (layer0_outputs(1805));
    layer1_outputs(2970) <= (layer0_outputs(706)) or (layer0_outputs(66));
    layer1_outputs(2971) <= (layer0_outputs(1931)) and not (layer0_outputs(880));
    layer1_outputs(2972) <= not(layer0_outputs(3826)) or (layer0_outputs(7664));
    layer1_outputs(2973) <= (layer0_outputs(2412)) and (layer0_outputs(241));
    layer1_outputs(2974) <= layer0_outputs(3941);
    layer1_outputs(2975) <= layer0_outputs(6202);
    layer1_outputs(2976) <= not(layer0_outputs(5872)) or (layer0_outputs(7407));
    layer1_outputs(2977) <= (layer0_outputs(6984)) and not (layer0_outputs(5579));
    layer1_outputs(2978) <= '0';
    layer1_outputs(2979) <= not(layer0_outputs(5327));
    layer1_outputs(2980) <= layer0_outputs(10130);
    layer1_outputs(2981) <= layer0_outputs(1229);
    layer1_outputs(2982) <= (layer0_outputs(35)) and (layer0_outputs(1892));
    layer1_outputs(2983) <= not(layer0_outputs(2057));
    layer1_outputs(2984) <= (layer0_outputs(4864)) and not (layer0_outputs(9380));
    layer1_outputs(2985) <= not((layer0_outputs(2323)) or (layer0_outputs(1188)));
    layer1_outputs(2986) <= not(layer0_outputs(3153)) or (layer0_outputs(12359));
    layer1_outputs(2987) <= (layer0_outputs(7191)) xor (layer0_outputs(7799));
    layer1_outputs(2988) <= (layer0_outputs(11801)) and not (layer0_outputs(90));
    layer1_outputs(2989) <= layer0_outputs(456);
    layer1_outputs(2990) <= not(layer0_outputs(9103)) or (layer0_outputs(6678));
    layer1_outputs(2991) <= not(layer0_outputs(2042)) or (layer0_outputs(488));
    layer1_outputs(2992) <= layer0_outputs(1104);
    layer1_outputs(2993) <= (layer0_outputs(9148)) and (layer0_outputs(9515));
    layer1_outputs(2994) <= not((layer0_outputs(8343)) xor (layer0_outputs(419)));
    layer1_outputs(2995) <= not((layer0_outputs(8925)) or (layer0_outputs(11502)));
    layer1_outputs(2996) <= not((layer0_outputs(4217)) and (layer0_outputs(7421)));
    layer1_outputs(2997) <= layer0_outputs(9229);
    layer1_outputs(2998) <= not(layer0_outputs(12400));
    layer1_outputs(2999) <= not((layer0_outputs(11570)) xor (layer0_outputs(6744)));
    layer1_outputs(3000) <= not(layer0_outputs(2884));
    layer1_outputs(3001) <= layer0_outputs(2792);
    layer1_outputs(3002) <= layer0_outputs(6709);
    layer1_outputs(3003) <= not((layer0_outputs(5933)) xor (layer0_outputs(11850)));
    layer1_outputs(3004) <= not(layer0_outputs(5564));
    layer1_outputs(3005) <= (layer0_outputs(7217)) and not (layer0_outputs(10927));
    layer1_outputs(3006) <= not(layer0_outputs(11159));
    layer1_outputs(3007) <= not(layer0_outputs(12324)) or (layer0_outputs(3576));
    layer1_outputs(3008) <= (layer0_outputs(3597)) and not (layer0_outputs(11498));
    layer1_outputs(3009) <= layer0_outputs(11250);
    layer1_outputs(3010) <= not((layer0_outputs(3010)) or (layer0_outputs(7211)));
    layer1_outputs(3011) <= '0';
    layer1_outputs(3012) <= (layer0_outputs(12169)) and (layer0_outputs(3656));
    layer1_outputs(3013) <= (layer0_outputs(6156)) and not (layer0_outputs(6463));
    layer1_outputs(3014) <= not(layer0_outputs(3017)) or (layer0_outputs(10013));
    layer1_outputs(3015) <= (layer0_outputs(11094)) and not (layer0_outputs(3784));
    layer1_outputs(3016) <= (layer0_outputs(8844)) and not (layer0_outputs(12479));
    layer1_outputs(3017) <= not((layer0_outputs(935)) or (layer0_outputs(7785)));
    layer1_outputs(3018) <= layer0_outputs(11372);
    layer1_outputs(3019) <= not(layer0_outputs(9050)) or (layer0_outputs(8385));
    layer1_outputs(3020) <= (layer0_outputs(1209)) and not (layer0_outputs(1511));
    layer1_outputs(3021) <= not(layer0_outputs(3379));
    layer1_outputs(3022) <= not(layer0_outputs(10576));
    layer1_outputs(3023) <= not(layer0_outputs(325));
    layer1_outputs(3024) <= not(layer0_outputs(7086)) or (layer0_outputs(11463));
    layer1_outputs(3025) <= (layer0_outputs(10294)) and not (layer0_outputs(2484));
    layer1_outputs(3026) <= (layer0_outputs(8865)) or (layer0_outputs(8421));
    layer1_outputs(3027) <= (layer0_outputs(4692)) and (layer0_outputs(7300));
    layer1_outputs(3028) <= (layer0_outputs(5572)) and (layer0_outputs(2427));
    layer1_outputs(3029) <= (layer0_outputs(5963)) and not (layer0_outputs(12754));
    layer1_outputs(3030) <= (layer0_outputs(12132)) xor (layer0_outputs(2713));
    layer1_outputs(3031) <= not((layer0_outputs(6725)) and (layer0_outputs(6740)));
    layer1_outputs(3032) <= not(layer0_outputs(3494)) or (layer0_outputs(5568));
    layer1_outputs(3033) <= not((layer0_outputs(1961)) or (layer0_outputs(9566)));
    layer1_outputs(3034) <= layer0_outputs(5161);
    layer1_outputs(3035) <= not((layer0_outputs(2720)) xor (layer0_outputs(316)));
    layer1_outputs(3036) <= layer0_outputs(8397);
    layer1_outputs(3037) <= not((layer0_outputs(7183)) xor (layer0_outputs(11519)));
    layer1_outputs(3038) <= not(layer0_outputs(9788));
    layer1_outputs(3039) <= (layer0_outputs(4535)) or (layer0_outputs(3956));
    layer1_outputs(3040) <= not(layer0_outputs(4352));
    layer1_outputs(3041) <= not((layer0_outputs(2164)) or (layer0_outputs(1947)));
    layer1_outputs(3042) <= (layer0_outputs(6403)) and not (layer0_outputs(10577));
    layer1_outputs(3043) <= not((layer0_outputs(4673)) xor (layer0_outputs(530)));
    layer1_outputs(3044) <= not(layer0_outputs(10434));
    layer1_outputs(3045) <= (layer0_outputs(4718)) and (layer0_outputs(8904));
    layer1_outputs(3046) <= not((layer0_outputs(2915)) or (layer0_outputs(8149)));
    layer1_outputs(3047) <= (layer0_outputs(10085)) and not (layer0_outputs(613));
    layer1_outputs(3048) <= not(layer0_outputs(7261));
    layer1_outputs(3049) <= layer0_outputs(9146);
    layer1_outputs(3050) <= layer0_outputs(7034);
    layer1_outputs(3051) <= '0';
    layer1_outputs(3052) <= (layer0_outputs(5094)) and not (layer0_outputs(1307));
    layer1_outputs(3053) <= layer0_outputs(2283);
    layer1_outputs(3054) <= not((layer0_outputs(11599)) or (layer0_outputs(5776)));
    layer1_outputs(3055) <= not(layer0_outputs(5902));
    layer1_outputs(3056) <= not(layer0_outputs(5036));
    layer1_outputs(3057) <= layer0_outputs(403);
    layer1_outputs(3058) <= (layer0_outputs(10909)) xor (layer0_outputs(11961));
    layer1_outputs(3059) <= not((layer0_outputs(6249)) xor (layer0_outputs(5596)));
    layer1_outputs(3060) <= not(layer0_outputs(1434)) or (layer0_outputs(5067));
    layer1_outputs(3061) <= not((layer0_outputs(8445)) or (layer0_outputs(4341)));
    layer1_outputs(3062) <= layer0_outputs(4605);
    layer1_outputs(3063) <= '1';
    layer1_outputs(3064) <= not((layer0_outputs(9316)) and (layer0_outputs(6559)));
    layer1_outputs(3065) <= layer0_outputs(8889);
    layer1_outputs(3066) <= not(layer0_outputs(1275));
    layer1_outputs(3067) <= layer0_outputs(722);
    layer1_outputs(3068) <= '1';
    layer1_outputs(3069) <= (layer0_outputs(6305)) xor (layer0_outputs(4283));
    layer1_outputs(3070) <= not(layer0_outputs(10016));
    layer1_outputs(3071) <= (layer0_outputs(1903)) and (layer0_outputs(3772));
    layer1_outputs(3072) <= not((layer0_outputs(12268)) or (layer0_outputs(11632)));
    layer1_outputs(3073) <= not(layer0_outputs(6958));
    layer1_outputs(3074) <= (layer0_outputs(11442)) xor (layer0_outputs(572));
    layer1_outputs(3075) <= '1';
    layer1_outputs(3076) <= not((layer0_outputs(8076)) or (layer0_outputs(2306)));
    layer1_outputs(3077) <= layer0_outputs(12295);
    layer1_outputs(3078) <= not((layer0_outputs(8847)) and (layer0_outputs(11969)));
    layer1_outputs(3079) <= not((layer0_outputs(3015)) xor (layer0_outputs(10446)));
    layer1_outputs(3080) <= not(layer0_outputs(4651)) or (layer0_outputs(7384));
    layer1_outputs(3081) <= not((layer0_outputs(1919)) and (layer0_outputs(8177)));
    layer1_outputs(3082) <= not(layer0_outputs(4337));
    layer1_outputs(3083) <= not(layer0_outputs(5193));
    layer1_outputs(3084) <= not(layer0_outputs(5772));
    layer1_outputs(3085) <= (layer0_outputs(397)) and not (layer0_outputs(10972));
    layer1_outputs(3086) <= not(layer0_outputs(7503)) or (layer0_outputs(12748));
    layer1_outputs(3087) <= not(layer0_outputs(11942));
    layer1_outputs(3088) <= (layer0_outputs(6893)) and not (layer0_outputs(6878));
    layer1_outputs(3089) <= (layer0_outputs(10955)) and not (layer0_outputs(6185));
    layer1_outputs(3090) <= layer0_outputs(11100);
    layer1_outputs(3091) <= (layer0_outputs(10069)) or (layer0_outputs(9587));
    layer1_outputs(3092) <= not(layer0_outputs(9560)) or (layer0_outputs(6615));
    layer1_outputs(3093) <= layer0_outputs(1152);
    layer1_outputs(3094) <= not(layer0_outputs(12215));
    layer1_outputs(3095) <= (layer0_outputs(8523)) and (layer0_outputs(10474));
    layer1_outputs(3096) <= not(layer0_outputs(9212));
    layer1_outputs(3097) <= (layer0_outputs(592)) and not (layer0_outputs(7710));
    layer1_outputs(3098) <= (layer0_outputs(444)) and (layer0_outputs(2434));
    layer1_outputs(3099) <= not(layer0_outputs(11308)) or (layer0_outputs(10919));
    layer1_outputs(3100) <= not(layer0_outputs(6934)) or (layer0_outputs(373));
    layer1_outputs(3101) <= not(layer0_outputs(8381)) or (layer0_outputs(6659));
    layer1_outputs(3102) <= not((layer0_outputs(12604)) and (layer0_outputs(8080)));
    layer1_outputs(3103) <= not((layer0_outputs(6772)) xor (layer0_outputs(5077)));
    layer1_outputs(3104) <= '1';
    layer1_outputs(3105) <= not(layer0_outputs(11794)) or (layer0_outputs(3911));
    layer1_outputs(3106) <= not((layer0_outputs(4472)) xor (layer0_outputs(4618)));
    layer1_outputs(3107) <= (layer0_outputs(12181)) and (layer0_outputs(4547));
    layer1_outputs(3108) <= not(layer0_outputs(6273));
    layer1_outputs(3109) <= '0';
    layer1_outputs(3110) <= not(layer0_outputs(6578));
    layer1_outputs(3111) <= not((layer0_outputs(7653)) or (layer0_outputs(1643)));
    layer1_outputs(3112) <= not(layer0_outputs(7223));
    layer1_outputs(3113) <= (layer0_outputs(2197)) or (layer0_outputs(7722));
    layer1_outputs(3114) <= (layer0_outputs(6480)) and (layer0_outputs(2538));
    layer1_outputs(3115) <= layer0_outputs(7136);
    layer1_outputs(3116) <= not((layer0_outputs(4669)) or (layer0_outputs(5051)));
    layer1_outputs(3117) <= not(layer0_outputs(9300));
    layer1_outputs(3118) <= (layer0_outputs(6578)) xor (layer0_outputs(2785));
    layer1_outputs(3119) <= not(layer0_outputs(11893));
    layer1_outputs(3120) <= not(layer0_outputs(11056)) or (layer0_outputs(3438));
    layer1_outputs(3121) <= '0';
    layer1_outputs(3122) <= layer0_outputs(5891);
    layer1_outputs(3123) <= layer0_outputs(3532);
    layer1_outputs(3124) <= not(layer0_outputs(4868)) or (layer0_outputs(10134));
    layer1_outputs(3125) <= layer0_outputs(12059);
    layer1_outputs(3126) <= (layer0_outputs(1975)) and (layer0_outputs(8637));
    layer1_outputs(3127) <= (layer0_outputs(3185)) xor (layer0_outputs(1470));
    layer1_outputs(3128) <= (layer0_outputs(10812)) and (layer0_outputs(6612));
    layer1_outputs(3129) <= layer0_outputs(8613);
    layer1_outputs(3130) <= not((layer0_outputs(7136)) or (layer0_outputs(5377)));
    layer1_outputs(3131) <= not(layer0_outputs(2841));
    layer1_outputs(3132) <= '1';
    layer1_outputs(3133) <= not((layer0_outputs(12140)) or (layer0_outputs(1484)));
    layer1_outputs(3134) <= not((layer0_outputs(5953)) and (layer0_outputs(67)));
    layer1_outputs(3135) <= layer0_outputs(10971);
    layer1_outputs(3136) <= not(layer0_outputs(11785));
    layer1_outputs(3137) <= (layer0_outputs(7106)) or (layer0_outputs(7960));
    layer1_outputs(3138) <= not(layer0_outputs(4232)) or (layer0_outputs(12549));
    layer1_outputs(3139) <= not((layer0_outputs(6293)) or (layer0_outputs(7882)));
    layer1_outputs(3140) <= not((layer0_outputs(2293)) or (layer0_outputs(1154)));
    layer1_outputs(3141) <= layer0_outputs(1299);
    layer1_outputs(3142) <= (layer0_outputs(10998)) and not (layer0_outputs(12076));
    layer1_outputs(3143) <= not((layer0_outputs(2795)) or (layer0_outputs(4814)));
    layer1_outputs(3144) <= (layer0_outputs(2850)) and not (layer0_outputs(7636));
    layer1_outputs(3145) <= (layer0_outputs(478)) xor (layer0_outputs(12348));
    layer1_outputs(3146) <= not((layer0_outputs(11741)) xor (layer0_outputs(7269)));
    layer1_outputs(3147) <= '1';
    layer1_outputs(3148) <= (layer0_outputs(10362)) and not (layer0_outputs(5748));
    layer1_outputs(3149) <= not(layer0_outputs(222));
    layer1_outputs(3150) <= not(layer0_outputs(325));
    layer1_outputs(3151) <= (layer0_outputs(2990)) and not (layer0_outputs(9480));
    layer1_outputs(3152) <= not(layer0_outputs(1384));
    layer1_outputs(3153) <= not(layer0_outputs(3874));
    layer1_outputs(3154) <= not(layer0_outputs(9979));
    layer1_outputs(3155) <= layer0_outputs(10217);
    layer1_outputs(3156) <= layer0_outputs(12100);
    layer1_outputs(3157) <= (layer0_outputs(12061)) or (layer0_outputs(2119));
    layer1_outputs(3158) <= not(layer0_outputs(9030));
    layer1_outputs(3159) <= (layer0_outputs(12038)) xor (layer0_outputs(10853));
    layer1_outputs(3160) <= (layer0_outputs(5673)) and (layer0_outputs(8141));
    layer1_outputs(3161) <= not(layer0_outputs(8495)) or (layer0_outputs(4744));
    layer1_outputs(3162) <= layer0_outputs(10731);
    layer1_outputs(3163) <= '0';
    layer1_outputs(3164) <= (layer0_outputs(4588)) xor (layer0_outputs(1854));
    layer1_outputs(3165) <= (layer0_outputs(9530)) and (layer0_outputs(9124));
    layer1_outputs(3166) <= not(layer0_outputs(3869));
    layer1_outputs(3167) <= layer0_outputs(5761);
    layer1_outputs(3168) <= not((layer0_outputs(2740)) xor (layer0_outputs(7028)));
    layer1_outputs(3169) <= (layer0_outputs(5813)) and not (layer0_outputs(194));
    layer1_outputs(3170) <= layer0_outputs(7344);
    layer1_outputs(3171) <= (layer0_outputs(1507)) xor (layer0_outputs(9238));
    layer1_outputs(3172) <= not((layer0_outputs(7376)) xor (layer0_outputs(5636)));
    layer1_outputs(3173) <= (layer0_outputs(10596)) and not (layer0_outputs(6148));
    layer1_outputs(3174) <= not(layer0_outputs(3333));
    layer1_outputs(3175) <= (layer0_outputs(4507)) and (layer0_outputs(443));
    layer1_outputs(3176) <= not(layer0_outputs(11185)) or (layer0_outputs(7060));
    layer1_outputs(3177) <= not((layer0_outputs(12476)) xor (layer0_outputs(3298)));
    layer1_outputs(3178) <= not(layer0_outputs(4456));
    layer1_outputs(3179) <= layer0_outputs(1649);
    layer1_outputs(3180) <= not((layer0_outputs(9948)) or (layer0_outputs(4440)));
    layer1_outputs(3181) <= (layer0_outputs(2078)) and (layer0_outputs(8133));
    layer1_outputs(3182) <= not(layer0_outputs(1685)) or (layer0_outputs(2513));
    layer1_outputs(3183) <= '0';
    layer1_outputs(3184) <= not((layer0_outputs(6200)) and (layer0_outputs(10091)));
    layer1_outputs(3185) <= (layer0_outputs(8986)) or (layer0_outputs(5593));
    layer1_outputs(3186) <= layer0_outputs(7201);
    layer1_outputs(3187) <= not(layer0_outputs(12162));
    layer1_outputs(3188) <= '0';
    layer1_outputs(3189) <= not((layer0_outputs(9485)) xor (layer0_outputs(796)));
    layer1_outputs(3190) <= not((layer0_outputs(11757)) and (layer0_outputs(8757)));
    layer1_outputs(3191) <= layer0_outputs(2694);
    layer1_outputs(3192) <= not((layer0_outputs(2919)) or (layer0_outputs(3170)));
    layer1_outputs(3193) <= (layer0_outputs(2652)) or (layer0_outputs(6104));
    layer1_outputs(3194) <= (layer0_outputs(6915)) and (layer0_outputs(6822));
    layer1_outputs(3195) <= not(layer0_outputs(4810)) or (layer0_outputs(6835));
    layer1_outputs(3196) <= (layer0_outputs(3684)) xor (layer0_outputs(8121));
    layer1_outputs(3197) <= layer0_outputs(9571);
    layer1_outputs(3198) <= not(layer0_outputs(2591));
    layer1_outputs(3199) <= layer0_outputs(4681);
    layer1_outputs(3200) <= not((layer0_outputs(7210)) or (layer0_outputs(11305)));
    layer1_outputs(3201) <= not(layer0_outputs(11280)) or (layer0_outputs(10040));
    layer1_outputs(3202) <= layer0_outputs(10529);
    layer1_outputs(3203) <= not((layer0_outputs(2979)) and (layer0_outputs(53)));
    layer1_outputs(3204) <= (layer0_outputs(2220)) and not (layer0_outputs(259));
    layer1_outputs(3205) <= not((layer0_outputs(11321)) or (layer0_outputs(10038)));
    layer1_outputs(3206) <= layer0_outputs(2399);
    layer1_outputs(3207) <= not(layer0_outputs(12282));
    layer1_outputs(3208) <= layer0_outputs(7911);
    layer1_outputs(3209) <= not(layer0_outputs(1877));
    layer1_outputs(3210) <= not((layer0_outputs(6181)) xor (layer0_outputs(709)));
    layer1_outputs(3211) <= not(layer0_outputs(6164)) or (layer0_outputs(12256));
    layer1_outputs(3212) <= not(layer0_outputs(2084)) or (layer0_outputs(4980));
    layer1_outputs(3213) <= not(layer0_outputs(9097));
    layer1_outputs(3214) <= (layer0_outputs(913)) and not (layer0_outputs(7791));
    layer1_outputs(3215) <= layer0_outputs(1119);
    layer1_outputs(3216) <= not((layer0_outputs(4340)) and (layer0_outputs(7323)));
    layer1_outputs(3217) <= layer0_outputs(2546);
    layer1_outputs(3218) <= not(layer0_outputs(8246)) or (layer0_outputs(10339));
    layer1_outputs(3219) <= not((layer0_outputs(489)) and (layer0_outputs(10084)));
    layer1_outputs(3220) <= layer0_outputs(10782);
    layer1_outputs(3221) <= layer0_outputs(8047);
    layer1_outputs(3222) <= (layer0_outputs(8507)) xor (layer0_outputs(8254));
    layer1_outputs(3223) <= not(layer0_outputs(4602));
    layer1_outputs(3224) <= (layer0_outputs(8336)) xor (layer0_outputs(1171));
    layer1_outputs(3225) <= not(layer0_outputs(6819));
    layer1_outputs(3226) <= (layer0_outputs(2366)) or (layer0_outputs(11094));
    layer1_outputs(3227) <= not(layer0_outputs(7017));
    layer1_outputs(3228) <= not((layer0_outputs(9529)) or (layer0_outputs(677)));
    layer1_outputs(3229) <= (layer0_outputs(6123)) or (layer0_outputs(4560));
    layer1_outputs(3230) <= (layer0_outputs(1263)) xor (layer0_outputs(2669));
    layer1_outputs(3231) <= (layer0_outputs(593)) or (layer0_outputs(805));
    layer1_outputs(3232) <= not(layer0_outputs(8147));
    layer1_outputs(3233) <= not(layer0_outputs(2639)) or (layer0_outputs(2356));
    layer1_outputs(3234) <= not((layer0_outputs(876)) xor (layer0_outputs(5775)));
    layer1_outputs(3235) <= (layer0_outputs(10063)) and not (layer0_outputs(6476));
    layer1_outputs(3236) <= not(layer0_outputs(5286));
    layer1_outputs(3237) <= layer0_outputs(824);
    layer1_outputs(3238) <= not(layer0_outputs(5867));
    layer1_outputs(3239) <= not(layer0_outputs(12496)) or (layer0_outputs(11386));
    layer1_outputs(3240) <= (layer0_outputs(9219)) and not (layer0_outputs(10257));
    layer1_outputs(3241) <= not((layer0_outputs(11877)) and (layer0_outputs(10949)));
    layer1_outputs(3242) <= not((layer0_outputs(6275)) or (layer0_outputs(11445)));
    layer1_outputs(3243) <= not(layer0_outputs(4469));
    layer1_outputs(3244) <= (layer0_outputs(12326)) xor (layer0_outputs(4645));
    layer1_outputs(3245) <= not(layer0_outputs(9108));
    layer1_outputs(3246) <= layer0_outputs(1218);
    layer1_outputs(3247) <= not(layer0_outputs(6540));
    layer1_outputs(3248) <= (layer0_outputs(9508)) and not (layer0_outputs(11406));
    layer1_outputs(3249) <= layer0_outputs(948);
    layer1_outputs(3250) <= not(layer0_outputs(290));
    layer1_outputs(3251) <= (layer0_outputs(3277)) and not (layer0_outputs(8900));
    layer1_outputs(3252) <= not((layer0_outputs(9191)) and (layer0_outputs(7097)));
    layer1_outputs(3253) <= layer0_outputs(647);
    layer1_outputs(3254) <= (layer0_outputs(10268)) and not (layer0_outputs(8648));
    layer1_outputs(3255) <= (layer0_outputs(6990)) and not (layer0_outputs(5533));
    layer1_outputs(3256) <= layer0_outputs(6637);
    layer1_outputs(3257) <= not(layer0_outputs(7574));
    layer1_outputs(3258) <= not(layer0_outputs(11177));
    layer1_outputs(3259) <= not((layer0_outputs(9280)) xor (layer0_outputs(3467)));
    layer1_outputs(3260) <= layer0_outputs(4349);
    layer1_outputs(3261) <= not((layer0_outputs(3842)) or (layer0_outputs(481)));
    layer1_outputs(3262) <= (layer0_outputs(801)) and not (layer0_outputs(1232));
    layer1_outputs(3263) <= not((layer0_outputs(4105)) or (layer0_outputs(9136)));
    layer1_outputs(3264) <= '0';
    layer1_outputs(3265) <= layer0_outputs(3153);
    layer1_outputs(3266) <= (layer0_outputs(4821)) and not (layer0_outputs(10357));
    layer1_outputs(3267) <= not((layer0_outputs(11651)) and (layer0_outputs(12703)));
    layer1_outputs(3268) <= not(layer0_outputs(6016));
    layer1_outputs(3269) <= not(layer0_outputs(11598)) or (layer0_outputs(10641));
    layer1_outputs(3270) <= (layer0_outputs(10937)) and not (layer0_outputs(10147));
    layer1_outputs(3271) <= (layer0_outputs(102)) and not (layer0_outputs(4681));
    layer1_outputs(3272) <= (layer0_outputs(9325)) and not (layer0_outputs(9838));
    layer1_outputs(3273) <= not(layer0_outputs(2348)) or (layer0_outputs(1160));
    layer1_outputs(3274) <= not((layer0_outputs(8628)) or (layer0_outputs(9177)));
    layer1_outputs(3275) <= layer0_outputs(934);
    layer1_outputs(3276) <= '1';
    layer1_outputs(3277) <= not(layer0_outputs(54)) or (layer0_outputs(7709));
    layer1_outputs(3278) <= layer0_outputs(1602);
    layer1_outputs(3279) <= (layer0_outputs(6580)) and not (layer0_outputs(3315));
    layer1_outputs(3280) <= not(layer0_outputs(10083)) or (layer0_outputs(10618));
    layer1_outputs(3281) <= layer0_outputs(12444);
    layer1_outputs(3282) <= (layer0_outputs(7556)) xor (layer0_outputs(2143));
    layer1_outputs(3283) <= layer0_outputs(11766);
    layer1_outputs(3284) <= layer0_outputs(1402);
    layer1_outputs(3285) <= layer0_outputs(12239);
    layer1_outputs(3286) <= not((layer0_outputs(10051)) or (layer0_outputs(1123)));
    layer1_outputs(3287) <= layer0_outputs(4577);
    layer1_outputs(3288) <= layer0_outputs(9355);
    layer1_outputs(3289) <= not((layer0_outputs(3329)) and (layer0_outputs(7764)));
    layer1_outputs(3290) <= not(layer0_outputs(7277));
    layer1_outputs(3291) <= layer0_outputs(5815);
    layer1_outputs(3292) <= (layer0_outputs(7079)) xor (layer0_outputs(705));
    layer1_outputs(3293) <= not(layer0_outputs(1834)) or (layer0_outputs(6115));
    layer1_outputs(3294) <= not((layer0_outputs(9700)) and (layer0_outputs(2445)));
    layer1_outputs(3295) <= not((layer0_outputs(6416)) or (layer0_outputs(11200)));
    layer1_outputs(3296) <= (layer0_outputs(1420)) xor (layer0_outputs(11198));
    layer1_outputs(3297) <= layer0_outputs(770);
    layer1_outputs(3298) <= (layer0_outputs(3917)) or (layer0_outputs(9921));
    layer1_outputs(3299) <= not(layer0_outputs(12102));
    layer1_outputs(3300) <= layer0_outputs(4141);
    layer1_outputs(3301) <= not((layer0_outputs(3672)) and (layer0_outputs(847)));
    layer1_outputs(3302) <= not((layer0_outputs(8430)) or (layer0_outputs(4457)));
    layer1_outputs(3303) <= not((layer0_outputs(8469)) xor (layer0_outputs(10381)));
    layer1_outputs(3304) <= layer0_outputs(10287);
    layer1_outputs(3305) <= (layer0_outputs(4953)) or (layer0_outputs(12180));
    layer1_outputs(3306) <= layer0_outputs(6322);
    layer1_outputs(3307) <= (layer0_outputs(11226)) or (layer0_outputs(8758));
    layer1_outputs(3308) <= (layer0_outputs(4825)) xor (layer0_outputs(8443));
    layer1_outputs(3309) <= not(layer0_outputs(8949));
    layer1_outputs(3310) <= not(layer0_outputs(7268)) or (layer0_outputs(8033));
    layer1_outputs(3311) <= layer0_outputs(2530);
    layer1_outputs(3312) <= '1';
    layer1_outputs(3313) <= (layer0_outputs(8049)) or (layer0_outputs(10573));
    layer1_outputs(3314) <= not((layer0_outputs(2390)) xor (layer0_outputs(3236)));
    layer1_outputs(3315) <= not((layer0_outputs(2950)) xor (layer0_outputs(4699)));
    layer1_outputs(3316) <= layer0_outputs(5204);
    layer1_outputs(3317) <= (layer0_outputs(5128)) and not (layer0_outputs(424));
    layer1_outputs(3318) <= (layer0_outputs(11348)) or (layer0_outputs(9111));
    layer1_outputs(3319) <= not(layer0_outputs(2766));
    layer1_outputs(3320) <= (layer0_outputs(4682)) and not (layer0_outputs(4358));
    layer1_outputs(3321) <= not((layer0_outputs(4789)) and (layer0_outputs(9360)));
    layer1_outputs(3322) <= not(layer0_outputs(2783));
    layer1_outputs(3323) <= layer0_outputs(11849);
    layer1_outputs(3324) <= not(layer0_outputs(7115)) or (layer0_outputs(7454));
    layer1_outputs(3325) <= not(layer0_outputs(8466));
    layer1_outputs(3326) <= not((layer0_outputs(6752)) or (layer0_outputs(5905)));
    layer1_outputs(3327) <= layer0_outputs(3495);
    layer1_outputs(3328) <= not(layer0_outputs(9411)) or (layer0_outputs(62));
    layer1_outputs(3329) <= layer0_outputs(3051);
    layer1_outputs(3330) <= not(layer0_outputs(11062)) or (layer0_outputs(8265));
    layer1_outputs(3331) <= not(layer0_outputs(11479)) or (layer0_outputs(3427));
    layer1_outputs(3332) <= (layer0_outputs(6103)) xor (layer0_outputs(9451));
    layer1_outputs(3333) <= not(layer0_outputs(2940)) or (layer0_outputs(1801));
    layer1_outputs(3334) <= not(layer0_outputs(1248));
    layer1_outputs(3335) <= not(layer0_outputs(6560));
    layer1_outputs(3336) <= '1';
    layer1_outputs(3337) <= not((layer0_outputs(461)) and (layer0_outputs(4951)));
    layer1_outputs(3338) <= (layer0_outputs(12522)) or (layer0_outputs(2240));
    layer1_outputs(3339) <= not(layer0_outputs(2695));
    layer1_outputs(3340) <= layer0_outputs(8701);
    layer1_outputs(3341) <= layer0_outputs(9673);
    layer1_outputs(3342) <= not(layer0_outputs(12635)) or (layer0_outputs(3144));
    layer1_outputs(3343) <= (layer0_outputs(11436)) and (layer0_outputs(10563));
    layer1_outputs(3344) <= not(layer0_outputs(12361)) or (layer0_outputs(2765));
    layer1_outputs(3345) <= not((layer0_outputs(6185)) or (layer0_outputs(11236)));
    layer1_outputs(3346) <= layer0_outputs(3502);
    layer1_outputs(3347) <= not(layer0_outputs(9159));
    layer1_outputs(3348) <= layer0_outputs(1609);
    layer1_outputs(3349) <= (layer0_outputs(5291)) or (layer0_outputs(901));
    layer1_outputs(3350) <= not((layer0_outputs(12091)) xor (layer0_outputs(1301)));
    layer1_outputs(3351) <= layer0_outputs(8022);
    layer1_outputs(3352) <= not(layer0_outputs(4374)) or (layer0_outputs(875));
    layer1_outputs(3353) <= not(layer0_outputs(11309));
    layer1_outputs(3354) <= not((layer0_outputs(6826)) or (layer0_outputs(9709)));
    layer1_outputs(3355) <= not((layer0_outputs(2308)) or (layer0_outputs(2019)));
    layer1_outputs(3356) <= not(layer0_outputs(1361));
    layer1_outputs(3357) <= (layer0_outputs(2864)) and (layer0_outputs(3623));
    layer1_outputs(3358) <= (layer0_outputs(12195)) and not (layer0_outputs(11771));
    layer1_outputs(3359) <= not((layer0_outputs(3187)) or (layer0_outputs(8707)));
    layer1_outputs(3360) <= layer0_outputs(11368);
    layer1_outputs(3361) <= (layer0_outputs(6121)) xor (layer0_outputs(8464));
    layer1_outputs(3362) <= not(layer0_outputs(4075));
    layer1_outputs(3363) <= (layer0_outputs(1266)) and not (layer0_outputs(4658));
    layer1_outputs(3364) <= not((layer0_outputs(251)) xor (layer0_outputs(2101)));
    layer1_outputs(3365) <= not((layer0_outputs(5437)) or (layer0_outputs(9216)));
    layer1_outputs(3366) <= layer0_outputs(4180);
    layer1_outputs(3367) <= not((layer0_outputs(1271)) or (layer0_outputs(9210)));
    layer1_outputs(3368) <= not(layer0_outputs(2628));
    layer1_outputs(3369) <= (layer0_outputs(933)) and not (layer0_outputs(12763));
    layer1_outputs(3370) <= not(layer0_outputs(6088));
    layer1_outputs(3371) <= layer0_outputs(10889);
    layer1_outputs(3372) <= (layer0_outputs(7076)) and not (layer0_outputs(4812));
    layer1_outputs(3373) <= (layer0_outputs(9260)) and (layer0_outputs(4763));
    layer1_outputs(3374) <= layer0_outputs(9858);
    layer1_outputs(3375) <= (layer0_outputs(3961)) xor (layer0_outputs(9427));
    layer1_outputs(3376) <= not((layer0_outputs(4545)) and (layer0_outputs(9031)));
    layer1_outputs(3377) <= layer0_outputs(4151);
    layer1_outputs(3378) <= not(layer0_outputs(5136));
    layer1_outputs(3379) <= (layer0_outputs(6575)) or (layer0_outputs(183));
    layer1_outputs(3380) <= not(layer0_outputs(5749));
    layer1_outputs(3381) <= not((layer0_outputs(3402)) or (layer0_outputs(12005)));
    layer1_outputs(3382) <= not((layer0_outputs(11135)) xor (layer0_outputs(7650)));
    layer1_outputs(3383) <= (layer0_outputs(883)) xor (layer0_outputs(392));
    layer1_outputs(3384) <= not(layer0_outputs(11683)) or (layer0_outputs(10994));
    layer1_outputs(3385) <= not(layer0_outputs(2252));
    layer1_outputs(3386) <= not(layer0_outputs(9975));
    layer1_outputs(3387) <= layer0_outputs(9003);
    layer1_outputs(3388) <= '0';
    layer1_outputs(3389) <= not(layer0_outputs(9497));
    layer1_outputs(3390) <= (layer0_outputs(9568)) and (layer0_outputs(3741));
    layer1_outputs(3391) <= layer0_outputs(6111);
    layer1_outputs(3392) <= not(layer0_outputs(7429));
    layer1_outputs(3393) <= (layer0_outputs(11283)) and not (layer0_outputs(6956));
    layer1_outputs(3394) <= not((layer0_outputs(528)) xor (layer0_outputs(1241)));
    layer1_outputs(3395) <= not(layer0_outputs(10282));
    layer1_outputs(3396) <= (layer0_outputs(7241)) and not (layer0_outputs(9883));
    layer1_outputs(3397) <= not(layer0_outputs(12497));
    layer1_outputs(3398) <= (layer0_outputs(3686)) and not (layer0_outputs(5846));
    layer1_outputs(3399) <= not((layer0_outputs(3580)) and (layer0_outputs(5066)));
    layer1_outputs(3400) <= (layer0_outputs(1842)) and (layer0_outputs(11314));
    layer1_outputs(3401) <= layer0_outputs(4341);
    layer1_outputs(3402) <= (layer0_outputs(5766)) or (layer0_outputs(9759));
    layer1_outputs(3403) <= (layer0_outputs(8267)) and not (layer0_outputs(9959));
    layer1_outputs(3404) <= not(layer0_outputs(10897)) or (layer0_outputs(10728));
    layer1_outputs(3405) <= layer0_outputs(12703);
    layer1_outputs(3406) <= not(layer0_outputs(7370)) or (layer0_outputs(8086));
    layer1_outputs(3407) <= (layer0_outputs(9849)) or (layer0_outputs(2942));
    layer1_outputs(3408) <= (layer0_outputs(10754)) and not (layer0_outputs(4616));
    layer1_outputs(3409) <= not((layer0_outputs(8731)) xor (layer0_outputs(832)));
    layer1_outputs(3410) <= (layer0_outputs(5834)) and (layer0_outputs(10165));
    layer1_outputs(3411) <= layer0_outputs(12011);
    layer1_outputs(3412) <= '0';
    layer1_outputs(3413) <= not(layer0_outputs(7075));
    layer1_outputs(3414) <= not(layer0_outputs(7144)) or (layer0_outputs(10784));
    layer1_outputs(3415) <= not((layer0_outputs(1568)) and (layer0_outputs(3562)));
    layer1_outputs(3416) <= (layer0_outputs(6155)) and not (layer0_outputs(12784));
    layer1_outputs(3417) <= not(layer0_outputs(4352));
    layer1_outputs(3418) <= not(layer0_outputs(7288)) or (layer0_outputs(10004));
    layer1_outputs(3419) <= not(layer0_outputs(7337)) or (layer0_outputs(6118));
    layer1_outputs(3420) <= not(layer0_outputs(4193)) or (layer0_outputs(12588));
    layer1_outputs(3421) <= layer0_outputs(604);
    layer1_outputs(3422) <= not(layer0_outputs(4245));
    layer1_outputs(3423) <= not((layer0_outputs(12527)) and (layer0_outputs(1571)));
    layer1_outputs(3424) <= not(layer0_outputs(8137)) or (layer0_outputs(11909));
    layer1_outputs(3425) <= not(layer0_outputs(2532));
    layer1_outputs(3426) <= not((layer0_outputs(9255)) xor (layer0_outputs(9762)));
    layer1_outputs(3427) <= (layer0_outputs(130)) xor (layer0_outputs(6419));
    layer1_outputs(3428) <= not(layer0_outputs(11150)) or (layer0_outputs(8547));
    layer1_outputs(3429) <= layer0_outputs(11574);
    layer1_outputs(3430) <= layer0_outputs(1258);
    layer1_outputs(3431) <= not(layer0_outputs(656)) or (layer0_outputs(11199));
    layer1_outputs(3432) <= layer0_outputs(1531);
    layer1_outputs(3433) <= not((layer0_outputs(833)) and (layer0_outputs(5028)));
    layer1_outputs(3434) <= (layer0_outputs(6593)) and (layer0_outputs(5796));
    layer1_outputs(3435) <= not((layer0_outputs(10006)) and (layer0_outputs(2168)));
    layer1_outputs(3436) <= not(layer0_outputs(7929));
    layer1_outputs(3437) <= not((layer0_outputs(11975)) xor (layer0_outputs(6437)));
    layer1_outputs(3438) <= (layer0_outputs(2010)) and (layer0_outputs(5633));
    layer1_outputs(3439) <= layer0_outputs(8458);
    layer1_outputs(3440) <= (layer0_outputs(6128)) and (layer0_outputs(2832));
    layer1_outputs(3441) <= '1';
    layer1_outputs(3442) <= not(layer0_outputs(12053));
    layer1_outputs(3443) <= not(layer0_outputs(6652)) or (layer0_outputs(7306));
    layer1_outputs(3444) <= not(layer0_outputs(1679));
    layer1_outputs(3445) <= not(layer0_outputs(7626));
    layer1_outputs(3446) <= (layer0_outputs(4020)) or (layer0_outputs(285));
    layer1_outputs(3447) <= (layer0_outputs(11609)) and (layer0_outputs(10722));
    layer1_outputs(3448) <= not(layer0_outputs(8854));
    layer1_outputs(3449) <= (layer0_outputs(2308)) and not (layer0_outputs(6539));
    layer1_outputs(3450) <= layer0_outputs(3765);
    layer1_outputs(3451) <= (layer0_outputs(1290)) and not (layer0_outputs(1618));
    layer1_outputs(3452) <= not(layer0_outputs(984)) or (layer0_outputs(8073));
    layer1_outputs(3453) <= layer0_outputs(918);
    layer1_outputs(3454) <= not((layer0_outputs(275)) or (layer0_outputs(6290)));
    layer1_outputs(3455) <= not(layer0_outputs(9153));
    layer1_outputs(3456) <= layer0_outputs(9740);
    layer1_outputs(3457) <= '0';
    layer1_outputs(3458) <= not(layer0_outputs(6803));
    layer1_outputs(3459) <= (layer0_outputs(9827)) and (layer0_outputs(4242));
    layer1_outputs(3460) <= not(layer0_outputs(1679));
    layer1_outputs(3461) <= not((layer0_outputs(9154)) or (layer0_outputs(5627)));
    layer1_outputs(3462) <= not((layer0_outputs(1483)) xor (layer0_outputs(2799)));
    layer1_outputs(3463) <= not(layer0_outputs(5950));
    layer1_outputs(3464) <= not((layer0_outputs(4969)) and (layer0_outputs(8380)));
    layer1_outputs(3465) <= layer0_outputs(6673);
    layer1_outputs(3466) <= layer0_outputs(9654);
    layer1_outputs(3467) <= (layer0_outputs(7462)) and not (layer0_outputs(6282));
    layer1_outputs(3468) <= not(layer0_outputs(4539));
    layer1_outputs(3469) <= (layer0_outputs(8392)) or (layer0_outputs(3915));
    layer1_outputs(3470) <= not(layer0_outputs(9749));
    layer1_outputs(3471) <= not((layer0_outputs(2922)) xor (layer0_outputs(1562)));
    layer1_outputs(3472) <= layer0_outputs(12122);
    layer1_outputs(3473) <= (layer0_outputs(2023)) and not (layer0_outputs(5147));
    layer1_outputs(3474) <= layer0_outputs(2319);
    layer1_outputs(3475) <= (layer0_outputs(2661)) or (layer0_outputs(8745));
    layer1_outputs(3476) <= (layer0_outputs(480)) and not (layer0_outputs(3246));
    layer1_outputs(3477) <= (layer0_outputs(10089)) and not (layer0_outputs(3767));
    layer1_outputs(3478) <= not(layer0_outputs(2074)) or (layer0_outputs(10969));
    layer1_outputs(3479) <= not(layer0_outputs(2404));
    layer1_outputs(3480) <= not((layer0_outputs(10580)) or (layer0_outputs(12709)));
    layer1_outputs(3481) <= (layer0_outputs(9586)) and not (layer0_outputs(6037));
    layer1_outputs(3482) <= not((layer0_outputs(3372)) or (layer0_outputs(4607)));
    layer1_outputs(3483) <= layer0_outputs(8742);
    layer1_outputs(3484) <= not(layer0_outputs(1218));
    layer1_outputs(3485) <= (layer0_outputs(9270)) and not (layer0_outputs(2839));
    layer1_outputs(3486) <= (layer0_outputs(3670)) and not (layer0_outputs(2818));
    layer1_outputs(3487) <= layer0_outputs(4848);
    layer1_outputs(3488) <= (layer0_outputs(10754)) and not (layer0_outputs(9256));
    layer1_outputs(3489) <= not((layer0_outputs(3069)) and (layer0_outputs(6478)));
    layer1_outputs(3490) <= '1';
    layer1_outputs(3491) <= not(layer0_outputs(9250)) or (layer0_outputs(6761));
    layer1_outputs(3492) <= not(layer0_outputs(2919));
    layer1_outputs(3493) <= not(layer0_outputs(6314)) or (layer0_outputs(463));
    layer1_outputs(3494) <= (layer0_outputs(12776)) xor (layer0_outputs(1004));
    layer1_outputs(3495) <= layer0_outputs(4277);
    layer1_outputs(3496) <= (layer0_outputs(8518)) xor (layer0_outputs(9221));
    layer1_outputs(3497) <= (layer0_outputs(3026)) and not (layer0_outputs(4803));
    layer1_outputs(3498) <= not((layer0_outputs(11802)) xor (layer0_outputs(11861)));
    layer1_outputs(3499) <= (layer0_outputs(5947)) and not (layer0_outputs(8384));
    layer1_outputs(3500) <= not((layer0_outputs(8376)) and (layer0_outputs(8004)));
    layer1_outputs(3501) <= not((layer0_outputs(4511)) or (layer0_outputs(1184)));
    layer1_outputs(3502) <= layer0_outputs(10252);
    layer1_outputs(3503) <= (layer0_outputs(12277)) or (layer0_outputs(3146));
    layer1_outputs(3504) <= (layer0_outputs(4615)) and not (layer0_outputs(10921));
    layer1_outputs(3505) <= layer0_outputs(2251);
    layer1_outputs(3506) <= '1';
    layer1_outputs(3507) <= (layer0_outputs(4986)) and (layer0_outputs(763));
    layer1_outputs(3508) <= (layer0_outputs(3114)) and (layer0_outputs(1546));
    layer1_outputs(3509) <= (layer0_outputs(12711)) xor (layer0_outputs(11532));
    layer1_outputs(3510) <= not(layer0_outputs(7489)) or (layer0_outputs(10433));
    layer1_outputs(3511) <= (layer0_outputs(6187)) and not (layer0_outputs(76));
    layer1_outputs(3512) <= (layer0_outputs(4027)) or (layer0_outputs(10195));
    layer1_outputs(3513) <= (layer0_outputs(3860)) and (layer0_outputs(8629));
    layer1_outputs(3514) <= layer0_outputs(1661);
    layer1_outputs(3515) <= (layer0_outputs(3601)) and not (layer0_outputs(867));
    layer1_outputs(3516) <= (layer0_outputs(9954)) or (layer0_outputs(5842));
    layer1_outputs(3517) <= '0';
    layer1_outputs(3518) <= '0';
    layer1_outputs(3519) <= not((layer0_outputs(2371)) or (layer0_outputs(1439)));
    layer1_outputs(3520) <= (layer0_outputs(2242)) xor (layer0_outputs(4508));
    layer1_outputs(3521) <= not((layer0_outputs(5293)) or (layer0_outputs(4238)));
    layer1_outputs(3522) <= (layer0_outputs(10015)) xor (layer0_outputs(8587));
    layer1_outputs(3523) <= not(layer0_outputs(4364)) or (layer0_outputs(2130));
    layer1_outputs(3524) <= layer0_outputs(7139);
    layer1_outputs(3525) <= (layer0_outputs(5406)) and (layer0_outputs(1268));
    layer1_outputs(3526) <= not(layer0_outputs(810));
    layer1_outputs(3527) <= layer0_outputs(12711);
    layer1_outputs(3528) <= (layer0_outputs(3683)) and not (layer0_outputs(7808));
    layer1_outputs(3529) <= layer0_outputs(6959);
    layer1_outputs(3530) <= not(layer0_outputs(11027)) or (layer0_outputs(10177));
    layer1_outputs(3531) <= not(layer0_outputs(10362));
    layer1_outputs(3532) <= not(layer0_outputs(5121)) or (layer0_outputs(9994));
    layer1_outputs(3533) <= '1';
    layer1_outputs(3534) <= not(layer0_outputs(4993));
    layer1_outputs(3535) <= '0';
    layer1_outputs(3536) <= '1';
    layer1_outputs(3537) <= not((layer0_outputs(2268)) and (layer0_outputs(10681)));
    layer1_outputs(3538) <= layer0_outputs(10404);
    layer1_outputs(3539) <= (layer0_outputs(12019)) xor (layer0_outputs(766));
    layer1_outputs(3540) <= not((layer0_outputs(1222)) xor (layer0_outputs(7493)));
    layer1_outputs(3541) <= (layer0_outputs(11393)) and (layer0_outputs(4505));
    layer1_outputs(3542) <= not((layer0_outputs(1797)) xor (layer0_outputs(12318)));
    layer1_outputs(3543) <= layer0_outputs(3245);
    layer1_outputs(3544) <= not(layer0_outputs(12648)) or (layer0_outputs(5646));
    layer1_outputs(3545) <= layer0_outputs(3659);
    layer1_outputs(3546) <= not((layer0_outputs(1193)) xor (layer0_outputs(316)));
    layer1_outputs(3547) <= (layer0_outputs(11322)) and (layer0_outputs(516));
    layer1_outputs(3548) <= not((layer0_outputs(7936)) xor (layer0_outputs(2845)));
    layer1_outputs(3549) <= not((layer0_outputs(11088)) and (layer0_outputs(10395)));
    layer1_outputs(3550) <= not(layer0_outputs(3825));
    layer1_outputs(3551) <= not(layer0_outputs(6730));
    layer1_outputs(3552) <= not(layer0_outputs(7231));
    layer1_outputs(3553) <= layer0_outputs(3674);
    layer1_outputs(3554) <= (layer0_outputs(9583)) or (layer0_outputs(10598));
    layer1_outputs(3555) <= '0';
    layer1_outputs(3556) <= layer0_outputs(11593);
    layer1_outputs(3557) <= (layer0_outputs(4240)) or (layer0_outputs(1109));
    layer1_outputs(3558) <= (layer0_outputs(3442)) and (layer0_outputs(4513));
    layer1_outputs(3559) <= not(layer0_outputs(5260)) or (layer0_outputs(2305));
    layer1_outputs(3560) <= not((layer0_outputs(6367)) xor (layer0_outputs(3041)));
    layer1_outputs(3561) <= (layer0_outputs(3577)) or (layer0_outputs(1518));
    layer1_outputs(3562) <= (layer0_outputs(5771)) and (layer0_outputs(8580));
    layer1_outputs(3563) <= layer0_outputs(1808);
    layer1_outputs(3564) <= not(layer0_outputs(18));
    layer1_outputs(3565) <= not(layer0_outputs(11605));
    layer1_outputs(3566) <= '1';
    layer1_outputs(3567) <= not(layer0_outputs(2152));
    layer1_outputs(3568) <= not((layer0_outputs(1844)) or (layer0_outputs(6747)));
    layer1_outputs(3569) <= (layer0_outputs(566)) xor (layer0_outputs(8024));
    layer1_outputs(3570) <= layer0_outputs(6782);
    layer1_outputs(3571) <= layer0_outputs(2500);
    layer1_outputs(3572) <= layer0_outputs(1530);
    layer1_outputs(3573) <= not(layer0_outputs(7683));
    layer1_outputs(3574) <= (layer0_outputs(1115)) xor (layer0_outputs(2599));
    layer1_outputs(3575) <= (layer0_outputs(7897)) and not (layer0_outputs(11195));
    layer1_outputs(3576) <= not(layer0_outputs(8375)) or (layer0_outputs(11676));
    layer1_outputs(3577) <= (layer0_outputs(7993)) or (layer0_outputs(99));
    layer1_outputs(3578) <= layer0_outputs(5911);
    layer1_outputs(3579) <= layer0_outputs(9618);
    layer1_outputs(3580) <= (layer0_outputs(7123)) and not (layer0_outputs(1100));
    layer1_outputs(3581) <= (layer0_outputs(10356)) or (layer0_outputs(8467));
    layer1_outputs(3582) <= (layer0_outputs(2050)) and (layer0_outputs(2218));
    layer1_outputs(3583) <= '0';
    layer1_outputs(3584) <= layer0_outputs(9455);
    layer1_outputs(3585) <= (layer0_outputs(8308)) xor (layer0_outputs(2773));
    layer1_outputs(3586) <= not((layer0_outputs(11277)) xor (layer0_outputs(894)));
    layer1_outputs(3587) <= not(layer0_outputs(12429));
    layer1_outputs(3588) <= not(layer0_outputs(6709)) or (layer0_outputs(8585));
    layer1_outputs(3589) <= not(layer0_outputs(10527));
    layer1_outputs(3590) <= layer0_outputs(9595);
    layer1_outputs(3591) <= not(layer0_outputs(8888)) or (layer0_outputs(4706));
    layer1_outputs(3592) <= (layer0_outputs(2112)) and (layer0_outputs(8537));
    layer1_outputs(3593) <= layer0_outputs(10104);
    layer1_outputs(3594) <= (layer0_outputs(4322)) and (layer0_outputs(7440));
    layer1_outputs(3595) <= (layer0_outputs(3000)) xor (layer0_outputs(11937));
    layer1_outputs(3596) <= not(layer0_outputs(1775)) or (layer0_outputs(11750));
    layer1_outputs(3597) <= not((layer0_outputs(12794)) xor (layer0_outputs(7630)));
    layer1_outputs(3598) <= (layer0_outputs(6288)) or (layer0_outputs(11848));
    layer1_outputs(3599) <= (layer0_outputs(7105)) and (layer0_outputs(945));
    layer1_outputs(3600) <= (layer0_outputs(12468)) and (layer0_outputs(6303));
    layer1_outputs(3601) <= not(layer0_outputs(830));
    layer1_outputs(3602) <= not((layer0_outputs(12054)) and (layer0_outputs(8468)));
    layer1_outputs(3603) <= (layer0_outputs(4067)) or (layer0_outputs(11237));
    layer1_outputs(3604) <= not(layer0_outputs(4560)) or (layer0_outputs(9553));
    layer1_outputs(3605) <= '0';
    layer1_outputs(3606) <= layer0_outputs(8215);
    layer1_outputs(3607) <= layer0_outputs(11637);
    layer1_outputs(3608) <= (layer0_outputs(2891)) xor (layer0_outputs(10396));
    layer1_outputs(3609) <= not((layer0_outputs(6239)) xor (layer0_outputs(6053)));
    layer1_outputs(3610) <= not(layer0_outputs(5382)) or (layer0_outputs(3811));
    layer1_outputs(3611) <= not(layer0_outputs(1078)) or (layer0_outputs(7970));
    layer1_outputs(3612) <= layer0_outputs(10788);
    layer1_outputs(3613) <= not((layer0_outputs(6337)) and (layer0_outputs(7917)));
    layer1_outputs(3614) <= layer0_outputs(8550);
    layer1_outputs(3615) <= not((layer0_outputs(10956)) xor (layer0_outputs(9570)));
    layer1_outputs(3616) <= layer0_outputs(10890);
    layer1_outputs(3617) <= layer0_outputs(8144);
    layer1_outputs(3618) <= (layer0_outputs(3230)) or (layer0_outputs(9756));
    layer1_outputs(3619) <= not(layer0_outputs(9495)) or (layer0_outputs(7188));
    layer1_outputs(3620) <= '1';
    layer1_outputs(3621) <= layer0_outputs(4425);
    layer1_outputs(3622) <= (layer0_outputs(1145)) or (layer0_outputs(1111));
    layer1_outputs(3623) <= not((layer0_outputs(5924)) and (layer0_outputs(2707)));
    layer1_outputs(3624) <= layer0_outputs(5923);
    layer1_outputs(3625) <= (layer0_outputs(4904)) and not (layer0_outputs(337));
    layer1_outputs(3626) <= (layer0_outputs(4695)) and not (layer0_outputs(10990));
    layer1_outputs(3627) <= not(layer0_outputs(2651));
    layer1_outputs(3628) <= layer0_outputs(7073);
    layer1_outputs(3629) <= not(layer0_outputs(10747));
    layer1_outputs(3630) <= layer0_outputs(4121);
    layer1_outputs(3631) <= (layer0_outputs(2344)) or (layer0_outputs(3085));
    layer1_outputs(3632) <= not(layer0_outputs(9278));
    layer1_outputs(3633) <= (layer0_outputs(6676)) xor (layer0_outputs(5498));
    layer1_outputs(3634) <= layer0_outputs(8638);
    layer1_outputs(3635) <= not((layer0_outputs(4393)) and (layer0_outputs(10035)));
    layer1_outputs(3636) <= not(layer0_outputs(10323));
    layer1_outputs(3637) <= '1';
    layer1_outputs(3638) <= layer0_outputs(10901);
    layer1_outputs(3639) <= '0';
    layer1_outputs(3640) <= not(layer0_outputs(551)) or (layer0_outputs(5132));
    layer1_outputs(3641) <= not(layer0_outputs(6343));
    layer1_outputs(3642) <= (layer0_outputs(7134)) and (layer0_outputs(1698));
    layer1_outputs(3643) <= not((layer0_outputs(3802)) and (layer0_outputs(10531)));
    layer1_outputs(3644) <= not(layer0_outputs(7941)) or (layer0_outputs(9937));
    layer1_outputs(3645) <= (layer0_outputs(6496)) or (layer0_outputs(2598));
    layer1_outputs(3646) <= not((layer0_outputs(7668)) xor (layer0_outputs(4434)));
    layer1_outputs(3647) <= not(layer0_outputs(11701));
    layer1_outputs(3648) <= not((layer0_outputs(12658)) xor (layer0_outputs(10039)));
    layer1_outputs(3649) <= not((layer0_outputs(2665)) or (layer0_outputs(5865)));
    layer1_outputs(3650) <= layer0_outputs(4934);
    layer1_outputs(3651) <= not((layer0_outputs(4465)) and (layer0_outputs(10309)));
    layer1_outputs(3652) <= not(layer0_outputs(10710));
    layer1_outputs(3653) <= not((layer0_outputs(12790)) xor (layer0_outputs(11858)));
    layer1_outputs(3654) <= (layer0_outputs(12570)) or (layer0_outputs(4132));
    layer1_outputs(3655) <= (layer0_outputs(2657)) xor (layer0_outputs(6050));
    layer1_outputs(3656) <= not(layer0_outputs(6845));
    layer1_outputs(3657) <= (layer0_outputs(5369)) xor (layer0_outputs(831));
    layer1_outputs(3658) <= (layer0_outputs(9835)) xor (layer0_outputs(4938));
    layer1_outputs(3659) <= layer0_outputs(63);
    layer1_outputs(3660) <= '0';
    layer1_outputs(3661) <= (layer0_outputs(2067)) and not (layer0_outputs(10605));
    layer1_outputs(3662) <= not(layer0_outputs(6040)) or (layer0_outputs(12515));
    layer1_outputs(3663) <= not(layer0_outputs(7558)) or (layer0_outputs(6142));
    layer1_outputs(3664) <= layer0_outputs(5658);
    layer1_outputs(3665) <= not(layer0_outputs(3748)) or (layer0_outputs(12503));
    layer1_outputs(3666) <= not((layer0_outputs(393)) and (layer0_outputs(9199)));
    layer1_outputs(3667) <= layer0_outputs(2503);
    layer1_outputs(3668) <= not((layer0_outputs(9110)) and (layer0_outputs(8452)));
    layer1_outputs(3669) <= layer0_outputs(868);
    layer1_outputs(3670) <= layer0_outputs(11687);
    layer1_outputs(3671) <= not(layer0_outputs(4664)) or (layer0_outputs(5023));
    layer1_outputs(3672) <= not(layer0_outputs(6500)) or (layer0_outputs(12017));
    layer1_outputs(3673) <= layer0_outputs(2362);
    layer1_outputs(3674) <= not(layer0_outputs(9855)) or (layer0_outputs(7805));
    layer1_outputs(3675) <= not((layer0_outputs(5096)) or (layer0_outputs(1161)));
    layer1_outputs(3676) <= layer0_outputs(822);
    layer1_outputs(3677) <= not(layer0_outputs(11649));
    layer1_outputs(3678) <= not(layer0_outputs(5950));
    layer1_outputs(3679) <= not((layer0_outputs(11600)) or (layer0_outputs(10844)));
    layer1_outputs(3680) <= not((layer0_outputs(5989)) and (layer0_outputs(12624)));
    layer1_outputs(3681) <= layer0_outputs(7145);
    layer1_outputs(3682) <= not((layer0_outputs(6940)) and (layer0_outputs(547)));
    layer1_outputs(3683) <= not(layer0_outputs(2297)) or (layer0_outputs(11435));
    layer1_outputs(3684) <= (layer0_outputs(3087)) or (layer0_outputs(3342));
    layer1_outputs(3685) <= not(layer0_outputs(11829));
    layer1_outputs(3686) <= not(layer0_outputs(8379));
    layer1_outputs(3687) <= not(layer0_outputs(1424)) or (layer0_outputs(4631));
    layer1_outputs(3688) <= (layer0_outputs(7132)) xor (layer0_outputs(5033));
    layer1_outputs(3689) <= not(layer0_outputs(4231)) or (layer0_outputs(5188));
    layer1_outputs(3690) <= (layer0_outputs(1915)) or (layer0_outputs(10770));
    layer1_outputs(3691) <= (layer0_outputs(3750)) and (layer0_outputs(5505));
    layer1_outputs(3692) <= not(layer0_outputs(10740)) or (layer0_outputs(8853));
    layer1_outputs(3693) <= layer0_outputs(11959);
    layer1_outputs(3694) <= not((layer0_outputs(7976)) xor (layer0_outputs(3165)));
    layer1_outputs(3695) <= layer0_outputs(8010);
    layer1_outputs(3696) <= not(layer0_outputs(213));
    layer1_outputs(3697) <= not(layer0_outputs(12005));
    layer1_outputs(3698) <= layer0_outputs(2433);
    layer1_outputs(3699) <= not(layer0_outputs(1713));
    layer1_outputs(3700) <= not(layer0_outputs(7980)) or (layer0_outputs(3862));
    layer1_outputs(3701) <= layer0_outputs(926);
    layer1_outputs(3702) <= '0';
    layer1_outputs(3703) <= not((layer0_outputs(5079)) xor (layer0_outputs(1223)));
    layer1_outputs(3704) <= (layer0_outputs(2638)) and (layer0_outputs(8227));
    layer1_outputs(3705) <= layer0_outputs(1255);
    layer1_outputs(3706) <= layer0_outputs(8601);
    layer1_outputs(3707) <= (layer0_outputs(7086)) and not (layer0_outputs(792));
    layer1_outputs(3708) <= layer0_outputs(10706);
    layer1_outputs(3709) <= not(layer0_outputs(908));
    layer1_outputs(3710) <= layer0_outputs(7886);
    layer1_outputs(3711) <= not(layer0_outputs(11895));
    layer1_outputs(3712) <= layer0_outputs(12545);
    layer1_outputs(3713) <= (layer0_outputs(384)) or (layer0_outputs(8340));
    layer1_outputs(3714) <= not(layer0_outputs(7727));
    layer1_outputs(3715) <= (layer0_outputs(3234)) or (layer0_outputs(10755));
    layer1_outputs(3716) <= layer0_outputs(6286);
    layer1_outputs(3717) <= not(layer0_outputs(3559));
    layer1_outputs(3718) <= not((layer0_outputs(6986)) and (layer0_outputs(5949)));
    layer1_outputs(3719) <= (layer0_outputs(1452)) xor (layer0_outputs(11792));
    layer1_outputs(3720) <= not(layer0_outputs(4031)) or (layer0_outputs(11001));
    layer1_outputs(3721) <= (layer0_outputs(8003)) xor (layer0_outputs(3157));
    layer1_outputs(3722) <= (layer0_outputs(12771)) and (layer0_outputs(10293));
    layer1_outputs(3723) <= not((layer0_outputs(4160)) xor (layer0_outputs(8462)));
    layer1_outputs(3724) <= (layer0_outputs(754)) xor (layer0_outputs(8326));
    layer1_outputs(3725) <= not((layer0_outputs(11571)) or (layer0_outputs(10746)));
    layer1_outputs(3726) <= not(layer0_outputs(11580));
    layer1_outputs(3727) <= (layer0_outputs(7830)) xor (layer0_outputs(1456));
    layer1_outputs(3728) <= (layer0_outputs(7591)) and not (layer0_outputs(5447));
    layer1_outputs(3729) <= layer0_outputs(10299);
    layer1_outputs(3730) <= layer0_outputs(7403);
    layer1_outputs(3731) <= '0';
    layer1_outputs(3732) <= not(layer0_outputs(3685));
    layer1_outputs(3733) <= '0';
    layer1_outputs(3734) <= not(layer0_outputs(47));
    layer1_outputs(3735) <= not((layer0_outputs(4358)) xor (layer0_outputs(11404)));
    layer1_outputs(3736) <= (layer0_outputs(1773)) or (layer0_outputs(2813));
    layer1_outputs(3737) <= not(layer0_outputs(6789));
    layer1_outputs(3738) <= not(layer0_outputs(1247));
    layer1_outputs(3739) <= (layer0_outputs(11029)) and not (layer0_outputs(12381));
    layer1_outputs(3740) <= not((layer0_outputs(2325)) and (layer0_outputs(8486)));
    layer1_outputs(3741) <= (layer0_outputs(10717)) xor (layer0_outputs(8794));
    layer1_outputs(3742) <= (layer0_outputs(12362)) and (layer0_outputs(1909));
    layer1_outputs(3743) <= not(layer0_outputs(1726)) or (layer0_outputs(2133));
    layer1_outputs(3744) <= '0';
    layer1_outputs(3745) <= layer0_outputs(6757);
    layer1_outputs(3746) <= layer0_outputs(2211);
    layer1_outputs(3747) <= (layer0_outputs(11649)) xor (layer0_outputs(3454));
    layer1_outputs(3748) <= not((layer0_outputs(10654)) or (layer0_outputs(6137)));
    layer1_outputs(3749) <= not((layer0_outputs(253)) xor (layer0_outputs(2798)));
    layer1_outputs(3750) <= (layer0_outputs(6256)) xor (layer0_outputs(11863));
    layer1_outputs(3751) <= (layer0_outputs(7718)) or (layer0_outputs(1021));
    layer1_outputs(3752) <= not(layer0_outputs(7526));
    layer1_outputs(3753) <= not((layer0_outputs(4753)) xor (layer0_outputs(3210)));
    layer1_outputs(3754) <= not((layer0_outputs(2273)) xor (layer0_outputs(6632)));
    layer1_outputs(3755) <= (layer0_outputs(8510)) and not (layer0_outputs(2688));
    layer1_outputs(3756) <= layer0_outputs(6304);
    layer1_outputs(3757) <= not(layer0_outputs(7598));
    layer1_outputs(3758) <= not((layer0_outputs(4624)) or (layer0_outputs(7708)));
    layer1_outputs(3759) <= not(layer0_outputs(3214));
    layer1_outputs(3760) <= '0';
    layer1_outputs(3761) <= not((layer0_outputs(1981)) xor (layer0_outputs(10973)));
    layer1_outputs(3762) <= layer0_outputs(11539);
    layer1_outputs(3763) <= layer0_outputs(10112);
    layer1_outputs(3764) <= (layer0_outputs(6391)) and not (layer0_outputs(11451));
    layer1_outputs(3765) <= not(layer0_outputs(6357));
    layer1_outputs(3766) <= not(layer0_outputs(11845));
    layer1_outputs(3767) <= not((layer0_outputs(2543)) or (layer0_outputs(11870)));
    layer1_outputs(3768) <= (layer0_outputs(3887)) and not (layer0_outputs(4835));
    layer1_outputs(3769) <= not(layer0_outputs(2008)) or (layer0_outputs(11904));
    layer1_outputs(3770) <= (layer0_outputs(10442)) and not (layer0_outputs(3760));
    layer1_outputs(3771) <= (layer0_outputs(2506)) and (layer0_outputs(8004));
    layer1_outputs(3772) <= (layer0_outputs(11962)) and not (layer0_outputs(5829));
    layer1_outputs(3773) <= (layer0_outputs(6958)) or (layer0_outputs(11459));
    layer1_outputs(3774) <= (layer0_outputs(94)) xor (layer0_outputs(992));
    layer1_outputs(3775) <= (layer0_outputs(3979)) xor (layer0_outputs(1980));
    layer1_outputs(3776) <= not(layer0_outputs(11141)) or (layer0_outputs(601));
    layer1_outputs(3777) <= layer0_outputs(7844);
    layer1_outputs(3778) <= (layer0_outputs(2)) and not (layer0_outputs(5379));
    layer1_outputs(3779) <= not((layer0_outputs(9643)) xor (layer0_outputs(6027)));
    layer1_outputs(3780) <= not(layer0_outputs(11111));
    layer1_outputs(3781) <= not(layer0_outputs(10656));
    layer1_outputs(3782) <= not(layer0_outputs(3173));
    layer1_outputs(3783) <= not(layer0_outputs(2856));
    layer1_outputs(3784) <= not(layer0_outputs(5605));
    layer1_outputs(3785) <= not(layer0_outputs(4535));
    layer1_outputs(3786) <= not((layer0_outputs(9253)) xor (layer0_outputs(387)));
    layer1_outputs(3787) <= not(layer0_outputs(10674)) or (layer0_outputs(1891));
    layer1_outputs(3788) <= layer0_outputs(5257);
    layer1_outputs(3789) <= not(layer0_outputs(6740));
    layer1_outputs(3790) <= layer0_outputs(6399);
    layer1_outputs(3791) <= (layer0_outputs(6188)) or (layer0_outputs(2918));
    layer1_outputs(3792) <= not(layer0_outputs(1038));
    layer1_outputs(3793) <= layer0_outputs(10791);
    layer1_outputs(3794) <= not(layer0_outputs(749)) or (layer0_outputs(7916));
    layer1_outputs(3795) <= layer0_outputs(8584);
    layer1_outputs(3796) <= (layer0_outputs(9744)) or (layer0_outputs(7409));
    layer1_outputs(3797) <= not((layer0_outputs(1080)) and (layer0_outputs(3463)));
    layer1_outputs(3798) <= '0';
    layer1_outputs(3799) <= (layer0_outputs(4800)) and (layer0_outputs(11963));
    layer1_outputs(3800) <= layer0_outputs(11737);
    layer1_outputs(3801) <= not(layer0_outputs(6444));
    layer1_outputs(3802) <= (layer0_outputs(519)) and not (layer0_outputs(1418));
    layer1_outputs(3803) <= layer0_outputs(4322);
    layer1_outputs(3804) <= '0';
    layer1_outputs(3805) <= (layer0_outputs(3155)) and not (layer0_outputs(4049));
    layer1_outputs(3806) <= layer0_outputs(4918);
    layer1_outputs(3807) <= not((layer0_outputs(1001)) xor (layer0_outputs(2384)));
    layer1_outputs(3808) <= layer0_outputs(1815);
    layer1_outputs(3809) <= not(layer0_outputs(3723));
    layer1_outputs(3810) <= not((layer0_outputs(9546)) and (layer0_outputs(1774)));
    layer1_outputs(3811) <= layer0_outputs(6638);
    layer1_outputs(3812) <= (layer0_outputs(7828)) or (layer0_outputs(10463));
    layer1_outputs(3813) <= (layer0_outputs(4640)) and not (layer0_outputs(5404));
    layer1_outputs(3814) <= layer0_outputs(9703);
    layer1_outputs(3815) <= not((layer0_outputs(2948)) and (layer0_outputs(1682)));
    layer1_outputs(3816) <= (layer0_outputs(7532)) and (layer0_outputs(5520));
    layer1_outputs(3817) <= layer0_outputs(9545);
    layer1_outputs(3818) <= not(layer0_outputs(12316));
    layer1_outputs(3819) <= not(layer0_outputs(12012));
    layer1_outputs(3820) <= not((layer0_outputs(3347)) or (layer0_outputs(11028)));
    layer1_outputs(3821) <= layer0_outputs(10045);
    layer1_outputs(3822) <= not(layer0_outputs(7809)) or (layer0_outputs(7344));
    layer1_outputs(3823) <= layer0_outputs(9302);
    layer1_outputs(3824) <= layer0_outputs(362);
    layer1_outputs(3825) <= not((layer0_outputs(7281)) or (layer0_outputs(9719)));
    layer1_outputs(3826) <= (layer0_outputs(300)) xor (layer0_outputs(9707));
    layer1_outputs(3827) <= not((layer0_outputs(2089)) xor (layer0_outputs(11912)));
    layer1_outputs(3828) <= not((layer0_outputs(7049)) and (layer0_outputs(860)));
    layer1_outputs(3829) <= (layer0_outputs(11334)) xor (layer0_outputs(3478));
    layer1_outputs(3830) <= not(layer0_outputs(7149));
    layer1_outputs(3831) <= not((layer0_outputs(10545)) xor (layer0_outputs(9033)));
    layer1_outputs(3832) <= not(layer0_outputs(4747)) or (layer0_outputs(7540));
    layer1_outputs(3833) <= not(layer0_outputs(1529));
    layer1_outputs(3834) <= not((layer0_outputs(8157)) and (layer0_outputs(10120)));
    layer1_outputs(3835) <= layer0_outputs(10246);
    layer1_outputs(3836) <= (layer0_outputs(12693)) and not (layer0_outputs(1525));
    layer1_outputs(3837) <= layer0_outputs(9730);
    layer1_outputs(3838) <= not((layer0_outputs(266)) and (layer0_outputs(8746)));
    layer1_outputs(3839) <= not(layer0_outputs(1318));
    layer1_outputs(3840) <= (layer0_outputs(11101)) or (layer0_outputs(12226));
    layer1_outputs(3841) <= not(layer0_outputs(12265)) or (layer0_outputs(9859));
    layer1_outputs(3842) <= (layer0_outputs(3044)) and not (layer0_outputs(2870));
    layer1_outputs(3843) <= layer0_outputs(826);
    layer1_outputs(3844) <= (layer0_outputs(10960)) and not (layer0_outputs(2171));
    layer1_outputs(3845) <= not(layer0_outputs(5712));
    layer1_outputs(3846) <= not((layer0_outputs(6420)) and (layer0_outputs(10021)));
    layer1_outputs(3847) <= layer0_outputs(6982);
    layer1_outputs(3848) <= (layer0_outputs(6971)) and (layer0_outputs(12431));
    layer1_outputs(3849) <= layer0_outputs(6607);
    layer1_outputs(3850) <= (layer0_outputs(4653)) and not (layer0_outputs(11146));
    layer1_outputs(3851) <= (layer0_outputs(2494)) and (layer0_outputs(4040));
    layer1_outputs(3852) <= (layer0_outputs(11506)) and (layer0_outputs(4942));
    layer1_outputs(3853) <= not(layer0_outputs(5445)) or (layer0_outputs(12663));
    layer1_outputs(3854) <= (layer0_outputs(642)) and not (layer0_outputs(10875));
    layer1_outputs(3855) <= (layer0_outputs(9049)) or (layer0_outputs(6702));
    layer1_outputs(3856) <= layer0_outputs(3481);
    layer1_outputs(3857) <= (layer0_outputs(449)) xor (layer0_outputs(4767));
    layer1_outputs(3858) <= not(layer0_outputs(10765));
    layer1_outputs(3859) <= (layer0_outputs(8212)) xor (layer0_outputs(1262));
    layer1_outputs(3860) <= layer0_outputs(12414);
    layer1_outputs(3861) <= not(layer0_outputs(3319)) or (layer0_outputs(3108));
    layer1_outputs(3862) <= not(layer0_outputs(4776)) or (layer0_outputs(8328));
    layer1_outputs(3863) <= not(layer0_outputs(3057));
    layer1_outputs(3864) <= layer0_outputs(8546);
    layer1_outputs(3865) <= not(layer0_outputs(3204)) or (layer0_outputs(11719));
    layer1_outputs(3866) <= not(layer0_outputs(1755));
    layer1_outputs(3867) <= (layer0_outputs(8609)) and not (layer0_outputs(4591));
    layer1_outputs(3868) <= (layer0_outputs(4456)) and (layer0_outputs(5895));
    layer1_outputs(3869) <= (layer0_outputs(11971)) and not (layer0_outputs(9868));
    layer1_outputs(3870) <= layer0_outputs(7098);
    layer1_outputs(3871) <= (layer0_outputs(12148)) xor (layer0_outputs(12719));
    layer1_outputs(3872) <= (layer0_outputs(12632)) and not (layer0_outputs(12420));
    layer1_outputs(3873) <= (layer0_outputs(582)) and (layer0_outputs(7884));
    layer1_outputs(3874) <= layer0_outputs(4108);
    layer1_outputs(3875) <= not((layer0_outputs(6624)) and (layer0_outputs(9506)));
    layer1_outputs(3876) <= not(layer0_outputs(8463));
    layer1_outputs(3877) <= layer0_outputs(12071);
    layer1_outputs(3878) <= not((layer0_outputs(1558)) xor (layer0_outputs(6969)));
    layer1_outputs(3879) <= (layer0_outputs(1742)) and not (layer0_outputs(8920));
    layer1_outputs(3880) <= '0';
    layer1_outputs(3881) <= not(layer0_outputs(7052));
    layer1_outputs(3882) <= not(layer0_outputs(10714));
    layer1_outputs(3883) <= not(layer0_outputs(11760));
    layer1_outputs(3884) <= not((layer0_outputs(5462)) and (layer0_outputs(10163)));
    layer1_outputs(3885) <= not(layer0_outputs(5287));
    layer1_outputs(3886) <= (layer0_outputs(4270)) and (layer0_outputs(4345));
    layer1_outputs(3887) <= not((layer0_outputs(2612)) and (layer0_outputs(11592)));
    layer1_outputs(3888) <= (layer0_outputs(2055)) and not (layer0_outputs(10649));
    layer1_outputs(3889) <= (layer0_outputs(9405)) or (layer0_outputs(5506));
    layer1_outputs(3890) <= not((layer0_outputs(5384)) xor (layer0_outputs(889)));
    layer1_outputs(3891) <= not((layer0_outputs(11035)) xor (layer0_outputs(780)));
    layer1_outputs(3892) <= not(layer0_outputs(964)) or (layer0_outputs(3134));
    layer1_outputs(3893) <= layer0_outputs(9595);
    layer1_outputs(3894) <= not(layer0_outputs(4704));
    layer1_outputs(3895) <= not(layer0_outputs(3535)) or (layer0_outputs(494));
    layer1_outputs(3896) <= not((layer0_outputs(8940)) xor (layer0_outputs(9115)));
    layer1_outputs(3897) <= not(layer0_outputs(1806));
    layer1_outputs(3898) <= (layer0_outputs(5268)) xor (layer0_outputs(1962));
    layer1_outputs(3899) <= not(layer0_outputs(1167));
    layer1_outputs(3900) <= (layer0_outputs(12117)) and not (layer0_outputs(12104));
    layer1_outputs(3901) <= layer0_outputs(814);
    layer1_outputs(3902) <= (layer0_outputs(3553)) and (layer0_outputs(2590));
    layer1_outputs(3903) <= not(layer0_outputs(8374));
    layer1_outputs(3904) <= (layer0_outputs(3839)) and not (layer0_outputs(2409));
    layer1_outputs(3905) <= not(layer0_outputs(10724)) or (layer0_outputs(9701));
    layer1_outputs(3906) <= not(layer0_outputs(5394)) or (layer0_outputs(6987));
    layer1_outputs(3907) <= (layer0_outputs(4103)) xor (layer0_outputs(11113));
    layer1_outputs(3908) <= layer0_outputs(3216);
    layer1_outputs(3909) <= not(layer0_outputs(4760));
    layer1_outputs(3910) <= not((layer0_outputs(12332)) or (layer0_outputs(2555)));
    layer1_outputs(3911) <= (layer0_outputs(2831)) or (layer0_outputs(5805));
    layer1_outputs(3912) <= not(layer0_outputs(9873)) or (layer0_outputs(9530));
    layer1_outputs(3913) <= (layer0_outputs(7121)) and (layer0_outputs(1958));
    layer1_outputs(3914) <= not(layer0_outputs(12612));
    layer1_outputs(3915) <= layer0_outputs(646);
    layer1_outputs(3916) <= (layer0_outputs(6299)) and not (layer0_outputs(7548));
    layer1_outputs(3917) <= (layer0_outputs(2148)) xor (layer0_outputs(804));
    layer1_outputs(3918) <= not((layer0_outputs(1736)) xor (layer0_outputs(10565)));
    layer1_outputs(3919) <= (layer0_outputs(12349)) xor (layer0_outputs(1627));
    layer1_outputs(3920) <= not(layer0_outputs(6100));
    layer1_outputs(3921) <= (layer0_outputs(2551)) or (layer0_outputs(7426));
    layer1_outputs(3922) <= not(layer0_outputs(4973));
    layer1_outputs(3923) <= not((layer0_outputs(545)) and (layer0_outputs(7274)));
    layer1_outputs(3924) <= not(layer0_outputs(160));
    layer1_outputs(3925) <= not((layer0_outputs(5984)) and (layer0_outputs(4430)));
    layer1_outputs(3926) <= not((layer0_outputs(10041)) xor (layer0_outputs(12586)));
    layer1_outputs(3927) <= (layer0_outputs(481)) and (layer0_outputs(10673));
    layer1_outputs(3928) <= not(layer0_outputs(7692));
    layer1_outputs(3929) <= not(layer0_outputs(1185));
    layer1_outputs(3930) <= not((layer0_outputs(5423)) and (layer0_outputs(8974)));
    layer1_outputs(3931) <= not((layer0_outputs(8760)) xor (layer0_outputs(8423)));
    layer1_outputs(3932) <= not(layer0_outputs(1658));
    layer1_outputs(3933) <= (layer0_outputs(3347)) and not (layer0_outputs(12183));
    layer1_outputs(3934) <= not((layer0_outputs(4937)) or (layer0_outputs(1836)));
    layer1_outputs(3935) <= not(layer0_outputs(12404));
    layer1_outputs(3936) <= (layer0_outputs(7394)) and not (layer0_outputs(7800));
    layer1_outputs(3937) <= layer0_outputs(9954);
    layer1_outputs(3938) <= '0';
    layer1_outputs(3939) <= (layer0_outputs(11296)) and (layer0_outputs(12035));
    layer1_outputs(3940) <= (layer0_outputs(2543)) or (layer0_outputs(9957));
    layer1_outputs(3941) <= not(layer0_outputs(484)) or (layer0_outputs(11041));
    layer1_outputs(3942) <= (layer0_outputs(4404)) and (layer0_outputs(3529));
    layer1_outputs(3943) <= not(layer0_outputs(3949));
    layer1_outputs(3944) <= not(layer0_outputs(283));
    layer1_outputs(3945) <= layer0_outputs(3035);
    layer1_outputs(3946) <= (layer0_outputs(1190)) and not (layer0_outputs(3840));
    layer1_outputs(3947) <= not((layer0_outputs(2333)) xor (layer0_outputs(6842)));
    layer1_outputs(3948) <= (layer0_outputs(324)) and not (layer0_outputs(5176));
    layer1_outputs(3949) <= not(layer0_outputs(6275)) or (layer0_outputs(9227));
    layer1_outputs(3950) <= (layer0_outputs(8569)) and not (layer0_outputs(3884));
    layer1_outputs(3951) <= (layer0_outputs(12789)) and not (layer0_outputs(6408));
    layer1_outputs(3952) <= (layer0_outputs(8203)) xor (layer0_outputs(3070));
    layer1_outputs(3953) <= not(layer0_outputs(7977));
    layer1_outputs(3954) <= (layer0_outputs(4902)) xor (layer0_outputs(6467));
    layer1_outputs(3955) <= (layer0_outputs(7039)) xor (layer0_outputs(1473));
    layer1_outputs(3956) <= not((layer0_outputs(914)) or (layer0_outputs(12283)));
    layer1_outputs(3957) <= (layer0_outputs(12245)) and not (layer0_outputs(5640));
    layer1_outputs(3958) <= layer0_outputs(1851);
    layer1_outputs(3959) <= not(layer0_outputs(7688));
    layer1_outputs(3960) <= (layer0_outputs(6360)) and not (layer0_outputs(7120));
    layer1_outputs(3961) <= (layer0_outputs(12535)) xor (layer0_outputs(12509));
    layer1_outputs(3962) <= not(layer0_outputs(6673));
    layer1_outputs(3963) <= not((layer0_outputs(1170)) or (layer0_outputs(12362)));
    layer1_outputs(3964) <= not(layer0_outputs(8478));
    layer1_outputs(3965) <= (layer0_outputs(6070)) and not (layer0_outputs(11344));
    layer1_outputs(3966) <= not((layer0_outputs(9323)) or (layer0_outputs(11244)));
    layer1_outputs(3967) <= not(layer0_outputs(6102)) or (layer0_outputs(5753));
    layer1_outputs(3968) <= not(layer0_outputs(7202));
    layer1_outputs(3969) <= layer0_outputs(4477);
    layer1_outputs(3970) <= not(layer0_outputs(9989)) or (layer0_outputs(11829));
    layer1_outputs(3971) <= layer0_outputs(10238);
    layer1_outputs(3972) <= (layer0_outputs(3621)) or (layer0_outputs(4417));
    layer1_outputs(3973) <= layer0_outputs(3763);
    layer1_outputs(3974) <= layer0_outputs(4025);
    layer1_outputs(3975) <= not(layer0_outputs(75));
    layer1_outputs(3976) <= (layer0_outputs(11910)) and not (layer0_outputs(1186));
    layer1_outputs(3977) <= not(layer0_outputs(3382)) or (layer0_outputs(7053));
    layer1_outputs(3978) <= '1';
    layer1_outputs(3979) <= not(layer0_outputs(10688));
    layer1_outputs(3980) <= (layer0_outputs(7012)) and not (layer0_outputs(3787));
    layer1_outputs(3981) <= not((layer0_outputs(1626)) or (layer0_outputs(5236)));
    layer1_outputs(3982) <= not((layer0_outputs(2158)) or (layer0_outputs(2572)));
    layer1_outputs(3983) <= '1';
    layer1_outputs(3984) <= not(layer0_outputs(2770)) or (layer0_outputs(12152));
    layer1_outputs(3985) <= not(layer0_outputs(2992));
    layer1_outputs(3986) <= layer0_outputs(6942);
    layer1_outputs(3987) <= '1';
    layer1_outputs(3988) <= layer0_outputs(6402);
    layer1_outputs(3989) <= not((layer0_outputs(3373)) and (layer0_outputs(7197)));
    layer1_outputs(3990) <= (layer0_outputs(10188)) or (layer0_outputs(7831));
    layer1_outputs(3991) <= not(layer0_outputs(11058)) or (layer0_outputs(4670));
    layer1_outputs(3992) <= not(layer0_outputs(3266)) or (layer0_outputs(753));
    layer1_outputs(3993) <= '0';
    layer1_outputs(3994) <= not(layer0_outputs(10596)) or (layer0_outputs(6724));
    layer1_outputs(3995) <= not(layer0_outputs(8603)) or (layer0_outputs(3335));
    layer1_outputs(3996) <= '0';
    layer1_outputs(3997) <= (layer0_outputs(7740)) and not (layer0_outputs(11751));
    layer1_outputs(3998) <= not((layer0_outputs(8579)) or (layer0_outputs(9672)));
    layer1_outputs(3999) <= layer0_outputs(4971);
    layer1_outputs(4000) <= layer0_outputs(6190);
    layer1_outputs(4001) <= not(layer0_outputs(12516));
    layer1_outputs(4002) <= (layer0_outputs(11559)) or (layer0_outputs(10576));
    layer1_outputs(4003) <= layer0_outputs(10097);
    layer1_outputs(4004) <= layer0_outputs(2053);
    layer1_outputs(4005) <= (layer0_outputs(12766)) or (layer0_outputs(208));
    layer1_outputs(4006) <= not((layer0_outputs(8886)) and (layer0_outputs(6287)));
    layer1_outputs(4007) <= not((layer0_outputs(681)) xor (layer0_outputs(2654)));
    layer1_outputs(4008) <= layer0_outputs(3137);
    layer1_outputs(4009) <= not(layer0_outputs(12164));
    layer1_outputs(4010) <= layer0_outputs(8651);
    layer1_outputs(4011) <= (layer0_outputs(627)) and not (layer0_outputs(8719));
    layer1_outputs(4012) <= not(layer0_outputs(1323));
    layer1_outputs(4013) <= not(layer0_outputs(769));
    layer1_outputs(4014) <= layer0_outputs(5925);
    layer1_outputs(4015) <= (layer0_outputs(12241)) and (layer0_outputs(12099));
    layer1_outputs(4016) <= (layer0_outputs(8364)) and (layer0_outputs(6410));
    layer1_outputs(4017) <= (layer0_outputs(7130)) and not (layer0_outputs(2235));
    layer1_outputs(4018) <= (layer0_outputs(9749)) and not (layer0_outputs(8453));
    layer1_outputs(4019) <= (layer0_outputs(9999)) or (layer0_outputs(10022));
    layer1_outputs(4020) <= not(layer0_outputs(8630));
    layer1_outputs(4021) <= layer0_outputs(5874);
    layer1_outputs(4022) <= (layer0_outputs(4893)) xor (layer0_outputs(12078));
    layer1_outputs(4023) <= not((layer0_outputs(970)) xor (layer0_outputs(3327)));
    layer1_outputs(4024) <= layer0_outputs(233);
    layer1_outputs(4025) <= not(layer0_outputs(3622));
    layer1_outputs(4026) <= (layer0_outputs(5828)) or (layer0_outputs(3588));
    layer1_outputs(4027) <= not((layer0_outputs(6779)) or (layer0_outputs(5044)));
    layer1_outputs(4028) <= not((layer0_outputs(3226)) and (layer0_outputs(818)));
    layer1_outputs(4029) <= not(layer0_outputs(11641)) or (layer0_outputs(8193));
    layer1_outputs(4030) <= layer0_outputs(5084);
    layer1_outputs(4031) <= not(layer0_outputs(5992)) or (layer0_outputs(2946));
    layer1_outputs(4032) <= not(layer0_outputs(2097));
    layer1_outputs(4033) <= not((layer0_outputs(4628)) and (layer0_outputs(5930)));
    layer1_outputs(4034) <= not(layer0_outputs(7955));
    layer1_outputs(4035) <= not(layer0_outputs(8652));
    layer1_outputs(4036) <= not(layer0_outputs(3025));
    layer1_outputs(4037) <= not((layer0_outputs(7608)) and (layer0_outputs(1287)));
    layer1_outputs(4038) <= layer0_outputs(5488);
    layer1_outputs(4039) <= (layer0_outputs(7822)) or (layer0_outputs(6940));
    layer1_outputs(4040) <= layer0_outputs(7445);
    layer1_outputs(4041) <= layer0_outputs(12603);
    layer1_outputs(4042) <= not(layer0_outputs(12451));
    layer1_outputs(4043) <= layer0_outputs(6418);
    layer1_outputs(4044) <= not(layer0_outputs(6220)) or (layer0_outputs(7863));
    layer1_outputs(4045) <= (layer0_outputs(8851)) xor (layer0_outputs(9014));
    layer1_outputs(4046) <= not(layer0_outputs(4065));
    layer1_outputs(4047) <= not(layer0_outputs(7311));
    layer1_outputs(4048) <= (layer0_outputs(9699)) xor (layer0_outputs(10519));
    layer1_outputs(4049) <= (layer0_outputs(9026)) and not (layer0_outputs(290));
    layer1_outputs(4050) <= not((layer0_outputs(7052)) and (layer0_outputs(7856)));
    layer1_outputs(4051) <= not(layer0_outputs(1625)) or (layer0_outputs(2421));
    layer1_outputs(4052) <= (layer0_outputs(3595)) and not (layer0_outputs(6765));
    layer1_outputs(4053) <= layer0_outputs(3643);
    layer1_outputs(4054) <= not((layer0_outputs(2807)) and (layer0_outputs(1764)));
    layer1_outputs(4055) <= (layer0_outputs(97)) and (layer0_outputs(4752));
    layer1_outputs(4056) <= not(layer0_outputs(3367));
    layer1_outputs(4057) <= layer0_outputs(16);
    layer1_outputs(4058) <= not(layer0_outputs(9026));
    layer1_outputs(4059) <= not((layer0_outputs(5844)) or (layer0_outputs(12163)));
    layer1_outputs(4060) <= not(layer0_outputs(896));
    layer1_outputs(4061) <= layer0_outputs(7877);
    layer1_outputs(4062) <= layer0_outputs(10666);
    layer1_outputs(4063) <= not(layer0_outputs(8990));
    layer1_outputs(4064) <= not((layer0_outputs(6952)) and (layer0_outputs(5598)));
    layer1_outputs(4065) <= (layer0_outputs(5839)) xor (layer0_outputs(2527));
    layer1_outputs(4066) <= (layer0_outputs(8733)) or (layer0_outputs(967));
    layer1_outputs(4067) <= not(layer0_outputs(10471));
    layer1_outputs(4068) <= not(layer0_outputs(1494));
    layer1_outputs(4069) <= not(layer0_outputs(6450));
    layer1_outputs(4070) <= (layer0_outputs(4606)) and (layer0_outputs(11524));
    layer1_outputs(4071) <= not(layer0_outputs(11354));
    layer1_outputs(4072) <= '0';
    layer1_outputs(4073) <= not(layer0_outputs(4419));
    layer1_outputs(4074) <= (layer0_outputs(10560)) and not (layer0_outputs(6634));
    layer1_outputs(4075) <= not(layer0_outputs(355));
    layer1_outputs(4076) <= not((layer0_outputs(6823)) or (layer0_outputs(9415)));
    layer1_outputs(4077) <= layer0_outputs(8643);
    layer1_outputs(4078) <= not(layer0_outputs(521)) or (layer0_outputs(3514));
    layer1_outputs(4079) <= '0';
    layer1_outputs(4080) <= layer0_outputs(5175);
    layer1_outputs(4081) <= (layer0_outputs(10833)) and not (layer0_outputs(5776));
    layer1_outputs(4082) <= not((layer0_outputs(8187)) xor (layer0_outputs(1524)));
    layer1_outputs(4083) <= layer0_outputs(1801);
    layer1_outputs(4084) <= layer0_outputs(503);
    layer1_outputs(4085) <= (layer0_outputs(1615)) or (layer0_outputs(8090));
    layer1_outputs(4086) <= '1';
    layer1_outputs(4087) <= layer0_outputs(10866);
    layer1_outputs(4088) <= not(layer0_outputs(710));
    layer1_outputs(4089) <= (layer0_outputs(12459)) and (layer0_outputs(8757));
    layer1_outputs(4090) <= layer0_outputs(5443);
    layer1_outputs(4091) <= (layer0_outputs(11612)) or (layer0_outputs(4657));
    layer1_outputs(4092) <= layer0_outputs(82);
    layer1_outputs(4093) <= not(layer0_outputs(8291)) or (layer0_outputs(5991));
    layer1_outputs(4094) <= (layer0_outputs(1737)) and not (layer0_outputs(4165));
    layer1_outputs(4095) <= not((layer0_outputs(3524)) or (layer0_outputs(5410)));
    layer1_outputs(4096) <= (layer0_outputs(11971)) xor (layer0_outputs(6737));
    layer1_outputs(4097) <= not(layer0_outputs(4536));
    layer1_outputs(4098) <= (layer0_outputs(365)) and not (layer0_outputs(12165));
    layer1_outputs(4099) <= not(layer0_outputs(9439));
    layer1_outputs(4100) <= (layer0_outputs(2511)) and (layer0_outputs(6308));
    layer1_outputs(4101) <= (layer0_outputs(2751)) and not (layer0_outputs(5031));
    layer1_outputs(4102) <= not(layer0_outputs(4030));
    layer1_outputs(4103) <= layer0_outputs(2138);
    layer1_outputs(4104) <= layer0_outputs(10965);
    layer1_outputs(4105) <= not(layer0_outputs(4036)) or (layer0_outputs(2596));
    layer1_outputs(4106) <= not(layer0_outputs(4222)) or (layer0_outputs(6832));
    layer1_outputs(4107) <= not(layer0_outputs(7860)) or (layer0_outputs(2312));
    layer1_outputs(4108) <= not(layer0_outputs(11260));
    layer1_outputs(4109) <= (layer0_outputs(5679)) and (layer0_outputs(11821));
    layer1_outputs(4110) <= not((layer0_outputs(5483)) and (layer0_outputs(9267)));
    layer1_outputs(4111) <= layer0_outputs(8877);
    layer1_outputs(4112) <= not((layer0_outputs(10309)) or (layer0_outputs(8503)));
    layer1_outputs(4113) <= (layer0_outputs(8422)) and (layer0_outputs(8651));
    layer1_outputs(4114) <= not((layer0_outputs(12469)) or (layer0_outputs(11773)));
    layer1_outputs(4115) <= '1';
    layer1_outputs(4116) <= (layer0_outputs(907)) and not (layer0_outputs(4254));
    layer1_outputs(4117) <= layer0_outputs(679);
    layer1_outputs(4118) <= not(layer0_outputs(2003));
    layer1_outputs(4119) <= layer0_outputs(1671);
    layer1_outputs(4120) <= layer0_outputs(408);
    layer1_outputs(4121) <= not((layer0_outputs(4602)) and (layer0_outputs(4967)));
    layer1_outputs(4122) <= '0';
    layer1_outputs(4123) <= (layer0_outputs(11886)) and not (layer0_outputs(9886));
    layer1_outputs(4124) <= not(layer0_outputs(5612)) or (layer0_outputs(10002));
    layer1_outputs(4125) <= (layer0_outputs(51)) and not (layer0_outputs(10365));
    layer1_outputs(4126) <= layer0_outputs(617);
    layer1_outputs(4127) <= not(layer0_outputs(3011)) or (layer0_outputs(2945));
    layer1_outputs(4128) <= layer0_outputs(9396);
    layer1_outputs(4129) <= (layer0_outputs(11165)) and not (layer0_outputs(12088));
    layer1_outputs(4130) <= not(layer0_outputs(4730));
    layer1_outputs(4131) <= not(layer0_outputs(12217)) or (layer0_outputs(5037));
    layer1_outputs(4132) <= (layer0_outputs(6006)) and (layer0_outputs(12379));
    layer1_outputs(4133) <= not((layer0_outputs(11434)) xor (layer0_outputs(8769)));
    layer1_outputs(4134) <= (layer0_outputs(11415)) and not (layer0_outputs(2338));
    layer1_outputs(4135) <= (layer0_outputs(4312)) and (layer0_outputs(5011));
    layer1_outputs(4136) <= not(layer0_outputs(10225)) or (layer0_outputs(2973));
    layer1_outputs(4137) <= (layer0_outputs(227)) and (layer0_outputs(4779));
    layer1_outputs(4138) <= layer0_outputs(106);
    layer1_outputs(4139) <= (layer0_outputs(193)) xor (layer0_outputs(5154));
    layer1_outputs(4140) <= layer0_outputs(5302);
    layer1_outputs(4141) <= not((layer0_outputs(10081)) xor (layer0_outputs(5832)));
    layer1_outputs(4142) <= not(layer0_outputs(942));
    layer1_outputs(4143) <= (layer0_outputs(8518)) and not (layer0_outputs(8764));
    layer1_outputs(4144) <= '0';
    layer1_outputs(4145) <= layer0_outputs(9368);
    layer1_outputs(4146) <= not(layer0_outputs(11172)) or (layer0_outputs(6517));
    layer1_outputs(4147) <= not(layer0_outputs(1687));
    layer1_outputs(4148) <= layer0_outputs(12075);
    layer1_outputs(4149) <= layer0_outputs(2166);
    layer1_outputs(4150) <= '1';
    layer1_outputs(4151) <= (layer0_outputs(5029)) xor (layer0_outputs(10686));
    layer1_outputs(4152) <= layer0_outputs(11945);
    layer1_outputs(4153) <= not(layer0_outputs(1292));
    layer1_outputs(4154) <= not((layer0_outputs(644)) xor (layer0_outputs(10915)));
    layer1_outputs(4155) <= not((layer0_outputs(12242)) or (layer0_outputs(5774)));
    layer1_outputs(4156) <= not(layer0_outputs(10247)) or (layer0_outputs(4988));
    layer1_outputs(4157) <= not(layer0_outputs(6238));
    layer1_outputs(4158) <= not((layer0_outputs(2390)) and (layer0_outputs(4106)));
    layer1_outputs(4159) <= not((layer0_outputs(8979)) and (layer0_outputs(812)));
    layer1_outputs(4160) <= not((layer0_outputs(2802)) or (layer0_outputs(4234)));
    layer1_outputs(4161) <= (layer0_outputs(12569)) or (layer0_outputs(11390));
    layer1_outputs(4162) <= not((layer0_outputs(276)) xor (layer0_outputs(5677)));
    layer1_outputs(4163) <= not(layer0_outputs(10124));
    layer1_outputs(4164) <= not((layer0_outputs(5690)) and (layer0_outputs(3346)));
    layer1_outputs(4165) <= not(layer0_outputs(5853)) or (layer0_outputs(9428));
    layer1_outputs(4166) <= not(layer0_outputs(7699));
    layer1_outputs(4167) <= (layer0_outputs(8785)) and (layer0_outputs(10354));
    layer1_outputs(4168) <= (layer0_outputs(12579)) and not (layer0_outputs(7412));
    layer1_outputs(4169) <= layer0_outputs(6595);
    layer1_outputs(4170) <= (layer0_outputs(11153)) or (layer0_outputs(6609));
    layer1_outputs(4171) <= not(layer0_outputs(974));
    layer1_outputs(4172) <= not(layer0_outputs(6526));
    layer1_outputs(4173) <= (layer0_outputs(5956)) or (layer0_outputs(11247));
    layer1_outputs(4174) <= layer0_outputs(7524);
    layer1_outputs(4175) <= not(layer0_outputs(3663));
    layer1_outputs(4176) <= not(layer0_outputs(4918));
    layer1_outputs(4177) <= (layer0_outputs(646)) and (layer0_outputs(4232));
    layer1_outputs(4178) <= not(layer0_outputs(4225));
    layer1_outputs(4179) <= not(layer0_outputs(12728));
    layer1_outputs(4180) <= (layer0_outputs(1629)) and not (layer0_outputs(4348));
    layer1_outputs(4181) <= not(layer0_outputs(9467)) or (layer0_outputs(4067));
    layer1_outputs(4182) <= layer0_outputs(7576);
    layer1_outputs(4183) <= layer0_outputs(7975);
    layer1_outputs(4184) <= not((layer0_outputs(5873)) and (layer0_outputs(0)));
    layer1_outputs(4185) <= not(layer0_outputs(865));
    layer1_outputs(4186) <= not(layer0_outputs(159));
    layer1_outputs(4187) <= (layer0_outputs(12232)) and not (layer0_outputs(5496));
    layer1_outputs(4188) <= (layer0_outputs(11089)) and not (layer0_outputs(12013));
    layer1_outputs(4189) <= not((layer0_outputs(9739)) and (layer0_outputs(6836)));
    layer1_outputs(4190) <= (layer0_outputs(7774)) or (layer0_outputs(7759));
    layer1_outputs(4191) <= (layer0_outputs(7613)) xor (layer0_outputs(517));
    layer1_outputs(4192) <= not(layer0_outputs(10252)) or (layer0_outputs(2104));
    layer1_outputs(4193) <= (layer0_outputs(1656)) or (layer0_outputs(8154));
    layer1_outputs(4194) <= not(layer0_outputs(3247));
    layer1_outputs(4195) <= layer0_outputs(12032);
    layer1_outputs(4196) <= '0';
    layer1_outputs(4197) <= layer0_outputs(2336);
    layer1_outputs(4198) <= (layer0_outputs(8457)) and (layer0_outputs(5658));
    layer1_outputs(4199) <= not(layer0_outputs(12748));
    layer1_outputs(4200) <= layer0_outputs(6092);
    layer1_outputs(4201) <= (layer0_outputs(11600)) or (layer0_outputs(9113));
    layer1_outputs(4202) <= not(layer0_outputs(3338)) or (layer0_outputs(2764));
    layer1_outputs(4203) <= layer0_outputs(3717);
    layer1_outputs(4204) <= (layer0_outputs(10631)) or (layer0_outputs(4738));
    layer1_outputs(4205) <= (layer0_outputs(5024)) and not (layer0_outputs(9967));
    layer1_outputs(4206) <= (layer0_outputs(2038)) and (layer0_outputs(792));
    layer1_outputs(4207) <= '0';
    layer1_outputs(4208) <= (layer0_outputs(6141)) and not (layer0_outputs(11960));
    layer1_outputs(4209) <= (layer0_outputs(1239)) xor (layer0_outputs(12137));
    layer1_outputs(4210) <= not((layer0_outputs(2416)) and (layer0_outputs(8584)));
    layer1_outputs(4211) <= not(layer0_outputs(2284)) or (layer0_outputs(11892));
    layer1_outputs(4212) <= (layer0_outputs(6239)) or (layer0_outputs(3053));
    layer1_outputs(4213) <= not((layer0_outputs(9085)) xor (layer0_outputs(6453)));
    layer1_outputs(4214) <= layer0_outputs(1069);
    layer1_outputs(4215) <= (layer0_outputs(6795)) and not (layer0_outputs(7641));
    layer1_outputs(4216) <= layer0_outputs(8072);
    layer1_outputs(4217) <= not((layer0_outputs(5846)) xor (layer0_outputs(11951)));
    layer1_outputs(4218) <= layer0_outputs(11171);
    layer1_outputs(4219) <= (layer0_outputs(12554)) and not (layer0_outputs(6949));
    layer1_outputs(4220) <= not(layer0_outputs(5735));
    layer1_outputs(4221) <= layer0_outputs(11597);
    layer1_outputs(4222) <= not(layer0_outputs(11747));
    layer1_outputs(4223) <= not(layer0_outputs(757));
    layer1_outputs(4224) <= not(layer0_outputs(11500));
    layer1_outputs(4225) <= (layer0_outputs(8671)) and not (layer0_outputs(12021));
    layer1_outputs(4226) <= not((layer0_outputs(4815)) or (layer0_outputs(9164)));
    layer1_outputs(4227) <= (layer0_outputs(2678)) and not (layer0_outputs(1850));
    layer1_outputs(4228) <= not(layer0_outputs(11604));
    layer1_outputs(4229) <= layer0_outputs(3060);
    layer1_outputs(4230) <= (layer0_outputs(5648)) or (layer0_outputs(6121));
    layer1_outputs(4231) <= not(layer0_outputs(10539));
    layer1_outputs(4232) <= not((layer0_outputs(3982)) or (layer0_outputs(357)));
    layer1_outputs(4233) <= (layer0_outputs(3495)) and (layer0_outputs(3794));
    layer1_outputs(4234) <= not(layer0_outputs(7071));
    layer1_outputs(4235) <= layer0_outputs(3459);
    layer1_outputs(4236) <= not(layer0_outputs(8661));
    layer1_outputs(4237) <= not(layer0_outputs(2070)) or (layer0_outputs(1186));
    layer1_outputs(4238) <= layer0_outputs(1029);
    layer1_outputs(4239) <= not(layer0_outputs(2695)) or (layer0_outputs(8714));
    layer1_outputs(4240) <= (layer0_outputs(9556)) xor (layer0_outputs(12540));
    layer1_outputs(4241) <= not((layer0_outputs(4224)) xor (layer0_outputs(12597)));
    layer1_outputs(4242) <= not((layer0_outputs(3721)) and (layer0_outputs(7864)));
    layer1_outputs(4243) <= not(layer0_outputs(11757));
    layer1_outputs(4244) <= (layer0_outputs(12437)) and not (layer0_outputs(6824));
    layer1_outputs(4245) <= (layer0_outputs(6572)) and not (layer0_outputs(2488));
    layer1_outputs(4246) <= '0';
    layer1_outputs(4247) <= not((layer0_outputs(11121)) xor (layer0_outputs(5845)));
    layer1_outputs(4248) <= not(layer0_outputs(1819)) or (layer0_outputs(1924));
    layer1_outputs(4249) <= not((layer0_outputs(9684)) and (layer0_outputs(1376)));
    layer1_outputs(4250) <= layer0_outputs(2881);
    layer1_outputs(4251) <= not(layer0_outputs(7902));
    layer1_outputs(4252) <= (layer0_outputs(5201)) and (layer0_outputs(2699));
    layer1_outputs(4253) <= not(layer0_outputs(3708));
    layer1_outputs(4254) <= not(layer0_outputs(2625));
    layer1_outputs(4255) <= not(layer0_outputs(9635));
    layer1_outputs(4256) <= (layer0_outputs(12778)) or (layer0_outputs(8539));
    layer1_outputs(4257) <= not((layer0_outputs(2001)) and (layer0_outputs(317)));
    layer1_outputs(4258) <= layer0_outputs(3687);
    layer1_outputs(4259) <= not((layer0_outputs(2840)) and (layer0_outputs(2977)));
    layer1_outputs(4260) <= layer0_outputs(1897);
    layer1_outputs(4261) <= not(layer0_outputs(4883));
    layer1_outputs(4262) <= not((layer0_outputs(11555)) and (layer0_outputs(5210)));
    layer1_outputs(4263) <= (layer0_outputs(9057)) and not (layer0_outputs(9202));
    layer1_outputs(4264) <= not(layer0_outputs(4782));
    layer1_outputs(4265) <= not((layer0_outputs(5306)) or (layer0_outputs(11308)));
    layer1_outputs(4266) <= not(layer0_outputs(11769));
    layer1_outputs(4267) <= not((layer0_outputs(10211)) xor (layer0_outputs(10003)));
    layer1_outputs(4268) <= (layer0_outputs(6817)) and not (layer0_outputs(7234));
    layer1_outputs(4269) <= (layer0_outputs(11033)) or (layer0_outputs(8222));
    layer1_outputs(4270) <= not(layer0_outputs(155)) or (layer0_outputs(607));
    layer1_outputs(4271) <= not(layer0_outputs(7625));
    layer1_outputs(4272) <= not(layer0_outputs(10280));
    layer1_outputs(4273) <= not(layer0_outputs(4343));
    layer1_outputs(4274) <= not((layer0_outputs(6069)) and (layer0_outputs(7446)));
    layer1_outputs(4275) <= (layer0_outputs(9915)) and not (layer0_outputs(8890));
    layer1_outputs(4276) <= not((layer0_outputs(2376)) xor (layer0_outputs(4541)));
    layer1_outputs(4277) <= (layer0_outputs(10265)) and not (layer0_outputs(9053));
    layer1_outputs(4278) <= layer0_outputs(7812);
    layer1_outputs(4279) <= layer0_outputs(2786);
    layer1_outputs(4280) <= not(layer0_outputs(7355));
    layer1_outputs(4281) <= layer0_outputs(1716);
    layer1_outputs(4282) <= layer0_outputs(11109);
    layer1_outputs(4283) <= layer0_outputs(6655);
    layer1_outputs(4284) <= (layer0_outputs(3493)) or (layer0_outputs(5668));
    layer1_outputs(4285) <= layer0_outputs(2939);
    layer1_outputs(4286) <= not(layer0_outputs(6161));
    layer1_outputs(4287) <= (layer0_outputs(5405)) xor (layer0_outputs(1459));
    layer1_outputs(4288) <= not(layer0_outputs(6393));
    layer1_outputs(4289) <= not(layer0_outputs(10391));
    layer1_outputs(4290) <= not((layer0_outputs(6384)) xor (layer0_outputs(708)));
    layer1_outputs(4291) <= not(layer0_outputs(7717));
    layer1_outputs(4292) <= not((layer0_outputs(5988)) and (layer0_outputs(8029)));
    layer1_outputs(4293) <= not(layer0_outputs(8265));
    layer1_outputs(4294) <= layer0_outputs(6362);
    layer1_outputs(4295) <= not(layer0_outputs(2175));
    layer1_outputs(4296) <= not(layer0_outputs(11228));
    layer1_outputs(4297) <= not((layer0_outputs(10838)) xor (layer0_outputs(5135)));
    layer1_outputs(4298) <= (layer0_outputs(5245)) xor (layer0_outputs(5663));
    layer1_outputs(4299) <= (layer0_outputs(6082)) and not (layer0_outputs(1046));
    layer1_outputs(4300) <= not((layer0_outputs(5712)) or (layer0_outputs(10179)));
    layer1_outputs(4301) <= layer0_outputs(7485);
    layer1_outputs(4302) <= (layer0_outputs(2972)) or (layer0_outputs(7516));
    layer1_outputs(4303) <= not(layer0_outputs(6676));
    layer1_outputs(4304) <= (layer0_outputs(10684)) or (layer0_outputs(11634));
    layer1_outputs(4305) <= (layer0_outputs(11426)) and not (layer0_outputs(4081));
    layer1_outputs(4306) <= not((layer0_outputs(11711)) or (layer0_outputs(11763)));
    layer1_outputs(4307) <= (layer0_outputs(12420)) xor (layer0_outputs(10420));
    layer1_outputs(4308) <= layer0_outputs(4447);
    layer1_outputs(4309) <= not(layer0_outputs(5232)) or (layer0_outputs(10037));
    layer1_outputs(4310) <= not(layer0_outputs(10936));
    layer1_outputs(4311) <= (layer0_outputs(11664)) xor (layer0_outputs(7250));
    layer1_outputs(4312) <= not(layer0_outputs(12593)) or (layer0_outputs(4554));
    layer1_outputs(4313) <= (layer0_outputs(9897)) xor (layer0_outputs(9286));
    layer1_outputs(4314) <= not((layer0_outputs(2493)) xor (layer0_outputs(6837)));
    layer1_outputs(4315) <= not(layer0_outputs(5149));
    layer1_outputs(4316) <= not((layer0_outputs(9247)) xor (layer0_outputs(8391)));
    layer1_outputs(4317) <= layer0_outputs(8301);
    layer1_outputs(4318) <= not(layer0_outputs(12657)) or (layer0_outputs(4391));
    layer1_outputs(4319) <= layer0_outputs(3462);
    layer1_outputs(4320) <= not((layer0_outputs(11425)) xor (layer0_outputs(4172)));
    layer1_outputs(4321) <= not((layer0_outputs(900)) or (layer0_outputs(10423)));
    layer1_outputs(4322) <= '1';
    layer1_outputs(4323) <= not(layer0_outputs(6220)) or (layer0_outputs(8738));
    layer1_outputs(4324) <= not(layer0_outputs(10793));
    layer1_outputs(4325) <= not((layer0_outputs(6135)) or (layer0_outputs(9652)));
    layer1_outputs(4326) <= layer0_outputs(4936);
    layer1_outputs(4327) <= not(layer0_outputs(10490)) or (layer0_outputs(11835));
    layer1_outputs(4328) <= (layer0_outputs(3931)) and (layer0_outputs(3100));
    layer1_outputs(4329) <= layer0_outputs(12430);
    layer1_outputs(4330) <= (layer0_outputs(10993)) and (layer0_outputs(9877));
    layer1_outputs(4331) <= layer0_outputs(5121);
    layer1_outputs(4332) <= not((layer0_outputs(6193)) and (layer0_outputs(7390)));
    layer1_outputs(4333) <= layer0_outputs(3606);
    layer1_outputs(4334) <= not((layer0_outputs(4736)) and (layer0_outputs(1219)));
    layer1_outputs(4335) <= not((layer0_outputs(3610)) xor (layer0_outputs(4943)));
    layer1_outputs(4336) <= not(layer0_outputs(5759));
    layer1_outputs(4337) <= not(layer0_outputs(5866));
    layer1_outputs(4338) <= (layer0_outputs(7379)) and (layer0_outputs(5005));
    layer1_outputs(4339) <= (layer0_outputs(6173)) xor (layer0_outputs(5969));
    layer1_outputs(4340) <= not(layer0_outputs(3675)) or (layer0_outputs(1771));
    layer1_outputs(4341) <= layer0_outputs(11814);
    layer1_outputs(4342) <= (layer0_outputs(60)) or (layer0_outputs(6552));
    layer1_outputs(4343) <= (layer0_outputs(12525)) and not (layer0_outputs(4198));
    layer1_outputs(4344) <= not(layer0_outputs(238)) or (layer0_outputs(1181));
    layer1_outputs(4345) <= not((layer0_outputs(2470)) or (layer0_outputs(3251)));
    layer1_outputs(4346) <= not(layer0_outputs(12779));
    layer1_outputs(4347) <= not(layer0_outputs(917));
    layer1_outputs(4348) <= not((layer0_outputs(12031)) or (layer0_outputs(11283)));
    layer1_outputs(4349) <= '0';
    layer1_outputs(4350) <= (layer0_outputs(2170)) and (layer0_outputs(8525));
    layer1_outputs(4351) <= layer0_outputs(9792);
    layer1_outputs(4352) <= not((layer0_outputs(5470)) xor (layer0_outputs(3019)));
    layer1_outputs(4353) <= not(layer0_outputs(8175)) or (layer0_outputs(6521));
    layer1_outputs(4354) <= not(layer0_outputs(9862));
    layer1_outputs(4355) <= (layer0_outputs(5687)) and not (layer0_outputs(1886));
    layer1_outputs(4356) <= not(layer0_outputs(4689)) or (layer0_outputs(5474));
    layer1_outputs(4357) <= '1';
    layer1_outputs(4358) <= not(layer0_outputs(960));
    layer1_outputs(4359) <= layer0_outputs(3878);
    layer1_outputs(4360) <= (layer0_outputs(12625)) and not (layer0_outputs(7324));
    layer1_outputs(4361) <= layer0_outputs(10584);
    layer1_outputs(4362) <= not((layer0_outputs(11775)) and (layer0_outputs(10581)));
    layer1_outputs(4363) <= (layer0_outputs(7998)) or (layer0_outputs(10932));
    layer1_outputs(4364) <= layer0_outputs(5630);
    layer1_outputs(4365) <= '0';
    layer1_outputs(4366) <= not((layer0_outputs(7568)) and (layer0_outputs(12751)));
    layer1_outputs(4367) <= not((layer0_outputs(5456)) or (layer0_outputs(5103)));
    layer1_outputs(4368) <= (layer0_outputs(11301)) and (layer0_outputs(5980));
    layer1_outputs(4369) <= (layer0_outputs(9504)) and not (layer0_outputs(12626));
    layer1_outputs(4370) <= layer0_outputs(3739);
    layer1_outputs(4371) <= not((layer0_outputs(4150)) xor (layer0_outputs(12084)));
    layer1_outputs(4372) <= not(layer0_outputs(6235));
    layer1_outputs(4373) <= layer0_outputs(2202);
    layer1_outputs(4374) <= not((layer0_outputs(10629)) or (layer0_outputs(9311)));
    layer1_outputs(4375) <= not(layer0_outputs(11466));
    layer1_outputs(4376) <= not(layer0_outputs(11342));
    layer1_outputs(4377) <= not(layer0_outputs(9298));
    layer1_outputs(4378) <= not((layer0_outputs(10996)) and (layer0_outputs(11640)));
    layer1_outputs(4379) <= not(layer0_outputs(11556));
    layer1_outputs(4380) <= not(layer0_outputs(5086));
    layer1_outputs(4381) <= not((layer0_outputs(1275)) and (layer0_outputs(10920)));
    layer1_outputs(4382) <= not(layer0_outputs(12089)) or (layer0_outputs(5052));
    layer1_outputs(4383) <= not((layer0_outputs(1760)) xor (layer0_outputs(12675)));
    layer1_outputs(4384) <= (layer0_outputs(597)) and not (layer0_outputs(6335));
    layer1_outputs(4385) <= layer0_outputs(9391);
    layer1_outputs(4386) <= not(layer0_outputs(7070)) or (layer0_outputs(7089));
    layer1_outputs(4387) <= layer0_outputs(894);
    layer1_outputs(4388) <= not((layer0_outputs(5908)) and (layer0_outputs(1743)));
    layer1_outputs(4389) <= not(layer0_outputs(5105));
    layer1_outputs(4390) <= not(layer0_outputs(9353));
    layer1_outputs(4391) <= not((layer0_outputs(7767)) or (layer0_outputs(9094)));
    layer1_outputs(4392) <= not(layer0_outputs(10056));
    layer1_outputs(4393) <= not(layer0_outputs(77)) or (layer0_outputs(5714));
    layer1_outputs(4394) <= '1';
    layer1_outputs(4395) <= layer0_outputs(2628);
    layer1_outputs(4396) <= (layer0_outputs(1121)) xor (layer0_outputs(12330));
    layer1_outputs(4397) <= layer0_outputs(2554);
    layer1_outputs(4398) <= layer0_outputs(5922);
    layer1_outputs(4399) <= not(layer0_outputs(11739));
    layer1_outputs(4400) <= layer0_outputs(3749);
    layer1_outputs(4401) <= layer0_outputs(12570);
    layer1_outputs(4402) <= (layer0_outputs(10675)) and not (layer0_outputs(1384));
    layer1_outputs(4403) <= not((layer0_outputs(9400)) or (layer0_outputs(9957)));
    layer1_outputs(4404) <= (layer0_outputs(6213)) xor (layer0_outputs(9042));
    layer1_outputs(4405) <= not((layer0_outputs(5202)) and (layer0_outputs(5594)));
    layer1_outputs(4406) <= layer0_outputs(9631);
    layer1_outputs(4407) <= layer0_outputs(10114);
    layer1_outputs(4408) <= not(layer0_outputs(2473));
    layer1_outputs(4409) <= layer0_outputs(11317);
    layer1_outputs(4410) <= layer0_outputs(3936);
    layer1_outputs(4411) <= not((layer0_outputs(9044)) or (layer0_outputs(7747)));
    layer1_outputs(4412) <= layer0_outputs(3976);
    layer1_outputs(4413) <= layer0_outputs(8399);
    layer1_outputs(4414) <= (layer0_outputs(4050)) and not (layer0_outputs(748));
    layer1_outputs(4415) <= not((layer0_outputs(8373)) xor (layer0_outputs(11167)));
    layer1_outputs(4416) <= not(layer0_outputs(10330));
    layer1_outputs(4417) <= not(layer0_outputs(4532));
    layer1_outputs(4418) <= not(layer0_outputs(11048));
    layer1_outputs(4419) <= layer0_outputs(5726);
    layer1_outputs(4420) <= layer0_outputs(8177);
    layer1_outputs(4421) <= (layer0_outputs(10860)) and not (layer0_outputs(8902));
    layer1_outputs(4422) <= not(layer0_outputs(6051)) or (layer0_outputs(10053));
    layer1_outputs(4423) <= not(layer0_outputs(7016)) or (layer0_outputs(12530));
    layer1_outputs(4424) <= layer0_outputs(4584);
    layer1_outputs(4425) <= not(layer0_outputs(9090)) or (layer0_outputs(1429));
    layer1_outputs(4426) <= (layer0_outputs(7444)) and not (layer0_outputs(4103));
    layer1_outputs(4427) <= not(layer0_outputs(4892)) or (layer0_outputs(7865));
    layer1_outputs(4428) <= not((layer0_outputs(10717)) or (layer0_outputs(9081)));
    layer1_outputs(4429) <= layer0_outputs(2693);
    layer1_outputs(4430) <= not((layer0_outputs(6041)) and (layer0_outputs(11100)));
    layer1_outputs(4431) <= (layer0_outputs(10346)) xor (layer0_outputs(6854));
    layer1_outputs(4432) <= (layer0_outputs(8694)) xor (layer0_outputs(6715));
    layer1_outputs(4433) <= layer0_outputs(3914);
    layer1_outputs(4434) <= layer0_outputs(2253);
    layer1_outputs(4435) <= (layer0_outputs(4280)) and not (layer0_outputs(5997));
    layer1_outputs(4436) <= (layer0_outputs(2880)) and (layer0_outputs(8001));
    layer1_outputs(4437) <= (layer0_outputs(4636)) and (layer0_outputs(11706));
    layer1_outputs(4438) <= layer0_outputs(2318);
    layer1_outputs(4439) <= layer0_outputs(10352);
    layer1_outputs(4440) <= not(layer0_outputs(1201));
    layer1_outputs(4441) <= (layer0_outputs(10157)) and (layer0_outputs(10601));
    layer1_outputs(4442) <= not(layer0_outputs(2440)) or (layer0_outputs(3428));
    layer1_outputs(4443) <= not(layer0_outputs(8394)) or (layer0_outputs(402));
    layer1_outputs(4444) <= not(layer0_outputs(699));
    layer1_outputs(4445) <= not(layer0_outputs(5453));
    layer1_outputs(4446) <= (layer0_outputs(7868)) or (layer0_outputs(4497));
    layer1_outputs(4447) <= layer0_outputs(9310);
    layer1_outputs(4448) <= (layer0_outputs(8763)) and not (layer0_outputs(1375));
    layer1_outputs(4449) <= (layer0_outputs(6011)) xor (layer0_outputs(6214));
    layer1_outputs(4450) <= not((layer0_outputs(2092)) or (layer0_outputs(3608)));
    layer1_outputs(4451) <= not(layer0_outputs(2266));
    layer1_outputs(4452) <= layer0_outputs(496);
    layer1_outputs(4453) <= not((layer0_outputs(11319)) or (layer0_outputs(4462)));
    layer1_outputs(4454) <= not((layer0_outputs(4988)) xor (layer0_outputs(8802)));
    layer1_outputs(4455) <= not((layer0_outputs(1821)) or (layer0_outputs(5729)));
    layer1_outputs(4456) <= not(layer0_outputs(3687));
    layer1_outputs(4457) <= layer0_outputs(10292);
    layer1_outputs(4458) <= not(layer0_outputs(12012)) or (layer0_outputs(9905));
    layer1_outputs(4459) <= '1';
    layer1_outputs(4460) <= (layer0_outputs(4201)) or (layer0_outputs(3224));
    layer1_outputs(4461) <= not(layer0_outputs(4419)) or (layer0_outputs(4985));
    layer1_outputs(4462) <= not(layer0_outputs(3878)) or (layer0_outputs(11343));
    layer1_outputs(4463) <= layer0_outputs(6375);
    layer1_outputs(4464) <= (layer0_outputs(2933)) and not (layer0_outputs(11343));
    layer1_outputs(4465) <= not((layer0_outputs(10741)) or (layer0_outputs(10515)));
    layer1_outputs(4466) <= not(layer0_outputs(2987)) or (layer0_outputs(7825));
    layer1_outputs(4467) <= not(layer0_outputs(7380));
    layer1_outputs(4468) <= '1';
    layer1_outputs(4469) <= (layer0_outputs(1995)) and not (layer0_outputs(4715));
    layer1_outputs(4470) <= not(layer0_outputs(4422)) or (layer0_outputs(9748));
    layer1_outputs(4471) <= (layer0_outputs(438)) and (layer0_outputs(1284));
    layer1_outputs(4472) <= layer0_outputs(4196);
    layer1_outputs(4473) <= (layer0_outputs(7037)) xor (layer0_outputs(11534));
    layer1_outputs(4474) <= not((layer0_outputs(4226)) xor (layer0_outputs(131)));
    layer1_outputs(4475) <= (layer0_outputs(7798)) or (layer0_outputs(6350));
    layer1_outputs(4476) <= not(layer0_outputs(6751)) or (layer0_outputs(6424));
    layer1_outputs(4477) <= not(layer0_outputs(11786)) or (layer0_outputs(9184));
    layer1_outputs(4478) <= (layer0_outputs(12654)) xor (layer0_outputs(10171));
    layer1_outputs(4479) <= layer0_outputs(359);
    layer1_outputs(4480) <= not(layer0_outputs(12442)) or (layer0_outputs(6685));
    layer1_outputs(4481) <= (layer0_outputs(12231)) or (layer0_outputs(2013));
    layer1_outputs(4482) <= not(layer0_outputs(12495)) or (layer0_outputs(12293));
    layer1_outputs(4483) <= not(layer0_outputs(2932)) or (layer0_outputs(6204));
    layer1_outputs(4484) <= (layer0_outputs(2658)) and not (layer0_outputs(9189));
    layer1_outputs(4485) <= layer0_outputs(11773);
    layer1_outputs(4486) <= layer0_outputs(1694);
    layer1_outputs(4487) <= (layer0_outputs(3196)) or (layer0_outputs(3515));
    layer1_outputs(4488) <= (layer0_outputs(9646)) and not (layer0_outputs(10152));
    layer1_outputs(4489) <= layer0_outputs(6682);
    layer1_outputs(4490) <= not((layer0_outputs(3324)) xor (layer0_outputs(3882)));
    layer1_outputs(4491) <= layer0_outputs(3229);
    layer1_outputs(4492) <= not((layer0_outputs(9106)) xor (layer0_outputs(7545)));
    layer1_outputs(4493) <= (layer0_outputs(12462)) or (layer0_outputs(3578));
    layer1_outputs(4494) <= layer0_outputs(12171);
    layer1_outputs(4495) <= (layer0_outputs(7642)) and (layer0_outputs(11789));
    layer1_outputs(4496) <= (layer0_outputs(9306)) and (layer0_outputs(1685));
    layer1_outputs(4497) <= not((layer0_outputs(7644)) and (layer0_outputs(12039)));
    layer1_outputs(4498) <= layer0_outputs(7657);
    layer1_outputs(4499) <= not((layer0_outputs(1712)) and (layer0_outputs(7353)));
    layer1_outputs(4500) <= (layer0_outputs(1007)) or (layer0_outputs(3097));
    layer1_outputs(4501) <= not((layer0_outputs(12142)) or (layer0_outputs(11968)));
    layer1_outputs(4502) <= not((layer0_outputs(8509)) and (layer0_outputs(557)));
    layer1_outputs(4503) <= not(layer0_outputs(3211)) or (layer0_outputs(7264));
    layer1_outputs(4504) <= (layer0_outputs(7296)) or (layer0_outputs(11279));
    layer1_outputs(4505) <= (layer0_outputs(12691)) and (layer0_outputs(6908));
    layer1_outputs(4506) <= not(layer0_outputs(4159));
    layer1_outputs(4507) <= (layer0_outputs(10679)) and not (layer0_outputs(686));
    layer1_outputs(4508) <= (layer0_outputs(8647)) and (layer0_outputs(9599));
    layer1_outputs(4509) <= (layer0_outputs(6280)) and (layer0_outputs(4498));
    layer1_outputs(4510) <= not(layer0_outputs(6708)) or (layer0_outputs(5138));
    layer1_outputs(4511) <= not((layer0_outputs(8598)) and (layer0_outputs(1952)));
    layer1_outputs(4512) <= not(layer0_outputs(8718));
    layer1_outputs(4513) <= (layer0_outputs(10807)) or (layer0_outputs(7242));
    layer1_outputs(4514) <= (layer0_outputs(7629)) or (layer0_outputs(2401));
    layer1_outputs(4515) <= (layer0_outputs(12622)) or (layer0_outputs(12108));
    layer1_outputs(4516) <= not(layer0_outputs(5702)) or (layer0_outputs(12176));
    layer1_outputs(4517) <= (layer0_outputs(128)) xor (layer0_outputs(6782));
    layer1_outputs(4518) <= (layer0_outputs(6136)) and (layer0_outputs(8772));
    layer1_outputs(4519) <= layer0_outputs(1057);
    layer1_outputs(4520) <= not((layer0_outputs(11800)) or (layer0_outputs(7925)));
    layer1_outputs(4521) <= (layer0_outputs(841)) xor (layer0_outputs(6439));
    layer1_outputs(4522) <= not(layer0_outputs(3107));
    layer1_outputs(4523) <= (layer0_outputs(6096)) and (layer0_outputs(9322));
    layer1_outputs(4524) <= not(layer0_outputs(1983)) or (layer0_outputs(11823));
    layer1_outputs(4525) <= not((layer0_outputs(6355)) and (layer0_outputs(2288)));
    layer1_outputs(4526) <= not(layer0_outputs(8227)) or (layer0_outputs(8643));
    layer1_outputs(4527) <= layer0_outputs(2972);
    layer1_outputs(4528) <= (layer0_outputs(6534)) and not (layer0_outputs(5151));
    layer1_outputs(4529) <= not(layer0_outputs(12296));
    layer1_outputs(4530) <= not((layer0_outputs(9839)) and (layer0_outputs(7339)));
    layer1_outputs(4531) <= (layer0_outputs(12353)) and not (layer0_outputs(3959));
    layer1_outputs(4532) <= not((layer0_outputs(8053)) and (layer0_outputs(1855)));
    layer1_outputs(4533) <= layer0_outputs(5285);
    layer1_outputs(4534) <= layer0_outputs(7886);
    layer1_outputs(4535) <= not(layer0_outputs(8631)) or (layer0_outputs(5369));
    layer1_outputs(4536) <= layer0_outputs(12449);
    layer1_outputs(4537) <= layer0_outputs(9860);
    layer1_outputs(4538) <= not((layer0_outputs(145)) or (layer0_outputs(1865)));
    layer1_outputs(4539) <= not(layer0_outputs(761)) or (layer0_outputs(9736));
    layer1_outputs(4540) <= not(layer0_outputs(9431));
    layer1_outputs(4541) <= not(layer0_outputs(3336));
    layer1_outputs(4542) <= (layer0_outputs(10381)) xor (layer0_outputs(3755));
    layer1_outputs(4543) <= layer0_outputs(5223);
    layer1_outputs(4544) <= layer0_outputs(4264);
    layer1_outputs(4545) <= not(layer0_outputs(9928));
    layer1_outputs(4546) <= (layer0_outputs(3263)) and not (layer0_outputs(2744));
    layer1_outputs(4547) <= not((layer0_outputs(275)) and (layer0_outputs(12563)));
    layer1_outputs(4548) <= not(layer0_outputs(5674));
    layer1_outputs(4549) <= (layer0_outputs(5644)) and not (layer0_outputs(1478));
    layer1_outputs(4550) <= (layer0_outputs(9586)) and (layer0_outputs(5563));
    layer1_outputs(4551) <= not(layer0_outputs(10395));
    layer1_outputs(4552) <= '1';
    layer1_outputs(4553) <= not((layer0_outputs(5295)) or (layer0_outputs(5900)));
    layer1_outputs(4554) <= layer0_outputs(7322);
    layer1_outputs(4555) <= not((layer0_outputs(1517)) or (layer0_outputs(8836)));
    layer1_outputs(4556) <= not((layer0_outputs(9368)) or (layer0_outputs(5944)));
    layer1_outputs(4557) <= (layer0_outputs(3678)) and (layer0_outputs(5752));
    layer1_outputs(4558) <= not(layer0_outputs(4495)) or (layer0_outputs(3334));
    layer1_outputs(4559) <= (layer0_outputs(1791)) and not (layer0_outputs(11855));
    layer1_outputs(4560) <= not((layer0_outputs(2282)) or (layer0_outputs(12667)));
    layer1_outputs(4561) <= not((layer0_outputs(893)) and (layer0_outputs(7667)));
    layer1_outputs(4562) <= not(layer0_outputs(11730)) or (layer0_outputs(11915));
    layer1_outputs(4563) <= not(layer0_outputs(8186));
    layer1_outputs(4564) <= layer0_outputs(1419);
    layer1_outputs(4565) <= not(layer0_outputs(12401));
    layer1_outputs(4566) <= not(layer0_outputs(1488)) or (layer0_outputs(2451));
    layer1_outputs(4567) <= (layer0_outputs(244)) and not (layer0_outputs(3873));
    layer1_outputs(4568) <= layer0_outputs(1741);
    layer1_outputs(4569) <= layer0_outputs(291);
    layer1_outputs(4570) <= not((layer0_outputs(9051)) and (layer0_outputs(5534)));
    layer1_outputs(4571) <= not((layer0_outputs(1002)) and (layer0_outputs(3483)));
    layer1_outputs(4572) <= layer0_outputs(5203);
    layer1_outputs(4573) <= layer0_outputs(2848);
    layer1_outputs(4574) <= (layer0_outputs(8365)) xor (layer0_outputs(1624));
    layer1_outputs(4575) <= not(layer0_outputs(6244));
    layer1_outputs(4576) <= (layer0_outputs(12516)) and not (layer0_outputs(9168));
    layer1_outputs(4577) <= not((layer0_outputs(10694)) or (layer0_outputs(2486)));
    layer1_outputs(4578) <= not(layer0_outputs(12043)) or (layer0_outputs(3183));
    layer1_outputs(4579) <= not(layer0_outputs(6640));
    layer1_outputs(4580) <= not((layer0_outputs(6837)) and (layer0_outputs(1778)));
    layer1_outputs(4581) <= layer0_outputs(12187);
    layer1_outputs(4582) <= not(layer0_outputs(5496)) or (layer0_outputs(11304));
    layer1_outputs(4583) <= not((layer0_outputs(694)) or (layer0_outputs(10535)));
    layer1_outputs(4584) <= (layer0_outputs(1501)) xor (layer0_outputs(117));
    layer1_outputs(4585) <= not(layer0_outputs(9211)) or (layer0_outputs(324));
    layer1_outputs(4586) <= layer0_outputs(12642);
    layer1_outputs(4587) <= layer0_outputs(7348);
    layer1_outputs(4588) <= not(layer0_outputs(4455));
    layer1_outputs(4589) <= layer0_outputs(1830);
    layer1_outputs(4590) <= (layer0_outputs(9307)) and not (layer0_outputs(9601));
    layer1_outputs(4591) <= not(layer0_outputs(10534)) or (layer0_outputs(8724));
    layer1_outputs(4592) <= not(layer0_outputs(459));
    layer1_outputs(4593) <= layer0_outputs(3604);
    layer1_outputs(4594) <= not(layer0_outputs(7288)) or (layer0_outputs(834));
    layer1_outputs(4595) <= not(layer0_outputs(3287));
    layer1_outputs(4596) <= layer0_outputs(10315);
    layer1_outputs(4597) <= (layer0_outputs(4486)) and not (layer0_outputs(4020));
    layer1_outputs(4598) <= not(layer0_outputs(5133));
    layer1_outputs(4599) <= not(layer0_outputs(2006)) or (layer0_outputs(10555));
    layer1_outputs(4600) <= not(layer0_outputs(3641));
    layer1_outputs(4601) <= not(layer0_outputs(8120));
    layer1_outputs(4602) <= not(layer0_outputs(5315)) or (layer0_outputs(2973));
    layer1_outputs(4603) <= layer0_outputs(8483);
    layer1_outputs(4604) <= not(layer0_outputs(2834)) or (layer0_outputs(2420));
    layer1_outputs(4605) <= not(layer0_outputs(6208));
    layer1_outputs(4606) <= (layer0_outputs(5118)) and (layer0_outputs(10971));
    layer1_outputs(4607) <= layer0_outputs(12415);
    layer1_outputs(4608) <= (layer0_outputs(7929)) or (layer0_outputs(11244));
    layer1_outputs(4609) <= layer0_outputs(4433);
    layer1_outputs(4610) <= (layer0_outputs(2022)) and (layer0_outputs(6541));
    layer1_outputs(4611) <= (layer0_outputs(7475)) and not (layer0_outputs(5926));
    layer1_outputs(4612) <= (layer0_outputs(6458)) xor (layer0_outputs(6672));
    layer1_outputs(4613) <= (layer0_outputs(1560)) and not (layer0_outputs(1796));
    layer1_outputs(4614) <= not(layer0_outputs(5213)) or (layer0_outputs(423));
    layer1_outputs(4615) <= (layer0_outputs(5688)) and (layer0_outputs(9448));
    layer1_outputs(4616) <= layer0_outputs(12580);
    layer1_outputs(4617) <= not(layer0_outputs(591)) or (layer0_outputs(6251));
    layer1_outputs(4618) <= layer0_outputs(10345);
    layer1_outputs(4619) <= (layer0_outputs(1132)) and not (layer0_outputs(3888));
    layer1_outputs(4620) <= not(layer0_outputs(9912));
    layer1_outputs(4621) <= not(layer0_outputs(4524)) or (layer0_outputs(11054));
    layer1_outputs(4622) <= not(layer0_outputs(9070)) or (layer0_outputs(5074));
    layer1_outputs(4623) <= not(layer0_outputs(7187));
    layer1_outputs(4624) <= not((layer0_outputs(3450)) or (layer0_outputs(2653)));
    layer1_outputs(4625) <= not(layer0_outputs(7294)) or (layer0_outputs(9253));
    layer1_outputs(4626) <= '1';
    layer1_outputs(4627) <= not(layer0_outputs(730));
    layer1_outputs(4628) <= (layer0_outputs(6886)) and not (layer0_outputs(9321));
    layer1_outputs(4629) <= layer0_outputs(1825);
    layer1_outputs(4630) <= not(layer0_outputs(2650));
    layer1_outputs(4631) <= not((layer0_outputs(3584)) and (layer0_outputs(912)));
    layer1_outputs(4632) <= not(layer0_outputs(8743));
    layer1_outputs(4633) <= (layer0_outputs(1293)) and (layer0_outputs(4373));
    layer1_outputs(4634) <= not((layer0_outputs(209)) or (layer0_outputs(8988)));
    layer1_outputs(4635) <= not(layer0_outputs(12060)) or (layer0_outputs(2255));
    layer1_outputs(4636) <= not((layer0_outputs(654)) xor (layer0_outputs(8583)));
    layer1_outputs(4637) <= (layer0_outputs(10643)) or (layer0_outputs(715));
    layer1_outputs(4638) <= not(layer0_outputs(630)) or (layer0_outputs(4995));
    layer1_outputs(4639) <= not((layer0_outputs(10704)) and (layer0_outputs(3488)));
    layer1_outputs(4640) <= not(layer0_outputs(9344));
    layer1_outputs(4641) <= (layer0_outputs(2491)) and not (layer0_outputs(9059));
    layer1_outputs(4642) <= not((layer0_outputs(2970)) xor (layer0_outputs(7999)));
    layer1_outputs(4643) <= '1';
    layer1_outputs(4644) <= layer0_outputs(294);
    layer1_outputs(4645) <= not((layer0_outputs(3819)) and (layer0_outputs(11550)));
    layer1_outputs(4646) <= not(layer0_outputs(5033)) or (layer0_outputs(222));
    layer1_outputs(4647) <= layer0_outputs(10745);
    layer1_outputs(4648) <= not(layer0_outputs(5784));
    layer1_outputs(4649) <= (layer0_outputs(6189)) and (layer0_outputs(6338));
    layer1_outputs(4650) <= not(layer0_outputs(4855));
    layer1_outputs(4651) <= (layer0_outputs(9765)) and not (layer0_outputs(3946));
    layer1_outputs(4652) <= '0';
    layer1_outputs(4653) <= layer0_outputs(16);
    layer1_outputs(4654) <= not(layer0_outputs(4175));
    layer1_outputs(4655) <= layer0_outputs(5202);
    layer1_outputs(4656) <= layer0_outputs(7003);
    layer1_outputs(4657) <= not(layer0_outputs(8176));
    layer1_outputs(4658) <= not((layer0_outputs(3222)) and (layer0_outputs(5318)));
    layer1_outputs(4659) <= layer0_outputs(3363);
    layer1_outputs(4660) <= '0';
    layer1_outputs(4661) <= (layer0_outputs(6371)) and not (layer0_outputs(11281));
    layer1_outputs(4662) <= (layer0_outputs(772)) or (layer0_outputs(5820));
    layer1_outputs(4663) <= not(layer0_outputs(6010));
    layer1_outputs(4664) <= not(layer0_outputs(11103));
    layer1_outputs(4665) <= not(layer0_outputs(6928));
    layer1_outputs(4666) <= (layer0_outputs(3168)) xor (layer0_outputs(8362));
    layer1_outputs(4667) <= layer0_outputs(170);
    layer1_outputs(4668) <= not(layer0_outputs(10700));
    layer1_outputs(4669) <= (layer0_outputs(11049)) and not (layer0_outputs(2565));
    layer1_outputs(4670) <= not(layer0_outputs(4882));
    layer1_outputs(4671) <= (layer0_outputs(5162)) and not (layer0_outputs(723));
    layer1_outputs(4672) <= not(layer0_outputs(9540)) or (layer0_outputs(7383));
    layer1_outputs(4673) <= (layer0_outputs(427)) and not (layer0_outputs(6618));
    layer1_outputs(4674) <= not(layer0_outputs(2045));
    layer1_outputs(4675) <= (layer0_outputs(2059)) xor (layer0_outputs(12363));
    layer1_outputs(4676) <= (layer0_outputs(7316)) xor (layer0_outputs(9051));
    layer1_outputs(4677) <= not((layer0_outputs(7827)) or (layer0_outputs(2700)));
    layer1_outputs(4678) <= not(layer0_outputs(6681)) or (layer0_outputs(1279));
    layer1_outputs(4679) <= not(layer0_outputs(11214));
    layer1_outputs(4680) <= not((layer0_outputs(4086)) and (layer0_outputs(8512)));
    layer1_outputs(4681) <= (layer0_outputs(8081)) and not (layer0_outputs(1706));
    layer1_outputs(4682) <= (layer0_outputs(8315)) and (layer0_outputs(3464));
    layer1_outputs(4683) <= not(layer0_outputs(11693)) or (layer0_outputs(2233));
    layer1_outputs(4684) <= layer0_outputs(8060);
    layer1_outputs(4685) <= layer0_outputs(2535);
    layer1_outputs(4686) <= layer0_outputs(5940);
    layer1_outputs(4687) <= not(layer0_outputs(8276));
    layer1_outputs(4688) <= not(layer0_outputs(7399));
    layer1_outputs(4689) <= not(layer0_outputs(6874));
    layer1_outputs(4690) <= '0';
    layer1_outputs(4691) <= not(layer0_outputs(693));
    layer1_outputs(4692) <= (layer0_outputs(10518)) and not (layer0_outputs(5281));
    layer1_outputs(4693) <= layer0_outputs(6168);
    layer1_outputs(4694) <= (layer0_outputs(2351)) and (layer0_outputs(4979));
    layer1_outputs(4695) <= (layer0_outputs(9040)) xor (layer0_outputs(12798));
    layer1_outputs(4696) <= (layer0_outputs(6077)) and not (layer0_outputs(12300));
    layer1_outputs(4697) <= (layer0_outputs(24)) and not (layer0_outputs(1260));
    layer1_outputs(4698) <= layer0_outputs(12419);
    layer1_outputs(4699) <= '1';
    layer1_outputs(4700) <= not(layer0_outputs(10916));
    layer1_outputs(4701) <= layer0_outputs(8080);
    layer1_outputs(4702) <= layer0_outputs(971);
    layer1_outputs(4703) <= not(layer0_outputs(3842)) or (layer0_outputs(8698));
    layer1_outputs(4704) <= not((layer0_outputs(9964)) xor (layer0_outputs(10172)));
    layer1_outputs(4705) <= (layer0_outputs(1996)) xor (layer0_outputs(4958));
    layer1_outputs(4706) <= not(layer0_outputs(11652));
    layer1_outputs(4707) <= not((layer0_outputs(4165)) or (layer0_outputs(9791)));
    layer1_outputs(4708) <= layer0_outputs(6485);
    layer1_outputs(4709) <= not((layer0_outputs(2905)) xor (layer0_outputs(2505)));
    layer1_outputs(4710) <= not(layer0_outputs(6551));
    layer1_outputs(4711) <= layer0_outputs(6114);
    layer1_outputs(4712) <= not(layer0_outputs(8123));
    layer1_outputs(4713) <= not((layer0_outputs(3964)) or (layer0_outputs(11990)));
    layer1_outputs(4714) <= not(layer0_outputs(4576));
    layer1_outputs(4715) <= not(layer0_outputs(7646));
    layer1_outputs(4716) <= not((layer0_outputs(8837)) xor (layer0_outputs(2514)));
    layer1_outputs(4717) <= (layer0_outputs(11053)) and (layer0_outputs(9445));
    layer1_outputs(4718) <= not((layer0_outputs(1191)) xor (layer0_outputs(65)));
    layer1_outputs(4719) <= (layer0_outputs(3038)) and not (layer0_outputs(10027));
    layer1_outputs(4720) <= layer0_outputs(5123);
    layer1_outputs(4721) <= not((layer0_outputs(8970)) or (layer0_outputs(6273)));
    layer1_outputs(4722) <= not((layer0_outputs(11955)) and (layer0_outputs(12128)));
    layer1_outputs(4723) <= '0';
    layer1_outputs(4724) <= (layer0_outputs(6731)) and not (layer0_outputs(124));
    layer1_outputs(4725) <= layer0_outputs(10721);
    layer1_outputs(4726) <= not((layer0_outputs(11086)) and (layer0_outputs(3253)));
    layer1_outputs(4727) <= (layer0_outputs(6307)) or (layer0_outputs(8808));
    layer1_outputs(4728) <= not(layer0_outputs(7219)) or (layer0_outputs(8747));
    layer1_outputs(4729) <= layer0_outputs(9455);
    layer1_outputs(4730) <= layer0_outputs(2800);
    layer1_outputs(4731) <= layer0_outputs(5870);
    layer1_outputs(4732) <= (layer0_outputs(11440)) and not (layer0_outputs(11974));
    layer1_outputs(4733) <= (layer0_outputs(12736)) and not (layer0_outputs(4520));
    layer1_outputs(4734) <= not((layer0_outputs(5488)) xor (layer0_outputs(4992)));
    layer1_outputs(4735) <= not((layer0_outputs(5386)) and (layer0_outputs(7497)));
    layer1_outputs(4736) <= not(layer0_outputs(2511)) or (layer0_outputs(1585));
    layer1_outputs(4737) <= not((layer0_outputs(1953)) xor (layer0_outputs(4739)));
    layer1_outputs(4738) <= (layer0_outputs(7723)) and not (layer0_outputs(11357));
    layer1_outputs(4739) <= layer0_outputs(1908);
    layer1_outputs(4740) <= not(layer0_outputs(11933));
    layer1_outputs(4741) <= not(layer0_outputs(10263)) or (layer0_outputs(11093));
    layer1_outputs(4742) <= not(layer0_outputs(3855)) or (layer0_outputs(5479));
    layer1_outputs(4743) <= layer0_outputs(6988);
    layer1_outputs(4744) <= not(layer0_outputs(3787)) or (layer0_outputs(1515));
    layer1_outputs(4745) <= not(layer0_outputs(9837));
    layer1_outputs(4746) <= (layer0_outputs(5282)) and (layer0_outputs(8025));
    layer1_outputs(4747) <= layer0_outputs(11383);
    layer1_outputs(4748) <= layer0_outputs(11194);
    layer1_outputs(4749) <= layer0_outputs(10887);
    layer1_outputs(4750) <= not(layer0_outputs(4909));
    layer1_outputs(4751) <= not(layer0_outputs(2358));
    layer1_outputs(4752) <= (layer0_outputs(6069)) and (layer0_outputs(5851));
    layer1_outputs(4753) <= not((layer0_outputs(5415)) and (layer0_outputs(2801)));
    layer1_outputs(4754) <= (layer0_outputs(3962)) and not (layer0_outputs(2814));
    layer1_outputs(4755) <= (layer0_outputs(100)) or (layer0_outputs(8572));
    layer1_outputs(4756) <= (layer0_outputs(8031)) and not (layer0_outputs(9216));
    layer1_outputs(4757) <= (layer0_outputs(34)) xor (layer0_outputs(6353));
    layer1_outputs(4758) <= not((layer0_outputs(4205)) xor (layer0_outputs(1373)));
    layer1_outputs(4759) <= layer0_outputs(7);
    layer1_outputs(4760) <= layer0_outputs(6212);
    layer1_outputs(4761) <= (layer0_outputs(4359)) and not (layer0_outputs(1450));
    layer1_outputs(4762) <= layer0_outputs(11382);
    layer1_outputs(4763) <= not(layer0_outputs(7474));
    layer1_outputs(4764) <= not(layer0_outputs(2442));
    layer1_outputs(4765) <= (layer0_outputs(5158)) or (layer0_outputs(3042));
    layer1_outputs(4766) <= not(layer0_outputs(2476)) or (layer0_outputs(11572));
    layer1_outputs(4767) <= (layer0_outputs(873)) or (layer0_outputs(10506));
    layer1_outputs(4768) <= not(layer0_outputs(8906));
    layer1_outputs(4769) <= (layer0_outputs(1185)) xor (layer0_outputs(4585));
    layer1_outputs(4770) <= layer0_outputs(12281);
    layer1_outputs(4771) <= (layer0_outputs(1871)) or (layer0_outputs(7073));
    layer1_outputs(4772) <= not(layer0_outputs(5409)) or (layer0_outputs(7009));
    layer1_outputs(4773) <= (layer0_outputs(7342)) and (layer0_outputs(12464));
    layer1_outputs(4774) <= (layer0_outputs(4362)) or (layer0_outputs(4582));
    layer1_outputs(4775) <= not(layer0_outputs(5329)) or (layer0_outputs(6341));
    layer1_outputs(4776) <= layer0_outputs(271);
    layer1_outputs(4777) <= (layer0_outputs(3281)) xor (layer0_outputs(11389));
    layer1_outputs(4778) <= layer0_outputs(8486);
    layer1_outputs(4779) <= not(layer0_outputs(11313));
    layer1_outputs(4780) <= not(layer0_outputs(5287));
    layer1_outputs(4781) <= (layer0_outputs(8594)) and not (layer0_outputs(3542));
    layer1_outputs(4782) <= layer0_outputs(852);
    layer1_outputs(4783) <= layer0_outputs(12547);
    layer1_outputs(4784) <= layer0_outputs(10585);
    layer1_outputs(4785) <= not(layer0_outputs(8969));
    layer1_outputs(4786) <= not((layer0_outputs(11016)) or (layer0_outputs(2581)));
    layer1_outputs(4787) <= (layer0_outputs(169)) xor (layer0_outputs(11478));
    layer1_outputs(4788) <= not(layer0_outputs(10933));
    layer1_outputs(4789) <= (layer0_outputs(3917)) and (layer0_outputs(4125));
    layer1_outputs(4790) <= layer0_outputs(11776);
    layer1_outputs(4791) <= not(layer0_outputs(11970)) or (layer0_outputs(3593));
    layer1_outputs(4792) <= (layer0_outputs(6620)) and not (layer0_outputs(12774));
    layer1_outputs(4793) <= not(layer0_outputs(361));
    layer1_outputs(4794) <= layer0_outputs(11449);
    layer1_outputs(4795) <= '1';
    layer1_outputs(4796) <= not(layer0_outputs(236)) or (layer0_outputs(4616));
    layer1_outputs(4797) <= layer0_outputs(9623);
    layer1_outputs(4798) <= (layer0_outputs(7485)) and not (layer0_outputs(4515));
    layer1_outputs(4799) <= not(layer0_outputs(11756));
    layer1_outputs(4800) <= (layer0_outputs(3407)) and not (layer0_outputs(2038));
    layer1_outputs(4801) <= not((layer0_outputs(9418)) or (layer0_outputs(1015)));
    layer1_outputs(4802) <= layer0_outputs(2150);
    layer1_outputs(4803) <= layer0_outputs(9880);
    layer1_outputs(4804) <= not((layer0_outputs(576)) and (layer0_outputs(9548)));
    layer1_outputs(4805) <= layer0_outputs(7208);
    layer1_outputs(4806) <= (layer0_outputs(5002)) and (layer0_outputs(5652));
    layer1_outputs(4807) <= not(layer0_outputs(4778));
    layer1_outputs(4808) <= not((layer0_outputs(6491)) xor (layer0_outputs(10939)));
    layer1_outputs(4809) <= (layer0_outputs(2419)) and not (layer0_outputs(587));
    layer1_outputs(4810) <= (layer0_outputs(12661)) or (layer0_outputs(2121));
    layer1_outputs(4811) <= (layer0_outputs(1647)) and not (layer0_outputs(11161));
    layer1_outputs(4812) <= (layer0_outputs(12057)) xor (layer0_outputs(9970));
    layer1_outputs(4813) <= not(layer0_outputs(6254));
    layer1_outputs(4814) <= (layer0_outputs(8902)) xor (layer0_outputs(1727));
    layer1_outputs(4815) <= (layer0_outputs(6402)) and (layer0_outputs(90));
    layer1_outputs(4816) <= not((layer0_outputs(7771)) and (layer0_outputs(3559)));
    layer1_outputs(4817) <= not(layer0_outputs(9688));
    layer1_outputs(4818) <= (layer0_outputs(6610)) and not (layer0_outputs(9439));
    layer1_outputs(4819) <= layer0_outputs(8005);
    layer1_outputs(4820) <= (layer0_outputs(1707)) and not (layer0_outputs(12298));
    layer1_outputs(4821) <= layer0_outputs(166);
    layer1_outputs(4822) <= (layer0_outputs(1458)) and not (layer0_outputs(279));
    layer1_outputs(4823) <= (layer0_outputs(10193)) and not (layer0_outputs(1669));
    layer1_outputs(4824) <= (layer0_outputs(4706)) and not (layer0_outputs(2135));
    layer1_outputs(4825) <= not((layer0_outputs(9462)) or (layer0_outputs(72)));
    layer1_outputs(4826) <= not(layer0_outputs(4452));
    layer1_outputs(4827) <= (layer0_outputs(10732)) or (layer0_outputs(4275));
    layer1_outputs(4828) <= not((layer0_outputs(1177)) or (layer0_outputs(814)));
    layer1_outputs(4829) <= layer0_outputs(1124);
    layer1_outputs(4830) <= not((layer0_outputs(2962)) or (layer0_outputs(9069)));
    layer1_outputs(4831) <= layer0_outputs(6122);
    layer1_outputs(4832) <= not(layer0_outputs(7390));
    layer1_outputs(4833) <= (layer0_outputs(3002)) or (layer0_outputs(12549));
    layer1_outputs(4834) <= (layer0_outputs(12596)) and (layer0_outputs(12184));
    layer1_outputs(4835) <= (layer0_outputs(2402)) and not (layer0_outputs(8759));
    layer1_outputs(4836) <= (layer0_outputs(8078)) and not (layer0_outputs(9775));
    layer1_outputs(4837) <= not(layer0_outputs(614)) or (layer0_outputs(7986));
    layer1_outputs(4838) <= not((layer0_outputs(11059)) or (layer0_outputs(6914)));
    layer1_outputs(4839) <= (layer0_outputs(12166)) and not (layer0_outputs(718));
    layer1_outputs(4840) <= (layer0_outputs(3159)) and not (layer0_outputs(6223));
    layer1_outputs(4841) <= not(layer0_outputs(491));
    layer1_outputs(4842) <= layer0_outputs(9648);
    layer1_outputs(4843) <= (layer0_outputs(9664)) or (layer0_outputs(8423));
    layer1_outputs(4844) <= not(layer0_outputs(6311));
    layer1_outputs(4845) <= (layer0_outputs(5190)) xor (layer0_outputs(768));
    layer1_outputs(4846) <= not((layer0_outputs(10336)) and (layer0_outputs(9539)));
    layer1_outputs(4847) <= layer0_outputs(639);
    layer1_outputs(4848) <= (layer0_outputs(5577)) or (layer0_outputs(6899));
    layer1_outputs(4849) <= not((layer0_outputs(2503)) and (layer0_outputs(9772)));
    layer1_outputs(4850) <= (layer0_outputs(10185)) and not (layer0_outputs(10903));
    layer1_outputs(4851) <= (layer0_outputs(471)) and not (layer0_outputs(11819));
    layer1_outputs(4852) <= not((layer0_outputs(6870)) xor (layer0_outputs(9257)));
    layer1_outputs(4853) <= '0';
    layer1_outputs(4854) <= layer0_outputs(11727);
    layer1_outputs(4855) <= '0';
    layer1_outputs(4856) <= not(layer0_outputs(9852));
    layer1_outputs(4857) <= (layer0_outputs(6598)) and (layer0_outputs(11401));
    layer1_outputs(4858) <= not(layer0_outputs(10356)) or (layer0_outputs(4107));
    layer1_outputs(4859) <= not(layer0_outputs(9281)) or (layer0_outputs(10410));
    layer1_outputs(4860) <= not((layer0_outputs(12635)) or (layer0_outputs(6250)));
    layer1_outputs(4861) <= not((layer0_outputs(3468)) or (layer0_outputs(11135)));
    layer1_outputs(4862) <= not(layer0_outputs(10075)) or (layer0_outputs(7845));
    layer1_outputs(4863) <= not(layer0_outputs(4631)) or (layer0_outputs(9012));
    layer1_outputs(4864) <= (layer0_outputs(1101)) and (layer0_outputs(12668));
    layer1_outputs(4865) <= layer0_outputs(9653);
    layer1_outputs(4866) <= not(layer0_outputs(5907));
    layer1_outputs(4867) <= layer0_outputs(6762);
    layer1_outputs(4868) <= not(layer0_outputs(11923));
    layer1_outputs(4869) <= not(layer0_outputs(1052));
    layer1_outputs(4870) <= not(layer0_outputs(261)) or (layer0_outputs(29));
    layer1_outputs(4871) <= '0';
    layer1_outputs(4872) <= not((layer0_outputs(6030)) xor (layer0_outputs(1441)));
    layer1_outputs(4873) <= not((layer0_outputs(2031)) and (layer0_outputs(9179)));
    layer1_outputs(4874) <= (layer0_outputs(9519)) xor (layer0_outputs(5376));
    layer1_outputs(4875) <= not(layer0_outputs(11136));
    layer1_outputs(4876) <= layer0_outputs(9804);
    layer1_outputs(4877) <= layer0_outputs(8555);
    layer1_outputs(4878) <= not((layer0_outputs(5276)) or (layer0_outputs(11646)));
    layer1_outputs(4879) <= (layer0_outputs(3812)) and (layer0_outputs(12522));
    layer1_outputs(4880) <= (layer0_outputs(5078)) and not (layer0_outputs(3480));
    layer1_outputs(4881) <= layer0_outputs(12132);
    layer1_outputs(4882) <= (layer0_outputs(3311)) or (layer0_outputs(4531));
    layer1_outputs(4883) <= not((layer0_outputs(3221)) or (layer0_outputs(11338)));
    layer1_outputs(4884) <= not(layer0_outputs(9188)) or (layer0_outputs(9117));
    layer1_outputs(4885) <= (layer0_outputs(11081)) and not (layer0_outputs(7174));
    layer1_outputs(4886) <= not(layer0_outputs(259));
    layer1_outputs(4887) <= not((layer0_outputs(7603)) or (layer0_outputs(1142)));
    layer1_outputs(4888) <= (layer0_outputs(916)) xor (layer0_outputs(8915));
    layer1_outputs(4889) <= not(layer0_outputs(10189));
    layer1_outputs(4890) <= not(layer0_outputs(7156));
    layer1_outputs(4891) <= (layer0_outputs(11070)) and not (layer0_outputs(10116));
    layer1_outputs(4892) <= not(layer0_outputs(1908)) or (layer0_outputs(3474));
    layer1_outputs(4893) <= not((layer0_outputs(2192)) and (layer0_outputs(10682)));
    layer1_outputs(4894) <= layer0_outputs(11758);
    layer1_outputs(4895) <= (layer0_outputs(12358)) and (layer0_outputs(3209));
    layer1_outputs(4896) <= not(layer0_outputs(5085));
    layer1_outputs(4897) <= (layer0_outputs(9024)) and not (layer0_outputs(1896));
    layer1_outputs(4898) <= not((layer0_outputs(9199)) or (layer0_outputs(1955)));
    layer1_outputs(4899) <= (layer0_outputs(3525)) or (layer0_outputs(4781));
    layer1_outputs(4900) <= (layer0_outputs(6178)) and not (layer0_outputs(7667));
    layer1_outputs(4901) <= not(layer0_outputs(108));
    layer1_outputs(4902) <= not((layer0_outputs(5696)) or (layer0_outputs(12465)));
    layer1_outputs(4903) <= not(layer0_outputs(9826));
    layer1_outputs(4904) <= not(layer0_outputs(9741));
    layer1_outputs(4905) <= not((layer0_outputs(7185)) or (layer0_outputs(5529)));
    layer1_outputs(4906) <= not(layer0_outputs(7087));
    layer1_outputs(4907) <= layer0_outputs(6021);
    layer1_outputs(4908) <= (layer0_outputs(1447)) and not (layer0_outputs(2966));
    layer1_outputs(4909) <= not((layer0_outputs(6474)) or (layer0_outputs(3344)));
    layer1_outputs(4910) <= not(layer0_outputs(8387));
    layer1_outputs(4911) <= not((layer0_outputs(11866)) xor (layer0_outputs(11160)));
    layer1_outputs(4912) <= not(layer0_outputs(7123));
    layer1_outputs(4913) <= (layer0_outputs(1690)) and (layer0_outputs(7476));
    layer1_outputs(4914) <= not(layer0_outputs(4167)) or (layer0_outputs(8483));
    layer1_outputs(4915) <= not(layer0_outputs(10070)) or (layer0_outputs(10692));
    layer1_outputs(4916) <= not(layer0_outputs(4840));
    layer1_outputs(4917) <= not((layer0_outputs(6446)) xor (layer0_outputs(2249)));
    layer1_outputs(4918) <= layer0_outputs(1205);
    layer1_outputs(4919) <= '0';
    layer1_outputs(4920) <= (layer0_outputs(5308)) or (layer0_outputs(3094));
    layer1_outputs(4921) <= layer0_outputs(711);
    layer1_outputs(4922) <= (layer0_outputs(12472)) or (layer0_outputs(9757));
    layer1_outputs(4923) <= not(layer0_outputs(2212));
    layer1_outputs(4924) <= not((layer0_outputs(1762)) or (layer0_outputs(7406)));
    layer1_outputs(4925) <= (layer0_outputs(532)) and not (layer0_outputs(1237));
    layer1_outputs(4926) <= (layer0_outputs(6473)) and not (layer0_outputs(5868));
    layer1_outputs(4927) <= not(layer0_outputs(1664)) or (layer0_outputs(10047));
    layer1_outputs(4928) <= not(layer0_outputs(10989));
    layer1_outputs(4929) <= layer0_outputs(7586);
    layer1_outputs(4930) <= not((layer0_outputs(2946)) and (layer0_outputs(2859)));
    layer1_outputs(4931) <= (layer0_outputs(3952)) or (layer0_outputs(11360));
    layer1_outputs(4932) <= not(layer0_outputs(4313));
    layer1_outputs(4933) <= not(layer0_outputs(11149)) or (layer0_outputs(8676));
    layer1_outputs(4934) <= (layer0_outputs(3984)) and (layer0_outputs(12652));
    layer1_outputs(4935) <= (layer0_outputs(6794)) xor (layer0_outputs(5205));
    layer1_outputs(4936) <= not(layer0_outputs(5057));
    layer1_outputs(4937) <= not(layer0_outputs(3215)) or (layer0_outputs(7249));
    layer1_outputs(4938) <= (layer0_outputs(5049)) and not (layer0_outputs(11925));
    layer1_outputs(4939) <= layer0_outputs(1400);
    layer1_outputs(4940) <= (layer0_outputs(10271)) xor (layer0_outputs(11616));
    layer1_outputs(4941) <= (layer0_outputs(5823)) xor (layer0_outputs(8005));
    layer1_outputs(4942) <= (layer0_outputs(11984)) and not (layer0_outputs(1407));
    layer1_outputs(4943) <= not(layer0_outputs(1609));
    layer1_outputs(4944) <= not(layer0_outputs(4011)) or (layer0_outputs(6700));
    layer1_outputs(4945) <= not(layer0_outputs(5311));
    layer1_outputs(4946) <= (layer0_outputs(3466)) and (layer0_outputs(4145));
    layer1_outputs(4947) <= (layer0_outputs(10841)) and not (layer0_outputs(8269));
    layer1_outputs(4948) <= (layer0_outputs(1633)) and not (layer0_outputs(9801));
    layer1_outputs(4949) <= (layer0_outputs(2983)) and (layer0_outputs(121));
    layer1_outputs(4950) <= (layer0_outputs(7358)) and not (layer0_outputs(9055));
    layer1_outputs(4951) <= (layer0_outputs(9498)) and not (layer0_outputs(7804));
    layer1_outputs(4952) <= (layer0_outputs(3201)) and not (layer0_outputs(3001));
    layer1_outputs(4953) <= not(layer0_outputs(826));
    layer1_outputs(4954) <= layer0_outputs(10582);
    layer1_outputs(4955) <= layer0_outputs(5251);
    layer1_outputs(4956) <= layer0_outputs(11384);
    layer1_outputs(4957) <= (layer0_outputs(3983)) or (layer0_outputs(7967));
    layer1_outputs(4958) <= (layer0_outputs(10949)) and (layer0_outputs(10547));
    layer1_outputs(4959) <= (layer0_outputs(1103)) and not (layer0_outputs(5692));
    layer1_outputs(4960) <= layer0_outputs(1127);
    layer1_outputs(4961) <= not(layer0_outputs(10500));
    layer1_outputs(4962) <= not((layer0_outputs(2892)) or (layer0_outputs(8430)));
    layer1_outputs(4963) <= layer0_outputs(2404);
    layer1_outputs(4964) <= not((layer0_outputs(11266)) and (layer0_outputs(927)));
    layer1_outputs(4965) <= not(layer0_outputs(3272));
    layer1_outputs(4966) <= not(layer0_outputs(7134)) or (layer0_outputs(3372));
    layer1_outputs(4967) <= (layer0_outputs(11636)) xor (layer0_outputs(4301));
    layer1_outputs(4968) <= layer0_outputs(11267);
    layer1_outputs(4969) <= not(layer0_outputs(5999)) or (layer0_outputs(11924));
    layer1_outputs(4970) <= not(layer0_outputs(11837));
    layer1_outputs(4971) <= (layer0_outputs(6482)) and not (layer0_outputs(12270));
    layer1_outputs(4972) <= (layer0_outputs(3496)) and not (layer0_outputs(12212));
    layer1_outputs(4973) <= not(layer0_outputs(10478));
    layer1_outputs(4974) <= not((layer0_outputs(1783)) or (layer0_outputs(11450)));
    layer1_outputs(4975) <= (layer0_outputs(2682)) and not (layer0_outputs(3765));
    layer1_outputs(4976) <= not(layer0_outputs(5158)) or (layer0_outputs(2583));
    layer1_outputs(4977) <= layer0_outputs(10214);
    layer1_outputs(4978) <= (layer0_outputs(12240)) or (layer0_outputs(6535));
    layer1_outputs(4979) <= layer0_outputs(11667);
    layer1_outputs(4980) <= (layer0_outputs(9024)) and not (layer0_outputs(4749));
    layer1_outputs(4981) <= not((layer0_outputs(3788)) xor (layer0_outputs(690)));
    layer1_outputs(4982) <= (layer0_outputs(11180)) and (layer0_outputs(5483));
    layer1_outputs(4983) <= (layer0_outputs(9129)) and not (layer0_outputs(1296));
    layer1_outputs(4984) <= not((layer0_outputs(3822)) xor (layer0_outputs(1494)));
    layer1_outputs(4985) <= not((layer0_outputs(12195)) and (layer0_outputs(10855)));
    layer1_outputs(4986) <= (layer0_outputs(968)) and (layer0_outputs(10747));
    layer1_outputs(4987) <= layer0_outputs(12679);
    layer1_outputs(4988) <= not(layer0_outputs(10300)) or (layer0_outputs(1022));
    layer1_outputs(4989) <= not(layer0_outputs(2927));
    layer1_outputs(4990) <= (layer0_outputs(7808)) or (layer0_outputs(11073));
    layer1_outputs(4991) <= layer0_outputs(7431);
    layer1_outputs(4992) <= not(layer0_outputs(6044));
    layer1_outputs(4993) <= (layer0_outputs(5548)) or (layer0_outputs(6779));
    layer1_outputs(4994) <= not(layer0_outputs(5721));
    layer1_outputs(4995) <= not(layer0_outputs(10570));
    layer1_outputs(4996) <= not(layer0_outputs(7004));
    layer1_outputs(4997) <= layer0_outputs(6972);
    layer1_outputs(4998) <= not(layer0_outputs(5619));
    layer1_outputs(4999) <= (layer0_outputs(3237)) or (layer0_outputs(2888));
    layer1_outputs(5000) <= not((layer0_outputs(1864)) or (layer0_outputs(1175)));
    layer1_outputs(5001) <= not(layer0_outputs(4081)) or (layer0_outputs(1085));
    layer1_outputs(5002) <= not(layer0_outputs(12489)) or (layer0_outputs(10498));
    layer1_outputs(5003) <= not(layer0_outputs(8493));
    layer1_outputs(5004) <= not(layer0_outputs(267));
    layer1_outputs(5005) <= not(layer0_outputs(1464));
    layer1_outputs(5006) <= layer0_outputs(9034);
    layer1_outputs(5007) <= not((layer0_outputs(5176)) and (layer0_outputs(11151)));
    layer1_outputs(5008) <= not(layer0_outputs(10778));
    layer1_outputs(5009) <= not(layer0_outputs(4296));
    layer1_outputs(5010) <= not(layer0_outputs(10768));
    layer1_outputs(5011) <= not((layer0_outputs(5748)) and (layer0_outputs(10040)));
    layer1_outputs(5012) <= layer0_outputs(11387);
    layer1_outputs(5013) <= not(layer0_outputs(7339));
    layer1_outputs(5014) <= not(layer0_outputs(9264)) or (layer0_outputs(400));
    layer1_outputs(5015) <= not(layer0_outputs(2197));
    layer1_outputs(5016) <= (layer0_outputs(8823)) and (layer0_outputs(2301));
    layer1_outputs(5017) <= (layer0_outputs(11345)) and not (layer0_outputs(7318));
    layer1_outputs(5018) <= not((layer0_outputs(12399)) and (layer0_outputs(5763)));
    layer1_outputs(5019) <= layer0_outputs(12168);
    layer1_outputs(5020) <= not(layer0_outputs(6564)) or (layer0_outputs(391));
    layer1_outputs(5021) <= layer0_outputs(10287);
    layer1_outputs(5022) <= (layer0_outputs(11804)) and (layer0_outputs(6470));
    layer1_outputs(5023) <= layer0_outputs(10201);
    layer1_outputs(5024) <= layer0_outputs(1575);
    layer1_outputs(5025) <= not(layer0_outputs(7029)) or (layer0_outputs(7878));
    layer1_outputs(5026) <= not(layer0_outputs(8037)) or (layer0_outputs(6942));
    layer1_outputs(5027) <= (layer0_outputs(2277)) or (layer0_outputs(8262));
    layer1_outputs(5028) <= not((layer0_outputs(4325)) or (layer0_outputs(8132)));
    layer1_outputs(5029) <= '0';
    layer1_outputs(5030) <= not(layer0_outputs(6766)) or (layer0_outputs(12172));
    layer1_outputs(5031) <= not(layer0_outputs(9689));
    layer1_outputs(5032) <= (layer0_outputs(6167)) or (layer0_outputs(4269));
    layer1_outputs(5033) <= layer0_outputs(4945);
    layer1_outputs(5034) <= not((layer0_outputs(11464)) or (layer0_outputs(2646)));
    layer1_outputs(5035) <= layer0_outputs(2212);
    layer1_outputs(5036) <= (layer0_outputs(7275)) and (layer0_outputs(5378));
    layer1_outputs(5037) <= (layer0_outputs(12366)) and not (layer0_outputs(1171));
    layer1_outputs(5038) <= (layer0_outputs(11288)) xor (layer0_outputs(565));
    layer1_outputs(5039) <= not((layer0_outputs(2294)) xor (layer0_outputs(5204)));
    layer1_outputs(5040) <= (layer0_outputs(4116)) and not (layer0_outputs(8886));
    layer1_outputs(5041) <= not(layer0_outputs(10192)) or (layer0_outputs(7466));
    layer1_outputs(5042) <= layer0_outputs(6127);
    layer1_outputs(5043) <= (layer0_outputs(982)) and not (layer0_outputs(6470));
    layer1_outputs(5044) <= layer0_outputs(3821);
    layer1_outputs(5045) <= not((layer0_outputs(10352)) or (layer0_outputs(1278)));
    layer1_outputs(5046) <= '0';
    layer1_outputs(5047) <= not((layer0_outputs(12573)) xor (layer0_outputs(3491)));
    layer1_outputs(5048) <= not((layer0_outputs(3689)) or (layer0_outputs(3416)));
    layer1_outputs(5049) <= not((layer0_outputs(8644)) or (layer0_outputs(11538)));
    layer1_outputs(5050) <= (layer0_outputs(3569)) and (layer0_outputs(7117));
    layer1_outputs(5051) <= layer0_outputs(5464);
    layer1_outputs(5052) <= (layer0_outputs(230)) and not (layer0_outputs(11931));
    layer1_outputs(5053) <= not((layer0_outputs(8118)) or (layer0_outputs(8)));
    layer1_outputs(5054) <= (layer0_outputs(3800)) or (layer0_outputs(6011));
    layer1_outputs(5055) <= (layer0_outputs(10902)) and (layer0_outputs(7732));
    layer1_outputs(5056) <= (layer0_outputs(3619)) and (layer0_outputs(5358));
    layer1_outputs(5057) <= not(layer0_outputs(4265)) or (layer0_outputs(2211));
    layer1_outputs(5058) <= not(layer0_outputs(11428));
    layer1_outputs(5059) <= (layer0_outputs(8416)) and (layer0_outputs(152));
    layer1_outputs(5060) <= not(layer0_outputs(5335)) or (layer0_outputs(1390));
    layer1_outputs(5061) <= not(layer0_outputs(10095)) or (layer0_outputs(6885));
    layer1_outputs(5062) <= layer0_outputs(9372);
    layer1_outputs(5063) <= (layer0_outputs(7714)) and not (layer0_outputs(689));
    layer1_outputs(5064) <= '1';
    layer1_outputs(5065) <= layer0_outputs(3804);
    layer1_outputs(5066) <= not(layer0_outputs(10153)) or (layer0_outputs(252));
    layer1_outputs(5067) <= (layer0_outputs(10273)) and not (layer0_outputs(5284));
    layer1_outputs(5068) <= (layer0_outputs(2957)) and (layer0_outputs(8933));
    layer1_outputs(5069) <= not(layer0_outputs(12167));
    layer1_outputs(5070) <= not(layer0_outputs(5458)) or (layer0_outputs(5980));
    layer1_outputs(5071) <= (layer0_outputs(7238)) and not (layer0_outputs(4373));
    layer1_outputs(5072) <= (layer0_outputs(835)) and not (layer0_outputs(9579));
    layer1_outputs(5073) <= layer0_outputs(6854);
    layer1_outputs(5074) <= not(layer0_outputs(11377)) or (layer0_outputs(1863));
    layer1_outputs(5075) <= (layer0_outputs(7932)) and not (layer0_outputs(5200));
    layer1_outputs(5076) <= layer0_outputs(2346);
    layer1_outputs(5077) <= (layer0_outputs(9956)) or (layer0_outputs(1308));
    layer1_outputs(5078) <= (layer0_outputs(4247)) and not (layer0_outputs(103));
    layer1_outputs(5079) <= not(layer0_outputs(11003)) or (layer0_outputs(6796));
    layer1_outputs(5080) <= (layer0_outputs(3295)) and not (layer0_outputs(3877));
    layer1_outputs(5081) <= not(layer0_outputs(8112)) or (layer0_outputs(6065));
    layer1_outputs(5082) <= layer0_outputs(4275);
    layer1_outputs(5083) <= not((layer0_outputs(1165)) and (layer0_outputs(4454)));
    layer1_outputs(5084) <= not(layer0_outputs(6377));
    layer1_outputs(5085) <= (layer0_outputs(4161)) and not (layer0_outputs(9708));
    layer1_outputs(5086) <= not((layer0_outputs(10060)) xor (layer0_outputs(784)));
    layer1_outputs(5087) <= not((layer0_outputs(9143)) and (layer0_outputs(3513)));
    layer1_outputs(5088) <= layer0_outputs(3103);
    layer1_outputs(5089) <= (layer0_outputs(550)) and not (layer0_outputs(11435));
    layer1_outputs(5090) <= '0';
    layer1_outputs(5091) <= layer0_outputs(6643);
    layer1_outputs(5092) <= (layer0_outputs(7968)) or (layer0_outputs(422));
    layer1_outputs(5093) <= (layer0_outputs(4815)) or (layer0_outputs(9161));
    layer1_outputs(5094) <= (layer0_outputs(6263)) and not (layer0_outputs(3172));
    layer1_outputs(5095) <= not(layer0_outputs(4527));
    layer1_outputs(5096) <= not(layer0_outputs(5799));
    layer1_outputs(5097) <= (layer0_outputs(3264)) and (layer0_outputs(6701));
    layer1_outputs(5098) <= not(layer0_outputs(8263));
    layer1_outputs(5099) <= not(layer0_outputs(4251)) or (layer0_outputs(1476));
    layer1_outputs(5100) <= not((layer0_outputs(425)) or (layer0_outputs(7524)));
    layer1_outputs(5101) <= not(layer0_outputs(3614)) or (layer0_outputs(2755));
    layer1_outputs(5102) <= '1';
    layer1_outputs(5103) <= not(layer0_outputs(8834));
    layer1_outputs(5104) <= not(layer0_outputs(7195));
    layer1_outputs(5105) <= (layer0_outputs(4751)) and not (layer0_outputs(2844));
    layer1_outputs(5106) <= (layer0_outputs(2395)) and (layer0_outputs(5601));
    layer1_outputs(5107) <= layer0_outputs(293);
    layer1_outputs(5108) <= layer0_outputs(4094);
    layer1_outputs(5109) <= (layer0_outputs(1550)) or (layer0_outputs(2557));
    layer1_outputs(5110) <= (layer0_outputs(11171)) and (layer0_outputs(6350));
    layer1_outputs(5111) <= (layer0_outputs(5961)) or (layer0_outputs(10102));
    layer1_outputs(5112) <= (layer0_outputs(4820)) and (layer0_outputs(520));
    layer1_outputs(5113) <= '0';
    layer1_outputs(5114) <= not(layer0_outputs(4512)) or (layer0_outputs(5869));
    layer1_outputs(5115) <= not((layer0_outputs(2272)) xor (layer0_outputs(1451)));
    layer1_outputs(5116) <= not((layer0_outputs(1469)) or (layer0_outputs(7019)));
    layer1_outputs(5117) <= not(layer0_outputs(6608)) or (layer0_outputs(12622));
    layer1_outputs(5118) <= not(layer0_outputs(1941));
    layer1_outputs(5119) <= (layer0_outputs(5692)) or (layer0_outputs(11188));
    layer1_outputs(5120) <= (layer0_outputs(6024)) and (layer0_outputs(9898));
    layer1_outputs(5121) <= not(layer0_outputs(4521));
    layer1_outputs(5122) <= not(layer0_outputs(2415));
    layer1_outputs(5123) <= (layer0_outputs(7970)) and (layer0_outputs(4207));
    layer1_outputs(5124) <= not(layer0_outputs(670));
    layer1_outputs(5125) <= not((layer0_outputs(3462)) and (layer0_outputs(11454)));
    layer1_outputs(5126) <= not((layer0_outputs(7719)) and (layer0_outputs(1443)));
    layer1_outputs(5127) <= layer0_outputs(4382);
    layer1_outputs(5128) <= not(layer0_outputs(7841)) or (layer0_outputs(3775));
    layer1_outputs(5129) <= not(layer0_outputs(12481));
    layer1_outputs(5130) <= (layer0_outputs(2932)) and (layer0_outputs(11455));
    layer1_outputs(5131) <= (layer0_outputs(4112)) xor (layer0_outputs(2073));
    layer1_outputs(5132) <= layer0_outputs(5650);
    layer1_outputs(5133) <= (layer0_outputs(4268)) and not (layer0_outputs(4556));
    layer1_outputs(5134) <= not(layer0_outputs(12713));
    layer1_outputs(5135) <= (layer0_outputs(3806)) and not (layer0_outputs(2352));
    layer1_outputs(5136) <= not((layer0_outputs(3222)) and (layer0_outputs(2673)));
    layer1_outputs(5137) <= (layer0_outputs(1053)) or (layer0_outputs(12623));
    layer1_outputs(5138) <= (layer0_outputs(8641)) and not (layer0_outputs(11722));
    layer1_outputs(5139) <= (layer0_outputs(1793)) or (layer0_outputs(12050));
    layer1_outputs(5140) <= not((layer0_outputs(9497)) or (layer0_outputs(4234)));
    layer1_outputs(5141) <= not(layer0_outputs(9819));
    layer1_outputs(5142) <= (layer0_outputs(4748)) and (layer0_outputs(1416));
    layer1_outputs(5143) <= (layer0_outputs(6269)) and (layer0_outputs(387));
    layer1_outputs(5144) <= (layer0_outputs(1198)) or (layer0_outputs(4201));
    layer1_outputs(5145) <= not(layer0_outputs(6385)) or (layer0_outputs(2241));
    layer1_outputs(5146) <= not(layer0_outputs(7922));
    layer1_outputs(5147) <= layer0_outputs(161);
    layer1_outputs(5148) <= layer0_outputs(8544);
    layer1_outputs(5149) <= layer0_outputs(4923);
    layer1_outputs(5150) <= (layer0_outputs(12548)) and not (layer0_outputs(4384));
    layer1_outputs(5151) <= '0';
    layer1_outputs(5152) <= layer0_outputs(10473);
    layer1_outputs(5153) <= (layer0_outputs(10320)) and not (layer0_outputs(10184));
    layer1_outputs(5154) <= (layer0_outputs(4642)) and not (layer0_outputs(1137));
    layer1_outputs(5155) <= layer0_outputs(6237);
    layer1_outputs(5156) <= not(layer0_outputs(10436));
    layer1_outputs(5157) <= layer0_outputs(11357);
    layer1_outputs(5158) <= (layer0_outputs(11795)) xor (layer0_outputs(8298));
    layer1_outputs(5159) <= (layer0_outputs(8057)) or (layer0_outputs(7954));
    layer1_outputs(5160) <= not((layer0_outputs(11684)) and (layer0_outputs(1448)));
    layer1_outputs(5161) <= not((layer0_outputs(10409)) or (layer0_outputs(4140)));
    layer1_outputs(5162) <= (layer0_outputs(5974)) and (layer0_outputs(11417));
    layer1_outputs(5163) <= not(layer0_outputs(3138));
    layer1_outputs(5164) <= not((layer0_outputs(10523)) or (layer0_outputs(10894)));
    layer1_outputs(5165) <= layer0_outputs(9974);
    layer1_outputs(5166) <= (layer0_outputs(4409)) and (layer0_outputs(10192));
    layer1_outputs(5167) <= (layer0_outputs(4529)) or (layer0_outputs(4879));
    layer1_outputs(5168) <= (layer0_outputs(8658)) and not (layer0_outputs(8337));
    layer1_outputs(5169) <= not(layer0_outputs(5968));
    layer1_outputs(5170) <= not(layer0_outputs(7905));
    layer1_outputs(5171) <= not((layer0_outputs(3921)) and (layer0_outputs(11901)));
    layer1_outputs(5172) <= not(layer0_outputs(10648)) or (layer0_outputs(2830));
    layer1_outputs(5173) <= (layer0_outputs(8174)) xor (layer0_outputs(5958));
    layer1_outputs(5174) <= layer0_outputs(6798);
    layer1_outputs(5175) <= not(layer0_outputs(1648));
    layer1_outputs(5176) <= (layer0_outputs(4883)) or (layer0_outputs(6830));
    layer1_outputs(5177) <= not(layer0_outputs(8789)) or (layer0_outputs(1272));
    layer1_outputs(5178) <= not((layer0_outputs(2623)) or (layer0_outputs(274)));
    layer1_outputs(5179) <= not((layer0_outputs(8429)) or (layer0_outputs(1271)));
    layer1_outputs(5180) <= not((layer0_outputs(2624)) and (layer0_outputs(5540)));
    layer1_outputs(5181) <= layer0_outputs(9016);
    layer1_outputs(5182) <= (layer0_outputs(8941)) and not (layer0_outputs(6906));
    layer1_outputs(5183) <= not(layer0_outputs(765)) or (layer0_outputs(10809));
    layer1_outputs(5184) <= not(layer0_outputs(6383));
    layer1_outputs(5185) <= layer0_outputs(1512);
    layer1_outputs(5186) <= not((layer0_outputs(2870)) xor (layer0_outputs(7521)));
    layer1_outputs(5187) <= not(layer0_outputs(7497));
    layer1_outputs(5188) <= not(layer0_outputs(5816)) or (layer0_outputs(8771));
    layer1_outputs(5189) <= not(layer0_outputs(8884));
    layer1_outputs(5190) <= (layer0_outputs(492)) or (layer0_outputs(12486));
    layer1_outputs(5191) <= not(layer0_outputs(7869)) or (layer0_outputs(11977));
    layer1_outputs(5192) <= '0';
    layer1_outputs(5193) <= '1';
    layer1_outputs(5194) <= not(layer0_outputs(3087)) or (layer0_outputs(10440));
    layer1_outputs(5195) <= not(layer0_outputs(1035));
    layer1_outputs(5196) <= (layer0_outputs(6514)) xor (layer0_outputs(8393));
    layer1_outputs(5197) <= not(layer0_outputs(4080));
    layer1_outputs(5198) <= (layer0_outputs(11550)) and (layer0_outputs(9396));
    layer1_outputs(5199) <= layer0_outputs(5504);
    layer1_outputs(5200) <= layer0_outputs(6863);
    layer1_outputs(5201) <= not(layer0_outputs(8278));
    layer1_outputs(5202) <= (layer0_outputs(498)) and (layer0_outputs(5169));
    layer1_outputs(5203) <= (layer0_outputs(683)) and not (layer0_outputs(5858));
    layer1_outputs(5204) <= not((layer0_outputs(7478)) and (layer0_outputs(2969)));
    layer1_outputs(5205) <= (layer0_outputs(4158)) and not (layer0_outputs(2173));
    layer1_outputs(5206) <= layer0_outputs(7001);
    layer1_outputs(5207) <= (layer0_outputs(199)) and not (layer0_outputs(5151));
    layer1_outputs(5208) <= not((layer0_outputs(12267)) xor (layer0_outputs(3642)));
    layer1_outputs(5209) <= not(layer0_outputs(1244));
    layer1_outputs(5210) <= not((layer0_outputs(9817)) or (layer0_outputs(5058)));
    layer1_outputs(5211) <= not((layer0_outputs(7701)) or (layer0_outputs(11625)));
    layer1_outputs(5212) <= not((layer0_outputs(9884)) or (layer0_outputs(10508)));
    layer1_outputs(5213) <= not(layer0_outputs(11827));
    layer1_outputs(5214) <= layer0_outputs(286);
    layer1_outputs(5215) <= layer0_outputs(11159);
    layer1_outputs(5216) <= (layer0_outputs(12389)) or (layer0_outputs(12300));
    layer1_outputs(5217) <= not(layer0_outputs(2520)) or (layer0_outputs(2864));
    layer1_outputs(5218) <= (layer0_outputs(12304)) xor (layer0_outputs(10389));
    layer1_outputs(5219) <= not(layer0_outputs(7454));
    layer1_outputs(5220) <= not(layer0_outputs(12346));
    layer1_outputs(5221) <= not(layer0_outputs(5385)) or (layer0_outputs(467));
    layer1_outputs(5222) <= not(layer0_outputs(10122)) or (layer0_outputs(5460));
    layer1_outputs(5223) <= (layer0_outputs(9500)) or (layer0_outputs(7557));
    layer1_outputs(5224) <= not(layer0_outputs(9817));
    layer1_outputs(5225) <= '1';
    layer1_outputs(5226) <= not(layer0_outputs(1206));
    layer1_outputs(5227) <= not((layer0_outputs(9068)) or (layer0_outputs(9125)));
    layer1_outputs(5228) <= (layer0_outputs(6335)) and not (layer0_outputs(12206));
    layer1_outputs(5229) <= not(layer0_outputs(10471)) or (layer0_outputs(8252));
    layer1_outputs(5230) <= not(layer0_outputs(2480));
    layer1_outputs(5231) <= not(layer0_outputs(2593));
    layer1_outputs(5232) <= layer0_outputs(1879);
    layer1_outputs(5233) <= layer0_outputs(4191);
    layer1_outputs(5234) <= (layer0_outputs(7006)) xor (layer0_outputs(11143));
    layer1_outputs(5235) <= layer0_outputs(12079);
    layer1_outputs(5236) <= layer0_outputs(12273);
    layer1_outputs(5237) <= not(layer0_outputs(9943)) or (layer0_outputs(375));
    layer1_outputs(5238) <= not(layer0_outputs(7987));
    layer1_outputs(5239) <= not(layer0_outputs(9070));
    layer1_outputs(5240) <= (layer0_outputs(1556)) and not (layer0_outputs(2975));
    layer1_outputs(5241) <= layer0_outputs(262);
    layer1_outputs(5242) <= (layer0_outputs(4242)) and not (layer0_outputs(9767));
    layer1_outputs(5243) <= layer0_outputs(3780);
    layer1_outputs(5244) <= not((layer0_outputs(9674)) and (layer0_outputs(7187)));
    layer1_outputs(5245) <= not(layer0_outputs(10987));
    layer1_outputs(5246) <= not((layer0_outputs(10064)) xor (layer0_outputs(2796)));
    layer1_outputs(5247) <= not(layer0_outputs(3204)) or (layer0_outputs(3212));
    layer1_outputs(5248) <= not(layer0_outputs(9498));
    layer1_outputs(5249) <= not(layer0_outputs(11658)) or (layer0_outputs(10620));
    layer1_outputs(5250) <= not(layer0_outputs(9812)) or (layer0_outputs(9325));
    layer1_outputs(5251) <= not(layer0_outputs(9019)) or (layer0_outputs(1455));
    layer1_outputs(5252) <= not((layer0_outputs(6876)) or (layer0_outputs(12445)));
    layer1_outputs(5253) <= not(layer0_outputs(10854));
    layer1_outputs(5254) <= not(layer0_outputs(1633)) or (layer0_outputs(1399));
    layer1_outputs(5255) <= not(layer0_outputs(11366));
    layer1_outputs(5256) <= (layer0_outputs(5363)) or (layer0_outputs(9830));
    layer1_outputs(5257) <= not(layer0_outputs(11681)) or (layer0_outputs(10377));
    layer1_outputs(5258) <= '1';
    layer1_outputs(5259) <= not(layer0_outputs(7375)) or (layer0_outputs(7211));
    layer1_outputs(5260) <= (layer0_outputs(254)) and not (layer0_outputs(382));
    layer1_outputs(5261) <= not(layer0_outputs(86));
    layer1_outputs(5262) <= not((layer0_outputs(2195)) or (layer0_outputs(5942)));
    layer1_outputs(5263) <= not((layer0_outputs(2453)) and (layer0_outputs(2301)));
    layer1_outputs(5264) <= (layer0_outputs(1841)) xor (layer0_outputs(11585));
    layer1_outputs(5265) <= (layer0_outputs(11872)) xor (layer0_outputs(2787));
    layer1_outputs(5266) <= (layer0_outputs(11156)) xor (layer0_outputs(9504));
    layer1_outputs(5267) <= not(layer0_outputs(665));
    layer1_outputs(5268) <= (layer0_outputs(10556)) and not (layer0_outputs(7989));
    layer1_outputs(5269) <= not(layer0_outputs(9624));
    layer1_outputs(5270) <= (layer0_outputs(2464)) and not (layer0_outputs(3366));
    layer1_outputs(5271) <= layer0_outputs(585);
    layer1_outputs(5272) <= not(layer0_outputs(360)) or (layer0_outputs(567));
    layer1_outputs(5273) <= (layer0_outputs(5745)) and not (layer0_outputs(12206));
    layer1_outputs(5274) <= not(layer0_outputs(7705));
    layer1_outputs(5275) <= not(layer0_outputs(10276)) or (layer0_outputs(5657));
    layer1_outputs(5276) <= layer0_outputs(6851);
    layer1_outputs(5277) <= not(layer0_outputs(4557));
    layer1_outputs(5278) <= layer0_outputs(4672);
    layer1_outputs(5279) <= layer0_outputs(3064);
    layer1_outputs(5280) <= not(layer0_outputs(12210));
    layer1_outputs(5281) <= layer0_outputs(7395);
    layer1_outputs(5282) <= not(layer0_outputs(7368)) or (layer0_outputs(4082));
    layer1_outputs(5283) <= '0';
    layer1_outputs(5284) <= not(layer0_outputs(2067)) or (layer0_outputs(2464));
    layer1_outputs(5285) <= not(layer0_outputs(5796));
    layer1_outputs(5286) <= not(layer0_outputs(12023)) or (layer0_outputs(8935));
    layer1_outputs(5287) <= layer0_outputs(6486);
    layer1_outputs(5288) <= layer0_outputs(8212);
    layer1_outputs(5289) <= layer0_outputs(7240);
    layer1_outputs(5290) <= '1';
    layer1_outputs(5291) <= layer0_outputs(11544);
    layer1_outputs(5292) <= not(layer0_outputs(1606)) or (layer0_outputs(10142));
    layer1_outputs(5293) <= not(layer0_outputs(2910));
    layer1_outputs(5294) <= not((layer0_outputs(7002)) or (layer0_outputs(5507)));
    layer1_outputs(5295) <= not((layer0_outputs(10883)) xor (layer0_outputs(10895)));
    layer1_outputs(5296) <= (layer0_outputs(7589)) xor (layer0_outputs(8337));
    layer1_outputs(5297) <= not((layer0_outputs(3074)) or (layer0_outputs(6934)));
    layer1_outputs(5298) <= not(layer0_outputs(1733));
    layer1_outputs(5299) <= not(layer0_outputs(9921)) or (layer0_outputs(11916));
    layer1_outputs(5300) <= not(layer0_outputs(304));
    layer1_outputs(5301) <= (layer0_outputs(5225)) and not (layer0_outputs(9482));
    layer1_outputs(5302) <= not((layer0_outputs(7543)) xor (layer0_outputs(12242)));
    layer1_outputs(5303) <= not(layer0_outputs(5020)) or (layer0_outputs(5109));
    layer1_outputs(5304) <= (layer0_outputs(2378)) and not (layer0_outputs(2542));
    layer1_outputs(5305) <= layer0_outputs(12497);
    layer1_outputs(5306) <= not(layer0_outputs(10131));
    layer1_outputs(5307) <= (layer0_outputs(8909)) and not (layer0_outputs(5860));
    layer1_outputs(5308) <= layer0_outputs(8245);
    layer1_outputs(5309) <= layer0_outputs(6543);
    layer1_outputs(5310) <= (layer0_outputs(299)) and not (layer0_outputs(1238));
    layer1_outputs(5311) <= layer0_outputs(1448);
    layer1_outputs(5312) <= not(layer0_outputs(5999));
    layer1_outputs(5313) <= (layer0_outputs(9569)) xor (layer0_outputs(8797));
    layer1_outputs(5314) <= not(layer0_outputs(7481)) or (layer0_outputs(12762));
    layer1_outputs(5315) <= not(layer0_outputs(3283)) or (layer0_outputs(8038));
    layer1_outputs(5316) <= (layer0_outputs(3174)) xor (layer0_outputs(8708));
    layer1_outputs(5317) <= not(layer0_outputs(8822));
    layer1_outputs(5318) <= not(layer0_outputs(6414));
    layer1_outputs(5319) <= layer0_outputs(1426);
    layer1_outputs(5320) <= not(layer0_outputs(6152));
    layer1_outputs(5321) <= (layer0_outputs(7601)) or (layer0_outputs(7963));
    layer1_outputs(5322) <= (layer0_outputs(5763)) and not (layer0_outputs(9982));
    layer1_outputs(5323) <= '0';
    layer1_outputs(5324) <= layer0_outputs(4802);
    layer1_outputs(5325) <= not((layer0_outputs(773)) and (layer0_outputs(11509)));
    layer1_outputs(5326) <= not(layer0_outputs(11666));
    layer1_outputs(5327) <= (layer0_outputs(2206)) or (layer0_outputs(11712));
    layer1_outputs(5328) <= not(layer0_outputs(182));
    layer1_outputs(5329) <= (layer0_outputs(10261)) and (layer0_outputs(10995));
    layer1_outputs(5330) <= (layer0_outputs(3208)) or (layer0_outputs(5921));
    layer1_outputs(5331) <= (layer0_outputs(5958)) and not (layer0_outputs(7373));
    layer1_outputs(5332) <= not(layer0_outputs(2182)) or (layer0_outputs(1587));
    layer1_outputs(5333) <= not((layer0_outputs(4475)) or (layer0_outputs(5799)));
    layer1_outputs(5334) <= layer0_outputs(1585);
    layer1_outputs(5335) <= layer0_outputs(10633);
    layer1_outputs(5336) <= not(layer0_outputs(7309));
    layer1_outputs(5337) <= (layer0_outputs(8649)) and not (layer0_outputs(12724));
    layer1_outputs(5338) <= layer0_outputs(7350);
    layer1_outputs(5339) <= '1';
    layer1_outputs(5340) <= not((layer0_outputs(6649)) or (layer0_outputs(6547)));
    layer1_outputs(5341) <= layer0_outputs(4984);
    layer1_outputs(5342) <= (layer0_outputs(11575)) xor (layer0_outputs(6859));
    layer1_outputs(5343) <= layer0_outputs(939);
    layer1_outputs(5344) <= not((layer0_outputs(1033)) and (layer0_outputs(8610)));
    layer1_outputs(5345) <= layer0_outputs(6435);
    layer1_outputs(5346) <= layer0_outputs(5330);
    layer1_outputs(5347) <= not(layer0_outputs(3439));
    layer1_outputs(5348) <= not(layer0_outputs(6611));
    layer1_outputs(5349) <= layer0_outputs(4333);
    layer1_outputs(5350) <= (layer0_outputs(10009)) and (layer0_outputs(7842));
    layer1_outputs(5351) <= layer0_outputs(7008);
    layer1_outputs(5352) <= layer0_outputs(8182);
    layer1_outputs(5353) <= layer0_outputs(10822);
    layer1_outputs(5354) <= '0';
    layer1_outputs(5355) <= not(layer0_outputs(5081));
    layer1_outputs(5356) <= not(layer0_outputs(10275));
    layer1_outputs(5357) <= layer0_outputs(781);
    layer1_outputs(5358) <= (layer0_outputs(8074)) and not (layer0_outputs(2667));
    layer1_outputs(5359) <= (layer0_outputs(12061)) and not (layer0_outputs(7131));
    layer1_outputs(5360) <= (layer0_outputs(8788)) or (layer0_outputs(3639));
    layer1_outputs(5361) <= layer0_outputs(7939);
    layer1_outputs(5362) <= not((layer0_outputs(6240)) or (layer0_outputs(9089)));
    layer1_outputs(5363) <= not(layer0_outputs(8223));
    layer1_outputs(5364) <= layer0_outputs(5309);
    layer1_outputs(5365) <= layer0_outputs(7133);
    layer1_outputs(5366) <= not(layer0_outputs(6527));
    layer1_outputs(5367) <= not(layer0_outputs(11297)) or (layer0_outputs(8806));
    layer1_outputs(5368) <= (layer0_outputs(1099)) and (layer0_outputs(6684));
    layer1_outputs(5369) <= not(layer0_outputs(3963));
    layer1_outputs(5370) <= layer0_outputs(1977);
    layer1_outputs(5371) <= not(layer0_outputs(1743));
    layer1_outputs(5372) <= not((layer0_outputs(3328)) or (layer0_outputs(7649)));
    layer1_outputs(5373) <= not((layer0_outputs(11284)) or (layer0_outputs(6792)));
    layer1_outputs(5374) <= not(layer0_outputs(1192));
    layer1_outputs(5375) <= (layer0_outputs(7368)) xor (layer0_outputs(9298));
    layer1_outputs(5376) <= not(layer0_outputs(6760));
    layer1_outputs(5377) <= not(layer0_outputs(1827)) or (layer0_outputs(5235));
    layer1_outputs(5378) <= not((layer0_outputs(4396)) or (layer0_outputs(1040)));
    layer1_outputs(5379) <= layer0_outputs(10004);
    layer1_outputs(5380) <= (layer0_outputs(9160)) xor (layer0_outputs(7161));
    layer1_outputs(5381) <= layer0_outputs(1924);
    layer1_outputs(5382) <= layer0_outputs(2777);
    layer1_outputs(5383) <= not(layer0_outputs(4355));
    layer1_outputs(5384) <= not(layer0_outputs(10886)) or (layer0_outputs(6147));
    layer1_outputs(5385) <= not((layer0_outputs(2275)) or (layer0_outputs(10850)));
    layer1_outputs(5386) <= not(layer0_outputs(8181)) or (layer0_outputs(10829));
    layer1_outputs(5387) <= not(layer0_outputs(11350)) or (layer0_outputs(6292));
    layer1_outputs(5388) <= layer0_outputs(11186);
    layer1_outputs(5389) <= layer0_outputs(12690);
    layer1_outputs(5390) <= (layer0_outputs(10454)) and (layer0_outputs(11699));
    layer1_outputs(5391) <= not((layer0_outputs(10228)) and (layer0_outputs(512)));
    layer1_outputs(5392) <= layer0_outputs(4441);
    layer1_outputs(5393) <= not(layer0_outputs(6408)) or (layer0_outputs(5859));
    layer1_outputs(5394) <= not((layer0_outputs(4193)) and (layer0_outputs(3414)));
    layer1_outputs(5395) <= (layer0_outputs(8026)) and not (layer0_outputs(10364));
    layer1_outputs(5396) <= not((layer0_outputs(5279)) and (layer0_outputs(4091)));
    layer1_outputs(5397) <= not(layer0_outputs(5101));
    layer1_outputs(5398) <= (layer0_outputs(888)) xor (layer0_outputs(388));
    layer1_outputs(5399) <= layer0_outputs(11957);
    layer1_outputs(5400) <= not(layer0_outputs(10558));
    layer1_outputs(5401) <= layer0_outputs(2379);
    layer1_outputs(5402) <= layer0_outputs(9465);
    layer1_outputs(5403) <= not((layer0_outputs(4292)) or (layer0_outputs(12672)));
    layer1_outputs(5404) <= layer0_outputs(5639);
    layer1_outputs(5405) <= layer0_outputs(6219);
    layer1_outputs(5406) <= (layer0_outputs(9983)) or (layer0_outputs(5106));
    layer1_outputs(5407) <= not(layer0_outputs(10687)) or (layer0_outputs(4517));
    layer1_outputs(5408) <= not(layer0_outputs(5197));
    layer1_outputs(5409) <= layer0_outputs(6981);
    layer1_outputs(5410) <= not(layer0_outputs(828)) or (layer0_outputs(4079));
    layer1_outputs(5411) <= layer0_outputs(5091);
    layer1_outputs(5412) <= not(layer0_outputs(9773));
    layer1_outputs(5413) <= '0';
    layer1_outputs(5414) <= not((layer0_outputs(510)) or (layer0_outputs(4296)));
    layer1_outputs(5415) <= (layer0_outputs(10848)) and (layer0_outputs(7700));
    layer1_outputs(5416) <= '1';
    layer1_outputs(5417) <= not(layer0_outputs(7075));
    layer1_outputs(5418) <= not(layer0_outputs(4684));
    layer1_outputs(5419) <= '1';
    layer1_outputs(5420) <= not(layer0_outputs(8313));
    layer1_outputs(5421) <= (layer0_outputs(12194)) and (layer0_outputs(1587));
    layer1_outputs(5422) <= not(layer0_outputs(6728)) or (layer0_outputs(5841));
    layer1_outputs(5423) <= not((layer0_outputs(9142)) and (layer0_outputs(5401)));
    layer1_outputs(5424) <= layer0_outputs(6049);
    layer1_outputs(5425) <= not(layer0_outputs(7020));
    layer1_outputs(5426) <= layer0_outputs(10867);
    layer1_outputs(5427) <= not(layer0_outputs(843)) or (layer0_outputs(4069));
    layer1_outputs(5428) <= layer0_outputs(9392);
    layer1_outputs(5429) <= layer0_outputs(4134);
    layer1_outputs(5430) <= (layer0_outputs(7267)) and not (layer0_outputs(10575));
    layer1_outputs(5431) <= not(layer0_outputs(10567));
    layer1_outputs(5432) <= '1';
    layer1_outputs(5433) <= layer0_outputs(6019);
    layer1_outputs(5434) <= not(layer0_outputs(1216));
    layer1_outputs(5435) <= not((layer0_outputs(4677)) and (layer0_outputs(7140)));
    layer1_outputs(5436) <= layer0_outputs(1928);
    layer1_outputs(5437) <= not((layer0_outputs(6767)) and (layer0_outputs(1048)));
    layer1_outputs(5438) <= not(layer0_outputs(11783)) or (layer0_outputs(5000));
    layer1_outputs(5439) <= not((layer0_outputs(5899)) xor (layer0_outputs(3757)));
    layer1_outputs(5440) <= (layer0_outputs(9913)) and not (layer0_outputs(6592));
    layer1_outputs(5441) <= not(layer0_outputs(1474)) or (layer0_outputs(321));
    layer1_outputs(5442) <= not(layer0_outputs(4074));
    layer1_outputs(5443) <= not((layer0_outputs(2140)) xor (layer0_outputs(3102)));
    layer1_outputs(5444) <= (layer0_outputs(3126)) xor (layer0_outputs(1156));
    layer1_outputs(5445) <= not(layer0_outputs(10746)) or (layer0_outputs(6391));
    layer1_outputs(5446) <= not(layer0_outputs(5745)) or (layer0_outputs(4959));
    layer1_outputs(5447) <= layer0_outputs(10181);
    layer1_outputs(5448) <= (layer0_outputs(2200)) and not (layer0_outputs(490));
    layer1_outputs(5449) <= not(layer0_outputs(4999)) or (layer0_outputs(2131));
    layer1_outputs(5450) <= not(layer0_outputs(5374)) or (layer0_outputs(11708));
    layer1_outputs(5451) <= (layer0_outputs(2291)) and not (layer0_outputs(9201));
    layer1_outputs(5452) <= (layer0_outputs(758)) or (layer0_outputs(3152));
    layer1_outputs(5453) <= layer0_outputs(8039);
    layer1_outputs(5454) <= not(layer0_outputs(1560));
    layer1_outputs(5455) <= not(layer0_outputs(8409));
    layer1_outputs(5456) <= not(layer0_outputs(7891));
    layer1_outputs(5457) <= (layer0_outputs(3005)) xor (layer0_outputs(7459));
    layer1_outputs(5458) <= not(layer0_outputs(4280));
    layer1_outputs(5459) <= layer0_outputs(1073);
    layer1_outputs(5460) <= (layer0_outputs(11160)) and not (layer0_outputs(2788));
    layer1_outputs(5461) <= (layer0_outputs(9573)) xor (layer0_outputs(8575));
    layer1_outputs(5462) <= not((layer0_outputs(2674)) xor (layer0_outputs(3194)));
    layer1_outputs(5463) <= not(layer0_outputs(745));
    layer1_outputs(5464) <= layer0_outputs(6688);
    layer1_outputs(5465) <= not(layer0_outputs(12513));
    layer1_outputs(5466) <= (layer0_outputs(443)) and not (layer0_outputs(4899));
    layer1_outputs(5467) <= (layer0_outputs(8189)) and not (layer0_outputs(2434));
    layer1_outputs(5468) <= layer0_outputs(10270);
    layer1_outputs(5469) <= not(layer0_outputs(7192)) or (layer0_outputs(8127));
    layer1_outputs(5470) <= (layer0_outputs(6451)) and (layer0_outputs(2847));
    layer1_outputs(5471) <= layer0_outputs(3239);
    layer1_outputs(5472) <= layer0_outputs(4231);
    layer1_outputs(5473) <= (layer0_outputs(7995)) and not (layer0_outputs(8531));
    layer1_outputs(5474) <= not(layer0_outputs(3191)) or (layer0_outputs(2641));
    layer1_outputs(5475) <= layer0_outputs(1676);
    layer1_outputs(5476) <= not(layer0_outputs(1882));
    layer1_outputs(5477) <= not(layer0_outputs(7494));
    layer1_outputs(5478) <= (layer0_outputs(6785)) and not (layer0_outputs(7796));
    layer1_outputs(5479) <= '1';
    layer1_outputs(5480) <= not(layer0_outputs(1786)) or (layer0_outputs(8634));
    layer1_outputs(5481) <= not(layer0_outputs(12162)) or (layer0_outputs(11223));
    layer1_outputs(5482) <= (layer0_outputs(1695)) and not (layer0_outputs(1440));
    layer1_outputs(5483) <= (layer0_outputs(3880)) and not (layer0_outputs(1027));
    layer1_outputs(5484) <= not(layer0_outputs(1338)) or (layer0_outputs(3564));
    layer1_outputs(5485) <= layer0_outputs(5418);
    layer1_outputs(5486) <= (layer0_outputs(10306)) and not (layer0_outputs(2015));
    layer1_outputs(5487) <= not(layer0_outputs(864));
    layer1_outputs(5488) <= layer0_outputs(1965);
    layer1_outputs(5489) <= not((layer0_outputs(902)) or (layer0_outputs(11393)));
    layer1_outputs(5490) <= not(layer0_outputs(8377)) or (layer0_outputs(9993));
    layer1_outputs(5491) <= layer0_outputs(5155);
    layer1_outputs(5492) <= not(layer0_outputs(6407)) or (layer0_outputs(2442));
    layer1_outputs(5493) <= (layer0_outputs(1552)) and not (layer0_outputs(2899));
    layer1_outputs(5494) <= (layer0_outputs(8190)) and not (layer0_outputs(6939));
    layer1_outputs(5495) <= not(layer0_outputs(2400));
    layer1_outputs(5496) <= (layer0_outputs(11619)) and not (layer0_outputs(10977));
    layer1_outputs(5497) <= layer0_outputs(5444);
    layer1_outputs(5498) <= (layer0_outputs(2640)) and not (layer0_outputs(3050));
    layer1_outputs(5499) <= (layer0_outputs(11755)) and not (layer0_outputs(1369));
    layer1_outputs(5500) <= not(layer0_outputs(6951));
    layer1_outputs(5501) <= not(layer0_outputs(11530)) or (layer0_outputs(6623));
    layer1_outputs(5502) <= (layer0_outputs(915)) and not (layer0_outputs(3071));
    layer1_outputs(5503) <= not((layer0_outputs(2254)) and (layer0_outputs(5434)));
    layer1_outputs(5504) <= not((layer0_outputs(5586)) or (layer0_outputs(3669)));
    layer1_outputs(5505) <= not(layer0_outputs(12447));
    layer1_outputs(5506) <= not(layer0_outputs(2332)) or (layer0_outputs(3607));
    layer1_outputs(5507) <= (layer0_outputs(8034)) and not (layer0_outputs(10931));
    layer1_outputs(5508) <= layer0_outputs(3596);
    layer1_outputs(5509) <= (layer0_outputs(4657)) and not (layer0_outputs(4084));
    layer1_outputs(5510) <= (layer0_outputs(953)) or (layer0_outputs(6546));
    layer1_outputs(5511) <= (layer0_outputs(2550)) xor (layer0_outputs(1351));
    layer1_outputs(5512) <= layer0_outputs(12255);
    layer1_outputs(5513) <= not(layer0_outputs(2731));
    layer1_outputs(5514) <= not(layer0_outputs(11811)) or (layer0_outputs(3588));
    layer1_outputs(5515) <= layer0_outputs(12354);
    layer1_outputs(5516) <= layer0_outputs(7420);
    layer1_outputs(5517) <= layer0_outputs(10047);
    layer1_outputs(5518) <= not(layer0_outputs(5858)) or (layer0_outputs(4609));
    layer1_outputs(5519) <= (layer0_outputs(12457)) and (layer0_outputs(10236));
    layer1_outputs(5520) <= (layer0_outputs(3086)) or (layer0_outputs(911));
    layer1_outputs(5521) <= (layer0_outputs(9546)) and not (layer0_outputs(6116));
    layer1_outputs(5522) <= not((layer0_outputs(4839)) or (layer0_outputs(746)));
    layer1_outputs(5523) <= (layer0_outputs(1226)) or (layer0_outputs(6292));
    layer1_outputs(5524) <= not((layer0_outputs(8248)) xor (layer0_outputs(7958)));
    layer1_outputs(5525) <= not(layer0_outputs(6822));
    layer1_outputs(5526) <= layer0_outputs(8488);
    layer1_outputs(5527) <= not((layer0_outputs(6513)) and (layer0_outputs(5672)));
    layer1_outputs(5528) <= layer0_outputs(12322);
    layer1_outputs(5529) <= layer0_outputs(4566);
    layer1_outputs(5530) <= (layer0_outputs(4206)) or (layer0_outputs(5526));
    layer1_outputs(5531) <= layer0_outputs(5556);
    layer1_outputs(5532) <= not(layer0_outputs(11741));
    layer1_outputs(5533) <= (layer0_outputs(12410)) or (layer0_outputs(8045));
    layer1_outputs(5534) <= not(layer0_outputs(10699));
    layer1_outputs(5535) <= not(layer0_outputs(9509));
    layer1_outputs(5536) <= (layer0_outputs(8136)) xor (layer0_outputs(1603));
    layer1_outputs(5537) <= layer0_outputs(3438);
    layer1_outputs(5538) <= (layer0_outputs(8356)) and not (layer0_outputs(3148));
    layer1_outputs(5539) <= not(layer0_outputs(7408));
    layer1_outputs(5540) <= (layer0_outputs(12412)) and not (layer0_outputs(1245));
    layer1_outputs(5541) <= layer0_outputs(7400);
    layer1_outputs(5542) <= not(layer0_outputs(3314));
    layer1_outputs(5543) <= '1';
    layer1_outputs(5544) <= (layer0_outputs(1581)) xor (layer0_outputs(6591));
    layer1_outputs(5545) <= not(layer0_outputs(7090));
    layer1_outputs(5546) <= layer0_outputs(3341);
    layer1_outputs(5547) <= (layer0_outputs(8438)) or (layer0_outputs(5527));
    layer1_outputs(5548) <= layer0_outputs(1327);
    layer1_outputs(5549) <= (layer0_outputs(5348)) xor (layer0_outputs(1881));
    layer1_outputs(5550) <= not(layer0_outputs(5186));
    layer1_outputs(5551) <= not((layer0_outputs(2478)) or (layer0_outputs(11479)));
    layer1_outputs(5552) <= not((layer0_outputs(2498)) and (layer0_outputs(1163)));
    layer1_outputs(5553) <= '0';
    layer1_outputs(5554) <= (layer0_outputs(8508)) or (layer0_outputs(1150));
    layer1_outputs(5555) <= not((layer0_outputs(12090)) and (layer0_outputs(764)));
    layer1_outputs(5556) <= not((layer0_outputs(10916)) and (layer0_outputs(5323)));
    layer1_outputs(5557) <= '1';
    layer1_outputs(5558) <= not(layer0_outputs(10229));
    layer1_outputs(5559) <= not(layer0_outputs(1062)) or (layer0_outputs(11363));
    layer1_outputs(5560) <= layer0_outputs(6146);
    layer1_outputs(5561) <= not(layer0_outputs(11620)) or (layer0_outputs(3167));
    layer1_outputs(5562) <= not(layer0_outputs(2866)) or (layer0_outputs(12233));
    layer1_outputs(5563) <= layer0_outputs(7500);
    layer1_outputs(5564) <= (layer0_outputs(11848)) and not (layer0_outputs(8381));
    layer1_outputs(5565) <= not((layer0_outputs(383)) or (layer0_outputs(10698)));
    layer1_outputs(5566) <= (layer0_outputs(6321)) and (layer0_outputs(12190));
    layer1_outputs(5567) <= not((layer0_outputs(8014)) xor (layer0_outputs(8347)));
    layer1_outputs(5568) <= (layer0_outputs(6744)) and not (layer0_outputs(11076));
    layer1_outputs(5569) <= not(layer0_outputs(8408)) or (layer0_outputs(8129));
    layer1_outputs(5570) <= not(layer0_outputs(768));
    layer1_outputs(5571) <= not((layer0_outputs(11269)) and (layer0_outputs(12546)));
    layer1_outputs(5572) <= not((layer0_outputs(12689)) and (layer0_outputs(3702)));
    layer1_outputs(5573) <= not(layer0_outputs(12131));
    layer1_outputs(5574) <= (layer0_outputs(5266)) and (layer0_outputs(10407));
    layer1_outputs(5575) <= (layer0_outputs(10428)) or (layer0_outputs(2949));
    layer1_outputs(5576) <= layer0_outputs(7565);
    layer1_outputs(5577) <= not((layer0_outputs(6499)) xor (layer0_outputs(784)));
    layer1_outputs(5578) <= layer0_outputs(11477);
    layer1_outputs(5579) <= not((layer0_outputs(8822)) or (layer0_outputs(4252)));
    layer1_outputs(5580) <= not(layer0_outputs(10368)) or (layer0_outputs(12325));
    layer1_outputs(5581) <= layer0_outputs(5676);
    layer1_outputs(5582) <= not(layer0_outputs(6752)) or (layer0_outputs(7035));
    layer1_outputs(5583) <= layer0_outputs(12237);
    layer1_outputs(5584) <= not(layer0_outputs(11603));
    layer1_outputs(5585) <= '1';
    layer1_outputs(5586) <= (layer0_outputs(12381)) and not (layer0_outputs(11843));
    layer1_outputs(5587) <= not((layer0_outputs(11450)) and (layer0_outputs(1380)));
    layer1_outputs(5588) <= layer0_outputs(5060);
    layer1_outputs(5589) <= not(layer0_outputs(105));
    layer1_outputs(5590) <= layer0_outputs(12777);
    layer1_outputs(5591) <= layer0_outputs(8746);
    layer1_outputs(5592) <= '1';
    layer1_outputs(5593) <= (layer0_outputs(4939)) xor (layer0_outputs(8020));
    layer1_outputs(5594) <= not(layer0_outputs(11602));
    layer1_outputs(5595) <= (layer0_outputs(11099)) or (layer0_outputs(9193));
    layer1_outputs(5596) <= not(layer0_outputs(12783)) or (layer0_outputs(8628));
    layer1_outputs(5597) <= layer0_outputs(3377);
    layer1_outputs(5598) <= layer0_outputs(7488);
    layer1_outputs(5599) <= (layer0_outputs(104)) xor (layer0_outputs(8003));
    layer1_outputs(5600) <= not(layer0_outputs(4650));
    layer1_outputs(5601) <= not((layer0_outputs(6504)) and (layer0_outputs(5588)));
    layer1_outputs(5602) <= layer0_outputs(2775);
    layer1_outputs(5603) <= not(layer0_outputs(12368));
    layer1_outputs(5604) <= (layer0_outputs(5030)) and (layer0_outputs(3546));
    layer1_outputs(5605) <= not(layer0_outputs(1577));
    layer1_outputs(5606) <= layer0_outputs(10012);
    layer1_outputs(5607) <= layer0_outputs(1204);
    layer1_outputs(5608) <= not((layer0_outputs(8446)) xor (layer0_outputs(6441)));
    layer1_outputs(5609) <= layer0_outputs(6227);
    layer1_outputs(5610) <= not(layer0_outputs(11179));
    layer1_outputs(5611) <= '1';
    layer1_outputs(5612) <= (layer0_outputs(6977)) and not (layer0_outputs(1929));
    layer1_outputs(5613) <= not(layer0_outputs(9866)) or (layer0_outputs(1199));
    layer1_outputs(5614) <= (layer0_outputs(6083)) and (layer0_outputs(7071));
    layer1_outputs(5615) <= '1';
    layer1_outputs(5616) <= not(layer0_outputs(3666)) or (layer0_outputs(4707));
    layer1_outputs(5617) <= layer0_outputs(3415);
    layer1_outputs(5618) <= not((layer0_outputs(3)) xor (layer0_outputs(1104)));
    layer1_outputs(5619) <= layer0_outputs(7099);
    layer1_outputs(5620) <= layer0_outputs(11168);
    layer1_outputs(5621) <= (layer0_outputs(3575)) or (layer0_outputs(2912));
    layer1_outputs(5622) <= layer0_outputs(10630);
    layer1_outputs(5623) <= '0';
    layer1_outputs(5624) <= (layer0_outputs(1266)) and not (layer0_outputs(1916));
    layer1_outputs(5625) <= not((layer0_outputs(4346)) or (layer0_outputs(8958)));
    layer1_outputs(5626) <= not(layer0_outputs(10839)) or (layer0_outputs(9116));
    layer1_outputs(5627) <= not(layer0_outputs(7205));
    layer1_outputs(5628) <= not((layer0_outputs(5304)) xor (layer0_outputs(7874)));
    layer1_outputs(5629) <= layer0_outputs(9060);
    layer1_outputs(5630) <= not((layer0_outputs(4123)) or (layer0_outputs(12729)));
    layer1_outputs(5631) <= layer0_outputs(3579);
    layer1_outputs(5632) <= (layer0_outputs(9189)) xor (layer0_outputs(219));
    layer1_outputs(5633) <= not(layer0_outputs(5463));
    layer1_outputs(5634) <= layer0_outputs(9430);
    layer1_outputs(5635) <= not((layer0_outputs(9071)) or (layer0_outputs(11714)));
    layer1_outputs(5636) <= layer0_outputs(2024);
    layer1_outputs(5637) <= not(layer0_outputs(10175));
    layer1_outputs(5638) <= not(layer0_outputs(3849));
    layer1_outputs(5639) <= not(layer0_outputs(6773)) or (layer0_outputs(6191));
    layer1_outputs(5640) <= layer0_outputs(11718);
    layer1_outputs(5641) <= not((layer0_outputs(312)) xor (layer0_outputs(2978)));
    layer1_outputs(5642) <= not(layer0_outputs(7704)) or (layer0_outputs(4847));
    layer1_outputs(5643) <= not(layer0_outputs(2920)) or (layer0_outputs(617));
    layer1_outputs(5644) <= not(layer0_outputs(3551)) or (layer0_outputs(11465));
    layer1_outputs(5645) <= (layer0_outputs(1518)) and not (layer0_outputs(3107));
    layer1_outputs(5646) <= not(layer0_outputs(12115));
    layer1_outputs(5647) <= not(layer0_outputs(9095));
    layer1_outputs(5648) <= (layer0_outputs(7196)) and not (layer0_outputs(5647));
    layer1_outputs(5649) <= layer0_outputs(5473);
    layer1_outputs(5650) <= not(layer0_outputs(1370));
    layer1_outputs(5651) <= (layer0_outputs(3853)) or (layer0_outputs(4522));
    layer1_outputs(5652) <= (layer0_outputs(10031)) xor (layer0_outputs(2827));
    layer1_outputs(5653) <= not(layer0_outputs(1261));
    layer1_outputs(5654) <= not((layer0_outputs(11669)) xor (layer0_outputs(11894)));
    layer1_outputs(5655) <= not((layer0_outputs(1882)) and (layer0_outputs(2663)));
    layer1_outputs(5656) <= not(layer0_outputs(9387));
    layer1_outputs(5657) <= not((layer0_outputs(2859)) xor (layer0_outputs(8027)));
    layer1_outputs(5658) <= '0';
    layer1_outputs(5659) <= '1';
    layer1_outputs(5660) <= not(layer0_outputs(12716)) or (layer0_outputs(2164));
    layer1_outputs(5661) <= not((layer0_outputs(2080)) or (layer0_outputs(3725)));
    layer1_outputs(5662) <= not(layer0_outputs(6398));
    layer1_outputs(5663) <= not(layer0_outputs(3791)) or (layer0_outputs(2893));
    layer1_outputs(5664) <= (layer0_outputs(7680)) and not (layer0_outputs(9623));
    layer1_outputs(5665) <= layer0_outputs(11921);
    layer1_outputs(5666) <= (layer0_outputs(9733)) and (layer0_outputs(4173));
    layer1_outputs(5667) <= not(layer0_outputs(5324));
    layer1_outputs(5668) <= layer0_outputs(129);
    layer1_outputs(5669) <= layer0_outputs(4042);
    layer1_outputs(5670) <= not(layer0_outputs(8157)) or (layer0_outputs(6694));
    layer1_outputs(5671) <= layer0_outputs(4945);
    layer1_outputs(5672) <= layer0_outputs(4474);
    layer1_outputs(5673) <= layer0_outputs(2371);
    layer1_outputs(5674) <= (layer0_outputs(4391)) and not (layer0_outputs(6823));
    layer1_outputs(5675) <= (layer0_outputs(10813)) and (layer0_outputs(9134));
    layer1_outputs(5676) <= not((layer0_outputs(8062)) xor (layer0_outputs(6468)));
    layer1_outputs(5677) <= not((layer0_outputs(4780)) and (layer0_outputs(5148)));
    layer1_outputs(5678) <= layer0_outputs(1839);
    layer1_outputs(5679) <= (layer0_outputs(5685)) xor (layer0_outputs(9394));
    layer1_outputs(5680) <= not((layer0_outputs(4705)) xor (layer0_outputs(12655)));
    layer1_outputs(5681) <= (layer0_outputs(9823)) or (layer0_outputs(2819));
    layer1_outputs(5682) <= not(layer0_outputs(364));
    layer1_outputs(5683) <= not(layer0_outputs(7333));
    layer1_outputs(5684) <= not(layer0_outputs(9584));
    layer1_outputs(5685) <= not((layer0_outputs(4168)) or (layer0_outputs(4392)));
    layer1_outputs(5686) <= layer0_outputs(8491);
    layer1_outputs(5687) <= not(layer0_outputs(3343));
    layer1_outputs(5688) <= layer0_outputs(479);
    layer1_outputs(5689) <= layer0_outputs(11593);
    layer1_outputs(5690) <= layer0_outputs(3504);
    layer1_outputs(5691) <= (layer0_outputs(9656)) and not (layer0_outputs(3040));
    layer1_outputs(5692) <= layer0_outputs(10787);
    layer1_outputs(5693) <= '0';
    layer1_outputs(5694) <= not(layer0_outputs(6876)) or (layer0_outputs(7516));
    layer1_outputs(5695) <= (layer0_outputs(9174)) and not (layer0_outputs(6585));
    layer1_outputs(5696) <= layer0_outputs(9691);
    layer1_outputs(5697) <= not(layer0_outputs(3670));
    layer1_outputs(5698) <= not((layer0_outputs(6669)) xor (layer0_outputs(5279)));
    layer1_outputs(5699) <= not((layer0_outputs(1664)) or (layer0_outputs(5603)));
    layer1_outputs(5700) <= layer0_outputs(9445);
    layer1_outputs(5701) <= not(layer0_outputs(5982)) or (layer0_outputs(10460));
    layer1_outputs(5702) <= layer0_outputs(4121);
    layer1_outputs(5703) <= not((layer0_outputs(4559)) and (layer0_outputs(8517)));
    layer1_outputs(5704) <= not((layer0_outputs(2705)) xor (layer0_outputs(8086)));
    layer1_outputs(5705) <= not(layer0_outputs(1740));
    layer1_outputs(5706) <= layer0_outputs(1353);
    layer1_outputs(5707) <= layer0_outputs(4544);
    layer1_outputs(5708) <= not((layer0_outputs(10779)) xor (layer0_outputs(5522)));
    layer1_outputs(5709) <= layer0_outputs(3911);
    layer1_outputs(5710) <= (layer0_outputs(3097)) and not (layer0_outputs(11711));
    layer1_outputs(5711) <= not(layer0_outputs(2512));
    layer1_outputs(5712) <= not((layer0_outputs(7603)) and (layer0_outputs(11417)));
    layer1_outputs(5713) <= not((layer0_outputs(7229)) xor (layer0_outputs(8016)));
    layer1_outputs(5714) <= not(layer0_outputs(1345));
    layer1_outputs(5715) <= (layer0_outputs(4596)) and not (layer0_outputs(10306));
    layer1_outputs(5716) <= not((layer0_outputs(12796)) xor (layer0_outputs(7445)));
    layer1_outputs(5717) <= layer0_outputs(9554);
    layer1_outputs(5718) <= layer0_outputs(9329);
    layer1_outputs(5719) <= (layer0_outputs(4807)) or (layer0_outputs(5726));
    layer1_outputs(5720) <= not(layer0_outputs(3067));
    layer1_outputs(5721) <= not(layer0_outputs(8300));
    layer1_outputs(5722) <= not(layer0_outputs(2076));
    layer1_outputs(5723) <= not(layer0_outputs(3069));
    layer1_outputs(5724) <= not((layer0_outputs(2047)) xor (layer0_outputs(10759)));
    layer1_outputs(5725) <= not((layer0_outputs(7442)) xor (layer0_outputs(1591)));
    layer1_outputs(5726) <= '1';
    layer1_outputs(5727) <= layer0_outputs(5339);
    layer1_outputs(5728) <= not((layer0_outputs(6689)) xor (layer0_outputs(3061)));
    layer1_outputs(5729) <= (layer0_outputs(7387)) or (layer0_outputs(3776));
    layer1_outputs(5730) <= not(layer0_outputs(4135));
    layer1_outputs(5731) <= not(layer0_outputs(12072)) or (layer0_outputs(3543));
    layer1_outputs(5732) <= not((layer0_outputs(12668)) or (layer0_outputs(12553)));
    layer1_outputs(5733) <= layer0_outputs(11918);
    layer1_outputs(5734) <= not((layer0_outputs(6736)) and (layer0_outputs(6135)));
    layer1_outputs(5735) <= not(layer0_outputs(5550));
    layer1_outputs(5736) <= (layer0_outputs(9600)) and not (layer0_outputs(7513));
    layer1_outputs(5737) <= (layer0_outputs(10104)) and not (layer0_outputs(7763));
    layer1_outputs(5738) <= not(layer0_outputs(8911)) or (layer0_outputs(1540));
    layer1_outputs(5739) <= layer0_outputs(10696);
    layer1_outputs(5740) <= not(layer0_outputs(3590));
    layer1_outputs(5741) <= not(layer0_outputs(3348));
    layer1_outputs(5742) <= not(layer0_outputs(2443));
    layer1_outputs(5743) <= (layer0_outputs(7307)) or (layer0_outputs(11978));
    layer1_outputs(5744) <= (layer0_outputs(3424)) xor (layer0_outputs(9589));
    layer1_outputs(5745) <= not(layer0_outputs(7304));
    layer1_outputs(5746) <= (layer0_outputs(3655)) and not (layer0_outputs(12793));
    layer1_outputs(5747) <= layer0_outputs(11013);
    layer1_outputs(5748) <= '0';
    layer1_outputs(5749) <= not(layer0_outputs(2223));
    layer1_outputs(5750) <= (layer0_outputs(767)) xor (layer0_outputs(8691));
    layer1_outputs(5751) <= (layer0_outputs(2879)) xor (layer0_outputs(2017));
    layer1_outputs(5752) <= not(layer0_outputs(5322)) or (layer0_outputs(9525));
    layer1_outputs(5753) <= layer0_outputs(1644);
    layer1_outputs(5754) <= layer0_outputs(9183);
    layer1_outputs(5755) <= not((layer0_outputs(1637)) or (layer0_outputs(7846)));
    layer1_outputs(5756) <= not(layer0_outputs(4923)) or (layer0_outputs(8980));
    layer1_outputs(5757) <= not((layer0_outputs(1189)) xor (layer0_outputs(6223)));
    layer1_outputs(5758) <= (layer0_outputs(9254)) or (layer0_outputs(1888));
    layer1_outputs(5759) <= not((layer0_outputs(2875)) and (layer0_outputs(6640)));
    layer1_outputs(5760) <= not((layer0_outputs(5913)) and (layer0_outputs(3100)));
    layer1_outputs(5761) <= (layer0_outputs(460)) and (layer0_outputs(10492));
    layer1_outputs(5762) <= not((layer0_outputs(690)) or (layer0_outputs(7924)));
    layer1_outputs(5763) <= (layer0_outputs(10647)) and (layer0_outputs(10427));
    layer1_outputs(5764) <= (layer0_outputs(744)) or (layer0_outputs(468));
    layer1_outputs(5765) <= (layer0_outputs(6786)) xor (layer0_outputs(8792));
    layer1_outputs(5766) <= layer0_outputs(2865);
    layer1_outputs(5767) <= (layer0_outputs(10211)) xor (layer0_outputs(5339));
    layer1_outputs(5768) <= not((layer0_outputs(8393)) xor (layer0_outputs(5821)));
    layer1_outputs(5769) <= '0';
    layer1_outputs(5770) <= (layer0_outputs(12069)) or (layer0_outputs(12442));
    layer1_outputs(5771) <= layer0_outputs(5000);
    layer1_outputs(5772) <= layer0_outputs(5239);
    layer1_outputs(5773) <= not(layer0_outputs(8187));
    layer1_outputs(5774) <= '0';
    layer1_outputs(5775) <= not((layer0_outputs(10181)) xor (layer0_outputs(3260)));
    layer1_outputs(5776) <= layer0_outputs(4383);
    layer1_outputs(5777) <= not(layer0_outputs(2447)) or (layer0_outputs(9282));
    layer1_outputs(5778) <= (layer0_outputs(991)) or (layer0_outputs(1201));
    layer1_outputs(5779) <= not(layer0_outputs(8422));
    layer1_outputs(5780) <= not(layer0_outputs(6606)) or (layer0_outputs(12193));
    layer1_outputs(5781) <= '1';
    layer1_outputs(5782) <= (layer0_outputs(11221)) and not (layer0_outputs(7567));
    layer1_outputs(5783) <= not(layer0_outputs(3548));
    layer1_outputs(5784) <= '0';
    layer1_outputs(5785) <= (layer0_outputs(4803)) and not (layer0_outputs(8565));
    layer1_outputs(5786) <= layer0_outputs(6035);
    layer1_outputs(5787) <= not(layer0_outputs(650));
    layer1_outputs(5788) <= (layer0_outputs(12594)) or (layer0_outputs(5174));
    layer1_outputs(5789) <= (layer0_outputs(4467)) and (layer0_outputs(7337));
    layer1_outputs(5790) <= layer0_outputs(6365);
    layer1_outputs(5791) <= not((layer0_outputs(1554)) and (layer0_outputs(4501)));
    layer1_outputs(5792) <= not(layer0_outputs(1588));
    layer1_outputs(5793) <= (layer0_outputs(12610)) and (layer0_outputs(3681));
    layer1_outputs(5794) <= layer0_outputs(9127);
    layer1_outputs(5795) <= not(layer0_outputs(2544));
    layer1_outputs(5796) <= (layer0_outputs(11286)) and not (layer0_outputs(1855));
    layer1_outputs(5797) <= layer0_outputs(417);
    layer1_outputs(5798) <= not(layer0_outputs(8720));
    layer1_outputs(5799) <= (layer0_outputs(12608)) and not (layer0_outputs(245));
    layer1_outputs(5800) <= (layer0_outputs(12460)) xor (layer0_outputs(575));
    layer1_outputs(5801) <= not(layer0_outputs(2548)) or (layer0_outputs(8632));
    layer1_outputs(5802) <= not(layer0_outputs(242));
    layer1_outputs(5803) <= not(layer0_outputs(2781));
    layer1_outputs(5804) <= (layer0_outputs(12416)) and not (layer0_outputs(9794));
    layer1_outputs(5805) <= (layer0_outputs(9149)) and (layer0_outputs(597));
    layer1_outputs(5806) <= (layer0_outputs(8489)) and not (layer0_outputs(1085));
    layer1_outputs(5807) <= not(layer0_outputs(7805)) or (layer0_outputs(2937));
    layer1_outputs(5808) <= (layer0_outputs(11868)) xor (layer0_outputs(601));
    layer1_outputs(5809) <= not((layer0_outputs(7613)) xor (layer0_outputs(10694)));
    layer1_outputs(5810) <= not(layer0_outputs(2549)) or (layer0_outputs(2194));
    layer1_outputs(5811) <= not(layer0_outputs(9764)) or (layer0_outputs(1412));
    layer1_outputs(5812) <= not((layer0_outputs(12131)) or (layer0_outputs(9409)));
    layer1_outputs(5813) <= (layer0_outputs(8614)) and (layer0_outputs(11729));
    layer1_outputs(5814) <= not(layer0_outputs(2604));
    layer1_outputs(5815) <= (layer0_outputs(4570)) and not (layer0_outputs(9315));
    layer1_outputs(5816) <= not(layer0_outputs(4315)) or (layer0_outputs(8645));
    layer1_outputs(5817) <= not(layer0_outputs(5058));
    layer1_outputs(5818) <= not(layer0_outputs(3120)) or (layer0_outputs(8627));
    layer1_outputs(5819) <= not(layer0_outputs(8102));
    layer1_outputs(5820) <= layer0_outputs(2544);
    layer1_outputs(5821) <= not(layer0_outputs(12261));
    layer1_outputs(5822) <= (layer0_outputs(4809)) and (layer0_outputs(3336));
    layer1_outputs(5823) <= not(layer0_outputs(6735));
    layer1_outputs(5824) <= not(layer0_outputs(12433));
    layer1_outputs(5825) <= (layer0_outputs(11533)) xor (layer0_outputs(9239));
    layer1_outputs(5826) <= '0';
    layer1_outputs(5827) <= not((layer0_outputs(1502)) xor (layer0_outputs(5331)));
    layer1_outputs(5828) <= (layer0_outputs(95)) and (layer0_outputs(5190));
    layer1_outputs(5829) <= layer0_outputs(432);
    layer1_outputs(5830) <= '0';
    layer1_outputs(5831) <= not(layer0_outputs(10642)) or (layer0_outputs(12029));
    layer1_outputs(5832) <= not(layer0_outputs(7409)) or (layer0_outputs(4770));
    layer1_outputs(5833) <= layer0_outputs(9427);
    layer1_outputs(5834) <= layer0_outputs(1480);
    layer1_outputs(5835) <= (layer0_outputs(11777)) and not (layer0_outputs(1531));
    layer1_outputs(5836) <= not(layer0_outputs(2051));
    layer1_outputs(5837) <= (layer0_outputs(9400)) xor (layer0_outputs(2401));
    layer1_outputs(5838) <= not(layer0_outputs(1912));
    layer1_outputs(5839) <= not(layer0_outputs(9800)) or (layer0_outputs(4475));
    layer1_outputs(5840) <= not(layer0_outputs(12077));
    layer1_outputs(5841) <= layer0_outputs(5465);
    layer1_outputs(5842) <= not((layer0_outputs(8712)) or (layer0_outputs(7230)));
    layer1_outputs(5843) <= (layer0_outputs(10554)) and not (layer0_outputs(2232));
    layer1_outputs(5844) <= layer0_outputs(4518);
    layer1_outputs(5845) <= not((layer0_outputs(11933)) and (layer0_outputs(2826)));
    layer1_outputs(5846) <= (layer0_outputs(6434)) and not (layer0_outputs(5320));
    layer1_outputs(5847) <= not((layer0_outputs(11957)) xor (layer0_outputs(11542)));
    layer1_outputs(5848) <= not((layer0_outputs(11624)) or (layer0_outputs(8596)));
    layer1_outputs(5849) <= '1';
    layer1_outputs(5850) <= not(layer0_outputs(12317)) or (layer0_outputs(12424));
    layer1_outputs(5851) <= not(layer0_outputs(3382));
    layer1_outputs(5852) <= (layer0_outputs(4643)) and not (layer0_outputs(10978));
    layer1_outputs(5853) <= (layer0_outputs(3034)) and not (layer0_outputs(5615));
    layer1_outputs(5854) <= (layer0_outputs(3647)) and not (layer0_outputs(9474));
    layer1_outputs(5855) <= layer0_outputs(4532);
    layer1_outputs(5856) <= layer0_outputs(11894);
    layer1_outputs(5857) <= not((layer0_outputs(6242)) xor (layer0_outputs(6721)));
    layer1_outputs(5858) <= not((layer0_outputs(6339)) xor (layer0_outputs(5422)));
    layer1_outputs(5859) <= (layer0_outputs(192)) or (layer0_outputs(9033));
    layer1_outputs(5860) <= not(layer0_outputs(11212));
    layer1_outputs(5861) <= not(layer0_outputs(9188));
    layer1_outputs(5862) <= (layer0_outputs(5928)) and not (layer0_outputs(1746));
    layer1_outputs(5863) <= (layer0_outputs(8808)) and not (layer0_outputs(6267));
    layer1_outputs(5864) <= not(layer0_outputs(2310));
    layer1_outputs(5865) <= (layer0_outputs(8232)) and (layer0_outputs(7943));
    layer1_outputs(5866) <= (layer0_outputs(7058)) and (layer0_outputs(1113));
    layer1_outputs(5867) <= not(layer0_outputs(6494));
    layer1_outputs(5868) <= layer0_outputs(6283);
    layer1_outputs(5869) <= not(layer0_outputs(3307));
    layer1_outputs(5870) <= (layer0_outputs(595)) or (layer0_outputs(7624));
    layer1_outputs(5871) <= layer0_outputs(8514);
    layer1_outputs(5872) <= layer0_outputs(5509);
    layer1_outputs(5873) <= not(layer0_outputs(2657));
    layer1_outputs(5874) <= not(layer0_outputs(6409));
    layer1_outputs(5875) <= (layer0_outputs(12259)) and not (layer0_outputs(9883));
    layer1_outputs(5876) <= layer0_outputs(3754);
    layer1_outputs(5877) <= not((layer0_outputs(7343)) or (layer0_outputs(11835)));
    layer1_outputs(5878) <= not(layer0_outputs(12398));
    layer1_outputs(5879) <= (layer0_outputs(11032)) xor (layer0_outputs(8410));
    layer1_outputs(5880) <= not(layer0_outputs(10936));
    layer1_outputs(5881) <= layer0_outputs(7269);
    layer1_outputs(5882) <= not(layer0_outputs(1618));
    layer1_outputs(5883) <= (layer0_outputs(544)) or (layer0_outputs(9755));
    layer1_outputs(5884) <= not(layer0_outputs(6570));
    layer1_outputs(5885) <= not(layer0_outputs(10763));
    layer1_outputs(5886) <= layer0_outputs(8211);
    layer1_outputs(5887) <= not((layer0_outputs(3925)) or (layer0_outputs(2536)));
    layer1_outputs(5888) <= (layer0_outputs(8402)) and not (layer0_outputs(1988));
    layer1_outputs(5889) <= '0';
    layer1_outputs(5890) <= not((layer0_outputs(147)) and (layer0_outputs(11632)));
    layer1_outputs(5891) <= (layer0_outputs(12157)) and not (layer0_outputs(12068));
    layer1_outputs(5892) <= (layer0_outputs(9115)) xor (layer0_outputs(5362));
    layer1_outputs(5893) <= layer0_outputs(11086);
    layer1_outputs(5894) <= (layer0_outputs(12169)) or (layer0_outputs(1941));
    layer1_outputs(5895) <= not(layer0_outputs(3903)) or (layer0_outputs(5132));
    layer1_outputs(5896) <= layer0_outputs(10659);
    layer1_outputs(5897) <= (layer0_outputs(75)) and (layer0_outputs(8792));
    layer1_outputs(5898) <= layer0_outputs(3632);
    layer1_outputs(5899) <= not(layer0_outputs(7129)) or (layer0_outputs(8695));
    layer1_outputs(5900) <= not(layer0_outputs(9618));
    layer1_outputs(5901) <= not((layer0_outputs(5475)) xor (layer0_outputs(4479)));
    layer1_outputs(5902) <= not((layer0_outputs(4990)) or (layer0_outputs(11645)));
    layer1_outputs(5903) <= not(layer0_outputs(10098));
    layer1_outputs(5904) <= (layer0_outputs(67)) and not (layer0_outputs(2951));
    layer1_outputs(5905) <= not(layer0_outputs(12177));
    layer1_outputs(5906) <= not(layer0_outputs(130));
    layer1_outputs(5907) <= not(layer0_outputs(2698));
    layer1_outputs(5908) <= not(layer0_outputs(1635)) or (layer0_outputs(2119));
    layer1_outputs(5909) <= layer0_outputs(4346);
    layer1_outputs(5910) <= not(layer0_outputs(4095));
    layer1_outputs(5911) <= (layer0_outputs(5234)) and not (layer0_outputs(12369));
    layer1_outputs(5912) <= not(layer0_outputs(8924)) or (layer0_outputs(9334));
    layer1_outputs(5913) <= (layer0_outputs(957)) and (layer0_outputs(12014));
    layer1_outputs(5914) <= not(layer0_outputs(5334));
    layer1_outputs(5915) <= (layer0_outputs(5782)) or (layer0_outputs(5707));
    layer1_outputs(5916) <= not(layer0_outputs(1358));
    layer1_outputs(5917) <= (layer0_outputs(10363)) and not (layer0_outputs(7254));
    layer1_outputs(5918) <= not(layer0_outputs(1724));
    layer1_outputs(5919) <= (layer0_outputs(1573)) xor (layer0_outputs(4691));
    layer1_outputs(5920) <= (layer0_outputs(5473)) and (layer0_outputs(7972));
    layer1_outputs(5921) <= not(layer0_outputs(4937));
    layer1_outputs(5922) <= not(layer0_outputs(7341)) or (layer0_outputs(4729));
    layer1_outputs(5923) <= (layer0_outputs(10571)) or (layer0_outputs(9607));
    layer1_outputs(5924) <= layer0_outputs(565);
    layer1_outputs(5925) <= not((layer0_outputs(12065)) xor (layer0_outputs(9207)));
    layer1_outputs(5926) <= not(layer0_outputs(4287));
    layer1_outputs(5927) <= not(layer0_outputs(5539));
    layer1_outputs(5928) <= (layer0_outputs(10623)) and not (layer0_outputs(7988));
    layer1_outputs(5929) <= not(layer0_outputs(2467)) or (layer0_outputs(7815));
    layer1_outputs(5930) <= layer0_outputs(6965);
    layer1_outputs(5931) <= not((layer0_outputs(9869)) or (layer0_outputs(5934)));
    layer1_outputs(5932) <= layer0_outputs(19);
    layer1_outputs(5933) <= not((layer0_outputs(3767)) and (layer0_outputs(1567)));
    layer1_outputs(5934) <= not((layer0_outputs(10317)) and (layer0_outputs(10615)));
    layer1_outputs(5935) <= not((layer0_outputs(4590)) and (layer0_outputs(6829)));
    layer1_outputs(5936) <= not(layer0_outputs(12045));
    layer1_outputs(5937) <= not(layer0_outputs(9044));
    layer1_outputs(5938) <= not(layer0_outputs(8013)) or (layer0_outputs(8547));
    layer1_outputs(5939) <= (layer0_outputs(9289)) and not (layer0_outputs(5817));
    layer1_outputs(5940) <= not((layer0_outputs(2307)) xor (layer0_outputs(12617)));
    layer1_outputs(5941) <= layer0_outputs(5829);
    layer1_outputs(5942) <= (layer0_outputs(7096)) xor (layer0_outputs(10547));
    layer1_outputs(5943) <= not((layer0_outputs(8748)) xor (layer0_outputs(5051)));
    layer1_outputs(5944) <= not(layer0_outputs(4575));
    layer1_outputs(5945) <= not(layer0_outputs(8854)) or (layer0_outputs(4759));
    layer1_outputs(5946) <= layer0_outputs(5179);
    layer1_outputs(5947) <= layer0_outputs(5708);
    layer1_outputs(5948) <= (layer0_outputs(6643)) or (layer0_outputs(5981));
    layer1_outputs(5949) <= (layer0_outputs(5384)) and (layer0_outputs(297));
    layer1_outputs(5950) <= (layer0_outputs(8527)) and (layer0_outputs(10769));
    layer1_outputs(5951) <= not(layer0_outputs(4668));
    layer1_outputs(5952) <= layer0_outputs(3118);
    layer1_outputs(5953) <= not(layer0_outputs(4306));
    layer1_outputs(5954) <= layer0_outputs(11482);
    layer1_outputs(5955) <= not(layer0_outputs(4202));
    layer1_outputs(5956) <= not(layer0_outputs(6977));
    layer1_outputs(5957) <= (layer0_outputs(8318)) xor (layer0_outputs(380));
    layer1_outputs(5958) <= (layer0_outputs(8293)) and not (layer0_outputs(1095));
    layer1_outputs(5959) <= (layer0_outputs(7575)) and not (layer0_outputs(7214));
    layer1_outputs(5960) <= layer0_outputs(3848);
    layer1_outputs(5961) <= not(layer0_outputs(5278));
    layer1_outputs(5962) <= not((layer0_outputs(11540)) xor (layer0_outputs(12554)));
    layer1_outputs(5963) <= not(layer0_outputs(10858)) or (layer0_outputs(5264));
    layer1_outputs(5964) <= (layer0_outputs(11098)) xor (layer0_outputs(1174));
    layer1_outputs(5965) <= layer0_outputs(12356);
    layer1_outputs(5966) <= (layer0_outputs(2244)) xor (layer0_outputs(9627));
    layer1_outputs(5967) <= (layer0_outputs(7836)) and not (layer0_outputs(12425));
    layer1_outputs(5968) <= (layer0_outputs(352)) and not (layer0_outputs(8225));
    layer1_outputs(5969) <= not(layer0_outputs(2718)) or (layer0_outputs(6145));
    layer1_outputs(5970) <= not((layer0_outputs(2818)) and (layer0_outputs(7990)));
    layer1_outputs(5971) <= not(layer0_outputs(6585));
    layer1_outputs(5972) <= (layer0_outputs(805)) xor (layer0_outputs(9825));
    layer1_outputs(5973) <= (layer0_outputs(6234)) xor (layer0_outputs(7686));
    layer1_outputs(5974) <= layer0_outputs(6592);
    layer1_outputs(5975) <= layer0_outputs(10168);
    layer1_outputs(5976) <= (layer0_outputs(4407)) and (layer0_outputs(8980));
    layer1_outputs(5977) <= (layer0_outputs(8398)) and not (layer0_outputs(9979));
    layer1_outputs(5978) <= (layer0_outputs(9470)) and not (layer0_outputs(9365));
    layer1_outputs(5979) <= not(layer0_outputs(80)) or (layer0_outputs(9269));
    layer1_outputs(5980) <= not(layer0_outputs(8894)) or (layer0_outputs(5596));
    layer1_outputs(5981) <= layer0_outputs(8501);
    layer1_outputs(5982) <= (layer0_outputs(1152)) or (layer0_outputs(635));
    layer1_outputs(5983) <= layer0_outputs(8625);
    layer1_outputs(5984) <= layer0_outputs(5570);
    layer1_outputs(5985) <= not(layer0_outputs(10220)) or (layer0_outputs(1542));
    layer1_outputs(5986) <= (layer0_outputs(9834)) and (layer0_outputs(12331));
    layer1_outputs(5987) <= (layer0_outputs(1604)) and not (layer0_outputs(11138));
    layer1_outputs(5988) <= (layer0_outputs(11311)) and not (layer0_outputs(4772));
    layer1_outputs(5989) <= (layer0_outputs(10994)) xor (layer0_outputs(6967));
    layer1_outputs(5990) <= not((layer0_outputs(3006)) and (layer0_outputs(4445)));
    layer1_outputs(5991) <= (layer0_outputs(3327)) xor (layer0_outputs(5843));
    layer1_outputs(5992) <= (layer0_outputs(5104)) and not (layer0_outputs(435));
    layer1_outputs(5993) <= (layer0_outputs(5046)) and not (layer0_outputs(10489));
    layer1_outputs(5994) <= not(layer0_outputs(1606)) or (layer0_outputs(1522));
    layer1_outputs(5995) <= not(layer0_outputs(4019));
    layer1_outputs(5996) <= layer0_outputs(171);
    layer1_outputs(5997) <= not(layer0_outputs(5231)) or (layer0_outputs(8153));
    layer1_outputs(5998) <= (layer0_outputs(12207)) and not (layer0_outputs(10802));
    layer1_outputs(5999) <= not(layer0_outputs(144)) or (layer0_outputs(5375));
    layer1_outputs(6000) <= layer0_outputs(8528);
    layer1_outputs(6001) <= not((layer0_outputs(12358)) and (layer0_outputs(9507)));
    layer1_outputs(6002) <= layer0_outputs(8720);
    layer1_outputs(6003) <= (layer0_outputs(366)) xor (layer0_outputs(12396));
    layer1_outputs(6004) <= not((layer0_outputs(11473)) or (layer0_outputs(6304)));
    layer1_outputs(6005) <= layer0_outputs(6551);
    layer1_outputs(6006) <= (layer0_outputs(2839)) and not (layer0_outputs(5296));
    layer1_outputs(6007) <= (layer0_outputs(4070)) and (layer0_outputs(12486));
    layer1_outputs(6008) <= layer0_outputs(3342);
    layer1_outputs(6009) <= not((layer0_outputs(4402)) and (layer0_outputs(9146)));
    layer1_outputs(6010) <= (layer0_outputs(1373)) and not (layer0_outputs(4436));
    layer1_outputs(6011) <= layer0_outputs(7304);
    layer1_outputs(6012) <= not(layer0_outputs(7302));
    layer1_outputs(6013) <= layer0_outputs(4448);
    layer1_outputs(6014) <= (layer0_outputs(10199)) xor (layer0_outputs(8559));
    layer1_outputs(6015) <= not((layer0_outputs(7357)) xor (layer0_outputs(4443)));
    layer1_outputs(6016) <= (layer0_outputs(9536)) and not (layer0_outputs(5542));
    layer1_outputs(6017) <= (layer0_outputs(2732)) or (layer0_outputs(8152));
    layer1_outputs(6018) <= (layer0_outputs(2337)) and not (layer0_outputs(1909));
    layer1_outputs(6019) <= (layer0_outputs(10065)) xor (layer0_outputs(4062));
    layer1_outputs(6020) <= not((layer0_outputs(74)) xor (layer0_outputs(12115)));
    layer1_outputs(6021) <= not(layer0_outputs(1719));
    layer1_outputs(6022) <= not((layer0_outputs(11080)) or (layer0_outputs(5518)));
    layer1_outputs(6023) <= (layer0_outputs(11213)) and (layer0_outputs(1195));
    layer1_outputs(6024) <= not((layer0_outputs(4749)) and (layer0_outputs(7028)));
    layer1_outputs(6025) <= not(layer0_outputs(7300));
    layer1_outputs(6026) <= (layer0_outputs(4617)) and (layer0_outputs(11847));
    layer1_outputs(6027) <= not(layer0_outputs(12675));
    layer1_outputs(6028) <= layer0_outputs(3584);
    layer1_outputs(6029) <= not((layer0_outputs(11658)) xor (layer0_outputs(1959)));
    layer1_outputs(6030) <= not((layer0_outputs(1748)) and (layer0_outputs(4317)));
    layer1_outputs(6031) <= not(layer0_outputs(5861)) or (layer0_outputs(9460));
    layer1_outputs(6032) <= (layer0_outputs(10778)) xor (layer0_outputs(8863));
    layer1_outputs(6033) <= (layer0_outputs(2851)) or (layer0_outputs(7410));
    layer1_outputs(6034) <= (layer0_outputs(10890)) and not (layer0_outputs(10061));
    layer1_outputs(6035) <= layer0_outputs(9725);
    layer1_outputs(6036) <= not(layer0_outputs(4414)) or (layer0_outputs(5002));
    layer1_outputs(6037) <= not(layer0_outputs(11432));
    layer1_outputs(6038) <= layer0_outputs(9550);
    layer1_outputs(6039) <= (layer0_outputs(10816)) and (layer0_outputs(10194));
    layer1_outputs(6040) <= not(layer0_outputs(7334));
    layer1_outputs(6041) <= (layer0_outputs(6421)) and not (layer0_outputs(3843));
    layer1_outputs(6042) <= '1';
    layer1_outputs(6043) <= not((layer0_outputs(4898)) or (layer0_outputs(1346)));
    layer1_outputs(6044) <= not((layer0_outputs(4494)) and (layer0_outputs(9594)));
    layer1_outputs(6045) <= not(layer0_outputs(3764)) or (layer0_outputs(8721));
    layer1_outputs(6046) <= not((layer0_outputs(3686)) or (layer0_outputs(9486)));
    layer1_outputs(6047) <= not((layer0_outputs(3521)) or (layer0_outputs(12151)));
    layer1_outputs(6048) <= not(layer0_outputs(4921));
    layer1_outputs(6049) <= layer0_outputs(3164);
    layer1_outputs(6050) <= (layer0_outputs(6460)) or (layer0_outputs(7207));
    layer1_outputs(6051) <= not(layer0_outputs(96));
    layer1_outputs(6052) <= (layer0_outputs(1589)) and not (layer0_outputs(1070));
    layer1_outputs(6053) <= (layer0_outputs(3712)) xor (layer0_outputs(807));
    layer1_outputs(6054) <= not(layer0_outputs(8159));
    layer1_outputs(6055) <= layer0_outputs(9984);
    layer1_outputs(6056) <= '0';
    layer1_outputs(6057) <= layer0_outputs(9995);
    layer1_outputs(6058) <= (layer0_outputs(11296)) and not (layer0_outputs(12634));
    layer1_outputs(6059) <= (layer0_outputs(2071)) xor (layer0_outputs(562));
    layer1_outputs(6060) <= not(layer0_outputs(11809)) or (layer0_outputs(11791));
    layer1_outputs(6061) <= not(layer0_outputs(3340));
    layer1_outputs(6062) <= not(layer0_outputs(9260)) or (layer0_outputs(6418));
    layer1_outputs(6063) <= not(layer0_outputs(871));
    layer1_outputs(6064) <= not(layer0_outputs(3941));
    layer1_outputs(6065) <= layer0_outputs(8924);
    layer1_outputs(6066) <= (layer0_outputs(10531)) and not (layer0_outputs(2997));
    layer1_outputs(6067) <= '0';
    layer1_outputs(6068) <= (layer0_outputs(10408)) and not (layer0_outputs(5751));
    layer1_outputs(6069) <= (layer0_outputs(7143)) or (layer0_outputs(5));
    layer1_outputs(6070) <= layer0_outputs(12353);
    layer1_outputs(6071) <= layer0_outputs(7675);
    layer1_outputs(6072) <= layer0_outputs(7821);
    layer1_outputs(6073) <= (layer0_outputs(10842)) or (layer0_outputs(11484));
    layer1_outputs(6074) <= not(layer0_outputs(5146));
    layer1_outputs(6075) <= not(layer0_outputs(8871)) or (layer0_outputs(10636));
    layer1_outputs(6076) <= layer0_outputs(12629);
    layer1_outputs(6077) <= (layer0_outputs(7813)) xor (layer0_outputs(3598));
    layer1_outputs(6078) <= layer0_outputs(2081);
    layer1_outputs(6079) <= (layer0_outputs(7424)) and not (layer0_outputs(4436));
    layer1_outputs(6080) <= not(layer0_outputs(7612));
    layer1_outputs(6081) <= (layer0_outputs(12223)) or (layer0_outputs(12361));
    layer1_outputs(6082) <= (layer0_outputs(10215)) xor (layer0_outputs(3430));
    layer1_outputs(6083) <= (layer0_outputs(5630)) or (layer0_outputs(3740));
    layer1_outputs(6084) <= (layer0_outputs(1039)) xor (layer0_outputs(6441));
    layer1_outputs(6085) <= not(layer0_outputs(8556)) or (layer0_outputs(12723));
    layer1_outputs(6086) <= (layer0_outputs(7128)) or (layer0_outputs(3657));
    layer1_outputs(6087) <= (layer0_outputs(10878)) and not (layer0_outputs(5046));
    layer1_outputs(6088) <= not(layer0_outputs(8620));
    layer1_outputs(6089) <= (layer0_outputs(12049)) xor (layer0_outputs(5364));
    layer1_outputs(6090) <= not((layer0_outputs(3866)) and (layer0_outputs(2276)));
    layer1_outputs(6091) <= layer0_outputs(9337);
    layer1_outputs(6092) <= (layer0_outputs(516)) or (layer0_outputs(5392));
    layer1_outputs(6093) <= not(layer0_outputs(5492));
    layer1_outputs(6094) <= layer0_outputs(4797);
    layer1_outputs(6095) <= not(layer0_outputs(10575)) or (layer0_outputs(8193));
    layer1_outputs(6096) <= '1';
    layer1_outputs(6097) <= not(layer0_outputs(2136)) or (layer0_outputs(4317));
    layer1_outputs(6098) <= layer0_outputs(12133);
    layer1_outputs(6099) <= not(layer0_outputs(6727));
    layer1_outputs(6100) <= (layer0_outputs(6091)) and (layer0_outputs(6386));
    layer1_outputs(6101) <= not(layer0_outputs(2124));
    layer1_outputs(6102) <= (layer0_outputs(11746)) xor (layer0_outputs(6182));
    layer1_outputs(6103) <= layer0_outputs(2639);
    layer1_outputs(6104) <= (layer0_outputs(6671)) and (layer0_outputs(2769));
    layer1_outputs(6105) <= (layer0_outputs(2814)) or (layer0_outputs(4488));
    layer1_outputs(6106) <= (layer0_outputs(10861)) or (layer0_outputs(4877));
    layer1_outputs(6107) <= '1';
    layer1_outputs(6108) <= not(layer0_outputs(6236));
    layer1_outputs(6109) <= not(layer0_outputs(9477));
    layer1_outputs(6110) <= not(layer0_outputs(6452));
    layer1_outputs(6111) <= (layer0_outputs(11734)) and (layer0_outputs(2682));
    layer1_outputs(6112) <= not((layer0_outputs(3556)) xor (layer0_outputs(3451)));
    layer1_outputs(6113) <= not(layer0_outputs(9770));
    layer1_outputs(6114) <= (layer0_outputs(3910)) or (layer0_outputs(4897));
    layer1_outputs(6115) <= (layer0_outputs(9505)) and not (layer0_outputs(2479));
    layer1_outputs(6116) <= not(layer0_outputs(9990));
    layer1_outputs(6117) <= layer0_outputs(12105);
    layer1_outputs(6118) <= layer0_outputs(8357);
    layer1_outputs(6119) <= layer0_outputs(12049);
    layer1_outputs(6120) <= (layer0_outputs(736)) and (layer0_outputs(1223));
    layer1_outputs(6121) <= layer0_outputs(7163);
    layer1_outputs(6122) <= not((layer0_outputs(4379)) or (layer0_outputs(11192)));
    layer1_outputs(6123) <= not(layer0_outputs(2329)) or (layer0_outputs(12523));
    layer1_outputs(6124) <= (layer0_outputs(12515)) and not (layer0_outputs(2187));
    layer1_outputs(6125) <= (layer0_outputs(11852)) and (layer0_outputs(32));
    layer1_outputs(6126) <= (layer0_outputs(1943)) or (layer0_outputs(3572));
    layer1_outputs(6127) <= layer0_outputs(11778);
    layer1_outputs(6128) <= (layer0_outputs(9319)) or (layer0_outputs(4905));
    layer1_outputs(6129) <= (layer0_outputs(11557)) and not (layer0_outputs(9584));
    layer1_outputs(6130) <= not((layer0_outputs(7031)) and (layer0_outputs(12198)));
    layer1_outputs(6131) <= not((layer0_outputs(11020)) and (layer0_outputs(12557)));
    layer1_outputs(6132) <= (layer0_outputs(142)) or (layer0_outputs(2646));
    layer1_outputs(6133) <= '1';
    layer1_outputs(6134) <= not(layer0_outputs(2846));
    layer1_outputs(6135) <= not(layer0_outputs(4899));
    layer1_outputs(6136) <= layer0_outputs(554);
    layer1_outputs(6137) <= layer0_outputs(4857);
    layer1_outputs(6138) <= not(layer0_outputs(10273)) or (layer0_outputs(5905));
    layer1_outputs(6139) <= (layer0_outputs(10190)) or (layer0_outputs(1511));
    layer1_outputs(6140) <= (layer0_outputs(5594)) or (layer0_outputs(8160));
    layer1_outputs(6141) <= layer0_outputs(5159);
    layer1_outputs(6142) <= not((layer0_outputs(4010)) or (layer0_outputs(6536)));
    layer1_outputs(6143) <= (layer0_outputs(12620)) and (layer0_outputs(6472));
    layer1_outputs(6144) <= not((layer0_outputs(7855)) and (layer0_outputs(6834)));
    layer1_outputs(6145) <= layer0_outputs(7857);
    layer1_outputs(6146) <= not((layer0_outputs(12342)) xor (layer0_outputs(1978)));
    layer1_outputs(6147) <= layer0_outputs(10340);
    layer1_outputs(6148) <= not(layer0_outputs(6130));
    layer1_outputs(6149) <= not(layer0_outputs(2586));
    layer1_outputs(6150) <= (layer0_outputs(1090)) and not (layer0_outputs(9152));
    layer1_outputs(6151) <= '0';
    layer1_outputs(6152) <= (layer0_outputs(10373)) and not (layer0_outputs(10453));
    layer1_outputs(6153) <= (layer0_outputs(10870)) and (layer0_outputs(4058));
    layer1_outputs(6154) <= (layer0_outputs(7893)) and not (layer0_outputs(9613));
    layer1_outputs(6155) <= not((layer0_outputs(11248)) xor (layer0_outputs(6297)));
    layer1_outputs(6156) <= not(layer0_outputs(5512));
    layer1_outputs(6157) <= '0';
    layer1_outputs(6158) <= not((layer0_outputs(9459)) or (layer0_outputs(10787)));
    layer1_outputs(6159) <= not(layer0_outputs(3391)) or (layer0_outputs(2343));
    layer1_outputs(6160) <= layer0_outputs(986);
    layer1_outputs(6161) <= '0';
    layer1_outputs(6162) <= not(layer0_outputs(6412)) or (layer0_outputs(12699));
    layer1_outputs(6163) <= not((layer0_outputs(4309)) xor (layer0_outputs(9512)));
    layer1_outputs(6164) <= (layer0_outputs(9978)) xor (layer0_outputs(6276));
    layer1_outputs(6165) <= not((layer0_outputs(1002)) and (layer0_outputs(8506)));
    layer1_outputs(6166) <= not(layer0_outputs(4660)) or (layer0_outputs(5824));
    layer1_outputs(6167) <= (layer0_outputs(11471)) or (layer0_outputs(6815));
    layer1_outputs(6168) <= (layer0_outputs(2226)) and not (layer0_outputs(2518));
    layer1_outputs(6169) <= layer0_outputs(1878);
    layer1_outputs(6170) <= not(layer0_outputs(2246)) or (layer0_outputs(6622));
    layer1_outputs(6171) <= not(layer0_outputs(5026));
    layer1_outputs(6172) <= not((layer0_outputs(9130)) xor (layer0_outputs(11486)));
    layer1_outputs(6173) <= layer0_outputs(7248);
    layer1_outputs(6174) <= not((layer0_outputs(128)) or (layer0_outputs(1207)));
    layer1_outputs(6175) <= not(layer0_outputs(12423));
    layer1_outputs(6176) <= (layer0_outputs(2791)) and not (layer0_outputs(11729));
    layer1_outputs(6177) <= not(layer0_outputs(6459)) or (layer0_outputs(8462));
    layer1_outputs(6178) <= layer0_outputs(8926);
    layer1_outputs(6179) <= layer0_outputs(2855);
    layer1_outputs(6180) <= (layer0_outputs(4047)) and not (layer0_outputs(5218));
    layer1_outputs(6181) <= not(layer0_outputs(3151));
    layer1_outputs(6182) <= (layer0_outputs(1697)) or (layer0_outputs(1617));
    layer1_outputs(6183) <= not((layer0_outputs(7108)) and (layer0_outputs(4514)));
    layer1_outputs(6184) <= layer0_outputs(8110);
    layer1_outputs(6185) <= not((layer0_outputs(2712)) xor (layer0_outputs(1957)));
    layer1_outputs(6186) <= layer0_outputs(11637);
    layer1_outputs(6187) <= (layer0_outputs(1902)) and not (layer0_outputs(2437));
    layer1_outputs(6188) <= not((layer0_outputs(8372)) xor (layer0_outputs(4728)));
    layer1_outputs(6189) <= not(layer0_outputs(8781));
    layer1_outputs(6190) <= (layer0_outputs(4017)) and not (layer0_outputs(12373));
    layer1_outputs(6191) <= layer0_outputs(6572);
    layer1_outputs(6192) <= layer0_outputs(12704);
    layer1_outputs(6193) <= layer0_outputs(10805);
    layer1_outputs(6194) <= not((layer0_outputs(11528)) or (layer0_outputs(1749)));
    layer1_outputs(6195) <= layer0_outputs(1319);
    layer1_outputs(6196) <= (layer0_outputs(7810)) or (layer0_outputs(394));
    layer1_outputs(6197) <= not(layer0_outputs(12246));
    layer1_outputs(6198) <= not(layer0_outputs(7330));
    layer1_outputs(6199) <= (layer0_outputs(9853)) xor (layer0_outputs(2036));
    layer1_outputs(6200) <= (layer0_outputs(1738)) and not (layer0_outputs(497));
    layer1_outputs(6201) <= layer0_outputs(2091);
    layer1_outputs(6202) <= layer0_outputs(9494);
    layer1_outputs(6203) <= not((layer0_outputs(12676)) or (layer0_outputs(656)));
    layer1_outputs(6204) <= not(layer0_outputs(4492));
    layer1_outputs(6205) <= not((layer0_outputs(6210)) and (layer0_outputs(7826)));
    layer1_outputs(6206) <= layer0_outputs(2418);
    layer1_outputs(6207) <= not((layer0_outputs(9238)) and (layer0_outputs(2664)));
    layer1_outputs(6208) <= not(layer0_outputs(7953));
    layer1_outputs(6209) <= not(layer0_outputs(4269));
    layer1_outputs(6210) <= layer0_outputs(12297);
    layer1_outputs(6211) <= (layer0_outputs(6221)) and not (layer0_outputs(4245));
    layer1_outputs(6212) <= not(layer0_outputs(4399));
    layer1_outputs(6213) <= (layer0_outputs(7492)) and not (layer0_outputs(1822));
    layer1_outputs(6214) <= not(layer0_outputs(7579));
    layer1_outputs(6215) <= (layer0_outputs(569)) xor (layer0_outputs(2006));
    layer1_outputs(6216) <= not((layer0_outputs(11253)) or (layer0_outputs(4845)));
    layer1_outputs(6217) <= not((layer0_outputs(4438)) xor (layer0_outputs(6023)));
    layer1_outputs(6218) <= not((layer0_outputs(12792)) or (layer0_outputs(9015)));
    layer1_outputs(6219) <= layer0_outputs(4495);
    layer1_outputs(6220) <= (layer0_outputs(5101)) xor (layer0_outputs(9326));
    layer1_outputs(6221) <= (layer0_outputs(12543)) and not (layer0_outputs(7538));
    layer1_outputs(6222) <= (layer0_outputs(466)) xor (layer0_outputs(110));
    layer1_outputs(6223) <= layer0_outputs(8038);
    layer1_outputs(6224) <= not((layer0_outputs(8104)) xor (layer0_outputs(9091)));
    layer1_outputs(6225) <= not(layer0_outputs(11182));
    layer1_outputs(6226) <= (layer0_outputs(5589)) and not (layer0_outputs(6143));
    layer1_outputs(6227) <= (layer0_outputs(2417)) and (layer0_outputs(6679));
    layer1_outputs(6228) <= (layer0_outputs(3370)) and not (layer0_outputs(9692));
    layer1_outputs(6229) <= '0';
    layer1_outputs(6230) <= not(layer0_outputs(11351)) or (layer0_outputs(10200));
    layer1_outputs(6231) <= not(layer0_outputs(97));
    layer1_outputs(6232) <= layer0_outputs(9912);
    layer1_outputs(6233) <= layer0_outputs(7683);
    layer1_outputs(6234) <= '0';
    layer1_outputs(6235) <= (layer0_outputs(10952)) and not (layer0_outputs(5102));
    layer1_outputs(6236) <= layer0_outputs(10751);
    layer1_outputs(6237) <= layer0_outputs(1200);
    layer1_outputs(6238) <= layer0_outputs(12604);
    layer1_outputs(6239) <= (layer0_outputs(10979)) and (layer0_outputs(8921));
    layer1_outputs(6240) <= not((layer0_outputs(6843)) xor (layer0_outputs(8297)));
    layer1_outputs(6241) <= (layer0_outputs(6433)) and not (layer0_outputs(5392));
    layer1_outputs(6242) <= not((layer0_outputs(12263)) or (layer0_outputs(1815)));
    layer1_outputs(6243) <= (layer0_outputs(3795)) and not (layer0_outputs(8128));
    layer1_outputs(6244) <= (layer0_outputs(2394)) xor (layer0_outputs(9133));
    layer1_outputs(6245) <= not(layer0_outputs(193));
    layer1_outputs(6246) <= (layer0_outputs(1813)) xor (layer0_outputs(10982));
    layer1_outputs(6247) <= layer0_outputs(1243);
    layer1_outputs(6248) <= not(layer0_outputs(3675));
    layer1_outputs(6249) <= not((layer0_outputs(2556)) and (layer0_outputs(5198)));
    layer1_outputs(6250) <= not((layer0_outputs(287)) or (layer0_outputs(11299)));
    layer1_outputs(6251) <= (layer0_outputs(2912)) and (layer0_outputs(1012));
    layer1_outputs(6252) <= '1';
    layer1_outputs(6253) <= not(layer0_outputs(2731));
    layer1_outputs(6254) <= layer0_outputs(4287);
    layer1_outputs(6255) <= not((layer0_outputs(7268)) xor (layer0_outputs(12591)));
    layer1_outputs(6256) <= not(layer0_outputs(10505));
    layer1_outputs(6257) <= (layer0_outputs(11630)) and not (layer0_outputs(9769));
    layer1_outputs(6258) <= layer0_outputs(10107);
    layer1_outputs(6259) <= not(layer0_outputs(12112));
    layer1_outputs(6260) <= layer0_outputs(10768);
    layer1_outputs(6261) <= (layer0_outputs(2237)) and (layer0_outputs(6103));
    layer1_outputs(6262) <= not((layer0_outputs(5951)) and (layer0_outputs(973)));
    layer1_outputs(6263) <= layer0_outputs(9936);
    layer1_outputs(6264) <= not((layer0_outputs(4571)) and (layer0_outputs(380)));
    layer1_outputs(6265) <= layer0_outputs(12734);
    layer1_outputs(6266) <= layer0_outputs(6953);
    layer1_outputs(6267) <= not((layer0_outputs(9513)) and (layer0_outputs(5601)));
    layer1_outputs(6268) <= layer0_outputs(8576);
    layer1_outputs(6269) <= '1';
    layer1_outputs(6270) <= (layer0_outputs(8704)) and not (layer0_outputs(4007));
    layer1_outputs(6271) <= layer0_outputs(9693);
    layer1_outputs(6272) <= not(layer0_outputs(5664));
    layer1_outputs(6273) <= not((layer0_outputs(8228)) and (layer0_outputs(7543)));
    layer1_outputs(6274) <= (layer0_outputs(4288)) xor (layer0_outputs(9523));
    layer1_outputs(6275) <= layer0_outputs(12296);
    layer1_outputs(6276) <= layer0_outputs(1449);
    layer1_outputs(6277) <= '1';
    layer1_outputs(6278) <= layer0_outputs(7819);
    layer1_outputs(6279) <= not(layer0_outputs(7544)) or (layer0_outputs(7691));
    layer1_outputs(6280) <= (layer0_outputs(10795)) and not (layer0_outputs(7596));
    layer1_outputs(6281) <= (layer0_outputs(9711)) and not (layer0_outputs(10871));
    layer1_outputs(6282) <= (layer0_outputs(120)) and not (layer0_outputs(7606));
    layer1_outputs(6283) <= not(layer0_outputs(2991));
    layer1_outputs(6284) <= (layer0_outputs(3243)) xor (layer0_outputs(4164));
    layer1_outputs(6285) <= (layer0_outputs(7716)) or (layer0_outputs(6199));
    layer1_outputs(6286) <= layer0_outputs(12028);
    layer1_outputs(6287) <= not(layer0_outputs(4960));
    layer1_outputs(6288) <= layer0_outputs(9962);
    layer1_outputs(6289) <= not(layer0_outputs(10595)) or (layer0_outputs(9809));
    layer1_outputs(6290) <= (layer0_outputs(4987)) and (layer0_outputs(6862));
    layer1_outputs(6291) <= (layer0_outputs(9435)) xor (layer0_outputs(4051));
    layer1_outputs(6292) <= not(layer0_outputs(12774));
    layer1_outputs(6293) <= not(layer0_outputs(11162));
    layer1_outputs(6294) <= layer0_outputs(7427);
    layer1_outputs(6295) <= not((layer0_outputs(7918)) or (layer0_outputs(7616)));
    layer1_outputs(6296) <= (layer0_outputs(10684)) and not (layer0_outputs(6618));
    layer1_outputs(6297) <= not((layer0_outputs(8497)) or (layer0_outputs(6801)));
    layer1_outputs(6298) <= (layer0_outputs(11420)) and not (layer0_outputs(9259));
    layer1_outputs(6299) <= not(layer0_outputs(753));
    layer1_outputs(6300) <= layer0_outputs(3467);
    layer1_outputs(6301) <= layer0_outputs(7803);
    layer1_outputs(6302) <= not(layer0_outputs(12202)) or (layer0_outputs(10129));
    layer1_outputs(6303) <= not(layer0_outputs(8243)) or (layer0_outputs(6241));
    layer1_outputs(6304) <= (layer0_outputs(5944)) and (layer0_outputs(8570));
    layer1_outputs(6305) <= not(layer0_outputs(7714));
    layer1_outputs(6306) <= (layer0_outputs(9913)) or (layer0_outputs(4711));
    layer1_outputs(6307) <= (layer0_outputs(5753)) or (layer0_outputs(9443));
    layer1_outputs(6308) <= not(layer0_outputs(6896));
    layer1_outputs(6309) <= (layer0_outputs(11908)) and (layer0_outputs(8847));
    layer1_outputs(6310) <= layer0_outputs(3942);
    layer1_outputs(6311) <= (layer0_outputs(651)) or (layer0_outputs(9710));
    layer1_outputs(6312) <= (layer0_outputs(6062)) or (layer0_outputs(5969));
    layer1_outputs(6313) <= not((layer0_outputs(12471)) and (layer0_outputs(4611)));
    layer1_outputs(6314) <= layer0_outputs(7510);
    layer1_outputs(6315) <= not(layer0_outputs(9122));
    layer1_outputs(6316) <= layer0_outputs(2853);
    layer1_outputs(6317) <= not(layer0_outputs(4919)) or (layer0_outputs(3582));
    layer1_outputs(6318) <= (layer0_outputs(2315)) or (layer0_outputs(10689));
    layer1_outputs(6319) <= not(layer0_outputs(7522));
    layer1_outputs(6320) <= not(layer0_outputs(1642)) or (layer0_outputs(99));
    layer1_outputs(6321) <= not(layer0_outputs(1149)) or (layer0_outputs(11547));
    layer1_outputs(6322) <= not(layer0_outputs(7948));
    layer1_outputs(6323) <= not((layer0_outputs(2292)) and (layer0_outputs(1491)));
    layer1_outputs(6324) <= not(layer0_outputs(9213)) or (layer0_outputs(8832));
    layer1_outputs(6325) <= not(layer0_outputs(10232));
    layer1_outputs(6326) <= not(layer0_outputs(20));
    layer1_outputs(6327) <= not((layer0_outputs(7825)) and (layer0_outputs(6657)));
    layer1_outputs(6328) <= layer0_outputs(6320);
    layer1_outputs(6329) <= not(layer0_outputs(136)) or (layer0_outputs(5777));
    layer1_outputs(6330) <= not(layer0_outputs(8149)) or (layer0_outputs(8713));
    layer1_outputs(6331) <= not(layer0_outputs(3772));
    layer1_outputs(6332) <= (layer0_outputs(8680)) or (layer0_outputs(3707));
    layer1_outputs(6333) <= not((layer0_outputs(9782)) or (layer0_outputs(4422)));
    layer1_outputs(6334) <= not((layer0_outputs(12539)) and (layer0_outputs(3536)));
    layer1_outputs(6335) <= (layer0_outputs(11326)) or (layer0_outputs(11446));
    layer1_outputs(6336) <= (layer0_outputs(1381)) and not (layer0_outputs(10534));
    layer1_outputs(6337) <= (layer0_outputs(10665)) and (layer0_outputs(11452));
    layer1_outputs(6338) <= layer0_outputs(12186);
    layer1_outputs(6339) <= (layer0_outputs(6602)) and not (layer0_outputs(12299));
    layer1_outputs(6340) <= (layer0_outputs(12199)) xor (layer0_outputs(418));
    layer1_outputs(6341) <= layer0_outputs(7694);
    layer1_outputs(6342) <= not(layer0_outputs(10556)) or (layer0_outputs(6149));
    layer1_outputs(6343) <= not((layer0_outputs(5194)) xor (layer0_outputs(4451)));
    layer1_outputs(6344) <= (layer0_outputs(10554)) or (layer0_outputs(1675));
    layer1_outputs(6345) <= not(layer0_outputs(6046)) or (layer0_outputs(2387));
    layer1_outputs(6346) <= (layer0_outputs(4972)) and not (layer0_outputs(38));
    layer1_outputs(6347) <= not(layer0_outputs(2003)) or (layer0_outputs(1991));
    layer1_outputs(6348) <= (layer0_outputs(5920)) and not (layer0_outputs(1172));
    layer1_outputs(6349) <= not(layer0_outputs(449)) or (layer0_outputs(825));
    layer1_outputs(6350) <= not((layer0_outputs(228)) or (layer0_outputs(12543)));
    layer1_outputs(6351) <= not(layer0_outputs(858)) or (layer0_outputs(12407));
    layer1_outputs(6352) <= not(layer0_outputs(11771)) or (layer0_outputs(8065));
    layer1_outputs(6353) <= not((layer0_outputs(10600)) xor (layer0_outputs(5425)));
    layer1_outputs(6354) <= layer0_outputs(1720);
    layer1_outputs(6355) <= not(layer0_outputs(11462)) or (layer0_outputs(5812));
    layer1_outputs(6356) <= not(layer0_outputs(2654)) or (layer0_outputs(8082));
    layer1_outputs(6357) <= not(layer0_outputs(3010));
    layer1_outputs(6358) <= not(layer0_outputs(3700));
    layer1_outputs(6359) <= layer0_outputs(11698);
    layer1_outputs(6360) <= layer0_outputs(570);
    layer1_outputs(6361) <= not(layer0_outputs(6129));
    layer1_outputs(6362) <= not(layer0_outputs(4450));
    layer1_outputs(6363) <= (layer0_outputs(5248)) and not (layer0_outputs(9786));
    layer1_outputs(6364) <= not((layer0_outputs(4321)) and (layer0_outputs(3242)));
    layer1_outputs(6365) <= not((layer0_outputs(4974)) or (layer0_outputs(7897)));
    layer1_outputs(6366) <= (layer0_outputs(12121)) and (layer0_outputs(1824));
    layer1_outputs(6367) <= not(layer0_outputs(5235));
    layer1_outputs(6368) <= layer0_outputs(3331);
    layer1_outputs(6369) <= not(layer0_outputs(7863)) or (layer0_outputs(5768));
    layer1_outputs(6370) <= not((layer0_outputs(11622)) and (layer0_outputs(6506)));
    layer1_outputs(6371) <= not(layer0_outputs(4637));
    layer1_outputs(6372) <= (layer0_outputs(11612)) and not (layer0_outputs(7563));
    layer1_outputs(6373) <= not(layer0_outputs(9932));
    layer1_outputs(6374) <= (layer0_outputs(1203)) xor (layer0_outputs(1105));
    layer1_outputs(6375) <= (layer0_outputs(8331)) or (layer0_outputs(11825));
    layer1_outputs(6376) <= layer0_outputs(5003);
    layer1_outputs(6377) <= (layer0_outputs(8620)) and (layer0_outputs(11395));
    layer1_outputs(6378) <= '1';
    layer1_outputs(6379) <= (layer0_outputs(10867)) and (layer0_outputs(8892));
    layer1_outputs(6380) <= not(layer0_outputs(1317)) or (layer0_outputs(8665));
    layer1_outputs(6381) <= layer0_outputs(7690);
    layer1_outputs(6382) <= not((layer0_outputs(273)) and (layer0_outputs(5832)));
    layer1_outputs(6383) <= layer0_outputs(3611);
    layer1_outputs(6384) <= not(layer0_outputs(11304));
    layer1_outputs(6385) <= not((layer0_outputs(7931)) and (layer0_outputs(10559)));
    layer1_outputs(6386) <= not(layer0_outputs(2064)) or (layer0_outputs(8539));
    layer1_outputs(6387) <= layer0_outputs(11907);
    layer1_outputs(6388) <= (layer0_outputs(1289)) and not (layer0_outputs(10668));
    layer1_outputs(6389) <= not((layer0_outputs(5096)) xor (layer0_outputs(8729)));
    layer1_outputs(6390) <= not(layer0_outputs(8918)) or (layer0_outputs(4920));
    layer1_outputs(6391) <= not(layer0_outputs(10050));
    layer1_outputs(6392) <= (layer0_outputs(6437)) and not (layer0_outputs(1960));
    layer1_outputs(6393) <= not(layer0_outputs(10943)) or (layer0_outputs(1670));
    layer1_outputs(6394) <= not(layer0_outputs(5451)) or (layer0_outputs(11628));
    layer1_outputs(6395) <= layer0_outputs(5808);
    layer1_outputs(6396) <= (layer0_outputs(8130)) and not (layer0_outputs(9324));
    layer1_outputs(6397) <= not(layer0_outputs(9032));
    layer1_outputs(6398) <= (layer0_outputs(10425)) or (layer0_outputs(3249));
    layer1_outputs(6399) <= not(layer0_outputs(7842));
    layer1_outputs(6400) <= (layer0_outputs(1709)) xor (layer0_outputs(9307));
    layer1_outputs(6401) <= layer0_outputs(1438);
    layer1_outputs(6402) <= (layer0_outputs(9563)) and not (layer0_outputs(4534));
    layer1_outputs(6403) <= layer0_outputs(6209);
    layer1_outputs(6404) <= not(layer0_outputs(2011));
    layer1_outputs(6405) <= not((layer0_outputs(9805)) and (layer0_outputs(4062)));
    layer1_outputs(6406) <= (layer0_outputs(7276)) xor (layer0_outputs(8241));
    layer1_outputs(6407) <= layer0_outputs(6010);
    layer1_outputs(6408) <= layer0_outputs(10750);
    layer1_outputs(6409) <= (layer0_outputs(2510)) or (layer0_outputs(4362));
    layer1_outputs(6410) <= not(layer0_outputs(296)) or (layer0_outputs(10270));
    layer1_outputs(6411) <= layer0_outputs(9241);
    layer1_outputs(6412) <= not(layer0_outputs(12463)) or (layer0_outputs(1026));
    layer1_outputs(6413) <= (layer0_outputs(9248)) or (layer0_outputs(26));
    layer1_outputs(6414) <= layer0_outputs(134);
    layer1_outputs(6415) <= not((layer0_outputs(6139)) and (layer0_outputs(5326)));
    layer1_outputs(6416) <= layer0_outputs(3060);
    layer1_outputs(6417) <= not((layer0_outputs(8351)) or (layer0_outputs(5115)));
    layer1_outputs(6418) <= not(layer0_outputs(9657));
    layer1_outputs(6419) <= (layer0_outputs(4041)) and not (layer0_outputs(11985));
    layer1_outputs(6420) <= not(layer0_outputs(7750));
    layer1_outputs(6421) <= (layer0_outputs(8297)) xor (layer0_outputs(2115));
    layer1_outputs(6422) <= '0';
    layer1_outputs(6423) <= not((layer0_outputs(5431)) or (layer0_outputs(2149)));
    layer1_outputs(6424) <= not(layer0_outputs(797));
    layer1_outputs(6425) <= (layer0_outputs(8831)) and not (layer0_outputs(5615));
    layer1_outputs(6426) <= not(layer0_outputs(12437)) or (layer0_outputs(2541));
    layer1_outputs(6427) <= not(layer0_outputs(3536));
    layer1_outputs(6428) <= layer0_outputs(486);
    layer1_outputs(6429) <= layer0_outputs(11836);
    layer1_outputs(6430) <= (layer0_outputs(10353)) and not (layer0_outputs(8799));
    layer1_outputs(6431) <= layer0_outputs(895);
    layer1_outputs(6432) <= not(layer0_outputs(4659)) or (layer0_outputs(2278));
    layer1_outputs(6433) <= not((layer0_outputs(11008)) xor (layer0_outputs(11532)));
    layer1_outputs(6434) <= layer0_outputs(2609);
    layer1_outputs(6435) <= not(layer0_outputs(3743));
    layer1_outputs(6436) <= layer0_outputs(10158);
    layer1_outputs(6437) <= (layer0_outputs(9850)) or (layer0_outputs(368));
    layer1_outputs(6438) <= not(layer0_outputs(1949));
    layer1_outputs(6439) <= not((layer0_outputs(3912)) and (layer0_outputs(9198)));
    layer1_outputs(6440) <= not(layer0_outputs(7433)) or (layer0_outputs(5061));
    layer1_outputs(6441) <= not((layer0_outputs(4486)) or (layer0_outputs(1285)));
    layer1_outputs(6442) <= not(layer0_outputs(2408)) or (layer0_outputs(9658));
    layer1_outputs(6443) <= not(layer0_outputs(6738)) or (layer0_outputs(10720));
    layer1_outputs(6444) <= layer0_outputs(7465);
    layer1_outputs(6445) <= (layer0_outputs(8091)) and (layer0_outputs(9701));
    layer1_outputs(6446) <= layer0_outputs(1787);
    layer1_outputs(6447) <= not(layer0_outputs(12620));
    layer1_outputs(6448) <= not(layer0_outputs(10203));
    layer1_outputs(6449) <= (layer0_outputs(4588)) and not (layer0_outputs(12752));
    layer1_outputs(6450) <= (layer0_outputs(10514)) and not (layer0_outputs(6445));
    layer1_outputs(6451) <= (layer0_outputs(295)) or (layer0_outputs(6824));
    layer1_outputs(6452) <= (layer0_outputs(9413)) and (layer0_outputs(9284));
    layer1_outputs(6453) <= not((layer0_outputs(8771)) and (layer0_outputs(7076)));
    layer1_outputs(6454) <= (layer0_outputs(8348)) and not (layer0_outputs(9815));
    layer1_outputs(6455) <= layer0_outputs(5209);
    layer1_outputs(6456) <= not((layer0_outputs(11081)) xor (layer0_outputs(2993)));
    layer1_outputs(6457) <= (layer0_outputs(12768)) and not (layer0_outputs(136));
    layer1_outputs(6458) <= (layer0_outputs(8774)) and not (layer0_outputs(987));
    layer1_outputs(6459) <= layer0_outputs(1020);
    layer1_outputs(6460) <= not(layer0_outputs(12023)) or (layer0_outputs(561));
    layer1_outputs(6461) <= not(layer0_outputs(1031));
    layer1_outputs(6462) <= (layer0_outputs(1114)) and not (layer0_outputs(2533));
    layer1_outputs(6463) <= layer0_outputs(5559);
    layer1_outputs(6464) <= layer0_outputs(7822);
    layer1_outputs(6465) <= layer0_outputs(1699);
    layer1_outputs(6466) <= not(layer0_outputs(9713));
    layer1_outputs(6467) <= (layer0_outputs(6973)) or (layer0_outputs(9340));
    layer1_outputs(6468) <= (layer0_outputs(9014)) xor (layer0_outputs(10137));
    layer1_outputs(6469) <= not(layer0_outputs(12026));
    layer1_outputs(6470) <= not(layer0_outputs(5861)) or (layer0_outputs(6363));
    layer1_outputs(6471) <= not((layer0_outputs(7406)) and (layer0_outputs(3706)));
    layer1_outputs(6472) <= not(layer0_outputs(1205));
    layer1_outputs(6473) <= not(layer0_outputs(8065));
    layer1_outputs(6474) <= not((layer0_outputs(7170)) or (layer0_outputs(5224)));
    layer1_outputs(6475) <= not((layer0_outputs(7133)) and (layer0_outputs(3666)));
    layer1_outputs(6476) <= (layer0_outputs(3485)) and not (layer0_outputs(11061));
    layer1_outputs(6477) <= (layer0_outputs(7114)) or (layer0_outputs(8087));
    layer1_outputs(6478) <= (layer0_outputs(3392)) or (layer0_outputs(8887));
    layer1_outputs(6479) <= (layer0_outputs(3872)) xor (layer0_outputs(11662));
    layer1_outputs(6480) <= not(layer0_outputs(1016)) or (layer0_outputs(11137));
    layer1_outputs(6481) <= '1';
    layer1_outputs(6482) <= not(layer0_outputs(6012)) or (layer0_outputs(4691));
    layer1_outputs(6483) <= not((layer0_outputs(5640)) xor (layer0_outputs(3747)));
    layer1_outputs(6484) <= '1';
    layer1_outputs(6485) <= not(layer0_outputs(1049));
    layer1_outputs(6486) <= layer0_outputs(1544);
    layer1_outputs(6487) <= (layer0_outputs(2030)) and (layer0_outputs(2545));
    layer1_outputs(6488) <= not((layer0_outputs(6505)) xor (layer0_outputs(1076)));
    layer1_outputs(6489) <= not(layer0_outputs(5555));
    layer1_outputs(6490) <= not(layer0_outputs(4073));
    layer1_outputs(6491) <= not(layer0_outputs(11889));
    layer1_outputs(6492) <= (layer0_outputs(1243)) and not (layer0_outputs(9958));
    layer1_outputs(6493) <= not(layer0_outputs(347)) or (layer0_outputs(8285));
    layer1_outputs(6494) <= not(layer0_outputs(8610));
    layer1_outputs(6495) <= (layer0_outputs(8740)) and not (layer0_outputs(8857));
    layer1_outputs(6496) <= not(layer0_outputs(9756));
    layer1_outputs(6497) <= not(layer0_outputs(6455)) or (layer0_outputs(2637));
    layer1_outputs(6498) <= (layer0_outputs(12214)) xor (layer0_outputs(3205));
    layer1_outputs(6499) <= not(layer0_outputs(6512));
    layer1_outputs(6500) <= not(layer0_outputs(3612));
    layer1_outputs(6501) <= (layer0_outputs(1188)) and not (layer0_outputs(3143));
    layer1_outputs(6502) <= layer0_outputs(11134);
    layer1_outputs(6503) <= layer0_outputs(1230);
    layer1_outputs(6504) <= (layer0_outputs(5886)) and not (layer0_outputs(8405));
    layer1_outputs(6505) <= not(layer0_outputs(3498));
    layer1_outputs(6506) <= not(layer0_outputs(9));
    layer1_outputs(6507) <= layer0_outputs(5871);
    layer1_outputs(6508) <= (layer0_outputs(8606)) or (layer0_outputs(1901));
    layer1_outputs(6509) <= (layer0_outputs(8774)) and not (layer0_outputs(9888));
    layer1_outputs(6510) <= not(layer0_outputs(7758));
    layer1_outputs(6511) <= not((layer0_outputs(8487)) xor (layer0_outputs(1603)));
    layer1_outputs(6512) <= not(layer0_outputs(5479));
    layer1_outputs(6513) <= layer0_outputs(10836);
    layer1_outputs(6514) <= (layer0_outputs(9663)) and not (layer0_outputs(10475));
    layer1_outputs(6515) <= (layer0_outputs(7223)) and not (layer0_outputs(5673));
    layer1_outputs(6516) <= not(layer0_outputs(11642)) or (layer0_outputs(6613));
    layer1_outputs(6517) <= (layer0_outputs(9113)) and not (layer0_outputs(7959));
    layer1_outputs(6518) <= not(layer0_outputs(4066));
    layer1_outputs(6519) <= (layer0_outputs(11412)) xor (layer0_outputs(3235));
    layer1_outputs(6520) <= layer0_outputs(5583);
    layer1_outputs(6521) <= not((layer0_outputs(2811)) xor (layer0_outputs(269)));
    layer1_outputs(6522) <= (layer0_outputs(4514)) or (layer0_outputs(9963));
    layer1_outputs(6523) <= layer0_outputs(5451);
    layer1_outputs(6524) <= layer0_outputs(12704);
    layer1_outputs(6525) <= not(layer0_outputs(9156));
    layer1_outputs(6526) <= layer0_outputs(4694);
    layer1_outputs(6527) <= (layer0_outputs(12765)) and (layer0_outputs(807));
    layer1_outputs(6528) <= not((layer0_outputs(1231)) or (layer0_outputs(2328)));
    layer1_outputs(6529) <= (layer0_outputs(11469)) and not (layer0_outputs(8479));
    layer1_outputs(6530) <= '0';
    layer1_outputs(6531) <= (layer0_outputs(878)) and (layer0_outputs(8287));
    layer1_outputs(6532) <= not((layer0_outputs(4609)) and (layer0_outputs(1521)));
    layer1_outputs(6533) <= not(layer0_outputs(12591));
    layer1_outputs(6534) <= (layer0_outputs(4100)) and not (layer0_outputs(2575));
    layer1_outputs(6535) <= (layer0_outputs(12245)) and (layer0_outputs(6463));
    layer1_outputs(6536) <= not((layer0_outputs(6124)) or (layer0_outputs(9240)));
    layer1_outputs(6537) <= (layer0_outputs(6373)) and not (layer0_outputs(184));
    layer1_outputs(6538) <= not((layer0_outputs(869)) and (layer0_outputs(11924)));
    layer1_outputs(6539) <= layer0_outputs(10479);
    layer1_outputs(6540) <= not((layer0_outputs(10691)) and (layer0_outputs(8070)));
    layer1_outputs(6541) <= not((layer0_outputs(5244)) xor (layer0_outputs(6107)));
    layer1_outputs(6542) <= not(layer0_outputs(12791)) or (layer0_outputs(4220));
    layer1_outputs(6543) <= layer0_outputs(1215);
    layer1_outputs(6544) <= layer0_outputs(3075);
    layer1_outputs(6545) <= layer0_outputs(6042);
    layer1_outputs(6546) <= not((layer0_outputs(1023)) or (layer0_outputs(6628)));
    layer1_outputs(6547) <= not((layer0_outputs(342)) or (layer0_outputs(11527)));
    layer1_outputs(6548) <= layer0_outputs(11626);
    layer1_outputs(6549) <= '0';
    layer1_outputs(6550) <= layer0_outputs(4673);
    layer1_outputs(6551) <= (layer0_outputs(3699)) xor (layer0_outputs(10785));
    layer1_outputs(6552) <= not((layer0_outputs(12025)) and (layer0_outputs(2518)));
    layer1_outputs(6553) <= '1';
    layer1_outputs(6554) <= layer0_outputs(300);
    layer1_outputs(6555) <= (layer0_outputs(1213)) or (layer0_outputs(9479));
    layer1_outputs(6556) <= (layer0_outputs(8850)) and not (layer0_outputs(751));
    layer1_outputs(6557) <= not((layer0_outputs(6976)) and (layer0_outputs(9637)));
    layer1_outputs(6558) <= (layer0_outputs(11403)) and not (layer0_outputs(9162));
    layer1_outputs(6559) <= (layer0_outputs(10218)) xor (layer0_outputs(8099));
    layer1_outputs(6560) <= (layer0_outputs(938)) and not (layer0_outputs(8067));
    layer1_outputs(6561) <= (layer0_outputs(5760)) and not (layer0_outputs(94));
    layer1_outputs(6562) <= not(layer0_outputs(9353));
    layer1_outputs(6563) <= not(layer0_outputs(460)) or (layer0_outputs(10897));
    layer1_outputs(6564) <= layer0_outputs(8436);
    layer1_outputs(6565) <= (layer0_outputs(2209)) and not (layer0_outputs(4900));
    layer1_outputs(6566) <= layer0_outputs(3964);
    layer1_outputs(6567) <= not(layer0_outputs(9016));
    layer1_outputs(6568) <= (layer0_outputs(12008)) or (layer0_outputs(985));
    layer1_outputs(6569) <= layer0_outputs(9716);
    layer1_outputs(6570) <= not((layer0_outputs(7297)) or (layer0_outputs(7824)));
    layer1_outputs(6571) <= not(layer0_outputs(12347));
    layer1_outputs(6572) <= layer0_outputs(9666);
    layer1_outputs(6573) <= not(layer0_outputs(8967));
    layer1_outputs(6574) <= (layer0_outputs(1692)) and not (layer0_outputs(3828));
    layer1_outputs(6575) <= not((layer0_outputs(5887)) or (layer0_outputs(8815)));
    layer1_outputs(6576) <= (layer0_outputs(6872)) and not (layer0_outputs(7541));
    layer1_outputs(6577) <= (layer0_outputs(2049)) and not (layer0_outputs(336));
    layer1_outputs(6578) <= not((layer0_outputs(5856)) and (layer0_outputs(1744)));
    layer1_outputs(6579) <= layer0_outputs(10307);
    layer1_outputs(6580) <= layer0_outputs(12150);
    layer1_outputs(6581) <= not((layer0_outputs(7638)) and (layer0_outputs(6703)));
    layer1_outputs(6582) <= not(layer0_outputs(5724));
    layer1_outputs(6583) <= not(layer0_outputs(4954)) or (layer0_outputs(9098));
    layer1_outputs(6584) <= (layer0_outputs(8342)) xor (layer0_outputs(10409));
    layer1_outputs(6585) <= layer0_outputs(10404);
    layer1_outputs(6586) <= not(layer0_outputs(512)) or (layer0_outputs(1809));
    layer1_outputs(6587) <= (layer0_outputs(5971)) or (layer0_outputs(4574));
    layer1_outputs(6588) <= layer0_outputs(6390);
    layer1_outputs(6589) <= not((layer0_outputs(10619)) or (layer0_outputs(12326)));
    layer1_outputs(6590) <= not(layer0_outputs(3927)) or (layer0_outputs(11697));
    layer1_outputs(6591) <= not(layer0_outputs(6447)) or (layer0_outputs(2383));
    layer1_outputs(6592) <= (layer0_outputs(9149)) or (layer0_outputs(9392));
    layer1_outputs(6593) <= not(layer0_outputs(1224));
    layer1_outputs(6594) <= (layer0_outputs(4015)) xor (layer0_outputs(11785));
    layer1_outputs(6595) <= '1';
    layer1_outputs(6596) <= (layer0_outputs(11126)) and not (layer0_outputs(2615));
    layer1_outputs(6597) <= layer0_outputs(10259);
    layer1_outputs(6598) <= not((layer0_outputs(8685)) or (layer0_outputs(2090)));
    layer1_outputs(6599) <= layer0_outputs(10085);
    layer1_outputs(6600) <= (layer0_outputs(10383)) and not (layer0_outputs(11940));
    layer1_outputs(6601) <= layer0_outputs(751);
    layer1_outputs(6602) <= not(layer0_outputs(1655));
    layer1_outputs(6603) <= (layer0_outputs(4101)) xor (layer0_outputs(7659));
    layer1_outputs(6604) <= layer0_outputs(3244);
    layer1_outputs(6605) <= (layer0_outputs(6818)) or (layer0_outputs(410));
    layer1_outputs(6606) <= not(layer0_outputs(12405)) or (layer0_outputs(2345));
    layer1_outputs(6607) <= (layer0_outputs(3868)) xor (layer0_outputs(2110));
    layer1_outputs(6608) <= (layer0_outputs(10631)) xor (layer0_outputs(3282));
    layer1_outputs(6609) <= '1';
    layer1_outputs(6610) <= layer0_outputs(3900);
    layer1_outputs(6611) <= layer0_outputs(2752);
    layer1_outputs(6612) <= layer0_outputs(3963);
    layer1_outputs(6613) <= not(layer0_outputs(6966)) or (layer0_outputs(10351));
    layer1_outputs(6614) <= not(layer0_outputs(989));
    layer1_outputs(6615) <= layer0_outputs(11402);
    layer1_outputs(6616) <= not(layer0_outputs(1051)) or (layer0_outputs(626));
    layer1_outputs(6617) <= layer0_outputs(8613);
    layer1_outputs(6618) <= (layer0_outputs(10726)) and (layer0_outputs(3119));
    layer1_outputs(6619) <= (layer0_outputs(9195)) and (layer0_outputs(7713));
    layer1_outputs(6620) <= not((layer0_outputs(3797)) or (layer0_outputs(1453)));
    layer1_outputs(6621) <= not(layer0_outputs(1708));
    layer1_outputs(6622) <= not(layer0_outputs(2837));
    layer1_outputs(6623) <= not(layer0_outputs(7289));
    layer1_outputs(6624) <= layer0_outputs(6908);
    layer1_outputs(6625) <= '1';
    layer1_outputs(6626) <= not((layer0_outputs(2710)) xor (layer0_outputs(9596)));
    layer1_outputs(6627) <= (layer0_outputs(11587)) or (layer0_outputs(4365));
    layer1_outputs(6628) <= not(layer0_outputs(36)) or (layer0_outputs(9097));
    layer1_outputs(6629) <= not(layer0_outputs(4316)) or (layer0_outputs(2219));
    layer1_outputs(6630) <= not((layer0_outputs(4948)) or (layer0_outputs(6267)));
    layer1_outputs(6631) <= not(layer0_outputs(7119)) or (layer0_outputs(1616));
    layer1_outputs(6632) <= layer0_outputs(10680);
    layer1_outputs(6633) <= not(layer0_outputs(9476));
    layer1_outputs(6634) <= not(layer0_outputs(1040));
    layer1_outputs(6635) <= not(layer0_outputs(2575)) or (layer0_outputs(4858));
    layer1_outputs(6636) <= not(layer0_outputs(10325));
    layer1_outputs(6637) <= not(layer0_outputs(7398)) or (layer0_outputs(9603));
    layer1_outputs(6638) <= not((layer0_outputs(6552)) and (layer0_outputs(1939)));
    layer1_outputs(6639) <= (layer0_outputs(9893)) and (layer0_outputs(10052));
    layer1_outputs(6640) <= (layer0_outputs(3023)) or (layer0_outputs(3509));
    layer1_outputs(6641) <= layer0_outputs(6753);
    layer1_outputs(6642) <= not(layer0_outputs(8734)) or (layer0_outputs(355));
    layer1_outputs(6643) <= not(layer0_outputs(10565));
    layer1_outputs(6644) <= layer0_outputs(3206);
    layer1_outputs(6645) <= layer0_outputs(4033);
    layer1_outputs(6646) <= layer0_outputs(8992);
    layer1_outputs(6647) <= (layer0_outputs(7405)) or (layer0_outputs(8329));
    layer1_outputs(6648) <= not((layer0_outputs(3186)) and (layer0_outputs(11218)));
    layer1_outputs(6649) <= layer0_outputs(12386);
    layer1_outputs(6650) <= not((layer0_outputs(160)) and (layer0_outputs(6787)));
    layer1_outputs(6651) <= not(layer0_outputs(8437)) or (layer0_outputs(654));
    layer1_outputs(6652) <= '1';
    layer1_outputs(6653) <= layer0_outputs(6113);
    layer1_outputs(6654) <= not((layer0_outputs(7345)) and (layer0_outputs(5801)));
    layer1_outputs(6655) <= layer0_outputs(4421);
    layer1_outputs(6656) <= (layer0_outputs(9591)) xor (layer0_outputs(3727));
    layer1_outputs(6657) <= not((layer0_outputs(790)) and (layer0_outputs(6412)));
    layer1_outputs(6658) <= not((layer0_outputs(6026)) or (layer0_outputs(5343)));
    layer1_outputs(6659) <= not(layer0_outputs(8752));
    layer1_outputs(6660) <= not((layer0_outputs(5994)) and (layer0_outputs(3901)));
    layer1_outputs(6661) <= not((layer0_outputs(2582)) or (layer0_outputs(10634)));
    layer1_outputs(6662) <= not(layer0_outputs(4930));
    layer1_outputs(6663) <= not((layer0_outputs(5323)) xor (layer0_outputs(2088)));
    layer1_outputs(6664) <= not(layer0_outputs(11344));
    layer1_outputs(6665) <= (layer0_outputs(988)) and not (layer0_outputs(1853));
    layer1_outputs(6666) <= layer0_outputs(372);
    layer1_outputs(6667) <= (layer0_outputs(8133)) xor (layer0_outputs(4530));
    layer1_outputs(6668) <= (layer0_outputs(1861)) and not (layer0_outputs(2507));
    layer1_outputs(6669) <= '0';
    layer1_outputs(6670) <= layer0_outputs(12572);
    layer1_outputs(6671) <= layer0_outputs(6075);
    layer1_outputs(6672) <= layer0_outputs(11352);
    layer1_outputs(6673) <= not((layer0_outputs(2670)) and (layer0_outputs(12027)));
    layer1_outputs(6674) <= not((layer0_outputs(9358)) and (layer0_outputs(938)));
    layer1_outputs(6675) <= not(layer0_outputs(722));
    layer1_outputs(6676) <= layer0_outputs(4014);
    layer1_outputs(6677) <= layer0_outputs(5183);
    layer1_outputs(6678) <= layer0_outputs(638);
    layer1_outputs(6679) <= not(layer0_outputs(328)) or (layer0_outputs(1559));
    layer1_outputs(6680) <= not(layer0_outputs(12505)) or (layer0_outputs(6255));
    layer1_outputs(6681) <= (layer0_outputs(12414)) xor (layer0_outputs(1175));
    layer1_outputs(6682) <= (layer0_outputs(8109)) and (layer0_outputs(10699));
    layer1_outputs(6683) <= (layer0_outputs(256)) and (layer0_outputs(3037));
    layer1_outputs(6684) <= not((layer0_outputs(11538)) xor (layer0_outputs(5223)));
    layer1_outputs(6685) <= not(layer0_outputs(9179));
    layer1_outputs(6686) <= (layer0_outputs(10526)) and not (layer0_outputs(11965));
    layer1_outputs(6687) <= layer0_outputs(2824);
    layer1_outputs(6688) <= (layer0_outputs(10072)) and not (layer0_outputs(11042));
    layer1_outputs(6689) <= (layer0_outputs(5635)) and not (layer0_outputs(12678));
    layer1_outputs(6690) <= (layer0_outputs(5261)) and (layer0_outputs(8696));
    layer1_outputs(6691) <= not((layer0_outputs(7736)) and (layer0_outputs(6694)));
    layer1_outputs(6692) <= not(layer0_outputs(21)) or (layer0_outputs(3908));
    layer1_outputs(6693) <= not(layer0_outputs(1730));
    layer1_outputs(6694) <= (layer0_outputs(1393)) or (layer0_outputs(12441));
    layer1_outputs(6695) <= layer0_outputs(6800);
    layer1_outputs(6696) <= not((layer0_outputs(4396)) or (layer0_outputs(2854)));
    layer1_outputs(6697) <= layer0_outputs(2427);
    layer1_outputs(6698) <= not(layer0_outputs(4196));
    layer1_outputs(6699) <= '0';
    layer1_outputs(6700) <= not((layer0_outputs(10748)) or (layer0_outputs(2901)));
    layer1_outputs(6701) <= not(layer0_outputs(7152));
    layer1_outputs(6702) <= (layer0_outputs(8432)) or (layer0_outputs(9304));
    layer1_outputs(6703) <= layer0_outputs(11144);
    layer1_outputs(6704) <= (layer0_outputs(9347)) and (layer0_outputs(146));
    layer1_outputs(6705) <= not((layer0_outputs(3144)) xor (layer0_outputs(850)));
    layer1_outputs(6706) <= (layer0_outputs(1716)) or (layer0_outputs(8959));
    layer1_outputs(6707) <= not(layer0_outputs(5250)) or (layer0_outputs(10267));
    layer1_outputs(6708) <= not(layer0_outputs(9141));
    layer1_outputs(6709) <= (layer0_outputs(8565)) and (layer0_outputs(3381));
    layer1_outputs(6710) <= not((layer0_outputs(12098)) or (layer0_outputs(6406)));
    layer1_outputs(6711) <= (layer0_outputs(2035)) and (layer0_outputs(619));
    layer1_outputs(6712) <= not(layer0_outputs(9420));
    layer1_outputs(6713) <= (layer0_outputs(7169)) and (layer0_outputs(9626));
    layer1_outputs(6714) <= layer0_outputs(6786);
    layer1_outputs(6715) <= layer0_outputs(11095);
    layer1_outputs(6716) <= (layer0_outputs(12445)) xor (layer0_outputs(4382));
    layer1_outputs(6717) <= layer0_outputs(8253);
    layer1_outputs(6718) <= layer0_outputs(10086);
    layer1_outputs(6719) <= layer0_outputs(2833);
    layer1_outputs(6720) <= (layer0_outputs(1770)) xor (layer0_outputs(6644));
    layer1_outputs(6721) <= not(layer0_outputs(8210));
    layer1_outputs(6722) <= not((layer0_outputs(666)) and (layer0_outputs(9769)));
    layer1_outputs(6723) <= (layer0_outputs(10918)) and not (layer0_outputs(8333));
    layer1_outputs(6724) <= not((layer0_outputs(9697)) xor (layer0_outputs(6933)));
    layer1_outputs(6725) <= (layer0_outputs(12298)) or (layer0_outputs(8505));
    layer1_outputs(6726) <= not((layer0_outputs(11232)) and (layer0_outputs(3444)));
    layer1_outputs(6727) <= layer0_outputs(527);
    layer1_outputs(6728) <= (layer0_outputs(11277)) and not (layer0_outputs(3574));
    layer1_outputs(6729) <= (layer0_outputs(2299)) and (layer0_outputs(11221));
    layer1_outputs(6730) <= layer0_outputs(10002);
    layer1_outputs(6731) <= not(layer0_outputs(413));
    layer1_outputs(6732) <= (layer0_outputs(10258)) and not (layer0_outputs(7274));
    layer1_outputs(6733) <= layer0_outputs(26);
    layer1_outputs(6734) <= not(layer0_outputs(3009));
    layer1_outputs(6735) <= not(layer0_outputs(11680)) or (layer0_outputs(3627));
    layer1_outputs(6736) <= (layer0_outputs(11483)) or (layer0_outputs(9166));
    layer1_outputs(6737) <= not(layer0_outputs(1586));
    layer1_outputs(6738) <= not(layer0_outputs(3624)) or (layer0_outputs(8002));
    layer1_outputs(6739) <= (layer0_outputs(1121)) and (layer0_outputs(1206));
    layer1_outputs(6740) <= (layer0_outputs(7849)) and not (layer0_outputs(12409));
    layer1_outputs(6741) <= layer0_outputs(3313);
    layer1_outputs(6742) <= layer0_outputs(1816);
    layer1_outputs(6743) <= not(layer0_outputs(11219)) or (layer0_outputs(9436));
    layer1_outputs(6744) <= not((layer0_outputs(451)) or (layer0_outputs(2282)));
    layer1_outputs(6745) <= (layer0_outputs(794)) or (layer0_outputs(3909));
    layer1_outputs(6746) <= '1';
    layer1_outputs(6747) <= not(layer0_outputs(9758)) or (layer0_outputs(12548));
    layer1_outputs(6748) <= not((layer0_outputs(5116)) xor (layer0_outputs(10998)));
    layer1_outputs(6749) <= not(layer0_outputs(477));
    layer1_outputs(6750) <= (layer0_outputs(2897)) and not (layer0_outputs(680));
    layer1_outputs(6751) <= layer0_outputs(2828);
    layer1_outputs(6752) <= (layer0_outputs(3534)) or (layer0_outputs(1612));
    layer1_outputs(6753) <= not(layer0_outputs(4174));
    layer1_outputs(6754) <= not(layer0_outputs(4832));
    layer1_outputs(6755) <= (layer0_outputs(9224)) or (layer0_outputs(1210));
    layer1_outputs(6756) <= (layer0_outputs(3137)) xor (layer0_outputs(7212));
    layer1_outputs(6757) <= not(layer0_outputs(5227)) or (layer0_outputs(5739));
    layer1_outputs(6758) <= (layer0_outputs(10856)) and (layer0_outputs(10415));
    layer1_outputs(6759) <= layer0_outputs(8848);
    layer1_outputs(6760) <= (layer0_outputs(11941)) and not (layer0_outputs(5561));
    layer1_outputs(6761) <= (layer0_outputs(10254)) or (layer0_outputs(10442));
    layer1_outputs(6762) <= not(layer0_outputs(8530)) or (layer0_outputs(12717));
    layer1_outputs(6763) <= (layer0_outputs(3854)) or (layer0_outputs(11834));
    layer1_outputs(6764) <= layer0_outputs(3114);
    layer1_outputs(6765) <= layer0_outputs(5422);
    layer1_outputs(6766) <= (layer0_outputs(8288)) and not (layer0_outputs(7231));
    layer1_outputs(6767) <= (layer0_outputs(9215)) and (layer0_outputs(2722));
    layer1_outputs(6768) <= (layer0_outputs(6667)) xor (layer0_outputs(7866));
    layer1_outputs(6769) <= not(layer0_outputs(11130)) or (layer0_outputs(3644));
    layer1_outputs(6770) <= '0';
    layer1_outputs(6771) <= not(layer0_outputs(10443)) or (layer0_outputs(9688));
    layer1_outputs(6772) <= not((layer0_outputs(6795)) and (layer0_outputs(3421)));
    layer1_outputs(6773) <= (layer0_outputs(313)) and (layer0_outputs(5171));
    layer1_outputs(6774) <= not(layer0_outputs(10603));
    layer1_outputs(6775) <= layer0_outputs(3032);
    layer1_outputs(6776) <= layer0_outputs(4117);
    layer1_outputs(6777) <= layer0_outputs(12471);
    layer1_outputs(6778) <= not(layer0_outputs(545));
    layer1_outputs(6779) <= layer0_outputs(1926);
    layer1_outputs(6780) <= not((layer0_outputs(924)) and (layer0_outputs(1037)));
    layer1_outputs(6781) <= not(layer0_outputs(3179)) or (layer0_outputs(2311));
    layer1_outputs(6782) <= not(layer0_outputs(5637));
    layer1_outputs(6783) <= layer0_outputs(6683);
    layer1_outputs(6784) <= not(layer0_outputs(7885));
    layer1_outputs(6785) <= layer0_outputs(10069);
    layer1_outputs(6786) <= not((layer0_outputs(5935)) or (layer0_outputs(2040)));
    layer1_outputs(6787) <= (layer0_outputs(12528)) and not (layer0_outputs(5863));
    layer1_outputs(6788) <= layer0_outputs(5431);
    layer1_outputs(6789) <= (layer0_outputs(5783)) and (layer0_outputs(2131));
    layer1_outputs(6790) <= not(layer0_outputs(1264)) or (layer0_outputs(5356));
    layer1_outputs(6791) <= (layer0_outputs(9617)) xor (layer0_outputs(5455));
    layer1_outputs(6792) <= not((layer0_outputs(11891)) and (layer0_outputs(8814)));
    layer1_outputs(6793) <= (layer0_outputs(837)) xor (layer0_outputs(10698));
    layer1_outputs(6794) <= layer0_outputs(3089);
    layer1_outputs(6795) <= not(layer0_outputs(425));
    layer1_outputs(6796) <= not(layer0_outputs(1058));
    layer1_outputs(6797) <= not(layer0_outputs(4444));
    layer1_outputs(6798) <= layer0_outputs(3394);
    layer1_outputs(6799) <= not(layer0_outputs(11123));
    layer1_outputs(6800) <= not(layer0_outputs(6357));
    layer1_outputs(6801) <= not(layer0_outputs(767));
    layer1_outputs(6802) <= (layer0_outputs(653)) and not (layer0_outputs(899));
    layer1_outputs(6803) <= (layer0_outputs(12572)) and not (layer0_outputs(6784));
    layer1_outputs(6804) <= not(layer0_outputs(3098));
    layer1_outputs(6805) <= (layer0_outputs(53)) and not (layer0_outputs(9872));
    layer1_outputs(6806) <= (layer0_outputs(4274)) or (layer0_outputs(8135));
    layer1_outputs(6807) <= layer0_outputs(1221);
    layer1_outputs(6808) <= layer0_outputs(10950);
    layer1_outputs(6809) <= not(layer0_outputs(2934));
    layer1_outputs(6810) <= layer0_outputs(8563);
    layer1_outputs(6811) <= not(layer0_outputs(9641));
    layer1_outputs(6812) <= (layer0_outputs(7051)) and (layer0_outputs(7742));
    layer1_outputs(6813) <= not((layer0_outputs(9005)) or (layer0_outputs(9205)));
    layer1_outputs(6814) <= (layer0_outputs(4224)) xor (layer0_outputs(772));
    layer1_outputs(6815) <= not(layer0_outputs(7901));
    layer1_outputs(6816) <= layer0_outputs(8667);
    layer1_outputs(6817) <= (layer0_outputs(7477)) and not (layer0_outputs(2072));
    layer1_outputs(6818) <= (layer0_outputs(8103)) and not (layer0_outputs(5885));
    layer1_outputs(6819) <= layer0_outputs(2679);
    layer1_outputs(6820) <= not(layer0_outputs(2354));
    layer1_outputs(6821) <= not(layer0_outputs(6537));
    layer1_outputs(6822) <= (layer0_outputs(3672)) and not (layer0_outputs(6369));
    layer1_outputs(6823) <= not(layer0_outputs(3642));
    layer1_outputs(6824) <= (layer0_outputs(6481)) and (layer0_outputs(7486));
    layer1_outputs(6825) <= not((layer0_outputs(9932)) and (layer0_outputs(839)));
    layer1_outputs(6826) <= not(layer0_outputs(7589));
    layer1_outputs(6827) <= layer0_outputs(9165);
    layer1_outputs(6828) <= not(layer0_outputs(9488)) or (layer0_outputs(5641));
    layer1_outputs(6829) <= (layer0_outputs(6177)) or (layer0_outputs(4186));
    layer1_outputs(6830) <= not(layer0_outputs(2742));
    layer1_outputs(6831) <= not(layer0_outputs(10948)) or (layer0_outputs(2020));
    layer1_outputs(6832) <= (layer0_outputs(750)) xor (layer0_outputs(10718));
    layer1_outputs(6833) <= not((layer0_outputs(6668)) and (layer0_outputs(2396)));
    layer1_outputs(6834) <= not(layer0_outputs(9615));
    layer1_outputs(6835) <= not((layer0_outputs(8870)) or (layer0_outputs(652)));
    layer1_outputs(6836) <= not(layer0_outputs(603)) or (layer0_outputs(5508));
    layer1_outputs(6837) <= not(layer0_outputs(11419)) or (layer0_outputs(7044));
    layer1_outputs(6838) <= not(layer0_outputs(3339));
    layer1_outputs(6839) <= not(layer0_outputs(2116)) or (layer0_outputs(11364));
    layer1_outputs(6840) <= not(layer0_outputs(7912)) or (layer0_outputs(7879));
    layer1_outputs(6841) <= not(layer0_outputs(9696)) or (layer0_outputs(5894));
    layer1_outputs(6842) <= not(layer0_outputs(2524)) or (layer0_outputs(7579));
    layer1_outputs(6843) <= layer0_outputs(8041);
    layer1_outputs(6844) <= (layer0_outputs(5721)) and (layer0_outputs(1796));
    layer1_outputs(6845) <= (layer0_outputs(3870)) xor (layer0_outputs(8542));
    layer1_outputs(6846) <= not(layer0_outputs(539)) or (layer0_outputs(9038));
    layer1_outputs(6847) <= (layer0_outputs(12352)) or (layer0_outputs(2480));
    layer1_outputs(6848) <= not((layer0_outputs(850)) or (layer0_outputs(1050)));
    layer1_outputs(6849) <= not(layer0_outputs(3300));
    layer1_outputs(6850) <= not(layer0_outputs(6565));
    layer1_outputs(6851) <= (layer0_outputs(6868)) or (layer0_outputs(6805));
    layer1_outputs(6852) <= (layer0_outputs(11421)) and not (layer0_outputs(5439));
    layer1_outputs(6853) <= not(layer0_outputs(1572)) or (layer0_outputs(9395));
    layer1_outputs(6854) <= not((layer0_outputs(10880)) and (layer0_outputs(12575)));
    layer1_outputs(6855) <= layer0_outputs(10682);
    layer1_outputs(6856) <= (layer0_outputs(3637)) and not (layer0_outputs(12009));
    layer1_outputs(6857) <= layer0_outputs(7000);
    layer1_outputs(6858) <= not(layer0_outputs(11724));
    layer1_outputs(6859) <= not((layer0_outputs(11896)) and (layer0_outputs(9531)));
    layer1_outputs(6860) <= '0';
    layer1_outputs(6861) <= layer0_outputs(6828);
    layer1_outputs(6862) <= (layer0_outputs(11758)) and not (layer0_outputs(9714));
    layer1_outputs(6863) <= not((layer0_outputs(8451)) and (layer0_outputs(9002)));
    layer1_outputs(6864) <= not(layer0_outputs(8343));
    layer1_outputs(6865) <= layer0_outputs(2159);
    layer1_outputs(6866) <= not(layer0_outputs(8855)) or (layer0_outputs(1516));
    layer1_outputs(6867) <= not(layer0_outputs(10311));
    layer1_outputs(6868) <= layer0_outputs(9640);
    layer1_outputs(6869) <= layer0_outputs(8754);
    layer1_outputs(6870) <= (layer0_outputs(1192)) and (layer0_outputs(8460));
    layer1_outputs(6871) <= layer0_outputs(875);
    layer1_outputs(6872) <= not(layer0_outputs(1125));
    layer1_outputs(6873) <= (layer0_outputs(6968)) or (layer0_outputs(10344));
    layer1_outputs(6874) <= not(layer0_outputs(8353)) or (layer0_outputs(11480));
    layer1_outputs(6875) <= not(layer0_outputs(7652)) or (layer0_outputs(9766));
    layer1_outputs(6876) <= (layer0_outputs(3893)) and not (layer0_outputs(6207));
    layer1_outputs(6877) <= not(layer0_outputs(12294));
    layer1_outputs(6878) <= not((layer0_outputs(7639)) and (layer0_outputs(1674)));
    layer1_outputs(6879) <= (layer0_outputs(8765)) or (layer0_outputs(5257));
    layer1_outputs(6880) <= layer0_outputs(6426);
    layer1_outputs(6881) <= (layer0_outputs(4493)) and not (layer0_outputs(9296));
    layer1_outputs(6882) <= not(layer0_outputs(1253)) or (layer0_outputs(7041));
    layer1_outputs(6883) <= not(layer0_outputs(4149)) or (layer0_outputs(9415));
    layer1_outputs(6884) <= (layer0_outputs(9064)) and not (layer0_outputs(6783));
    layer1_outputs(6885) <= not((layer0_outputs(5578)) xor (layer0_outputs(2643)));
    layer1_outputs(6886) <= (layer0_outputs(9378)) or (layer0_outputs(10836));
    layer1_outputs(6887) <= not((layer0_outputs(12713)) xor (layer0_outputs(3571)));
    layer1_outputs(6888) <= not((layer0_outputs(5843)) and (layer0_outputs(7634)));
    layer1_outputs(6889) <= (layer0_outputs(10140)) and not (layer0_outputs(7158));
    layer1_outputs(6890) <= not((layer0_outputs(2685)) or (layer0_outputs(1032)));
    layer1_outputs(6891) <= not(layer0_outputs(4095));
    layer1_outputs(6892) <= not(layer0_outputs(10437));
    layer1_outputs(6893) <= not(layer0_outputs(5975));
    layer1_outputs(6894) <= not(layer0_outputs(11877));
    layer1_outputs(6895) <= layer0_outputs(1110);
    layer1_outputs(6896) <= layer0_outputs(8501);
    layer1_outputs(6897) <= (layer0_outputs(4768)) or (layer0_outputs(1108));
    layer1_outputs(6898) <= (layer0_outputs(4851)) xor (layer0_outputs(9336));
    layer1_outputs(6899) <= layer0_outputs(10048);
    layer1_outputs(6900) <= not(layer0_outputs(2745));
    layer1_outputs(6901) <= not((layer0_outputs(4392)) and (layer0_outputs(4921)));
    layer1_outputs(6902) <= layer0_outputs(5350);
    layer1_outputs(6903) <= not((layer0_outputs(3757)) or (layer0_outputs(52)));
    layer1_outputs(6904) <= not(layer0_outputs(9727)) or (layer0_outputs(442));
    layer1_outputs(6905) <= '0';
    layer1_outputs(6906) <= (layer0_outputs(7035)) and not (layer0_outputs(3749));
    layer1_outputs(6907) <= layer0_outputs(11768);
    layer1_outputs(6908) <= not((layer0_outputs(8880)) or (layer0_outputs(12280)));
    layer1_outputs(6909) <= (layer0_outputs(12323)) xor (layer0_outputs(5962));
    layer1_outputs(6910) <= layer0_outputs(229);
    layer1_outputs(6911) <= (layer0_outputs(7994)) and (layer0_outputs(12357));
    layer1_outputs(6912) <= not((layer0_outputs(6992)) or (layer0_outputs(1110)));
    layer1_outputs(6913) <= not(layer0_outputs(7005)) or (layer0_outputs(12448));
    layer1_outputs(6914) <= (layer0_outputs(6891)) and (layer0_outputs(12639));
    layer1_outputs(6915) <= not((layer0_outputs(9326)) and (layer0_outputs(11936)));
    layer1_outputs(6916) <= (layer0_outputs(5977)) or (layer0_outputs(1395));
    layer1_outputs(6917) <= not((layer0_outputs(7332)) xor (layer0_outputs(8732)));
    layer1_outputs(6918) <= layer0_outputs(4686);
    layer1_outputs(6919) <= (layer0_outputs(10278)) and not (layer0_outputs(10950));
    layer1_outputs(6920) <= (layer0_outputs(1071)) and not (layer0_outputs(6980));
    layer1_outputs(6921) <= not(layer0_outputs(3990));
    layer1_outputs(6922) <= not((layer0_outputs(3177)) or (layer0_outputs(6787)));
    layer1_outputs(6923) <= layer0_outputs(8796);
    layer1_outputs(6924) <= layer0_outputs(10445);
    layer1_outputs(6925) <= not((layer0_outputs(8124)) and (layer0_outputs(7042)));
    layer1_outputs(6926) <= not(layer0_outputs(10248));
    layer1_outputs(6927) <= not(layer0_outputs(2671));
    layer1_outputs(6928) <= layer0_outputs(7770);
    layer1_outputs(6929) <= (layer0_outputs(1309)) xor (layer0_outputs(3086));
    layer1_outputs(6930) <= not((layer0_outputs(10056)) and (layer0_outputs(8151)));
    layer1_outputs(6931) <= not((layer0_outputs(11206)) xor (layer0_outputs(7505)));
    layer1_outputs(6932) <= not((layer0_outputs(12761)) and (layer0_outputs(8296)));
    layer1_outputs(6933) <= not((layer0_outputs(3940)) xor (layer0_outputs(1314)));
    layer1_outputs(6934) <= not(layer0_outputs(6897)) or (layer0_outputs(11227));
    layer1_outputs(6935) <= layer0_outputs(8951);
    layer1_outputs(6936) <= not(layer0_outputs(4775));
    layer1_outputs(6937) <= not(layer0_outputs(502));
    layer1_outputs(6938) <= '1';
    layer1_outputs(6939) <= layer0_outputs(1481);
    layer1_outputs(6940) <= not(layer0_outputs(1923)) or (layer0_outputs(8015));
    layer1_outputs(6941) <= (layer0_outputs(2132)) or (layer0_outputs(11414));
    layer1_outputs(6942) <= (layer0_outputs(2309)) xor (layer0_outputs(11307));
    layer1_outputs(6943) <= (layer0_outputs(8374)) and not (layer0_outputs(12178));
    layer1_outputs(6944) <= '1';
    layer1_outputs(6945) <= not(layer0_outputs(10978)) or (layer0_outputs(1138));
    layer1_outputs(6946) <= not(layer0_outputs(10467)) or (layer0_outputs(10272));
    layer1_outputs(6947) <= not(layer0_outputs(3766));
    layer1_outputs(6948) <= not((layer0_outputs(9782)) and (layer0_outputs(1151)));
    layer1_outputs(6949) <= not((layer0_outputs(7680)) and (layer0_outputs(7701)));
    layer1_outputs(6950) <= not(layer0_outputs(7633));
    layer1_outputs(6951) <= not((layer0_outputs(11303)) or (layer0_outputs(9190)));
    layer1_outputs(6952) <= (layer0_outputs(1643)) and not (layer0_outputs(1870));
    layer1_outputs(6953) <= not(layer0_outputs(12787));
    layer1_outputs(6954) <= (layer0_outputs(2620)) and not (layer0_outputs(5671));
    layer1_outputs(6955) <= layer0_outputs(4528);
    layer1_outputs(6956) <= not((layer0_outputs(4243)) and (layer0_outputs(2520)));
    layer1_outputs(6957) <= not(layer0_outputs(11302));
    layer1_outputs(6958) <= (layer0_outputs(3497)) and (layer0_outputs(11579));
    layer1_outputs(6959) <= (layer0_outputs(9218)) xor (layer0_outputs(2180));
    layer1_outputs(6960) <= (layer0_outputs(8102)) and not (layer0_outputs(11437));
    layer1_outputs(6961) <= (layer0_outputs(10057)) and (layer0_outputs(10265));
    layer1_outputs(6962) <= not((layer0_outputs(11832)) and (layer0_outputs(4013)));
    layer1_outputs(6963) <= '0';
    layer1_outputs(6964) <= '1';
    layer1_outputs(6965) <= (layer0_outputs(4858)) and (layer0_outputs(2002));
    layer1_outputs(6966) <= not(layer0_outputs(8883));
    layer1_outputs(6967) <= layer0_outputs(11644);
    layer1_outputs(6968) <= not(layer0_outputs(4834)) or (layer0_outputs(12770));
    layer1_outputs(6969) <= layer0_outputs(10071);
    layer1_outputs(6970) <= (layer0_outputs(12183)) and not (layer0_outputs(10274));
    layer1_outputs(6971) <= (layer0_outputs(6965)) xor (layer0_outputs(7099));
    layer1_outputs(6972) <= (layer0_outputs(4628)) xor (layer0_outputs(2426));
    layer1_outputs(6973) <= layer0_outputs(5631);
    layer1_outputs(6974) <= (layer0_outputs(4246)) or (layer0_outputs(396));
    layer1_outputs(6975) <= (layer0_outputs(7582)) and not (layer0_outputs(11995));
    layer1_outputs(6976) <= (layer0_outputs(12127)) xor (layer0_outputs(8657));
    layer1_outputs(6977) <= not((layer0_outputs(4875)) xor (layer0_outputs(9975)));
    layer1_outputs(6978) <= (layer0_outputs(10543)) and not (layer0_outputs(4045));
    layer1_outputs(6979) <= not(layer0_outputs(12578)) or (layer0_outputs(8686));
    layer1_outputs(6980) <= not(layer0_outputs(2248)) or (layer0_outputs(6014));
    layer1_outputs(6981) <= not(layer0_outputs(10363));
    layer1_outputs(6982) <= (layer0_outputs(11405)) and not (layer0_outputs(6586));
    layer1_outputs(6983) <= '0';
    layer1_outputs(6984) <= (layer0_outputs(1530)) xor (layer0_outputs(5577));
    layer1_outputs(6985) <= not((layer0_outputs(4835)) or (layer0_outputs(614)));
    layer1_outputs(6986) <= not(layer0_outputs(4157));
    layer1_outputs(6987) <= (layer0_outputs(10430)) and not (layer0_outputs(2179));
    layer1_outputs(6988) <= not((layer0_outputs(10113)) and (layer0_outputs(1892)));
    layer1_outputs(6989) <= not((layer0_outputs(9128)) or (layer0_outputs(3718)));
    layer1_outputs(6990) <= (layer0_outputs(11779)) and (layer0_outputs(5282));
    layer1_outputs(6991) <= (layer0_outputs(10317)) and not (layer0_outputs(3184));
    layer1_outputs(6992) <= (layer0_outputs(5420)) and not (layer0_outputs(11821));
    layer1_outputs(6993) <= (layer0_outputs(2201)) and not (layer0_outputs(10824));
    layer1_outputs(6994) <= (layer0_outputs(7439)) and not (layer0_outputs(9847));
    layer1_outputs(6995) <= not(layer0_outputs(10563));
    layer1_outputs(6996) <= (layer0_outputs(6593)) and not (layer0_outputs(10043));
    layer1_outputs(6997) <= (layer0_outputs(8112)) and (layer0_outputs(9018));
    layer1_outputs(6998) <= (layer0_outputs(12421)) xor (layer0_outputs(7151));
    layer1_outputs(6999) <= not(layer0_outputs(4566));
    layer1_outputs(7000) <= (layer0_outputs(5252)) and not (layer0_outputs(6884));
    layer1_outputs(7001) <= not((layer0_outputs(9643)) or (layer0_outputs(6925)));
    layer1_outputs(7002) <= not(layer0_outputs(7491));
    layer1_outputs(7003) <= not(layer0_outputs(11784));
    layer1_outputs(7004) <= not((layer0_outputs(8562)) and (layer0_outputs(10714)));
    layer1_outputs(7005) <= layer0_outputs(3619);
    layer1_outputs(7006) <= layer0_outputs(1897);
    layer1_outputs(7007) <= '0';
    layer1_outputs(7008) <= not(layer0_outputs(2815));
    layer1_outputs(7009) <= not(layer0_outputs(3969));
    layer1_outputs(7010) <= not((layer0_outputs(12586)) and (layer0_outputs(2150)));
    layer1_outputs(7011) <= not(layer0_outputs(2855));
    layer1_outputs(7012) <= (layer0_outputs(5743)) and not (layer0_outputs(11704));
    layer1_outputs(7013) <= (layer0_outputs(8807)) and (layer0_outputs(519));
    layer1_outputs(7014) <= (layer0_outputs(9076)) or (layer0_outputs(9143));
    layer1_outputs(7015) <= not(layer0_outputs(4133)) or (layer0_outputs(6976));
    layer1_outputs(7016) <= not(layer0_outputs(5166)) or (layer0_outputs(1288));
    layer1_outputs(7017) <= (layer0_outputs(3119)) or (layer0_outputs(3652));
    layer1_outputs(7018) <= not((layer0_outputs(6889)) xor (layer0_outputs(10709)));
    layer1_outputs(7019) <= layer0_outputs(6006);
    layer1_outputs(7020) <= layer0_outputs(6760);
    layer1_outputs(7021) <= not((layer0_outputs(5993)) or (layer0_outputs(11071)));
    layer1_outputs(7022) <= (layer0_outputs(11631)) and (layer0_outputs(9774));
    layer1_outputs(7023) <= (layer0_outputs(1240)) and not (layer0_outputs(5486));
    layer1_outputs(7024) <= not(layer0_outputs(2205));
    layer1_outputs(7025) <= not(layer0_outputs(7343));
    layer1_outputs(7026) <= not((layer0_outputs(11169)) and (layer0_outputs(11594)));
    layer1_outputs(7027) <= (layer0_outputs(4213)) and not (layer0_outputs(2689));
    layer1_outputs(7028) <= (layer0_outputs(498)) or (layer0_outputs(9257));
    layer1_outputs(7029) <= (layer0_outputs(10588)) and not (layer0_outputs(4603));
    layer1_outputs(7030) <= (layer0_outputs(11425)) and (layer0_outputs(1256));
    layer1_outputs(7031) <= not(layer0_outputs(12274));
    layer1_outputs(7032) <= not(layer0_outputs(2635));
    layer1_outputs(7033) <= layer0_outputs(5587);
    layer1_outputs(7034) <= not(layer0_outputs(6641));
    layer1_outputs(7035) <= '0';
    layer1_outputs(7036) <= not(layer0_outputs(2261)) or (layer0_outputs(1286));
    layer1_outputs(7037) <= layer0_outputs(12480);
    layer1_outputs(7038) <= (layer0_outputs(7924)) and not (layer0_outputs(1645));
    layer1_outputs(7039) <= not(layer0_outputs(2749)) or (layer0_outputs(10644));
    layer1_outputs(7040) <= (layer0_outputs(7252)) and not (layer0_outputs(10125));
    layer1_outputs(7041) <= not(layer0_outputs(11077));
    layer1_outputs(7042) <= (layer0_outputs(9355)) and not (layer0_outputs(787));
    layer1_outputs(7043) <= (layer0_outputs(12289)) and not (layer0_outputs(3788));
    layer1_outputs(7044) <= layer0_outputs(3117);
    layer1_outputs(7045) <= layer0_outputs(4064);
    layer1_outputs(7046) <= layer0_outputs(11845);
    layer1_outputs(7047) <= layer0_outputs(3074);
    layer1_outputs(7048) <= layer0_outputs(1790);
    layer1_outputs(7049) <= (layer0_outputs(6379)) and not (layer0_outputs(3849));
    layer1_outputs(7050) <= not(layer0_outputs(6798)) or (layer0_outputs(911));
    layer1_outputs(7051) <= not((layer0_outputs(7537)) or (layer0_outputs(8458)));
    layer1_outputs(7052) <= not(layer0_outputs(2235)) or (layer0_outputs(10987));
    layer1_outputs(7053) <= not(layer0_outputs(3055)) or (layer0_outputs(8075));
    layer1_outputs(7054) <= (layer0_outputs(1003)) and (layer0_outputs(3817));
    layer1_outputs(7055) <= not(layer0_outputs(2675)) or (layer0_outputs(10375));
    layer1_outputs(7056) <= '1';
    layer1_outputs(7057) <= (layer0_outputs(6112)) or (layer0_outputs(978));
    layer1_outputs(7058) <= not(layer0_outputs(4485));
    layer1_outputs(7059) <= layer0_outputs(8983);
    layer1_outputs(7060) <= (layer0_outputs(7949)) or (layer0_outputs(10564));
    layer1_outputs(7061) <= not(layer0_outputs(1803));
    layer1_outputs(7062) <= not(layer0_outputs(8329)) or (layer0_outputs(10852));
    layer1_outputs(7063) <= layer0_outputs(11026);
    layer1_outputs(7064) <= not((layer0_outputs(3321)) xor (layer0_outputs(1372)));
    layer1_outputs(7065) <= not(layer0_outputs(1631));
    layer1_outputs(7066) <= not(layer0_outputs(6553));
    layer1_outputs(7067) <= (layer0_outputs(3233)) and (layer0_outputs(1935));
    layer1_outputs(7068) <= not(layer0_outputs(7089));
    layer1_outputs(7069) <= not(layer0_outputs(4753));
    layer1_outputs(7070) <= (layer0_outputs(11235)) and (layer0_outputs(5385));
    layer1_outputs(7071) <= (layer0_outputs(10578)) and not (layer0_outputs(3296));
    layer1_outputs(7072) <= not(layer0_outputs(748));
    layer1_outputs(7073) <= not((layer0_outputs(8072)) xor (layer0_outputs(4607)));
    layer1_outputs(7074) <= not(layer0_outputs(7867)) or (layer0_outputs(4833));
    layer1_outputs(7075) <= layer0_outputs(4504);
    layer1_outputs(7076) <= (layer0_outputs(1158)) and not (layer0_outputs(2145));
    layer1_outputs(7077) <= layer0_outputs(6582);
    layer1_outputs(7078) <= not((layer0_outputs(6375)) xor (layer0_outputs(930)));
    layer1_outputs(7079) <= not((layer0_outputs(4959)) xor (layer0_outputs(6836)));
    layer1_outputs(7080) <= layer0_outputs(2193);
    layer1_outputs(7081) <= not(layer0_outputs(8936)) or (layer0_outputs(12697));
    layer1_outputs(7082) <= (layer0_outputs(6948)) and (layer0_outputs(8654));
    layer1_outputs(7083) <= not(layer0_outputs(5528)) or (layer0_outputs(9120));
    layer1_outputs(7084) <= layer0_outputs(8472);
    layer1_outputs(7085) <= (layer0_outputs(6873)) and not (layer0_outputs(11954));
    layer1_outputs(7086) <= layer0_outputs(6061);
    layer1_outputs(7087) <= not(layer0_outputs(7887));
    layer1_outputs(7088) <= '0';
    layer1_outputs(7089) <= not(layer0_outputs(3109));
    layer1_outputs(7090) <= (layer0_outputs(8579)) and not (layer0_outputs(8864));
    layer1_outputs(7091) <= not((layer0_outputs(5801)) and (layer0_outputs(7735)));
    layer1_outputs(7092) <= (layer0_outputs(2270)) and not (layer0_outputs(9085));
    layer1_outputs(7093) <= not(layer0_outputs(9175));
    layer1_outputs(7094) <= not((layer0_outputs(1874)) xor (layer0_outputs(107)));
    layer1_outputs(7095) <= not(layer0_outputs(5125)) or (layer0_outputs(7115));
    layer1_outputs(7096) <= layer0_outputs(9538);
    layer1_outputs(7097) <= not((layer0_outputs(1043)) and (layer0_outputs(10880)));
    layer1_outputs(7098) <= not((layer0_outputs(10727)) xor (layer0_outputs(1729)));
    layer1_outputs(7099) <= not(layer0_outputs(10842));
    layer1_outputs(7100) <= not(layer0_outputs(9751));
    layer1_outputs(7101) <= (layer0_outputs(5375)) and not (layer0_outputs(3406));
    layer1_outputs(7102) <= not((layer0_outputs(7434)) xor (layer0_outputs(507)));
    layer1_outputs(7103) <= not((layer0_outputs(12651)) xor (layer0_outputs(7239)));
    layer1_outputs(7104) <= '0';
    layer1_outputs(7105) <= (layer0_outputs(3486)) xor (layer0_outputs(10863));
    layer1_outputs(7106) <= (layer0_outputs(8830)) or (layer0_outputs(3401));
    layer1_outputs(7107) <= layer0_outputs(12357);
    layer1_outputs(7108) <= '1';
    layer1_outputs(7109) <= layer0_outputs(8068);
    layer1_outputs(7110) <= not(layer0_outputs(224));
    layer1_outputs(7111) <= not(layer0_outputs(1500)) or (layer0_outputs(8455));
    layer1_outputs(7112) <= (layer0_outputs(5222)) and not (layer0_outputs(10087));
    layer1_outputs(7113) <= layer0_outputs(6258);
    layer1_outputs(7114) <= not(layer0_outputs(5360));
    layer1_outputs(7115) <= not((layer0_outputs(8960)) or (layer0_outputs(11679)));
    layer1_outputs(7116) <= (layer0_outputs(5180)) and not (layer0_outputs(4769));
    layer1_outputs(7117) <= not(layer0_outputs(5111));
    layer1_outputs(7118) <= (layer0_outputs(5666)) and (layer0_outputs(12209));
    layer1_outputs(7119) <= layer0_outputs(10302);
    layer1_outputs(7120) <= (layer0_outputs(3030)) xor (layer0_outputs(3326));
    layer1_outputs(7121) <= not(layer0_outputs(12208));
    layer1_outputs(7122) <= not(layer0_outputs(6719));
    layer1_outputs(7123) <= not(layer0_outputs(1402));
    layer1_outputs(7124) <= layer0_outputs(5281);
    layer1_outputs(7125) <= not(layer0_outputs(4147));
    layer1_outputs(7126) <= not(layer0_outputs(11272)) or (layer0_outputs(4010));
    layer1_outputs(7127) <= layer0_outputs(1839);
    layer1_outputs(7128) <= not(layer0_outputs(1899));
    layer1_outputs(7129) <= layer0_outputs(27);
    layer1_outputs(7130) <= layer0_outputs(2431);
    layer1_outputs(7131) <= not(layer0_outputs(11381));
    layer1_outputs(7132) <= not(layer0_outputs(7984)) or (layer0_outputs(1654));
    layer1_outputs(7133) <= (layer0_outputs(812)) and (layer0_outputs(9030));
    layer1_outputs(7134) <= (layer0_outputs(11536)) and not (layer0_outputs(6987));
    layer1_outputs(7135) <= not(layer0_outputs(5090)) or (layer0_outputs(8242));
    layer1_outputs(7136) <= (layer0_outputs(6138)) xor (layer0_outputs(6236));
    layer1_outputs(7137) <= not(layer0_outputs(2685)) or (layer0_outputs(4089));
    layer1_outputs(7138) <= (layer0_outputs(9676)) and not (layer0_outputs(1660));
    layer1_outputs(7139) <= layer0_outputs(12573);
    layer1_outputs(7140) <= not((layer0_outputs(3158)) xor (layer0_outputs(12246)));
    layer1_outputs(7141) <= not(layer0_outputs(6999));
    layer1_outputs(7142) <= (layer0_outputs(11707)) and not (layer0_outputs(3957));
    layer1_outputs(7143) <= layer0_outputs(5955);
    layer1_outputs(7144) <= layer0_outputs(2162);
    layer1_outputs(7145) <= layer0_outputs(4793);
    layer1_outputs(7146) <= not((layer0_outputs(9112)) and (layer0_outputs(12613)));
    layer1_outputs(7147) <= not(layer0_outputs(8629));
    layer1_outputs(7148) <= (layer0_outputs(11415)) xor (layer0_outputs(9261));
    layer1_outputs(7149) <= (layer0_outputs(10088)) xor (layer0_outputs(12374));
    layer1_outputs(7150) <= not((layer0_outputs(7919)) or (layer0_outputs(6758)));
    layer1_outputs(7151) <= not(layer0_outputs(1396)) or (layer0_outputs(3844));
    layer1_outputs(7152) <= layer0_outputs(3374);
    layer1_outputs(7153) <= not((layer0_outputs(282)) and (layer0_outputs(12630)));
    layer1_outputs(7154) <= not(layer0_outputs(1083)) or (layer0_outputs(1994));
    layer1_outputs(7155) <= layer0_outputs(10183);
    layer1_outputs(7156) <= not(layer0_outputs(2987)) or (layer0_outputs(10644));
    layer1_outputs(7157) <= (layer0_outputs(1722)) and (layer0_outputs(7054));
    layer1_outputs(7158) <= not((layer0_outputs(1641)) or (layer0_outputs(4523)));
    layer1_outputs(7159) <= not(layer0_outputs(2708));
    layer1_outputs(7160) <= not(layer0_outputs(833));
    layer1_outputs(7161) <= layer0_outputs(6597);
    layer1_outputs(7162) <= not(layer0_outputs(12527)) or (layer0_outputs(12166));
    layer1_outputs(7163) <= (layer0_outputs(8705)) and not (layer0_outputs(8541));
    layer1_outputs(7164) <= (layer0_outputs(9364)) and not (layer0_outputs(5127));
    layer1_outputs(7165) <= not(layer0_outputs(7623)) or (layer0_outputs(8164));
    layer1_outputs(7166) <= layer0_outputs(9357);
    layer1_outputs(7167) <= not(layer0_outputs(12680));
    layer1_outputs(7168) <= not(layer0_outputs(3781));
    layer1_outputs(7169) <= (layer0_outputs(11496)) or (layer0_outputs(9622));
    layer1_outputs(7170) <= (layer0_outputs(7732)) and not (layer0_outputs(6875));
    layer1_outputs(7171) <= not(layer0_outputs(11752));
    layer1_outputs(7172) <= not(layer0_outputs(1405));
    layer1_outputs(7173) <= (layer0_outputs(9636)) xor (layer0_outputs(9096));
    layer1_outputs(7174) <= layer0_outputs(7622);
    layer1_outputs(7175) <= (layer0_outputs(7519)) xor (layer0_outputs(5009));
    layer1_outputs(7176) <= not((layer0_outputs(10740)) or (layer0_outputs(1736)));
    layer1_outputs(7177) <= (layer0_outputs(1745)) and not (layer0_outputs(6401));
    layer1_outputs(7178) <= '0';
    layer1_outputs(7179) <= not((layer0_outputs(8608)) xor (layer0_outputs(11936)));
    layer1_outputs(7180) <= (layer0_outputs(2324)) and (layer0_outputs(2547));
    layer1_outputs(7181) <= not(layer0_outputs(6079));
    layer1_outputs(7182) <= not(layer0_outputs(9872)) or (layer0_outputs(4110));
    layer1_outputs(7183) <= layer0_outputs(7730);
    layer1_outputs(7184) <= not(layer0_outputs(7509));
    layer1_outputs(7185) <= '0';
    layer1_outputs(7186) <= not(layer0_outputs(11826));
    layer1_outputs(7187) <= (layer0_outputs(3305)) xor (layer0_outputs(8756));
    layer1_outputs(7188) <= not(layer0_outputs(4478));
    layer1_outputs(7189) <= (layer0_outputs(7743)) or (layer0_outputs(3346));
    layer1_outputs(7190) <= (layer0_outputs(11817)) or (layer0_outputs(7529));
    layer1_outputs(7191) <= layer0_outputs(11115);
    layer1_outputs(7192) <= (layer0_outputs(2808)) and not (layer0_outputs(12605));
    layer1_outputs(7193) <= not((layer0_outputs(9944)) or (layer0_outputs(11935)));
    layer1_outputs(7194) <= not(layer0_outputs(10286)) or (layer0_outputs(163));
    layer1_outputs(7195) <= not((layer0_outputs(11400)) or (layer0_outputs(12266)));
    layer1_outputs(7196) <= not(layer0_outputs(10486)) or (layer0_outputs(5634));
    layer1_outputs(7197) <= not(layer0_outputs(1111));
    layer1_outputs(7198) <= layer0_outputs(1542);
    layer1_outputs(7199) <= layer0_outputs(3577);
    layer1_outputs(7200) <= (layer0_outputs(2909)) or (layer0_outputs(4087));
    layer1_outputs(7201) <= layer0_outputs(11832);
    layer1_outputs(7202) <= (layer0_outputs(12799)) and not (layer0_outputs(7299));
    layer1_outputs(7203) <= layer0_outputs(4204);
    layer1_outputs(7204) <= (layer0_outputs(3833)) and not (layer0_outputs(3919));
    layer1_outputs(7205) <= layer0_outputs(8222);
    layer1_outputs(7206) <= (layer0_outputs(3865)) and not (layer0_outputs(1144));
    layer1_outputs(7207) <= not((layer0_outputs(8228)) and (layer0_outputs(11455)));
    layer1_outputs(7208) <= layer0_outputs(1166);
    layer1_outputs(7209) <= (layer0_outputs(12112)) or (layer0_outputs(12221));
    layer1_outputs(7210) <= not((layer0_outputs(4902)) or (layer0_outputs(7094)));
    layer1_outputs(7211) <= (layer0_outputs(9567)) and not (layer0_outputs(10394));
    layer1_outputs(7212) <= not((layer0_outputs(8583)) or (layer0_outputs(10674)));
    layer1_outputs(7213) <= (layer0_outputs(3442)) or (layer0_outputs(11118));
    layer1_outputs(7214) <= not((layer0_outputs(10681)) and (layer0_outputs(4859)));
    layer1_outputs(7215) <= '1';
    layer1_outputs(7216) <= not((layer0_outputs(12643)) and (layer0_outputs(7771)));
    layer1_outputs(7217) <= not(layer0_outputs(11886));
    layer1_outputs(7218) <= (layer0_outputs(203)) and not (layer0_outputs(12438));
    layer1_outputs(7219) <= layer0_outputs(6152);
    layer1_outputs(7220) <= not((layer0_outputs(1401)) or (layer0_outputs(2761)));
    layer1_outputs(7221) <= (layer0_outputs(2832)) or (layer0_outputs(4592));
    layer1_outputs(7222) <= layer0_outputs(12102);
    layer1_outputs(7223) <= layer0_outputs(587);
    layer1_outputs(7224) <= not(layer0_outputs(5273));
    layer1_outputs(7225) <= layer0_outputs(4573);
    layer1_outputs(7226) <= layer0_outputs(5308);
    layer1_outputs(7227) <= not(layer0_outputs(8278)) or (layer0_outputs(5045));
    layer1_outputs(7228) <= (layer0_outputs(8703)) and not (layer0_outputs(4853));
    layer1_outputs(7229) <= not((layer0_outputs(3910)) or (layer0_outputs(3502)));
    layer1_outputs(7230) <= not(layer0_outputs(1100));
    layer1_outputs(7231) <= not(layer0_outputs(1777));
    layer1_outputs(7232) <= (layer0_outputs(5214)) and (layer0_outputs(3938));
    layer1_outputs(7233) <= (layer0_outputs(10929)) or (layer0_outputs(10449));
    layer1_outputs(7234) <= not(layer0_outputs(12683));
    layer1_outputs(7235) <= layer0_outputs(4431);
    layer1_outputs(7236) <= not(layer0_outputs(3400)) or (layer0_outputs(8319));
    layer1_outputs(7237) <= layer0_outputs(12742);
    layer1_outputs(7238) <= not((layer0_outputs(5833)) xor (layer0_outputs(12094)));
    layer1_outputs(7239) <= (layer0_outputs(9327)) or (layer0_outputs(4481));
    layer1_outputs(7240) <= not(layer0_outputs(2162)) or (layer0_outputs(8572));
    layer1_outputs(7241) <= (layer0_outputs(7956)) and not (layer0_outputs(5562));
    layer1_outputs(7242) <= (layer0_outputs(2512)) xor (layer0_outputs(4489));
    layer1_outputs(7243) <= layer0_outputs(4952);
    layer1_outputs(7244) <= layer0_outputs(11077);
    layer1_outputs(7245) <= not((layer0_outputs(9607)) or (layer0_outputs(8989)));
    layer1_outputs(7246) <= not(layer0_outputs(887));
    layer1_outputs(7247) <= layer0_outputs(5528);
    layer1_outputs(7248) <= '0';
    layer1_outputs(7249) <= not(layer0_outputs(11201)) or (layer0_outputs(4818));
    layer1_outputs(7250) <= (layer0_outputs(11864)) and (layer0_outputs(10135));
    layer1_outputs(7251) <= layer0_outputs(6301);
    layer1_outputs(7252) <= not(layer0_outputs(9614));
    layer1_outputs(7253) <= (layer0_outputs(10438)) xor (layer0_outputs(7404));
    layer1_outputs(7254) <= not((layer0_outputs(9291)) xor (layer0_outputs(5518)));
    layer1_outputs(7255) <= layer0_outputs(3822);
    layer1_outputs(7256) <= layer0_outputs(8856);
    layer1_outputs(7257) <= layer0_outputs(9802);
    layer1_outputs(7258) <= (layer0_outputs(10985)) and not (layer0_outputs(476));
    layer1_outputs(7259) <= (layer0_outputs(9100)) and not (layer0_outputs(9220));
    layer1_outputs(7260) <= not((layer0_outputs(1811)) and (layer0_outputs(12204)));
    layer1_outputs(7261) <= layer0_outputs(2586);
    layer1_outputs(7262) <= not(layer0_outputs(8820)) or (layer0_outputs(2154));
    layer1_outputs(7263) <= not(layer0_outputs(206));
    layer1_outputs(7264) <= (layer0_outputs(5211)) xor (layer0_outputs(433));
    layer1_outputs(7265) <= not(layer0_outputs(4527));
    layer1_outputs(7266) <= not((layer0_outputs(6800)) and (layer0_outputs(849)));
    layer1_outputs(7267) <= not(layer0_outputs(5215));
    layer1_outputs(7268) <= not((layer0_outputs(1274)) xor (layer0_outputs(3353)));
    layer1_outputs(7269) <= not((layer0_outputs(5378)) xor (layer0_outputs(7226)));
    layer1_outputs(7270) <= layer0_outputs(10701);
    layer1_outputs(7271) <= layer0_outputs(8404);
    layer1_outputs(7272) <= (layer0_outputs(9924)) or (layer0_outputs(11588));
    layer1_outputs(7273) <= not(layer0_outputs(965)) or (layer0_outputs(3455));
    layer1_outputs(7274) <= (layer0_outputs(11197)) and not (layer0_outputs(11037));
    layer1_outputs(7275) <= '1';
    layer1_outputs(7276) <= not(layer0_outputs(1514));
    layer1_outputs(7277) <= layer0_outputs(1526);
    layer1_outputs(7278) <= (layer0_outputs(7349)) xor (layer0_outputs(799));
    layer1_outputs(7279) <= (layer0_outputs(4569)) and not (layer0_outputs(4796));
    layer1_outputs(7280) <= not((layer0_outputs(1244)) xor (layer0_outputs(10782)));
    layer1_outputs(7281) <= (layer0_outputs(7008)) and not (layer0_outputs(5864));
    layer1_outputs(7282) <= not(layer0_outputs(11311));
    layer1_outputs(7283) <= not(layer0_outputs(891)) or (layer0_outputs(5735));
    layer1_outputs(7284) <= (layer0_outputs(9675)) and not (layer0_outputs(12455));
    layer1_outputs(7285) <= (layer0_outputs(6896)) and not (layer0_outputs(6775));
    layer1_outputs(7286) <= not((layer0_outputs(2952)) or (layer0_outputs(1576)));
    layer1_outputs(7287) <= '0';
    layer1_outputs(7288) <= (layer0_outputs(2208)) and (layer0_outputs(7973));
    layer1_outputs(7289) <= not((layer0_outputs(8094)) xor (layer0_outputs(11245)));
    layer1_outputs(7290) <= not(layer0_outputs(8342)) or (layer0_outputs(7697));
    layer1_outputs(7291) <= layer0_outputs(332);
    layer1_outputs(7292) <= layer0_outputs(9185);
    layer1_outputs(7293) <= not((layer0_outputs(3422)) or (layer0_outputs(6351)));
    layer1_outputs(7294) <= (layer0_outputs(7819)) xor (layer0_outputs(4410));
    layer1_outputs(7295) <= not((layer0_outputs(2603)) or (layer0_outputs(4060)));
    layer1_outputs(7296) <= layer0_outputs(12056);
    layer1_outputs(7297) <= not(layer0_outputs(10330));
    layer1_outputs(7298) <= not(layer0_outputs(10873)) or (layer0_outputs(11329));
    layer1_outputs(7299) <= not(layer0_outputs(4056));
    layer1_outputs(7300) <= layer0_outputs(11887);
    layer1_outputs(7301) <= (layer0_outputs(4886)) and (layer0_outputs(8007));
    layer1_outputs(7302) <= not(layer0_outputs(4526));
    layer1_outputs(7303) <= layer0_outputs(2659);
    layer1_outputs(7304) <= not(layer0_outputs(10894));
    layer1_outputs(7305) <= not(layer0_outputs(10590)) or (layer0_outputs(11249));
    layer1_outputs(7306) <= not((layer0_outputs(5909)) or (layer0_outputs(3078)));
    layer1_outputs(7307) <= (layer0_outputs(2349)) or (layer0_outputs(9373));
    layer1_outputs(7308) <= (layer0_outputs(8879)) and not (layer0_outputs(7899));
    layer1_outputs(7309) <= (layer0_outputs(5546)) or (layer0_outputs(7082));
    layer1_outputs(7310) <= not(layer0_outputs(4411));
    layer1_outputs(7311) <= (layer0_outputs(11398)) and not (layer0_outputs(3648));
    layer1_outputs(7312) <= (layer0_outputs(6382)) and not (layer0_outputs(6646));
    layer1_outputs(7313) <= not(layer0_outputs(11972));
    layer1_outputs(7314) <= '1';
    layer1_outputs(7315) <= (layer0_outputs(6087)) or (layer0_outputs(6171));
    layer1_outputs(7316) <= (layer0_outputs(12055)) or (layer0_outputs(12599));
    layer1_outputs(7317) <= layer0_outputs(7852);
    layer1_outputs(7318) <= not(layer0_outputs(7528));
    layer1_outputs(7319) <= layer0_outputs(864);
    layer1_outputs(7320) <= not((layer0_outputs(10194)) or (layer0_outputs(11700)));
    layer1_outputs(7321) <= not(layer0_outputs(12637));
    layer1_outputs(7322) <= not((layer0_outputs(11207)) and (layer0_outputs(7614)));
    layer1_outputs(7323) <= not(layer0_outputs(5563));
    layer1_outputs(7324) <= (layer0_outputs(3759)) and (layer0_outputs(6651));
    layer1_outputs(7325) <= not(layer0_outputs(6498)) or (layer0_outputs(8948));
    layer1_outputs(7326) <= layer0_outputs(7502);
    layer1_outputs(7327) <= not(layer0_outputs(10635));
    layer1_outputs(7328) <= (layer0_outputs(12550)) and not (layer0_outputs(12629));
    layer1_outputs(7329) <= not(layer0_outputs(9891)) or (layer0_outputs(10383));
    layer1_outputs(7330) <= (layer0_outputs(6224)) and not (layer0_outputs(5241));
    layer1_outputs(7331) <= not(layer0_outputs(1499));
    layer1_outputs(7332) <= (layer0_outputs(10221)) xor (layer0_outputs(1710));
    layer1_outputs(7333) <= not(layer0_outputs(1553)) or (layer0_outputs(2379));
    layer1_outputs(7334) <= (layer0_outputs(3225)) and not (layer0_outputs(5211));
    layer1_outputs(7335) <= layer0_outputs(2191);
    layer1_outputs(7336) <= not(layer0_outputs(8355)) or (layer0_outputs(5164));
    layer1_outputs(7337) <= (layer0_outputs(12741)) and not (layer0_outputs(9352));
    layer1_outputs(7338) <= not((layer0_outputs(7726)) xor (layer0_outputs(11113)));
    layer1_outputs(7339) <= (layer0_outputs(12287)) and not (layer0_outputs(7508));
    layer1_outputs(7340) <= not((layer0_outputs(3266)) or (layer0_outputs(252)));
    layer1_outputs(7341) <= (layer0_outputs(9303)) xor (layer0_outputs(7904));
    layer1_outputs(7342) <= not(layer0_outputs(2744)) or (layer0_outputs(4276));
    layer1_outputs(7343) <= not(layer0_outputs(776)) or (layer0_outputs(12653));
    layer1_outputs(7344) <= layer0_outputs(4417);
    layer1_outputs(7345) <= not(layer0_outputs(284)) or (layer0_outputs(2606));
    layer1_outputs(7346) <= not((layer0_outputs(8606)) or (layer0_outputs(334)));
    layer1_outputs(7347) <= layer0_outputs(11863);
    layer1_outputs(7348) <= (layer0_outputs(8634)) or (layer0_outputs(5));
    layer1_outputs(7349) <= (layer0_outputs(12536)) or (layer0_outputs(3583));
    layer1_outputs(7350) <= not(layer0_outputs(8084)) or (layer0_outputs(8387));
    layer1_outputs(7351) <= not(layer0_outputs(11290));
    layer1_outputs(7352) <= (layer0_outputs(5146)) and (layer0_outputs(12498));
    layer1_outputs(7353) <= not(layer0_outputs(2094)) or (layer0_outputs(7696));
    layer1_outputs(7354) <= (layer0_outputs(11856)) and not (layer0_outputs(6781));
    layer1_outputs(7355) <= not(layer0_outputs(12707));
    layer1_outputs(7356) <= not((layer0_outputs(4389)) xor (layer0_outputs(1292)));
    layer1_outputs(7357) <= not(layer0_outputs(633));
    layer1_outputs(7358) <= layer0_outputs(2293);
    layer1_outputs(7359) <= not(layer0_outputs(3405));
    layer1_outputs(7360) <= not(layer0_outputs(2118));
    layer1_outputs(7361) <= (layer0_outputs(1084)) and not (layer0_outputs(2044));
    layer1_outputs(7362) <= (layer0_outputs(2627)) and (layer0_outputs(2100));
    layer1_outputs(7363) <= (layer0_outputs(9526)) and (layer0_outputs(11915));
    layer1_outputs(7364) <= layer0_outputs(5171);
    layer1_outputs(7365) <= not(layer0_outputs(10913));
    layer1_outputs(7366) <= not((layer0_outputs(10243)) or (layer0_outputs(4082)));
    layer1_outputs(7367) <= (layer0_outputs(2492)) and (layer0_outputs(2627));
    layer1_outputs(7368) <= not((layer0_outputs(11433)) xor (layer0_outputs(3021)));
    layer1_outputs(7369) <= layer0_outputs(6422);
    layer1_outputs(7370) <= not((layer0_outputs(11688)) xor (layer0_outputs(7327)));
    layer1_outputs(7371) <= not(layer0_outputs(10503));
    layer1_outputs(7372) <= not((layer0_outputs(12597)) and (layer0_outputs(9435)));
    layer1_outputs(7373) <= not(layer0_outputs(10154)) or (layer0_outputs(4288));
    layer1_outputs(7374) <= (layer0_outputs(119)) and (layer0_outputs(3075));
    layer1_outputs(7375) <= layer0_outputs(3122);
    layer1_outputs(7376) <= not(layer0_outputs(1873)) or (layer0_outputs(3897));
    layer1_outputs(7377) <= not((layer0_outputs(10702)) xor (layer0_outputs(7492)));
    layer1_outputs(7378) <= not((layer0_outputs(3501)) or (layer0_outputs(2725)));
    layer1_outputs(7379) <= not((layer0_outputs(1858)) and (layer0_outputs(9331)));
    layer1_outputs(7380) <= layer0_outputs(3108);
    layer1_outputs(7381) <= (layer0_outputs(8650)) and (layer0_outputs(6460));
    layer1_outputs(7382) <= layer0_outputs(9424);
    layer1_outputs(7383) <= not((layer0_outputs(4828)) or (layer0_outputs(8508)));
    layer1_outputs(7384) <= layer0_outputs(12463);
    layer1_outputs(7385) <= not(layer0_outputs(9226)) or (layer0_outputs(7908));
    layer1_outputs(7386) <= layer0_outputs(6647);
    layer1_outputs(7387) <= layer0_outputs(5742);
    layer1_outputs(7388) <= not((layer0_outputs(10761)) and (layer0_outputs(7665)));
    layer1_outputs(7389) <= not(layer0_outputs(11636));
    layer1_outputs(7390) <= not((layer0_outputs(4980)) or (layer0_outputs(1952)));
    layer1_outputs(7391) <= not((layer0_outputs(5098)) or (layer0_outputs(2267)));
    layer1_outputs(7392) <= not(layer0_outputs(51));
    layer1_outputs(7393) <= layer0_outputs(1160);
    layer1_outputs(7394) <= not(layer0_outputs(1690)) or (layer0_outputs(3647));
    layer1_outputs(7395) <= (layer0_outputs(9144)) or (layer0_outputs(10360));
    layer1_outputs(7396) <= '0';
    layer1_outputs(7397) <= not((layer0_outputs(11932)) or (layer0_outputs(3970)));
    layer1_outputs(7398) <= layer0_outputs(1894);
    layer1_outputs(7399) <= (layer0_outputs(7612)) and (layer0_outputs(6468));
    layer1_outputs(7400) <= not(layer0_outputs(7728));
    layer1_outputs(7401) <= layer0_outputs(12304);
    layer1_outputs(7402) <= not(layer0_outputs(4156));
    layer1_outputs(7403) <= not((layer0_outputs(3618)) and (layer0_outputs(9526)));
    layer1_outputs(7404) <= (layer0_outputs(6722)) and not (layer0_outputs(2185));
    layer1_outputs(7405) <= not((layer0_outputs(5249)) and (layer0_outputs(5094)));
    layer1_outputs(7406) <= layer0_outputs(6957);
    layer1_outputs(7407) <= (layer0_outputs(12447)) and not (layer0_outputs(8012));
    layer1_outputs(7408) <= (layer0_outputs(7995)) xor (layer0_outputs(2104));
    layer1_outputs(7409) <= layer0_outputs(3875);
    layer1_outputs(7410) <= not(layer0_outputs(6675));
    layer1_outputs(7411) <= not(layer0_outputs(10484)) or (layer0_outputs(919));
    layer1_outputs(7412) <= not(layer0_outputs(5714));
    layer1_outputs(7413) <= not(layer0_outputs(12232));
    layer1_outputs(7414) <= (layer0_outputs(8385)) xor (layer0_outputs(5226));
    layer1_outputs(7415) <= not(layer0_outputs(11121));
    layer1_outputs(7416) <= layer0_outputs(12672);
    layer1_outputs(7417) <= not(layer0_outputs(1673)) or (layer0_outputs(10551));
    layer1_outputs(7418) <= not((layer0_outputs(3713)) and (layer0_outputs(10847)));
    layer1_outputs(7419) <= not(layer0_outputs(12200));
    layer1_outputs(7420) <= layer0_outputs(4710);
    layer1_outputs(7421) <= not((layer0_outputs(9972)) or (layer0_outputs(11183)));
    layer1_outputs(7422) <= layer0_outputs(464);
    layer1_outputs(7423) <= layer0_outputs(11740);
    layer1_outputs(7424) <= (layer0_outputs(1599)) and not (layer0_outputs(10419));
    layer1_outputs(7425) <= (layer0_outputs(1998)) or (layer0_outputs(6201));
    layer1_outputs(7426) <= not(layer0_outputs(846));
    layer1_outputs(7427) <= (layer0_outputs(11457)) and not (layer0_outputs(7188));
    layer1_outputs(7428) <= not(layer0_outputs(736)) or (layer0_outputs(9996));
    layer1_outputs(7429) <= not((layer0_outputs(2504)) and (layer0_outputs(8927)));
    layer1_outputs(7430) <= (layer0_outputs(10815)) and not (layer0_outputs(7388));
    layer1_outputs(7431) <= not(layer0_outputs(12177)) or (layer0_outputs(5357));
    layer1_outputs(7432) <= (layer0_outputs(1250)) and not (layer0_outputs(2280));
    layer1_outputs(7433) <= not((layer0_outputs(6494)) xor (layer0_outputs(1251)));
    layer1_outputs(7434) <= not(layer0_outputs(3306)) or (layer0_outputs(8677));
    layer1_outputs(7435) <= not(layer0_outputs(3433)) or (layer0_outputs(1339));
    layer1_outputs(7436) <= (layer0_outputs(12406)) xor (layer0_outputs(11216));
    layer1_outputs(7437) <= layer0_outputs(2086);
    layer1_outputs(7438) <= layer0_outputs(7523);
    layer1_outputs(7439) <= not(layer0_outputs(7964)) or (layer0_outputs(12235));
    layer1_outputs(7440) <= (layer0_outputs(3399)) and (layer0_outputs(11703));
    layer1_outputs(7441) <= (layer0_outputs(8192)) or (layer0_outputs(6697));
    layer1_outputs(7442) <= layer0_outputs(3322);
    layer1_outputs(7443) <= layer0_outputs(881);
    layer1_outputs(7444) <= (layer0_outputs(1442)) and not (layer0_outputs(4989));
    layer1_outputs(7445) <= not(layer0_outputs(12666)) or (layer0_outputs(12016));
    layer1_outputs(7446) <= (layer0_outputs(1527)) and (layer0_outputs(9692));
    layer1_outputs(7447) <= not((layer0_outputs(10803)) xor (layer0_outputs(3435)));
    layer1_outputs(7448) <= layer0_outputs(2487);
    layer1_outputs(7449) <= layer0_outputs(154);
    layer1_outputs(7450) <= layer0_outputs(2754);
    layer1_outputs(7451) <= not(layer0_outputs(452));
    layer1_outputs(7452) <= not((layer0_outputs(6187)) xor (layer0_outputs(2930)));
    layer1_outputs(7453) <= not(layer0_outputs(3477));
    layer1_outputs(7454) <= not(layer0_outputs(2534)) or (layer0_outputs(9339));
    layer1_outputs(7455) <= '1';
    layer1_outputs(7456) <= not(layer0_outputs(10266)) or (layer0_outputs(12028));
    layer1_outputs(7457) <= (layer0_outputs(1865)) xor (layer0_outputs(12308));
    layer1_outputs(7458) <= (layer0_outputs(3337)) and not (layer0_outputs(2334));
    layer1_outputs(7459) <= not((layer0_outputs(6124)) and (layer0_outputs(4152)));
    layer1_outputs(7460) <= not(layer0_outputs(1916)) or (layer0_outputs(5877));
    layer1_outputs(7461) <= not(layer0_outputs(2399)) or (layer0_outputs(2236));
    layer1_outputs(7462) <= (layer0_outputs(11568)) and (layer0_outputs(12397));
    layer1_outputs(7463) <= (layer0_outputs(9083)) xor (layer0_outputs(5167));
    layer1_outputs(7464) <= layer0_outputs(9388);
    layer1_outputs(7465) <= not(layer0_outputs(2822));
    layer1_outputs(7466) <= not(layer0_outputs(10773)) or (layer0_outputs(9906));
    layer1_outputs(7467) <= not(layer0_outputs(1880));
    layer1_outputs(7468) <= not(layer0_outputs(1147));
    layer1_outputs(7469) <= layer0_outputs(11861);
    layer1_outputs(7470) <= not(layer0_outputs(12544)) or (layer0_outputs(6557));
    layer1_outputs(7471) <= (layer0_outputs(10795)) and not (layer0_outputs(6373));
    layer1_outputs(7472) <= not((layer0_outputs(8898)) and (layer0_outputs(9140)));
    layer1_outputs(7473) <= (layer0_outputs(4109)) and not (layer0_outputs(1829));
    layer1_outputs(7474) <= not(layer0_outputs(2649)) or (layer0_outputs(11191));
    layer1_outputs(7475) <= not((layer0_outputs(10413)) xor (layer0_outputs(2174)));
    layer1_outputs(7476) <= (layer0_outputs(7034)) or (layer0_outputs(899));
    layer1_outputs(7477) <= not(layer0_outputs(3403));
    layer1_outputs(7478) <= (layer0_outputs(11855)) and not (layer0_outputs(2391));
    layer1_outputs(7479) <= (layer0_outputs(11927)) and (layer0_outputs(480));
    layer1_outputs(7480) <= '0';
    layer1_outputs(7481) <= (layer0_outputs(3550)) and (layer0_outputs(1613));
    layer1_outputs(7482) <= not((layer0_outputs(7184)) and (layer0_outputs(6170)));
    layer1_outputs(7483) <= '1';
    layer1_outputs(7484) <= (layer0_outputs(6991)) or (layer0_outputs(8324));
    layer1_outputs(7485) <= not((layer0_outputs(8503)) xor (layer0_outputs(2767)));
    layer1_outputs(7486) <= (layer0_outputs(10546)) and (layer0_outputs(12731));
    layer1_outputs(7487) <= layer0_outputs(5099);
    layer1_outputs(7488) <= (layer0_outputs(1322)) and (layer0_outputs(3398));
    layer1_outputs(7489) <= not((layer0_outputs(10044)) or (layer0_outputs(108)));
    layer1_outputs(7490) <= not(layer0_outputs(11085));
    layer1_outputs(7491) <= not(layer0_outputs(5276)) or (layer0_outputs(931));
    layer1_outputs(7492) <= (layer0_outputs(10318)) and not (layer0_outputs(6031));
    layer1_outputs(7493) <= not((layer0_outputs(315)) or (layer0_outputs(10735)));
    layer1_outputs(7494) <= not(layer0_outputs(5347)) or (layer0_outputs(3737));
    layer1_outputs(7495) <= not(layer0_outputs(5013));
    layer1_outputs(7496) <= layer0_outputs(406);
    layer1_outputs(7497) <= layer0_outputs(4732);
    layer1_outputs(7498) <= not((layer0_outputs(11790)) xor (layer0_outputs(5113)));
    layer1_outputs(7499) <= not(layer0_outputs(3578));
    layer1_outputs(7500) <= (layer0_outputs(5010)) or (layer0_outputs(3332));
    layer1_outputs(7501) <= layer0_outputs(9456);
    layer1_outputs(7502) <= not(layer0_outputs(4114));
    layer1_outputs(7503) <= (layer0_outputs(6737)) or (layer0_outputs(9230));
    layer1_outputs(7504) <= not(layer0_outputs(11950));
    layer1_outputs(7505) <= not(layer0_outputs(6588));
    layer1_outputs(7506) <= not((layer0_outputs(5517)) and (layer0_outputs(6758)));
    layer1_outputs(7507) <= (layer0_outputs(4766)) or (layer0_outputs(5575));
    layer1_outputs(7508) <= (layer0_outputs(9681)) or (layer0_outputs(10451));
    layer1_outputs(7509) <= not(layer0_outputs(12308)) or (layer0_outputs(4515));
    layer1_outputs(7510) <= (layer0_outputs(5009)) xor (layer0_outputs(1911));
    layer1_outputs(7511) <= (layer0_outputs(8064)) or (layer0_outputs(11108));
    layer1_outputs(7512) <= '1';
    layer1_outputs(7513) <= layer0_outputs(9800);
    layer1_outputs(7514) <= not(layer0_outputs(12197)) or (layer0_outputs(8500));
    layer1_outputs(7515) <= not(layer0_outputs(7737));
    layer1_outputs(7516) <= not(layer0_outputs(776));
    layer1_outputs(7517) <= '0';
    layer1_outputs(7518) <= layer0_outputs(7372);
    layer1_outputs(7519) <= not((layer0_outputs(12683)) and (layer0_outputs(11918)));
    layer1_outputs(7520) <= (layer0_outputs(3801)) or (layer0_outputs(11328));
    layer1_outputs(7521) <= not(layer0_outputs(12303));
    layer1_outputs(7522) <= not((layer0_outputs(4735)) xor (layer0_outputs(3879)));
    layer1_outputs(7523) <= not(layer0_outputs(4272));
    layer1_outputs(7524) <= '0';
    layer1_outputs(7525) <= not((layer0_outputs(3413)) xor (layer0_outputs(5871)));
    layer1_outputs(7526) <= (layer0_outputs(9554)) or (layer0_outputs(197));
    layer1_outputs(7527) <= layer0_outputs(12271);
    layer1_outputs(7528) <= (layer0_outputs(12260)) and not (layer0_outputs(11744));
    layer1_outputs(7529) <= not((layer0_outputs(4138)) xor (layer0_outputs(10833)));
    layer1_outputs(7530) <= not(layer0_outputs(9585)) or (layer0_outputs(192));
    layer1_outputs(7531) <= not((layer0_outputs(9693)) xor (layer0_outputs(7546)));
    layer1_outputs(7532) <= not(layer0_outputs(139));
    layer1_outputs(7533) <= (layer0_outputs(429)) and (layer0_outputs(6180));
    layer1_outputs(7534) <= layer0_outputs(5676);
    layer1_outputs(7535) <= (layer0_outputs(1481)) and (layer0_outputs(2447));
    layer1_outputs(7536) <= layer0_outputs(662);
    layer1_outputs(7537) <= not((layer0_outputs(7826)) and (layer0_outputs(7991)));
    layer1_outputs(7538) <= (layer0_outputs(5125)) or (layer0_outputs(7495));
    layer1_outputs(7539) <= (layer0_outputs(3579)) xor (layer0_outputs(7594));
    layer1_outputs(7540) <= (layer0_outputs(9186)) xor (layer0_outputs(3104));
    layer1_outputs(7541) <= (layer0_outputs(7312)) xor (layer0_outputs(12236));
    layer1_outputs(7542) <= layer0_outputs(7621);
    layer1_outputs(7543) <= not((layer0_outputs(12499)) xor (layer0_outputs(11728)));
    layer1_outputs(7544) <= not((layer0_outputs(2608)) or (layer0_outputs(3404)));
    layer1_outputs(7545) <= (layer0_outputs(2004)) and not (layer0_outputs(8073));
    layer1_outputs(7546) <= not((layer0_outputs(8678)) xor (layer0_outputs(8210)));
    layer1_outputs(7547) <= layer0_outputs(2549);
    layer1_outputs(7548) <= (layer0_outputs(5316)) or (layer0_outputs(12523));
    layer1_outputs(7549) <= not(layer0_outputs(8295));
    layer1_outputs(7550) <= not(layer0_outputs(7870));
    layer1_outputs(7551) <= not(layer0_outputs(9910));
    layer1_outputs(7552) <= layer0_outputs(2885);
    layer1_outputs(7553) <= (layer0_outputs(9302)) or (layer0_outputs(1478));
    layer1_outputs(7554) <= (layer0_outputs(7569)) and not (layer0_outputs(11993));
    layer1_outputs(7555) <= (layer0_outputs(6759)) and not (layer0_outputs(10373));
    layer1_outputs(7556) <= (layer0_outputs(4134)) and not (layer0_outputs(6743));
    layer1_outputs(7557) <= not((layer0_outputs(7414)) xor (layer0_outputs(11091)));
    layer1_outputs(7558) <= not(layer0_outputs(9976));
    layer1_outputs(7559) <= not(layer0_outputs(8846));
    layer1_outputs(7560) <= not(layer0_outputs(655));
    layer1_outputs(7561) <= (layer0_outputs(11286)) or (layer0_outputs(10267));
    layer1_outputs(7562) <= layer0_outputs(3223);
    layer1_outputs(7563) <= layer0_outputs(2462);
    layer1_outputs(7564) <= not(layer0_outputs(3264));
    layer1_outputs(7565) <= layer0_outputs(9909);
    layer1_outputs(7566) <= layer0_outputs(4238);
    layer1_outputs(7567) <= not(layer0_outputs(8100));
    layer1_outputs(7568) <= not(layer0_outputs(1368)) or (layer0_outputs(1500));
    layer1_outputs(7569) <= not(layer0_outputs(8699)) or (layer0_outputs(4655));
    layer1_outputs(7570) <= not(layer0_outputs(1807));
    layer1_outputs(7571) <= not(layer0_outputs(6295)) or (layer0_outputs(11124));
    layer1_outputs(7572) <= not(layer0_outputs(5230));
    layer1_outputs(7573) <= (layer0_outputs(1789)) and not (layer0_outputs(8567));
    layer1_outputs(7574) <= layer0_outputs(4634);
    layer1_outputs(7575) <= layer0_outputs(10760);
    layer1_outputs(7576) <= layer0_outputs(6802);
    layer1_outputs(7577) <= (layer0_outputs(2980)) xor (layer0_outputs(9718));
    layer1_outputs(7578) <= (layer0_outputs(11473)) xor (layer0_outputs(11034));
    layer1_outputs(7579) <= '1';
    layer1_outputs(7580) <= (layer0_outputs(11043)) xor (layer0_outputs(6038));
    layer1_outputs(7581) <= not(layer0_outputs(10361));
    layer1_outputs(7582) <= layer0_outputs(6073);
    layer1_outputs(7583) <= (layer0_outputs(12151)) and not (layer0_outputs(11331));
    layer1_outputs(7584) <= not(layer0_outputs(6092));
    layer1_outputs(7585) <= not(layer0_outputs(4836));
    layer1_outputs(7586) <= layer0_outputs(4991);
    layer1_outputs(7587) <= not(layer0_outputs(9989)) or (layer0_outputs(7693));
    layer1_outputs(7588) <= (layer0_outputs(3488)) xor (layer0_outputs(5597));
    layer1_outputs(7589) <= layer0_outputs(3724);
    layer1_outputs(7590) <= not(layer0_outputs(913));
    layer1_outputs(7591) <= not(layer0_outputs(552));
    layer1_outputs(7592) <= not(layer0_outputs(12123));
    layer1_outputs(7593) <= (layer0_outputs(10177)) and (layer0_outputs(8515));
    layer1_outputs(7594) <= not((layer0_outputs(3132)) and (layer0_outputs(1343)));
    layer1_outputs(7595) <= layer0_outputs(8995);
    layer1_outputs(7596) <= not((layer0_outputs(3517)) xor (layer0_outputs(6317)));
    layer1_outputs(7597) <= (layer0_outputs(2885)) and not (layer0_outputs(11526));
    layer1_outputs(7598) <= not(layer0_outputs(8469)) or (layer0_outputs(11102));
    layer1_outputs(7599) <= (layer0_outputs(7719)) xor (layer0_outputs(8310));
    layer1_outputs(7600) <= layer0_outputs(4574);
    layer1_outputs(7601) <= layer0_outputs(2806);
    layer1_outputs(7602) <= not(layer0_outputs(2664)) or (layer0_outputs(5480));
    layer1_outputs(7603) <= layer0_outputs(317);
    layer1_outputs(7604) <= layer0_outputs(6323);
    layer1_outputs(7605) <= not(layer0_outputs(11938));
    layer1_outputs(7606) <= layer0_outputs(6955);
    layer1_outputs(7607) <= (layer0_outputs(8335)) and (layer0_outputs(3057));
    layer1_outputs(7608) <= not(layer0_outputs(10713)) or (layer0_outputs(11341));
    layer1_outputs(7609) <= not((layer0_outputs(7054)) and (layer0_outputs(3843)));
    layer1_outputs(7610) <= not(layer0_outputs(6743));
    layer1_outputs(7611) <= (layer0_outputs(3084)) or (layer0_outputs(2678));
    layer1_outputs(7612) <= not((layer0_outputs(11898)) or (layer0_outputs(9940)));
    layer1_outputs(7613) <= layer0_outputs(4085);
    layer1_outputs(7614) <= (layer0_outputs(836)) and not (layer0_outputs(8180));
    layer1_outputs(7615) <= (layer0_outputs(7130)) and (layer0_outputs(5970));
    layer1_outputs(7616) <= (layer0_outputs(9210)) or (layer0_outputs(10445));
    layer1_outputs(7617) <= not(layer0_outputs(7594));
    layer1_outputs(7618) <= not((layer0_outputs(6067)) and (layer0_outputs(673)));
    layer1_outputs(7619) <= layer0_outputs(2825);
    layer1_outputs(7620) <= not(layer0_outputs(4633));
    layer1_outputs(7621) <= (layer0_outputs(12107)) and (layer0_outputs(7763));
    layer1_outputs(7622) <= not((layer0_outputs(4363)) xor (layer0_outputs(6108)));
    layer1_outputs(7623) <= layer0_outputs(9471);
    layer1_outputs(7624) <= (layer0_outputs(4038)) xor (layer0_outputs(10838));
    layer1_outputs(7625) <= (layer0_outputs(10622)) and (layer0_outputs(10781));
    layer1_outputs(7626) <= not((layer0_outputs(8947)) or (layer0_outputs(7479)));
    layer1_outputs(7627) <= (layer0_outputs(1828)) and not (layer0_outputs(7393));
    layer1_outputs(7628) <= layer0_outputs(11177);
    layer1_outputs(7629) <= not((layer0_outputs(3419)) and (layer0_outputs(4630)));
    layer1_outputs(7630) <= not(layer0_outputs(3070));
    layer1_outputs(7631) <= not(layer0_outputs(3654)) or (layer0_outputs(3071));
    layer1_outputs(7632) <= (layer0_outputs(4187)) and not (layer0_outputs(4004));
    layer1_outputs(7633) <= not((layer0_outputs(11671)) and (layer0_outputs(4562)));
    layer1_outputs(7634) <= not(layer0_outputs(10048));
    layer1_outputs(7635) <= not((layer0_outputs(2806)) xor (layer0_outputs(2328)));
    layer1_outputs(7636) <= (layer0_outputs(8205)) and not (layer0_outputs(3277));
    layer1_outputs(7637) <= (layer0_outputs(188)) or (layer0_outputs(4551));
    layer1_outputs(7638) <= not(layer0_outputs(307)) or (layer0_outputs(1763));
    layer1_outputs(7639) <= not(layer0_outputs(5620));
    layer1_outputs(7640) <= not((layer0_outputs(11775)) and (layer0_outputs(12146)));
    layer1_outputs(7641) <= not(layer0_outputs(7780)) or (layer0_outputs(7422));
    layer1_outputs(7642) <= not((layer0_outputs(5476)) or (layer0_outputs(8884)));
    layer1_outputs(7643) <= not(layer0_outputs(7724));
    layer1_outputs(7644) <= (layer0_outputs(3685)) or (layer0_outputs(12688));
    layer1_outputs(7645) <= (layer0_outputs(8194)) xor (layer0_outputs(1267));
    layer1_outputs(7646) <= layer0_outputs(6639);
    layer1_outputs(7647) <= (layer0_outputs(459)) xor (layer0_outputs(1227));
    layer1_outputs(7648) <= (layer0_outputs(9346)) and not (layer0_outputs(711));
    layer1_outputs(7649) <= (layer0_outputs(7607)) and not (layer0_outputs(10332));
    layer1_outputs(7650) <= layer0_outputs(7820);
    layer1_outputs(7651) <= not(layer0_outputs(914));
    layer1_outputs(7652) <= not((layer0_outputs(10962)) xor (layer0_outputs(11101)));
    layer1_outputs(7653) <= not(layer0_outputs(7397));
    layer1_outputs(7654) <= not((layer0_outputs(12129)) xor (layer0_outputs(7103)));
    layer1_outputs(7655) <= (layer0_outputs(9846)) xor (layer0_outputs(4831));
    layer1_outputs(7656) <= not((layer0_outputs(4072)) and (layer0_outputs(2960)));
    layer1_outputs(7657) <= not(layer0_outputs(11982));
    layer1_outputs(7658) <= '1';
    layer1_outputs(7659) <= layer0_outputs(10297);
    layer1_outputs(7660) <= not(layer0_outputs(4910));
    layer1_outputs(7661) <= (layer0_outputs(118)) xor (layer0_outputs(604));
    layer1_outputs(7662) <= not(layer0_outputs(310)) or (layer0_outputs(8743));
    layer1_outputs(7663) <= not(layer0_outputs(5275));
    layer1_outputs(7664) <= layer0_outputs(9185);
    layer1_outputs(7665) <= '0';
    layer1_outputs(7666) <= (layer0_outputs(9169)) and not (layer0_outputs(3291));
    layer1_outputs(7667) <= layer0_outputs(7599);
    layer1_outputs(7668) <= not(layer0_outputs(785));
    layer1_outputs(7669) <= (layer0_outputs(8332)) and not (layer0_outputs(9308));
    layer1_outputs(7670) <= (layer0_outputs(4716)) and (layer0_outputs(9785));
    layer1_outputs(7671) <= (layer0_outputs(10151)) and not (layer0_outputs(1168));
    layer1_outputs(7672) <= (layer0_outputs(12392)) xor (layer0_outputs(6012));
    layer1_outputs(7673) <= not((layer0_outputs(11647)) xor (layer0_outputs(1423)));
    layer1_outputs(7674) <= not(layer0_outputs(5818)) or (layer0_outputs(9442));
    layer1_outputs(7675) <= not(layer0_outputs(2925)) or (layer0_outputs(5758));
    layer1_outputs(7676) <= layer0_outputs(2102);
    layer1_outputs(7677) <= (layer0_outputs(9398)) and not (layer0_outputs(4415));
    layer1_outputs(7678) <= not(layer0_outputs(27));
    layer1_outputs(7679) <= layer0_outputs(3831);
    layer1_outputs(7680) <= (layer0_outputs(9011)) and not (layer0_outputs(2734));
    layer1_outputs(7681) <= not(layer0_outputs(9694)) or (layer0_outputs(5912));
    layer1_outputs(7682) <= not(layer0_outputs(7782)) or (layer0_outputs(7128));
    layer1_outputs(7683) <= not((layer0_outputs(12133)) or (layer0_outputs(739)));
    layer1_outputs(7684) <= (layer0_outputs(6120)) and not (layer0_outputs(9418));
    layer1_outputs(7685) <= not(layer0_outputs(803)) or (layer0_outputs(5600));
    layer1_outputs(7686) <= not((layer0_outputs(9182)) and (layer0_outputs(11695)));
    layer1_outputs(7687) <= (layer0_outputs(618)) and not (layer0_outputs(9297));
    layer1_outputs(7688) <= (layer0_outputs(11468)) and not (layer0_outputs(4247));
    layer1_outputs(7689) <= not(layer0_outputs(8600));
    layer1_outputs(7690) <= not((layer0_outputs(917)) and (layer0_outputs(7644)));
    layer1_outputs(7691) <= not(layer0_outputs(6735)) or (layer0_outputs(1650));
    layer1_outputs(7692) <= (layer0_outputs(5059)) or (layer0_outputs(10799));
    layer1_outputs(7693) <= (layer0_outputs(11934)) or (layer0_outputs(6568));
    layer1_outputs(7694) <= not(layer0_outputs(9818));
    layer1_outputs(7695) <= not(layer0_outputs(11630));
    layer1_outputs(7696) <= not(layer0_outputs(8593));
    layer1_outputs(7697) <= not(layer0_outputs(420));
    layer1_outputs(7698) <= not((layer0_outputs(4597)) or (layer0_outputs(5408)));
    layer1_outputs(7699) <= (layer0_outputs(5554)) or (layer0_outputs(762));
    layer1_outputs(7700) <= not(layer0_outputs(5571));
    layer1_outputs(7701) <= not((layer0_outputs(369)) xor (layer0_outputs(4880)));
    layer1_outputs(7702) <= not(layer0_outputs(10327));
    layer1_outputs(7703) <= (layer0_outputs(1930)) and not (layer0_outputs(5015));
    layer1_outputs(7704) <= not((layer0_outputs(5960)) or (layer0_outputs(3626)));
    layer1_outputs(7705) <= not((layer0_outputs(2887)) and (layer0_outputs(6039)));
    layer1_outputs(7706) <= (layer0_outputs(9466)) and not (layer0_outputs(3385));
    layer1_outputs(7707) <= not(layer0_outputs(11888)) or (layer0_outputs(10347));
    layer1_outputs(7708) <= '1';
    layer1_outputs(7709) <= (layer0_outputs(2708)) and (layer0_outputs(2078));
    layer1_outputs(7710) <= layer0_outputs(2418);
    layer1_outputs(7711) <= layer0_outputs(437);
    layer1_outputs(7712) <= not(layer0_outputs(2921));
    layer1_outputs(7713) <= not(layer0_outputs(2706));
    layer1_outputs(7714) <= (layer0_outputs(2388)) or (layer0_outputs(10984));
    layer1_outputs(7715) <= not(layer0_outputs(10166)) or (layer0_outputs(6186));
    layer1_outputs(7716) <= (layer0_outputs(11116)) and not (layer0_outputs(5010));
    layer1_outputs(7717) <= layer0_outputs(10240);
    layer1_outputs(7718) <= layer0_outputs(8687);
    layer1_outputs(7719) <= not(layer0_outputs(1883));
    layer1_outputs(7720) <= not((layer0_outputs(12789)) xor (layer0_outputs(10311)));
    layer1_outputs(7721) <= not((layer0_outputs(8633)) or (layer0_outputs(8703)));
    layer1_outputs(7722) <= not(layer0_outputs(3865)) or (layer0_outputs(9642));
    layer1_outputs(7723) <= not(layer0_outputs(9470)) or (layer0_outputs(8593));
    layer1_outputs(7724) <= '0';
    layer1_outputs(7725) <= not(layer0_outputs(7741)) or (layer0_outputs(6131));
    layer1_outputs(7726) <= (layer0_outputs(950)) and (layer0_outputs(12092));
    layer1_outputs(7727) <= not((layer0_outputs(1031)) or (layer0_outputs(3250)));
    layer1_outputs(7728) <= not(layer0_outputs(4092));
    layer1_outputs(7729) <= (layer0_outputs(5117)) and not (layer0_outputs(5529));
    layer1_outputs(7730) <= not(layer0_outputs(5689)) or (layer0_outputs(8194));
    layer1_outputs(7731) <= not((layer0_outputs(3354)) xor (layer0_outputs(2875)));
    layer1_outputs(7732) <= not(layer0_outputs(9537)) or (layer0_outputs(5080));
    layer1_outputs(7733) <= layer0_outputs(10430);
    layer1_outputs(7734) <= not(layer0_outputs(11231));
    layer1_outputs(7735) <= layer0_outputs(4122);
    layer1_outputs(7736) <= not(layer0_outputs(4488));
    layer1_outputs(7737) <= (layer0_outputs(3210)) and not (layer0_outputs(4688));
    layer1_outputs(7738) <= not(layer0_outputs(8801)) or (layer0_outputs(350));
    layer1_outputs(7739) <= not(layer0_outputs(6395)) or (layer0_outputs(6916));
    layer1_outputs(7740) <= layer0_outputs(4656);
    layer1_outputs(7741) <= not(layer0_outputs(10325)) or (layer0_outputs(546));
    layer1_outputs(7742) <= not(layer0_outputs(8286)) or (layer0_outputs(3729));
    layer1_outputs(7743) <= not((layer0_outputs(6995)) or (layer0_outputs(11379)));
    layer1_outputs(7744) <= (layer0_outputs(10628)) and (layer0_outputs(2485));
    layer1_outputs(7745) <= not((layer0_outputs(6167)) or (layer0_outputs(340)));
    layer1_outputs(7746) <= (layer0_outputs(488)) and not (layer0_outputs(6968));
    layer1_outputs(7747) <= '1';
    layer1_outputs(7748) <= not(layer0_outputs(7554));
    layer1_outputs(7749) <= layer0_outputs(8938);
    layer1_outputs(7750) <= not(layer0_outputs(10114));
    layer1_outputs(7751) <= (layer0_outputs(8664)) and (layer0_outputs(657));
    layer1_outputs(7752) <= not(layer0_outputs(2683));
    layer1_outputs(7753) <= not(layer0_outputs(2545));
    layer1_outputs(7754) <= not(layer0_outputs(782));
    layer1_outputs(7755) <= not(layer0_outputs(4711));
    layer1_outputs(7756) <= not((layer0_outputs(3864)) or (layer0_outputs(7365)));
    layer1_outputs(7757) <= (layer0_outputs(38)) and not (layer0_outputs(1814));
    layer1_outputs(7758) <= layer0_outputs(2584);
    layer1_outputs(7759) <= not((layer0_outputs(3540)) and (layer0_outputs(836)));
    layer1_outputs(7760) <= layer0_outputs(840);
    layer1_outputs(7761) <= '1';
    layer1_outputs(7762) <= (layer0_outputs(886)) and not (layer0_outputs(12382));
    layer1_outputs(7763) <= (layer0_outputs(7395)) and (layer0_outputs(12705));
    layer1_outputs(7764) <= not((layer0_outputs(7247)) and (layer0_outputs(2663)));
    layer1_outputs(7765) <= not((layer0_outputs(7539)) or (layer0_outputs(6432)));
    layer1_outputs(7766) <= (layer0_outputs(12467)) xor (layer0_outputs(2091));
    layer1_outputs(7767) <= not(layer0_outputs(8401)) or (layer0_outputs(1533));
    layer1_outputs(7768) <= not(layer0_outputs(11191));
    layer1_outputs(7769) <= (layer0_outputs(3131)) or (layer0_outputs(7639));
    layer1_outputs(7770) <= '1';
    layer1_outputs(7771) <= not(layer0_outputs(1136));
    layer1_outputs(7772) <= (layer0_outputs(1145)) and not (layer0_outputs(3133));
    layer1_outputs(7773) <= not((layer0_outputs(10938)) or (layer0_outputs(499)));
    layer1_outputs(7774) <= (layer0_outputs(7881)) or (layer0_outputs(12365));
    layer1_outputs(7775) <= layer0_outputs(1543);
    layer1_outputs(7776) <= not((layer0_outputs(358)) or (layer0_outputs(9750)));
    layer1_outputs(7777) <= (layer0_outputs(8659)) xor (layer0_outputs(7832));
    layer1_outputs(7778) <= not(layer0_outputs(7890));
    layer1_outputs(7779) <= layer0_outputs(12145);
    layer1_outputs(7780) <= not(layer0_outputs(6611));
    layer1_outputs(7781) <= (layer0_outputs(5395)) and (layer0_outputs(583));
    layer1_outputs(7782) <= (layer0_outputs(10375)) and not (layer0_outputs(6902));
    layer1_outputs(7783) <= not(layer0_outputs(3413)) or (layer0_outputs(6204));
    layer1_outputs(7784) <= not(layer0_outputs(7794));
    layer1_outputs(7785) <= layer0_outputs(6719);
    layer1_outputs(7786) <= not(layer0_outputs(10163)) or (layer0_outputs(9052));
    layer1_outputs(7787) <= (layer0_outputs(2933)) and (layer0_outputs(8358));
    layer1_outputs(7788) <= layer0_outputs(9778);
    layer1_outputs(7789) <= (layer0_outputs(4962)) xor (layer0_outputs(8277));
    layer1_outputs(7790) <= (layer0_outputs(5313)) and (layer0_outputs(5900));
    layer1_outputs(7791) <= not(layer0_outputs(7835)) or (layer0_outputs(1258));
    layer1_outputs(7792) <= not((layer0_outputs(9135)) xor (layer0_outputs(11012)));
    layer1_outputs(7793) <= (layer0_outputs(691)) and (layer0_outputs(6784));
    layer1_outputs(7794) <= not(layer0_outputs(3200));
    layer1_outputs(7795) <= not(layer0_outputs(6015)) or (layer0_outputs(3615));
    layer1_outputs(7796) <= not(layer0_outputs(3899));
    layer1_outputs(7797) <= not(layer0_outputs(9147));
    layer1_outputs(7798) <= layer0_outputs(12154);
    layer1_outputs(7799) <= not(layer0_outputs(10500));
    layer1_outputs(7800) <= not(layer0_outputs(6409));
    layer1_outputs(7801) <= (layer0_outputs(2568)) and not (layer0_outputs(5041));
    layer1_outputs(7802) <= layer0_outputs(11140);
    layer1_outputs(7803) <= (layer0_outputs(195)) and not (layer0_outputs(5481));
    layer1_outputs(7804) <= layer0_outputs(6848);
    layer1_outputs(7805) <= (layer0_outputs(6444)) and not (layer0_outputs(7235));
    layer1_outputs(7806) <= not(layer0_outputs(9367)) or (layer0_outputs(5571));
    layer1_outputs(7807) <= not(layer0_outputs(2537));
    layer1_outputs(7808) <= not(layer0_outputs(10673));
    layer1_outputs(7809) <= not(layer0_outputs(1568));
    layer1_outputs(7810) <= (layer0_outputs(84)) or (layer0_outputs(11867));
    layer1_outputs(7811) <= layer0_outputs(960);
    layer1_outputs(7812) <= not(layer0_outputs(3846)) or (layer0_outputs(10629));
    layer1_outputs(7813) <= layer0_outputs(8070);
    layer1_outputs(7814) <= layer0_outputs(11040);
    layer1_outputs(7815) <= not(layer0_outputs(9625));
    layer1_outputs(7816) <= layer0_outputs(12718);
    layer1_outputs(7817) <= not(layer0_outputs(7630));
    layer1_outputs(7818) <= (layer0_outputs(12351)) and not (layer0_outputs(1436));
    layer1_outputs(7819) <= not((layer0_outputs(12735)) and (layer0_outputs(5405)));
    layer1_outputs(7820) <= not(layer0_outputs(5238)) or (layer0_outputs(4492));
    layer1_outputs(7821) <= not(layer0_outputs(4327)) or (layer0_outputs(5400));
    layer1_outputs(7822) <= layer0_outputs(12118);
    layer1_outputs(7823) <= layer0_outputs(256);
    layer1_outputs(7824) <= layer0_outputs(11668);
    layer1_outputs(7825) <= (layer0_outputs(7653)) and not (layer0_outputs(8566));
    layer1_outputs(7826) <= (layer0_outputs(11015)) and not (layer0_outputs(1753));
    layer1_outputs(7827) <= not(layer0_outputs(6064));
    layer1_outputs(7828) <= not((layer0_outputs(6693)) and (layer0_outputs(10049)));
    layer1_outputs(7829) <= not(layer0_outputs(7244));
    layer1_outputs(7830) <= (layer0_outputs(6138)) and not (layer0_outputs(11258));
    layer1_outputs(7831) <= not(layer0_outputs(3509)) or (layer0_outputs(72));
    layer1_outputs(7832) <= layer0_outputs(10808);
    layer1_outputs(7833) <= not(layer0_outputs(10449));
    layer1_outputs(7834) <= not(layer0_outputs(10390));
    layer1_outputs(7835) <= not(layer0_outputs(7499));
    layer1_outputs(7836) <= layer0_outputs(10415);
    layer1_outputs(7837) <= (layer0_outputs(448)) xor (layer0_outputs(8602));
    layer1_outputs(7838) <= not(layer0_outputs(9170)) or (layer0_outputs(5248));
    layer1_outputs(7839) <= not(layer0_outputs(6382)) or (layer0_outputs(2552));
    layer1_outputs(7840) <= (layer0_outputs(3147)) and (layer0_outputs(2262));
    layer1_outputs(7841) <= layer0_outputs(8109);
    layer1_outputs(7842) <= not(layer0_outputs(9613)) or (layer0_outputs(2128));
    layer1_outputs(7843) <= not((layer0_outputs(7657)) xor (layer0_outputs(11055)));
    layer1_outputs(7844) <= not(layer0_outputs(2439));
    layer1_outputs(7845) <= not(layer0_outputs(5628));
    layer1_outputs(7846) <= not((layer0_outputs(8083)) or (layer0_outputs(7758)));
    layer1_outputs(7847) <= layer0_outputs(4754);
    layer1_outputs(7848) <= not(layer0_outputs(824));
    layer1_outputs(7849) <= layer0_outputs(7966);
    layer1_outputs(7850) <= '0';
    layer1_outputs(7851) <= not(layer0_outputs(2765));
    layer1_outputs(7852) <= not(layer0_outputs(5102));
    layer1_outputs(7853) <= (layer0_outputs(3644)) and not (layer0_outputs(1241));
    layer1_outputs(7854) <= not(layer0_outputs(12108)) or (layer0_outputs(4867));
    layer1_outputs(7855) <= not(layer0_outputs(12139));
    layer1_outputs(7856) <= not(layer0_outputs(1157));
    layer1_outputs(7857) <= not(layer0_outputs(1979));
    layer1_outputs(7858) <= not(layer0_outputs(6415));
    layer1_outputs(7859) <= layer0_outputs(11960);
    layer1_outputs(7860) <= not(layer0_outputs(2670));
    layer1_outputs(7861) <= '0';
    layer1_outputs(7862) <= not(layer0_outputs(2463));
    layer1_outputs(7863) <= layer0_outputs(11709);
    layer1_outputs(7864) <= not((layer0_outputs(8)) and (layer0_outputs(11953)));
    layer1_outputs(7865) <= not(layer0_outputs(11413));
    layer1_outputs(7866) <= (layer0_outputs(8568)) xor (layer0_outputs(6996));
    layer1_outputs(7867) <= not(layer0_outputs(150)) or (layer0_outputs(3863));
    layer1_outputs(7868) <= (layer0_outputs(5538)) and not (layer0_outputs(12734));
    layer1_outputs(7869) <= not(layer0_outputs(2570));
    layer1_outputs(7870) <= not(layer0_outputs(5608));
    layer1_outputs(7871) <= not((layer0_outputs(4158)) and (layer0_outputs(12454)));
    layer1_outputs(7872) <= not(layer0_outputs(811));
    layer1_outputs(7873) <= (layer0_outputs(2396)) or (layer0_outputs(8594));
    layer1_outputs(7874) <= not(layer0_outputs(944));
    layer1_outputs(7875) <= not(layer0_outputs(2413)) or (layer0_outputs(11554));
    layer1_outputs(7876) <= not(layer0_outputs(11852));
    layer1_outputs(7877) <= (layer0_outputs(4161)) xor (layer0_outputs(3284));
    layer1_outputs(7878) <= not((layer0_outputs(4308)) and (layer0_outputs(4145)));
    layer1_outputs(7879) <= layer0_outputs(3485);
    layer1_outputs(7880) <= not((layer0_outputs(227)) and (layer0_outputs(5242)));
    layer1_outputs(7881) <= not(layer0_outputs(10057)) or (layer0_outputs(1793));
    layer1_outputs(7882) <= (layer0_outputs(1833)) and (layer0_outputs(5565));
    layer1_outputs(7883) <= not((layer0_outputs(10014)) or (layer0_outputs(11919)));
    layer1_outputs(7884) <= (layer0_outputs(11611)) xor (layer0_outputs(11881));
    layer1_outputs(7885) <= layer0_outputs(10716);
    layer1_outputs(7886) <= layer0_outputs(549);
    layer1_outputs(7887) <= layer0_outputs(9351);
    layer1_outputs(7888) <= '0';
    layer1_outputs(7889) <= not((layer0_outputs(3156)) and (layer0_outputs(11551)));
    layer1_outputs(7890) <= (layer0_outputs(9463)) and (layer0_outputs(2022));
    layer1_outputs(7891) <= not(layer0_outputs(3059));
    layer1_outputs(7892) <= not((layer0_outputs(6922)) xor (layer0_outputs(12384)));
    layer1_outputs(7893) <= (layer0_outputs(10210)) and (layer0_outputs(11625));
    layer1_outputs(7894) <= not(layer0_outputs(1102)) or (layer0_outputs(671));
    layer1_outputs(7895) <= (layer0_outputs(172)) and not (layer0_outputs(6091));
    layer1_outputs(7896) <= not((layer0_outputs(5365)) and (layer0_outputs(7580)));
    layer1_outputs(7897) <= not((layer0_outputs(1506)) and (layer0_outputs(11136)));
    layer1_outputs(7898) <= (layer0_outputs(8261)) and not (layer0_outputs(2903));
    layer1_outputs(7899) <= '0';
    layer1_outputs(7900) <= (layer0_outputs(168)) or (layer0_outputs(10324));
    layer1_outputs(7901) <= '1';
    layer1_outputs(7902) <= (layer0_outputs(2728)) and (layer0_outputs(5300));
    layer1_outputs(7903) <= (layer0_outputs(5833)) and not (layer0_outputs(2780));
    layer1_outputs(7904) <= not(layer0_outputs(11608)) or (layer0_outputs(12314));
    layer1_outputs(7905) <= layer0_outputs(3239);
    layer1_outputs(7906) <= layer0_outputs(2472);
    layer1_outputs(7907) <= (layer0_outputs(1489)) or (layer0_outputs(12340));
    layer1_outputs(7908) <= (layer0_outputs(5949)) and not (layer0_outputs(2737));
    layer1_outputs(7909) <= not(layer0_outputs(10440));
    layer1_outputs(7910) <= not((layer0_outputs(10961)) and (layer0_outputs(4344)));
    layer1_outputs(7911) <= layer0_outputs(729);
    layer1_outputs(7912) <= not((layer0_outputs(6523)) or (layer0_outputs(8397)));
    layer1_outputs(7913) <= not((layer0_outputs(1955)) or (layer0_outputs(10917)));
    layer1_outputs(7914) <= (layer0_outputs(11981)) xor (layer0_outputs(2176));
    layer1_outputs(7915) <= not(layer0_outputs(9290));
    layer1_outputs(7916) <= (layer0_outputs(12347)) and not (layer0_outputs(1248));
    layer1_outputs(7917) <= layer0_outputs(10406);
    layer1_outputs(7918) <= layer0_outputs(11698);
    layer1_outputs(7919) <= '1';
    layer1_outputs(7920) <= layer0_outputs(7369);
    layer1_outputs(7921) <= (layer0_outputs(3189)) or (layer0_outputs(10322));
    layer1_outputs(7922) <= (layer0_outputs(3851)) and (layer0_outputs(1634));
    layer1_outputs(7923) <= (layer0_outputs(6347)) or (layer0_outputs(8671));
    layer1_outputs(7924) <= not(layer0_outputs(9385));
    layer1_outputs(7925) <= layer0_outputs(8876);
    layer1_outputs(7926) <= not(layer0_outputs(3599)) or (layer0_outputs(5770));
    layer1_outputs(7927) <= layer0_outputs(10703);
    layer1_outputs(7928) <= (layer0_outputs(5857)) xor (layer0_outputs(8195));
    layer1_outputs(7929) <= not((layer0_outputs(8912)) and (layer0_outputs(2984)));
    layer1_outputs(7930) <= layer0_outputs(9920);
    layer1_outputs(7931) <= not((layer0_outputs(9824)) xor (layer0_outputs(10092)));
    layer1_outputs(7932) <= not((layer0_outputs(10910)) or (layer0_outputs(1640)));
    layer1_outputs(7933) <= not(layer0_outputs(606));
    layer1_outputs(7934) <= not(layer0_outputs(2443)) or (layer0_outputs(1337));
    layer1_outputs(7935) <= not((layer0_outputs(4202)) or (layer0_outputs(11434)));
    layer1_outputs(7936) <= not(layer0_outputs(10384)) or (layer0_outputs(3951));
    layer1_outputs(7937) <= layer0_outputs(6489);
    layer1_outputs(7938) <= not(layer0_outputs(6821));
    layer1_outputs(7939) <= (layer0_outputs(11204)) xor (layer0_outputs(6626));
    layer1_outputs(7940) <= (layer0_outputs(11476)) or (layer0_outputs(816));
    layer1_outputs(7941) <= layer0_outputs(3353);
    layer1_outputs(7942) <= (layer0_outputs(10237)) or (layer0_outputs(11989));
    layer1_outputs(7943) <= layer0_outputs(9288);
    layer1_outputs(7944) <= not(layer0_outputs(11917)) or (layer0_outputs(4938));
    layer1_outputs(7945) <= not((layer0_outputs(5324)) or (layer0_outputs(12058)));
    layer1_outputs(7946) <= not(layer0_outputs(3895));
    layer1_outputs(7947) <= not(layer0_outputs(9285)) or (layer0_outputs(7766));
    layer1_outputs(7948) <= layer0_outputs(11679);
    layer1_outputs(7949) <= not((layer0_outputs(11992)) xor (layer0_outputs(3774)));
    layer1_outputs(7950) <= not(layer0_outputs(7681)) or (layer0_outputs(11904));
    layer1_outputs(7951) <= not(layer0_outputs(6930));
    layer1_outputs(7952) <= layer0_outputs(6106);
    layer1_outputs(7953) <= not((layer0_outputs(10100)) and (layer0_outputs(8383)));
    layer1_outputs(7954) <= not(layer0_outputs(5221)) or (layer0_outputs(1857));
    layer1_outputs(7955) <= (layer0_outputs(3047)) xor (layer0_outputs(12401));
    layer1_outputs(7956) <= layer0_outputs(12601);
    layer1_outputs(7957) <= layer0_outputs(6613);
    layer1_outputs(7958) <= not(layer0_outputs(5076));
    layer1_outputs(7959) <= layer0_outputs(5398);
    layer1_outputs(7960) <= not((layer0_outputs(5653)) xor (layer0_outputs(11050)));
    layer1_outputs(7961) <= layer0_outputs(863);
    layer1_outputs(7962) <= (layer0_outputs(8723)) xor (layer0_outputs(2127));
    layer1_outputs(7963) <= layer0_outputs(12656);
    layer1_outputs(7964) <= not(layer0_outputs(7065)) or (layer0_outputs(12025));
    layer1_outputs(7965) <= not((layer0_outputs(2564)) or (layer0_outputs(8424)));
    layer1_outputs(7966) <= layer0_outputs(5156);
    layer1_outputs(7967) <= not(layer0_outputs(8067));
    layer1_outputs(7968) <= (layer0_outputs(2533)) xor (layer0_outputs(11762));
    layer1_outputs(7969) <= (layer0_outputs(1747)) and (layer0_outputs(8877));
    layer1_outputs(7970) <= not((layer0_outputs(5902)) xor (layer0_outputs(7025)));
    layer1_outputs(7971) <= not((layer0_outputs(3562)) and (layer0_outputs(5383)));
    layer1_outputs(7972) <= (layer0_outputs(8950)) or (layer0_outputs(3716));
    layer1_outputs(7973) <= (layer0_outputs(7692)) and (layer0_outputs(12780));
    layer1_outputs(7974) <= not(layer0_outputs(2640)) or (layer0_outputs(7298));
    layer1_outputs(7975) <= not(layer0_outputs(7382));
    layer1_outputs(7976) <= not(layer0_outputs(10777));
    layer1_outputs(7977) <= layer0_outputs(9075);
    layer1_outputs(7978) <= not(layer0_outputs(1316));
    layer1_outputs(7979) <= not(layer0_outputs(9417)) or (layer0_outputs(7275));
    layer1_outputs(7980) <= (layer0_outputs(12084)) and (layer0_outputs(4294));
    layer1_outputs(7981) <= (layer0_outputs(6461)) xor (layer0_outputs(3290));
    layer1_outputs(7982) <= (layer0_outputs(1394)) xor (layer0_outputs(2790));
    layer1_outputs(7983) <= not(layer0_outputs(7892));
    layer1_outputs(7984) <= not(layer0_outputs(7117));
    layer1_outputs(7985) <= not(layer0_outputs(7791));
    layer1_outputs(7986) <= (layer0_outputs(9458)) and (layer0_outputs(2428));
    layer1_outputs(7987) <= not(layer0_outputs(8601)) or (layer0_outputs(9639));
    layer1_outputs(7988) <= layer0_outputs(10198);
    layer1_outputs(7989) <= '0';
    layer1_outputs(7990) <= (layer0_outputs(8180)) and not (layer0_outputs(12085));
    layer1_outputs(7991) <= layer0_outputs(3048);
    layer1_outputs(7992) <= not((layer0_outputs(1666)) or (layer0_outputs(2658)));
    layer1_outputs(7993) <= not(layer0_outputs(8762));
    layer1_outputs(7994) <= (layer0_outputs(250)) and (layer0_outputs(3998));
    layer1_outputs(7995) <= layer0_outputs(7480);
    layer1_outputs(7996) <= not(layer0_outputs(10139));
    layer1_outputs(7997) <= not(layer0_outputs(12600)) or (layer0_outputs(7165));
    layer1_outputs(7998) <= not(layer0_outputs(8689));
    layer1_outputs(7999) <= (layer0_outputs(7750)) xor (layer0_outputs(916));
    layer1_outputs(8000) <= not((layer0_outputs(478)) or (layer0_outputs(7637)));
    layer1_outputs(8001) <= layer0_outputs(2373);
    layer1_outputs(8002) <= (layer0_outputs(2215)) xor (layer0_outputs(2804));
    layer1_outputs(8003) <= (layer0_outputs(10633)) and not (layer0_outputs(11372));
    layer1_outputs(8004) <= layer0_outputs(6935);
    layer1_outputs(8005) <= layer0_outputs(10374);
    layer1_outputs(8006) <= layer0_outputs(11158);
    layer1_outputs(8007) <= (layer0_outputs(2032)) xor (layer0_outputs(7487));
    layer1_outputs(8008) <= layer0_outputs(9335);
    layer1_outputs(8009) <= (layer0_outputs(537)) and not (layer0_outputs(10703));
    layer1_outputs(8010) <= not(layer0_outputs(7746));
    layer1_outputs(8011) <= not(layer0_outputs(3448)) or (layer0_outputs(9815));
    layer1_outputs(8012) <= not((layer0_outputs(5723)) and (layer0_outputs(4695)));
    layer1_outputs(8013) <= (layer0_outputs(10041)) and not (layer0_outputs(1885));
    layer1_outputs(8014) <= not(layer0_outputs(7552));
    layer1_outputs(8015) <= not(layer0_outputs(10752)) or (layer0_outputs(6254));
    layer1_outputs(8016) <= not(layer0_outputs(3396));
    layer1_outputs(8017) <= layer0_outputs(7302);
    layer1_outputs(8018) <= not(layer0_outputs(9583));
    layer1_outputs(8019) <= not(layer0_outputs(2214));
    layer1_outputs(8020) <= layer0_outputs(7194);
    layer1_outputs(8021) <= (layer0_outputs(8538)) and not (layer0_outputs(7032));
    layer1_outputs(8022) <= not((layer0_outputs(12101)) xor (layer0_outputs(5386)));
    layer1_outputs(8023) <= (layer0_outputs(856)) and not (layer0_outputs(6313));
    layer1_outputs(8024) <= not(layer0_outputs(2515));
    layer1_outputs(8025) <= (layer0_outputs(7559)) and not (layer0_outputs(10434));
    layer1_outputs(8026) <= layer0_outputs(5812);
    layer1_outputs(8027) <= layer0_outputs(7625);
    layer1_outputs(8028) <= layer0_outputs(2405);
    layer1_outputs(8029) <= '1';
    layer1_outputs(8030) <= (layer0_outputs(4131)) and not (layer0_outputs(5754));
    layer1_outputs(8031) <= (layer0_outputs(1127)) and not (layer0_outputs(2632));
    layer1_outputs(8032) <= layer0_outputs(4248);
    layer1_outputs(8033) <= not(layer0_outputs(6289));
    layer1_outputs(8034) <= (layer0_outputs(568)) and (layer0_outputs(1065));
    layer1_outputs(8035) <= not((layer0_outputs(11332)) and (layer0_outputs(6387)));
    layer1_outputs(8036) <= not((layer0_outputs(11930)) and (layer0_outputs(1115)));
    layer1_outputs(8037) <= layer0_outputs(6506);
    layer1_outputs(8038) <= not((layer0_outputs(7587)) xor (layer0_outputs(1619)));
    layer1_outputs(8039) <= not(layer0_outputs(5478));
    layer1_outputs(8040) <= not(layer0_outputs(738)) or (layer0_outputs(1503));
    layer1_outputs(8041) <= layer0_outputs(2239);
    layer1_outputs(8042) <= (layer0_outputs(308)) and (layer0_outputs(11299));
    layer1_outputs(8043) <= not(layer0_outputs(9905));
    layer1_outputs(8044) <= (layer0_outputs(5284)) and not (layer0_outputs(1315));
    layer1_outputs(8045) <= layer0_outputs(4623);
    layer1_outputs(8046) <= not(layer0_outputs(1781)) or (layer0_outputs(2350));
    layer1_outputs(8047) <= not((layer0_outputs(6675)) or (layer0_outputs(12518)));
    layer1_outputs(8048) <= not(layer0_outputs(3649));
    layer1_outputs(8049) <= not((layer0_outputs(2500)) xor (layer0_outputs(10331)));
    layer1_outputs(8050) <= not((layer0_outputs(1907)) or (layer0_outputs(1905)));
    layer1_outputs(8051) <= (layer0_outputs(8571)) xor (layer0_outputs(1543));
    layer1_outputs(8052) <= '1';
    layer1_outputs(8053) <= not(layer0_outputs(12000));
    layer1_outputs(8054) <= layer0_outputs(7571);
    layer1_outputs(8055) <= not((layer0_outputs(6603)) and (layer0_outputs(7859)));
    layer1_outputs(8056) <= not((layer0_outputs(9639)) or (layer0_outputs(7490)));
    layer1_outputs(8057) <= not((layer0_outputs(8117)) and (layer0_outputs(8938)));
    layer1_outputs(8058) <= not((layer0_outputs(7655)) xor (layer0_outputs(3867)));
    layer1_outputs(8059) <= layer0_outputs(4840);
    layer1_outputs(8060) <= not((layer0_outputs(6842)) and (layer0_outputs(5882)));
    layer1_outputs(8061) <= (layer0_outputs(11897)) and (layer0_outputs(176));
    layer1_outputs(8062) <= not(layer0_outputs(3894));
    layer1_outputs(8063) <= (layer0_outputs(6687)) and (layer0_outputs(5260));
    layer1_outputs(8064) <= (layer0_outputs(10847)) and (layer0_outputs(4393));
    layer1_outputs(8065) <= layer0_outputs(624);
    layer1_outputs(8066) <= not(layer0_outputs(9571));
    layer1_outputs(8067) <= (layer0_outputs(11752)) or (layer0_outputs(10541));
    layer1_outputs(8068) <= not((layer0_outputs(1441)) xor (layer0_outputs(9505)));
    layer1_outputs(8069) <= not(layer0_outputs(10835)) or (layer0_outputs(11759));
    layer1_outputs(8070) <= layer0_outputs(8270);
    layer1_outputs(8071) <= (layer0_outputs(9009)) xor (layer0_outputs(538));
    layer1_outputs(8072) <= layer0_outputs(9807);
    layer1_outputs(8073) <= (layer0_outputs(123)) xor (layer0_outputs(4545));
    layer1_outputs(8074) <= (layer0_outputs(7354)) and (layer0_outputs(8753));
    layer1_outputs(8075) <= not(layer0_outputs(2618)) or (layer0_outputs(5788));
    layer1_outputs(8076) <= layer0_outputs(4595);
    layer1_outputs(8077) <= layer0_outputs(9419);
    layer1_outputs(8078) <= (layer0_outputs(6309)) and (layer0_outputs(10609));
    layer1_outputs(8079) <= not(layer0_outputs(10272));
    layer1_outputs(8080) <= not(layer0_outputs(1788)) or (layer0_outputs(3435));
    layer1_outputs(8081) <= not(layer0_outputs(9334)) or (layer0_outputs(5717));
    layer1_outputs(8082) <= not((layer0_outputs(440)) and (layer0_outputs(8991)));
    layer1_outputs(8083) <= (layer0_outputs(1154)) xor (layer0_outputs(2415));
    layer1_outputs(8084) <= layer0_outputs(5952);
    layer1_outputs(8085) <= not(layer0_outputs(956)) or (layer0_outputs(2702));
    layer1_outputs(8086) <= not((layer0_outputs(9600)) and (layer0_outputs(9945)));
    layer1_outputs(8087) <= not(layer0_outputs(1750)) or (layer0_outputs(6557));
    layer1_outputs(8088) <= not(layer0_outputs(7014)) or (layer0_outputs(10665));
    layer1_outputs(8089) <= layer0_outputs(3905);
    layer1_outputs(8090) <= not(layer0_outputs(11907));
    layer1_outputs(8091) <= layer0_outputs(10174);
    layer1_outputs(8092) <= (layer0_outputs(12682)) and (layer0_outputs(976));
    layer1_outputs(8093) <= (layer0_outputs(8867)) xor (layer0_outputs(844));
    layer1_outputs(8094) <= not((layer0_outputs(7352)) and (layer0_outputs(1887)));
    layer1_outputs(8095) <= not(layer0_outputs(6978));
    layer1_outputs(8096) <= layer0_outputs(8931);
    layer1_outputs(8097) <= not((layer0_outputs(10824)) or (layer0_outputs(11010)));
    layer1_outputs(8098) <= layer0_outputs(9318);
    layer1_outputs(8099) <= layer0_outputs(10139);
    layer1_outputs(8100) <= (layer0_outputs(8826)) and not (layer0_outputs(6145));
    layer1_outputs(8101) <= not((layer0_outputs(1112)) and (layer0_outputs(1984)));
    layer1_outputs(8102) <= not(layer0_outputs(5157)) or (layer0_outputs(700));
    layer1_outputs(8103) <= (layer0_outputs(1937)) and (layer0_outputs(5607));
    layer1_outputs(8104) <= layer0_outputs(5853);
    layer1_outputs(8105) <= (layer0_outputs(12440)) and (layer0_outputs(6004));
    layer1_outputs(8106) <= (layer0_outputs(3683)) and not (layer0_outputs(8357));
    layer1_outputs(8107) <= not(layer0_outputs(44));
    layer1_outputs(8108) <= not(layer0_outputs(9616));
    layer1_outputs(8109) <= (layer0_outputs(3694)) or (layer0_outputs(6869));
    layer1_outputs(8110) <= layer0_outputs(7583);
    layer1_outputs(8111) <= not((layer0_outputs(5195)) xor (layer0_outputs(4112)));
    layer1_outputs(8112) <= layer0_outputs(8990);
    layer1_outputs(8113) <= '1';
    layer1_outputs(8114) <= not(layer0_outputs(3067));
    layer1_outputs(8115) <= (layer0_outputs(9558)) and (layer0_outputs(1426));
    layer1_outputs(8116) <= not(layer0_outputs(12258)) or (layer0_outputs(8908));
    layer1_outputs(8117) <= not((layer0_outputs(1686)) or (layer0_outputs(10774)));
    layer1_outputs(8118) <= not((layer0_outputs(6160)) and (layer0_outputs(1840)));
    layer1_outputs(8119) <= not(layer0_outputs(4029));
    layer1_outputs(8120) <= (layer0_outputs(3573)) and (layer0_outputs(7935));
    layer1_outputs(8121) <= not(layer0_outputs(8433));
    layer1_outputs(8122) <= layer0_outputs(420);
    layer1_outputs(8123) <= not(layer0_outputs(9277));
    layer1_outputs(8124) <= layer0_outputs(5840);
    layer1_outputs(8125) <= (layer0_outputs(7958)) and not (layer0_outputs(3188));
    layer1_outputs(8126) <= layer0_outputs(4381);
    layer1_outputs(8127) <= not(layer0_outputs(3921));
    layer1_outputs(8128) <= not((layer0_outputs(6051)) xor (layer0_outputs(5499)));
    layer1_outputs(8129) <= not((layer0_outputs(2260)) and (layer0_outputs(241)));
    layer1_outputs(8130) <= not(layer0_outputs(4819)) or (layer0_outputs(10017));
    layer1_outputs(8131) <= not(layer0_outputs(5967));
    layer1_outputs(8132) <= layer0_outputs(6322);
    layer1_outputs(8133) <= not(layer0_outputs(4191));
    layer1_outputs(8134) <= (layer0_outputs(10193)) xor (layer0_outputs(3975));
    layer1_outputs(8135) <= layer0_outputs(1259);
    layer1_outputs(8136) <= not(layer0_outputs(7437));
    layer1_outputs(8137) <= (layer0_outputs(4790)) and not (layer0_outputs(3874));
    layer1_outputs(8138) <= not(layer0_outputs(5787));
    layer1_outputs(8139) <= layer0_outputs(920);
    layer1_outputs(8140) <= (layer0_outputs(10591)) or (layer0_outputs(8875));
    layer1_outputs(8141) <= layer0_outputs(11196);
    layer1_outputs(8142) <= not(layer0_outputs(11298));
    layer1_outputs(8143) <= layer0_outputs(1385);
    layer1_outputs(8144) <= not((layer0_outputs(5237)) and (layer0_outputs(11788)));
    layer1_outputs(8145) <= not(layer0_outputs(6576));
    layer1_outputs(8146) <= not(layer0_outputs(528));
    layer1_outputs(8147) <= not(layer0_outputs(7738));
    layer1_outputs(8148) <= layer0_outputs(12099);
    layer1_outputs(8149) <= not(layer0_outputs(3289));
    layer1_outputs(8150) <= layer0_outputs(9902);
    layer1_outputs(8151) <= not((layer0_outputs(31)) or (layer0_outputs(4077)));
    layer1_outputs(8152) <= layer0_outputs(9956);
    layer1_outputs(8153) <= not((layer0_outputs(3840)) xor (layer0_outputs(6745)));
    layer1_outputs(8154) <= (layer0_outputs(5320)) and not (layer0_outputs(10353));
    layer1_outputs(8155) <= layer0_outputs(127);
    layer1_outputs(8156) <= not((layer0_outputs(10305)) and (layer0_outputs(1818)));
    layer1_outputs(8157) <= not(layer0_outputs(1772)) or (layer0_outputs(4413));
    layer1_outputs(8158) <= layer0_outputs(9423);
    layer1_outputs(8159) <= not(layer0_outputs(12712));
    layer1_outputs(8160) <= not(layer0_outputs(697));
    layer1_outputs(8161) <= layer0_outputs(2340);
    layer1_outputs(8162) <= (layer0_outputs(1683)) and not (layer0_outputs(2762));
    layer1_outputs(8163) <= not(layer0_outputs(8717));
    layer1_outputs(8164) <= not(layer0_outputs(1008));
    layer1_outputs(8165) <= (layer0_outputs(6754)) or (layer0_outputs(4621));
    layer1_outputs(8166) <= '0';
    layer1_outputs(8167) <= (layer0_outputs(11922)) xor (layer0_outputs(4401));
    layer1_outputs(8168) <= (layer0_outputs(5674)) and (layer0_outputs(4805));
    layer1_outputs(8169) <= layer0_outputs(11990);
    layer1_outputs(8170) <= not(layer0_outputs(9163));
    layer1_outputs(8171) <= (layer0_outputs(3220)) and not (layer0_outputs(10403));
    layer1_outputs(8172) <= not(layer0_outputs(740));
    layer1_outputs(8173) <= (layer0_outputs(11956)) and (layer0_outputs(2704));
    layer1_outputs(8174) <= not((layer0_outputs(11326)) or (layer0_outputs(6799)));
    layer1_outputs(8175) <= layer0_outputs(4990);
    layer1_outputs(8176) <= not(layer0_outputs(167));
    layer1_outputs(8177) <= (layer0_outputs(2417)) and (layer0_outputs(6970));
    layer1_outputs(8178) <= (layer0_outputs(9249)) or (layer0_outputs(9029));
    layer1_outputs(8179) <= not((layer0_outputs(2322)) or (layer0_outputs(2553)));
    layer1_outputs(8180) <= not(layer0_outputs(1884)) or (layer0_outputs(5018));
    layer1_outputs(8181) <= (layer0_outputs(5632)) xor (layer0_outputs(2587));
    layer1_outputs(8182) <= '1';
    layer1_outputs(8183) <= (layer0_outputs(3396)) and not (layer0_outputs(7160));
    layer1_outputs(8184) <= not(layer0_outputs(2858));
    layer1_outputs(8185) <= not((layer0_outputs(7272)) or (layer0_outputs(12793)));
    layer1_outputs(8186) <= layer0_outputs(7698);
    layer1_outputs(8187) <= layer0_outputs(5185);
    layer1_outputs(8188) <= (layer0_outputs(326)) and not (layer0_outputs(9829));
    layer1_outputs(8189) <= not(layer0_outputs(3512));
    layer1_outputs(8190) <= layer0_outputs(8106);
    layer1_outputs(8191) <= not(layer0_outputs(21)) or (layer0_outputs(8839));
    layer1_outputs(8192) <= layer0_outputs(4349);
    layer1_outputs(8193) <= (layer0_outputs(7316)) xor (layer0_outputs(3021));
    layer1_outputs(8194) <= layer0_outputs(10785);
    layer1_outputs(8195) <= not(layer0_outputs(9453));
    layer1_outputs(8196) <= not(layer0_outputs(3320));
    layer1_outputs(8197) <= (layer0_outputs(6918)) and (layer0_outputs(4853));
    layer1_outputs(8198) <= not((layer0_outputs(6501)) xor (layer0_outputs(5208)));
    layer1_outputs(8199) <= not(layer0_outputs(2770));
    layer1_outputs(8200) <= (layer0_outputs(4410)) and not (layer0_outputs(7544));
    layer1_outputs(8201) <= '0';
    layer1_outputs(8202) <= (layer0_outputs(1273)) xor (layer0_outputs(1055));
    layer1_outputs(8203) <= layer0_outputs(3980);
    layer1_outputs(8204) <= layer0_outputs(906);
    layer1_outputs(8205) <= '0';
    layer1_outputs(8206) <= not(layer0_outputs(12130)) or (layer0_outputs(9281));
    layer1_outputs(8207) <= not(layer0_outputs(10321));
    layer1_outputs(8208) <= not(layer0_outputs(3847));
    layer1_outputs(8209) <= not((layer0_outputs(5304)) or (layer0_outputs(8676)));
    layer1_outputs(8210) <= not(layer0_outputs(405));
    layer1_outputs(8211) <= not(layer0_outputs(9464)) or (layer0_outputs(9947));
    layer1_outputs(8212) <= (layer0_outputs(3904)) and not (layer0_outputs(8705));
    layer1_outputs(8213) <= (layer0_outputs(11857)) and not (layer0_outputs(718));
    layer1_outputs(8214) <= not((layer0_outputs(2869)) and (layer0_outputs(7468)));
    layer1_outputs(8215) <= (layer0_outputs(1367)) or (layer0_outputs(2065));
    layer1_outputs(8216) <= not(layer0_outputs(10870));
    layer1_outputs(8217) <= not((layer0_outputs(11717)) or (layer0_outputs(6096)));
    layer1_outputs(8218) <= '0';
    layer1_outputs(8219) <= (layer0_outputs(10186)) and (layer0_outputs(6633));
    layer1_outputs(8220) <= not(layer0_outputs(9169));
    layer1_outputs(8221) <= layer0_outputs(2333);
    layer1_outputs(8222) <= not(layer0_outputs(1894));
    layer1_outputs(8223) <= not((layer0_outputs(2982)) xor (layer0_outputs(84)));
    layer1_outputs(8224) <= '0';
    layer1_outputs(8225) <= layer0_outputs(12611);
    layer1_outputs(8226) <= (layer0_outputs(10809)) or (layer0_outputs(4804));
    layer1_outputs(8227) <= not(layer0_outputs(4946)) or (layer0_outputs(12135));
    layer1_outputs(8228) <= not(layer0_outputs(10705));
    layer1_outputs(8229) <= not(layer0_outputs(6905));
    layer1_outputs(8230) <= not(layer0_outputs(12018));
    layer1_outputs(8231) <= (layer0_outputs(3490)) or (layer0_outputs(7249));
    layer1_outputs(8232) <= layer0_outputs(6359);
    layer1_outputs(8233) <= (layer0_outputs(8407)) and not (layer0_outputs(1677));
    layer1_outputs(8234) <= not(layer0_outputs(5270)) or (layer0_outputs(12048));
    layer1_outputs(8235) <= layer0_outputs(5070);
    layer1_outputs(8236) <= not(layer0_outputs(8544));
    layer1_outputs(8237) <= not((layer0_outputs(8110)) xor (layer0_outputs(10707)));
    layer1_outputs(8238) <= (layer0_outputs(4767)) and not (layer0_outputs(6284));
    layer1_outputs(8239) <= not((layer0_outputs(6018)) or (layer0_outputs(8440)));
    layer1_outputs(8240) <= not((layer0_outputs(3891)) xor (layer0_outputs(12109)));
    layer1_outputs(8241) <= layer0_outputs(1913);
    layer1_outputs(8242) <= layer0_outputs(9629);
    layer1_outputs(8243) <= '1';
    layer1_outputs(8244) <= not(layer0_outputs(7030)) or (layer0_outputs(3751));
    layer1_outputs(8245) <= not(layer0_outputs(10113));
    layer1_outputs(8246) <= layer0_outputs(6845);
    layer1_outputs(8247) <= layer0_outputs(11942);
    layer1_outputs(8248) <= not((layer0_outputs(5122)) xor (layer0_outputs(8794)));
    layer1_outputs(8249) <= layer0_outputs(9739);
    layer1_outputs(8250) <= layer0_outputs(8398);
    layer1_outputs(8251) <= (layer0_outputs(10730)) and (layer0_outputs(6808));
    layer1_outputs(8252) <= not(layer0_outputs(3681));
    layer1_outputs(8253) <= not(layer0_outputs(4526)) or (layer0_outputs(11333));
    layer1_outputs(8254) <= (layer0_outputs(5785)) and not (layer0_outputs(5327));
    layer1_outputs(8255) <= not((layer0_outputs(4647)) xor (layer0_outputs(5590)));
    layer1_outputs(8256) <= '1';
    layer1_outputs(8257) <= (layer0_outputs(7165)) and (layer0_outputs(11922));
    layer1_outputs(8258) <= not(layer0_outputs(9069));
    layer1_outputs(8259) <= not((layer0_outputs(11208)) or (layer0_outputs(11134)));
    layer1_outputs(8260) <= not((layer0_outputs(3004)) and (layer0_outputs(2996)));
    layer1_outputs(8261) <= not(layer0_outputs(8249)) or (layer0_outputs(3321));
    layer1_outputs(8262) <= layer0_outputs(11039);
    layer1_outputs(8263) <= not(layer0_outputs(3360)) or (layer0_outputs(3420));
    layer1_outputs(8264) <= not((layer0_outputs(8043)) and (layer0_outputs(755)));
    layer1_outputs(8265) <= not((layer0_outputs(4924)) or (layer0_outputs(6939)));
    layer1_outputs(8266) <= not((layer0_outputs(215)) xor (layer0_outputs(5083)));
    layer1_outputs(8267) <= not((layer0_outputs(113)) and (layer0_outputs(2482)));
    layer1_outputs(8268) <= (layer0_outputs(466)) xor (layer0_outputs(6993));
    layer1_outputs(8269) <= not((layer0_outputs(1313)) xor (layer0_outputs(6438)));
    layer1_outputs(8270) <= not(layer0_outputs(4359)) or (layer0_outputs(12293));
    layer1_outputs(8271) <= (layer0_outputs(8089)) and (layer0_outputs(7837));
    layer1_outputs(8272) <= not((layer0_outputs(12492)) xor (layer0_outputs(2279)));
    layer1_outputs(8273) <= not(layer0_outputs(7446)) or (layer0_outputs(1329));
    layer1_outputs(8274) <= not(layer0_outputs(9964)) or (layer0_outputs(10402));
    layer1_outputs(8275) <= not(layer0_outputs(7738));
    layer1_outputs(8276) <= not((layer0_outputs(4115)) or (layer0_outputs(11571)));
    layer1_outputs(8277) <= (layer0_outputs(9908)) and (layer0_outputs(4027));
    layer1_outputs(8278) <= '0';
    layer1_outputs(8279) <= layer0_outputs(6810);
    layer1_outputs(8280) <= (layer0_outputs(248)) and not (layer0_outputs(6360));
    layer1_outputs(8281) <= layer0_outputs(9197);
    layer1_outputs(8282) <= layer0_outputs(1385);
    layer1_outputs(8283) <= (layer0_outputs(7408)) and not (layer0_outputs(6892));
    layer1_outputs(8284) <= (layer0_outputs(2370)) xor (layer0_outputs(11482));
    layer1_outputs(8285) <= not(layer0_outputs(8895));
    layer1_outputs(8286) <= not(layer0_outputs(12334)) or (layer0_outputs(9438));
    layer1_outputs(8287) <= (layer0_outputs(11085)) and (layer0_outputs(7580));
    layer1_outputs(8288) <= (layer0_outputs(3594)) and (layer0_outputs(6264));
    layer1_outputs(8289) <= not(layer0_outputs(1792));
    layer1_outputs(8290) <= layer0_outputs(4754);
    layer1_outputs(8291) <= layer0_outputs(2604);
    layer1_outputs(8292) <= (layer0_outputs(2759)) and not (layer0_outputs(11215));
    layer1_outputs(8293) <= not((layer0_outputs(7974)) or (layer0_outputs(12)));
    layer1_outputs(8294) <= not(layer0_outputs(11747));
    layer1_outputs(8295) <= (layer0_outputs(8825)) xor (layer0_outputs(6255));
    layer1_outputs(8296) <= not(layer0_outputs(6057));
    layer1_outputs(8297) <= (layer0_outputs(7007)) and not (layer0_outputs(10508));
    layer1_outputs(8298) <= not(layer0_outputs(6029));
    layer1_outputs(8299) <= not(layer0_outputs(10256));
    layer1_outputs(8300) <= not(layer0_outputs(9492));
    layer1_outputs(8301) <= '1';
    layer1_outputs(8302) <= not((layer0_outputs(11305)) xor (layer0_outputs(7087)));
    layer1_outputs(8303) <= not(layer0_outputs(2600));
    layer1_outputs(8304) <= layer0_outputs(3661);
    layer1_outputs(8305) <= not((layer0_outputs(5372)) or (layer0_outputs(957)));
    layer1_outputs(8306) <= layer0_outputs(7879);
    layer1_outputs(8307) <= layer0_outputs(11370);
    layer1_outputs(8308) <= (layer0_outputs(7429)) and not (layer0_outputs(10422));
    layer1_outputs(8309) <= not(layer0_outputs(10993));
    layer1_outputs(8310) <= layer0_outputs(9792);
    layer1_outputs(8311) <= not(layer0_outputs(564));
    layer1_outputs(8312) <= not(layer0_outputs(64));
    layer1_outputs(8313) <= layer0_outputs(5458);
    layer1_outputs(8314) <= layer0_outputs(11359);
    layer1_outputs(8315) <= layer0_outputs(92);
    layer1_outputs(8316) <= (layer0_outputs(3993)) or (layer0_outputs(2186));
    layer1_outputs(8317) <= not(layer0_outputs(11194));
    layer1_outputs(8318) <= layer0_outputs(4839);
    layer1_outputs(8319) <= layer0_outputs(10466);
    layer1_outputs(8320) <= not(layer0_outputs(9035));
    layer1_outputs(8321) <= (layer0_outputs(8082)) xor (layer0_outputs(11157));
    layer1_outputs(8322) <= (layer0_outputs(5987)) or (layer0_outputs(740));
    layer1_outputs(8323) <= not(layer0_outputs(7649));
    layer1_outputs(8324) <= not(layer0_outputs(7930));
    layer1_outputs(8325) <= not(layer0_outputs(268));
    layer1_outputs(8326) <= not(layer0_outputs(2493));
    layer1_outputs(8327) <= not((layer0_outputs(1794)) xor (layer0_outputs(12261)));
    layer1_outputs(8328) <= (layer0_outputs(5182)) and not (layer0_outputs(9875));
    layer1_outputs(8329) <= not(layer0_outputs(10689)) or (layer0_outputs(11929));
    layer1_outputs(8330) <= not((layer0_outputs(1390)) or (layer0_outputs(4538)));
    layer1_outputs(8331) <= (layer0_outputs(7698)) and not (layer0_outputs(12037));
    layer1_outputs(8332) <= (layer0_outputs(6963)) and not (layer0_outputs(12074));
    layer1_outputs(8333) <= not(layer0_outputs(11988));
    layer1_outputs(8334) <= not(layer0_outputs(5068));
    layer1_outputs(8335) <= not(layer0_outputs(3437)) or (layer0_outputs(7443));
    layer1_outputs(8336) <= not(layer0_outputs(7027));
    layer1_outputs(8337) <= layer0_outputs(10221);
    layer1_outputs(8338) <= (layer0_outputs(5996)) and not (layer0_outputs(3668));
    layer1_outputs(8339) <= (layer0_outputs(7679)) or (layer0_outputs(11656));
    layer1_outputs(8340) <= (layer0_outputs(5716)) or (layer0_outputs(12777));
    layer1_outputs(8341) <= not(layer0_outputs(6761)) or (layer0_outputs(12377));
    layer1_outputs(8342) <= not((layer0_outputs(6095)) or (layer0_outputs(11219)));
    layer1_outputs(8343) <= (layer0_outputs(4843)) and not (layer0_outputs(494));
    layer1_outputs(8344) <= not(layer0_outputs(12644)) or (layer0_outputs(8403));
    layer1_outputs(8345) <= (layer0_outputs(11731)) and not (layer0_outputs(11623));
    layer1_outputs(8346) <= layer0_outputs(2666);
    layer1_outputs(8347) <= not((layer0_outputs(3890)) and (layer0_outputs(5212)));
    layer1_outputs(8348) <= not(layer0_outputs(1648)) or (layer0_outputs(9087));
    layer1_outputs(8349) <= not((layer0_outputs(5039)) xor (layer0_outputs(10884)));
    layer1_outputs(8350) <= not(layer0_outputs(427));
    layer1_outputs(8351) <= not(layer0_outputs(12168)) or (layer0_outputs(6895));
    layer1_outputs(8352) <= not(layer0_outputs(10380));
    layer1_outputs(8353) <= (layer0_outputs(9502)) and not (layer0_outputs(9724));
    layer1_outputs(8354) <= layer0_outputs(7226);
    layer1_outputs(8355) <= layer0_outputs(7491);
    layer1_outputs(8356) <= layer0_outputs(8851);
    layer1_outputs(8357) <= not(layer0_outputs(10683));
    layer1_outputs(8358) <= not((layer0_outputs(11214)) and (layer0_outputs(7167)));
    layer1_outputs(8359) <= (layer0_outputs(2147)) and not (layer0_outputs(12590));
    layer1_outputs(8360) <= (layer0_outputs(10403)) and (layer0_outputs(10514));
    layer1_outputs(8361) <= layer0_outputs(7691);
    layer1_outputs(8362) <= not(layer0_outputs(7709));
    layer1_outputs(8363) <= not(layer0_outputs(10773));
    layer1_outputs(8364) <= not(layer0_outputs(6519));
    layer1_outputs(8365) <= layer0_outputs(11190);
    layer1_outputs(8366) <= (layer0_outputs(10561)) and (layer0_outputs(452));
    layer1_outputs(8367) <= layer0_outputs(4332);
    layer1_outputs(8368) <= not(layer0_outputs(6176));
    layer1_outputs(8369) <= layer0_outputs(2257);
    layer1_outputs(8370) <= not(layer0_outputs(2238));
    layer1_outputs(8371) <= (layer0_outputs(10453)) and (layer0_outputs(1605));
    layer1_outputs(8372) <= not(layer0_outputs(6499));
    layer1_outputs(8373) <= not(layer0_outputs(6773)) or (layer0_outputs(7839));
    layer1_outputs(8374) <= not(layer0_outputs(7253));
    layer1_outputs(8375) <= not((layer0_outputs(4033)) and (layer0_outputs(6625)));
    layer1_outputs(8376) <= not(layer0_outputs(12129)) or (layer0_outputs(11525));
    layer1_outputs(8377) <= (layer0_outputs(8199)) and not (layer0_outputs(11678));
    layer1_outputs(8378) <= layer0_outputs(11167);
    layer1_outputs(8379) <= not((layer0_outputs(11765)) or (layer0_outputs(10959)));
    layer1_outputs(8380) <= not(layer0_outputs(4499));
    layer1_outputs(8381) <= not(layer0_outputs(3121)) or (layer0_outputs(5859));
    layer1_outputs(8382) <= (layer0_outputs(9021)) and not (layer0_outputs(2729));
    layer1_outputs(8383) <= not(layer0_outputs(7802)) or (layer0_outputs(6619));
    layer1_outputs(8384) <= not((layer0_outputs(10958)) xor (layer0_outputs(6032)));
    layer1_outputs(8385) <= layer0_outputs(12558);
    layer1_outputs(8386) <= layer0_outputs(7935);
    layer1_outputs(8387) <= (layer0_outputs(11031)) or (layer0_outputs(10074));
    layer1_outputs(8388) <= layer0_outputs(11022);
    layer1_outputs(8389) <= not(layer0_outputs(2599));
    layer1_outputs(8390) <= (layer0_outputs(6410)) and not (layer0_outputs(7832));
    layer1_outputs(8391) <= (layer0_outputs(9939)) and not (layer0_outputs(1859));
    layer1_outputs(8392) <= '0';
    layer1_outputs(8393) <= not((layer0_outputs(2509)) xor (layer0_outputs(8591)));
    layer1_outputs(8394) <= '1';
    layer1_outputs(8395) <= '0';
    layer1_outputs(8396) <= not((layer0_outputs(9567)) xor (layer0_outputs(10913)));
    layer1_outputs(8397) <= (layer0_outputs(963)) and not (layer0_outputs(1023));
    layer1_outputs(8398) <= not(layer0_outputs(8641));
    layer1_outputs(8399) <= layer0_outputs(7453);
    layer1_outputs(8400) <= not(layer0_outputs(1779));
    layer1_outputs(8401) <= not(layer0_outputs(10023)) or (layer0_outputs(1683));
    layer1_outputs(8402) <= not((layer0_outputs(10452)) and (layer0_outputs(5351)));
    layer1_outputs(8403) <= layer0_outputs(5460);
    layer1_outputs(8404) <= not(layer0_outputs(4388)) or (layer0_outputs(8612));
    layer1_outputs(8405) <= (layer0_outputs(3262)) and (layer0_outputs(2411));
    layer1_outputs(8406) <= (layer0_outputs(12317)) and not (layer0_outputs(2502));
    layer1_outputs(8407) <= layer0_outputs(12589);
    layer1_outputs(8408) <= layer0_outputs(9718);
    layer1_outputs(8409) <= (layer0_outputs(4896)) or (layer0_outputs(5038));
    layer1_outputs(8410) <= not((layer0_outputs(45)) and (layer0_outputs(8828)));
    layer1_outputs(8411) <= (layer0_outputs(9918)) and not (layer0_outputs(8642));
    layer1_outputs(8412) <= not((layer0_outputs(5380)) xor (layer0_outputs(1180)));
    layer1_outputs(8413) <= layer0_outputs(349);
    layer1_outputs(8414) <= layer0_outputs(12229);
    layer1_outputs(8415) <= (layer0_outputs(9667)) xor (layer0_outputs(9783));
    layer1_outputs(8416) <= not((layer0_outputs(6071)) and (layer0_outputs(1852)));
    layer1_outputs(8417) <= not(layer0_outputs(1130));
    layer1_outputs(8418) <= layer0_outputs(6840);
    layer1_outputs(8419) <= (layer0_outputs(3673)) and (layer0_outputs(7963));
    layer1_outputs(8420) <= (layer0_outputs(7356)) and (layer0_outputs(7940));
    layer1_outputs(8421) <= not(layer0_outputs(747)) or (layer0_outputs(5197));
    layer1_outputs(8422) <= (layer0_outputs(181)) and not (layer0_outputs(4429));
    layer1_outputs(8423) <= (layer0_outputs(1943)) xor (layer0_outputs(5655));
    layer1_outputs(8424) <= layer0_outputs(9147);
    layer1_outputs(8425) <= layer0_outputs(2753);
    layer1_outputs(8426) <= (layer0_outputs(602)) and not (layer0_outputs(5550));
    layer1_outputs(8427) <= not((layer0_outputs(6864)) xor (layer0_outputs(157)));
    layer1_outputs(8428) <= not((layer0_outputs(10174)) and (layer0_outputs(168)));
    layer1_outputs(8429) <= not((layer0_outputs(9312)) xor (layer0_outputs(11129)));
    layer1_outputs(8430) <= (layer0_outputs(3827)) or (layer0_outputs(8010));
    layer1_outputs(8431) <= (layer0_outputs(1146)) and not (layer0_outputs(10234));
    layer1_outputs(8432) <= not(layer0_outputs(9429));
    layer1_outputs(8433) <= (layer0_outputs(8582)) and (layer0_outputs(7039));
    layer1_outputs(8434) <= layer0_outputs(11790);
    layer1_outputs(8435) <= (layer0_outputs(1019)) and (layer0_outputs(12456));
    layer1_outputs(8436) <= not(layer0_outputs(7907));
    layer1_outputs(8437) <= layer0_outputs(6149);
    layer1_outputs(8438) <= (layer0_outputs(2938)) and (layer0_outputs(1359));
    layer1_outputs(8439) <= (layer0_outputs(10573)) or (layer0_outputs(10202));
    layer1_outputs(8440) <= not(layer0_outputs(645)) or (layer0_outputs(1010));
    layer1_outputs(8441) <= (layer0_outputs(3371)) and not (layer0_outputs(2603));
    layer1_outputs(8442) <= not(layer0_outputs(8366));
    layer1_outputs(8443) <= layer0_outputs(322);
    layer1_outputs(8444) <= layer0_outputs(10672);
    layer1_outputs(8445) <= not(layer0_outputs(12517));
    layer1_outputs(8446) <= not((layer0_outputs(7881)) or (layer0_outputs(8595)));
    layer1_outputs(8447) <= not(layer0_outputs(6868));
    layer1_outputs(8448) <= (layer0_outputs(591)) and (layer0_outputs(2028));
    layer1_outputs(8449) <= layer0_outputs(9231);
    layer1_outputs(8450) <= not(layer0_outputs(1488));
    layer1_outputs(8451) <= not((layer0_outputs(8432)) and (layer0_outputs(6059)));
    layer1_outputs(8452) <= (layer0_outputs(9674)) and not (layer0_outputs(9763));
    layer1_outputs(8453) <= (layer0_outputs(4931)) and (layer0_outputs(112));
    layer1_outputs(8454) <= layer0_outputs(4459);
    layer1_outputs(8455) <= (layer0_outputs(1415)) and (layer0_outputs(5906));
    layer1_outputs(8456) <= not(layer0_outputs(3955));
    layer1_outputs(8457) <= layer0_outputs(2042);
    layer1_outputs(8458) <= layer0_outputs(5361);
    layer1_outputs(8459) <= layer0_outputs(11200);
    layer1_outputs(8460) <= layer0_outputs(4625);
    layer1_outputs(8461) <= not((layer0_outputs(1365)) or (layer0_outputs(7310)));
    layer1_outputs(8462) <= (layer0_outputs(6656)) and not (layer0_outputs(11458));
    layer1_outputs(8463) <= (layer0_outputs(2380)) and (layer0_outputs(10290));
    layer1_outputs(8464) <= not((layer0_outputs(10156)) and (layer0_outputs(12457)));
    layer1_outputs(8465) <= layer0_outputs(10966);
    layer1_outputs(8466) <= layer0_outputs(5232);
    layer1_outputs(8467) <= not((layer0_outputs(9998)) xor (layer0_outputs(12662)));
    layer1_outputs(8468) <= (layer0_outputs(8457)) and (layer0_outputs(2907));
    layer1_outputs(8469) <= not(layer0_outputs(12388));
    layer1_outputs(8470) <= not((layer0_outputs(3433)) and (layer0_outputs(10992)));
    layer1_outputs(8471) <= not((layer0_outputs(11092)) and (layer0_outputs(7717)));
    layer1_outputs(8472) <= layer0_outputs(3814);
    layer1_outputs(8473) <= layer0_outputs(1574);
    layer1_outputs(8474) <= layer0_outputs(5848);
    layer1_outputs(8475) <= layer0_outputs(12531);
    layer1_outputs(8476) <= not(layer0_outputs(6362)) or (layer0_outputs(3461));
    layer1_outputs(8477) <= not((layer0_outputs(6986)) or (layer0_outputs(3671)));
    layer1_outputs(8478) <= (layer0_outputs(450)) and not (layer0_outputs(7507));
    layer1_outputs(8479) <= layer0_outputs(11361);
    layer1_outputs(8480) <= not(layer0_outputs(2287)) or (layer0_outputs(12017));
    layer1_outputs(8481) <= (layer0_outputs(2483)) or (layer0_outputs(2437));
    layer1_outputs(8482) <= not(layer0_outputs(11280)) or (layer0_outputs(5538));
    layer1_outputs(8483) <= not(layer0_outputs(7695));
    layer1_outputs(8484) <= not(layer0_outputs(2713)) or (layer0_outputs(8895));
    layer1_outputs(8485) <= not(layer0_outputs(990));
    layer1_outputs(8486) <= not(layer0_outputs(5153)) or (layer0_outputs(8241));
    layer1_outputs(8487) <= (layer0_outputs(12654)) xor (layer0_outputs(3805));
    layer1_outputs(8488) <= not((layer0_outputs(3861)) or (layer0_outputs(1294)));
    layer1_outputs(8489) <= (layer0_outputs(9104)) or (layer0_outputs(7197));
    layer1_outputs(8490) <= not((layer0_outputs(5704)) or (layer0_outputs(5077)));
    layer1_outputs(8491) <= layer0_outputs(4166);
    layer1_outputs(8492) <= not(layer0_outputs(7045));
    layer1_outputs(8493) <= (layer0_outputs(4324)) and not (layer0_outputs(2108));
    layer1_outputs(8494) <= layer0_outputs(5396);
    layer1_outputs(8495) <= layer0_outputs(8543);
    layer1_outputs(8496) <= not(layer0_outputs(2681));
    layer1_outputs(8497) <= not(layer0_outputs(7564));
    layer1_outputs(8498) <= not((layer0_outputs(1059)) and (layer0_outputs(4032)));
    layer1_outputs(8499) <= not(layer0_outputs(3139)) or (layer0_outputs(9610));
    layer1_outputs(8500) <= not((layer0_outputs(10313)) xor (layer0_outputs(11315)));
    layer1_outputs(8501) <= layer0_outputs(5441);
    layer1_outputs(8502) <= not(layer0_outputs(2087));
    layer1_outputs(8503) <= (layer0_outputs(8937)) xor (layer0_outputs(12485));
    layer1_outputs(8504) <= not(layer0_outputs(9667));
    layer1_outputs(8505) <= not(layer0_outputs(3625));
    layer1_outputs(8506) <= not(layer0_outputs(9726));
    layer1_outputs(8507) <= not(layer0_outputs(6326));
    layer1_outputs(8508) <= not(layer0_outputs(10545));
    layer1_outputs(8509) <= not(layer0_outputs(11648));
    layer1_outputs(8510) <= not((layer0_outputs(7729)) and (layer0_outputs(11045)));
    layer1_outputs(8511) <= layer0_outputs(3225);
    layer1_outputs(8512) <= not((layer0_outputs(1132)) and (layer0_outputs(2085)));
    layer1_outputs(8513) <= not(layer0_outputs(3854)) or (layer0_outputs(2384));
    layer1_outputs(8514) <= not((layer0_outputs(1074)) and (layer0_outputs(4213)));
    layer1_outputs(8515) <= not(layer0_outputs(5844));
    layer1_outputs(8516) <= not(layer0_outputs(8619));
    layer1_outputs(8517) <= not(layer0_outputs(11580));
    layer1_outputs(8518) <= (layer0_outputs(12426)) and not (layer0_outputs(8953));
    layer1_outputs(8519) <= not((layer0_outputs(10281)) and (layer0_outputs(6434)));
    layer1_outputs(8520) <= not((layer0_outputs(4914)) or (layer0_outputs(1680)));
    layer1_outputs(8521) <= not(layer0_outputs(6556));
    layer1_outputs(8522) <= (layer0_outputs(10026)) or (layer0_outputs(1133));
    layer1_outputs(8523) <= (layer0_outputs(2687)) and not (layer0_outputs(7785));
    layer1_outputs(8524) <= not((layer0_outputs(2129)) or (layer0_outputs(7591)));
    layer1_outputs(8525) <= (layer0_outputs(12521)) or (layer0_outputs(6376));
    layer1_outputs(8526) <= layer0_outputs(7426);
    layer1_outputs(8527) <= (layer0_outputs(7531)) xor (layer0_outputs(11313));
    layer1_outputs(8528) <= (layer0_outputs(8431)) and not (layer0_outputs(10024));
    layer1_outputs(8529) <= (layer0_outputs(319)) and not (layer0_outputs(351));
    layer1_outputs(8530) <= (layer0_outputs(9328)) and not (layer0_outputs(2561));
    layer1_outputs(8531) <= not((layer0_outputs(6061)) and (layer0_outputs(6853)));
    layer1_outputs(8532) <= layer0_outputs(8185);
    layer1_outputs(8533) <= (layer0_outputs(11373)) and not (layer0_outputs(1723));
    layer1_outputs(8534) <= not(layer0_outputs(12665));
    layer1_outputs(8535) <= layer0_outputs(12026);
    layer1_outputs(8536) <= not(layer0_outputs(7369));
    layer1_outputs(8537) <= not(layer0_outputs(6413)) or (layer0_outputs(9300));
    layer1_outputs(8538) <= not((layer0_outputs(9386)) xor (layer0_outputs(8932)));
    layer1_outputs(8539) <= layer0_outputs(4968);
    layer1_outputs(8540) <= not(layer0_outputs(9111));
    layer1_outputs(8541) <= not((layer0_outputs(4538)) xor (layer0_outputs(750)));
    layer1_outputs(8542) <= layer0_outputs(9524);
    layer1_outputs(8543) <= layer0_outputs(7876);
    layer1_outputs(8544) <= not(layer0_outputs(2189));
    layer1_outputs(8545) <= layer0_outputs(2084);
    layer1_outputs(8546) <= layer0_outputs(3358);
    layer1_outputs(8547) <= not(layer0_outputs(2984));
    layer1_outputs(8548) <= (layer0_outputs(3750)) and not (layer0_outputs(12359));
    layer1_outputs(8549) <= not(layer0_outputs(1536));
    layer1_outputs(8550) <= (layer0_outputs(7870)) and not (layer0_outputs(129));
    layer1_outputs(8551) <= not((layer0_outputs(11620)) or (layer0_outputs(8273)));
    layer1_outputs(8552) <= not(layer0_outputs(1148));
    layer1_outputs(8553) <= not(layer0_outputs(4085)) or (layer0_outputs(7787));
    layer1_outputs(8554) <= not((layer0_outputs(8126)) and (layer0_outputs(10302)));
    layer1_outputs(8555) <= layer0_outputs(7634);
    layer1_outputs(8556) <= not((layer0_outputs(5894)) xor (layer0_outputs(10549)));
    layer1_outputs(8557) <= (layer0_outputs(6068)) and not (layer0_outputs(4433));
    layer1_outputs(8558) <= not(layer0_outputs(1167));
    layer1_outputs(8559) <= (layer0_outputs(6632)) xor (layer0_outputs(10488));
    layer1_outputs(8560) <= (layer0_outputs(6485)) and (layer0_outputs(463));
    layer1_outputs(8561) <= not(layer0_outputs(8345));
    layer1_outputs(8562) <= (layer0_outputs(12248)) and not (layer0_outputs(4696));
    layer1_outputs(8563) <= not(layer0_outputs(10504));
    layer1_outputs(8564) <= not((layer0_outputs(4794)) and (layer0_outputs(9008)));
    layer1_outputs(8565) <= layer0_outputs(2347);
    layer1_outputs(8566) <= layer0_outputs(10520);
    layer1_outputs(8567) <= not(layer0_outputs(6166)) or (layer0_outputs(1357));
    layer1_outputs(8568) <= not(layer0_outputs(8229));
    layer1_outputs(8569) <= not(layer0_outputs(9213)) or (layer0_outputs(2889));
    layer1_outputs(8570) <= not(layer0_outputs(2199));
    layer1_outputs(8571) <= not((layer0_outputs(9994)) and (layer0_outputs(8291)));
    layer1_outputs(8572) <= not(layer0_outputs(2452));
    layer1_outputs(8573) <= not(layer0_outputs(11156));
    layer1_outputs(8574) <= not(layer0_outputs(11365)) or (layer0_outputs(175));
    layer1_outputs(8575) <= layer0_outputs(11817);
    layer1_outputs(8576) <= layer0_outputs(9926);
    layer1_outputs(8577) <= not(layer0_outputs(7503));
    layer1_outputs(8578) <= not((layer0_outputs(1601)) or (layer0_outputs(286)));
    layer1_outputs(8579) <= (layer0_outputs(2259)) or (layer0_outputs(12010));
    layer1_outputs(8580) <= layer0_outputs(1252);
    layer1_outputs(8581) <= layer0_outputs(6838);
    layer1_outputs(8582) <= (layer0_outputs(12323)) xor (layer0_outputs(339));
    layer1_outputs(8583) <= not(layer0_outputs(638));
    layer1_outputs(8584) <= (layer0_outputs(8218)) and (layer0_outputs(1598));
    layer1_outputs(8585) <= not((layer0_outputs(7262)) and (layer0_outputs(7164)));
    layer1_outputs(8586) <= layer0_outputs(1816);
    layer1_outputs(8587) <= not(layer0_outputs(2943)) or (layer0_outputs(4001));
    layer1_outputs(8588) <= (layer0_outputs(7002)) and (layer0_outputs(4432));
    layer1_outputs(8589) <= not(layer0_outputs(7583));
    layer1_outputs(8590) <= not((layer0_outputs(5800)) xor (layer0_outputs(240)));
    layer1_outputs(8591) <= not(layer0_outputs(8627));
    layer1_outputs(8592) <= not(layer0_outputs(8542));
    layer1_outputs(8593) <= not(layer0_outputs(10227)) or (layer0_outputs(11373));
    layer1_outputs(8594) <= not(layer0_outputs(9100)) or (layer0_outputs(6763));
    layer1_outputs(8595) <= not(layer0_outputs(10357));
    layer1_outputs(8596) <= layer0_outputs(4068);
    layer1_outputs(8597) <= '1';
    layer1_outputs(8598) <= (layer0_outputs(3575)) and not (layer0_outputs(6024));
    layer1_outputs(8599) <= layer0_outputs(10290);
    layer1_outputs(8600) <= not(layer0_outputs(4665)) or (layer0_outputs(5544));
    layer1_outputs(8601) <= not((layer0_outputs(7792)) and (layer0_outputs(7411)));
    layer1_outputs(8602) <= not(layer0_outputs(5193)) or (layer0_outputs(11537));
    layer1_outputs(8603) <= (layer0_outputs(4006)) xor (layer0_outputs(3431));
    layer1_outputs(8604) <= layer0_outputs(9393);
    layer1_outputs(8605) <= not(layer0_outputs(8789));
    layer1_outputs(8606) <= layer0_outputs(4162);
    layer1_outputs(8607) <= (layer0_outputs(4823)) and (layer0_outputs(234));
    layer1_outputs(8608) <= (layer0_outputs(8221)) and not (layer0_outputs(3593));
    layer1_outputs(8609) <= (layer0_outputs(6607)) or (layer0_outputs(7609));
    layer1_outputs(8610) <= layer0_outputs(6310);
    layer1_outputs(8611) <= not(layer0_outputs(8781));
    layer1_outputs(8612) <= not(layer0_outputs(1300)) or (layer0_outputs(7620));
    layer1_outputs(8613) <= not(layer0_outputs(6474));
    layer1_outputs(8614) <= (layer0_outputs(11623)) xor (layer0_outputs(11098));
    layer1_outputs(8615) <= (layer0_outputs(147)) xor (layer0_outputs(1514));
    layer1_outputs(8616) <= (layer0_outputs(4297)) and (layer0_outputs(6186));
    layer1_outputs(8617) <= not((layer0_outputs(731)) xor (layer0_outputs(8048)));
    layer1_outputs(8618) <= not(layer0_outputs(9483));
    layer1_outputs(8619) <= layer0_outputs(10039);
    layer1_outputs(8620) <= (layer0_outputs(12576)) and (layer0_outputs(8235));
    layer1_outputs(8621) <= layer0_outputs(2322);
    layer1_outputs(8622) <= layer0_outputs(6366);
    layer1_outputs(8623) <= not(layer0_outputs(9484)) or (layer0_outputs(12257));
    layer1_outputs(8624) <= (layer0_outputs(12322)) and not (layer0_outputs(3530));
    layer1_outputs(8625) <= (layer0_outputs(9839)) and not (layer0_outputs(1249));
    layer1_outputs(8626) <= not(layer0_outputs(558)) or (layer0_outputs(6911));
    layer1_outputs(8627) <= '0';
    layer1_outputs(8628) <= not(layer0_outputs(12274)) or (layer0_outputs(5680));
    layer1_outputs(8629) <= (layer0_outputs(3062)) or (layer0_outputs(4302));
    layer1_outputs(8630) <= layer0_outputs(9117);
    layer1_outputs(8631) <= not((layer0_outputs(4713)) or (layer0_outputs(9101)));
    layer1_outputs(8632) <= not((layer0_outputs(7513)) and (layer0_outputs(2653)));
    layer1_outputs(8633) <= not(layer0_outputs(11601)) or (layer0_outputs(10618));
    layer1_outputs(8634) <= layer0_outputs(1204);
    layer1_outputs(8635) <= not((layer0_outputs(1228)) and (layer0_outputs(7107)));
    layer1_outputs(8636) <= not(layer0_outputs(5342));
    layer1_outputs(8637) <= not(layer0_outputs(3881));
    layer1_outputs(8638) <= (layer0_outputs(8675)) xor (layer0_outputs(920));
    layer1_outputs(8639) <= layer0_outputs(9606);
    layer1_outputs(8640) <= (layer0_outputs(5669)) and not (layer0_outputs(8309));
    layer1_outputs(8641) <= (layer0_outputs(10239)) and not (layer0_outputs(12568));
    layer1_outputs(8642) <= not(layer0_outputs(7937));
    layer1_outputs(8643) <= not(layer0_outputs(5680));
    layer1_outputs(8644) <= not(layer0_outputs(9293)) or (layer0_outputs(4267));
    layer1_outputs(8645) <= (layer0_outputs(4485)) and (layer0_outputs(1592));
    layer1_outputs(8646) <= not(layer0_outputs(9825));
    layer1_outputs(8647) <= not((layer0_outputs(10400)) xor (layer0_outputs(4026)));
    layer1_outputs(8648) <= not(layer0_outputs(12340)) or (layer0_outputs(2123));
    layer1_outputs(8649) <= layer0_outputs(4697);
    layer1_outputs(8650) <= layer0_outputs(11075);
    layer1_outputs(8651) <= layer0_outputs(1739);
    layer1_outputs(8652) <= layer0_outputs(7794);
    layer1_outputs(8653) <= layer0_outputs(12533);
    layer1_outputs(8654) <= not((layer0_outputs(6780)) xor (layer0_outputs(11096)));
    layer1_outputs(8655) <= layer0_outputs(9804);
    layer1_outputs(8656) <= not(layer0_outputs(2799)) or (layer0_outputs(3746));
    layer1_outputs(8657) <= (layer0_outputs(4644)) and not (layer0_outputs(4021));
    layer1_outputs(8658) <= layer0_outputs(5290);
    layer1_outputs(8659) <= (layer0_outputs(3232)) and (layer0_outputs(4940));
    layer1_outputs(8660) <= (layer0_outputs(10401)) and (layer0_outputs(1005));
    layer1_outputs(8661) <= layer0_outputs(9538);
    layer1_outputs(8662) <= layer0_outputs(243);
    layer1_outputs(8663) <= layer0_outputs(2943);
    layer1_outputs(8664) <= not(layer0_outputs(12482));
    layer1_outputs(8665) <= layer0_outputs(6491);
    layer1_outputs(8666) <= not(layer0_outputs(6014));
    layer1_outputs(8667) <= (layer0_outputs(5842)) and not (layer0_outputs(9000));
    layer1_outputs(8668) <= '1';
    layer1_outputs(8669) <= not(layer0_outputs(2529));
    layer1_outputs(8670) <= (layer0_outputs(9848)) xor (layer0_outputs(4168));
    layer1_outputs(8671) <= layer0_outputs(820);
    layer1_outputs(8672) <= not((layer0_outputs(2531)) and (layer0_outputs(3974)));
    layer1_outputs(8673) <= (layer0_outputs(1825)) and (layer0_outputs(2393));
    layer1_outputs(8674) <= '0';
    layer1_outputs(8675) <= layer0_outputs(5663);
    layer1_outputs(8676) <= (layer0_outputs(12067)) and not (layer0_outputs(3658));
    layer1_outputs(8677) <= (layer0_outputs(5662)) and not (layer0_outputs(179));
    layer1_outputs(8678) <= '0';
    layer1_outputs(8679) <= not(layer0_outputs(10467));
    layer1_outputs(8680) <= not(layer0_outputs(367));
    layer1_outputs(8681) <= not(layer0_outputs(1007)) or (layer0_outputs(12192));
    layer1_outputs(8682) <= layer0_outputs(9854);
    layer1_outputs(8683) <= not(layer0_outputs(1893)) or (layer0_outputs(9678));
    layer1_outputs(8684) <= not(layer0_outputs(928)) or (layer0_outputs(11497));
    layer1_outputs(8685) <= not((layer0_outputs(6909)) or (layer0_outputs(4842)));
    layer1_outputs(8686) <= not(layer0_outputs(370));
    layer1_outputs(8687) <= (layer0_outputs(15)) xor (layer0_outputs(6601));
    layer1_outputs(8688) <= not(layer0_outputs(345));
    layer1_outputs(8689) <= not((layer0_outputs(5095)) xor (layer0_outputs(9218)));
    layer1_outputs(8690) <= not(layer0_outputs(6630)) or (layer0_outputs(10431));
    layer1_outputs(8691) <= layer0_outputs(11281);
    layer1_outputs(8692) <= layer0_outputs(3380);
    layer1_outputs(8693) <= not(layer0_outputs(10337)) or (layer0_outputs(4363));
    layer1_outputs(8694) <= not(layer0_outputs(9031)) or (layer0_outputs(3312));
    layer1_outputs(8695) <= layer0_outputs(12072);
    layer1_outputs(8696) <= not(layer0_outputs(6256));
    layer1_outputs(8697) <= (layer0_outputs(1811)) xor (layer0_outputs(426));
    layer1_outputs(8698) <= (layer0_outputs(10389)) xor (layer0_outputs(6573));
    layer1_outputs(8699) <= layer0_outputs(6120);
    layer1_outputs(8700) <= (layer0_outputs(8818)) or (layer0_outputs(3508));
    layer1_outputs(8701) <= not((layer0_outputs(6432)) or (layer0_outputs(1972)));
    layer1_outputs(8702) <= layer0_outputs(2242);
    layer1_outputs(8703) <= layer0_outputs(3476);
    layer1_outputs(8704) <= not(layer0_outputs(3044));
    layer1_outputs(8705) <= not(layer0_outputs(3479));
    layer1_outputs(8706) <= (layer0_outputs(5140)) and (layer0_outputs(474));
    layer1_outputs(8707) <= layer0_outputs(1177);
    layer1_outputs(8708) <= not(layer0_outputs(5004));
    layer1_outputs(8709) <= not(layer0_outputs(4926)) or (layer0_outputs(7861));
    layer1_outputs(8710) <= (layer0_outputs(7510)) or (layer0_outputs(7960));
    layer1_outputs(8711) <= (layer0_outputs(6286)) and (layer0_outputs(2893));
    layer1_outputs(8712) <= not((layer0_outputs(9080)) and (layer0_outputs(8474)));
    layer1_outputs(8713) <= not(layer0_outputs(9985));
    layer1_outputs(8714) <= not((layer0_outputs(10372)) xor (layer0_outputs(2923)));
    layer1_outputs(8715) <= not(layer0_outputs(4209));
    layer1_outputs(8716) <= (layer0_outputs(11489)) and not (layer0_outputs(3477));
    layer1_outputs(8717) <= layer0_outputs(3232);
    layer1_outputs(8718) <= not(layer0_outputs(2574)) or (layer0_outputs(4339));
    layer1_outputs(8719) <= not(layer0_outputs(1638));
    layer1_outputs(8720) <= not((layer0_outputs(5280)) or (layer0_outputs(8582)));
    layer1_outputs(8721) <= not(layer0_outputs(11006));
    layer1_outputs(8722) <= layer0_outputs(6996);
    layer1_outputs(8723) <= (layer0_outputs(4088)) or (layer0_outputs(8025));
    layer1_outputs(8724) <= not(layer0_outputs(8391));
    layer1_outputs(8725) <= (layer0_outputs(262)) and not (layer0_outputs(5296));
    layer1_outputs(8726) <= layer0_outputs(8406);
    layer1_outputs(8727) <= (layer0_outputs(10343)) and not (layer0_outputs(3875));
    layer1_outputs(8728) <= layer0_outputs(11430);
    layer1_outputs(8729) <= not(layer0_outputs(7940));
    layer1_outputs(8730) <= not((layer0_outputs(7373)) xor (layer0_outputs(12045)));
    layer1_outputs(8731) <= not(layer0_outputs(8009)) or (layer0_outputs(10840));
    layer1_outputs(8732) <= not(layer0_outputs(2005));
    layer1_outputs(8733) <= not(layer0_outputs(3019));
    layer1_outputs(8734) <= (layer0_outputs(627)) and not (layer0_outputs(4500));
    layer1_outputs(8735) <= not(layer0_outputs(4911));
    layer1_outputs(8736) <= layer0_outputs(5610);
    layer1_outputs(8737) <= (layer0_outputs(3295)) or (layer0_outputs(8202));
    layer1_outputs(8738) <= not((layer0_outputs(583)) xor (layer0_outputs(9960)));
    layer1_outputs(8739) <= layer0_outputs(6211);
    layer1_outputs(8740) <= '1';
    layer1_outputs(8741) <= layer0_outputs(11647);
    layer1_outputs(8742) <= not(layer0_outputs(7036)) or (layer0_outputs(11947));
    layer1_outputs(8743) <= not((layer0_outputs(9676)) and (layer0_outputs(1126)));
    layer1_outputs(8744) <= not(layer0_outputs(6036));
    layer1_outputs(8745) <= not(layer0_outputs(9421));
    layer1_outputs(8746) <= not((layer0_outputs(11452)) and (layer0_outputs(10803)));
    layer1_outputs(8747) <= layer0_outputs(9256);
    layer1_outputs(8748) <= (layer0_outputs(11958)) and (layer0_outputs(6057));
    layer1_outputs(8749) <= not((layer0_outputs(8427)) or (layer0_outputs(9137)));
    layer1_outputs(8750) <= not(layer0_outputs(6086));
    layer1_outputs(8751) <= (layer0_outputs(11534)) and (layer0_outputs(696));
    layer1_outputs(8752) <= '0';
    layer1_outputs(8753) <= not(layer0_outputs(6584));
    layer1_outputs(8754) <= not(layer0_outputs(226));
    layer1_outputs(8755) <= not((layer0_outputs(1555)) or (layer0_outputs(1490)));
    layer1_outputs(8756) <= not((layer0_outputs(12380)) and (layer0_outputs(5442)));
    layer1_outputs(8757) <= layer0_outputs(959);
    layer1_outputs(8758) <= (layer0_outputs(3482)) or (layer0_outputs(5100));
    layer1_outputs(8759) <= (layer0_outputs(5497)) or (layer0_outputs(4932));
    layer1_outputs(8760) <= layer0_outputs(7868);
    layer1_outputs(8761) <= not(layer0_outputs(1975));
    layer1_outputs(8762) <= not(layer0_outputs(5145)) or (layer0_outputs(6961));
    layer1_outputs(8763) <= (layer0_outputs(10335)) and (layer0_outputs(508));
    layer1_outputs(8764) <= layer0_outputs(12191);
    layer1_outputs(8765) <= not(layer0_outputs(8707));
    layer1_outputs(8766) <= not(layer0_outputs(11092));
    layer1_outputs(8767) <= '0';
    layer1_outputs(8768) <= (layer0_outputs(12218)) and not (layer0_outputs(1055));
    layer1_outputs(8769) <= not((layer0_outputs(2819)) or (layer0_outputs(6354)));
    layer1_outputs(8770) <= layer0_outputs(5376);
    layer1_outputs(8771) <= not(layer0_outputs(7483));
    layer1_outputs(8772) <= (layer0_outputs(8496)) and not (layer0_outputs(3268));
    layer1_outputs(8773) <= layer0_outputs(1659);
    layer1_outputs(8774) <= not(layer0_outputs(1417)) or (layer0_outputs(12002));
    layer1_outputs(8775) <= (layer0_outputs(2868)) xor (layer0_outputs(9371));
    layer1_outputs(8776) <= not((layer0_outputs(7665)) or (layer0_outputs(10323)));
    layer1_outputs(8777) <= (layer0_outputs(10586)) or (layer0_outputs(3250));
    layer1_outputs(8778) <= not((layer0_outputs(7687)) and (layer0_outputs(356)));
    layer1_outputs(8779) <= (layer0_outputs(1732)) and not (layer0_outputs(8958));
    layer1_outputs(8780) <= (layer0_outputs(6126)) and (layer0_outputs(8292));
    layer1_outputs(8781) <= (layer0_outputs(2897)) and (layer0_outputs(10438));
    layer1_outputs(8782) <= (layer0_outputs(10595)) or (layer0_outputs(2954));
    layer1_outputs(8783) <= not((layer0_outputs(283)) or (layer0_outputs(4503)));
    layer1_outputs(8784) <= (layer0_outputs(2077)) and not (layer0_outputs(5024));
    layer1_outputs(8785) <= not((layer0_outputs(11103)) xor (layer0_outputs(11599)));
    layer1_outputs(8786) <= not(layer0_outputs(4811)) or (layer0_outputs(2966));
    layer1_outputs(8787) <= (layer0_outputs(8925)) and (layer0_outputs(4542));
    layer1_outputs(8788) <= '1';
    layer1_outputs(8789) <= (layer0_outputs(3554)) xor (layer0_outputs(4580));
    layer1_outputs(8790) <= not(layer0_outputs(2785));
    layer1_outputs(8791) <= not(layer0_outputs(1486)) or (layer0_outputs(8243));
    layer1_outputs(8792) <= not((layer0_outputs(4093)) xor (layer0_outputs(1687)));
    layer1_outputs(8793) <= not((layer0_outputs(5186)) and (layer0_outputs(10654)));
    layer1_outputs(8794) <= not(layer0_outputs(4022));
    layer1_outputs(8795) <= '0';
    layer1_outputs(8796) <= not(layer0_outputs(6532)) or (layer0_outputs(3530));
    layer1_outputs(8797) <= not((layer0_outputs(374)) xor (layer0_outputs(10015)));
    layer1_outputs(8798) <= not(layer0_outputs(3500)) or (layer0_outputs(6306));
    layer1_outputs(8799) <= not(layer0_outputs(3650)) or (layer0_outputs(4578));
    layer1_outputs(8800) <= not((layer0_outputs(5018)) and (layer0_outputs(7313)));
    layer1_outputs(8801) <= not(layer0_outputs(5917));
    layer1_outputs(8802) <= (layer0_outputs(3197)) and (layer0_outputs(5739));
    layer1_outputs(8803) <= not((layer0_outputs(1388)) xor (layer0_outputs(8043)));
    layer1_outputs(8804) <= not(layer0_outputs(9785));
    layer1_outputs(8805) <= layer0_outputs(12741);
    layer1_outputs(8806) <= (layer0_outputs(7949)) xor (layer0_outputs(1697));
    layer1_outputs(8807) <= (layer0_outputs(3129)) and not (layer0_outputs(4632));
    layer1_outputs(8808) <= (layer0_outputs(5400)) or (layer0_outputs(10013));
    layer1_outputs(8809) <= (layer0_outputs(12547)) or (layer0_outputs(1006));
    layer1_outputs(8810) <= not(layer0_outputs(2079)) or (layer0_outputs(4687));
    layer1_outputs(8811) <= (layer0_outputs(8339)) and not (layer0_outputs(1705));
    layer1_outputs(8812) <= not(layer0_outputs(3945));
    layer1_outputs(8813) <= not((layer0_outputs(3634)) xor (layer0_outputs(5338)));
    layer1_outputs(8814) <= layer0_outputs(9997);
    layer1_outputs(8815) <= (layer0_outputs(7290)) or (layer0_outputs(12368));
    layer1_outputs(8816) <= layer0_outputs(7835);
    layer1_outputs(8817) <= not((layer0_outputs(2472)) or (layer0_outputs(10744)));
    layer1_outputs(8818) <= not((layer0_outputs(1700)) or (layer0_outputs(704)));
    layer1_outputs(8819) <= (layer0_outputs(3465)) or (layer0_outputs(5075));
    layer1_outputs(8820) <= not((layer0_outputs(12506)) xor (layer0_outputs(5943)));
    layer1_outputs(8821) <= not((layer0_outputs(7766)) xor (layer0_outputs(8390)));
    layer1_outputs(8822) <= (layer0_outputs(7812)) and not (layer0_outputs(10908));
    layer1_outputs(8823) <= not((layer0_outputs(1513)) and (layer0_outputs(6745)));
    layer1_outputs(8824) <= not(layer0_outputs(6569));
    layer1_outputs(8825) <= not(layer0_outputs(4360)) or (layer0_outputs(3286));
    layer1_outputs(8826) <= layer0_outputs(3785);
    layer1_outputs(8827) <= (layer0_outputs(1261)) and (layer0_outputs(2126));
    layer1_outputs(8828) <= not((layer0_outputs(7753)) xor (layer0_outputs(7484)));
    layer1_outputs(8829) <= not(layer0_outputs(6200));
    layer1_outputs(8830) <= not(layer0_outputs(11166));
    layer1_outputs(8831) <= not(layer0_outputs(5890)) or (layer0_outputs(12065));
    layer1_outputs(8832) <= layer0_outputs(8947);
    layer1_outputs(8833) <= '1';
    layer1_outputs(8834) <= not(layer0_outputs(8244));
    layer1_outputs(8835) <= (layer0_outputs(2217)) or (layer0_outputs(261));
    layer1_outputs(8836) <= (layer0_outputs(7884)) and not (layer0_outputs(12240));
    layer1_outputs(8837) <= not(layer0_outputs(7733)) or (layer0_outputs(10366));
    layer1_outputs(8838) <= (layer0_outputs(2454)) and not (layer0_outputs(10752));
    layer1_outputs(8839) <= not((layer0_outputs(8612)) xor (layer0_outputs(10150)));
    layer1_outputs(8840) <= '0';
    layer1_outputs(8841) <= layer0_outputs(8931);
    layer1_outputs(8842) <= not(layer0_outputs(6969));
    layer1_outputs(8843) <= not(layer0_outputs(10097)) or (layer0_outputs(5671));
    layer1_outputs(8844) <= layer0_outputs(445);
    layer1_outputs(8845) <= layer0_outputs(9223);
    layer1_outputs(8846) <= (layer0_outputs(12224)) and not (layer0_outputs(11498));
    layer1_outputs(8847) <= not(layer0_outputs(5530));
    layer1_outputs(8848) <= not(layer0_outputs(606));
    layer1_outputs(8849) <= not(layer0_outputs(1427)) or (layer0_outputs(2706));
    layer1_outputs(8850) <= not((layer0_outputs(9192)) and (layer0_outputs(7192)));
    layer1_outputs(8851) <= not((layer0_outputs(1920)) xor (layer0_outputs(968)));
    layer1_outputs(8852) <= (layer0_outputs(10229)) and not (layer0_outputs(4641));
    layer1_outputs(8853) <= (layer0_outputs(3711)) and not (layer0_outputs(3167));
    layer1_outputs(8854) <= not(layer0_outputs(10031)) or (layer0_outputs(8076));
    layer1_outputs(8855) <= not(layer0_outputs(184));
    layer1_outputs(8856) <= not(layer0_outputs(5004));
    layer1_outputs(8857) <= (layer0_outputs(3748)) and not (layer0_outputs(7638));
    layer1_outputs(8858) <= (layer0_outputs(10660)) and (layer0_outputs(10891));
    layer1_outputs(8859) <= layer0_outputs(7584);
    layer1_outputs(8860) <= not(layer0_outputs(5939));
    layer1_outputs(8861) <= (layer0_outputs(1624)) or (layer0_outputs(778));
    layer1_outputs(8862) <= (layer0_outputs(568)) and (layer0_outputs(12483));
    layer1_outputs(8863) <= not(layer0_outputs(9242)) or (layer0_outputs(7044));
    layer1_outputs(8864) <= (layer0_outputs(523)) and not (layer0_outputs(6346));
    layer1_outputs(8865) <= not(layer0_outputs(11567));
    layer1_outputs(8866) <= not(layer0_outputs(12397));
    layer1_outputs(8867) <= (layer0_outputs(2347)) and (layer0_outputs(3760));
    layer1_outputs(8868) <= not((layer0_outputs(7979)) or (layer0_outputs(502)));
    layer1_outputs(8869) <= (layer0_outputs(5523)) and not (layer0_outputs(5099));
    layer1_outputs(8870) <= (layer0_outputs(4709)) and not (layer0_outputs(9522));
    layer1_outputs(8871) <= '0';
    layer1_outputs(8872) <= (layer0_outputs(1895)) and not (layer0_outputs(9666));
    layer1_outputs(8873) <= layer0_outputs(11602);
    layer1_outputs(8874) <= (layer0_outputs(6450)) and not (layer0_outputs(5345));
    layer1_outputs(8875) <= '0';
    layer1_outputs(8876) <= layer0_outputs(817);
    layer1_outputs(8877) <= layer0_outputs(5187);
    layer1_outputs(8878) <= not(layer0_outputs(10976));
    layer1_outputs(8879) <= not((layer0_outputs(79)) and (layer0_outputs(7380)));
    layer1_outputs(8880) <= not((layer0_outputs(1312)) and (layer0_outputs(5126)));
    layer1_outputs(8881) <= (layer0_outputs(3674)) and not (layer0_outputs(4769));
    layer1_outputs(8882) <= not(layer0_outputs(8011)) or (layer0_outputs(12602));
    layer1_outputs(8883) <= not(layer0_outputs(4174));
    layer1_outputs(8884) <= not(layer0_outputs(6312));
    layer1_outputs(8885) <= (layer0_outputs(4525)) and not (layer0_outputs(7872));
    layer1_outputs(8886) <= '1';
    layer1_outputs(8887) <= not(layer0_outputs(3325));
    layer1_outputs(8888) <= not((layer0_outputs(119)) xor (layer0_outputs(6948)));
    layer1_outputs(8889) <= '1';
    layer1_outputs(8890) <= not(layer0_outputs(7555)) or (layer0_outputs(2958));
    layer1_outputs(8891) <= (layer0_outputs(7581)) and not (layer0_outputs(9743));
    layer1_outputs(8892) <= not(layer0_outputs(10084)) or (layer0_outputs(4119));
    layer1_outputs(8893) <= (layer0_outputs(7131)) and not (layer0_outputs(5332));
    layer1_outputs(8894) <= (layer0_outputs(11892)) and not (layer0_outputs(11744));
    layer1_outputs(8895) <= layer0_outputs(3152);
    layer1_outputs(8896) <= '0';
    layer1_outputs(8897) <= (layer0_outputs(7005)) and not (layer0_outputs(11576));
    layer1_outputs(8898) <= '0';
    layer1_outputs(8899) <= not(layer0_outputs(11671));
    layer1_outputs(8900) <= not(layer0_outputs(2676));
    layer1_outputs(8901) <= (layer0_outputs(6923)) and not (layer0_outputs(1305));
    layer1_outputs(8902) <= layer0_outputs(11216);
    layer1_outputs(8903) <= (layer0_outputs(11766)) or (layer0_outputs(9105));
    layer1_outputs(8904) <= not(layer0_outputs(11931)) or (layer0_outputs(9245));
    layer1_outputs(8905) <= layer0_outputs(5337);
    layer1_outputs(8906) <= '1';
    layer1_outputs(8907) <= not(layer0_outputs(12487));
    layer1_outputs(8908) <= not(layer0_outputs(8445)) or (layer0_outputs(2209));
    layer1_outputs(8909) <= layer0_outputs(1338);
    layer1_outputs(8910) <= '0';
    layer1_outputs(8911) <= not(layer0_outputs(9404)) or (layer0_outputs(11127));
    layer1_outputs(8912) <= (layer0_outputs(8058)) and (layer0_outputs(1386));
    layer1_outputs(8913) <= not(layer0_outputs(7565)) or (layer0_outputs(3948));
    layer1_outputs(8914) <= not(layer0_outputs(847));
    layer1_outputs(8915) <= not(layer0_outputs(4126));
    layer1_outputs(8916) <= not(layer0_outputs(4701));
    layer1_outputs(8917) <= not((layer0_outputs(2683)) and (layer0_outputs(4233)));
    layer1_outputs(8918) <= not((layer0_outputs(5265)) and (layer0_outputs(12370)));
    layer1_outputs(8919) <= layer0_outputs(8412);
    layer1_outputs(8920) <= layer0_outputs(2018);
    layer1_outputs(8921) <= (layer0_outputs(6937)) xor (layer0_outputs(3475));
    layer1_outputs(8922) <= not(layer0_outputs(3580));
    layer1_outputs(8923) <= layer0_outputs(124);
    layer1_outputs(8924) <= layer0_outputs(8852);
    layer1_outputs(8925) <= (layer0_outputs(11021)) and not (layer0_outputs(7481));
    layer1_outputs(8926) <= not((layer0_outputs(2257)) and (layer0_outputs(4621)));
    layer1_outputs(8927) <= (layer0_outputs(5807)) and not (layer0_outputs(3830));
    layer1_outputs(8928) <= (layer0_outputs(11713)) or (layer0_outputs(8148));
    layer1_outputs(8929) <= (layer0_outputs(1323)) and (layer0_outputs(10083));
    layer1_outputs(8930) <= not(layer0_outputs(2841)) or (layer0_outputs(1878));
    layer1_outputs(8931) <= (layer0_outputs(975)) xor (layer0_outputs(8079));
    layer1_outputs(8932) <= not(layer0_outputs(7220));
    layer1_outputs(8933) <= not((layer0_outputs(3329)) or (layer0_outputs(6271)));
    layer1_outputs(8934) <= layer0_outputs(12623);
    layer1_outputs(8935) <= (layer0_outputs(12138)) or (layer0_outputs(11201));
    layer1_outputs(8936) <= (layer0_outputs(246)) and not (layer0_outputs(2323));
    layer1_outputs(8937) <= (layer0_outputs(4721)) and not (layer0_outputs(3937));
    layer1_outputs(8938) <= (layer0_outputs(10291)) or (layer0_outputs(5765));
    layer1_outputs(8939) <= not(layer0_outputs(1492)) or (layer0_outputs(2099));
    layer1_outputs(8940) <= (layer0_outputs(5346)) xor (layer0_outputs(7600));
    layer1_outputs(8941) <= not((layer0_outputs(2147)) and (layer0_outputs(4799)));
    layer1_outputs(8942) <= not(layer0_outputs(9597)) or (layer0_outputs(7710));
    layer1_outputs(8943) <= not(layer0_outputs(3706));
    layer1_outputs(8944) <= '0';
    layer1_outputs(8945) <= layer0_outputs(2354);
    layer1_outputs(8946) <= not(layer0_outputs(8660)) or (layer0_outputs(9246));
    layer1_outputs(8947) <= not(layer0_outputs(11715)) or (layer0_outputs(10816));
    layer1_outputs(8948) <= (layer0_outputs(1995)) or (layer0_outputs(4712));
    layer1_outputs(8949) <= not((layer0_outputs(6062)) xor (layer0_outputs(8833)));
    layer1_outputs(8950) <= (layer0_outputs(8471)) and not (layer0_outputs(10258));
    layer1_outputs(8951) <= not(layer0_outputs(4113));
    layer1_outputs(8952) <= layer0_outputs(7506);
    layer1_outputs(8953) <= not(layer0_outputs(2428)) or (layer0_outputs(10723));
    layer1_outputs(8954) <= not(layer0_outputs(7362));
    layer1_outputs(8955) <= layer0_outputs(11034);
    layer1_outputs(8956) <= not((layer0_outputs(3617)) and (layer0_outputs(6078)));
    layer1_outputs(8957) <= not(layer0_outputs(4920));
    layer1_outputs(8958) <= not(layer0_outputs(8530));
    layer1_outputs(8959) <= not(layer0_outputs(2844));
    layer1_outputs(8960) <= not((layer0_outputs(3125)) xor (layer0_outputs(3968)));
    layer1_outputs(8961) <= (layer0_outputs(1352)) and not (layer0_outputs(4089));
    layer1_outputs(8962) <= not((layer0_outputs(12336)) or (layer0_outputs(3080)));
    layer1_outputs(8963) <= not((layer0_outputs(4226)) and (layer0_outputs(7590)));
    layer1_outputs(8964) <= not(layer0_outputs(2931)) or (layer0_outputs(4218));
    layer1_outputs(8965) <= not(layer0_outputs(12776)) or (layer0_outputs(6165));
    layer1_outputs(8966) <= not(layer0_outputs(4335)) or (layer0_outputs(12329));
    layer1_outputs(8967) <= not(layer0_outputs(1835));
    layer1_outputs(8968) <= layer0_outputs(12665);
    layer1_outputs(8969) <= not((layer0_outputs(8353)) or (layer0_outputs(4109)));
    layer1_outputs(8970) <= (layer0_outputs(4051)) or (layer0_outputs(8017));
    layer1_outputs(8971) <= (layer0_outputs(4575)) or (layer0_outputs(11139));
    layer1_outputs(8972) <= (layer0_outputs(9450)) and (layer0_outputs(12011));
    layer1_outputs(8973) <= layer0_outputs(5654);
    layer1_outputs(8974) <= layer0_outputs(5436);
    layer1_outputs(8975) <= (layer0_outputs(3192)) and not (layer0_outputs(6568));
    layer1_outputs(8976) <= layer0_outputs(10973);
    layer1_outputs(8977) <= not(layer0_outputs(9576)) or (layer0_outputs(2135));
    layer1_outputs(8978) <= not((layer0_outputs(6329)) xor (layer0_outputs(6052)));
    layer1_outputs(8979) <= not(layer0_outputs(11334)) or (layer0_outputs(2185));
    layer1_outputs(8980) <= not((layer0_outputs(10058)) xor (layer0_outputs(3447)));
    layer1_outputs(8981) <= layer0_outputs(2035);
    layer1_outputs(8982) <= '0';
    layer1_outputs(8983) <= (layer0_outputs(6998)) and not (layer0_outputs(3631));
    layer1_outputs(8984) <= (layer0_outputs(7444)) or (layer0_outputs(2020));
    layer1_outputs(8985) <= (layer0_outputs(3437)) and not (layer0_outputs(10861));
    layer1_outputs(8986) <= (layer0_outputs(2151)) or (layer0_outputs(4148));
    layer1_outputs(8987) <= (layer0_outputs(1422)) and not (layer0_outputs(5957));
    layer1_outputs(8988) <= not(layer0_outputs(474)) or (layer0_outputs(8161));
    layer1_outputs(8989) <= not(layer0_outputs(11724)) or (layer0_outputs(3630));
    layer1_outputs(8990) <= (layer0_outputs(10080)) and not (layer0_outputs(3184));
    layer1_outputs(8991) <= not(layer0_outputs(12191));
    layer1_outputs(8992) <= '0';
    layer1_outputs(8993) <= not(layer0_outputs(10288));
    layer1_outputs(8994) <= layer0_outputs(10686);
    layer1_outputs(8995) <= not((layer0_outputs(6525)) and (layer0_outputs(11857)));
    layer1_outputs(8996) <= not(layer0_outputs(1197));
    layer1_outputs(8997) <= not((layer0_outputs(2877)) and (layer0_outputs(9770)));
    layer1_outputs(8998) <= not(layer0_outputs(4155)) or (layer0_outputs(1252));
    layer1_outputs(8999) <= layer0_outputs(2075);
    layer1_outputs(9000) <= not(layer0_outputs(9243));
    layer1_outputs(9001) <= not(layer0_outputs(1983));
    layer1_outputs(9002) <= layer0_outputs(11474);
    layer1_outputs(9003) <= (layer0_outputs(3218)) and not (layer0_outputs(3091));
    layer1_outputs(9004) <= layer0_outputs(5353);
    layer1_outputs(9005) <= not(layer0_outputs(1071)) or (layer0_outputs(12029));
    layer1_outputs(9006) <= not(layer0_outputs(4735));
    layer1_outputs(9007) <= not((layer0_outputs(608)) and (layer0_outputs(8260)));
    layer1_outputs(9008) <= not(layer0_outputs(5258));
    layer1_outputs(9009) <= (layer0_outputs(3177)) xor (layer0_outputs(9107));
    layer1_outputs(9010) <= layer0_outputs(6377);
    layer1_outputs(9011) <= (layer0_outputs(5103)) and (layer0_outputs(9946));
    layer1_outputs(9012) <= (layer0_outputs(11009)) xor (layer0_outputs(578));
    layer1_outputs(9013) <= (layer0_outputs(6056)) xor (layer0_outputs(7040));
    layer1_outputs(9014) <= (layer0_outputs(3110)) and (layer0_outputs(12394));
    layer1_outputs(9015) <= not(layer0_outputs(11225));
    layer1_outputs(9016) <= not((layer0_outputs(8708)) xor (layer0_outputs(8604)));
    layer1_outputs(9017) <= (layer0_outputs(1106)) xor (layer0_outputs(3301));
    layer1_outputs(9018) <= layer0_outputs(1612);
    layer1_outputs(9019) <= '1';
    layer1_outputs(9020) <= (layer0_outputs(2422)) xor (layer0_outputs(8928));
    layer1_outputs(9021) <= not(layer0_outputs(4898));
    layer1_outputs(9022) <= not((layer0_outputs(7271)) and (layer0_outputs(50)));
    layer1_outputs(9023) <= (layer0_outputs(7120)) and not (layer0_outputs(6270));
    layer1_outputs(9024) <= layer0_outputs(10155);
    layer1_outputs(9025) <= not(layer0_outputs(663)) or (layer0_outputs(12476));
    layer1_outputs(9026) <= not(layer0_outputs(3041));
    layer1_outputs(9027) <= not(layer0_outputs(7279));
    layer1_outputs(9028) <= not((layer0_outputs(2410)) and (layer0_outputs(10786)));
    layer1_outputs(9029) <= (layer0_outputs(2329)) and (layer0_outputs(8448));
    layer1_outputs(9030) <= not((layer0_outputs(5678)) or (layer0_outputs(2465)));
    layer1_outputs(9031) <= layer0_outputs(12702);
    layer1_outputs(9032) <= not(layer0_outputs(8849));
    layer1_outputs(9033) <= not(layer0_outputs(5299)) or (layer0_outputs(3375));
    layer1_outputs(9034) <= layer0_outputs(6813);
    layer1_outputs(9035) <= not((layer0_outputs(5143)) or (layer0_outputs(11023)));
    layer1_outputs(9036) <= not((layer0_outputs(10169)) or (layer0_outputs(11585)));
    layer1_outputs(9037) <= not(layer0_outputs(9220));
    layer1_outputs(9038) <= (layer0_outputs(28)) or (layer0_outputs(5649));
    layer1_outputs(9039) <= (layer0_outputs(7592)) xor (layer0_outputs(7564));
    layer1_outputs(9040) <= layer0_outputs(9874);
    layer1_outputs(9041) <= not(layer0_outputs(12280));
    layer1_outputs(9042) <= layer0_outputs(10313);
    layer1_outputs(9043) <= '0';
    layer1_outputs(9044) <= layer0_outputs(10580);
    layer1_outputs(9045) <= not(layer0_outputs(200));
    layer1_outputs(9046) <= not(layer0_outputs(8201));
    layer1_outputs(9047) <= (layer0_outputs(1400)) and not (layer0_outputs(9896));
    layer1_outputs(9048) <= layer0_outputs(9457);
    layer1_outputs(9049) <= not((layer0_outputs(195)) and (layer0_outputs(10204)));
    layer1_outputs(9050) <= not(layer0_outputs(7601));
    layer1_outputs(9051) <= (layer0_outputs(1976)) and not (layer0_outputs(8179));
    layer1_outputs(9052) <= not((layer0_outputs(7977)) or (layer0_outputs(7920)));
    layer1_outputs(9053) <= (layer0_outputs(1886)) and not (layer0_outputs(4124));
    layer1_outputs(9054) <= not(layer0_outputs(1868));
    layer1_outputs(9055) <= (layer0_outputs(535)) and not (layer0_outputs(1959));
    layer1_outputs(9056) <= '1';
    layer1_outputs(9057) <= not(layer0_outputs(2539));
    layer1_outputs(9058) <= not(layer0_outputs(260)) or (layer0_outputs(1842));
    layer1_outputs(9059) <= (layer0_outputs(310)) and (layer0_outputs(2925));
    layer1_outputs(9060) <= (layer0_outputs(4987)) and not (layer0_outputs(5087));
    layer1_outputs(9061) <= not(layer0_outputs(4126)) or (layer0_outputs(9790));
    layer1_outputs(9062) <= (layer0_outputs(7384)) and not (layer0_outputs(1540));
    layer1_outputs(9063) <= '0';
    layer1_outputs(9064) <= not(layer0_outputs(9290)) or (layer0_outputs(9087));
    layer1_outputs(9065) <= layer0_outputs(1532);
    layer1_outputs(9066) <= not(layer0_outputs(7622)) or (layer0_outputs(4332));
    layer1_outputs(9067) <= not((layer0_outputs(7299)) and (layer0_outputs(8449)));
    layer1_outputs(9068) <= '0';
    layer1_outputs(9069) <= layer0_outputs(1787);
    layer1_outputs(9070) <= layer0_outputs(1378);
    layer1_outputs(9071) <= (layer0_outputs(6756)) or (layer0_outputs(11780));
    layer1_outputs(9072) <= layer0_outputs(2609);
    layer1_outputs(9073) <= (layer0_outputs(9880)) and (layer0_outputs(10812));
    layer1_outputs(9074) <= layer0_outputs(5926);
    layer1_outputs(9075) <= not((layer0_outputs(2778)) or (layer0_outputs(817)));
    layer1_outputs(9076) <= not((layer0_outputs(9084)) and (layer0_outputs(2206)));
    layer1_outputs(9077) <= layer0_outputs(5330);
    layer1_outputs(9078) <= not(layer0_outputs(8499));
    layer1_outputs(9079) <= not(layer0_outputs(3969));
    layer1_outputs(9080) <= not(layer0_outputs(10507));
    layer1_outputs(9081) <= not(layer0_outputs(9276));
    layer1_outputs(9082) <= not((layer0_outputs(2482)) and (layer0_outputs(12567)));
    layer1_outputs(9083) <= not(layer0_outputs(12418));
    layer1_outputs(9084) <= not((layer0_outputs(4573)) xor (layer0_outputs(4889)));
    layer1_outputs(9085) <= layer0_outputs(3470);
    layer1_outputs(9086) <= (layer0_outputs(11269)) or (layer0_outputs(6831));
    layer1_outputs(9087) <= not(layer0_outputs(9669));
    layer1_outputs(9088) <= not((layer0_outputs(3426)) xor (layer0_outputs(1217)));
    layer1_outputs(9089) <= (layer0_outputs(10233)) xor (layer0_outputs(7359));
    layer1_outputs(9090) <= not((layer0_outputs(7418)) xor (layer0_outputs(3645)));
    layer1_outputs(9091) <= (layer0_outputs(11122)) and (layer0_outputs(7080));
    layer1_outputs(9092) <= (layer0_outputs(2594)) and not (layer0_outputs(11148));
    layer1_outputs(9093) <= not(layer0_outputs(5793));
    layer1_outputs(9094) <= not((layer0_outputs(11815)) and (layer0_outputs(11681)));
    layer1_outputs(9095) <= (layer0_outputs(1179)) xor (layer0_outputs(12490));
    layer1_outputs(9096) <= not(layer0_outputs(3808));
    layer1_outputs(9097) <= layer0_outputs(1519);
    layer1_outputs(9098) <= layer0_outputs(4600);
    layer1_outputs(9099) <= (layer0_outputs(5459)) xor (layer0_outputs(536));
    layer1_outputs(9100) <= layer0_outputs(3937);
    layer1_outputs(9101) <= layer0_outputs(12448);
    layer1_outputs(9102) <= (layer0_outputs(2915)) or (layer0_outputs(7880));
    layer1_outputs(9103) <= not(layer0_outputs(2816)) or (layer0_outputs(5983));
    layer1_outputs(9104) <= not(layer0_outputs(10493));
    layer1_outputs(9105) <= (layer0_outputs(3985)) and not (layer0_outputs(11859));
    layer1_outputs(9106) <= not((layer0_outputs(5255)) xor (layer0_outputs(5424)));
    layer1_outputs(9107) <= (layer0_outputs(9869)) and (layer0_outputs(3992));
    layer1_outputs(9108) <= not((layer0_outputs(3770)) and (layer0_outputs(5321)));
    layer1_outputs(9109) <= (layer0_outputs(6201)) and not (layer0_outputs(522));
    layer1_outputs(9110) <= not(layer0_outputs(10429));
    layer1_outputs(9111) <= (layer0_outputs(176)) or (layer0_outputs(5054));
    layer1_outputs(9112) <= not((layer0_outputs(7674)) or (layer0_outputs(8844)));
    layer1_outputs(9113) <= not(layer0_outputs(2626)) or (layer0_outputs(12736));
    layer1_outputs(9114) <= not(layer0_outputs(5267)) or (layer0_outputs(6725));
    layer1_outputs(9115) <= not(layer0_outputs(12782));
    layer1_outputs(9116) <= not((layer0_outputs(12740)) or (layer0_outputs(8044)));
    layer1_outputs(9117) <= '1';
    layer1_outputs(9118) <= not(layer0_outputs(12505)) or (layer0_outputs(2662));
    layer1_outputs(9119) <= not(layer0_outputs(12345));
    layer1_outputs(9120) <= not(layer0_outputs(11740));
    layer1_outputs(9121) <= layer0_outputs(4890);
    layer1_outputs(9122) <= (layer0_outputs(10255)) and not (layer0_outputs(6535));
    layer1_outputs(9123) <= (layer0_outputs(11596)) xor (layer0_outputs(11716));
    layer1_outputs(9124) <= not((layer0_outputs(12652)) or (layer0_outputs(10296)));
    layer1_outputs(9125) <= not((layer0_outputs(11226)) and (layer0_outputs(9547)));
    layer1_outputs(9126) <= not(layer0_outputs(9132));
    layer1_outputs(9127) <= not(layer0_outputs(2996));
    layer1_outputs(9128) <= not(layer0_outputs(9581)) or (layer0_outputs(12239));
    layer1_outputs(9129) <= (layer0_outputs(3778)) xor (layer0_outputs(8498));
    layer1_outputs(9130) <= not(layer0_outputs(378));
    layer1_outputs(9131) <= not(layer0_outputs(4810)) or (layer0_outputs(3570));
    layer1_outputs(9132) <= not((layer0_outputs(5690)) xor (layer0_outputs(9177)));
    layer1_outputs(9133) <= not(layer0_outputs(4356));
    layer1_outputs(9134) <= (layer0_outputs(5389)) and not (layer0_outputs(3939));
    layer1_outputs(9135) <= (layer0_outputs(9632)) and not (layer0_outputs(2063));
    layer1_outputs(9136) <= (layer0_outputs(7382)) or (layer0_outputs(8354));
    layer1_outputs(9137) <= (layer0_outputs(10082)) and not (layer0_outputs(3728));
    layer1_outputs(9138) <= not(layer0_outputs(5557));
    layer1_outputs(9139) <= layer0_outputs(3980);
    layer1_outputs(9140) <= not(layer0_outputs(7456));
    layer1_outputs(9141) <= (layer0_outputs(4387)) and not (layer0_outputs(6665));
    layer1_outputs(9142) <= (layer0_outputs(3360)) and (layer0_outputs(3542));
    layer1_outputs(9143) <= not(layer0_outputs(7222));
    layer1_outputs(9144) <= (layer0_outputs(12747)) or (layer0_outputs(7072));
    layer1_outputs(9145) <= not(layer0_outputs(3658));
    layer1_outputs(9146) <= not(layer0_outputs(9020));
    layer1_outputs(9147) <= layer0_outputs(8519);
    layer1_outputs(9148) <= not((layer0_outputs(12282)) or (layer0_outputs(9237)));
    layer1_outputs(9149) <= not(layer0_outputs(2916));
    layer1_outputs(9150) <= (layer0_outputs(11797)) and (layer0_outputs(854));
    layer1_outputs(9151) <= not(layer0_outputs(11995)) or (layer0_outputs(12130));
    layer1_outputs(9152) <= layer0_outputs(4250);
    layer1_outputs(9153) <= not((layer0_outputs(4943)) or (layer0_outputs(6067)));
    layer1_outputs(9154) <= not(layer0_outputs(4879));
    layer1_outputs(9155) <= not((layer0_outputs(8429)) or (layer0_outputs(4798)));
    layer1_outputs(9156) <= layer0_outputs(2156);
    layer1_outputs(9157) <= not(layer0_outputs(11691));
    layer1_outputs(9158) <= layer0_outputs(4594);
    layer1_outputs(9159) <= layer0_outputs(7765);
    layer1_outputs(9160) <= not((layer0_outputs(8059)) or (layer0_outputs(2057)));
    layer1_outputs(9161) <= not(layer0_outputs(4237));
    layer1_outputs(9162) <= layer0_outputs(4461);
    layer1_outputs(9163) <= layer0_outputs(12491);
    layer1_outputs(9164) <= not(layer0_outputs(4470)) or (layer0_outputs(12528));
    layer1_outputs(9165) <= not((layer0_outputs(1843)) or (layer0_outputs(1768)));
    layer1_outputs(9166) <= not(layer0_outputs(1776)) or (layer0_outputs(980));
    layer1_outputs(9167) <= (layer0_outputs(10396)) xor (layer0_outputs(7084));
    layer1_outputs(9168) <= not(layer0_outputs(10494));
    layer1_outputs(9169) <= not(layer0_outputs(7397)) or (layer0_outputs(8049));
    layer1_outputs(9170) <= '0';
    layer1_outputs(9171) <= (layer0_outputs(10282)) and (layer0_outputs(9670));
    layer1_outputs(9172) <= not((layer0_outputs(3309)) and (layer0_outputs(9406)));
    layer1_outputs(9173) <= '0';
    layer1_outputs(9174) <= not(layer0_outputs(8021)) or (layer0_outputs(7792));
    layer1_outputs(9175) <= not((layer0_outputs(4480)) xor (layer0_outputs(5574)));
    layer1_outputs(9176) <= not(layer0_outputs(3538));
    layer1_outputs(9177) <= not((layer0_outputs(11297)) xor (layer0_outputs(9005)));
    layer1_outputs(9178) <= not(layer0_outputs(3453));
    layer1_outputs(9179) <= not(layer0_outputs(9283));
    layer1_outputs(9180) <= not(layer0_outputs(12491)) or (layer0_outputs(9677));
    layer1_outputs(9181) <= layer0_outputs(8670);
    layer1_outputs(9182) <= layer0_outputs(1320);
    layer1_outputs(9183) <= not(layer0_outputs(6420));
    layer1_outputs(9184) <= (layer0_outputs(1306)) and (layer0_outputs(2610));
    layer1_outputs(9185) <= layer0_outputs(163);
    layer1_outputs(9186) <= not((layer0_outputs(6938)) or (layer0_outputs(6218)));
    layer1_outputs(9187) <= (layer0_outputs(9716)) or (layer0_outputs(857));
    layer1_outputs(9188) <= not(layer0_outputs(7030)) or (layer0_outputs(7909));
    layer1_outputs(9189) <= layer0_outputs(8233);
    layer1_outputs(9190) <= not(layer0_outputs(1971));
    layer1_outputs(9191) <= not(layer0_outputs(6862));
    layer1_outputs(9192) <= layer0_outputs(2760);
    layer1_outputs(9193) <= (layer0_outputs(827)) and not (layer0_outputs(987));
    layer1_outputs(9194) <= not((layer0_outputs(1270)) or (layer0_outputs(4295)));
    layer1_outputs(9195) <= (layer0_outputs(1056)) and not (layer0_outputs(6569));
    layer1_outputs(9196) <= '1';
    layer1_outputs(9197) <= (layer0_outputs(10722)) xor (layer0_outputs(6411));
    layer1_outputs(9198) <= layer0_outputs(12489);
    layer1_outputs(9199) <= (layer0_outputs(8153)) and not (layer0_outputs(11355));
    layer1_outputs(9200) <= (layer0_outputs(2483)) and not (layer0_outputs(1627));
    layer1_outputs(9201) <= layer0_outputs(1849);
    layer1_outputs(9202) <= not(layer0_outputs(6944));
    layer1_outputs(9203) <= layer0_outputs(8552);
    layer1_outputs(9204) <= layer0_outputs(11706);
    layer1_outputs(9205) <= layer0_outputs(2144);
    layer1_outputs(9206) <= not((layer0_outputs(8314)) or (layer0_outputs(9052)));
    layer1_outputs(9207) <= layer0_outputs(4528);
    layer1_outputs(9208) <= (layer0_outputs(4380)) and not (layer0_outputs(1885));
    layer1_outputs(9209) <= not(layer0_outputs(3951)) or (layer0_outputs(2758));
    layer1_outputs(9210) <= not(layer0_outputs(4078));
    layer1_outputs(9211) <= not(layer0_outputs(9288));
    layer1_outputs(9212) <= not(layer0_outputs(1863));
    layer1_outputs(9213) <= not((layer0_outputs(9449)) or (layer0_outputs(1979)));
    layer1_outputs(9214) <= not((layer0_outputs(9340)) xor (layer0_outputs(4144)));
    layer1_outputs(9215) <= not(layer0_outputs(8156)) or (layer0_outputs(3024));
    layer1_outputs(9216) <= (layer0_outputs(11890)) and not (layer0_outputs(11302));
    layer1_outputs(9217) <= (layer0_outputs(4894)) and (layer0_outputs(12307));
    layer1_outputs(9218) <= layer0_outputs(9831);
    layer1_outputs(9219) <= layer0_outputs(7775);
    layer1_outputs(9220) <= layer0_outputs(12772);
    layer1_outputs(9221) <= not(layer0_outputs(3392)) or (layer0_outputs(11903));
    layer1_outputs(9222) <= not(layer0_outputs(1987));
    layer1_outputs(9223) <= (layer0_outputs(3441)) or (layer0_outputs(109));
    layer1_outputs(9224) <= not(layer0_outputs(10388)) or (layer0_outputs(9472));
    layer1_outputs(9225) <= not(layer0_outputs(11306));
    layer1_outputs(9226) <= layer0_outputs(11871);
    layer1_outputs(9227) <= (layer0_outputs(12458)) and (layer0_outputs(1213));
    layer1_outputs(9228) <= (layer0_outputs(5052)) and not (layer0_outputs(10884));
    layer1_outputs(9229) <= (layer0_outputs(7712)) and not (layer0_outputs(9814));
    layer1_outputs(9230) <= not((layer0_outputs(9317)) or (layer0_outputs(146)));
    layer1_outputs(9231) <= layer0_outputs(6207);
    layer1_outputs(9232) <= not(layer0_outputs(7922)) or (layer0_outputs(4365));
    layer1_outputs(9233) <= (layer0_outputs(485)) or (layer0_outputs(2971));
    layer1_outputs(9234) <= (layer0_outputs(10106)) or (layer0_outputs(619));
    layer1_outputs(9235) <= layer0_outputs(10459);
    layer1_outputs(9236) <= not((layer0_outputs(7945)) and (layer0_outputs(11071)));
    layer1_outputs(9237) <= (layer0_outputs(8341)) xor (layer0_outputs(3520));
    layer1_outputs(9238) <= (layer0_outputs(3123)) and (layer0_outputs(8982));
    layer1_outputs(9239) <= layer0_outputs(10619);
    layer1_outputs(9240) <= (layer0_outputs(8745)) or (layer0_outputs(93));
    layer1_outputs(9241) <= not(layer0_outputs(8077));
    layer1_outputs(9242) <= layer0_outputs(1738);
    layer1_outputs(9243) <= not(layer0_outputs(6598));
    layer1_outputs(9244) <= (layer0_outputs(1325)) or (layer0_outputs(9680));
    layer1_outputs(9245) <= not((layer0_outputs(9411)) or (layer0_outputs(8872)));
    layer1_outputs(9246) <= layer0_outputs(8690);
    layer1_outputs(9247) <= not((layer0_outputs(336)) or (layer0_outputs(11639)));
    layer1_outputs(9248) <= layer0_outputs(930);
    layer1_outputs(9249) <= not(layer0_outputs(6294)) or (layer0_outputs(7400));
    layer1_outputs(9250) <= not((layer0_outputs(7100)) xor (layer0_outputs(8425)));
    layer1_outputs(9251) <= not(layer0_outputs(9985));
    layer1_outputs(9252) <= layer0_outputs(8588);
    layer1_outputs(9253) <= not(layer0_outputs(3130));
    layer1_outputs(9254) <= (layer0_outputs(4309)) xor (layer0_outputs(11899));
    layer1_outputs(9255) <= not(layer0_outputs(8607));
    layer1_outputs(9256) <= not((layer0_outputs(6620)) or (layer0_outputs(4814)));
    layer1_outputs(9257) <= layer0_outputs(4297);
    layer1_outputs(9258) <= not((layer0_outputs(4344)) xor (layer0_outputs(12175)));
    layer1_outputs(9259) <= not(layer0_outputs(1945));
    layer1_outputs(9260) <= (layer0_outputs(4652)) and not (layer0_outputs(5078));
    layer1_outputs(9261) <= not(layer0_outputs(3138));
    layer1_outputs(9262) <= (layer0_outputs(4069)) xor (layer0_outputs(11562));
    layer1_outputs(9263) <= not((layer0_outputs(5068)) and (layer0_outputs(6931)));
    layer1_outputs(9264) <= not(layer0_outputs(4241));
    layer1_outputs(9265) <= (layer0_outputs(11202)) or (layer0_outputs(409));
    layer1_outputs(9266) <= not(layer0_outputs(4480));
    layer1_outputs(9267) <= layer0_outputs(8303);
    layer1_outputs(9268) <= not(layer0_outputs(205)) or (layer0_outputs(9063));
    layer1_outputs(9269) <= (layer0_outputs(9995)) and not (layer0_outputs(7854));
    layer1_outputs(9270) <= not(layer0_outputs(73)) or (layer0_outputs(48));
    layer1_outputs(9271) <= not(layer0_outputs(852));
    layer1_outputs(9272) <= layer0_outputs(6264);
    layer1_outputs(9273) <= not(layer0_outputs(9702)) or (layer0_outputs(3292));
    layer1_outputs(9274) <= layer0_outputs(1621);
    layer1_outputs(9275) <= (layer0_outputs(8767)) or (layer0_outputs(3175));
    layer1_outputs(9276) <= not((layer0_outputs(10730)) xor (layer0_outputs(6715)));
    layer1_outputs(9277) <= layer0_outputs(11068);
    layer1_outputs(9278) <= not(layer0_outputs(487));
    layer1_outputs(9279) <= layer0_outputs(12610);
    layer1_outputs(9280) <= not(layer0_outputs(6332));
    layer1_outputs(9281) <= not(layer0_outputs(997)) or (layer0_outputs(12710));
    layer1_outputs(9282) <= (layer0_outputs(2432)) and (layer0_outputs(5322));
    layer1_outputs(9283) <= not((layer0_outputs(12664)) xor (layer0_outputs(181)));
    layer1_outputs(9284) <= not(layer0_outputs(7871)) or (layer0_outputs(5918));
    layer1_outputs(9285) <= (layer0_outputs(9309)) and (layer0_outputs(143));
    layer1_outputs(9286) <= layer0_outputs(12701);
    layer1_outputs(9287) <= not(layer0_outputs(630));
    layer1_outputs(9288) <= not((layer0_outputs(10963)) xor (layer0_outputs(10230)));
    layer1_outputs(9289) <= not(layer0_outputs(2573));
    layer1_outputs(9290) <= not(layer0_outputs(6516));
    layer1_outputs(9291) <= layer0_outputs(7672);
    layer1_outputs(9292) <= not(layer0_outputs(3855));
    layer1_outputs(9293) <= '1';
    layer1_outputs(9294) <= (layer0_outputs(10176)) and (layer0_outputs(2988));
    layer1_outputs(9295) <= (layer0_outputs(7938)) xor (layer0_outputs(11765));
    layer1_outputs(9296) <= not(layer0_outputs(11025));
    layer1_outputs(9297) <= not(layer0_outputs(8191)) or (layer0_outputs(6013));
    layer1_outputs(9298) <= (layer0_outputs(4612)) xor (layer0_outputs(224));
    layer1_outputs(9299) <= (layer0_outputs(186)) and not (layer0_outputs(5954));
    layer1_outputs(9300) <= (layer0_outputs(3355)) xor (layer0_outputs(10269));
    layer1_outputs(9301) <= not(layer0_outputs(3417));
    layer1_outputs(9302) <= not(layer0_outputs(8206));
    layer1_outputs(9303) <= not(layer0_outputs(9091)) or (layer0_outputs(353));
    layer1_outputs(9304) <= not(layer0_outputs(5786));
    layer1_outputs(9305) <= (layer0_outputs(6428)) and not (layer0_outputs(6416));
    layer1_outputs(9306) <= (layer0_outputs(3514)) and (layer0_outputs(10892));
    layer1_outputs(9307) <= layer0_outputs(11128);
    layer1_outputs(9308) <= layer0_outputs(9000);
    layer1_outputs(9309) <= not(layer0_outputs(10557));
    layer1_outputs(9310) <= not(layer0_outputs(12510));
    layer1_outputs(9311) <= not((layer0_outputs(4559)) or (layer0_outputs(8981)));
    layer1_outputs(9312) <= not(layer0_outputs(2873));
    layer1_outputs(9313) <= layer0_outputs(10522);
    layer1_outputs(9314) <= not(layer0_outputs(7520));
    layer1_outputs(9315) <= not(layer0_outputs(6704));
    layer1_outputs(9316) <= (layer0_outputs(1471)) and not (layer0_outputs(434));
    layer1_outputs(9317) <= not(layer0_outputs(4397)) or (layer0_outputs(4506));
    layer1_outputs(9318) <= (layer0_outputs(10341)) and not (layer0_outputs(1493));
    layer1_outputs(9319) <= (layer0_outputs(8591)) or (layer0_outputs(5124));
    layer1_outputs(9320) <= (layer0_outputs(8911)) and (layer0_outputs(821));
    layer1_outputs(9321) <= not(layer0_outputs(11541)) or (layer0_outputs(10756));
    layer1_outputs(9322) <= (layer0_outputs(11895)) or (layer0_outputs(11013));
    layer1_outputs(9323) <= '1';
    layer1_outputs(9324) <= layer0_outputs(2941);
    layer1_outputs(9325) <= '0';
    layer1_outputs(9326) <= (layer0_outputs(6564)) and (layer0_outputs(5841));
    layer1_outputs(9327) <= (layer0_outputs(8023)) xor (layer0_outputs(1312));
    layer1_outputs(9328) <= layer0_outputs(12496);
    layer1_outputs(9329) <= not(layer0_outputs(7383));
    layer1_outputs(9330) <= not(layer0_outputs(10426));
    layer1_outputs(9331) <= (layer0_outputs(526)) or (layer0_outputs(6125));
    layer1_outputs(9332) <= not((layer0_outputs(7751)) and (layer0_outputs(3118)));
    layer1_outputs(9333) <= (layer0_outputs(4083)) and not (layer0_outputs(8685));
    layer1_outputs(9334) <= layer0_outputs(12);
    layer1_outputs(9335) <= (layer0_outputs(2043)) and not (layer0_outputs(8198));
    layer1_outputs(9336) <= (layer0_outputs(2538)) and (layer0_outputs(9679));
    layer1_outputs(9337) <= not(layer0_outputs(3261)) or (layer0_outputs(12393));
    layer1_outputs(9338) <= layer0_outputs(2325);
    layer1_outputs(9339) <= not(layer0_outputs(856)) or (layer0_outputs(12756));
    layer1_outputs(9340) <= not(layer0_outputs(8996));
    layer1_outputs(9341) <= not((layer0_outputs(3183)) xor (layer0_outputs(4649)));
    layer1_outputs(9342) <= not(layer0_outputs(2484));
    layer1_outputs(9343) <= not(layer0_outputs(243)) or (layer0_outputs(1456));
    layer1_outputs(9344) <= (layer0_outputs(5220)) xor (layer0_outputs(9092));
    layer1_outputs(9345) <= (layer0_outputs(6170)) and not (layer0_outputs(3483));
    layer1_outputs(9346) <= (layer0_outputs(6669)) and (layer0_outputs(8842));
    layer1_outputs(9347) <= not(layer0_outputs(12093));
    layer1_outputs(9348) <= layer0_outputs(7968);
    layer1_outputs(9349) <= not(layer0_outputs(2436));
    layer1_outputs(9350) <= layer0_outputs(11787);
    layer1_outputs(9351) <= not(layer0_outputs(11573));
    layer1_outputs(9352) <= '1';
    layer1_outputs(9353) <= (layer0_outputs(6936)) or (layer0_outputs(377));
    layer1_outputs(9354) <= not(layer0_outputs(3699)) or (layer0_outputs(8411));
    layer1_outputs(9355) <= (layer0_outputs(3981)) xor (layer0_outputs(1884));
    layer1_outputs(9356) <= not((layer0_outputs(10128)) and (layer0_outputs(12349)));
    layer1_outputs(9357) <= layer0_outputs(3193);
    layer1_outputs(9358) <= layer0_outputs(5819);
    layer1_outputs(9359) <= not((layer0_outputs(8903)) and (layer0_outputs(2264)));
    layer1_outputs(9360) <= (layer0_outputs(10851)) and not (layer0_outputs(8475));
    layer1_outputs(9361) <= not(layer0_outputs(10656)) or (layer0_outputs(6692));
    layer1_outputs(9362) <= layer0_outputs(12760);
    layer1_outputs(9363) <= (layer0_outputs(11276)) and not (layer0_outputs(4002));
    layer1_outputs(9364) <= (layer0_outputs(3720)) or (layer0_outputs(11050));
    layer1_outputs(9365) <= not(layer0_outputs(118)) or (layer0_outputs(2430));
    layer1_outputs(9366) <= (layer0_outputs(6680)) and (layer0_outputs(10641));
    layer1_outputs(9367) <= layer0_outputs(5896);
    layer1_outputs(9368) <= not(layer0_outputs(11822));
    layer1_outputs(9369) <= not((layer0_outputs(10208)) and (layer0_outputs(2222)));
    layer1_outputs(9370) <= (layer0_outputs(3125)) and not (layer0_outputs(2494));
    layer1_outputs(9371) <= not(layer0_outputs(8561)) or (layer0_outputs(4887));
    layer1_outputs(9372) <= not(layer0_outputs(8322));
    layer1_outputs(9373) <= not(layer0_outputs(2772)) or (layer0_outputs(2343));
    layer1_outputs(9374) <= (layer0_outputs(10446)) and (layer0_outputs(11763));
    layer1_outputs(9375) <= layer0_outputs(874);
    layer1_outputs(9376) <= '1';
    layer1_outputs(9377) <= not(layer0_outputs(8968));
    layer1_outputs(9378) <= not((layer0_outputs(7781)) xor (layer0_outputs(1584)));
    layer1_outputs(9379) <= layer0_outputs(932);
    layer1_outputs(9380) <= (layer0_outputs(11976)) or (layer0_outputs(6465));
    layer1_outputs(9381) <= layer0_outputs(6144);
    layer1_outputs(9382) <= (layer0_outputs(6164)) and (layer0_outputs(8446));
    layer1_outputs(9383) <= not(layer0_outputs(1429));
    layer1_outputs(9384) <= not((layer0_outputs(7500)) xor (layer0_outputs(155)));
    layer1_outputs(9385) <= not(layer0_outputs(4394)) or (layer0_outputs(12106));
    layer1_outputs(9386) <= not((layer0_outputs(5402)) or (layer0_outputs(3015)));
    layer1_outputs(9387) <= (layer0_outputs(10248)) and (layer0_outputs(4876));
    layer1_outputs(9388) <= (layer0_outputs(912)) and (layer0_outputs(8481));
    layer1_outputs(9389) <= not((layer0_outputs(7246)) and (layer0_outputs(6904)));
    layer1_outputs(9390) <= (layer0_outputs(2246)) and (layer0_outputs(4491));
    layer1_outputs(9391) <= layer0_outputs(9966);
    layer1_outputs(9392) <= (layer0_outputs(9081)) or (layer0_outputs(7595));
    layer1_outputs(9393) <= layer0_outputs(6799);
    layer1_outputs(9394) <= layer0_outputs(190);
    layer1_outputs(9395) <= not(layer0_outputs(9349));
    layer1_outputs(9396) <= not(layer0_outputs(7604)) or (layer0_outputs(8172));
    layer1_outputs(9397) <= (layer0_outputs(10597)) or (layer0_outputs(7059));
    layer1_outputs(9398) <= not((layer0_outputs(8347)) and (layer0_outputs(272)));
    layer1_outputs(9399) <= not(layer0_outputs(9649)) or (layer0_outputs(9449));
    layer1_outputs(9400) <= layer0_outputs(8913);
    layer1_outputs(9401) <= (layer0_outputs(7823)) and (layer0_outputs(9156));
    layer1_outputs(9402) <= (layer0_outputs(6022)) or (layer0_outputs(4240));
    layer1_outputs(9403) <= layer0_outputs(6427);
    layer1_outputs(9404) <= layer0_outputs(8307);
    layer1_outputs(9405) <= (layer0_outputs(5997)) and not (layer0_outputs(9108));
    layer1_outputs(9406) <= (layer0_outputs(23)) and not (layer0_outputs(11400));
    layer1_outputs(9407) <= layer0_outputs(5466);
    layer1_outputs(9408) <= not(layer0_outputs(4086));
    layer1_outputs(9409) <= layer0_outputs(8843);
    layer1_outputs(9410) <= not((layer0_outputs(11849)) and (layer0_outputs(2016)));
    layer1_outputs(9411) <= (layer0_outputs(10059)) or (layer0_outputs(2648));
    layer1_outputs(9412) <= not(layer0_outputs(1267));
    layer1_outputs(9413) <= not((layer0_outputs(3698)) or (layer0_outputs(3774)));
    layer1_outputs(9414) <= (layer0_outputs(2079)) and (layer0_outputs(1234));
    layer1_outputs(9415) <= '1';
    layer1_outputs(9416) <= '1';
    layer1_outputs(9417) <= layer0_outputs(981);
    layer1_outputs(9418) <= not(layer0_outputs(5986));
    layer1_outputs(9419) <= (layer0_outputs(7392)) and not (layer0_outputs(5579));
    layer1_outputs(9420) <= layer0_outputs(10456);
    layer1_outputs(9421) <= not(layer0_outputs(3659)) or (layer0_outputs(3636));
    layer1_outputs(9422) <= not((layer0_outputs(8787)) or (layer0_outputs(2109)));
    layer1_outputs(9423) <= (layer0_outputs(12081)) and not (layer0_outputs(1620));
    layer1_outputs(9424) <= (layer0_outputs(8679)) or (layer0_outputs(6804));
    layer1_outputs(9425) <= not(layer0_outputs(4361));
    layer1_outputs(9426) <= (layer0_outputs(10465)) and (layer0_outputs(10120));
    layer1_outputs(9427) <= (layer0_outputs(4330)) or (layer0_outputs(596));
    layer1_outputs(9428) <= (layer0_outputs(2668)) xor (layer0_outputs(12314));
    layer1_outputs(9429) <= not(layer0_outputs(869)) or (layer0_outputs(1940));
    layer1_outputs(9430) <= not((layer0_outputs(11813)) or (layer0_outputs(6082)));
    layer1_outputs(9431) <= not(layer0_outputs(925));
    layer1_outputs(9432) <= layer0_outputs(10961);
    layer1_outputs(9433) <= not(layer0_outputs(9702));
    layer1_outputs(9434) <= not(layer0_outputs(682));
    layer1_outputs(9435) <= '1';
    layer1_outputs(9436) <= (layer0_outputs(11536)) and (layer0_outputs(3661));
    layer1_outputs(9437) <= not(layer0_outputs(6726));
    layer1_outputs(9438) <= not((layer0_outputs(12785)) xor (layer0_outputs(12786)));
    layer1_outputs(9439) <= layer0_outputs(5426);
    layer1_outputs(9440) <= (layer0_outputs(1483)) and not (layer0_outputs(9202));
    layer1_outputs(9441) <= layer0_outputs(7885);
    layer1_outputs(9442) <= not(layer0_outputs(5625));
    layer1_outputs(9443) <= layer0_outputs(2492);
    layer1_outputs(9444) <= not(layer0_outputs(3698));
    layer1_outputs(9445) <= not(layer0_outputs(12720)) or (layer0_outputs(8224));
    layer1_outputs(9446) <= not(layer0_outputs(7687)) or (layer0_outputs(1067));
    layer1_outputs(9447) <= layer0_outputs(4939);
    layer1_outputs(9448) <= (layer0_outputs(4323)) and not (layer0_outputs(2924));
    layer1_outputs(9449) <= not((layer0_outputs(11082)) and (layer0_outputs(12520)));
    layer1_outputs(9450) <= (layer0_outputs(8460)) and not (layer0_outputs(4149));
    layer1_outputs(9451) <= layer0_outputs(6168);
    layer1_outputs(9452) <= (layer0_outputs(544)) or (layer0_outputs(3544));
    layer1_outputs(9453) <= (layer0_outputs(388)) and (layer0_outputs(435));
    layer1_outputs(9454) <= not(layer0_outputs(9416)) or (layer0_outputs(8600));
    layer1_outputs(9455) <= not(layer0_outputs(977));
    layer1_outputs(9456) <= (layer0_outputs(1981)) or (layer0_outputs(3930));
    layer1_outputs(9457) <= not((layer0_outputs(3609)) xor (layer0_outputs(2537)));
    layer1_outputs(9458) <= not(layer0_outputs(6151)) or (layer0_outputs(1239));
    layer1_outputs(9459) <= not((layer0_outputs(11020)) xor (layer0_outputs(8982)));
    layer1_outputs(9460) <= (layer0_outputs(5165)) and not (layer0_outputs(1294));
    layer1_outputs(9461) <= (layer0_outputs(10651)) and (layer0_outputs(3080));
    layer1_outputs(9462) <= not((layer0_outputs(6367)) and (layer0_outputs(8480)));
    layer1_outputs(9463) <= (layer0_outputs(3481)) xor (layer0_outputs(6894));
    layer1_outputs(9464) <= not(layer0_outputs(4736)) or (layer0_outputs(8313));
    layer1_outputs(9465) <= '0';
    layer1_outputs(9466) <= not(layer0_outputs(9428));
    layer1_outputs(9467) <= (layer0_outputs(6004)) or (layer0_outputs(1377));
    layer1_outputs(9468) <= not(layer0_outputs(8799));
    layer1_outputs(9469) <= (layer0_outputs(11123)) and not (layer0_outputs(3425));
    layer1_outputs(9470) <= (layer0_outputs(11735)) and (layer0_outputs(410));
    layer1_outputs(9471) <= layer0_outputs(7731);
    layer1_outputs(9472) <= not(layer0_outputs(3916)) or (layer0_outputs(1317));
    layer1_outputs(9473) <= layer0_outputs(11047);
    layer1_outputs(9474) <= not(layer0_outputs(8464)) or (layer0_outputs(8463));
    layer1_outputs(9475) <= not(layer0_outputs(12148));
    layer1_outputs(9476) <= not(layer0_outputs(2655)) or (layer0_outputs(12171));
    layer1_outputs(9477) <= (layer0_outputs(4589)) xor (layer0_outputs(3202));
    layer1_outputs(9478) <= not(layer0_outputs(10197)) or (layer0_outputs(8256));
    layer1_outputs(9479) <= layer0_outputs(3798);
    layer1_outputs(9480) <= (layer0_outputs(2407)) and not (layer0_outputs(8441));
    layer1_outputs(9481) <= layer0_outputs(10899);
    layer1_outputs(9482) <= not(layer0_outputs(5734)) or (layer0_outputs(10312));
    layer1_outputs(9483) <= '1';
    layer1_outputs(9484) <= not(layer0_outputs(1784)) or (layer0_outputs(9555));
    layer1_outputs(9485) <= not(layer0_outputs(9132));
    layer1_outputs(9486) <= not(layer0_outputs(2874)) or (layer0_outputs(8186));
    layer1_outputs(9487) <= not((layer0_outputs(5756)) xor (layer0_outputs(10905)));
    layer1_outputs(9488) <= layer0_outputs(3092);
    layer1_outputs(9489) <= (layer0_outputs(2455)) and not (layer0_outputs(8715));
    layer1_outputs(9490) <= not(layer0_outputs(6495));
    layer1_outputs(9491) <= layer0_outputs(10608);
    layer1_outputs(9492) <= not(layer0_outputs(2143));
    layer1_outputs(9493) <= not(layer0_outputs(3359)) or (layer0_outputs(5432));
    layer1_outputs(9494) <= not((layer0_outputs(1216)) or (layer0_outputs(4303)));
    layer1_outputs(9495) <= not((layer0_outputs(8655)) and (layer0_outputs(2552)));
    layer1_outputs(9496) <= (layer0_outputs(8791)) or (layer0_outputs(11756));
    layer1_outputs(9497) <= not((layer0_outputs(3405)) or (layer0_outputs(11764)));
    layer1_outputs(9498) <= not(layer0_outputs(7670));
    layer1_outputs(9499) <= (layer0_outputs(6510)) and not (layer0_outputs(1965));
    layer1_outputs(9500) <= layer0_outputs(5489);
    layer1_outputs(9501) <= (layer0_outputs(9572)) and not (layer0_outputs(6388));
    layer1_outputs(9502) <= not(layer0_outputs(10086));
    layer1_outputs(9503) <= not(layer0_outputs(9403));
    layer1_outputs(9504) <= not(layer0_outputs(10481));
    layer1_outputs(9505) <= not((layer0_outputs(6866)) or (layer0_outputs(4376)));
    layer1_outputs(9506) <= not((layer0_outputs(1356)) or (layer0_outputs(9487)));
    layer1_outputs(9507) <= '0';
    layer1_outputs(9508) <= not(layer0_outputs(4390));
    layer1_outputs(9509) <= (layer0_outputs(1524)) or (layer0_outputs(9514));
    layer1_outputs(9510) <= not(layer0_outputs(7329)) or (layer0_outputs(4524));
    layer1_outputs(9511) <= layer0_outputs(3912);
    layer1_outputs(9512) <= (layer0_outputs(10828)) and not (layer0_outputs(6973));
    layer1_outputs(9513) <= (layer0_outputs(563)) xor (layer0_outputs(5053));
    layer1_outputs(9514) <= not((layer0_outputs(6356)) and (layer0_outputs(3376)));
    layer1_outputs(9515) <= not((layer0_outputs(1949)) and (layer0_outputs(1810)));
    layer1_outputs(9516) <= (layer0_outputs(4284)) xor (layer0_outputs(7046));
    layer1_outputs(9517) <= not(layer0_outputs(11951));
    layer1_outputs(9518) <= (layer0_outputs(3615)) or (layer0_outputs(3503));
    layer1_outputs(9519) <= not((layer0_outputs(923)) or (layer0_outputs(109)));
    layer1_outputs(9520) <= (layer0_outputs(3928)) or (layer0_outputs(9379));
    layer1_outputs(9521) <= '0';
    layer1_outputs(9522) <= '1';
    layer1_outputs(9523) <= not((layer0_outputs(1926)) or (layer0_outputs(11606)));
    layer1_outputs(9524) <= (layer0_outputs(2085)) xor (layer0_outputs(6163));
    layer1_outputs(9525) <= not(layer0_outputs(5459)) or (layer0_outputs(10789));
    layer1_outputs(9526) <= (layer0_outputs(3596)) and not (layer0_outputs(5254));
    layer1_outputs(9527) <= layer0_outputs(3122);
    layer1_outputs(9528) <= layer0_outputs(2917);
    layer1_outputs(9529) <= (layer0_outputs(8560)) and not (layer0_outputs(2155));
    layer1_outputs(9530) <= (layer0_outputs(7417)) and not (layer0_outputs(9980));
    layer1_outputs(9531) <= not((layer0_outputs(10068)) xor (layer0_outputs(2093)));
    layer1_outputs(9532) <= layer0_outputs(12753);
    layer1_outputs(9533) <= (layer0_outputs(1282)) and not (layer0_outputs(6034));
    layer1_outputs(9534) <= not((layer0_outputs(7239)) and (layer0_outputs(37)));
    layer1_outputs(9535) <= not((layer0_outputs(8240)) and (layer0_outputs(5335)));
    layer1_outputs(9536) <= not(layer0_outputs(8054));
    layer1_outputs(9537) <= not(layer0_outputs(11356));
    layer1_outputs(9538) <= (layer0_outputs(11195)) and not (layer0_outputs(12478));
    layer1_outputs(9539) <= not(layer0_outputs(6329));
    layer1_outputs(9540) <= not((layer0_outputs(11288)) xor (layer0_outputs(4997)));
    layer1_outputs(9541) <= (layer0_outputs(1467)) and not (layer0_outputs(3640));
    layer1_outputs(9542) <= not(layer0_outputs(6790)) or (layer0_outputs(504));
    layer1_outputs(9543) <= not((layer0_outputs(10035)) and (layer0_outputs(5974)));
    layer1_outputs(9544) <= (layer0_outputs(5614)) or (layer0_outputs(6901));
    layer1_outputs(9545) <= not((layer0_outputs(7752)) xor (layer0_outputs(8811)));
    layer1_outputs(9546) <= (layer0_outputs(4871)) and not (layer0_outputs(10095));
    layer1_outputs(9547) <= layer0_outputs(6443);
    layer1_outputs(9548) <= layer0_outputs(2058);
    layer1_outputs(9549) <= (layer0_outputs(8096)) and (layer0_outputs(3521));
    layer1_outputs(9550) <= not((layer0_outputs(5645)) xor (layer0_outputs(542)));
    layer1_outputs(9551) <= (layer0_outputs(5530)) and not (layer0_outputs(4763));
    layer1_outputs(9552) <= (layer0_outputs(5649)) and not (layer0_outputs(1435));
    layer1_outputs(9553) <= not((layer0_outputs(7470)) and (layer0_outputs(6427)));
    layer1_outputs(9554) <= '0';
    layer1_outputs(9555) <= not((layer0_outputs(8413)) xor (layer0_outputs(11726)));
    layer1_outputs(9556) <= not(layer0_outputs(9339)) or (layer0_outputs(3076));
    layer1_outputs(9557) <= (layer0_outputs(7778)) and not (layer0_outputs(7297));
    layer1_outputs(9558) <= layer0_outputs(6330);
    layer1_outputs(9559) <= (layer0_outputs(9192)) and not (layer0_outputs(5691));
    layer1_outputs(9560) <= not((layer0_outputs(1580)) or (layer0_outputs(9720)));
    layer1_outputs(9561) <= (layer0_outputs(4517)) and not (layer0_outputs(12698));
    layer1_outputs(9562) <= not((layer0_outputs(5722)) or (layer0_outputs(6860)));
    layer1_outputs(9563) <= not((layer0_outputs(4483)) or (layer0_outputs(3745)));
    layer1_outputs(9564) <= (layer0_outputs(2184)) and (layer0_outputs(4016));
    layer1_outputs(9565) <= not(layer0_outputs(8929)) or (layer0_outputs(4911));
    layer1_outputs(9566) <= (layer0_outputs(8489)) and not (layer0_outputs(11075));
    layer1_outputs(9567) <= not(layer0_outputs(11469)) or (layer0_outputs(5168));
    layer1_outputs(9568) <= not(layer0_outputs(12555)) or (layer0_outputs(4432));
    layer1_outputs(9569) <= not(layer0_outputs(2782)) or (layer0_outputs(1388));
    layer1_outputs(9570) <= not((layer0_outputs(12502)) or (layer0_outputs(12530)));
    layer1_outputs(9571) <= (layer0_outputs(783)) xor (layer0_outputs(1092));
    layer1_outputs(9572) <= not((layer0_outputs(10947)) or (layer0_outputs(3995)));
    layer1_outputs(9573) <= layer0_outputs(9387);
    layer1_outputs(9574) <= (layer0_outputs(8470)) and (layer0_outputs(4963));
    layer1_outputs(9575) <= not(layer0_outputs(68)) or (layer0_outputs(451));
    layer1_outputs(9576) <= (layer0_outputs(5869)) and not (layer0_outputs(10021));
    layer1_outputs(9577) <= layer0_outputs(9675);
    layer1_outputs(9578) <= not(layer0_outputs(3269)) or (layer0_outputs(2716));
    layer1_outputs(9579) <= not(layer0_outputs(10779));
    layer1_outputs(9580) <= layer0_outputs(2857);
    layer1_outputs(9581) <= not(layer0_outputs(4104));
    layer1_outputs(9582) <= (layer0_outputs(521)) xor (layer0_outputs(7172));
    layer1_outputs(9583) <= (layer0_outputs(696)) and (layer0_outputs(10188));
    layer1_outputs(9584) <= not(layer0_outputs(7438)) or (layer0_outputs(2025));
    layer1_outputs(9585) <= not(layer0_outputs(3605)) or (layer0_outputs(3365));
    layer1_outputs(9586) <= (layer0_outputs(8997)) xor (layer0_outputs(10071));
    layer1_outputs(9587) <= '0';
    layer1_outputs(9588) <= not((layer0_outputs(7428)) or (layer0_outputs(649)));
    layer1_outputs(9589) <= layer0_outputs(5413);
    layer1_outputs(9590) <= not(layer0_outputs(8683)) or (layer0_outputs(4011));
    layer1_outputs(9591) <= not((layer0_outputs(3784)) or (layer0_outputs(9671)));
    layer1_outputs(9592) <= not(layer0_outputs(1457));
    layer1_outputs(9593) <= '1';
    layer1_outputs(9594) <= (layer0_outputs(8672)) xor (layer0_outputs(8108));
    layer1_outputs(9595) <= layer0_outputs(3424);
    layer1_outputs(9596) <= not((layer0_outputs(1550)) and (layer0_outputs(1780)));
    layer1_outputs(9597) <= not(layer0_outputs(12583));
    layer1_outputs(9598) <= layer0_outputs(10007);
    layer1_outputs(9599) <= (layer0_outputs(1276)) xor (layer0_outputs(11328));
    layer1_outputs(9600) <= not(layer0_outputs(4489));
    layer1_outputs(9601) <= (layer0_outputs(1399)) xor (layer0_outputs(5882));
    layer1_outputs(9602) <= (layer0_outputs(3403)) and (layer0_outputs(3778));
    layer1_outputs(9603) <= not((layer0_outputs(7906)) or (layer0_outputs(3885)));
    layer1_outputs(9604) <= (layer0_outputs(7829)) xor (layer0_outputs(3120));
    layer1_outputs(9605) <= (layer0_outputs(9951)) and (layer0_outputs(11926));
    layer1_outputs(9606) <= layer0_outputs(3708);
    layer1_outputs(9607) <= not((layer0_outputs(8129)) and (layer0_outputs(3653)));
    layer1_outputs(9608) <= not(layer0_outputs(8549));
    layer1_outputs(9609) <= not(layer0_outputs(2490));
    layer1_outputs(9610) <= layer0_outputs(2203);
    layer1_outputs(9611) <= not(layer0_outputs(10345));
    layer1_outputs(9612) <= not(layer0_outputs(534)) or (layer0_outputs(11402));
    layer1_outputs(9613) <= layer0_outputs(10786);
    layer1_outputs(9614) <= (layer0_outputs(909)) xor (layer0_outputs(4903));
    layer1_outputs(9615) <= not(layer0_outputs(2746));
    layer1_outputs(9616) <= (layer0_outputs(7703)) and not (layer0_outputs(7488));
    layer1_outputs(9617) <= not(layer0_outputs(7074));
    layer1_outputs(9618) <= layer0_outputs(1389);
    layer1_outputs(9619) <= layer0_outputs(3881);
    layer1_outputs(9620) <= (layer0_outputs(10023)) and not (layer0_outputs(3421));
    layer1_outputs(9621) <= (layer0_outputs(2656)) and not (layer0_outputs(11065));
    layer1_outputs(9622) <= (layer0_outputs(10525)) and not (layer0_outputs(2485));
    layer1_outputs(9623) <= (layer0_outputs(5143)) and not (layer0_outputs(9150));
    layer1_outputs(9624) <= not((layer0_outputs(430)) or (layer0_outputs(8681)));
    layer1_outputs(9625) <= layer0_outputs(2341);
    layer1_outputs(9626) <= not((layer0_outputs(8897)) or (layer0_outputs(11142)));
    layer1_outputs(9627) <= layer0_outputs(2222);
    layer1_outputs(9628) <= not((layer0_outputs(8181)) or (layer0_outputs(11805)));
    layer1_outputs(9629) <= (layer0_outputs(7180)) or (layer0_outputs(1179));
    layer1_outputs(9630) <= layer0_outputs(2327);
    layer1_outputs(9631) <= layer0_outputs(4916);
    layer1_outputs(9632) <= not((layer0_outputs(4221)) or (layer0_outputs(7122)));
    layer1_outputs(9633) <= not(layer0_outputs(5661));
    layer1_outputs(9634) <= (layer0_outputs(11204)) and not (layer0_outputs(6894));
    layer1_outputs(9635) <= layer0_outputs(3256);
    layer1_outputs(9636) <= not(layer0_outputs(12176));
    layer1_outputs(9637) <= not(layer0_outputs(838));
    layer1_outputs(9638) <= not(layer0_outputs(5624));
    layer1_outputs(9639) <= not(layer0_outputs(8097)) or (layer0_outputs(5379));
    layer1_outputs(9640) <= layer0_outputs(6261);
    layer1_outputs(9641) <= layer0_outputs(7648);
    layer1_outputs(9642) <= not((layer0_outputs(3408)) or (layer0_outputs(5347)));
    layer1_outputs(9643) <= not(layer0_outputs(2687)) or (layer0_outputs(4907));
    layer1_outputs(9644) <= not(layer0_outputs(10757));
    layer1_outputs(9645) <= not((layer0_outputs(1712)) or (layer0_outputs(10444)));
    layer1_outputs(9646) <= (layer0_outputs(1693)) and not (layer0_outputs(6021));
    layer1_outputs(9647) <= (layer0_outputs(10895)) and not (layer0_outputs(3572));
    layer1_outputs(9648) <= layer0_outputs(221);
    layer1_outputs(9649) <= not(layer0_outputs(2645));
    layer1_outputs(9650) <= not((layer0_outputs(3274)) or (layer0_outputs(2767)));
    layer1_outputs(9651) <= (layer0_outputs(3005)) xor (layer0_outputs(8024));
    layer1_outputs(9652) <= (layer0_outputs(12788)) and (layer0_outputs(6086));
    layer1_outputs(9653) <= (layer0_outputs(12134)) and not (layer0_outputs(2136));
    layer1_outputs(9654) <= not(layer0_outputs(2370));
    layer1_outputs(9655) <= (layer0_outputs(12034)) and not (layer0_outputs(12700));
    layer1_outputs(9656) <= layer0_outputs(5435);
    layer1_outputs(9657) <= not(layer0_outputs(3461)) or (layer0_outputs(11496));
    layer1_outputs(9658) <= (layer0_outputs(2177)) and not (layer0_outputs(10695));
    layer1_outputs(9659) <= not((layer0_outputs(11733)) xor (layer0_outputs(6340)));
    layer1_outputs(9660) <= not(layer0_outputs(2976)) or (layer0_outputs(4962));
    layer1_outputs(9661) <= (layer0_outputs(8258)) xor (layer0_outputs(2820));
    layer1_outputs(9662) <= not(layer0_outputs(7734));
    layer1_outputs(9663) <= (layer0_outputs(668)) and not (layer0_outputs(3535));
    layer1_outputs(9664) <= not((layer0_outputs(9336)) xor (layer0_outputs(5325)));
    layer1_outputs(9665) <= not(layer0_outputs(11310)) or (layer0_outputs(11376));
    layer1_outputs(9666) <= (layer0_outputs(5417)) and not (layer0_outputs(10574));
    layer1_outputs(9667) <= not(layer0_outputs(247)) or (layer0_outputs(1046));
    layer1_outputs(9668) <= '1';
    layer1_outputs(9669) <= layer0_outputs(11865);
    layer1_outputs(9670) <= layer0_outputs(2123);
    layer1_outputs(9671) <= not((layer0_outputs(5194)) xor (layer0_outputs(10450)));
    layer1_outputs(9672) <= not(layer0_outputs(1615)) or (layer0_outputs(9553));
    layer1_outputs(9673) <= (layer0_outputs(9214)) and not (layer0_outputs(11794));
    layer1_outputs(9674) <= layer0_outputs(7318);
    layer1_outputs(9675) <= (layer0_outputs(0)) and not (layer0_outputs(10486));
    layer1_outputs(9676) <= layer0_outputs(10602);
    layer1_outputs(9677) <= not((layer0_outputs(3734)) or (layer0_outputs(8087)));
    layer1_outputs(9678) <= not((layer0_outputs(2560)) or (layer0_outputs(4179)));
    layer1_outputs(9679) <= (layer0_outputs(5111)) or (layer0_outputs(8079));
    layer1_outputs(9680) <= (layer0_outputs(5341)) and (layer0_outputs(5364));
    layer1_outputs(9681) <= not(layer0_outputs(6642));
    layer1_outputs(9682) <= not(layer0_outputs(8012));
    layer1_outputs(9683) <= not((layer0_outputs(3340)) xor (layer0_outputs(7820)));
    layer1_outputs(9684) <= (layer0_outputs(11468)) and not (layer0_outputs(7137));
    layer1_outputs(9685) <= not(layer0_outputs(9071)) or (layer0_outputs(8350));
    layer1_outputs(9686) <= not(layer0_outputs(7900));
    layer1_outputs(9687) <= not(layer0_outputs(8395)) or (layer0_outputs(10480));
    layer1_outputs(9688) <= not(layer0_outputs(7888));
    layer1_outputs(9689) <= layer0_outputs(7447);
    layer1_outputs(9690) <= not(layer0_outputs(3367));
    layer1_outputs(9691) <= not(layer0_outputs(7350)) or (layer0_outputs(4541));
    layer1_outputs(9692) <= (layer0_outputs(726)) and not (layer0_outputs(8188));
    layer1_outputs(9693) <= (layer0_outputs(12354)) xor (layer0_outputs(115));
    layer1_outputs(9694) <= not((layer0_outputs(2029)) or (layer0_outputs(4304)));
    layer1_outputs(9695) <= layer0_outputs(7330);
    layer1_outputs(9696) <= not((layer0_outputs(2798)) and (layer0_outputs(5552)));
    layer1_outputs(9697) <= (layer0_outputs(7561)) and not (layer0_outputs(4257));
    layer1_outputs(9698) <= not(layer0_outputs(5904));
    layer1_outputs(9699) <= layer0_outputs(6852);
    layer1_outputs(9700) <= not(layer0_outputs(6935)) or (layer0_outputs(3207));
    layer1_outputs(9701) <= (layer0_outputs(623)) and not (layer0_outputs(6017));
    layer1_outputs(9702) <= not(layer0_outputs(9318));
    layer1_outputs(9703) <= not((layer0_outputs(4154)) xor (layer0_outputs(7116)));
    layer1_outputs(9704) <= (layer0_outputs(7496)) xor (layer0_outputs(2576));
    layer1_outputs(9705) <= (layer0_outputs(3833)) and not (layer0_outputs(6289));
    layer1_outputs(9706) <= layer0_outputs(6637);
    layer1_outputs(9707) <= (layer0_outputs(7847)) and not (layer0_outputs(7797));
    layer1_outputs(9708) <= not((layer0_outputs(9760)) and (layer0_outputs(9797)));
    layer1_outputs(9709) <= not((layer0_outputs(5866)) and (layer0_outputs(1487)));
    layer1_outputs(9710) <= (layer0_outputs(9317)) or (layer0_outputs(2026));
    layer1_outputs(9711) <= '1';
    layer1_outputs(9712) <= not(layer0_outputs(6161));
    layer1_outputs(9713) <= (layer0_outputs(10099)) and (layer0_outputs(11104));
    layer1_outputs(9714) <= not((layer0_outputs(7801)) xor (layer0_outputs(7777)));
    layer1_outputs(9715) <= not((layer0_outputs(8145)) xor (layer0_outputs(994)));
    layer1_outputs(9716) <= not(layer0_outputs(5888));
    layer1_outputs(9717) <= not((layer0_outputs(4048)) or (layer0_outputs(970)));
    layer1_outputs(9718) <= not(layer0_outputs(8379));
    layer1_outputs(9719) <= layer0_outputs(10517);
    layer1_outputs(9720) <= not(layer0_outputs(10506)) or (layer0_outputs(10295));
    layer1_outputs(9721) <= (layer0_outputs(10376)) and not (layer0_outputs(5142));
    layer1_outputs(9722) <= layer0_outputs(5290);
    layer1_outputs(9723) <= not(layer0_outputs(2935));
    layer1_outputs(9724) <= not(layer0_outputs(2327));
    layer1_outputs(9725) <= layer0_outputs(4375);
    layer1_outputs(9726) <= layer0_outputs(3508);
    layer1_outputs(9727) <= '1';
    layer1_outputs(9728) <= (layer0_outputs(7696)) and not (layer0_outputs(5112));
    layer1_outputs(9729) <= not((layer0_outputs(10094)) and (layer0_outputs(7014)));
    layer1_outputs(9730) <= not(layer0_outputs(774)) or (layer0_outputs(10399));
    layer1_outputs(9731) <= layer0_outputs(12730);
    layer1_outputs(9732) <= not(layer0_outputs(10390));
    layer1_outputs(9733) <= layer0_outputs(1663);
    layer1_outputs(9734) <= not(layer0_outputs(3038));
    layer1_outputs(9735) <= not((layer0_outputs(4272)) xor (layer0_outputs(4281)));
    layer1_outputs(9736) <= not(layer0_outputs(6005));
    layer1_outputs(9737) <= (layer0_outputs(202)) and (layer0_outputs(8793));
    layer1_outputs(9738) <= not(layer0_outputs(10392)) or (layer0_outputs(12392));
    layer1_outputs(9739) <= (layer0_outputs(197)) and not (layer0_outputs(4965));
    layer1_outputs(9740) <= layer0_outputs(4220);
    layer1_outputs(9741) <= (layer0_outputs(3271)) and (layer0_outputs(2125));
    layer1_outputs(9742) <= not(layer0_outputs(7923));
    layer1_outputs(9743) <= not(layer0_outputs(9865));
    layer1_outputs(9744) <= layer0_outputs(6181);
    layer1_outputs(9745) <= (layer0_outputs(9323)) and not (layer0_outputs(4922));
    layer1_outputs(9746) <= not((layer0_outputs(7021)) xor (layer0_outputs(7795)));
    layer1_outputs(9747) <= not(layer0_outputs(3844));
    layer1_outputs(9748) <= not(layer0_outputs(8893)) or (layer0_outputs(2208));
    layer1_outputs(9749) <= not((layer0_outputs(4812)) and (layer0_outputs(9977)));
    layer1_outputs(9750) <= layer0_outputs(11695);
    layer1_outputs(9751) <= layer0_outputs(1861);
    layer1_outputs(9752) <= (layer0_outputs(11490)) and (layer0_outputs(5085));
    layer1_outputs(9753) <= not(layer0_outputs(9930));
    layer1_outputs(9754) <= not(layer0_outputs(9698)) or (layer0_outputs(10011));
    layer1_outputs(9755) <= '1';
    layer1_outputs(9756) <= layer0_outputs(4228);
    layer1_outputs(9757) <= (layer0_outputs(5017)) and (layer0_outputs(7890));
    layer1_outputs(9758) <= not(layer0_outputs(5710));
    layer1_outputs(9759) <= layer0_outputs(4277);
    layer1_outputs(9760) <= not((layer0_outputs(9349)) xor (layer0_outputs(319)));
    layer1_outputs(9761) <= not(layer0_outputs(11911));
    layer1_outputs(9762) <= (layer0_outputs(4827)) xor (layer0_outputs(11007));
    layer1_outputs(9763) <= not(layer0_outputs(1363));
    layer1_outputs(9764) <= not(layer0_outputs(1291));
    layer1_outputs(9765) <= (layer0_outputs(12201)) or (layer0_outputs(3557));
    layer1_outputs(9766) <= (layer0_outputs(1906)) xor (layer0_outputs(7861));
    layer1_outputs(9767) <= not(layer0_outputs(6399)) or (layer0_outputs(5129));
    layer1_outputs(9768) <= (layer0_outputs(10162)) or (layer0_outputs(8465));
    layer1_outputs(9769) <= (layer0_outputs(2118)) and not (layer0_outputs(4750));
    layer1_outputs(9770) <= (layer0_outputs(8899)) and not (layer0_outputs(4627));
    layer1_outputs(9771) <= not(layer0_outputs(4912)) or (layer0_outputs(658));
    layer1_outputs(9772) <= not(layer0_outputs(8307));
    layer1_outputs(9773) <= layer0_outputs(6599);
    layer1_outputs(9774) <= not((layer0_outputs(11093)) or (layer0_outputs(1491)));
    layer1_outputs(9775) <= not(layer0_outputs(3857)) or (layer0_outputs(7645));
    layer1_outputs(9776) <= not(layer0_outputs(6196));
    layer1_outputs(9777) <= (layer0_outputs(11954)) or (layer0_outputs(4424));
    layer1_outputs(9778) <= not((layer0_outputs(10536)) and (layer0_outputs(8061)));
    layer1_outputs(9779) <= (layer0_outputs(1141)) or (layer0_outputs(4863));
    layer1_outputs(9780) <= not(layer0_outputs(12159));
    layer1_outputs(9781) <= not((layer0_outputs(1852)) and (layer0_outputs(7363)));
    layer1_outputs(9782) <= layer0_outputs(2302);
    layer1_outputs(9783) <= layer0_outputs(10983);
    layer1_outputs(9784) <= layer0_outputs(11018);
    layer1_outputs(9785) <= (layer0_outputs(1577)) and (layer0_outputs(1369));
    layer1_outputs(9786) <= not((layer0_outputs(2773)) xor (layer0_outputs(10898)));
    layer1_outputs(9787) <= not(layer0_outputs(6627));
    layer1_outputs(9788) <= (layer0_outputs(8255)) xor (layer0_outputs(2274));
    layer1_outputs(9789) <= '0';
    layer1_outputs(9790) <= layer0_outputs(5383);
    layer1_outputs(9791) <= not(layer0_outputs(4697)) or (layer0_outputs(8506));
    layer1_outputs(9792) <= layer0_outputs(10148);
    layer1_outputs(9793) <= layer0_outputs(4473);
    layer1_outputs(9794) <= (layer0_outputs(1032)) and not (layer0_outputs(8952));
    layer1_outputs(9795) <= layer0_outputs(10780);
    layer1_outputs(9796) <= (layer0_outputs(2044)) and (layer0_outputs(892));
    layer1_outputs(9797) <= layer0_outputs(2794);
    layer1_outputs(9798) <= not(layer0_outputs(10090));
    layer1_outputs(9799) <= not((layer0_outputs(10099)) or (layer0_outputs(12238)));
    layer1_outputs(9800) <= (layer0_outputs(10942)) and (layer0_outputs(6099));
    layer1_outputs(9801) <= not(layer0_outputs(10387)) or (layer0_outputs(10018));
    layer1_outputs(9802) <= not(layer0_outputs(12487));
    layer1_outputs(9803) <= layer0_outputs(6768);
    layer1_outputs(9804) <= (layer0_outputs(2159)) and not (layer0_outputs(5686));
    layer1_outputs(9805) <= (layer0_outputs(2564)) and not (layer0_outputs(9056));
    layer1_outputs(9806) <= (layer0_outputs(946)) and not (layer0_outputs(4170));
    layer1_outputs(9807) <= layer0_outputs(1187);
    layer1_outputs(9808) <= not((layer0_outputs(6180)) or (layer0_outputs(2975)));
    layer1_outputs(9809) <= not((layer0_outputs(2847)) and (layer0_outputs(105)));
    layer1_outputs(9810) <= (layer0_outputs(11582)) and (layer0_outputs(1168));
    layer1_outputs(9811) <= (layer0_outputs(454)) and (layer0_outputs(5892));
    layer1_outputs(9812) <= not(layer0_outputs(621));
    layer1_outputs(9813) <= not(layer0_outputs(12335));
    layer1_outputs(9814) <= not(layer0_outputs(8185));
    layer1_outputs(9815) <= not(layer0_outputs(6403)) or (layer0_outputs(8061));
    layer1_outputs(9816) <= not((layer0_outputs(755)) and (layer0_outputs(10368)));
    layer1_outputs(9817) <= not(layer0_outputs(10180));
    layer1_outputs(9818) <= not(layer0_outputs(3397));
    layer1_outputs(9819) <= layer0_outputs(12729);
    layer1_outputs(9820) <= not(layer0_outputs(9039)) or (layer0_outputs(3294));
    layer1_outputs(9821) <= layer0_outputs(11560);
    layer1_outputs(9822) <= layer0_outputs(788);
    layer1_outputs(9823) <= not(layer0_outputs(3085)) or (layer0_outputs(1854));
    layer1_outputs(9824) <= not(layer0_outputs(6754)) or (layer0_outputs(2183));
    layer1_outputs(9825) <= layer0_outputs(11355);
    layer1_outputs(9826) <= not(layer0_outputs(4199));
    layer1_outputs(9827) <= not((layer0_outputs(5039)) xor (layer0_outputs(3527)));
    layer1_outputs(9828) <= not((layer0_outputs(7422)) xor (layer0_outputs(7463)));
    layer1_outputs(9829) <= layer0_outputs(9904);
    layer1_outputs(9830) <= not(layer0_outputs(6042));
    layer1_outputs(9831) <= (layer0_outputs(3298)) and not (layer0_outputs(12367));
    layer1_outputs(9832) <= layer0_outputs(10424);
    layer1_outputs(9833) <= (layer0_outputs(10813)) and (layer0_outputs(7742));
    layer1_outputs(9834) <= layer0_outputs(9843);
    layer1_outputs(9835) <= layer0_outputs(7725);
    layer1_outputs(9836) <= not((layer0_outputs(5720)) xor (layer0_outputs(7320)));
    layer1_outputs(9837) <= layer0_outputs(9784);
    layer1_outputs(9838) <= (layer0_outputs(9468)) and not (layer0_outputs(8363));
    layer1_outputs(9839) <= (layer0_outputs(9973)) and not (layer0_outputs(4589));
    layer1_outputs(9840) <= not(layer0_outputs(9359));
    layer1_outputs(9841) <= not(layer0_outputs(6503)) or (layer0_outputs(9393));
    layer1_outputs(9842) <= (layer0_outputs(1668)) xor (layer0_outputs(11312));
    layer1_outputs(9843) <= layer0_outputs(7365);
    layer1_outputs(9844) <= layer0_outputs(6247);
    layer1_outputs(9845) <= not(layer0_outputs(2934));
    layer1_outputs(9846) <= not(layer0_outputs(2723)) or (layer0_outputs(7169));
    layer1_outputs(9847) <= layer0_outputs(11980);
    layer1_outputs(9848) <= not((layer0_outputs(11672)) and (layer0_outputs(1936)));
    layer1_outputs(9849) <= layer0_outputs(10498);
    layer1_outputs(9850) <= not(layer0_outputs(1383)) or (layer0_outputs(3499));
    layer1_outputs(9851) <= not(layer0_outputs(14));
    layer1_outputs(9852) <= '0';
    layer1_outputs(9853) <= not((layer0_outputs(12511)) xor (layer0_outputs(1256)));
    layer1_outputs(9854) <= '0';
    layer1_outputs(9855) <= layer0_outputs(8280);
    layer1_outputs(9856) <= layer0_outputs(3146);
    layer1_outputs(9857) <= '0';
    layer1_outputs(9858) <= not(layer0_outputs(7258));
    layer1_outputs(9859) <= (layer0_outputs(4383)) and not (layer0_outputs(278));
    layer1_outputs(9860) <= not((layer0_outputs(9585)) or (layer0_outputs(7942)));
    layer1_outputs(9861) <= layer0_outputs(3801);
    layer1_outputs(9862) <= layer0_outputs(7110);
    layer1_outputs(9863) <= layer0_outputs(1974);
    layer1_outputs(9864) <= (layer0_outputs(5756)) or (layer0_outputs(3215));
    layer1_outputs(9865) <= not(layer0_outputs(8336));
    layer1_outputs(9866) <= (layer0_outputs(1731)) xor (layer0_outputs(1537));
    layer1_outputs(9867) <= (layer0_outputs(10154)) xor (layer0_outputs(8768));
    layer1_outputs(9868) <= not(layer0_outputs(11796)) or (layer0_outputs(1835));
    layer1_outputs(9869) <= layer0_outputs(954);
    layer1_outputs(9870) <= not(layer0_outputs(3092)) or (layer0_outputs(2809));
    layer1_outputs(9871) <= layer0_outputs(8838);
    layer1_outputs(9872) <= (layer0_outputs(7032)) and not (layer0_outputs(7457));
    layer1_outputs(9873) <= not(layer0_outputs(8882)) or (layer0_outputs(8427));
    layer1_outputs(9874) <= layer0_outputs(1548);
    layer1_outputs(9875) <= (layer0_outputs(12583)) and (layer0_outputs(829));
    layer1_outputs(9876) <= layer0_outputs(1653);
    layer1_outputs(9877) <= (layer0_outputs(2054)) and (layer0_outputs(4239));
    layer1_outputs(9878) <= not(layer0_outputs(10253));
    layer1_outputs(9879) <= layer0_outputs(1918);
    layer1_outputs(9880) <= layer0_outputs(2629);
    layer1_outputs(9881) <= layer0_outputs(11896);
    layer1_outputs(9882) <= layer0_outputs(4934);
    layer1_outputs(9883) <= not((layer0_outputs(3616)) or (layer0_outputs(88)));
    layer1_outputs(9884) <= (layer0_outputs(12088)) xor (layer0_outputs(10164));
    layer1_outputs(9885) <= (layer0_outputs(11660)) and not (layer0_outputs(6803));
    layer1_outputs(9886) <= not((layer0_outputs(2048)) or (layer0_outputs(7788)));
    layer1_outputs(9887) <= not(layer0_outputs(775));
    layer1_outputs(9888) <= not(layer0_outputs(11441));
    layer1_outputs(9889) <= not(layer0_outputs(4387));
    layer1_outputs(9890) <= layer0_outputs(7222);
    layer1_outputs(9891) <= (layer0_outputs(11116)) and not (layer0_outputs(2730));
    layer1_outputs(9892) <= not(layer0_outputs(4808));
    layer1_outputs(9893) <= (layer0_outputs(1257)) and not (layer0_outputs(9594));
    layer1_outputs(9894) <= not(layer0_outputs(4761)) or (layer0_outputs(8028));
    layer1_outputs(9895) <= layer0_outputs(4552);
    layer1_outputs(9896) <= layer0_outputs(3213);
    layer1_outputs(9897) <= not(layer0_outputs(11459));
    layer1_outputs(9898) <= not((layer0_outputs(1020)) or (layer0_outputs(5713)));
    layer1_outputs(9899) <= not((layer0_outputs(10662)) or (layer0_outputs(6997)));
    layer1_outputs(9900) <= layer0_outputs(866);
    layer1_outputs(9901) <= not(layer0_outputs(11618));
    layer1_outputs(9902) <= not(layer0_outputs(12390));
    layer1_outputs(9903) <= not((layer0_outputs(8298)) xor (layer0_outputs(11793)));
    layer1_outputs(9904) <= not((layer0_outputs(1471)) xor (layer0_outputs(11128)));
    layer1_outputs(9905) <= (layer0_outputs(3039)) and not (layer0_outputs(8417));
    layer1_outputs(9906) <= not(layer0_outputs(3029));
    layer1_outputs(9907) <= not(layer0_outputs(9242));
    layer1_outputs(9908) <= layer0_outputs(12698);
    layer1_outputs(9909) <= not(layer0_outputs(6833));
    layer1_outputs(9910) <= (layer0_outputs(1649)) and not (layer0_outputs(1423));
    layer1_outputs(9911) <= layer0_outputs(9137);
    layer1_outputs(9912) <= not(layer0_outputs(10010));
    layer1_outputs(9913) <= layer0_outputs(5169);
    layer1_outputs(9914) <= (layer0_outputs(7069)) and not (layer0_outputs(482));
    layer1_outputs(9915) <= '1';
    layer1_outputs(9916) <= (layer0_outputs(6326)) xor (layer0_outputs(3722));
    layer1_outputs(9917) <= layer0_outputs(2981);
    layer1_outputs(9918) <= not((layer0_outputs(11252)) or (layer0_outputs(1087)));
    layer1_outputs(9919) <= not((layer0_outputs(11176)) xor (layer0_outputs(10160)));
    layer1_outputs(9920) <= (layer0_outputs(6633)) and not (layer0_outputs(2558));
    layer1_outputs(9921) <= (layer0_outputs(2068)) and not (layer0_outputs(10797));
    layer1_outputs(9922) <= not(layer0_outputs(2161));
    layer1_outputs(9923) <= not(layer0_outputs(7598));
    layer1_outputs(9924) <= layer0_outputs(7379);
    layer1_outputs(9925) <= not(layer0_outputs(7693));
    layer1_outputs(9926) <= not(layer0_outputs(11846));
    layer1_outputs(9927) <= (layer0_outputs(10043)) and not (layer0_outputs(8872));
    layer1_outputs(9928) <= layer0_outputs(6240);
    layer1_outputs(9929) <= not(layer0_outputs(5301));
    layer1_outputs(9930) <= not(layer0_outputs(976)) or (layer0_outputs(8762));
    layer1_outputs(9931) <= not(layer0_outputs(3304));
    layer1_outputs(9932) <= '0';
    layer1_outputs(9933) <= (layer0_outputs(8173)) and (layer0_outputs(17));
    layer1_outputs(9934) <= (layer0_outputs(11463)) and (layer0_outputs(4965));
    layer1_outputs(9935) <= '0';
    layer1_outputs(9936) <= not(layer0_outputs(3254));
    layer1_outputs(9937) <= layer0_outputs(5465);
    layer1_outputs(9938) <= not(layer0_outputs(1133));
    layer1_outputs(9939) <= layer0_outputs(12307);
    layer1_outputs(9940) <= not(layer0_outputs(1817));
    layer1_outputs(9941) <= (layer0_outputs(1436)) and (layer0_outputs(12495));
    layer1_outputs(9942) <= not(layer0_outputs(4440)) or (layer0_outputs(10900));
    layer1_outputs(9943) <= not((layer0_outputs(3376)) xor (layer0_outputs(7415)));
    layer1_outputs(9944) <= layer0_outputs(12450);
    layer1_outputs(9945) <= not(layer0_outputs(10718)) or (layer0_outputs(12475));
    layer1_outputs(9946) <= not((layer0_outputs(1089)) or (layer0_outputs(3783)));
    layer1_outputs(9947) <= not((layer0_outputs(335)) xor (layer0_outputs(6385)));
    layer1_outputs(9948) <= layer0_outputs(6336);
    layer1_outputs(9949) <= not(layer0_outputs(6045)) or (layer0_outputs(4088));
    layer1_outputs(9950) <= layer0_outputs(341);
    layer1_outputs(9951) <= (layer0_outputs(5973)) and not (layer0_outputs(5901));
    layer1_outputs(9952) <= not(layer0_outputs(5494));
    layer1_outputs(9953) <= layer0_outputs(3227);
    layer1_outputs(9954) <= not(layer0_outputs(5262)) or (layer0_outputs(1942));
    layer1_outputs(9955) <= (layer0_outputs(8075)) and (layer0_outputs(8975));
    layer1_outputs(9956) <= layer0_outputs(11627);
    layer1_outputs(9957) <= (layer0_outputs(349)) and not (layer0_outputs(1391));
    layer1_outputs(9958) <= not(layer0_outputs(940));
    layer1_outputs(9959) <= (layer0_outputs(3089)) and (layer0_outputs(6423));
    layer1_outputs(9960) <= (layer0_outputs(6458)) xor (layer0_outputs(2407));
    layer1_outputs(9961) <= not((layer0_outputs(1379)) xor (layer0_outputs(7309)));
    layer1_outputs(9962) <= (layer0_outputs(3914)) xor (layer0_outputs(5110));
    layer1_outputs(9963) <= not(layer0_outputs(5862)) or (layer0_outputs(4768));
    layer1_outputs(9964) <= (layer0_outputs(8839)) and (layer0_outputs(1800));
    layer1_outputs(9965) <= (layer0_outputs(7062)) and (layer0_outputs(4933));
    layer1_outputs(9966) <= (layer0_outputs(12682)) xor (layer0_outputs(10000));
    layer1_outputs(9967) <= not((layer0_outputs(11018)) xor (layer0_outputs(4481)));
    layer1_outputs(9968) <= not((layer0_outputs(1290)) or (layer0_outputs(11748)));
    layer1_outputs(9969) <= not(layer0_outputs(848));
    layer1_outputs(9970) <= (layer0_outputs(7078)) and (layer0_outputs(9992));
    layer1_outputs(9971) <= (layer0_outputs(7109)) and not (layer0_outputs(10821));
    layer1_outputs(9972) <= layer0_outputs(5264);
    layer1_outputs(9973) <= (layer0_outputs(6208)) and not (layer0_outputs(4914));
    layer1_outputs(9974) <= not(layer0_outputs(2618));
    layer1_outputs(9975) <= (layer0_outputs(5986)) or (layer0_outputs(5816));
    layer1_outputs(9976) <= not(layer0_outputs(4708));
    layer1_outputs(9977) <= layer0_outputs(11386);
    layer1_outputs(9978) <= not(layer0_outputs(3140)) or (layer0_outputs(8272));
    layer1_outputs(9979) <= (layer0_outputs(4017)) and (layer0_outputs(6528));
    layer1_outputs(9980) <= not(layer0_outputs(1134));
    layer1_outputs(9981) <= not((layer0_outputs(3568)) xor (layer0_outputs(5502)));
    layer1_outputs(9982) <= layer0_outputs(9174);
    layer1_outputs(9983) <= (layer0_outputs(10869)) and not (layer0_outputs(4438));
    layer1_outputs(9984) <= not((layer0_outputs(7287)) or (layer0_outputs(6650)));
    layer1_outputs(9985) <= not((layer0_outputs(2081)) and (layer0_outputs(9753)));
    layer1_outputs(9986) <= not((layer0_outputs(12664)) and (layer0_outputs(10178)));
    layer1_outputs(9987) <= (layer0_outputs(12287)) and not (layer0_outputs(11225));
    layer1_outputs(9988) <= not(layer0_outputs(9552));
    layer1_outputs(9989) <= not((layer0_outputs(734)) xor (layer0_outputs(11546)));
    layer1_outputs(9990) <= (layer0_outputs(3260)) or (layer0_outputs(6123));
    layer1_outputs(9991) <= layer0_outputs(4306);
    layer1_outputs(9992) <= not(layer0_outputs(9741)) or (layer0_outputs(4219));
    layer1_outputs(9993) <= (layer0_outputs(5216)) or (layer0_outputs(9372));
    layer1_outputs(9994) <= layer0_outputs(2588);
    layer1_outputs(9995) <= not((layer0_outputs(6686)) and (layer0_outputs(6913)));
    layer1_outputs(9996) <= (layer0_outputs(12595)) and not (layer0_outputs(4448));
    layer1_outputs(9997) <= not(layer0_outputs(7892));
    layer1_outputs(9998) <= not(layer0_outputs(2237)) or (layer0_outputs(5414));
    layer1_outputs(9999) <= not(layer0_outputs(10657)) or (layer0_outputs(5448));
    layer1_outputs(10000) <= (layer0_outputs(1652)) and not (layer0_outputs(5875));
    layer1_outputs(10001) <= layer0_outputs(7726);
    layer1_outputs(10002) <= layer0_outputs(11667);
    layer1_outputs(10003) <= (layer0_outputs(5955)) and not (layer0_outputs(7505));
    layer1_outputs(10004) <= (layer0_outputs(9788)) and (layer0_outputs(11379));
    layer1_outputs(10005) <= not((layer0_outputs(7347)) and (layer0_outputs(1678)));
    layer1_outputs(10006) <= (layer0_outputs(10450)) or (layer0_outputs(2913));
    layer1_outputs(10007) <= not((layer0_outputs(9806)) or (layer0_outputs(5800)));
    layer1_outputs(10008) <= (layer0_outputs(11412)) or (layer0_outputs(7587));
    layer1_outputs(10009) <= not(layer0_outputs(365));
    layer1_outputs(10010) <= (layer0_outputs(7263)) xor (layer0_outputs(1537));
    layer1_outputs(10011) <= '1';
    layer1_outputs(10012) <= not(layer0_outputs(8860));
    layer1_outputs(10013) <= not((layer0_outputs(6342)) or (layer0_outputs(9230)));
    layer1_outputs(10014) <= layer0_outputs(12479);
    layer1_outputs(10015) <= not(layer0_outputs(9190));
    layer1_outputs(10016) <= not(layer0_outputs(4342));
    layer1_outputs(10017) <= layer0_outputs(4738);
    layer1_outputs(10018) <= (layer0_outputs(997)) or (layer0_outputs(809));
    layer1_outputs(10019) <= not(layer0_outputs(6901));
    layer1_outputs(10020) <= not(layer0_outputs(10896)) or (layer0_outputs(2278));
    layer1_outputs(10021) <= not(layer0_outputs(8456)) or (layer0_outputs(6687));
    layer1_outputs(10022) <= (layer0_outputs(8276)) and not (layer0_outputs(10830));
    layer1_outputs(10023) <= layer0_outputs(10846);
    layer1_outputs(10024) <= not(layer0_outputs(6621));
    layer1_outputs(10025) <= (layer0_outputs(4892)) and not (layer0_outputs(668));
    layer1_outputs(10026) <= not(layer0_outputs(7244)) or (layer0_outputs(12787));
    layer1_outputs(10027) <= layer0_outputs(7982);
    layer1_outputs(10028) <= layer0_outputs(12117);
    layer1_outputs(10029) <= layer0_outputs(1608);
    layer1_outputs(10030) <= (layer0_outputs(7056)) or (layer0_outputs(4058));
    layer1_outputs(10031) <= layer0_outputs(4519);
    layer1_outputs(10032) <= not(layer0_outputs(2108));
    layer1_outputs(10033) <= (layer0_outputs(3434)) and not (layer0_outputs(11154));
    layer1_outputs(10034) <= '1';
    layer1_outputs(10035) <= '1';
    layer1_outputs(10036) <= (layer0_outputs(4223)) or (layer0_outputs(11853));
    layer1_outputs(10037) <= not(layer0_outputs(8404));
    layer1_outputs(10038) <= layer0_outputs(2595);
    layer1_outputs(10039) <= not(layer0_outputs(11851));
    layer1_outputs(10040) <= not((layer0_outputs(12758)) or (layer0_outputs(12119)));
    layer1_outputs(10041) <= layer0_outputs(5063);
    layer1_outputs(10042) <= not(layer0_outputs(3357)) or (layer0_outputs(8311));
    layer1_outputs(10043) <= not((layer0_outputs(12161)) or (layer0_outputs(7112)));
    layer1_outputs(10044) <= '0';
    layer1_outputs(10045) <= not(layer0_outputs(7036));
    layer1_outputs(10046) <= not((layer0_outputs(676)) or (layer0_outputs(9102)));
    layer1_outputs(10047) <= not((layer0_outputs(8418)) xor (layer0_outputs(5880)));
    layer1_outputs(10048) <= not(layer0_outputs(9425)) or (layer0_outputs(5983));
    layer1_outputs(10049) <= layer0_outputs(433);
    layer1_outputs(10050) <= not(layer0_outputs(8889)) or (layer0_outputs(8778));
    layer1_outputs(10051) <= not((layer0_outputs(8182)) or (layer0_outputs(2567)));
    layer1_outputs(10052) <= not(layer0_outputs(9942));
    layer1_outputs(10053) <= not(layer0_outputs(778)) or (layer0_outputs(11662));
    layer1_outputs(10054) <= (layer0_outputs(3629)) and not (layer0_outputs(1155));
    layer1_outputs(10055) <= not(layer0_outputs(10589)) or (layer0_outputs(4013));
    layer1_outputs(10056) <= not(layer0_outputs(2423));
    layer1_outputs(10057) <= not(layer0_outputs(6945));
    layer1_outputs(10058) <= '0';
    layer1_outputs(10059) <= not(layer0_outputs(5855)) or (layer0_outputs(4757));
    layer1_outputs(10060) <= not(layer0_outputs(3573));
    layer1_outputs(10061) <= (layer0_outputs(5407)) xor (layer0_outputs(2199));
    layer1_outputs(10062) <= not((layer0_outputs(7553)) and (layer0_outputs(7252)));
    layer1_outputs(10063) <= not(layer0_outputs(6809));
    layer1_outputs(10064) <= not((layer0_outputs(8840)) or (layer0_outputs(3420)));
    layer1_outputs(10065) <= layer0_outputs(7009);
    layer1_outputs(10066) <= '0';
    layer1_outputs(10067) <= layer0_outputs(9347);
    layer1_outputs(10068) <= layer0_outputs(1434);
    layer1_outputs(10069) <= not(layer0_outputs(4717)) or (layer0_outputs(3541));
    layer1_outputs(10070) <= not((layer0_outputs(2191)) xor (layer0_outputs(1765)));
    layer1_outputs(10071) <= not(layer0_outputs(5047));
    layer1_outputs(10072) <= not((layer0_outputs(7875)) and (layer0_outputs(10170)));
    layer1_outputs(10073) <= (layer0_outputs(625)) xor (layer0_outputs(1485));
    layer1_outputs(10074) <= not((layer0_outputs(2245)) and (layer0_outputs(6291)));
    layer1_outputs(10075) <= not((layer0_outputs(9559)) or (layer0_outputs(4806)));
    layer1_outputs(10076) <= layer0_outputs(2391);
    layer1_outputs(10077) <= not((layer0_outputs(10159)) and (layer0_outputs(11812)));
    layer1_outputs(10078) <= (layer0_outputs(2607)) and not (layer0_outputs(7019));
    layer1_outputs(10079) <= layer0_outputs(3065);
    layer1_outputs(10080) <= not(layer0_outputs(5612)) or (layer0_outputs(7916));
    layer1_outputs(10081) <= (layer0_outputs(2364)) and (layer0_outputs(8240));
    layer1_outputs(10082) <= (layer0_outputs(7442)) and not (layer0_outputs(9351));
    layer1_outputs(10083) <= not(layer0_outputs(5131));
    layer1_outputs(10084) <= not(layer0_outputs(10075));
    layer1_outputs(10085) <= not(layer0_outputs(3753)) or (layer0_outputs(8768));
    layer1_outputs(10086) <= layer0_outputs(1906);
    layer1_outputs(10087) <= not(layer0_outputs(9074)) or (layer0_outputs(1303));
    layer1_outputs(10088) <= layer0_outputs(1128);
    layer1_outputs(10089) <= layer0_outputs(12485);
    layer1_outputs(10090) <= (layer0_outputs(12797)) and not (layer0_outputs(4722));
    layer1_outputs(10091) <= (layer0_outputs(4930)) and (layer0_outputs(4613));
    layer1_outputs(10092) <= (layer0_outputs(843)) and not (layer0_outputs(9494));
    layer1_outputs(10093) <= not((layer0_outputs(5559)) or (layer0_outputs(701)));
    layer1_outputs(10094) <= (layer0_outputs(5074)) xor (layer0_outputs(1097));
    layer1_outputs(10095) <= not(layer0_outputs(6698));
    layer1_outputs(10096) <= not((layer0_outputs(12512)) and (layer0_outputs(6248)));
    layer1_outputs(10097) <= not(layer0_outputs(2662)) or (layer0_outputs(11338));
    layer1_outputs(10098) <= not(layer0_outputs(12751));
    layer1_outputs(10099) <= (layer0_outputs(9138)) or (layer0_outputs(9158));
    layer1_outputs(10100) <= layer0_outputs(8545);
    layer1_outputs(10101) <= (layer0_outputs(3506)) and not (layer0_outputs(2724));
    layer1_outputs(10102) <= (layer0_outputs(9279)) and not (layer0_outputs(6653));
    layer1_outputs(10103) <= not((layer0_outputs(12618)) xor (layer0_outputs(5321)));
    layer1_outputs(10104) <= (layer0_outputs(1985)) and not (layer0_outputs(7175));
    layer1_outputs(10105) <= layer0_outputs(4372);
    layer1_outputs(10106) <= (layer0_outputs(1759)) and not (layer0_outputs(10316));
    layer1_outputs(10107) <= not((layer0_outputs(1578)) or (layer0_outputs(11945)));
    layer1_outputs(10108) <= not((layer0_outputs(7936)) xor (layer0_outputs(12533)));
    layer1_outputs(10109) <= not(layer0_outputs(10497));
    layer1_outputs(10110) <= not(layer0_outputs(9563)) or (layer0_outputs(182));
    layer1_outputs(10111) <= (layer0_outputs(7648)) xor (layer0_outputs(8477));
    layer1_outputs(10112) <= (layer0_outputs(11781)) and (layer0_outputs(1696));
    layer1_outputs(10113) <= not((layer0_outputs(10364)) and (layer0_outputs(11736)));
    layer1_outputs(10114) <= not(layer0_outputs(694));
    layer1_outputs(10115) <= not(layer0_outputs(59));
    layer1_outputs(10116) <= (layer0_outputs(167)) xor (layer0_outputs(9631));
    layer1_outputs(10117) <= not((layer0_outputs(1629)) or (layer0_outputs(7243)));
    layer1_outputs(10118) <= not(layer0_outputs(3710));
    layer1_outputs(10119) <= (layer0_outputs(148)) and not (layer0_outputs(6520));
    layer1_outputs(10120) <= not(layer0_outputs(7952));
    layer1_outputs(10121) <= not(layer0_outputs(1277));
    layer1_outputs(10122) <= '1';
    layer1_outputs(10123) <= not((layer0_outputs(10957)) xor (layer0_outputs(11170)));
    layer1_outputs(10124) <= layer0_outputs(2874);
    layer1_outputs(10125) <= layer0_outputs(6955);
    layer1_outputs(10126) <= not(layer0_outputs(6648));
    layer1_outputs(10127) <= (layer0_outputs(7704)) and not (layer0_outputs(1330));
    layer1_outputs(10128) <= not(layer0_outputs(12109)) or (layer0_outputs(9173));
    layer1_outputs(10129) <= not((layer0_outputs(8159)) or (layer0_outputs(8438)));
    layer1_outputs(10130) <= layer0_outputs(2168);
    layer1_outputs(10131) <= not((layer0_outputs(4171)) and (layer0_outputs(3623)));
    layer1_outputs(10132) <= not(layer0_outputs(11337));
    layer1_outputs(10133) <= not((layer0_outputs(9180)) or (layer0_outputs(9397)));
    layer1_outputs(10134) <= (layer0_outputs(7151)) and not (layer0_outputs(2457));
    layer1_outputs(10135) <= not((layer0_outputs(11605)) and (layer0_outputs(6865)));
    layer1_outputs(10136) <= not((layer0_outputs(10019)) and (layer0_outputs(5020)));
    layer1_outputs(10137) <= (layer0_outputs(5830)) and not (layer0_outputs(8035));
    layer1_outputs(10138) <= not(layer0_outputs(1782));
    layer1_outputs(10139) <= (layer0_outputs(11527)) and not (layer0_outputs(11720));
    layer1_outputs(10140) <= layer0_outputs(7487);
    layer1_outputs(10141) <= layer0_outputs(4958);
    layer1_outputs(10142) <= not((layer0_outputs(10001)) or (layer0_outputs(4983)));
    layer1_outputs(10143) <= not(layer0_outputs(3088));
    layer1_outputs(10144) <= not(layer0_outputs(3694));
    layer1_outputs(10145) <= layer0_outputs(6080);
    layer1_outputs(10146) <= layer0_outputs(4188);
    layer1_outputs(10147) <= (layer0_outputs(6094)) xor (layer0_outputs(4865));
    layer1_outputs(10148) <= not(layer0_outputs(6276));
    layer1_outputs(10149) <= not(layer0_outputs(4700));
    layer1_outputs(10150) <= not((layer0_outputs(1570)) and (layer0_outputs(11518)));
    layer1_outputs(10151) <= not(layer0_outputs(4781));
    layer1_outputs(10152) <= (layer0_outputs(7144)) xor (layer0_outputs(264));
    layer1_outputs(10153) <= (layer0_outputs(11203)) xor (layer0_outputs(2784));
    layer1_outputs(10154) <= not((layer0_outputs(603)) or (layer0_outputs(10616)));
    layer1_outputs(10155) <= not((layer0_outputs(582)) and (layer0_outputs(7560)));
    layer1_outputs(10156) <= layer0_outputs(4338);
    layer1_outputs(10157) <= not((layer0_outputs(12227)) xor (layer0_outputs(855)));
    layer1_outputs(10158) <= layer0_outputs(8964);
    layer1_outputs(10159) <= (layer0_outputs(5179)) xor (layer0_outputs(9790));
    layer1_outputs(10160) <= (layer0_outputs(2565)) or (layer0_outputs(6334));
    layer1_outputs(10161) <= not((layer0_outputs(6233)) xor (layer0_outputs(3556)));
    layer1_outputs(10162) <= not((layer0_outputs(11119)) and (layer0_outputs(2137)));
    layer1_outputs(10163) <= layer0_outputs(8155);
    layer1_outputs(10164) <= not(layer0_outputs(7887));
    layer1_outputs(10165) <= (layer0_outputs(6881)) and not (layer0_outputs(11968));
    layer1_outputs(10166) <= not(layer0_outputs(4460));
    layer1_outputs(10167) <= not(layer0_outputs(632));
    layer1_outputs(10168) <= layer0_outputs(11987);
    layer1_outputs(10169) <= not((layer0_outputs(4388)) and (layer0_outputs(3178)));
    layer1_outputs(10170) <= layer0_outputs(3278);
    layer1_outputs(10171) <= not(layer0_outputs(11802)) or (layer0_outputs(12377));
    layer1_outputs(10172) <= layer0_outputs(7556);
    layer1_outputs(10173) <= not((layer0_outputs(9506)) or (layer0_outputs(6073)));
    layer1_outputs(10174) <= layer0_outputs(11533);
    layer1_outputs(10175) <= (layer0_outputs(3565)) or (layer0_outputs(6072));
    layer1_outputs(10176) <= (layer0_outputs(6132)) or (layer0_outputs(1628));
    layer1_outputs(10177) <= layer0_outputs(4442);
    layer1_outputs(10178) <= not((layer0_outputs(6058)) and (layer0_outputs(7229)));
    layer1_outputs(10179) <= layer0_outputs(8859);
    layer1_outputs(10180) <= not((layer0_outputs(946)) and (layer0_outputs(7319)));
    layer1_outputs(10181) <= (layer0_outputs(11577)) and not (layer0_outputs(11491));
    layer1_outputs(10182) <= layer0_outputs(3412);
    layer1_outputs(10183) <= (layer0_outputs(12007)) and not (layer0_outputs(11369));
    layer1_outputs(10184) <= (layer0_outputs(412)) and (layer0_outputs(306));
    layer1_outputs(10185) <= not(layer0_outputs(8971)) or (layer0_outputs(4141));
    layer1_outputs(10186) <= (layer0_outputs(5404)) xor (layer0_outputs(10333));
    layer1_outputs(10187) <= not(layer0_outputs(2833));
    layer1_outputs(10188) <= layer0_outputs(6764);
    layer1_outputs(10189) <= (layer0_outputs(9093)) xor (layer0_outputs(702));
    layer1_outputs(10190) <= (layer0_outputs(11491)) or (layer0_outputs(7399));
    layer1_outputs(10191) <= (layer0_outputs(6109)) and not (layer0_outputs(7553));
    layer1_outputs(10192) <= not((layer0_outputs(42)) and (layer0_outputs(7060)));
    layer1_outputs(10193) <= not(layer0_outputs(6028)) or (layer0_outputs(12726));
    layer1_outputs(10194) <= not(layer0_outputs(156));
    layer1_outputs(10195) <= (layer0_outputs(7551)) and (layer0_outputs(9007));
    layer1_outputs(10196) <= layer0_outputs(4685);
    layer1_outputs(10197) <= not((layer0_outputs(4712)) and (layer0_outputs(1176)));
    layer1_outputs(10198) <= (layer0_outputs(11708)) or (layer0_outputs(2539));
    layer1_outputs(10199) <= not((layer0_outputs(2455)) xor (layer0_outputs(4977)));
    layer1_outputs(10200) <= not(layer0_outputs(6153));
    layer1_outputs(10201) <= layer0_outputs(7872);
    layer1_outputs(10202) <= (layer0_outputs(6022)) and (layer0_outputs(2763));
    layer1_outputs(10203) <= (layer0_outputs(126)) and not (layer0_outputs(9062));
    layer1_outputs(10204) <= (layer0_outputs(7291)) and not (layer0_outputs(692));
    layer1_outputs(10205) <= layer0_outputs(139);
    layer1_outputs(10206) <= layer0_outputs(2317);
    layer1_outputs(10207) <= not(layer0_outputs(5655));
    layer1_outputs(10208) <= layer0_outputs(10205);
    layer1_outputs(10209) <= '1';
    layer1_outputs(10210) <= not((layer0_outputs(6225)) or (layer0_outputs(4765)));
    layer1_outputs(10211) <= layer0_outputs(3726);
    layer1_outputs(10212) <= '1';
    layer1_outputs(10213) <= (layer0_outputs(10249)) and not (layer0_outputs(7550));
    layer1_outputs(10214) <= not(layer0_outputs(9722)) or (layer0_outputs(8008));
    layer1_outputs(10215) <= not(layer0_outputs(3824));
    layer1_outputs(10216) <= not(layer0_outputs(7602));
    layer1_outputs(10217) <= (layer0_outputs(5438)) and (layer0_outputs(11169));
    layer1_outputs(10218) <= not((layer0_outputs(687)) and (layer0_outputs(6386)));
    layer1_outputs(10219) <= not(layer0_outputs(7432));
    layer1_outputs(10220) <= layer0_outputs(12737);
    layer1_outputs(10221) <= (layer0_outputs(4361)) or (layer0_outputs(10857));
    layer1_outputs(10222) <= layer0_outputs(490);
    layer1_outputs(10223) <= not(layer0_outputs(2015));
    layer1_outputs(10224) <= (layer0_outputs(4228)) xor (layer0_outputs(3633));
    layer1_outputs(10225) <= (layer0_outputs(5985)) and not (layer0_outputs(500));
    layer1_outputs(10226) <= (layer0_outputs(2630)) and not (layer0_outputs(1130));
    layer1_outputs(10227) <= '0';
    layer1_outputs(10228) <= not(layer0_outputs(9865)) or (layer0_outputs(861));
    layer1_outputs(10229) <= (layer0_outputs(2853)) xor (layer0_outputs(8722));
    layer1_outputs(10230) <= not(layer0_outputs(7377)) or (layer0_outputs(7004));
    layer1_outputs(10231) <= (layer0_outputs(5126)) and not (layer0_outputs(10));
    layer1_outputs(10232) <= layer0_outputs(11657);
    layer1_outputs(10233) <= not(layer0_outputs(12582)) or (layer0_outputs(4696));
    layer1_outputs(10234) <= not((layer0_outputs(11675)) or (layer0_outputs(3600)));
    layer1_outputs(10235) <= not((layer0_outputs(6110)) xor (layer0_outputs(11454)));
    layer1_outputs(10236) <= (layer0_outputs(2905)) xor (layer0_outputs(4817));
    layer1_outputs(10237) <= not(layer0_outputs(11346));
    layer1_outputs(10238) <= layer0_outputs(1468);
    layer1_outputs(10239) <= not(layer0_outputs(9284));
    layer1_outputs(10240) <= (layer0_outputs(5781)) and not (layer0_outputs(11145));
    layer1_outputs(10241) <= layer0_outputs(12076);
    layer1_outputs(10242) <= not(layer0_outputs(3377));
    layer1_outputs(10243) <= not(layer0_outputs(1311)) or (layer0_outputs(5688));
    layer1_outputs(10244) <= (layer0_outputs(1362)) and (layer0_outputs(11784));
    layer1_outputs(10245) <= layer0_outputs(12327);
    layer1_outputs(10246) <= not((layer0_outputs(5414)) or (layer0_outputs(851)));
    layer1_outputs(10247) <= not((layer0_outputs(8006)) xor (layer0_outputs(3986)));
    layer1_outputs(10248) <= (layer0_outputs(1086)) and not (layer0_outputs(6372));
    layer1_outputs(10249) <= layer0_outputs(6266);
    layer1_outputs(10250) <= (layer0_outputs(6512)) xor (layer0_outputs(5957));
    layer1_outputs(10251) <= not(layer0_outputs(3550));
    layer1_outputs(10252) <= not((layer0_outputs(2411)) or (layer0_outputs(8619)));
    layer1_outputs(10253) <= not(layer0_outputs(6148));
    layer1_outputs(10254) <= not(layer0_outputs(7748));
    layer1_outputs(10255) <= not(layer0_outputs(10310)) or (layer0_outputs(9589));
    layer1_outputs(10256) <= not((layer0_outputs(4421)) or (layer0_outputs(1019)));
    layer1_outputs(10257) <= layer0_outputs(8712);
    layer1_outputs(10258) <= not(layer0_outputs(8574)) or (layer0_outputs(10935));
    layer1_outputs(10259) <= (layer0_outputs(3648)) and not (layer0_outputs(1934));
    layer1_outputs(10260) <= not(layer0_outputs(8554));
    layer1_outputs(10261) <= not(layer0_outputs(3655));
    layer1_outputs(10262) <= (layer0_outputs(9958)) and not (layer0_outputs(9528));
    layer1_outputs(10263) <= not(layer0_outputs(9496));
    layer1_outputs(10264) <= (layer0_outputs(10874)) and not (layer0_outputs(11687));
    layer1_outputs(10265) <= not(layer0_outputs(1011));
    layer1_outputs(10266) <= (layer0_outputs(10264)) and not (layer0_outputs(12369));
    layer1_outputs(10267) <= not(layer0_outputs(1693));
    layer1_outputs(10268) <= not((layer0_outputs(1837)) xor (layer0_outputs(10587)));
    layer1_outputs(10269) <= not(layer0_outputs(703));
    layer1_outputs(10270) <= (layer0_outputs(5747)) and (layer0_outputs(2515));
    layer1_outputs(10271) <= (layer0_outputs(348)) or (layer0_outputs(6644));
    layer1_outputs(10272) <= not(layer0_outputs(12252));
    layer1_outputs(10273) <= not((layer0_outputs(8103)) and (layer0_outputs(2938)));
    layer1_outputs(10274) <= not(layer0_outputs(10465)) or (layer0_outputs(12073));
    layer1_outputs(10275) <= not(layer0_outputs(4976)) or (layer0_outputs(4809));
    layer1_outputs(10276) <= '1';
    layer1_outputs(10277) <= (layer0_outputs(3871)) and not (layer0_outputs(9988));
    layer1_outputs(10278) <= (layer0_outputs(7141)) and not (layer0_outputs(5946));
    layer1_outputs(10279) <= not((layer0_outputs(2243)) xor (layer0_outputs(8749)));
    layer1_outputs(10280) <= not((layer0_outputs(10918)) and (layer0_outputs(11914)));
    layer1_outputs(10281) <= (layer0_outputs(3891)) xor (layer0_outputs(4227));
    layer1_outputs(10282) <= not((layer0_outputs(11233)) xor (layer0_outputs(2479)));
    layer1_outputs(10283) <= layer0_outputs(7301);
    layer1_outputs(10284) <= layer0_outputs(12551);
    layer1_outputs(10285) <= layer0_outputs(3920);
    layer1_outputs(10286) <= not((layer0_outputs(8819)) or (layer0_outputs(6008)));
    layer1_outputs(10287) <= (layer0_outputs(10626)) and not (layer0_outputs(8491));
    layer1_outputs(10288) <= not(layer0_outputs(6589));
    layer1_outputs(10289) <= not((layer0_outputs(5990)) and (layer0_outputs(12674)));
    layer1_outputs(10290) <= not((layer0_outputs(7359)) xor (layer0_outputs(7011)));
    layer1_outputs(10291) <= (layer0_outputs(10926)) and not (layer0_outputs(5189));
    layer1_outputs(10292) <= not(layer0_outputs(6555)) or (layer0_outputs(2286));
    layer1_outputs(10293) <= (layer0_outputs(9444)) xor (layer0_outputs(7361));
    layer1_outputs(10294) <= '1';
    layer1_outputs(10295) <= not((layer0_outputs(7751)) or (layer0_outputs(1932)));
    layer1_outputs(10296) <= not((layer0_outputs(2032)) and (layer0_outputs(3208)));
    layer1_outputs(10297) <= layer0_outputs(2167);
    layer1_outputs(10298) <= layer0_outputs(8055);
    layer1_outputs(10299) <= not(layer0_outputs(1607));
    layer1_outputs(10300) <= (layer0_outputs(4476)) and not (layer0_outputs(3027));
    layer1_outputs(10301) <= not(layer0_outputs(11235));
    layer1_outputs(10302) <= not((layer0_outputs(1813)) xor (layer0_outputs(8533)));
    layer1_outputs(10303) <= not(layer0_outputs(9337));
    layer1_outputs(10304) <= layer0_outputs(10502);
    layer1_outputs(10305) <= not((layer0_outputs(2389)) or (layer0_outputs(844)));
    layer1_outputs(10306) <= '0';
    layer1_outputs(10307) <= not(layer0_outputs(61));
    layer1_outputs(10308) <= not((layer0_outputs(4863)) and (layer0_outputs(2871)));
    layer1_outputs(10309) <= not(layer0_outputs(9367));
    layer1_outputs(10310) <= layer0_outputs(1646);
    layer1_outputs(10311) <= not((layer0_outputs(6814)) xor (layer0_outputs(10700)));
    layer1_outputs(10312) <= (layer0_outputs(10865)) and (layer0_outputs(196));
    layer1_outputs(10313) <= layer0_outputs(4737);
    layer1_outputs(10314) <= not(layer0_outputs(11928));
    layer1_outputs(10315) <= not(layer0_outputs(5319));
    layer1_outputs(10316) <= (layer0_outputs(6214)) or (layer0_outputs(462));
    layer1_outputs(10317) <= not(layer0_outputs(1331)) or (layer0_outputs(7875));
    layer1_outputs(10318) <= (layer0_outputs(658)) and not (layer0_outputs(7125));
    layer1_outputs(10319) <= (layer0_outputs(329)) xor (layer0_outputs(3453));
    layer1_outputs(10320) <= not(layer0_outputs(4730));
    layer1_outputs(10321) <= (layer0_outputs(12475)) and (layer0_outputs(11166));
    layer1_outputs(10322) <= layer0_outputs(10969);
    layer1_outputs(10323) <= not(layer0_outputs(788));
    layer1_outputs(10324) <= (layer0_outputs(4741)) and not (layer0_outputs(5750));
    layer1_outputs(10325) <= (layer0_outputs(12324)) and not (layer0_outputs(10739));
    layer1_outputs(10326) <= layer0_outputs(379);
    layer1_outputs(10327) <= layer0_outputs(7818);
    layer1_outputs(10328) <= (layer0_outputs(4142)) and not (layer0_outputs(6713));
    layer1_outputs(10329) <= (layer0_outputs(11503)) and (layer0_outputs(5206));
    layer1_outputs(10330) <= not(layer0_outputs(7346));
    layer1_outputs(10331) <= not(layer0_outputs(7961));
    layer1_outputs(10332) <= not((layer0_outputs(10653)) xor (layer0_outputs(11546)));
    layer1_outputs(10333) <= not((layer0_outputs(9072)) xor (layer0_outputs(639)));
    layer1_outputs(10334) <= not((layer0_outputs(9297)) xor (layer0_outputs(11213)));
    layer1_outputs(10335) <= not(layer0_outputs(3816)) or (layer0_outputs(12426));
    layer1_outputs(10336) <= layer0_outputs(8092);
    layer1_outputs(10337) <= (layer0_outputs(6811)) and not (layer0_outputs(1523));
    layer1_outputs(10338) <= (layer0_outputs(11405)) or (layer0_outputs(10308));
    layer1_outputs(10339) <= (layer0_outputs(285)) and not (layer0_outputs(5695));
    layer1_outputs(10340) <= layer0_outputs(7851);
    layer1_outputs(10341) <= not(layer0_outputs(1472)) or (layer0_outputs(1476));
    layer1_outputs(10342) <= layer0_outputs(3446);
    layer1_outputs(10343) <= (layer0_outputs(6465)) or (layer0_outputs(8378));
    layer1_outputs(10344) <= (layer0_outputs(1233)) and (layer0_outputs(8862));
    layer1_outputs(10345) <= not((layer0_outputs(674)) or (layer0_outputs(7948)));
    layer1_outputs(10346) <= not(layer0_outputs(10672));
    layer1_outputs(10347) <= (layer0_outputs(9746)) xor (layer0_outputs(2149));
    layer1_outputs(10348) <= layer0_outputs(7512);
    layer1_outputs(10349) <= not(layer0_outputs(12311)) or (layer0_outputs(3971));
    layer1_outputs(10350) <= (layer0_outputs(8218)) and not (layer0_outputs(3233));
    layer1_outputs(10351) <= not(layer0_outputs(6936));
    layer1_outputs(10352) <= not(layer0_outputs(10617));
    layer1_outputs(10353) <= (layer0_outputs(4375)) and not (layer0_outputs(8698));
    layer1_outputs(10354) <= not(layer0_outputs(12228)) or (layer0_outputs(7469));
    layer1_outputs(10355) <= layer0_outputs(729);
    layer1_outputs(10356) <= not(layer0_outputs(9492)) or (layer0_outputs(7247));
    layer1_outputs(10357) <= (layer0_outputs(1217)) xor (layer0_outputs(4604));
    layer1_outputs(10358) <= layer0_outputs(7472);
    layer1_outputs(10359) <= layer0_outputs(802);
    layer1_outputs(10360) <= not(layer0_outputs(2065)) or (layer0_outputs(3310));
    layer1_outputs(10361) <= (layer0_outputs(3929)) xor (layer0_outputs(2203));
    layer1_outputs(10362) <= layer0_outputs(9083);
    layer1_outputs(10363) <= (layer0_outputs(3959)) and (layer0_outputs(10725));
    layer1_outputs(10364) <= (layer0_outputs(11005)) and (layer0_outputs(180));
    layer1_outputs(10365) <= '0';
    layer1_outputs(10366) <= (layer0_outputs(2958)) and (layer0_outputs(2672));
    layer1_outputs(10367) <= layer0_outputs(4582);
    layer1_outputs(10368) <= (layer0_outputs(2725)) xor (layer0_outputs(10772));
    layer1_outputs(10369) <= not(layer0_outputs(5611)) or (layer0_outputs(7663));
    layer1_outputs(10370) <= not(layer0_outputs(6793));
    layer1_outputs(10371) <= layer0_outputs(9338);
    layer1_outputs(10372) <= not((layer0_outputs(187)) and (layer0_outputs(1170)));
    layer1_outputs(10373) <= layer0_outputs(10172);
    layer1_outputs(10374) <= '0';
    layer1_outputs(10375) <= (layer0_outputs(11586)) xor (layer0_outputs(263));
    layer1_outputs(10376) <= not(layer0_outputs(892)) or (layer0_outputs(1704));
    layer1_outputs(10377) <= (layer0_outputs(6625)) and not (layer0_outputs(9837));
    layer1_outputs(10378) <= not(layer0_outputs(10663));
    layer1_outputs(10379) <= layer0_outputs(1740);
    layer1_outputs(10380) <= not((layer0_outputs(6066)) or (layer0_outputs(7671)));
    layer1_outputs(10381) <= not(layer0_outputs(7111)) or (layer0_outputs(9217));
    layer1_outputs(10382) <= layer0_outputs(1757);
    layer1_outputs(10383) <= '0';
    layer1_outputs(10384) <= not(layer0_outputs(12384));
    layer1_outputs(10385) <= not(layer0_outputs(8960));
    layer1_outputs(10386) <= not((layer0_outputs(10051)) or (layer0_outputs(12783)));
    layer1_outputs(10387) <= layer0_outputs(685);
    layer1_outputs(10388) <= layer0_outputs(3384);
    layer1_outputs(10389) <= (layer0_outputs(10276)) and not (layer0_outputs(1853));
    layer1_outputs(10390) <= (layer0_outputs(1604)) and not (layer0_outputs(4498));
    layer1_outputs(10391) <= layer0_outputs(2283);
    layer1_outputs(10392) <= (layer0_outputs(6137)) or (layer0_outputs(631));
    layer1_outputs(10393) <= (layer0_outputs(7749)) xor (layer0_outputs(3710));
    layer1_outputs(10394) <= (layer0_outputs(1433)) and (layer0_outputs(3563));
    layer1_outputs(10395) <= not(layer0_outputs(576)) or (layer0_outputs(10678));
    layer1_outputs(10396) <= (layer0_outputs(4283)) xor (layer0_outputs(739));
    layer1_outputs(10397) <= (layer0_outputs(5867)) and not (layer0_outputs(4278));
    layer1_outputs(10398) <= (layer0_outputs(5246)) or (layer0_outputs(12681));
    layer1_outputs(10399) <= layer0_outputs(9820);
    layer1_outputs(10400) <= not(layer0_outputs(4977));
    layer1_outputs(10401) <= (layer0_outputs(10033)) and (layer0_outputs(12337));
    layer1_outputs(10402) <= not(layer0_outputs(9001)) or (layer0_outputs(7179));
    layer1_outputs(10403) <= not(layer0_outputs(2829)) or (layer0_outputs(12618));
    layer1_outputs(10404) <= not((layer0_outputs(11935)) xor (layer0_outputs(10541)));
    layer1_outputs(10405) <= (layer0_outputs(2741)) xor (layer0_outputs(10197));
    layer1_outputs(10406) <= (layer0_outputs(12279)) or (layer0_outputs(3522));
    layer1_outputs(10407) <= not(layer0_outputs(4466)) or (layer0_outputs(9750));
    layer1_outputs(10408) <= not(layer0_outputs(10297));
    layer1_outputs(10409) <= (layer0_outputs(4788)) or (layer0_outputs(10935));
    layer1_outputs(10410) <= not(layer0_outputs(4374));
    layer1_outputs(10411) <= (layer0_outputs(10328)) and not (layer0_outputs(6971));
    layer1_outputs(10412) <= not(layer0_outputs(11548));
    layer1_outputs(10413) <= not(layer0_outputs(6917)) or (layer0_outputs(7664));
    layer1_outputs(10414) <= not((layer0_outputs(11375)) and (layer0_outputs(3769)));
    layer1_outputs(10415) <= (layer0_outputs(6093)) and not (layer0_outputs(10637));
    layer1_outputs(10416) <= layer0_outputs(5346);
    layer1_outputs(10417) <= not((layer0_outputs(2258)) or (layer0_outputs(11337)));
    layer1_outputs(10418) <= (layer0_outputs(12581)) xor (layer0_outputs(12179));
    layer1_outputs(10419) <= not(layer0_outputs(3236)) or (layer0_outputs(5698));
    layer1_outputs(10420) <= (layer0_outputs(9673)) and not (layer0_outputs(3928));
    layer1_outputs(10421) <= layer0_outputs(3427);
    layer1_outputs(10422) <= (layer0_outputs(1487)) and not (layer0_outputs(12684));
    layer1_outputs(10423) <= not((layer0_outputs(3294)) or (layer0_outputs(1260)));
    layer1_outputs(10424) <= (layer0_outputs(5779)) xor (layer0_outputs(7023));
    layer1_outputs(10425) <= not(layer0_outputs(1155)) or (layer0_outputs(4546));
    layer1_outputs(10426) <= layer0_outputs(13);
    layer1_outputs(10427) <= not((layer0_outputs(4230)) or (layer0_outputs(7902)));
    layer1_outputs(10428) <= not(layer0_outputs(8175));
    layer1_outputs(10429) <= not(layer0_outputs(11004)) or (layer0_outputs(2791));
    layer1_outputs(10430) <= not(layer0_outputs(4758)) or (layer0_outputs(10070));
    layer1_outputs(10431) <= not(layer0_outputs(5160)) or (layer0_outputs(7509));
    layer1_outputs(10432) <= (layer0_outputs(3474)) or (layer0_outputs(3022));
    layer1_outputs(10433) <= layer0_outputs(11689);
    layer1_outputs(10434) <= not((layer0_outputs(8292)) or (layer0_outputs(11589)));
    layer1_outputs(10435) <= layer0_outputs(11406);
    layer1_outputs(10436) <= not(layer0_outputs(5764));
    layer1_outputs(10437) <= not(layer0_outputs(2974));
    layer1_outputs(10438) <= not(layer0_outputs(4940));
    layer1_outputs(10439) <= (layer0_outputs(10231)) or (layer0_outputs(7706));
    layer1_outputs(10440) <= not((layer0_outputs(12178)) or (layer0_outputs(9573)));
    layer1_outputs(10441) <= (layer0_outputs(4326)) and not (layer0_outputs(2413));
    layer1_outputs(10442) <= layer0_outputs(10216);
    layer1_outputs(10443) <= layer0_outputs(4561);
    layer1_outputs(10444) <= not(layer0_outputs(5178)) or (layer0_outputs(10184));
    layer1_outputs(10445) <= layer0_outputs(5022);
    layer1_outputs(10446) <= layer0_outputs(2994);
    layer1_outputs(10447) <= layer0_outputs(2887);
    layer1_outputs(10448) <= not((layer0_outputs(2342)) or (layer0_outputs(9010)));
    layer1_outputs(10449) <= not((layer0_outputs(5927)) or (layer0_outputs(5959)));
    layer1_outputs(10450) <= '0';
    layer1_outputs(10451) <= (layer0_outputs(6841)) and (layer0_outputs(4494));
    layer1_outputs(10452) <= not(layer0_outputs(231));
    layer1_outputs(10453) <= not(layer0_outputs(9840));
    layer1_outputs(10454) <= (layer0_outputs(10553)) and not (layer0_outputs(394));
    layer1_outputs(10455) <= not(layer0_outputs(1492)) or (layer0_outputs(3348));
    layer1_outputs(10456) <= layer0_outputs(6176);
    layer1_outputs(10457) <= not(layer0_outputs(10466)) or (layer0_outputs(2052));
    layer1_outputs(10458) <= (layer0_outputs(2876)) or (layer0_outputs(1710));
    layer1_outputs(10459) <= not(layer0_outputs(7319));
    layer1_outputs(10460) <= (layer0_outputs(12374)) and (layer0_outputs(1495));
    layer1_outputs(10461) <= (layer0_outputs(6912)) and not (layer0_outputs(4877));
    layer1_outputs(10462) <= not(layer0_outputs(6299));
    layer1_outputs(10463) <= layer0_outputs(8063);
    layer1_outputs(10464) <= (layer0_outputs(9265)) xor (layer0_outputs(9320));
    layer1_outputs(10465) <= not((layer0_outputs(8833)) and (layer0_outputs(4253)));
    layer1_outputs(10466) <= (layer0_outputs(3216)) or (layer0_outputs(8511));
    layer1_outputs(10467) <= (layer0_outputs(7578)) and not (layer0_outputs(8370));
    layer1_outputs(10468) <= not(layer0_outputs(7786)) or (layer0_outputs(10370));
    layer1_outputs(10469) <= not((layer0_outputs(3465)) or (layer0_outputs(6629)));
    layer1_outputs(10470) <= not(layer0_outputs(9438)) or (layer0_outputs(8650));
    layer1_outputs(10471) <= layer0_outputs(247);
    layer1_outputs(10472) <= not(layer0_outputs(6394));
    layer1_outputs(10473) <= layer0_outputs(11854);
    layer1_outputs(10474) <= layer0_outputs(10951);
    layer1_outputs(10475) <= layer0_outputs(1662);
    layer1_outputs(10476) <= layer0_outputs(11500);
    layer1_outputs(10477) <= not(layer0_outputs(8411));
    layer1_outputs(10478) <= '0';
    layer1_outputs(10479) <= not((layer0_outputs(8107)) or (layer0_outputs(11247)));
    layer1_outputs(10480) <= (layer0_outputs(2816)) and not (layer0_outputs(9472));
    layer1_outputs(10481) <= '0';
    layer1_outputs(10482) <= layer0_outputs(8759);
    layer1_outputs(10483) <= layer0_outputs(7254);
    layer1_outputs(10484) <= (layer0_outputs(2218)) and (layer0_outputs(2908));
    layer1_outputs(10485) <= not(layer0_outputs(12749)) or (layer0_outputs(8277));
    layer1_outputs(10486) <= not((layer0_outputs(8014)) and (layer0_outputs(5929)));
    layer1_outputs(10487) <= not(layer0_outputs(11220));
    layer1_outputs(10488) <= not(layer0_outputs(8461));
    layer1_outputs(10489) <= (layer0_outputs(172)) and not (layer0_outputs(1966));
    layer1_outputs(10490) <= not((layer0_outputs(485)) xor (layer0_outputs(6755)));
    layer1_outputs(10491) <= not(layer0_outputs(600)) or (layer0_outputs(4705));
    layer1_outputs(10492) <= not((layer0_outputs(577)) xor (layer0_outputs(6002)));
    layer1_outputs(10493) <= (layer0_outputs(5598)) xor (layer0_outputs(9076));
    layer1_outputs(10494) <= not(layer0_outputs(1538));
    layer1_outputs(10495) <= not(layer0_outputs(1419)) or (layer0_outputs(10329));
    layer1_outputs(10496) <= not(layer0_outputs(4177));
    layer1_outputs(10497) <= not((layer0_outputs(11607)) or (layer0_outputs(3436)));
    layer1_outputs(10498) <= not(layer0_outputs(1563));
    layer1_outputs(10499) <= not(layer0_outputs(675)) or (layer0_outputs(4384));
    layer1_outputs(10500) <= layer0_outputs(5576);
    layer1_outputs(10501) <= not(layer0_outputs(9035));
    layer1_outputs(10502) <= not(layer0_outputs(6020));
    layer1_outputs(10503) <= not(layer0_outputs(6453)) or (layer0_outputs(3657));
    layer1_outputs(10504) <= (layer0_outputs(2636)) and not (layer0_outputs(5064));
    layer1_outputs(10505) <= not(layer0_outputs(2043));
    layer1_outputs(10506) <= layer0_outputs(9937);
    layer1_outputs(10507) <= (layer0_outputs(3737)) or (layer0_outputs(2466));
    layer1_outputs(10508) <= not(layer0_outputs(7588));
    layer1_outputs(10509) <= layer0_outputs(6561);
    layer1_outputs(10510) <= (layer0_outputs(7518)) and (layer0_outputs(563));
    layer1_outputs(10511) <= not((layer0_outputs(7527)) or (layer0_outputs(2660)));
    layer1_outputs(10512) <= '1';
    layer1_outputs(10513) <= (layer0_outputs(4982)) and not (layer0_outputs(8266));
    layer1_outputs(10514) <= (layer0_outputs(5462)) and (layer0_outputs(6341));
    layer1_outputs(10515) <= not(layer0_outputs(268));
    layer1_outputs(10516) <= not(layer0_outputs(3201)) or (layer0_outputs(5247));
    layer1_outputs(10517) <= not((layer0_outputs(7919)) or (layer0_outputs(1559)));
    layer1_outputs(10518) <= (layer0_outputs(2334)) and not (layer0_outputs(4437));
    layer1_outputs(10519) <= not(layer0_outputs(2061)) or (layer0_outputs(9440));
    layer1_outputs(10520) <= not(layer0_outputs(5819));
    layer1_outputs(10521) <= not((layer0_outputs(11174)) and (layer0_outputs(7381)));
    layer1_outputs(10522) <= (layer0_outputs(9292)) xor (layer0_outputs(1348));
    layer1_outputs(10523) <= (layer0_outputs(8262)) and not (layer0_outputs(1936));
    layer1_outputs(10524) <= not((layer0_outputs(9126)) or (layer0_outputs(9845)));
    layer1_outputs(10525) <= not(layer0_outputs(9103)) or (layer0_outputs(6781));
    layer1_outputs(10526) <= (layer0_outputs(2286)) and not (layer0_outputs(1731));
    layer1_outputs(10527) <= not(layer0_outputs(7856)) or (layer0_outputs(3202));
    layer1_outputs(10528) <= layer0_outputs(11439);
    layer1_outputs(10529) <= not((layer0_outputs(12730)) and (layer0_outputs(10636)));
    layer1_outputs(10530) <= layer0_outputs(1069);
    layer1_outputs(10531) <= (layer0_outputs(3176)) xor (layer0_outputs(9812));
    layer1_outputs(10532) <= not((layer0_outputs(11952)) and (layer0_outputs(234)));
    layer1_outputs(10533) <= (layer0_outputs(8896)) and not (layer0_outputs(9715));
    layer1_outputs(10534) <= not(layer0_outputs(8069));
    layer1_outputs(10535) <= not(layer0_outputs(2013));
    layer1_outputs(10536) <= layer0_outputs(6828);
    layer1_outputs(10537) <= not((layer0_outputs(6008)) or (layer0_outputs(1758)));
    layer1_outputs(10538) <= not(layer0_outputs(9403));
    layer1_outputs(10539) <= (layer0_outputs(4111)) xor (layer0_outputs(11652));
    layer1_outputs(10540) <= not(layer0_outputs(9136));
    layer1_outputs(10541) <= '1';
    layer1_outputs(10542) <= not((layer0_outputs(11798)) and (layer0_outputs(2196)));
    layer1_outputs(10543) <= (layer0_outputs(9155)) or (layer0_outputs(1775));
    layer1_outputs(10544) <= not((layer0_outputs(11300)) or (layer0_outputs(11456)));
    layer1_outputs(10545) <= (layer0_outputs(3763)) xor (layer0_outputs(9417));
    layer1_outputs(10546) <= layer0_outputs(5373);
    layer1_outputs(10547) <= (layer0_outputs(11125)) xor (layer0_outputs(270));
    layer1_outputs(10548) <= '0';
    layer1_outputs(10549) <= not(layer0_outputs(7910)) or (layer0_outputs(702));
    layer1_outputs(10550) <= (layer0_outputs(8922)) or (layer0_outputs(10326));
    layer1_outputs(10551) <= (layer0_outputs(7162)) xor (layer0_outputs(327));
    layer1_outputs(10552) <= (layer0_outputs(7236)) xor (layer0_outputs(9123));
    layer1_outputs(10553) <= not(layer0_outputs(11691));
    layer1_outputs(10554) <= not((layer0_outputs(4508)) and (layer0_outputs(7452)));
    layer1_outputs(10555) <= not(layer0_outputs(5888)) or (layer0_outputs(11378));
    layer1_outputs(10556) <= not(layer0_outputs(10794)) or (layer0_outputs(12701));
    layer1_outputs(10557) <= not(layer0_outputs(1215));
    layer1_outputs(10558) <= '0';
    layer1_outputs(10559) <= not((layer0_outputs(11443)) or (layer0_outputs(6068)));
    layer1_outputs(10560) <= (layer0_outputs(12204)) and not (layer0_outputs(2296));
    layer1_outputs(10561) <= (layer0_outputs(7260)) or (layer0_outputs(5780));
    layer1_outputs(10562) <= not(layer0_outputs(7617)) or (layer0_outputs(5724));
    layer1_outputs(10563) <= not(layer0_outputs(5123));
    layer1_outputs(10564) <= not(layer0_outputs(6882));
    layer1_outputs(10565) <= layer0_outputs(2296);
    layer1_outputs(10566) <= not(layer0_outputs(11287)) or (layer0_outputs(11854));
    layer1_outputs(10567) <= layer0_outputs(5152);
    layer1_outputs(10568) <= layer0_outputs(11345);
    layer1_outputs(10569) <= layer0_outputs(7413);
    layer1_outputs(10570) <= not(layer0_outputs(958));
    layer1_outputs(10571) <= (layer0_outputs(10558)) and not (layer0_outputs(3078));
    layer1_outputs(10572) <= (layer0_outputs(1025)) and not (layer0_outputs(3235));
    layer1_outputs(10573) <= not(layer0_outputs(10889)) or (layer0_outputs(7063));
    layer1_outputs(10574) <= not(layer0_outputs(9727)) or (layer0_outputs(3971));
    layer1_outputs(10575) <= (layer0_outputs(4507)) and (layer0_outputs(37));
    layer1_outputs(10576) <= not((layer0_outputs(11812)) and (layer0_outputs(8247)));
    layer1_outputs(10577) <= (layer0_outputs(2643)) or (layer0_outputs(7143));
    layer1_outputs(10578) <= '0';
    layer1_outputs(10579) <= not(layer0_outputs(12014));
    layer1_outputs(10580) <= layer0_outputs(3223);
    layer1_outputs(10581) <= not((layer0_outputs(3198)) and (layer0_outputs(3319)));
    layer1_outputs(10582) <= not(layer0_outputs(6584));
    layer1_outputs(10583) <= not((layer0_outputs(7149)) or (layer0_outputs(8630)));
    layer1_outputs(10584) <= not((layer0_outputs(4290)) xor (layer0_outputs(5362)));
    layer1_outputs(10585) <= layer0_outputs(1227);
    layer1_outputs(10586) <= layer0_outputs(3915);
    layer1_outputs(10587) <= not((layer0_outputs(3456)) xor (layer0_outputs(3862)));
    layer1_outputs(10588) <= layer0_outputs(1449);
    layer1_outputs(10589) <= (layer0_outputs(5643)) and not (layer0_outputs(7101));
    layer1_outputs(10590) <= not((layer0_outputs(9881)) or (layer0_outputs(3537)));
    layer1_outputs(10591) <= (layer0_outputs(7620)) xor (layer0_outputs(3275));
    layer1_outputs(10592) <= not((layer0_outputs(8465)) or (layer0_outputs(11769)));
    layer1_outputs(10593) <= not(layer0_outputs(7951)) or (layer0_outputs(8395));
    layer1_outputs(10594) <= not(layer0_outputs(4572));
    layer1_outputs(10595) <= layer0_outputs(9209);
    layer1_outputs(10596) <= not((layer0_outputs(1642)) and (layer0_outputs(685)));
    layer1_outputs(10597) <= not((layer0_outputs(10610)) or (layer0_outputs(7043)));
    layer1_outputs(10598) <= layer0_outputs(8305);
    layer1_outputs(10599) <= not(layer0_outputs(11755));
    layer1_outputs(10600) <= not(layer0_outputs(7241));
    layer1_outputs(10601) <= (layer0_outputs(9377)) and not (layer0_outputs(1406));
    layer1_outputs(10602) <= (layer0_outputs(1866)) and not (layer0_outputs(9591));
    layer1_outputs(10603) <= not(layer0_outputs(8281));
    layer1_outputs(10604) <= (layer0_outputs(10814)) and not (layer0_outputs(11063));
    layer1_outputs(10605) <= (layer0_outputs(10766)) and (layer0_outputs(6298));
    layer1_outputs(10606) <= layer0_outputs(5120);
    layer1_outputs(10607) <= not((layer0_outputs(8338)) or (layer0_outputs(10863)));
    layer1_outputs(10608) <= not(layer0_outputs(4008)) or (layer0_outputs(3023));
    layer1_outputs(10609) <= layer0_outputs(6627);
    layer1_outputs(10610) <= not(layer0_outputs(500));
    layer1_outputs(10611) <= not((layer0_outputs(4601)) xor (layer0_outputs(2723)));
    layer1_outputs(10612) <= layer0_outputs(5519);
    layer1_outputs(10613) <= (layer0_outputs(5307)) xor (layer0_outputs(4411));
    layer1_outputs(10614) <= layer0_outputs(10517);
    layer1_outputs(10615) <= not((layer0_outputs(5251)) or (layer0_outputs(1635)));
    layer1_outputs(10616) <= (layer0_outputs(6897)) and not (layer0_outputs(11331));
    layer1_outputs(10617) <= not(layer0_outputs(6579));
    layer1_outputs(10618) <= (layer0_outputs(581)) or (layer0_outputs(1333));
    layer1_outputs(10619) <= (layer0_outputs(6147)) or (layer0_outputs(8419));
    layer1_outputs(10620) <= layer0_outputs(2263);
    layer1_outputs(10621) <= layer0_outputs(4824);
    layer1_outputs(10622) <= not(layer0_outputs(9345)) or (layer0_outputs(6953));
    layer1_outputs(10623) <= (layer0_outputs(11289)) and not (layer0_outputs(6241));
    layer1_outputs(10624) <= not((layer0_outputs(1102)) or (layer0_outputs(4064)));
    layer1_outputs(10625) <= layer0_outputs(5887);
    layer1_outputs(10626) <= (layer0_outputs(2424)) xor (layer0_outputs(4005));
    layer1_outputs(10627) <= not((layer0_outputs(5363)) or (layer0_outputs(10074)));
    layer1_outputs(10628) <= '1';
    layer1_outputs(10629) <= not(layer0_outputs(8231)) or (layer0_outputs(1608));
    layer1_outputs(10630) <= (layer0_outputs(1786)) and not (layer0_outputs(6718));
    layer1_outputs(10631) <= not(layer0_outputs(220));
    layer1_outputs(10632) <= (layer0_outputs(2050)) xor (layer0_outputs(1360));
    layer1_outputs(10633) <= not((layer0_outputs(6001)) and (layer0_outputs(12275)));
    layer1_outputs(10634) <= layer0_outputs(10443);
    layer1_outputs(10635) <= not(layer0_outputs(5585));
    layer1_outputs(10636) <= (layer0_outputs(7191)) xor (layer0_outputs(5995));
    layer1_outputs(10637) <= layer0_outputs(12722);
    layer1_outputs(10638) <= not(layer0_outputs(4606));
    layer1_outputs(10639) <= not(layer0_outputs(10367));
    layer1_outputs(10640) <= not((layer0_outputs(9813)) xor (layer0_outputs(8127)));
    layer1_outputs(10641) <= not(layer0_outputs(6960)) or (layer0_outputs(4624));
    layer1_outputs(10642) <= not(layer0_outputs(1176));
    layer1_outputs(10643) <= not((layer0_outputs(11656)) and (layer0_outputs(5623)));
    layer1_outputs(10644) <= (layer0_outputs(12050)) and (layer0_outputs(9848));
    layer1_outputs(10645) <= not(layer0_outputs(3984));
    layer1_outputs(10646) <= (layer0_outputs(10883)) or (layer0_outputs(4390));
    layer1_outputs(10647) <= not(layer0_outputs(4216)) or (layer0_outputs(3832));
    layer1_outputs(10648) <= not((layer0_outputs(5377)) or (layer0_outputs(1620)));
    layer1_outputs(10649) <= not(layer0_outputs(8913));
    layer1_outputs(10650) <= not((layer0_outputs(11938)) or (layer0_outputs(10957)));
    layer1_outputs(10651) <= layer0_outputs(11461);
    layer1_outputs(10652) <= not(layer0_outputs(4413)) or (layer0_outputs(2571));
    layer1_outputs(10653) <= not(layer0_outputs(2165));
    layer1_outputs(10654) <= (layer0_outputs(6080)) xor (layer0_outputs(6587));
    layer1_outputs(10655) <= '0';
    layer1_outputs(10656) <= not(layer0_outputs(11582));
    layer1_outputs(10657) <= (layer0_outputs(4096)) and not (layer0_outputs(8608));
    layer1_outputs(10658) <= (layer0_outputs(11754)) and not (layer0_outputs(4423));
    layer1_outputs(10659) <= not(layer0_outputs(11003));
    layer1_outputs(10660) <= (layer0_outputs(9970)) or (layer0_outputs(9380));
    layer1_outputs(10661) <= not(layer0_outputs(3450)) or (layer0_outputs(7895));
    layer1_outputs(10662) <= not((layer0_outputs(4590)) or (layer0_outputs(4046)));
    layer1_outputs(10663) <= not((layer0_outputs(11070)) and (layer0_outputs(12715)));
    layer1_outputs(10664) <= not(layer0_outputs(610));
    layer1_outputs(10665) <= (layer0_outputs(994)) and not (layer0_outputs(679));
    layer1_outputs(10666) <= layer0_outputs(6516);
    layer1_outputs(10667) <= (layer0_outputs(11813)) or (layer0_outputs(9421));
    layer1_outputs(10668) <= not(layer0_outputs(7181)) or (layer0_outputs(6364));
    layer1_outputs(10669) <= not(layer0_outputs(6545));
    layer1_outputs(10670) <= (layer0_outputs(3256)) and not (layer0_outputs(4627));
    layer1_outputs(10671) <= (layer0_outputs(3198)) and not (layer0_outputs(10226));
    layer1_outputs(10672) <= (layer0_outputs(9121)) or (layer0_outputs(3552));
    layer1_outputs(10673) <= (layer0_outputs(5295)) and not (layer0_outputs(3894));
    layer1_outputs(10674) <= (layer0_outputs(8392)) xor (layer0_outputs(1309));
    layer1_outputs(10675) <= not(layer0_outputs(12612)) or (layer0_outputs(7743));
    layer1_outputs(10676) <= (layer0_outputs(3148)) and not (layer0_outputs(10482));
    layer1_outputs(10677) <= not((layer0_outputs(8196)) or (layer0_outputs(853)));
    layer1_outputs(10678) <= (layer0_outputs(11429)) xor (layer0_outputs(2998));
    layer1_outputs(10679) <= not((layer0_outputs(2247)) and (layer0_outputs(6381)));
    layer1_outputs(10680) <= (layer0_outputs(1151)) and not (layer0_outputs(7796));
    layer1_outputs(10681) <= layer0_outputs(39);
    layer1_outputs(10682) <= not(layer0_outputs(10821));
    layer1_outputs(10683) <= layer0_outputs(4003);
    layer1_outputs(10684) <= layer0_outputs(2141);
    layer1_outputs(10685) <= not(layer0_outputs(1335)) or (layer0_outputs(12649));
    layer1_outputs(10686) <= not((layer0_outputs(4059)) or (layer0_outputs(9203)));
    layer1_outputs(10687) <= not(layer0_outputs(9350));
    layer1_outputs(10688) <= (layer0_outputs(4567)) xor (layer0_outputs(11639));
    layer1_outputs(10689) <= not((layer0_outputs(7317)) or (layer0_outputs(3829)));
    layer1_outputs(10690) <= not((layer0_outputs(3162)) xor (layer0_outputs(7585)));
    layer1_outputs(10691) <= layer0_outputs(10808);
    layer1_outputs(10692) <= '1';
    layer1_outputs(10693) <= not(layer0_outputs(9379)) or (layer0_outputs(11676));
    layer1_outputs(10694) <= not(layer0_outputs(6638));
    layer1_outputs(10695) <= not((layer0_outputs(11739)) and (layer0_outputs(9171)));
    layer1_outputs(10696) <= not(layer0_outputs(60));
    layer1_outputs(10697) <= not(layer0_outputs(5358));
    layer1_outputs(10698) <= not(layer0_outputs(2470));
    layer1_outputs(10699) <= not((layer0_outputs(7673)) xor (layer0_outputs(8141)));
    layer1_outputs(10700) <= not((layer0_outputs(7593)) or (layer0_outputs(5602)));
    layer1_outputs(10701) <= (layer0_outputs(2526)) xor (layer0_outputs(12179));
    layer1_outputs(10702) <= (layer0_outputs(3561)) xor (layer0_outputs(8057));
    layer1_outputs(10703) <= (layer0_outputs(10801)) and (layer0_outputs(6960));
    layer1_outputs(10704) <= layer0_outputs(610);
    layer1_outputs(10705) <= not(layer0_outputs(11054)) or (layer0_outputs(11830));
    layer1_outputs(10706) <= not((layer0_outputs(1501)) and (layer0_outputs(2207)));
    layer1_outputs(10707) <= not(layer0_outputs(10572)) or (layer0_outputs(4632));
    layer1_outputs(10708) <= layer0_outputs(11551);
    layer1_outputs(10709) <= layer0_outputs(7340);
    layer1_outputs(10710) <= (layer0_outputs(6169)) xor (layer0_outputs(49));
    layer1_outputs(10711) <= (layer0_outputs(9644)) and not (layer0_outputs(5271));
    layer1_outputs(10712) <= not(layer0_outputs(1148));
    layer1_outputs(10713) <= layer0_outputs(9686);
    layer1_outputs(10714) <= not(layer0_outputs(10814));
    layer1_outputs(10715) <= not(layer0_outputs(8607));
    layer1_outputs(10716) <= not(layer0_outputs(12508));
    layer1_outputs(10717) <= not(layer0_outputs(6078));
    layer1_outputs(10718) <= (layer0_outputs(11091)) xor (layer0_outputs(12033));
    layer1_outputs(10719) <= not(layer0_outputs(11278));
    layer1_outputs(10720) <= not((layer0_outputs(2497)) and (layer0_outputs(7889)));
    layer1_outputs(10721) <= '0';
    layer1_outputs(10722) <= (layer0_outputs(5568)) and not (layer0_outputs(5868));
    layer1_outputs(10723) <= layer0_outputs(580);
    layer1_outputs(10724) <= '1';
    layer1_outputs(10725) <= not((layer0_outputs(1978)) or (layer0_outputs(11220)));
    layer1_outputs(10726) <= not((layer0_outputs(7236)) and (layer0_outputs(3589)));
    layer1_outputs(10727) <= not(layer0_outputs(11591));
    layer1_outputs(10728) <= not((layer0_outputs(3560)) or (layer0_outputs(7257)));
    layer1_outputs(10729) <= not(layer0_outputs(12318));
    layer1_outputs(10730) <= not(layer0_outputs(9249));
    layer1_outputs(10731) <= layer0_outputs(7574);
    layer1_outputs(10732) <= not(layer0_outputs(4519));
    layer1_outputs(10733) <= (layer0_outputs(10905)) and (layer0_outputs(6295));
    layer1_outputs(10734) <= layer0_outputs(1911);
    layer1_outputs(10735) <= layer0_outputs(9410);
    layer1_outputs(10736) <= not((layer0_outputs(12083)) and (layer0_outputs(8231)));
    layer1_outputs(10737) <= not((layer0_outputs(2718)) and (layer0_outputs(1060)));
    layer1_outputs(10738) <= (layer0_outputs(3280)) or (layer0_outputs(199));
    layer1_outputs(10739) <= not(layer0_outputs(12761));
    layer1_outputs(10740) <= layer0_outputs(3651);
    layer1_outputs(10741) <= not(layer0_outputs(3032));
    layer1_outputs(10742) <= layer0_outputs(1017);
    layer1_outputs(10743) <= (layer0_outputs(7388)) or (layer0_outputs(6840));
    layer1_outputs(10744) <= not((layer0_outputs(6904)) xor (layer0_outputs(5525)));
    layer1_outputs(10745) <= not((layer0_outputs(3422)) and (layer0_outputs(2928)));
    layer1_outputs(10746) <= layer0_outputs(3419);
    layer1_outputs(10747) <= layer0_outputs(11079);
    layer1_outputs(10748) <= (layer0_outputs(5399)) xor (layer0_outputs(1414));
    layer1_outputs(10749) <= (layer0_outputs(5407)) and (layer0_outputs(4986));
    layer1_outputs(10750) <= layer0_outputs(2105);
    layer1_outputs(10751) <= layer0_outputs(3707);
    layer1_outputs(10752) <= (layer0_outputs(3116)) and not (layer0_outputs(2597));
    layer1_outputs(10753) <= not(layer0_outputs(5145));
    layer1_outputs(10754) <= layer0_outputs(6378);
    layer1_outputs(10755) <= (layer0_outputs(6544)) and not (layer0_outputs(1202));
    layer1_outputs(10756) <= layer0_outputs(3831);
    layer1_outputs(10757) <= not(layer0_outputs(3059)) or (layer0_outputs(9255));
    layer1_outputs(10758) <= not((layer0_outputs(777)) and (layer0_outputs(5491)));
    layer1_outputs(10759) <= not(layer0_outputs(6549)) or (layer0_outputs(8954));
    layer1_outputs(10760) <= (layer0_outputs(5698)) or (layer0_outputs(8299));
    layer1_outputs(10761) <= not(layer0_outputs(11517));
    layer1_outputs(10762) <= not((layer0_outputs(8810)) xor (layer0_outputs(7546)));
    layer1_outputs(10763) <= not((layer0_outputs(1303)) or (layer0_outputs(8737)));
    layer1_outputs(10764) <= layer0_outputs(3117);
    layer1_outputs(10765) <= not(layer0_outputs(3518));
    layer1_outputs(10766) <= not((layer0_outputs(9215)) or (layer0_outputs(1875)));
    layer1_outputs(10767) <= not((layer0_outputs(9134)) xor (layer0_outputs(8692)));
    layer1_outputs(10768) <= '0';
    layer1_outputs(10769) <= not(layer0_outputs(7061));
    layer1_outputs(10770) <= (layer0_outputs(2803)) and (layer0_outputs(1960));
    layer1_outputs(10771) <= (layer0_outputs(1671)) and not (layer0_outputs(4279));
    layer1_outputs(10772) <= layer0_outputs(8548);
    layer1_outputs(10773) <= layer0_outputs(12603);
    layer1_outputs(10774) <= layer0_outputs(9514);
    layer1_outputs(10775) <= (layer0_outputs(8044)) and not (layer0_outputs(9376));
    layer1_outputs(10776) <= (layer0_outputs(11079)) or (layer0_outputs(8260));
    layer1_outputs(10777) <= not(layer0_outputs(9894)) or (layer0_outputs(10533));
    layer1_outputs(10778) <= not((layer0_outputs(8217)) and (layer0_outputs(10538)));
    layer1_outputs(10779) <= layer0_outputs(3423);
    layer1_outputs(10780) <= not((layer0_outputs(1961)) or (layer0_outputs(6949)));
    layer1_outputs(10781) <= (layer0_outputs(653)) and not (layer0_outputs(6262));
    layer1_outputs(10782) <= not(layer0_outputs(8204));
    layer1_outputs(10783) <= (layer0_outputs(10655)) and not (layer0_outputs(8415));
    layer1_outputs(10784) <= not(layer0_outputs(5778)) or (layer0_outputs(9043));
    layer1_outputs(10785) <= not(layer0_outputs(428));
    layer1_outputs(10786) <= layer0_outputs(11860);
    layer1_outputs(10787) <= (layer0_outputs(3505)) or (layer0_outputs(7257));
    layer1_outputs(10788) <= not(layer0_outputs(1722));
    layer1_outputs(10789) <= not(layer0_outputs(10255)) or (layer0_outputs(9422));
    layer1_outputs(10790) <= (layer0_outputs(3515)) and not (layer0_outputs(3627));
    layer1_outputs(10791) <= (layer0_outputs(4484)) and not (layer0_outputs(5600));
    layer1_outputs(10792) <= not(layer0_outputs(4694)) or (layer0_outputs(2263));
    layer1_outputs(10793) <= (layer0_outputs(12250)) and not (layer0_outputs(1220));
    layer1_outputs(10794) <= (layer0_outputs(7686)) and (layer0_outputs(1466));
    layer1_outputs(10795) <= (layer0_outputs(9401)) or (layer0_outputs(12338));
    layer1_outputs(10796) <= not((layer0_outputs(4435)) xor (layer0_outputs(10917)));
    layer1_outputs(10797) <= (layer0_outputs(9310)) and (layer0_outputs(5641));
    layer1_outputs(10798) <= not((layer0_outputs(7146)) xor (layer0_outputs(4178)));
    layer1_outputs(10799) <= layer0_outputs(3200);
    layer1_outputs(10800) <= not(layer0_outputs(10896));
    layer1_outputs(10801) <= (layer0_outputs(793)) or (layer0_outputs(3314));
    layer1_outputs(10802) <= layer0_outputs(1549);
    layer1_outputs(10803) <= not((layer0_outputs(6872)) or (layer0_outputs(9900)));
    layer1_outputs(10804) <= layer0_outputs(11271);
    layer1_outputs(10805) <= layer0_outputs(8791);
    layer1_outputs(10806) <= layer0_outputs(4327);
    layer1_outputs(10807) <= layer0_outputs(10898);
    layer1_outputs(10808) <= not(layer0_outputs(9414)) or (layer0_outputs(2251));
    layer1_outputs(10809) <= layer0_outputs(8639);
    layer1_outputs(10810) <= (layer0_outputs(10829)) xor (layer0_outputs(7325));
    layer1_outputs(10811) <= (layer0_outputs(5826)) and not (layer0_outputs(7540));
    layer1_outputs(10812) <= not(layer0_outputs(11874));
    layer1_outputs(10813) <= (layer0_outputs(10989)) xor (layer0_outputs(7828));
    layer1_outputs(10814) <= not(layer0_outputs(5371));
    layer1_outputs(10815) <= layer0_outputs(10370);
    layer1_outputs(10816) <= not((layer0_outputs(7050)) xor (layer0_outputs(30)));
    layer1_outputs(10817) <= not(layer0_outputs(11392));
    layer1_outputs(10818) <= not(layer0_outputs(7385));
    layer1_outputs(10819) <= not(layer0_outputs(2330)) or (layer0_outputs(4219));
    layer1_outputs(10820) <= (layer0_outputs(10571)) and not (layer0_outputs(6647));
    layer1_outputs(10821) <= not((layer0_outputs(2709)) or (layer0_outputs(10474)));
    layer1_outputs(10822) <= (layer0_outputs(1536)) xor (layer0_outputs(10551));
    layer1_outputs(10823) <= (layer0_outputs(6336)) and not (layer0_outputs(12599));
    layer1_outputs(10824) <= (layer0_outputs(637)) and not (layer0_outputs(1792));
    layer1_outputs(10825) <= not(layer0_outputs(589));
    layer1_outputs(10826) <= not(layer0_outputs(4791));
    layer1_outputs(10827) <= not(layer0_outputs(8178));
    layer1_outputs(10828) <= layer0_outputs(5648);
    layer1_outputs(10829) <= (layer0_outputs(385)) and not (layer0_outputs(992));
    layer1_outputs(10830) <= layer0_outputs(11229);
    layer1_outputs(10831) <= not(layer0_outputs(3546)) or (layer0_outputs(7283));
    layer1_outputs(10832) <= not(layer0_outputs(6690));
    layer1_outputs(10833) <= (layer0_outputs(7721)) and not (layer0_outputs(2137));
    layer1_outputs(10834) <= (layer0_outputs(11472)) and not (layer0_outputs(8135));
    layer1_outputs(10835) <= (layer0_outputs(7170)) or (layer0_outputs(2245));
    layer1_outputs(10836) <= not(layer0_outputs(11438)) or (layer0_outputs(6415));
    layer1_outputs(10837) <= not(layer0_outputs(9208));
    layer1_outputs(10838) <= layer0_outputs(11883);
    layer1_outputs(10839) <= not(layer0_outputs(12564)) or (layer0_outputs(10857));
    layer1_outputs(10840) <= not(layer0_outputs(4913)) or (layer0_outputs(1932));
    layer1_outputs(10841) <= (layer0_outputs(5391)) and not (layer0_outputs(2661));
    layer1_outputs(10842) <= not((layer0_outputs(9145)) and (layer0_outputs(7628)));
    layer1_outputs(10843) <= (layer0_outputs(12640)) and (layer0_outputs(2382));
    layer1_outputs(10844) <= '0';
    layer1_outputs(10845) <= not(layer0_outputs(7464));
    layer1_outputs(10846) <= not((layer0_outputs(12160)) and (layer0_outputs(7992)));
    layer1_outputs(10847) <= layer0_outputs(798);
    layer1_outputs(10848) <= (layer0_outputs(11155)) and not (layer0_outputs(406));
    layer1_outputs(10849) <= not(layer0_outputs(8700)) or (layer0_outputs(1741));
    layer1_outputs(10850) <= not(layer0_outputs(7097));
    layer1_outputs(10851) <= '0';
    layer1_outputs(10852) <= not(layer0_outputs(3819)) or (layer0_outputs(3090));
    layer1_outputs(10853) <= not(layer0_outputs(217));
    layer1_outputs(10854) <= not(layer0_outputs(5632));
    layer1_outputs(10855) <= (layer0_outputs(6484)) and not (layer0_outputs(2166));
    layer1_outputs(10856) <= not((layer0_outputs(9378)) or (layer0_outputs(5036)));
    layer1_outputs(10857) <= not(layer0_outputs(5299)) or (layer0_outputs(363));
    layer1_outputs(10858) <= (layer0_outputs(8522)) and (layer0_outputs(971));
    layer1_outputs(10859) <= not((layer0_outputs(11223)) and (layer0_outputs(12126)));
    layer1_outputs(10860) <= (layer0_outputs(11298)) and (layer0_outputs(6562));
    layer1_outputs(10861) <= not(layer0_outputs(5443));
    layer1_outputs(10862) <= not((layer0_outputs(849)) and (layer0_outputs(5071)));
    layer1_outputs(10863) <= (layer0_outputs(5162)) and (layer0_outputs(2082));
    layer1_outputs(10864) <= (layer0_outputs(2127)) and not (layer0_outputs(7048));
    layer1_outputs(10865) <= not(layer0_outputs(2783)) or (layer0_outputs(10518));
    layer1_outputs(10866) <= not(layer0_outputs(5787)) or (layer0_outputs(9892));
    layer1_outputs(10867) <= (layer0_outputs(12383)) and (layer0_outputs(3519));
    layer1_outputs(10868) <= (layer0_outputs(8363)) or (layer0_outputs(9413));
    layer1_outputs(10869) <= not(layer0_outputs(8899)) or (layer0_outputs(7992));
    layer1_outputs(10870) <= not((layer0_outputs(6818)) and (layer0_outputs(2559)));
    layer1_outputs(10871) <= (layer0_outputs(137)) or (layer0_outputs(7846));
    layer1_outputs(10872) <= '1';
    layer1_outputs(10873) <= not(layer0_outputs(1967));
    layer1_outputs(10874) <= not(layer0_outputs(5134)) or (layer0_outputs(8496));
    layer1_outputs(10875) <= not(layer0_outputs(5418));
    layer1_outputs(10876) <= (layer0_outputs(8167)) and not (layer0_outputs(4676));
    layer1_outputs(10877) <= not(layer0_outputs(10279)) or (layer0_outputs(637));
    layer1_outputs(10878) <= not(layer0_outputs(5956));
    layer1_outputs(10879) <= (layer0_outputs(3373)) and (layer0_outputs(7189));
    layer1_outputs(10880) <= (layer0_outputs(6665)) and not (layer0_outputs(9934));
    layer1_outputs(10881) <= not(layer0_outputs(10235)) or (layer0_outputs(3131));
    layer1_outputs(10882) <= (layer0_outputs(1750)) and not (layer0_outputs(8209));
    layer1_outputs(10883) <= layer0_outputs(9551);
    layer1_outputs(10884) <= not((layer0_outputs(3727)) and (layer0_outputs(30)));
    layer1_outputs(10885) <= layer0_outputs(1041);
    layer1_outputs(10886) <= not(layer0_outputs(4123)) or (layer0_outputs(1336));
    layer1_outputs(10887) <= (layer0_outputs(10530)) and not (layer0_outputs(11750));
    layer1_outputs(10888) <= not(layer0_outputs(11655));
    layer1_outputs(10889) <= not((layer0_outputs(5706)) xor (layer0_outputs(10146)));
    layer1_outputs(10890) <= layer0_outputs(6159);
    layer1_outputs(10891) <= not(layer0_outputs(2774)) or (layer0_outputs(1485));
    layer1_outputs(10892) <= not(layer0_outputs(10742));
    layer1_outputs(10893) <= not(layer0_outputs(12436)) or (layer0_outputs(7607));
    layer1_outputs(10894) <= (layer0_outputs(10256)) or (layer0_outputs(1122));
    layer1_outputs(10895) <= layer0_outputs(3626);
    layer1_outputs(10896) <= (layer0_outputs(2372)) and not (layer0_outputs(6985));
    layer1_outputs(10897) <= (layer0_outputs(10777)) and (layer0_outputs(11672));
    layer1_outputs(10898) <= not(layer0_outputs(7282));
    layer1_outputs(10899) <= not((layer0_outputs(12073)) or (layer0_outputs(11055)));
    layer1_outputs(10900) <= layer0_outputs(4378);
    layer1_outputs(10901) <= layer0_outputs(9027);
    layer1_outputs(10902) <= not(layer0_outputs(8666)) or (layer0_outputs(7721));
    layer1_outputs(10903) <= not((layer0_outputs(7195)) or (layer0_outputs(12771)));
    layer1_outputs(10904) <= layer0_outputs(8352);
    layer1_outputs(10905) <= not(layer0_outputs(2331)) or (layer0_outputs(5682));
    layer1_outputs(10906) <= not((layer0_outputs(2528)) xor (layer0_outputs(5312)));
    layer1_outputs(10907) <= not(layer0_outputs(11989));
    layer1_outputs(10908) <= '1';
    layer1_outputs(10909) <= layer0_outputs(2826);
    layer1_outputs(10910) <= not((layer0_outputs(11365)) and (layer0_outputs(265)));
    layer1_outputs(10911) <= not(layer0_outputs(8662));
    layer1_outputs(10912) <= (layer0_outputs(6379)) or (layer0_outputs(9244));
    layer1_outputs(10913) <= layer0_outputs(1966);
    layer1_outputs(10914) <= layer0_outputs(9124);
    layer1_outputs(10915) <= not((layer0_outputs(2139)) and (layer0_outputs(12577)));
    layer1_outputs(10916) <= (layer0_outputs(11262)) and not (layer0_outputs(3364));
    layer1_outputs(10917) <= (layer0_outputs(3190)) and (layer0_outputs(11511));
    layer1_outputs(10918) <= layer0_outputs(677);
    layer1_outputs(10919) <= (layer0_outputs(2383)) and not (layer0_outputs(5705));
    layer1_outputs(10920) <= layer0_outputs(5864);
    layer1_outputs(10921) <= '1';
    layer1_outputs(10922) <= layer0_outputs(11502);
    layer1_outputs(10923) <= (layer0_outputs(7712)) xor (layer0_outputs(10840));
    layer1_outputs(10924) <= not((layer0_outputs(5034)) and (layer0_outputs(4555)));
    layer1_outputs(10925) <= not(layer0_outputs(3136));
    layer1_outputs(10926) <= (layer0_outputs(10516)) and not (layer0_outputs(9437));
    layer1_outputs(10927) <= (layer0_outputs(11697)) xor (layer0_outputs(2461));
    layer1_outputs(10928) <= (layer0_outputs(4487)) xor (layer0_outputs(10198));
    layer1_outputs(10929) <= layer0_outputs(5073);
    layer1_outputs(10930) <= (layer0_outputs(12016)) and not (layer0_outputs(3274));
    layer1_outputs(10931) <= (layer0_outputs(5590)) and not (layer0_outputs(5359));
    layer1_outputs(10932) <= layer0_outputs(8183);
    layer1_outputs(10933) <= layer0_outputs(5865);
    layer1_outputs(10934) <= not(layer0_outputs(8555));
    layer1_outputs(10935) <= (layer0_outputs(4423)) xor (layer0_outputs(7203));
    layer1_outputs(10936) <= '0';
    layer1_outputs(10937) <= not((layer0_outputs(6071)) xor (layer0_outputs(3368)));
    layer1_outputs(10938) <= (layer0_outputs(7956)) and not (layer0_outputs(966));
    layer1_outputs(10939) <= (layer0_outputs(116)) or (layer0_outputs(5106));
    layer1_outputs(10940) <= layer0_outputs(2872);
    layer1_outputs(10941) <= layer0_outputs(5172);
    layer1_outputs(10942) <= (layer0_outputs(6631)) and not (layer0_outputs(7528));
    layer1_outputs(10943) <= not(layer0_outputs(11828)) or (layer0_outputs(2869));
    layer1_outputs(10944) <= (layer0_outputs(10974)) or (layer0_outputs(12213));
    layer1_outputs(10945) <= (layer0_outputs(12643)) or (layer0_outputs(1425));
    layer1_outputs(10946) <= not(layer0_outputs(12743));
    layer1_outputs(10947) <= (layer0_outputs(11448)) xor (layer0_outputs(6554));
    layer1_outputs(10948) <= layer0_outputs(1480);
    layer1_outputs(10949) <= not((layer0_outputs(4565)) and (layer0_outputs(9777)));
    layer1_outputs(10950) <= layer0_outputs(11106);
    layer1_outputs(10951) <= (layer0_outputs(10750)) or (layer0_outputs(11774));
    layer1_outputs(10952) <= (layer0_outputs(8099)) and (layer0_outputs(10308));
    layer1_outputs(10953) <= not((layer0_outputs(6486)) and (layer0_outputs(10876)));
    layer1_outputs(10954) <= not((layer0_outputs(3313)) and (layer0_outputs(5967)));
    layer1_outputs(10955) <= (layer0_outputs(10468)) and not (layer0_outputs(12024));
    layer1_outputs(10956) <= not(layer0_outputs(4620)) or (layer0_outputs(9633));
    layer1_outputs(10957) <= layer0_outputs(11962);
    layer1_outputs(10958) <= not(layer0_outputs(12403)) or (layer0_outputs(389));
    layer1_outputs(10959) <= (layer0_outputs(3400)) and not (layer0_outputs(8117));
    layer1_outputs(10960) <= (layer0_outputs(10142)) and not (layer0_outputs(10615));
    layer1_outputs(10961) <= layer0_outputs(8484);
    layer1_outputs(10962) <= not(layer0_outputs(4056));
    layer1_outputs(10963) <= '1';
    layer1_outputs(10964) <= layer0_outputs(7210);
    layer1_outputs(10965) <= (layer0_outputs(219)) and (layer0_outputs(5583));
    layer1_outputs(10966) <= not(layer0_outputs(8989));
    layer1_outputs(10967) <= not(layer0_outputs(12225));
    layer1_outputs(10968) <= not(layer0_outputs(7204));
    layer1_outputs(10969) <= not((layer0_outputs(9376)) and (layer0_outputs(3503)));
    layer1_outputs(10970) <= (layer0_outputs(5793)) or (layer0_outputs(8000));
    layer1_outputs(10971) <= not(layer0_outputs(3369));
    layer1_outputs(10972) <= (layer0_outputs(2504)) xor (layer0_outputs(9857));
    layer1_outputs(10973) <= not(layer0_outputs(7560));
    layer1_outputs(10974) <= layer0_outputs(7715);
    layer1_outputs(10975) <= layer0_outputs(688);
    layer1_outputs(10976) <= layer0_outputs(10528);
    layer1_outputs(10977) <= not((layer0_outputs(8945)) and (layer0_outputs(6950)));
    layer1_outputs(10978) <= (layer0_outputs(9863)) and (layer0_outputs(1788));
    layer1_outputs(10979) <= layer0_outputs(10532);
    layer1_outputs(10980) <= (layer0_outputs(9473)) or (layer0_outputs(9037));
    layer1_outputs(10981) <= layer0_outputs(3902);
    layer1_outputs(10982) <= (layer0_outputs(6811)) and not (layer0_outputs(2743));
    layer1_outputs(10983) <= not((layer0_outputs(6979)) xor (layer0_outputs(8050)));
    layer1_outputs(10984) <= not(layer0_outputs(3157));
    layer1_outputs(10985) <= layer0_outputs(1357);
    layer1_outputs(10986) <= not(layer0_outputs(5972));
    layer1_outputs(10987) <= (layer0_outputs(1847)) and not (layer0_outputs(5381));
    layer1_outputs(10988) <= not(layer0_outputs(11014));
    layer1_outputs(10989) <= not(layer0_outputs(1525));
    layer1_outputs(10990) <= (layer0_outputs(2860)) and (layer0_outputs(8549));
    layer1_outputs(10991) <= (layer0_outputs(4124)) and (layer0_outputs(8592));
    layer1_outputs(10992) <= layer0_outputs(1305);
    layer1_outputs(10993) <= (layer0_outputs(1444)) and not (layer0_outputs(11973));
    layer1_outputs(10994) <= not(layer0_outputs(10219));
    layer1_outputs(10995) <= not(layer0_outputs(9632));
    layer1_outputs(10996) <= not(layer0_outputs(4197)) or (layer0_outputs(9402));
    layer1_outputs(10997) <= (layer0_outputs(9171)) and not (layer0_outputs(4645));
    layer1_outputs(10998) <= not((layer0_outputs(1316)) or (layer0_outputs(1639)));
    layer1_outputs(10999) <= (layer0_outputs(2536)) and not (layer0_outputs(990));
    layer1_outputs(11000) <= not((layer0_outputs(5336)) xor (layer0_outputs(4127)));
    layer1_outputs(11001) <= not((layer0_outputs(3293)) xor (layer0_outputs(10094)));
    layer1_outputs(11002) <= not((layer0_outputs(5147)) xor (layer0_outputs(794)));
    layer1_outputs(11003) <= not(layer0_outputs(5925));
    layer1_outputs(11004) <= layer0_outputs(8695);
    layer1_outputs(11005) <= not(layer0_outputs(7065)) or (layer0_outputs(12602));
    layer1_outputs(11006) <= not((layer0_outputs(4844)) or (layer0_outputs(125)));
    layer1_outputs(11007) <= '1';
    layer1_outputs(11008) <= not((layer0_outputs(4190)) and (layer0_outputs(559)));
    layer1_outputs(11009) <= not(layer0_outputs(12562)) or (layer0_outputs(6541));
    layer1_outputs(11010) <= layer0_outputs(9736);
    layer1_outputs(11011) <= not((layer0_outputs(12786)) xor (layer0_outputs(7194)));
    layer1_outputs(11012) <= not(layer0_outputs(6806));
    layer1_outputs(11013) <= not((layer0_outputs(9518)) xor (layer0_outputs(5535)));
    layer1_outputs(11014) <= not(layer0_outputs(4772));
    layer1_outputs(11015) <= not((layer0_outputs(11819)) or (layer0_outputs(1129)));
    layer1_outputs(11016) <= not((layer0_outputs(12313)) and (layer0_outputs(5416)));
    layer1_outputs(11017) <= not(layer0_outputs(12343));
    layer1_outputs(11018) <= layer0_outputs(3714);
    layer1_outputs(11019) <= (layer0_outputs(3155)) and not (layer0_outputs(6244));
    layer1_outputs(11020) <= (layer0_outputs(6216)) and not (layer0_outputs(1173));
    layer1_outputs(11021) <= (layer0_outputs(1024)) xor (layer0_outputs(2762));
    layer1_outputs(11022) <= (layer0_outputs(6175)) or (layer0_outputs(3690));
    layer1_outputs(11023) <= (layer0_outputs(9086)) xor (layer0_outputs(11705));
    layer1_outputs(11024) <= layer0_outputs(11260);
    layer1_outputs(11025) <= '1';
    layer1_outputs(11026) <= not(layer0_outputs(10781));
    layer1_outputs(11027) <= (layer0_outputs(11949)) and not (layer0_outputs(5670));
    layer1_outputs(11028) <= (layer0_outputs(3510)) or (layer0_outputs(6532));
    layer1_outputs(11029) <= not(layer0_outputs(3463));
    layer1_outputs(11030) <= layer0_outputs(10772);
    layer1_outputs(11031) <= not((layer0_outputs(223)) and (layer0_outputs(2350)));
    layer1_outputs(11032) <= not((layer0_outputs(955)) xor (layer0_outputs(10386)));
    layer1_outputs(11033) <= not(layer0_outputs(3523));
    layer1_outputs(11034) <= (layer0_outputs(1403)) and (layer0_outputs(6839));
    layer1_outputs(11035) <= (layer0_outputs(7980)) and not (layer0_outputs(5240));
    layer1_outputs(11036) <= not((layer0_outputs(1374)) and (layer0_outputs(7398)));
    layer1_outputs(11037) <= not(layer0_outputs(339));
    layer1_outputs(11038) <= not(layer0_outputs(3818));
    layer1_outputs(11039) <= '1';
    layer1_outputs(11040) <= not(layer0_outputs(6469));
    layer1_outputs(11041) <= not(layer0_outputs(6338));
    layer1_outputs(11042) <= (layer0_outputs(11684)) or (layer0_outputs(12310));
    layer1_outputs(11043) <= (layer0_outputs(5298)) xor (layer0_outputs(3520));
    layer1_outputs(11044) <= not(layer0_outputs(12705));
    layer1_outputs(11045) <= (layer0_outputs(1999)) and not (layer0_outputs(11515));
    layer1_outputs(11046) <= (layer0_outputs(4629)) and (layer0_outputs(11392));
    layer1_outputs(11047) <= (layer0_outputs(5942)) and not (layer0_outputs(6183));
    layer1_outputs(11048) <= not(layer0_outputs(872)) or (layer0_outputs(10239));
    layer1_outputs(11049) <= layer0_outputs(7615);
    layer1_outputs(11050) <= layer0_outputs(503);
    layer1_outputs(11051) <= layer0_outputs(4321);
    layer1_outputs(11052) <= layer0_outputs(6380);
    layer1_outputs(11053) <= not(layer0_outputs(2669));
    layer1_outputs(11054) <= layer0_outputs(12619);
    layer1_outputs(11055) <= not((layer0_outputs(8987)) and (layer0_outputs(5522)));
    layer1_outputs(11056) <= not(layer0_outputs(1799));
    layer1_outputs(11057) <= not(layer0_outputs(10866));
    layer1_outputs(11058) <= (layer0_outputs(4026)) xor (layer0_outputs(11716));
    layer1_outputs(11059) <= not((layer0_outputs(3149)) or (layer0_outputs(4284)));
    layer1_outputs(11060) <= not(layer0_outputs(1018));
    layer1_outputs(11061) <= (layer0_outputs(3696)) xor (layer0_outputs(6724));
    layer1_outputs(11062) <= not(layer0_outputs(6582));
    layer1_outputs(11063) <= (layer0_outputs(2522)) or (layer0_outputs(10017));
    layer1_outputs(11064) <= (layer0_outputs(2444)) xor (layer0_outputs(802));
    layer1_outputs(11065) <= not(layer0_outputs(1584)) or (layer0_outputs(551));
    layer1_outputs(11066) <= (layer0_outputs(8739)) and not (layer0_outputs(2508));
    layer1_outputs(11067) <= not(layer0_outputs(4536));
    layer1_outputs(11068) <= not((layer0_outputs(6616)) and (layer0_outputs(5259)));
    layer1_outputs(11069) <= not(layer0_outputs(11705)) or (layer0_outputs(5262));
    layer1_outputs(11070) <= (layer0_outputs(81)) xor (layer0_outputs(8058));
    layer1_outputs(11071) <= (layer0_outputs(3845)) and (layer0_outputs(6595));
    layer1_outputs(11072) <= not((layer0_outputs(6550)) and (layer0_outputs(7733)));
    layer1_outputs(11073) <= not(layer0_outputs(4263));
    layer1_outputs(11074) <= not((layer0_outputs(11324)) xor (layer0_outputs(9361)));
    layer1_outputs(11075) <= (layer0_outputs(3832)) xor (layer0_outputs(11397));
    layer1_outputs(11076) <= layer0_outputs(10806);
    layer1_outputs(11077) <= (layer0_outputs(3885)) xor (layer0_outputs(12531));
    layer1_outputs(11078) <= (layer0_outputs(6277)) xor (layer0_outputs(8829));
    layer1_outputs(11079) <= not(layer0_outputs(8996));
    layer1_outputs(11080) <= not(layer0_outputs(3145)) or (layer0_outputs(7789));
    layer1_outputs(11081) <= (layer0_outputs(8113)) and not (layer0_outputs(9236));
    layer1_outputs(11082) <= (layer0_outputs(11152)) and not (layer0_outputs(8645));
    layer1_outputs(11083) <= not(layer0_outputs(7135));
    layer1_outputs(11084) <= '1';
    layer1_outputs(11085) <= layer0_outputs(3231);
    layer1_outputs(11086) <= not((layer0_outputs(8275)) and (layer0_outputs(11665)));
    layer1_outputs(11087) <= (layer0_outputs(10435)) and not (layer0_outputs(9510));
    layer1_outputs(11088) <= not(layer0_outputs(11408)) or (layer0_outputs(3009));
    layer1_outputs(11089) <= not(layer0_outputs(1090));
    layer1_outputs(11090) <= (layer0_outputs(7760)) and not (layer0_outputs(5732));
    layer1_outputs(11091) <= (layer0_outputs(10461)) and not (layer0_outputs(3128));
    layer1_outputs(11092) <= (layer0_outputs(10141)) and not (layer0_outputs(7432));
    layer1_outputs(11093) <= layer0_outputs(2045);
    layer1_outputs(11094) <= layer0_outputs(11825);
    layer1_outputs(11095) <= (layer0_outputs(1350)) xor (layer0_outputs(5995));
    layer1_outputs(11096) <= layer0_outputs(2775);
    layer1_outputs(11097) <= (layer0_outputs(10247)) xor (layer0_outputs(2315));
    layer1_outputs(11098) <= not(layer0_outputs(3088)) or (layer0_outputs(68));
    layer1_outputs(11099) <= layer0_outputs(10399);
    layer1_outputs(11100) <= layer0_outputs(12285);
    layer1_outputs(11101) <= layer0_outputs(5523);
    layer1_outputs(11102) <= not(layer0_outputs(7072)) or (layer0_outputs(11975));
    layer1_outputs(11103) <= (layer0_outputs(7079)) and not (layer0_outputs(1737));
    layer1_outputs(11104) <= (layer0_outputs(2735)) xor (layer0_outputs(4002));
    layer1_outputs(11105) <= not(layer0_outputs(3501));
    layer1_outputs(11106) <= layer0_outputs(9888);
    layer1_outputs(11107) <= layer0_outputs(10241);
    layer1_outputs(11108) <= not((layer0_outputs(2541)) xor (layer0_outputs(3478)));
    layer1_outputs(11109) <= not(layer0_outputs(7624)) or (layer0_outputs(9622));
    layer1_outputs(11110) <= not(layer0_outputs(8642)) or (layer0_outputs(10638));
    layer1_outputs(11111) <= not(layer0_outputs(939)) or (layer0_outputs(1408));
    layer1_outputs(11112) <= not(layer0_outputs(10042)) or (layer0_outputs(318));
    layer1_outputs(11113) <= (layer0_outputs(8351)) and (layer0_outputs(719));
    layer1_outputs(11114) <= not((layer0_outputs(10107)) xor (layer0_outputs(7435)));
    layer1_outputs(11115) <= not((layer0_outputs(3897)) xor (layer0_outputs(11371)));
    layer1_outputs(11116) <= not((layer0_outputs(1691)) and (layer0_outputs(7880)));
    layer1_outputs(11117) <= not(layer0_outputs(10052));
    layer1_outputs(11118) <= not(layer0_outputs(5551));
    layer1_outputs(11119) <= not(layer0_outputs(8955)) or (layer0_outputs(1138));
    layer1_outputs(11120) <= not((layer0_outputs(6052)) or (layer0_outputs(8511)));
    layer1_outputs(11121) <= (layer0_outputs(8798)) and not (layer0_outputs(9436));
    layer1_outputs(11122) <= (layer0_outputs(3860)) and not (layer0_outputs(10513));
    layer1_outputs(11123) <= layer0_outputs(104);
    layer1_outputs(11124) <= not((layer0_outputs(2120)) xor (layer0_outputs(7069)));
    layer1_outputs(11125) <= layer0_outputs(9686);
    layer1_outputs(11126) <= layer0_outputs(9537);
    layer1_outputs(11127) <= (layer0_outputs(11257)) and not (layer0_outputs(9060));
    layer1_outputs(11128) <= (layer0_outputs(2771)) and (layer0_outputs(10168));
    layer1_outputs(11129) <= not((layer0_outputs(10208)) and (layer0_outputs(7741)));
    layer1_outputs(11130) <= not(layer0_outputs(2262));
    layer1_outputs(11131) <= layer0_outputs(6448);
    layer1_outputs(11132) <= not(layer0_outputs(12439)) or (layer0_outputs(11325));
    layer1_outputs(11133) <= (layer0_outputs(6044)) or (layer0_outputs(10690));
    layer1_outputs(11134) <= not((layer0_outputs(292)) or (layer0_outputs(6097)));
    layer1_outputs(11135) <= layer0_outputs(11239);
    layer1_outputs(11136) <= (layer0_outputs(11202)) and (layer0_outputs(9723));
    layer1_outputs(11137) <= not((layer0_outputs(4302)) or (layer0_outputs(8176)));
    layer1_outputs(11138) <= not(layer0_outputs(6279)) or (layer0_outputs(10805));
    layer1_outputs(11139) <= (layer0_outputs(8056)) xor (layer0_outputs(4719));
    layer1_outputs(11140) <= (layer0_outputs(6677)) or (layer0_outputs(9986));
    layer1_outputs(11141) <= not(layer0_outputs(7525));
    layer1_outputs(11142) <= not(layer0_outputs(8504));
    layer1_outputs(11143) <= layer0_outputs(10210);
    layer1_outputs(11144) <= not(layer0_outputs(6029));
    layer1_outputs(11145) <= layer0_outputs(1013);
    layer1_outputs(11146) <= not((layer0_outputs(4979)) and (layer0_outputs(1557)));
    layer1_outputs(11147) <= layer0_outputs(3893);
    layer1_outputs(11148) <= (layer0_outputs(5233)) and not (layer0_outputs(9961));
    layer1_outputs(11149) <= (layer0_outputs(1739)) and not (layer0_outputs(2297));
    layer1_outputs(11150) <= not(layer0_outputs(10003));
    layer1_outputs(11151) <= (layer0_outputs(4209)) and not (layer0_outputs(10150));
    layer1_outputs(11152) <= (layer0_outputs(11109)) and not (layer0_outputs(12742));
    layer1_outputs(11153) <= not(layer0_outputs(3665));
    layer1_outputs(11154) <= (layer0_outputs(7202)) xor (layer0_outputs(9507));
    layer1_outputs(11155) <= not((layer0_outputs(9062)) xor (layer0_outputs(7042)));
    layer1_outputs(11156) <= layer0_outputs(8373);
    layer1_outputs(11157) <= not(layer0_outputs(6053));
    layer1_outputs(11158) <= not(layer0_outputs(6324));
    layer1_outputs(11159) <= not(layer0_outputs(8615)) or (layer0_outputs(10457));
    layer1_outputs(11160) <= (layer0_outputs(4493)) and (layer0_outputs(524));
    layer1_outputs(11161) <= layer0_outputs(2019);
    layer1_outputs(11162) <= not((layer0_outputs(10117)) or (layer0_outputs(8966)));
    layer1_outputs(11163) <= not(layer0_outputs(1977)) or (layer0_outputs(1482));
    layer1_outputs(11164) <= layer0_outputs(2542);
    layer1_outputs(11165) <= (layer0_outputs(9258)) and not (layer0_outputs(4881));
    layer1_outputs(11166) <= not((layer0_outputs(7533)) and (layer0_outputs(43)));
    layer1_outputs(11167) <= not(layer0_outputs(12559));
    layer1_outputs(11168) <= (layer0_outputs(4755)) and not (layer0_outputs(10830));
    layer1_outputs(11169) <= (layer0_outputs(11509)) and not (layer0_outputs(2321));
    layer1_outputs(11170) <= (layer0_outputs(11264)) or (layer0_outputs(9002));
    layer1_outputs(11171) <= not((layer0_outputs(1425)) and (layer0_outputs(3158)));
    layer1_outputs(11172) <= layer0_outputs(4106);
    layer1_outputs(11173) <= layer0_outputs(9730);
    layer1_outputs(11174) <= not(layer0_outputs(8454));
    layer1_outputs(11175) <= (layer0_outputs(12628)) and not (layer0_outputs(7450));
    layer1_outputs(11176) <= not(layer0_outputs(5329));
    layer1_outputs(11177) <= not(layer0_outputs(1661)) or (layer0_outputs(9599));
    layer1_outputs(11178) <= not((layer0_outputs(12212)) xor (layer0_outputs(1482)));
    layer1_outputs(11179) <= not((layer0_outputs(6198)) and (layer0_outputs(9073)));
    layer1_outputs(11180) <= layer0_outputs(3386);
    layer1_outputs(11181) <= '1';
    layer1_outputs(11182) <= (layer0_outputs(270)) xor (layer0_outputs(1308));
    layer1_outputs(11183) <= not(layer0_outputs(11403)) or (layer0_outputs(10121));
    layer1_outputs(11184) <= (layer0_outputs(4130)) and not (layer0_outputs(9496));
    layer1_outputs(11185) <= not(layer0_outputs(3797));
    layer1_outputs(11186) <= not(layer0_outputs(4838)) or (layer0_outputs(9273));
    layer1_outputs(11187) <= not((layer0_outputs(1475)) xor (layer0_outputs(9224)));
    layer1_outputs(11188) <= layer0_outputs(1052);
    layer1_outputs(11189) <= layer0_outputs(3471);
    layer1_outputs(11190) <= (layer0_outputs(6381)) or (layer0_outputs(11523));
    layer1_outputs(11191) <= not((layer0_outputs(12616)) or (layer0_outputs(11181)));
    layer1_outputs(11192) <= '0';
    layer1_outputs(11193) <= '1';
    layer1_outputs(11194) <= not((layer0_outputs(173)) xor (layer0_outputs(7797)));
    layer1_outputs(11195) <= not((layer0_outputs(10928)) or (layer0_outputs(2467)));
    layer1_outputs(11196) <= layer0_outputs(10447);
    layer1_outputs(11197) <= not((layer0_outputs(3063)) xor (layer0_outputs(11920)));
    layer1_outputs(11198) <= layer0_outputs(804);
    layer1_outputs(11199) <= (layer0_outputs(11736)) xor (layer0_outputs(4278));
    layer1_outputs(11200) <= (layer0_outputs(12251)) xor (layer0_outputs(9398));
    layer1_outputs(11201) <= (layer0_outputs(5659)) and not (layer0_outputs(12284));
    layer1_outputs(11202) <= not(layer0_outputs(3533)) or (layer0_outputs(634));
    layer1_outputs(11203) <= layer0_outputs(5071);
    layer1_outputs(11204) <= not(layer0_outputs(7173));
    layer1_outputs(11205) <= (layer0_outputs(9971)) and (layer0_outputs(2821));
    layer1_outputs(11206) <= not(layer0_outputs(1747)) or (layer0_outputs(4221));
    layer1_outputs(11207) <= '0';
    layer1_outputs(11208) <= not(layer0_outputs(5430));
    layer1_outputs(11209) <= not((layer0_outputs(2236)) xor (layer0_outputs(12750)));
    layer1_outputs(11210) <= not(layer0_outputs(10425));
    layer1_outputs(11211) <= (layer0_outputs(3691)) or (layer0_outputs(4418));
    layer1_outputs(11212) <= not((layer0_outputs(12764)) or (layer0_outputs(10839)));
    layer1_outputs(11213) <= not((layer0_outputs(6511)) or (layer0_outputs(8686)));
    layer1_outputs(11214) <= (layer0_outputs(6471)) or (layer0_outputs(1092));
    layer1_outputs(11215) <= not(layer0_outputs(8360));
    layer1_outputs(11216) <= layer0_outputs(4243);
    layer1_outputs(11217) <= '0';
    layer1_outputs(11218) <= not((layer0_outputs(3693)) and (layer0_outputs(11613)));
    layer1_outputs(11219) <= (layer0_outputs(6183)) or (layer0_outputs(9225));
    layer1_outputs(11220) <= not((layer0_outputs(4076)) and (layer0_outputs(7795)));
    layer1_outputs(11221) <= layer0_outputs(1836);
    layer1_outputs(11222) <= layer0_outputs(1420);
    layer1_outputs(11223) <= (layer0_outputs(10849)) and not (layer0_outputs(1744));
    layer1_outputs(11224) <= (layer0_outputs(2436)) or (layer0_outputs(5954));
    layer1_outputs(11225) <= not(layer0_outputs(6510));
    layer1_outputs(11226) <= (layer0_outputs(4479)) and (layer0_outputs(11436));
    layer1_outputs(11227) <= not((layer0_outputs(9931)) xor (layer0_outputs(220)));
    layer1_outputs(11228) <= '1';
    layer1_outputs(11229) <= (layer0_outputs(10088)) or (layer0_outputs(5175));
    layer1_outputs(11230) <= (layer0_outputs(2863)) xor (layer0_outputs(4849));
    layer1_outputs(11231) <= not(layer0_outputs(4744));
    layer1_outputs(11232) <= (layer0_outputs(7333)) and not (layer0_outputs(7328));
    layer1_outputs(11233) <= not(layer0_outputs(8975)) or (layer0_outputs(12164));
    layer1_outputs(11234) <= not(layer0_outputs(2600));
    layer1_outputs(11235) <= not(layer0_outputs(3736));
    layer1_outputs(11236) <= (layer0_outputs(1142)) and not (layer0_outputs(4400));
    layer1_outputs(11237) <= not(layer0_outputs(430));
    layer1_outputs(11238) <= not(layer0_outputs(8756)) or (layer0_outputs(12677));
    layer1_outputs(11239) <= (layer0_outputs(10470)) and not (layer0_outputs(7572));
    layer1_outputs(11240) <= layer0_outputs(11760);
    layer1_outputs(11241) <= not(layer0_outputs(6296));
    layer1_outputs(11242) <= not((layer0_outputs(9483)) or (layer0_outputs(3925)));
    layer1_outputs(11243) <= layer0_outputs(9984);
    layer1_outputs(11244) <= not(layer0_outputs(4340)) or (layer0_outputs(1295));
    layer1_outputs(11245) <= not(layer0_outputs(7964)) or (layer0_outputs(8783));
    layer1_outputs(11246) <= not((layer0_outputs(7700)) and (layer0_outputs(7448)));
    layer1_outputs(11247) <= not((layer0_outputs(8258)) or (layer0_outputs(2947)));
    layer1_outputs(11248) <= (layer0_outputs(3042)) xor (layer0_outputs(3901));
    layer1_outputs(11249) <= not(layer0_outputs(2929));
    layer1_outputs(11250) <= not(layer0_outputs(8941));
    layer1_outputs(11251) <= layer0_outputs(11316);
    layer1_outputs(11252) <= not(layer0_outputs(4870)) or (layer0_outputs(9845));
    layer1_outputs(11253) <= layer0_outputs(8208);
    layer1_outputs(11254) <= (layer0_outputs(1003)) or (layer0_outputs(7790));
    layer1_outputs(11255) <= (layer0_outputs(3498)) and not (layer0_outputs(12059));
    layer1_outputs(11256) <= layer0_outputs(8775);
    layer1_outputs(11257) <= (layer0_outputs(5604)) and not (layer0_outputs(11772));
    layer1_outputs(11258) <= layer0_outputs(2008);
    layer1_outputs(11259) <= not((layer0_outputs(9779)) and (layer0_outputs(8726)));
    layer1_outputs(11260) <= '1';
    layer1_outputs(11261) <= '0';
    layer1_outputs(11262) <= '1';
    layer1_outputs(11263) <= '0';
    layer1_outputs(11264) <= not(layer0_outputs(4250));
    layer1_outputs(11265) <= (layer0_outputs(11638)) or (layer0_outputs(8140));
    layer1_outputs(11266) <= not(layer0_outputs(6796));
    layer1_outputs(11267) <= layer0_outputs(12006);
    layer1_outputs(11268) <= not(layer0_outputs(5827)) or (layer0_outputs(10232));
    layer1_outputs(11269) <= layer0_outputs(7385);
    layer1_outputs(11270) <= (layer0_outputs(2440)) xor (layer0_outputs(10831));
    layer1_outputs(11271) <= not((layer0_outputs(419)) and (layer0_outputs(2429)));
    layer1_outputs(11272) <= not(layer0_outputs(3171));
    layer1_outputs(11273) <= (layer0_outputs(2344)) or (layer0_outputs(8868));
    layer1_outputs(11274) <= not((layer0_outputs(4200)) and (layer0_outputs(8164)));
    layer1_outputs(11275) <= (layer0_outputs(11943)) and not (layer0_outputs(7452));
    layer1_outputs(11276) <= (layer0_outputs(5446)) and not (layer0_outputs(7514));
    layer1_outputs(11277) <= (layer0_outputs(1951)) or (layer0_outputs(386));
    layer1_outputs(11278) <= not(layer0_outputs(395)) or (layer0_outputs(3582));
    layer1_outputs(11279) <= not(layer0_outputs(1520));
    layer1_outputs(11280) <= not(layer0_outputs(3064));
    layer1_outputs(11281) <= layer0_outputs(8942);
    layer1_outputs(11282) <= (layer0_outputs(10675)) and not (layer0_outputs(6810));
    layer1_outputs(11283) <= not(layer0_outputs(2572));
    layer1_outputs(11284) <= (layer0_outputs(1512)) xor (layer0_outputs(11761));
    layer1_outputs(11285) <= (layer0_outputs(7029)) or (layer0_outputs(8251));
    layer1_outputs(11286) <= not(layer0_outputs(7706));
    layer1_outputs(11287) <= not((layer0_outputs(3827)) and (layer0_outputs(4870)));
    layer1_outputs(11288) <= '0';
    layer1_outputs(11289) <= not(layer0_outputs(12003));
    layer1_outputs(11290) <= (layer0_outputs(4426)) or (layer0_outputs(11866));
    layer1_outputs(11291) <= not((layer0_outputs(616)) or (layer0_outputs(980)));
    layer1_outputs(11292) <= layer0_outputs(10319);
    layer1_outputs(11293) <= (layer0_outputs(3272)) and not (layer0_outputs(4557));
    layer1_outputs(11294) <= not((layer0_outputs(6716)) and (layer0_outputs(5889)));
    layer1_outputs(11295) <= (layer0_outputs(3929)) and not (layer0_outputs(5805));
    layer1_outputs(11296) <= (layer0_outputs(8602)) xor (layer0_outputs(4024));
    layer1_outputs(11297) <= layer0_outputs(6331);
    layer1_outputs(11298) <= (layer0_outputs(6084)) xor (layer0_outputs(1128));
    layer1_outputs(11299) <= '1';
    layer1_outputs(11300) <= not(layer0_outputs(1463)) or (layer0_outputs(2098));
    layer1_outputs(11301) <= not((layer0_outputs(383)) or (layer0_outputs(12143)));
    layer1_outputs(11302) <= '0';
    layer1_outputs(11303) <= not((layer0_outputs(8502)) xor (layer0_outputs(7850)));
    layer1_outputs(11304) <= (layer0_outputs(555)) or (layer0_outputs(10339));
    layer1_outputs(11305) <= (layer0_outputs(1118)) and not (layer0_outputs(3267));
    layer1_outputs(11306) <= not((layer0_outputs(7265)) and (layer0_outputs(8576)));
    layer1_outputs(11307) <= layer0_outputs(12216);
    layer1_outputs(11308) <= not((layer0_outputs(10858)) xor (layer0_outputs(10161)));
    layer1_outputs(11309) <= not((layer0_outputs(10704)) and (layer0_outputs(11078)));
    layer1_outputs(11310) <= not(layer0_outputs(10677));
    layer1_outputs(11311) <= (layer0_outputs(12513)) or (layer0_outputs(6216));
    layer1_outputs(11312) <= not(layer0_outputs(236)) or (layer0_outputs(7103));
    layer1_outputs(11313) <= (layer0_outputs(3095)) and not (layer0_outputs(1934));
    layer1_outputs(11314) <= (layer0_outputs(3199)) xor (layer0_outputs(2230));
    layer1_outputs(11315) <= (layer0_outputs(3219)) and not (layer0_outputs(1602));
    layer1_outputs(11316) <= (layer0_outputs(10919)) and not (layer0_outputs(10891));
    layer1_outputs(11317) <= not((layer0_outputs(11721)) or (layer0_outputs(1751)));
    layer1_outputs(11318) <= not(layer0_outputs(2092)) or (layer0_outputs(6661));
    layer1_outputs(11319) <= not(layer0_outputs(11051));
    layer1_outputs(11320) <= not((layer0_outputs(6081)) xor (layer0_outputs(9732)));
    layer1_outputs(11321) <= not(layer0_outputs(2129));
    layer1_outputs(11322) <= not(layer0_outputs(10749));
    layer1_outputs(11323) <= not((layer0_outputs(6849)) xor (layer0_outputs(8095)));
    layer1_outputs(11324) <= (layer0_outputs(3436)) xor (layer0_outputs(11275));
    layer1_outputs(11325) <= not(layer0_outputs(10954));
    layer1_outputs(11326) <= not(layer0_outputs(1235)) or (layer0_outputs(4185));
    layer1_outputs(11327) <= not(layer0_outputs(11011)) or (layer0_outputs(4947));
    layer1_outputs(11328) <= not(layer0_outputs(11980));
    layer1_outputs(11329) <= not((layer0_outputs(5961)) and (layer0_outputs(12588)));
    layer1_outputs(11330) <= layer0_outputs(9499);
    layer1_outputs(11331) <= (layer0_outputs(4148)) and not (layer0_outputs(9475));
    layer1_outputs(11332) <= not((layer0_outputs(9980)) or (layer0_outputs(3528)));
    layer1_outputs(11333) <= layer0_outputs(11887);
    layer1_outputs(11334) <= not(layer0_outputs(9776)) or (layer0_outputs(1078));
    layer1_outputs(11335) <= not((layer0_outputs(6405)) and (layer0_outputs(9655)));
    layer1_outputs(11336) <= (layer0_outputs(9061)) and not (layer0_outputs(1956));
    layer1_outputs(11337) <= not(layer0_outputs(2953));
    layer1_outputs(11338) <= (layer0_outputs(8455)) or (layer0_outputs(4014));
    layer1_outputs(11339) <= (layer0_outputs(6192)) and not (layer0_outputs(4463));
    layer1_outputs(11340) <= (layer0_outputs(2487)) and (layer0_outputs(11095));
    layer1_outputs(11341) <= layer0_outputs(5951);
    layer1_outputs(11342) <= layer0_outputs(8287);
    layer1_outputs(11343) <= (layer0_outputs(23)) and not (layer0_outputs(7753));
    layer1_outputs(11344) <= (layer0_outputs(8365)) and not (layer0_outputs(4312));
    layer1_outputs(11345) <= not((layer0_outputs(4131)) and (layer0_outputs(5536)));
    layer1_outputs(11346) <= layer0_outputs(3635);
    layer1_outputs(11347) <= not((layer0_outputs(4568)) or (layer0_outputs(8226)));
    layer1_outputs(11348) <= not(layer0_outputs(8230));
    layer1_outputs(11349) <= layer0_outputs(4796);
    layer1_outputs(11350) <= not(layer0_outputs(3331));
    layer1_outputs(11351) <= layer0_outputs(6989);
    layer1_outputs(11352) <= (layer0_outputs(1238)) or (layer0_outputs(8316));
    layer1_outputs(11353) <= not((layer0_outputs(9404)) and (layer0_outputs(4827)));
    layer1_outputs(11354) <= not((layer0_outputs(7436)) and (layer0_outputs(8069)));
    layer1_outputs(11355) <= not(layer0_outputs(7393));
    layer1_outputs(11356) <= not(layer0_outputs(301));
    layer1_outputs(11357) <= (layer0_outputs(10001)) xor (layer0_outputs(333));
    layer1_outputs(11358) <= (layer0_outputs(10038)) and not (layer0_outputs(5965));
    layer1_outputs(11359) <= layer0_outputs(10380);
    layer1_outputs(11360) <= not(layer0_outputs(2801));
    layer1_outputs(11361) <= not(layer0_outputs(738));
    layer1_outputs(11362) <= (layer0_outputs(9891)) xor (layer0_outputs(9965));
    layer1_outputs(11363) <= not((layer0_outputs(8406)) or (layer0_outputs(3817)));
    layer1_outputs(11364) <= layer0_outputs(6222);
    layer1_outputs(11365) <= '1';
    layer1_outputs(11366) <= (layer0_outputs(10651)) and not (layer0_outputs(4634));
    layer1_outputs(11367) <= (layer0_outputs(10643)) xor (layer0_outputs(9454));
    layer1_outputs(11368) <= (layer0_outputs(12473)) or (layer0_outputs(10925));
    layer1_outputs(11369) <= layer0_outputs(3318);
    layer1_outputs(11370) <= (layer0_outputs(11227)) and not (layer0_outputs(5130));
    layer1_outputs(11371) <= (layer0_outputs(10690)) xor (layer0_outputs(7221));
    layer1_outputs(11372) <= layer0_outputs(4510);
    layer1_outputs(11373) <= (layer0_outputs(4981)) xor (layer0_outputs(12116));
    layer1_outputs(11374) <= not(layer0_outputs(10614));
    layer1_outputs(11375) <= not(layer0_outputs(5886));
    layer1_outputs(11376) <= layer0_outputs(4260);
    layer1_outputs(11377) <= layer0_outputs(7125);
    layer1_outputs(11378) <= not(layer0_outputs(6922)) or (layer0_outputs(2890));
    layer1_outputs(11379) <= not(layer0_outputs(4083));
    layer1_outputs(11380) <= not(layer0_outputs(8066)) or (layer0_outputs(9168));
    layer1_outputs(11381) <= layer0_outputs(1822);
    layer1_outputs(11382) <= not(layer0_outputs(1567)) or (layer0_outputs(8500));
    layer1_outputs(11383) <= not((layer0_outputs(5606)) and (layer0_outputs(4128)));
    layer1_outputs(11384) <= (layer0_outputs(560)) and not (layer0_outputs(7551));
    layer1_outputs(11385) <= not(layer0_outputs(11027)) or (layer0_outputs(1974));
    layer1_outputs(11386) <= (layer0_outputs(6916)) and not (layer0_outputs(8978));
    layer1_outputs(11387) <= not(layer0_outputs(267)) or (layer0_outputs(10351));
    layer1_outputs(11388) <= (layer0_outputs(4319)) and not (layer0_outputs(8571));
    layer1_outputs(11389) <= '0';
    layer1_outputs(11390) <= (layer0_outputs(531)) and not (layer0_outputs(3594));
    layer1_outputs(11391) <= not((layer0_outputs(3846)) and (layer0_outputs(6253)));
    layer1_outputs(11392) <= not((layer0_outputs(6117)) or (layer0_outputs(3983)));
    layer1_outputs(11393) <= (layer0_outputs(4273)) or (layer0_outputs(6344));
    layer1_outputs(11394) <= layer0_outputs(8296);
    layer1_outputs(11395) <= '0';
    layer1_outputs(11396) <= not(layer0_outputs(6831));
    layer1_outputs(11397) <= (layer0_outputs(214)) and not (layer0_outputs(3083));
    layer1_outputs(11398) <= not((layer0_outputs(6174)) and (layer0_outputs(10801)));
    layer1_outputs(11399) <= layer0_outputs(12474);
    layer1_outputs(11400) <= (layer0_outputs(684)) and (layer0_outputs(8414));
    layer1_outputs(11401) <= layer0_outputs(11076);
    layer1_outputs(11402) <= (layer0_outputs(4757)) or (layer0_outputs(3366));
    layer1_outputs(11403) <= not((layer0_outputs(9176)) and (layer0_outputs(10044)));
    layer1_outputs(11404) <= layer0_outputs(7439);
    layer1_outputs(11405) <= not(layer0_outputs(1982));
    layer1_outputs(11406) <= '0';
    layer1_outputs(11407) <= layer0_outputs(8492);
    layer1_outputs(11408) <= not(layer0_outputs(8171)) or (layer0_outputs(12676));
    layer1_outputs(11409) <= not(layer0_outputs(11410)) or (layer0_outputs(11046));
    layer1_outputs(11410) <= not(layer0_outputs(7681));
    layer1_outputs(11411) <= layer0_outputs(5531);
    layer1_outputs(11412) <= (layer0_outputs(312)) and not (layer0_outputs(7570));
    layer1_outputs(11413) <= not(layer0_outputs(11181)) or (layer0_outputs(3790));
    layer1_outputs(11414) <= (layer0_outputs(216)) and not (layer0_outputs(4129));
    layer1_outputs(11415) <= not(layer0_outputs(8011)) or (layer0_outputs(3507));
    layer1_outputs(11416) <= (layer0_outputs(11569)) and not (layer0_outputs(12434));
    layer1_outputs(11417) <= not((layer0_outputs(6970)) xor (layer0_outputs(5481)));
    layer1_outputs(11418) <= (layer0_outputs(4601)) or (layer0_outputs(11628));
    layer1_outputs(11419) <= (layer0_outputs(3213)) and not (layer0_outputs(3470));
    layer1_outputs(11420) <= layer0_outputs(12114);
    layer1_outputs(11421) <= layer0_outputs(588);
    layer1_outputs(11422) <= not(layer0_outputs(2831));
    layer1_outputs(11423) <= (layer0_outputs(2300)) or (layer0_outputs(5709));
    layer1_outputs(11424) <= layer0_outputs(3079);
    layer1_outputs(11425) <= not(layer0_outputs(2573));
    layer1_outputs(11426) <= layer0_outputs(10157);
    layer1_outputs(11427) <= not((layer0_outputs(10336)) xor (layer0_outputs(4445)));
    layer1_outputs(11428) <= layer0_outputs(1219);
    layer1_outputs(11429) <= (layer0_outputs(143)) and not (layer0_outputs(11273));
    layer1_outputs(11430) <= layer0_outputs(4610);
    layer1_outputs(11431) <= not(layer0_outputs(7111)) or (layer0_outputs(12243));
    layer1_outputs(11432) <= (layer0_outputs(2899)) or (layer0_outputs(1453));
    layer1_outputs(11433) <= '0';
    layer1_outputs(11434) <= (layer0_outputs(11670)) and not (layer0_outputs(9875));
    layer1_outputs(11435) <= (layer0_outputs(3049)) and not (layer0_outputs(11349));
    layer1_outputs(11436) <= '1';
    layer1_outputs(11437) <= not(layer0_outputs(10455)) or (layer0_outputs(5064));
    layer1_outputs(11438) <= (layer0_outputs(4471)) xor (layer0_outputs(12342));
    layer1_outputs(11439) <= layer0_outputs(2562);
    layer1_outputs(11440) <= (layer0_outputs(10025)) and (layer0_outputs(5927));
    layer1_outputs(11441) <= layer0_outputs(2429);
    layer1_outputs(11442) <= layer0_outputs(752);
    layer1_outputs(11443) <= not((layer0_outputs(1234)) and (layer0_outputs(832)));
    layer1_outputs(11444) <= not(layer0_outputs(3548));
    layer1_outputs(11445) <= not(layer0_outputs(5107)) or (layer0_outputs(10670));
    layer1_outputs(11446) <= layer0_outputs(11972);
    layer1_outputs(11447) <= not(layer0_outputs(7168));
    layer1_outputs(11448) <= not(layer0_outputs(2547));
    layer1_outputs(11449) <= not(layer0_outputs(2425));
    layer1_outputs(11450) <= not(layer0_outputs(11506)) or (layer0_outputs(8787));
    layer1_outputs(11451) <= layer0_outputs(6105);
    layer1_outputs(11452) <= '0';
    layer1_outputs(11453) <= (layer0_outputs(6055)) and not (layer0_outputs(3961));
    layer1_outputs(11454) <= (layer0_outputs(10975)) and not (layer0_outputs(2918));
    layer1_outputs(11455) <= not(layer0_outputs(2529));
    layer1_outputs(11456) <= (layer0_outputs(4669)) or (layer0_outputs(6909));
    layer1_outputs(11457) <= '1';
    layer1_outputs(11458) <= (layer0_outputs(10046)) xor (layer0_outputs(3361));
    layer1_outputs(11459) <= not(layer0_outputs(11111));
    layer1_outputs(11460) <= not(layer0_outputs(1465)) or (layer0_outputs(10055));
    layer1_outputs(11461) <= not((layer0_outputs(11653)) or (layer0_outputs(5467)));
    layer1_outputs(11462) <= not((layer0_outputs(7673)) and (layer0_outputs(2940)));
    layer1_outputs(11463) <= not(layer0_outputs(1035)) or (layer0_outputs(7635));
    layer1_outputs(11464) <= (layer0_outputs(11983)) xor (layer0_outputs(8233));
    layer1_outputs(11465) <= not(layer0_outputs(10092));
    layer1_outputs(11466) <= (layer0_outputs(8116)) and not (layer0_outputs(4054));
    layer1_outputs(11467) <= not(layer0_outputs(7938)) or (layer0_outputs(12234));
    layer1_outputs(11468) <= not(layer0_outputs(6654));
    layer1_outputs(11469) <= (layer0_outputs(9319)) or (layer0_outputs(9084));
    layer1_outputs(11470) <= layer0_outputs(8976);
    layer1_outputs(11471) <= (layer0_outputs(4957)) and not (layer0_outputs(8862));
    layer1_outputs(11472) <= layer0_outputs(9572);
    layer1_outputs(11473) <= (layer0_outputs(4544)) xor (layer0_outputs(1862));
    layer1_outputs(11474) <= not(layer0_outputs(10800)) or (layer0_outputs(153));
    layer1_outputs(11475) <= not((layer0_outputs(12196)) xor (layer0_outputs(9294)));
    layer1_outputs(11476) <= layer0_outputs(5589);
    layer1_outputs(11477) <= layer0_outputs(6242);
    layer1_outputs(11478) <= layer0_outputs(1249);
    layer1_outputs(11479) <= (layer0_outputs(11723)) xor (layer0_outputs(8301));
    layer1_outputs(11480) <= not(layer0_outputs(6253));
    layer1_outputs(11481) <= not(layer0_outputs(922)) or (layer0_outputs(9950));
    layer1_outputs(11482) <= layer0_outputs(7658);
    layer1_outputs(11483) <= layer0_outputs(786);
    layer1_outputs(11484) <= (layer0_outputs(10879)) xor (layer0_outputs(9930));
    layer1_outputs(11485) <= (layer0_outputs(1042)) xor (layer0_outputs(8323));
    layer1_outputs(11486) <= not((layer0_outputs(4210)) and (layer0_outputs(8101)));
    layer1_outputs(11487) <= layer0_outputs(2410);
    layer1_outputs(11488) <= not(layer0_outputs(7147)) or (layer0_outputs(11614));
    layer1_outputs(11489) <= layer0_outputs(2517);
    layer1_outputs(11490) <= not((layer0_outputs(5802)) xor (layer0_outputs(2951)));
    layer1_outputs(11491) <= not(layer0_outputs(12075));
    layer1_outputs(11492) <= (layer0_outputs(9962)) and not (layer0_outputs(7745));
    layer1_outputs(11493) <= not(layer0_outputs(6764)) or (layer0_outputs(982));
    layer1_outputs(11494) <= not(layer0_outputs(4447));
    layer1_outputs(11495) <= not((layer0_outputs(1659)) xor (layer0_outputs(12687)));
    layer1_outputs(11496) <= (layer0_outputs(11782)) xor (layer0_outputs(467));
    layer1_outputs(11497) <= (layer0_outputs(1057)) and not (layer0_outputs(7331));
    layer1_outputs(11498) <= not(layer0_outputs(11234));
    layer1_outputs(11499) <= layer0_outputs(11354);
    layer1_outputs(11500) <= layer0_outputs(6234);
    layer1_outputs(11501) <= not((layer0_outputs(334)) xor (layer0_outputs(5498)));
    layer1_outputs(11502) <= not(layer0_outputs(7755)) or (layer0_outputs(835));
    layer1_outputs(11503) <= not(layer0_outputs(7489));
    layer1_outputs(11504) <= not(layer0_outputs(2738)) or (layer0_outputs(2989));
    layer1_outputs(11505) <= layer0_outputs(11382);
    layer1_outputs(11506) <= layer0_outputs(12291);
    layer1_outputs(11507) <= not(layer0_outputs(7062));
    layer1_outputs(11508) <= layer0_outputs(6670);
    layer1_outputs(11509) <= not(layer0_outputs(12378));
    layer1_outputs(11510) <= not((layer0_outputs(11293)) and (layer0_outputs(6370)));
    layer1_outputs(11511) <= (layer0_outputs(12764)) and not (layer0_outputs(3557));
    layer1_outputs(11512) <= (layer0_outputs(1157)) and (layer0_outputs(9918));
    layer1_outputs(11513) <= (layer0_outputs(12490)) xor (layer0_outputs(2314));
    layer1_outputs(11514) <= not(layer0_outputs(305)) or (layer0_outputs(9154));
    layer1_outputs(11515) <= (layer0_outputs(6509)) and not (layer0_outputs(12552));
    layer1_outputs(11516) <= layer0_outputs(7800);
    layer1_outputs(11517) <= '1';
    layer1_outputs(11518) <= '0';
    layer1_outputs(11519) <= (layer0_outputs(9698)) and not (layer0_outputs(11563));
    layer1_outputs(11520) <= layer0_outputs(2578);
    layer1_outputs(11521) <= not(layer0_outputs(1554));
    layer1_outputs(11522) <= (layer0_outputs(12033)) or (layer0_outputs(2304));
    layer1_outputs(11523) <= (layer0_outputs(4385)) and not (layer0_outputs(2527));
    layer1_outputs(11524) <= not((layer0_outputs(9668)) xor (layer0_outputs(1838)));
    layer1_outputs(11525) <= not(layer0_outputs(8359));
    layer1_outputs(11526) <= layer0_outputs(3323);
    layer1_outputs(11527) <= not(layer0_outputs(2195));
    layer1_outputs(11528) <= layer0_outputs(6064);
    layer1_outputs(11529) <= (layer0_outputs(1431)) or (layer0_outputs(7303));
    layer1_outputs(11530) <= (layer0_outputs(9808)) and not (layer0_outputs(859));
    layer1_outputs(11531) <= not(layer0_outputs(8389));
    layer1_outputs(11532) <= (layer0_outputs(2911)) or (layer0_outputs(5947));
    layer1_outputs(11533) <= not((layer0_outputs(810)) and (layer0_outputs(514)));
    layer1_outputs(11534) <= not(layer0_outputs(615)) or (layer0_outputs(2976));
    layer1_outputs(11535) <= not((layer0_outputs(1272)) and (layer0_outputs(12488)));
    layer1_outputs(11536) <= not((layer0_outputs(5736)) xor (layer0_outputs(5543)));
    layer1_outputs(11537) <= not((layer0_outputs(12732)) and (layer0_outputs(8444)));
    layer1_outputs(11538) <= not(layer0_outputs(8709));
    layer1_outputs(11539) <= not(layer0_outputs(9907)) or (layer0_outputs(9009));
    layer1_outputs(11540) <= not(layer0_outputs(169)) or (layer0_outputs(4000));
    layer1_outputs(11541) <= not(layer0_outputs(2830));
    layer1_outputs(11542) <= not((layer0_outputs(1684)) and (layer0_outputs(7182)));
    layer1_outputs(11543) <= layer0_outputs(9920);
    layer1_outputs(11544) <= not(layer0_outputs(7003)) or (layer0_outputs(9939));
    layer1_outputs(11545) <= not((layer0_outputs(320)) or (layer0_outputs(11780)));
    layer1_outputs(11546) <= layer0_outputs(7256);
    layer1_outputs(11547) <= not(layer0_outputs(8165));
    layer1_outputs(11548) <= layer0_outputs(669);
    layer1_outputs(11549) <= not((layer0_outputs(6009)) and (layer0_outputs(4966)));
    layer1_outputs(11550) <= not(layer0_outputs(5393));
    layer1_outputs(11551) <= not(layer0_outputs(5073));
    layer1_outputs(11552) <= not(layer0_outputs(8654));
    layer1_outputs(11553) <= not(layer0_outputs(4553));
    layer1_outputs(11554) <= (layer0_outputs(1745)) and not (layer0_outputs(9206));
    layer1_outputs(11555) <= layer0_outputs(6456);
    layer1_outputs(11556) <= not((layer0_outputs(1435)) xor (layer0_outputs(1970)));
    layer1_outputs(11557) <= not(layer0_outputs(5356)) or (layer0_outputs(9917));
    layer1_outputs(11558) <= (layer0_outputs(4181)) xor (layer0_outputs(6065));
    layer1_outputs(11559) <= not(layer0_outputs(4872));
    layer1_outputs(11560) <= layer0_outputs(11811);
    layer1_outputs(11561) <= not((layer0_outputs(3913)) and (layer0_outputs(1785)));
    layer1_outputs(11562) <= layer0_outputs(7404);
    layer1_outputs(11563) <= (layer0_outputs(4500)) or (layer0_outputs(8944));
    layer1_outputs(11564) <= not(layer0_outputs(1409));
    layer1_outputs(11565) <= (layer0_outputs(879)) or (layer0_outputs(3808));
    layer1_outputs(11566) <= (layer0_outputs(2221)) xor (layer0_outputs(7802));
    layer1_outputs(11567) <= (layer0_outputs(885)) and not (layer0_outputs(10061));
    layer1_outputs(11568) <= layer0_outputs(3303);
    layer1_outputs(11569) <= not((layer0_outputs(1558)) or (layer0_outputs(11732)));
    layer1_outputs(11570) <= not(layer0_outputs(1915)) or (layer0_outputs(12198));
    layer1_outputs(11571) <= not((layer0_outputs(6374)) or (layer0_outputs(8419)));
    layer1_outputs(11572) <= layer0_outputs(5881);
    layer1_outputs(11573) <= '0';
    layer1_outputs(11574) <= layer0_outputs(5482);
    layer1_outputs(11575) <= not((layer0_outputs(85)) xor (layer0_outputs(7789)));
    layer1_outputs(11576) <= layer0_outputs(7475);
    layer1_outputs(11577) <= (layer0_outputs(7150)) and (layer0_outputs(7973));
    layer1_outputs(11578) <= layer0_outputs(6113);
    layer1_outputs(11579) <= (layer0_outputs(10165)) or (layer0_outputs(11084));
    layer1_outputs(11580) <= layer0_outputs(6785);
    layer1_outputs(11581) <= (layer0_outputs(9330)) and (layer0_outputs(11293));
    layer1_outputs(11582) <= not((layer0_outputs(3933)) and (layer0_outputs(1714)));
    layer1_outputs(11583) <= not(layer0_outputs(5119));
    layer1_outputs(11584) <= not(layer0_outputs(7946));
    layer1_outputs(11585) <= (layer0_outputs(3545)) xor (layer0_outputs(5549));
    layer1_outputs(11586) <= (layer0_outputs(9721)) and (layer0_outputs(4118));
    layer1_outputs(11587) <= not((layer0_outputs(5979)) or (layer0_outputs(5660)));
    layer1_outputs(11588) <= layer0_outputs(929);
    layer1_outputs(11589) <= not(layer0_outputs(12555)) or (layer0_outputs(10671));
    layer1_outputs(11590) <= layer0_outputs(11408);
    layer1_outputs(11591) <= not(layer0_outputs(2076));
    layer1_outputs(11592) <= not((layer0_outputs(953)) or (layer0_outputs(7921)));
    layer1_outputs(11593) <= layer0_outputs(1696);
    layer1_outputs(11594) <= (layer0_outputs(4970)) and (layer0_outputs(12399));
    layer1_outputs(11595) <= not(layer0_outputs(1762));
    layer1_outputs(11596) <= (layer0_outputs(9272)) or (layer0_outputs(3966));
    layer1_outputs(11597) <= (layer0_outputs(10624)) xor (layer0_outputs(5943));
    layer1_outputs(11598) <= '0';
    layer1_outputs(11599) <= not((layer0_outputs(6074)) and (layer0_outputs(9484)));
    layer1_outputs(11600) <= (layer0_outputs(7242)) xor (layer0_outputs(10799));
    layer1_outputs(11601) <= (layer0_outputs(12532)) and (layer0_outputs(7793));
    layer1_outputs(11602) <= not((layer0_outputs(5463)) and (layer0_outputs(5592)));
    layer1_outputs(11603) <= layer0_outputs(3697);
    layer1_outputs(11604) <= not(layer0_outputs(3856)) or (layer0_outputs(5472));
    layer1_outputs(11605) <= (layer0_outputs(9503)) xor (layer0_outputs(8062));
    layer1_outputs(11606) <= (layer0_outputs(6102)) and not (layer0_outputs(2386));
    layer1_outputs(11607) <= (layer0_outputs(132)) and not (layer0_outputs(2585));
    layer1_outputs(11608) <= layer0_outputs(10492);
    layer1_outputs(11609) <= not((layer0_outputs(5695)) xor (layer0_outputs(4305)));
    layer1_outputs(11610) <= (layer0_outputs(10646)) and not (layer0_outputs(9581));
    layer1_outputs(11611) <= not(layer0_outputs(4404));
    layer1_outputs(11612) <= layer0_outputs(7346);
    layer1_outputs(11613) <= (layer0_outputs(12046)) xor (layer0_outputs(372));
    layer1_outputs(11614) <= (layer0_outputs(7314)) xor (layer0_outputs(12345));
    layer1_outputs(11615) <= not((layer0_outputs(5100)) xor (layer0_outputs(3063)));
    layer1_outputs(11616) <= layer0_outputs(1183);
    layer1_outputs(11617) <= (layer0_outputs(12671)) and not (layer0_outputs(6509));
    layer1_outputs(11618) <= not(layer0_outputs(3241));
    layer1_outputs(11619) <= not(layer0_outputs(8119));
    layer1_outputs(11620) <= not(layer0_outputs(10885));
    layer1_outputs(11621) <= (layer0_outputs(11089)) and not (layer0_outputs(6604));
    layer1_outputs(11622) <= not((layer0_outputs(1591)) and (layer0_outputs(233)));
    layer1_outputs(11623) <= not(layer0_outputs(10124));
    layer1_outputs(11624) <= not(layer0_outputs(709));
    layer1_outputs(11625) <= not((layer0_outputs(9489)) xor (layer0_outputs(10421)));
    layer1_outputs(11626) <= layer0_outputs(9079);
    layer1_outputs(11627) <= not((layer0_outputs(6692)) and (layer0_outputs(2053)));
    layer1_outputs(11628) <= layer0_outputs(4811);
    layer1_outputs(11629) <= layer0_outputs(11661);
    layer1_outputs(11630) <= not(layer0_outputs(6313));
    layer1_outputs(11631) <= layer0_outputs(8267);
    layer1_outputs(11632) <= layer0_outputs(1748);
    layer1_outputs(11633) <= (layer0_outputs(8723)) and not (layer0_outputs(4334));
    layer1_outputs(11634) <= (layer0_outputs(8918)) and not (layer0_outputs(11484));
    layer1_outputs(11635) <= not((layer0_outputs(6296)) or (layer0_outputs(6089)));
    layer1_outputs(11636) <= not(layer0_outputs(1795));
    layer1_outputs(11637) <= (layer0_outputs(3259)) and (layer0_outputs(5403));
    layer1_outputs(11638) <= (layer0_outputs(10266)) and not (layer0_outputs(8449));
    layer1_outputs(11639) <= layer0_outputs(3518);
    layer1_outputs(11640) <= not((layer0_outputs(4596)) xor (layer0_outputs(2733)));
    layer1_outputs(11641) <= (layer0_outputs(8147)) or (layer0_outputs(8963));
    layer1_outputs(11642) <= layer0_outputs(5978);
    layer1_outputs(11643) <= not(layer0_outputs(7459));
    layer1_outputs(11644) <= not(layer0_outputs(5199));
    layer1_outputs(11645) <= layer0_outputs(5789);
    layer1_outputs(11646) <= not((layer0_outputs(11396)) xor (layer0_outputs(4719)));
    layer1_outputs(11647) <= '0';
    layer1_outputs(11648) <= not(layer0_outputs(6392)) or (layer0_outputs(4511));
    layer1_outputs(11649) <= not(layer0_outputs(2157));
    layer1_outputs(11650) <= not(layer0_outputs(6457));
    layer1_outputs(11651) <= layer0_outputs(10406);
    layer1_outputs(11652) <= not((layer0_outputs(2337)) or (layer0_outputs(1551)));
    layer1_outputs(11653) <= not(layer0_outputs(3245));
    layer1_outputs(11654) <= not(layer0_outputs(14));
    layer1_outputs(11655) <= not(layer0_outputs(258));
    layer1_outputs(11656) <= not((layer0_outputs(343)) and (layer0_outputs(2689)));
    layer1_outputs(11657) <= not(layer0_outputs(2694));
    layer1_outputs(11658) <= not((layer0_outputs(11026)) xor (layer0_outputs(11422)));
    layer1_outputs(11659) <= layer0_outputs(1858);
    layer1_outputs(11660) <= layer0_outputs(1703);
    layer1_outputs(11661) <= not((layer0_outputs(5707)) and (layer0_outputs(4961)));
    layer1_outputs(11662) <= (layer0_outputs(8856)) xor (layer0_outputs(6982));
    layer1_outputs(11663) <= not(layer0_outputs(12042));
    layer1_outputs(11664) <= not(layer0_outputs(11579));
    layer1_outputs(11665) <= not((layer0_outputs(3777)) xor (layer0_outputs(12773)));
    layer1_outputs(11666) <= not(layer0_outputs(2771));
    layer1_outputs(11667) <= not(layer0_outputs(5365));
    layer1_outputs(11668) <= not(layer0_outputs(4935)) or (layer0_outputs(5343));
    layer1_outputs(11669) <= layer0_outputs(1421);
    layer1_outputs(11670) <= (layer0_outputs(12458)) and not (layer0_outputs(8878));
    layer1_outputs(11671) <= not((layer0_outputs(4626)) and (layer0_outputs(974)));
    layer1_outputs(11672) <= layer0_outputs(756);
    layer1_outputs(11673) <= not(layer0_outputs(1474));
    layer1_outputs(11674) <= layer0_outputs(2959);
    layer1_outputs(11675) <= layer0_outputs(11929);
    layer1_outputs(11676) <= layer0_outputs(1917);
    layer1_outputs(11677) <= not((layer0_outputs(7862)) or (layer0_outputs(2581)));
    layer1_outputs(11678) <= (layer0_outputs(9431)) and (layer0_outputs(1824));
    layer1_outputs(11679) <= not(layer0_outputs(141)) or (layer0_outputs(727));
    layer1_outputs(11680) <= not(layer0_outputs(2498));
    layer1_outputs(11681) <= (layer0_outputs(9588)) and (layer0_outputs(8169));
    layer1_outputs(11682) <= layer0_outputs(6747);
    layer1_outputs(11683) <= not((layer0_outputs(9131)) xor (layer0_outputs(2636)));
    layer1_outputs(11684) <= not(layer0_outputs(3850));
    layer1_outputs(11685) <= not((layer0_outputs(9227)) and (layer0_outputs(12250)));
    layer1_outputs(11686) <= (layer0_outputs(12450)) and not (layer0_outputs(8358));
    layer1_outputs(11687) <= not((layer0_outputs(10250)) and (layer0_outputs(9287)));
    layer1_outputs(11688) <= layer0_outputs(12036);
    layer1_outputs(11689) <= not(layer0_outputs(5285));
    layer1_outputs(11690) <= layer0_outputs(12551);
    layer1_outputs(11691) <= not(layer0_outputs(5311));
    layer1_outputs(11692) <= (layer0_outputs(2735)) or (layer0_outputs(2012));
    layer1_outputs(11693) <= layer0_outputs(8306);
    layer1_outputs(11694) <= not((layer0_outputs(4179)) xor (layer0_outputs(7351)));
    layer1_outputs(11695) <= (layer0_outputs(5245)) and (layer0_outputs(6421));
    layer1_outputs(11696) <= not(layer0_outputs(1597)) or (layer0_outputs(4750));
    layer1_outputs(11697) <= layer0_outputs(10495);
    layer1_outputs(11698) <= not(layer0_outputs(6309)) or (layer0_outputs(7833));
    layer1_outputs(11699) <= (layer0_outputs(4867)) or (layer0_outputs(5668));
    layer1_outputs(11700) <= (layer0_outputs(3896)) or (layer0_outputs(616));
    layer1_outputs(11701) <= not(layer0_outputs(1367));
    layer1_outputs(11702) <= layer0_outputs(12082);
    layer1_outputs(11703) <= not(layer0_outputs(9375));
    layer1_outputs(11704) <= not(layer0_outputs(9046)) or (layer0_outputs(2204));
    layer1_outputs(11705) <= not(layer0_outputs(11351));
    layer1_outputs(11706) <= layer0_outputs(7777);
    layer1_outputs(11707) <= not(layer0_outputs(455));
    layer1_outputs(11708) <= not(layer0_outputs(7356));
    layer1_outputs(11709) <= layer0_outputs(9760);
    layer1_outputs(11710) <= (layer0_outputs(11725)) and not (layer0_outputs(5380));
    layer1_outputs(11711) <= not(layer0_outputs(5786));
    layer1_outputs(11712) <= layer0_outputs(10965);
    layer1_outputs(11713) <= (layer0_outputs(9237)) and not (layer0_outputs(8617));
    layer1_outputs(11714) <= layer0_outputs(11641);
    layer1_outputs(11715) <= (layer0_outputs(8232)) xor (layer0_outputs(6712));
    layer1_outputs(11716) <= not((layer0_outputs(9897)) xor (layer0_outputs(9048)));
    layer1_outputs(11717) <= not(layer0_outputs(5366));
    layer1_outputs(11718) <= (layer0_outputs(6850)) and not (layer0_outputs(4227));
    layer1_outputs(11719) <= layer0_outputs(3334);
    layer1_outputs(11720) <= (layer0_outputs(5215)) and not (layer0_outputs(5541));
    layer1_outputs(11721) <= not(layer0_outputs(1597)) or (layer0_outputs(7817));
    layer1_outputs(11722) <= not((layer0_outputs(12402)) or (layer0_outputs(808)));
    layer1_outputs(11723) <= not(layer0_outputs(10511));
    layer1_outputs(11724) <= (layer0_outputs(3766)) and (layer0_outputs(2601));
    layer1_outputs(11725) <= layer0_outputs(2619);
    layer1_outputs(11726) <= (layer0_outputs(11416)) and not (layer0_outputs(3464));
    layer1_outputs(11727) <= layer0_outputs(4311);
    layer1_outputs(11728) <= (layer0_outputs(3522)) and not (layer0_outputs(8828));
    layer1_outputs(11729) <= layer0_outputs(12673);
    layer1_outputs(11730) <= (layer0_outputs(2279)) and (layer0_outputs(2834));
    layer1_outputs(11731) <= not(layer0_outputs(2589));
    layer1_outputs(11732) <= not(layer0_outputs(7232)) or (layer0_outputs(1114));
    layer1_outputs(11733) <= not((layer0_outputs(1137)) and (layer0_outputs(7022)));
    layer1_outputs(11734) <= not(layer0_outputs(3838)) or (layer0_outputs(1783));
    layer1_outputs(11735) <= not(layer0_outputs(1764)) or (layer0_outputs(8998));
    layer1_outputs(11736) <= layer0_outputs(10329);
    layer1_outputs(11737) <= not(layer0_outputs(3129)) or (layer0_outputs(876));
    layer1_outputs(11738) <= (layer0_outputs(11859)) or (layer0_outputs(4368));
    layer1_outputs(11739) <= not((layer0_outputs(4008)) xor (layer0_outputs(4721)));
    layer1_outputs(11740) <= (layer0_outputs(3315)) xor (layer0_outputs(8545));
    layer1_outputs(11741) <= (layer0_outputs(8578)) and (layer0_outputs(12333));
    layer1_outputs(11742) <= not((layer0_outputs(373)) xor (layer0_outputs(6804)));
    layer1_outputs(11743) <= (layer0_outputs(1351)) and not (layer0_outputs(8442));
    layer1_outputs(11744) <= not(layer0_outputs(8741));
    layer1_outputs(11745) <= layer0_outputs(4963);
    layer1_outputs(11746) <= (layer0_outputs(9251)) and not (layer0_outputs(5609));
    layer1_outputs(11747) <= not(layer0_outputs(3430)) or (layer0_outputs(3454));
    layer1_outputs(11748) <= layer0_outputs(8567);
    layer1_outputs(11749) <= not((layer0_outputs(12785)) xor (layer0_outputs(7744)));
    layer1_outputs(11750) <= (layer0_outputs(5173)) and (layer0_outputs(3605));
    layer1_outputs(11751) <= not(layer0_outputs(7407));
    layer1_outputs(11752) <= layer0_outputs(215);
    layer1_outputs(11753) <= not(layer0_outputs(8441)) or (layer0_outputs(5852));
    layer1_outputs(11754) <= not(layer0_outputs(6211));
    layer1_outputs(11755) <= not(layer0_outputs(9360)) or (layer0_outputs(7689));
    layer1_outputs(11756) <= not(layer0_outputs(10537)) or (layer0_outputs(3056));
    layer1_outputs(11757) <= not((layer0_outputs(2836)) xor (layer0_outputs(11576)));
    layer1_outputs(11758) <= not((layer0_outputs(2151)) or (layer0_outputs(6097)));
    layer1_outputs(11759) <= (layer0_outputs(1976)) and (layer0_outputs(2736));
    layer1_outputs(11760) <= '1';
    layer1_outputs(11761) <= not(layer0_outputs(11906)) or (layer0_outputs(6258));
    layer1_outputs(11762) <= layer0_outputs(3457);
    layer1_outputs(11763) <= not(layer0_outputs(3350));
    layer1_outputs(11764) <= layer0_outputs(11559);
    layer1_outputs(11765) <= not((layer0_outputs(5736)) and (layer0_outputs(86)));
    layer1_outputs(11766) <= not((layer0_outputs(1109)) xor (layer0_outputs(6077)));
    layer1_outputs(11767) <= layer0_outputs(10166);
    layer1_outputs(11768) <= not(layer0_outputs(4997));
    layer1_outputs(11769) <= not(layer0_outputs(5547)) or (layer0_outputs(7279));
    layer1_outputs(11770) <= not(layer0_outputs(9341));
    layer1_outputs(11771) <= not((layer0_outputs(8554)) or (layer0_outputs(7839)));
    layer1_outputs(11772) <= not(layer0_outputs(2805));
    layer1_outputs(11773) <= (layer0_outputs(6925)) and not (layer0_outputs(2796));
    layer1_outputs(11774) <= layer0_outputs(4975);
    layer1_outputs(11775) <= layer0_outputs(272);
    layer1_outputs(11776) <= layer0_outputs(10522);
    layer1_outputs(11777) <= '0';
    layer1_outputs(11778) <= (layer0_outputs(4556)) xor (layer0_outputs(4018));
    layer1_outputs(11779) <= layer0_outputs(7286);
    layer1_outputs(11780) <= not(layer0_outputs(7167)) or (layer0_outputs(2290));
    layer1_outputs(11781) <= layer0_outputs(9634);
    layer1_outputs(11782) <= (layer0_outputs(2763)) and not (layer0_outputs(10419));
    layer1_outputs(11783) <= not(layer0_outputs(11401));
    layer1_outputs(11784) <= (layer0_outputs(1254)) and not (layer0_outputs(346));
    layer1_outputs(11785) <= (layer0_outputs(11428)) xor (layer0_outputs(8885));
    layer1_outputs(11786) <= (layer0_outputs(8356)) and not (layer0_outputs(3457));
    layer1_outputs(11787) <= not(layer0_outputs(4675));
    layer1_outputs(11788) <= layer0_outputs(5008);
    layer1_outputs(11789) <= (layer0_outputs(10105)) and (layer0_outputs(64));
    layer1_outputs(11790) <= (layer0_outputs(4834)) or (layer0_outputs(12385));
    layer1_outputs(11791) <= not((layer0_outputs(7647)) xor (layer0_outputs(8573)));
    layer1_outputs(11792) <= (layer0_outputs(6318)) xor (layer0_outputs(11327));
    layer1_outputs(11793) <= (layer0_outputs(6226)) and not (layer0_outputs(4806));
    layer1_outputs(11794) <= (layer0_outputs(9974)) or (layer0_outputs(1925));
    layer1_outputs(11795) <= '1';
    layer1_outputs(11796) <= not((layer0_outputs(3054)) and (layer0_outputs(11021)));
    layer1_outputs(11797) <= layer0_outputs(6440);
    layer1_outputs(11798) <= (layer0_outputs(18)) and (layer0_outputs(8271));
    layer1_outputs(11799) <= layer0_outputs(4731);
    layer1_outputs(11800) <= not((layer0_outputs(8811)) or (layer0_outputs(5811)));
    layer1_outputs(11801) <= not(layer0_outputs(2033));
    layer1_outputs(11802) <= (layer0_outputs(7502)) or (layer0_outputs(8830));
    layer1_outputs(11803) <= not(layer0_outputs(7403));
    layer1_outputs(11804) <= layer0_outputs(1989);
    layer1_outputs(11805) <= (layer0_outputs(2857)) xor (layer0_outputs(122));
    layer1_outputs(11806) <= layer0_outputs(2228);
    layer1_outputs(11807) <= layer0_outputs(6271);
    layer1_outputs(11808) <= not((layer0_outputs(7199)) or (layer0_outputs(11653)));
    layer1_outputs(11809) <= layer0_outputs(12222);
    layer1_outputs(11810) <= not(layer0_outputs(11347));
    layer1_outputs(11811) <= not(layer0_outputs(9153)) or (layer0_outputs(2207));
    layer1_outputs(11812) <= not(layer0_outputs(6667)) or (layer0_outputs(2714));
    layer1_outputs(11813) <= layer0_outputs(7);
    layer1_outputs(11814) <= not((layer0_outputs(4405)) or (layer0_outputs(8281)));
    layer1_outputs(11815) <= (layer0_outputs(8467)) and not (layer0_outputs(10693));
    layer1_outputs(11816) <= not(layer0_outputs(9803)) or (layer0_outputs(4074));
    layer1_outputs(11817) <= not(layer0_outputs(7931));
    layer1_outputs(11818) <= not((layer0_outputs(3308)) xor (layer0_outputs(3871)));
    layer1_outputs(11819) <= not(layer0_outputs(9388));
    layer1_outputs(11820) <= (layer0_outputs(9270)) and not (layer0_outputs(10627));
    layer1_outputs(11821) <= not(layer0_outputs(803)) or (layer0_outputs(10332));
    layer1_outputs(11822) <= (layer0_outputs(1080)) or (layer0_outputs(3381));
    layer1_outputs(11823) <= layer0_outputs(4639);
    layer1_outputs(11824) <= not((layer0_outputs(9034)) or (layer0_outputs(309)));
    layer1_outputs(11825) <= (layer0_outputs(10669)) and not (layer0_outputs(2139));
    layer1_outputs(11826) <= (layer0_outputs(8764)) and not (layer0_outputs(6508));
    layer1_outputs(11827) <= layer0_outputs(5353);
    layer1_outputs(11828) <= layer0_outputs(225);
    layer1_outputs(11829) <= not((layer0_outputs(6150)) xor (layer0_outputs(11377)));
    layer1_outputs(11830) <= not(layer0_outputs(11976)) or (layer0_outputs(8779));
    layer1_outputs(11831) <= not(layer0_outputs(4595)) or (layer0_outputs(7482));
    layer1_outputs(11832) <= (layer0_outputs(12034)) and not (layer0_outputs(2734));
    layer1_outputs(11833) <= (layer0_outputs(10378)) and not (layer0_outputs(547));
    layer1_outputs(11834) <= not((layer0_outputs(548)) or (layer0_outputs(10108)));
    layer1_outputs(11835) <= '1';
    layer1_outputs(11836) <= not((layer0_outputs(4978)) or (layer0_outputs(12301)));
    layer1_outputs(11837) <= (layer0_outputs(114)) or (layer0_outputs(3679));
    layer1_outputs(11838) <= (layer0_outputs(6346)) and (layer0_outputs(9045));
    layer1_outputs(11839) <= (layer0_outputs(2519)) and not (layer0_outputs(10539));
    layer1_outputs(11840) <= not((layer0_outputs(10118)) or (layer0_outputs(1162)));
    layer1_outputs(11841) <= not((layer0_outputs(12541)) or (layer0_outputs(12408)));
    layer1_outputs(11842) <= not(layer0_outputs(4351)) or (layer0_outputs(2228));
    layer1_outputs(11843) <= not((layer0_outputs(6387)) and (layer0_outputs(8366)));
    layer1_outputs(11844) <= layer0_outputs(5015);
    layer1_outputs(11845) <= not((layer0_outputs(6233)) and (layer0_outputs(10510)));
    layer1_outputs(11846) <= not(layer0_outputs(11333));
    layer1_outputs(11847) <= layer0_outputs(5374);
    layer1_outputs(11848) <= layer0_outputs(2178);
    layer1_outputs(11849) <= (layer0_outputs(8407)) and not (layer0_outputs(8476));
    layer1_outputs(11850) <= (layer0_outputs(9384)) or (layer0_outputs(6567));
    layer1_outputs(11851) <= not(layer0_outputs(6175));
    layer1_outputs(11852) <= not((layer0_outputs(7760)) xor (layer0_outputs(5993)));
    layer1_outputs(11853) <= (layer0_outputs(4846)) and not (layer0_outputs(5621));
    layer1_outputs(11854) <= not((layer0_outputs(4502)) or (layer0_outputs(9028)));
    layer1_outputs(11855) <= not((layer0_outputs(7402)) and (layer0_outputs(6723)));
    layer1_outputs(11856) <= (layer0_outputs(6310)) or (layer0_outputs(10566));
    layer1_outputs(11857) <= not((layer0_outputs(4555)) and (layer0_outputs(5428)));
    layer1_outputs(11858) <= not(layer0_outputs(12175)) or (layer0_outputs(6783));
    layer1_outputs(11859) <= not(layer0_outputs(8951));
    layer1_outputs(11860) <= not((layer0_outputs(541)) or (layer0_outputs(3410)));
    layer1_outputs(11861) <= not((layer0_outputs(7074)) xor (layer0_outputs(1998)));
    layer1_outputs(11862) <= not((layer0_outputs(8905)) or (layer0_outputs(7559)));
    layer1_outputs(11863) <= (layer0_outputs(2710)) and (layer0_outputs(10715));
    layer1_outputs(11864) <= not(layer0_outputs(4080));
    layer1_outputs(11865) <= layer0_outputs(886);
    layer1_outputs(11866) <= (layer0_outputs(12062)) xor (layer0_outputs(6683));
    layer1_outputs(11867) <= not(layer0_outputs(712)) or (layer0_outputs(7780));
    layer1_outputs(11868) <= not(layer0_outputs(11060)) or (layer0_outputs(11670));
    layer1_outputs(11869) <= not((layer0_outputs(10997)) xor (layer0_outputs(8137)));
    layer1_outputs(11870) <= not(layer0_outputs(231)) or (layer0_outputs(2181));
    layer1_outputs(11871) <= (layer0_outputs(12172)) and (layer0_outputs(12152));
    layer1_outputs(11872) <= (layer0_outputs(3987)) or (layer0_outputs(10819));
    layer1_outputs(11873) <= (layer0_outputs(7530)) and not (layer0_outputs(1876));
    layer1_outputs(11874) <= layer0_outputs(634);
    layer1_outputs(11875) <= not((layer0_outputs(6597)) xor (layer0_outputs(5618)));
    layer1_outputs(11876) <= (layer0_outputs(3106)) or (layer0_outputs(5127));
    layer1_outputs(11877) <= not(layer0_outputs(296));
    layer1_outputs(11878) <= not(layer0_outputs(4603)) or (layer0_outputs(9580));
    layer1_outputs(11879) <= not((layer0_outputs(3022)) or (layer0_outputs(1452)));
    layer1_outputs(11880) <= not(layer0_outputs(9493));
    layer1_outputs(11881) <= not((layer0_outputs(3731)) and (layer0_outputs(3408)));
    layer1_outputs(11882) <= not(layer0_outputs(4286));
    layer1_outputs(11883) <= not(layer0_outputs(7413));
    layer1_outputs(11884) <= layer0_outputs(4316);
    layer1_outputs(11885) <= not(layer0_outputs(9433));
    layer1_outputs(11886) <= layer0_outputs(8815);
    layer1_outputs(11887) <= not((layer0_outputs(6972)) or (layer0_outputs(3754)));
    layer1_outputs(11888) <= layer0_outputs(11996);
    layer1_outputs(11889) <= not(layer0_outputs(11513));
    layer1_outputs(11890) <= layer0_outputs(7806);
    layer1_outputs(11891) <= not(layer0_outputs(4741)) or (layer0_outputs(6847));
    layer1_outputs(11892) <= (layer0_outputs(9927)) or (layer0_outputs(829));
    layer1_outputs(11893) <= not((layer0_outputs(6850)) xor (layer0_outputs(4584)));
    layer1_outputs(11894) <= (layer0_outputs(10691)) xor (layer0_outputs(546));
    layer1_outputs(11895) <= layer0_outputs(8515);
    layer1_outputs(11896) <= not(layer0_outputs(8410));
    layer1_outputs(11897) <= (layer0_outputs(5810)) or (layer0_outputs(5124));
    layer1_outputs(11898) <= (layer0_outputs(2356)) and not (layer0_outputs(5599));
    layer1_outputs(11899) <= (layer0_outputs(952)) and (layer0_outputs(8782));
    layer1_outputs(11900) <= (layer0_outputs(125)) and not (layer0_outputs(2435));
    layer1_outputs(11901) <= layer0_outputs(469);
    layer1_outputs(11902) <= layer0_outputs(11284);
    layer1_outputs(11903) <= not((layer0_outputs(8221)) and (layer0_outputs(79)));
    layer1_outputs(11904) <= layer0_outputs(1281);
    layer1_outputs(11905) <= not(layer0_outputs(10159));
    layer1_outputs(11906) <= not(layer0_outputs(4891));
    layer1_outputs(11907) <= not((layer0_outputs(12341)) or (layer0_outputs(9374)));
    layer1_outputs(11908) <= (layer0_outputs(8706)) and (layer0_outputs(12160));
    layer1_outputs(11909) <= (layer0_outputs(5968)) and not (layer0_outputs(5532));
    layer1_outputs(11910) <= not(layer0_outputs(940));
    layer1_outputs(11911) <= not(layer0_outputs(845));
    layer1_outputs(11912) <= not((layer0_outputs(7865)) or (layer0_outputs(6173)));
    layer1_outputs(11913) <= not(layer0_outputs(499));
    layer1_outputs(11914) <= layer0_outputs(11844);
    layer1_outputs(11915) <= (layer0_outputs(3449)) and not (layer0_outputs(1665));
    layer1_outputs(11916) <= layer0_outputs(10745);
    layer1_outputs(11917) <= not(layer0_outputs(9532));
    layer1_outputs(11918) <= not((layer0_outputs(3312)) xor (layer0_outputs(2089)));
    layer1_outputs(11919) <= not(layer0_outputs(9458));
    layer1_outputs(11920) <= not(layer0_outputs(4720)) or (layer0_outputs(6074));
    layer1_outputs(11921) <= not((layer0_outputs(9519)) and (layer0_outputs(1593)));
    layer1_outputs(11922) <= (layer0_outputs(6177)) and not (layer0_outputs(7367));
    layer1_outputs(11923) <= not(layer0_outputs(12524));
    layer1_outputs(11924) <= not(layer0_outputs(135)) or (layer0_outputs(8524));
    layer1_outputs(11925) <= layer0_outputs(2659);
    layer1_outputs(11926) <= (layer0_outputs(6389)) xor (layer0_outputs(3907));
    layer1_outputs(11927) <= not(layer0_outputs(827));
    layer1_outputs(11928) <= not(layer0_outputs(11754));
    layer1_outputs(11929) <= not((layer0_outputs(11475)) xor (layer0_outputs(5471)));
    layer1_outputs(11930) <= not(layer0_outputs(3354)) or (layer0_outputs(2134));
    layer1_outputs(11931) <= not(layer0_outputs(10032));
    layer1_outputs(11932) <= (layer0_outputs(5849)) xor (layer0_outputs(9138));
    layer1_outputs(11933) <= not(layer0_outputs(5919));
    layer1_outputs(11934) <= (layer0_outputs(465)) and not (layer0_outputs(7852));
    layer1_outputs(11935) <= not(layer0_outputs(1759)) or (layer0_outputs(8604));
    layer1_outputs(11936) <= '1';
    layer1_outputs(11937) <= not(layer0_outputs(4178));
    layer1_outputs(11938) <= not((layer0_outputs(7631)) and (layer0_outputs(12763)));
    layer1_outputs(11939) <= not((layer0_outputs(12114)) and (layer0_outputs(11114)));
    layer1_outputs(11940) <= not(layer0_outputs(6195));
    layer1_outputs(11941) <= (layer0_outputs(1477)) and not (layer0_outputs(8520));
    layer1_outputs(11942) <= not((layer0_outputs(1919)) and (layer0_outputs(11470)));
    layer1_outputs(11943) <= not(layer0_outputs(393));
    layer1_outputs(11944) <= layer0_outputs(10912);
    layer1_outputs(11945) <= (layer0_outputs(2269)) and not (layer0_outputs(8009));
    layer1_outputs(11946) <= layer0_outputs(2510);
    layer1_outputs(11947) <= (layer0_outputs(9587)) and not (layer0_outputs(7493));
    layer1_outputs(11948) <= not(layer0_outputs(3733));
    layer1_outputs(11949) <= layer0_outputs(8540);
    layer1_outputs(11950) <= not((layer0_outputs(9728)) or (layer0_outputs(3835)));
    layer1_outputs(11951) <= (layer0_outputs(469)) and not (layer0_outputs(1000));
    layer1_outputs(11952) <= (layer0_outputs(2449)) and not (layer0_outputs(4935));
    layer1_outputs(11953) <= layer0_outputs(11610);
    layer1_outputs(11954) <= (layer0_outputs(4732)) or (layer0_outputs(1047));
    layer1_outputs(11955) <= (layer0_outputs(11212)) and not (layer0_outputs(4635));
    layer1_outputs(11956) <= (layer0_outputs(1393)) and not (layer0_outputs(5331));
    layer1_outputs(11957) <= not((layer0_outputs(301)) or (layer0_outputs(7464)));
    layer1_outputs(11958) <= not(layer0_outputs(1169)) or (layer0_outputs(5435));
    layer1_outputs(11959) <= not(layer0_outputs(4251)) or (layer0_outputs(7656));
    layer1_outputs(11960) <= layer0_outputs(5558);
    layer1_outputs(11961) <= '0';
    layer1_outputs(11962) <= layer0_outputs(8403);
    layer1_outputs(11963) <= not(layer0_outputs(11688)) or (layer0_outputs(6685));
    layer1_outputs(11964) <= layer0_outputs(9414);
    layer1_outputs(11965) <= not(layer0_outputs(3981)) or (layer0_outputs(4012));
    layer1_outputs(11966) <= (layer0_outputs(771)) and not (layer0_outputs(8755));
    layer1_outputs(11967) <= layer0_outputs(11734);
    layer1_outputs(11968) <= not((layer0_outputs(735)) or (layer0_outputs(2895)));
    layer1_outputs(11969) <= not((layer0_outputs(1766)) or (layer0_outputs(5272)));
    layer1_outputs(11970) <= not(layer0_outputs(5672));
    layer1_outputs(11971) <= not((layer0_outputs(3926)) and (layer0_outputs(6352)));
    layer1_outputs(11972) <= (layer0_outputs(4677)) xor (layer0_outputs(156));
    layer1_outputs(11973) <= (layer0_outputs(5229)) and not (layer0_outputs(3570));
    layer1_outputs(11974) <= layer0_outputs(4504);
    layer1_outputs(11975) <= not((layer0_outputs(9077)) and (layer0_outputs(1565)));
    layer1_outputs(11976) <= not(layer0_outputs(12526));
    layer1_outputs(11977) <= layer0_outputs(1014);
    layer1_outputs(11978) <= not(layer0_outputs(6277));
    layer1_outputs(11979) <= layer0_outputs(7189);
    layer1_outputs(11980) <= layer0_outputs(1510);
    layer1_outputs(11981) <= layer0_outputs(12633);
    layer1_outputs(11982) <= not((layer0_outputs(3730)) or (layer0_outputs(5874)));
    layer1_outputs(11983) <= (layer0_outputs(3730)) or (layer0_outputs(9575));
    layer1_outputs(11984) <= (layer0_outputs(3497)) or (layer0_outputs(3993));
    layer1_outputs(11985) <= (layer0_outputs(1735)) and not (layer0_outputs(4708));
    layer1_outputs(11986) <= (layer0_outputs(2093)) and not (layer0_outputs(10642));
    layer1_outputs(11987) <= (layer0_outputs(3650)) and not (layer0_outputs(10826));
    layer1_outputs(11988) <= not((layer0_outputs(1922)) or (layer0_outputs(7627)));
    layer1_outputs(11989) <= layer0_outputs(9752);
    layer1_outputs(11990) <= not(layer0_outputs(9818)) or (layer0_outputs(2679));
    layer1_outputs(11991) <= not(layer0_outputs(11615));
    layer1_outputs(11992) <= not(layer0_outputs(10473)) or (layer0_outputs(10344));
    layer1_outputs(11993) <= not(layer0_outputs(279));
    layer1_outputs(11994) <= not(layer0_outputs(5403));
    layer1_outputs(11995) <= (layer0_outputs(11718)) and not (layer0_outputs(9119));
    layer1_outputs(11996) <= (layer0_outputs(5450)) and (layer0_outputs(1613));
    layer1_outputs(11997) <= (layer0_outputs(11846)) and (layer0_outputs(10661));
    layer1_outputs(11998) <= (layer0_outputs(9588)) and not (layer0_outputs(4885));
    layer1_outputs(11999) <= layer0_outputs(6967);
    layer1_outputs(12000) <= (layer0_outputs(7416)) and (layer0_outputs(719));
    layer1_outputs(12001) <= (layer0_outputs(12292)) and (layer0_outputs(5394));
    layer1_outputs(12002) <= not(layer0_outputs(12446));
    layer1_outputs(12003) <= (layer0_outputs(8556)) or (layer0_outputs(12439));
    layer1_outputs(12004) <= (layer0_outputs(12514)) and not (layer0_outputs(5513));
    layer1_outputs(12005) <= not((layer0_outputs(5507)) and (layer0_outputs(720)));
    layer1_outputs(12006) <= (layer0_outputs(12607)) xor (layer0_outputs(9853));
    layer1_outputs(12007) <= '1';
    layer1_outputs(12008) <= not(layer0_outputs(12477));
    layer1_outputs(12009) <= (layer0_outputs(10537)) and (layer0_outputs(806));
    layer1_outputs(12010) <= (layer0_outputs(6281)) xor (layer0_outputs(4917));
    layer1_outputs(12011) <= not(layer0_outputs(11240)) or (layer0_outputs(9738));
    layer1_outputs(12012) <= not((layer0_outputs(11521)) and (layer0_outputs(3027)));
    layer1_outputs(12013) <= not(layer0_outputs(10485));
    layer1_outputs(12014) <= not(layer0_outputs(6348));
    layer1_outputs(12015) <= not((layer0_outputs(8481)) or (layer0_outputs(7450)));
    layer1_outputs(12016) <= (layer0_outputs(4950)) or (layer0_outputs(7109));
    layer1_outputs(12017) <= (layer0_outputs(9661)) and not (layer0_outputs(11973));
    layer1_outputs(12018) <= not(layer0_outputs(6339));
    layer1_outputs(12019) <= not(layer0_outputs(11759)) or (layer0_outputs(10709));
    layer1_outputs(12020) <= not(layer0_outputs(3545)) or (layer0_outputs(2039));
    layer1_outputs(12021) <= not((layer0_outputs(536)) and (layer0_outputs(4120)));
    layer1_outputs(12022) <= '1';
    layer1_outputs(12023) <= layer0_outputs(1588);
    layer1_outputs(12024) <= not(layer0_outputs(12395));
    layer1_outputs(12025) <= not(layer0_outputs(4451));
    layer1_outputs(12026) <= not(layer0_outputs(7332));
    layer1_outputs(12027) <= not(layer0_outputs(10733));
    layer1_outputs(12028) <= '0';
    layer1_outputs(12029) <= layer0_outputs(12685);
    layer1_outputs(12030) <= (layer0_outputs(1354)) and not (layer0_outputs(12217));
    layer1_outputs(12031) <= not(layer0_outputs(11251));
    layer1_outputs(12032) <= (layer0_outputs(1545)) and not (layer0_outputs(6586));
    layer1_outputs(12033) <= (layer0_outputs(9495)) and not (layer0_outputs(9229));
    layer1_outputs(12034) <= layer0_outputs(9285);
    layer1_outputs(12035) <= layer0_outputs(12565);
    layer1_outputs(12036) <= layer0_outputs(2580);
    layer1_outputs(12037) <= (layer0_outputs(5334)) and not (layer0_outputs(6802));
    layer1_outputs(12038) <= (layer0_outputs(1616)) and not (layer0_outputs(7371));
    layer1_outputs(12039) <= (layer0_outputs(7611)) and (layer0_outputs(636));
    layer1_outputs(12040) <= (layer0_outputs(10133)) and not (layer0_outputs(10856));
    layer1_outputs(12041) <= layer0_outputs(3918);
    layer1_outputs(12042) <= not(layer0_outputs(881));
    layer1_outputs(12043) <= layer0_outputs(1135);
    layer1_outputs(12044) <= not(layer0_outputs(3406)) or (layer0_outputs(9831));
    layer1_outputs(12045) <= (layer0_outputs(517)) and not (layer0_outputs(5573));
    layer1_outputs(12046) <= (layer0_outputs(10388)) or (layer0_outputs(8936));
    layer1_outputs(12047) <= (layer0_outputs(3369)) and (layer0_outputs(11211));
    layer1_outputs(12048) <= not((layer0_outputs(7043)) and (layer0_outputs(9683)));
    layer1_outputs(12049) <= not(layer0_outputs(8750)) or (layer0_outputs(2501));
    layer1_outputs(12050) <= layer0_outputs(1094);
    layer1_outputs(12051) <= layer0_outputs(1372);
    layer1_outputs(12052) <= not(layer0_outputs(4804));
    layer1_outputs(12053) <= not((layer0_outputs(391)) or (layer0_outputs(5920)));
    layer1_outputs(12054) <= layer0_outputs(11789);
    layer1_outputs(12055) <= not(layer0_outputs(704));
    layer1_outputs(12056) <= not(layer0_outputs(11988));
    layer1_outputs(12057) <= not(layer0_outputs(12773));
    layer1_outputs(12058) <= not(layer0_outputs(8818));
    layer1_outputs(12059) <= not((layer0_outputs(2986)) and (layer0_outputs(509)));
    layer1_outputs(12060) <= not((layer0_outputs(11263)) xor (layer0_outputs(5238)));
    layer1_outputs(12061) <= layer0_outputs(10996);
    layer1_outputs(12062) <= not(layer0_outputs(3169)) or (layer0_outputs(11045));
    layer1_outputs(12063) <= not(layer0_outputs(2647));
    layer1_outputs(12064) <= not((layer0_outputs(8945)) and (layer0_outputs(7563)));
    layer1_outputs(12065) <= (layer0_outputs(2502)) or (layer0_outputs(6931));
    layer1_outputs(12066) <= (layer0_outputs(9710)) or (layer0_outputs(1538));
    layer1_outputs(12067) <= (layer0_outputs(5580)) and not (layer0_outputs(10049));
    layer1_outputs(12068) <= not((layer0_outputs(9814)) xor (layer0_outputs(11520)));
    layer1_outputs(12069) <= (layer0_outputs(25)) or (layer0_outputs(2917));
    layer1_outputs(12070) <= (layer0_outputs(4186)) xor (layer0_outputs(5141));
    layer1_outputs(12071) <= not(layer0_outputs(12140));
    layer1_outputs(12072) <= (layer0_outputs(4329)) and not (layer0_outputs(8130));
    layer1_outputs(12073) <= (layer0_outputs(6411)) or (layer0_outputs(10790));
    layer1_outputs(12074) <= (layer0_outputs(11782)) or (layer0_outputs(1470));
    layer1_outputs(12075) <= layer0_outputs(4398);
    layer1_outputs(12076) <= not(layer0_outputs(4516));
    layer1_outputs(12077) <= (layer0_outputs(362)) or (layer0_outputs(323));
    layer1_outputs(12078) <= (layer0_outputs(6734)) and (layer0_outputs(2941));
    layer1_outputs(12079) <= (layer0_outputs(6128)) xor (layer0_outputs(1159));
    layer1_outputs(12080) <= (layer0_outputs(3999)) xor (layer0_outputs(1651));
    layer1_outputs(12081) <= not(layer0_outputs(8201));
    layer1_outputs(12082) <= layer0_outputs(5940);
    layer1_outputs(12083) <= '1';
    layer1_outputs(12084) <= layer0_outputs(1869);
    layer1_outputs(12085) <= not((layer0_outputs(11346)) or (layer0_outputs(7814)));
    layer1_outputs(12086) <= layer0_outputs(11451);
    layer1_outputs(12087) <= not((layer0_outputs(12047)) xor (layer0_outputs(6101)));
    layer1_outputs(12088) <= not((layer0_outputs(314)) or (layer0_outputs(2101)));
    layer1_outputs(12089) <= not(layer0_outputs(11019)) or (layer0_outputs(2346));
    layer1_outputs(12090) <= (layer0_outputs(8937)) and not (layer0_outputs(7731));
    layer1_outputs(12091) <= '1';
    layer1_outputs(12092) <= (layer0_outputs(9566)) and not (layer0_outputs(760));
    layer1_outputs(12093) <= (layer0_outputs(11489)) and not (layer0_outputs(10110));
    layer1_outputs(12094) <= (layer0_outputs(5729)) and not (layer0_outputs(5715));
    layer1_outputs(12095) <= not((layer0_outputs(6630)) or (layer0_outputs(3224)));
    layer1_outputs(12096) <= layer0_outputs(8868);
    layer1_outputs(12097) <= not((layer0_outputs(2359)) or (layer0_outputs(7684)));
    layer1_outputs(12098) <= not(layer0_outputs(7329));
    layer1_outputs(12099) <= layer0_outputs(11173);
    layer1_outputs(12100) <= (layer0_outputs(482)) or (layer0_outputs(9063));
    layer1_outputs(12101) <= layer0_outputs(7078);
    layer1_outputs(12102) <= layer0_outputs(7788);
    layer1_outputs(12103) <= layer0_outputs(10734);
    layer1_outputs(12104) <= (layer0_outputs(1070)) or (layer0_outputs(5421));
    layer1_outputs(12105) <= layer0_outputs(7662);
    layer1_outputs(12106) <= (layer0_outputs(1533)) and not (layer0_outputs(5627));
    layer1_outputs(12107) <= layer0_outputs(5217);
    layer1_outputs(12108) <= (layer0_outputs(11350)) xor (layer0_outputs(10293));
    layer1_outputs(12109) <= layer0_outputs(6880);
    layer1_outputs(12110) <= not(layer0_outputs(1754)) or (layer0_outputs(7974));
    layer1_outputs(12111) <= (layer0_outputs(8533)) xor (layer0_outputs(9430));
    layer1_outputs(12112) <= '1';
    layer1_outputs(12113) <= not(layer0_outputs(8188));
    layer1_outputs(12114) <= (layer0_outputs(5038)) or (layer0_outputs(11015));
    layer1_outputs(12115) <= not(layer0_outputs(2034));
    layer1_outputs(12116) <= layer0_outputs(3241);
    layer1_outputs(12117) <= (layer0_outputs(5477)) and (layer0_outputs(5441));
    layer1_outputs(12118) <= not(layer0_outputs(8962));
    layer1_outputs(12119) <= not(layer0_outputs(4061)) or (layer0_outputs(4932));
    layer1_outputs(12120) <= not(layer0_outputs(12389));
    layer1_outputs(12121) <= not(layer0_outputs(10412));
    layer1_outputs(12122) <= layer0_outputs(4129);
    layer1_outputs(12123) <= not(layer0_outputs(4873));
    layer1_outputs(12124) <= not((layer0_outputs(12673)) xor (layer0_outputs(11581)));
    layer1_outputs(12125) <= not(layer0_outputs(8352));
    layer1_outputs(12126) <= (layer0_outputs(5184)) and (layer0_outputs(10647));
    layer1_outputs(12127) <= (layer0_outputs(7066)) and not (layer0_outputs(11492));
    layer1_outputs(12128) <= (layer0_outputs(4371)) or (layer0_outputs(5987));
    layer1_outputs(12129) <= layer0_outputs(2755);
    layer1_outputs(12130) <= (layer0_outputs(1780)) or (layer0_outputs(4889));
    layer1_outputs(12131) <= (layer0_outputs(6759)) and (layer0_outputs(8611));
    layer1_outputs(12132) <= (layer0_outputs(8063)) xor (layer0_outputs(11838));
    layer1_outputs(12133) <= layer0_outputs(1931);
    layer1_outputs(12134) <= not(layer0_outputs(12219)) or (layer0_outputs(7934));
    layer1_outputs(12135) <= (layer0_outputs(3221)) xor (layer0_outputs(2631));
    layer1_outputs(12136) <= not((layer0_outputs(2351)) and (layer0_outputs(6534)));
    layer1_outputs(12137) <= not(layer0_outputs(11650));
    layer1_outputs(12138) <= not((layer0_outputs(11953)) or (layer0_outputs(4996)));
    layer1_outputs(12139) <= layer0_outputs(1318);
    layer1_outputs(12140) <= not(layer0_outputs(12659));
    layer1_outputs(12141) <= not(layer0_outputs(9022));
    layer1_outputs(12142) <= not(layer0_outputs(4153));
    layer1_outputs(12143) <= not(layer0_outputs(8257)) or (layer0_outputs(4871));
    layer1_outputs(12144) <= not((layer0_outputs(3541)) xor (layer0_outputs(10110)));
    layer1_outputs(12145) <= layer0_outputs(783);
    layer1_outputs(12146) <= not((layer0_outputs(11885)) and (layer0_outputs(10688)));
    layer1_outputs(12147) <= (layer0_outputs(1330)) xor (layer0_outputs(11964));
    layer1_outputs(12148) <= (layer0_outputs(5492)) and not (layer0_outputs(6865));
    layer1_outputs(12149) <= layer0_outputs(7921);
    layer1_outputs(12150) <= (layer0_outputs(12163)) xor (layer0_outputs(10751));
    layer1_outputs(12151) <= not(layer0_outputs(7182)) or (layer0_outputs(961));
    layer1_outputs(12152) <= layer0_outputs(1969);
    layer1_outputs(12153) <= (layer0_outputs(6929)) and not (layer0_outputs(12376));
    layer1_outputs(12154) <= not((layer0_outputs(10378)) and (layer0_outputs(9893)));
    layer1_outputs(12155) <= not((layer0_outputs(10397)) and (layer0_outputs(3753)));
    layer1_outputs(12156) <= not(layer0_outputs(4016));
    layer1_outputs(12157) <= not(layer0_outputs(12580));
    layer1_outputs(12158) <= (layer0_outputs(12087)) xor (layer0_outputs(11010));
    layer1_outputs(12159) <= not(layer0_outputs(7904));
    layer1_outputs(12160) <= layer0_outputs(2768);
    layer1_outputs(12161) <= layer0_outputs(1621);
    layer1_outputs(12162) <= not((layer0_outputs(5065)) or (layer0_outputs(1667)));
    layer1_outputs(12163) <= (layer0_outputs(8684)) or (layer0_outputs(9176));
    layer1_outputs(12164) <= not(layer0_outputs(8219));
    layer1_outputs(12165) <= (layer0_outputs(6604)) and (layer0_outputs(10609));
    layer1_outputs(12166) <= not(layer0_outputs(11725));
    layer1_outputs(12167) <= layer0_outputs(8778);
    layer1_outputs(12168) <= layer0_outputs(3998);
    layer1_outputs(12169) <= not(layer0_outputs(8115));
    layer1_outputs(12170) <= (layer0_outputs(2792)) xor (layer0_outputs(8306));
    layer1_outputs(12171) <= '0';
    layer1_outputs(12172) <= (layer0_outputs(3820)) xor (layer0_outputs(7602));
    layer1_outputs(12173) <= (layer0_outputs(7224)) and not (layer0_outputs(11282));
    layer1_outputs(12174) <= not((layer0_outputs(10019)) and (layer0_outputs(1569)));
    layer1_outputs(12175) <= not((layer0_outputs(8631)) or (layer0_outputs(3533)));
    layer1_outputs(12176) <= (layer0_outputs(12669)) xor (layer0_outputs(2737));
    layer1_outputs(12177) <= not(layer0_outputs(5556)) or (layer0_outputs(2644));
    layer1_outputs(12178) <= not(layer0_outputs(7031));
    layer1_outputs(12179) <= not(layer0_outputs(5561));
    layer1_outputs(12180) <= layer0_outputs(2884);
    layer1_outputs(12181) <= not((layer0_outputs(11751)) and (layer0_outputs(12398)));
    layer1_outputs(12182) <= layer0_outputs(303);
    layer1_outputs(12183) <= not((layer0_outputs(2961)) and (layer0_outputs(1398)));
    layer1_outputs(12184) <= layer0_outputs(11196);
    layer1_outputs(12185) <= (layer0_outputs(608)) and (layer0_outputs(4291));
    layer1_outputs(12186) <= not(layer0_outputs(7684));
    layer1_outputs(12187) <= not(layer0_outputs(819)) or (layer0_outputs(8644));
    layer1_outputs(12188) <= layer0_outputs(5309);
    layer1_outputs(12189) <= layer0_outputs(2392);
    layer1_outputs(12190) <= (layer0_outputs(8435)) and (layer0_outputs(3338));
    layer1_outputs(12191) <= not(layer0_outputs(4452)) or (layer0_outputs(728));
    layer1_outputs(12192) <= layer0_outputs(11707);
    layer1_outputs(12193) <= not((layer0_outputs(1875)) xor (layer0_outputs(8963)));
    layer1_outputs(12194) <= (layer0_outputs(7352)) and (layer0_outputs(4259));
    layer1_outputs(12195) <= not(layer0_outputs(9419));
    layer1_outputs(12196) <= layer0_outputs(2637);
    layer1_outputs(12197) <= not((layer0_outputs(5860)) xor (layer0_outputs(8558)));
    layer1_outputs(12198) <= (layer0_outputs(2471)) and (layer0_outputs(8858));
    layer1_outputs(12199) <= (layer0_outputs(7883)) and not (layer0_outputs(7596));
    layer1_outputs(12200) <= (layer0_outputs(10599)) xor (layer0_outputs(5139));
    layer1_outputs(12201) <= not((layer0_outputs(7176)) and (layer0_outputs(3106)));
    layer1_outputs(12202) <= layer0_outputs(4534);
    layer1_outputs(12203) <= layer0_outputs(10160);
    layer1_outputs(12204) <= (layer0_outputs(9929)) or (layer0_outputs(4643));
    layer1_outputs(12205) <= not(layer0_outputs(4901));
    layer1_outputs(12206) <= not(layer0_outputs(10999));
    layer1_outputs(12207) <= not(layer0_outputs(9527));
    layer1_outputs(12208) <= (layer0_outputs(8319)) and (layer0_outputs(1029));
    layer1_outputs(12209) <= not((layer0_outputs(6893)) or (layer0_outputs(5629)));
    layer1_outputs(12210) <= not(layer0_outputs(82));
    layer1_outputs(12211) <= not((layer0_outputs(10798)) or (layer0_outputs(7153)));
    layer1_outputs(12212) <= not(layer0_outputs(3066));
    layer1_outputs(12213) <= not(layer0_outputs(421)) or (layer0_outputs(8742));
    layer1_outputs(12214) <= not((layer0_outputs(4896)) or (layer0_outputs(5230)));
    layer1_outputs(12215) <= not(layer0_outputs(3697));
    layer1_outputs(12216) <= not((layer0_outputs(4156)) or (layer0_outputs(9471)));
    layer1_outputs(12217) <= (layer0_outputs(11270)) and not (layer0_outputs(11965));
    layer1_outputs(12218) <= layer0_outputs(3569);
    layer1_outputs(12219) <= not(layer0_outputs(5675)) or (layer0_outputs(9019));
    layer1_outputs(12220) <= not(layer0_outputs(1888));
    layer1_outputs(12221) <= (layer0_outputs(12494)) or (layer0_outputs(4291));
    layer1_outputs(12222) <= not(layer0_outputs(3473));
    layer1_outputs(12223) <= not(layer0_outputs(8714)) or (layer0_outputs(1461));
    layer1_outputs(12224) <= not(layer0_outputs(6206));
    layer1_outputs(12225) <= not(layer0_outputs(320)) or (layer0_outputs(8015));
    layer1_outputs(12226) <= not(layer0_outputs(12243));
    layer1_outputs(12227) <= not(layer0_outputs(2821)) or (layer0_outputs(8316));
    layer1_outputs(12228) <= not(layer0_outputs(12145)) or (layer0_outputs(9654));
    layer1_outputs(12229) <= (layer0_outputs(571)) or (layer0_outputs(5286));
    layer1_outputs(12230) <= not(layer0_outputs(2756));
    layer1_outputs(12231) <= not(layer0_outputs(8040)) or (layer0_outputs(2385));
    layer1_outputs(12232) <= (layer0_outputs(4908)) or (layer0_outputs(1843));
    layer1_outputs(12233) <= not(layer0_outputs(12093)) or (layer0_outputs(4629));
    layer1_outputs(12234) <= layer0_outputs(8300);
    layer1_outputs(12235) <= not((layer0_outputs(4060)) or (layer0_outputs(6003)));
    layer1_outputs(12236) <= (layer0_outputs(11424)) xor (layer0_outputs(7495));
    layer1_outputs(12237) <= (layer0_outputs(8605)) xor (layer0_outputs(7889));
    layer1_outputs(12238) <= layer0_outputs(2936);
    layer1_outputs(12239) <= not((layer0_outputs(4461)) and (layer0_outputs(2133)));
    layer1_outputs(12240) <= (layer0_outputs(3446)) and (layer0_outputs(476));
    layer1_outputs(12241) <= not(layer0_outputs(12453));
    layer1_outputs(12242) <= (layer0_outputs(4868)) and (layer0_outputs(8754));
    layer1_outputs(12243) <= not(layer0_outputs(11666)) or (layer0_outputs(4487));
    layer1_outputs(12244) <= not(layer0_outputs(9240)) or (layer0_outputs(12199));
    layer1_outputs(12245) <= (layer0_outputs(5994)) or (layer0_outputs(6642));
    layer1_outputs(12246) <= (layer0_outputs(6657)) and (layer0_outputs(4402));
    layer1_outputs(12247) <= not((layer0_outputs(11878)) xor (layer0_outputs(7562)));
    layer1_outputs(12248) <= not(layer0_outputs(11172));
    layer1_outputs(12249) <= (layer0_outputs(386)) and (layer0_outputs(10141));
    layer1_outputs(12250) <= (layer0_outputs(9743)) and (layer0_outputs(2258));
    layer1_outputs(12251) <= layer0_outputs(9744);
    layer1_outputs(12252) <= not(layer0_outputs(6348));
    layer1_outputs(12253) <= not(layer0_outputs(5625));
    layer1_outputs(12254) <= (layer0_outputs(10837)) xor (layer0_outputs(4429));
    layer1_outputs(12255) <= not(layer0_outputs(3792));
    layer1_outputs(12256) <= '0';
    layer1_outputs(12257) <= (layer0_outputs(9167)) and (layer0_outputs(7093));
    layer1_outputs(12258) <= (layer0_outputs(9810)) and (layer0_outputs(10214));
    layer1_outputs(12259) <= not(layer0_outputs(6230));
    layer1_outputs(12260) <= not((layer0_outputs(377)) xor (layer0_outputs(9899)));
    layer1_outputs(12261) <= not(layer0_outputs(7386));
    layer1_outputs(12262) <= not(layer0_outputs(1466));
    layer1_outputs(12263) <= layer0_outputs(2088);
    layer1_outputs(12264) <= (layer0_outputs(3870)) and not (layer0_outputs(7573));
    layer1_outputs(12265) <= not(layer0_outputs(8817));
    layer1_outputs(12266) <= (layer0_outputs(4180)) xor (layer0_outputs(2667));
    layer1_outputs(12267) <= not(layer0_outputs(1134)) or (layer0_outputs(8150));
    layer1_outputs(12268) <= (layer0_outputs(11066)) or (layer0_outputs(3278));
    layer1_outputs(12269) <= (layer0_outputs(11023)) or (layer0_outputs(7047));
    layer1_outputs(12270) <= not(layer0_outputs(8744));
    layer1_outputs(12271) <= not(layer0_outputs(1636)) or (layer0_outputs(4581));
    layer1_outputs(12272) <= layer0_outputs(8114);
    layer1_outputs(12273) <= (layer0_outputs(8813)) or (layer0_outputs(7599));
    layer1_outputs(12274) <= not((layer0_outputs(1360)) xor (layer0_outputs(3390)));
    layer1_outputs(12275) <= (layer0_outputs(1860)) xor (layer0_outputs(6280));
    layer1_outputs(12276) <= (layer0_outputs(10000)) or (layer0_outputs(9068));
    layer1_outputs(12277) <= layer0_outputs(3716);
    layer1_outputs(12278) <= not(layer0_outputs(1946));
    layer1_outputs(12279) <= (layer0_outputs(11282)) and not (layer0_outputs(6635));
    layer1_outputs(12280) <= not((layer0_outputs(12546)) xor (layer0_outputs(305)));
    layer1_outputs(12281) <= layer0_outputs(4110);
    layer1_outputs(12282) <= layer0_outputs(149);
    layer1_outputs(12283) <= layer0_outputs(12553);
    layer1_outputs(12284) <= not(layer0_outputs(8728));
    layer1_outputs(12285) <= layer0_outputs(2201);
    layer1_outputs(12286) <= (layer0_outputs(10652)) or (layer0_outputs(11567));
    layer1_outputs(12287) <= not(layer0_outputs(3896));
    layer1_outputs(12288) <= (layer0_outputs(10078)) or (layer0_outputs(3267));
    layer1_outputs(12289) <= not(layer0_outputs(4773));
    layer1_outputs(12290) <= layer0_outputs(7152);
    layer1_outputs(12291) <= layer0_outputs(629);
    layer1_outputs(12292) <= not(layer0_outputs(501));
    layer1_outputs(12293) <= not(layer0_outputs(12600)) or (layer0_outputs(674));
    layer1_outputs(12294) <= layer0_outputs(2914);
    layer1_outputs(12295) <= (layer0_outputs(7479)) or (layer0_outputs(5093));
    layer1_outputs(12296) <= not((layer0_outputs(122)) and (layer0_outputs(4564)));
    layer1_outputs(12297) <= not(layer0_outputs(4263));
    layer1_outputs(12298) <= '0';
    layer1_outputs(12299) <= '1';
    layer1_outputs(12300) <= not((layer0_outputs(9725)) and (layer0_outputs(436)));
    layer1_outputs(12301) <= layer0_outputs(8537);
    layer1_outputs(12302) <= not(layer0_outputs(9605)) or (layer0_outputs(10710));
    layer1_outputs(12303) <= not(layer0_outputs(8134));
    layer1_outputs(12304) <= not((layer0_outputs(2335)) xor (layer0_outputs(11900)));
    layer1_outputs(12305) <= not(layer0_outputs(7172));
    layer1_outputs(12306) <= layer0_outputs(7348);
    layer1_outputs(12307) <= not(layer0_outputs(4936));
    layer1_outputs(12308) <= layer0_outputs(4872);
    layer1_outputs(12309) <= not(layer0_outputs(3116));
    layer1_outputs(12310) <= layer0_outputs(5592);
    layer1_outputs(12311) <= not(layer0_outputs(4915));
    layer1_outputs(12312) <= (layer0_outputs(3906)) xor (layer0_outputs(11199));
    layer1_outputs(12313) <= not(layer0_outputs(8852)) or (layer0_outputs(5918));
    layer1_outputs(12314) <= (layer0_outputs(1398)) xor (layer0_outputs(1214));
    layer1_outputs(12315) <= not((layer0_outputs(12143)) and (layer0_outputs(5730)));
    layer1_outputs(12316) <= layer0_outputs(1727);
    layer1_outputs(12317) <= not(layer0_outputs(5454)) or (layer0_outputs(4318));
    layer1_outputs(12318) <= not(layer0_outputs(8961));
    layer1_outputs(12319) <= layer0_outputs(1654);
    layer1_outputs(12320) <= not(layer0_outputs(6066));
    layer1_outputs(12321) <= (layer0_outputs(9638)) and not (layer0_outputs(7272));
    layer1_outputs(12322) <= (layer0_outputs(6856)) or (layer0_outputs(2906));
    layer1_outputs(12323) <= '1';
    layer1_outputs(12324) <= layer0_outputs(3048);
    layer1_outputs(12325) <= layer0_outputs(6565);
    layer1_outputs(12326) <= not(layer0_outputs(4021));
    layer1_outputs(12327) <= (layer0_outputs(7979)) and not (layer0_outputs(3923));
    layer1_outputs(12328) <= not(layer0_outputs(3561)) or (layer0_outputs(11329));
    layer1_outputs(12329) <= not(layer0_outputs(2264)) or (layer0_outputs(6820));
    layer1_outputs(12330) <= (layer0_outputs(3986)) and (layer0_outputs(4890));
    layer1_outputs(12331) <= not(layer0_outputs(8022));
    layer1_outputs(12332) <= (layer0_outputs(12582)) and (layer0_outputs(9465));
    layer1_outputs(12333) <= not((layer0_outputs(6488)) xor (layer0_outputs(7435)));
    layer1_outputs(12334) <= (layer0_outputs(12510)) or (layer0_outputs(10827));
    layer1_outputs(12335) <= (layer0_outputs(273)) or (layer0_outputs(4455));
    layer1_outputs(12336) <= (layer0_outputs(660)) and not (layer0_outputs(10859));
    layer1_outputs(12337) <= not((layer0_outputs(7782)) and (layer0_outputs(6318)));
    layer1_outputs(12338) <= layer0_outputs(248);
    layer1_outputs(12339) <= not(layer0_outputs(3255)) or (layer0_outputs(9886));
    layer1_outputs(12340) <= layer0_outputs(6649);
    layer1_outputs(12341) <= (layer0_outputs(2507)) and not (layer0_outputs(9878));
    layer1_outputs(12342) <= (layer0_outputs(10119)) or (layer0_outputs(9747));
    layer1_outputs(12343) <= not(layer0_outputs(8848));
    layer1_outputs(12344) <= not(layer0_outputs(2097)) or (layer0_outputs(5505));
    layer1_outputs(12345) <= not((layer0_outputs(12799)) and (layer0_outputs(4044)));
    layer1_outputs(12346) <= (layer0_outputs(7658)) and not (layer0_outputs(5326));
    layer1_outputs(12347) <= not(layer0_outputs(1072));
    layer1_outputs(12348) <= (layer0_outputs(7910)) and not (layer0_outputs(6115));
    layer1_outputs(12349) <= not(layer0_outputs(12080));
    layer1_outputs(12350) <= not((layer0_outputs(6076)) or (layer0_outputs(1990)));
    layer1_outputs(12351) <= not(layer0_outputs(1314)) or (layer0_outputs(10888));
    layer1_outputs(12352) <= not((layer0_outputs(9781)) or (layer0_outputs(10524)));
    layer1_outputs(12353) <= (layer0_outputs(901)) or (layer0_outputs(10175));
    layer1_outputs(12354) <= not(layer0_outputs(6954)) or (layer0_outputs(7864));
    layer1_outputs(12355) <= not(layer0_outputs(1304)) or (layer0_outputs(12343));
    layer1_outputs(12356) <= not(layer0_outputs(4672));
    layer1_outputs(12357) <= layer0_outputs(5547);
    layer1_outputs(12358) <= not(layer0_outputs(11358));
    layer1_outputs(12359) <= layer0_outputs(3934);
    layer1_outputs(12360) <= not(layer0_outputs(4466));
    layer1_outputs(12361) <= not((layer0_outputs(12759)) or (layer0_outputs(9066)));
    layer1_outputs(12362) <= (layer0_outputs(10515)) and not (layer0_outputs(863));
    layer1_outputs(12363) <= not(layer0_outputs(5855));
    layer1_outputs(12364) <= not(layer0_outputs(3759)) or (layer0_outputs(9816));
    layer1_outputs(12365) <= not(layer0_outputs(9751));
    layer1_outputs(12366) <= not((layer0_outputs(10125)) xor (layer0_outputs(4981)));
    layer1_outputs(12367) <= not(layer0_outputs(10335)) or (layer0_outputs(12188));
    layer1_outputs(12368) <= not(layer0_outputs(6616)) or (layer0_outputs(1342));
    layer1_outputs(12369) <= layer0_outputs(5521);
    layer1_outputs(12370) <= layer0_outputs(7313);
    layer1_outputs(12371) <= not(layer0_outputs(12053));
    layer1_outputs(12372) <= (layer0_outputs(12336)) or (layer0_outputs(402));
    layer1_outputs(12373) <= not((layer0_outputs(5913)) xor (layer0_outputs(3109)));
    layer1_outputs(12374) <= not(layer0_outputs(2244));
    layer1_outputs(12375) <= not(layer0_outputs(11838));
    layer1_outputs(12376) <= not(layer0_outputs(5042));
    layer1_outputs(12377) <= not(layer0_outputs(8023));
    layer1_outputs(12378) <= not(layer0_outputs(404));
    layer1_outputs(12379) <= not(layer0_outputs(10502));
    layer1_outputs(12380) <= layer0_outputs(9911);
    layer1_outputs(12381) <= not((layer0_outputs(12387)) xor (layer0_outputs(12552)));
    layer1_outputs(12382) <= (layer0_outputs(6480)) xor (layer0_outputs(5368));
    layer1_outputs(12383) <= not(layer0_outputs(730)) or (layer0_outputs(1947));
    layer1_outputs(12384) <= (layer0_outputs(1442)) and (layer0_outputs(2339));
    layer1_outputs(12385) <= not(layer0_outputs(7425));
    layer1_outputs(12386) <= layer0_outputs(5848);
    layer1_outputs(12387) <= not(layer0_outputs(6218)) or (layer0_outputs(922));
    layer1_outputs(12388) <= '0';
    layer1_outputs(12389) <= not((layer0_outputs(6178)) and (layer0_outputs(6324)));
    layer1_outputs(12390) <= not(layer0_outputs(11040)) or (layer0_outputs(2524));
    layer1_outputs(12391) <= not(layer0_outputs(10148));
    layer1_outputs(12392) <= not(layer0_outputs(5040));
    layer1_outputs(12393) <= layer0_outputs(5357);
    layer1_outputs(12394) <= (layer0_outputs(1702)) or (layer0_outputs(9661));
    layer1_outputs(12395) <= layer0_outputs(5515);
    layer1_outputs(12396) <= not(layer0_outputs(6815));
    layer1_outputs(12397) <= not(layer0_outputs(8478));
    layer1_outputs(12398) <= layer0_outputs(6431);
    layer1_outputs(12399) <= not((layer0_outputs(3310)) or (layer0_outputs(1548)));
    layer1_outputs(12400) <= layer0_outputs(10327);
    layer1_outputs(12401) <= (layer0_outputs(10608)) or (layer0_outputs(6599));
    layer1_outputs(12402) <= not(layer0_outputs(5216)) or (layer0_outputs(11799));
    layer1_outputs(12403) <= (layer0_outputs(8083)) and not (layer0_outputs(6484));
    layer1_outputs(12404) <= not(layer0_outputs(8095));
    layer1_outputs(12405) <= (layer0_outputs(11621)) and (layer0_outputs(11448));
    layer1_outputs(12406) <= not((layer0_outputs(2757)) xor (layer0_outputs(928)));
    layer1_outputs(12407) <= (layer0_outputs(8451)) or (layer0_outputs(5820));
    layer1_outputs(12408) <= (layer0_outputs(7461)) and not (layer0_outputs(12288));
    layer1_outputs(12409) <= (layer0_outputs(5897)) xor (layer0_outputs(12462));
    layer1_outputs(12410) <= not(layer0_outputs(5917));
    layer1_outputs(12411) <= (layer0_outputs(8952)) xor (layer0_outputs(8113));
    layer1_outputs(12412) <= not(layer0_outputs(3492));
    layer1_outputs(12413) <= not(layer0_outputs(6526));
    layer1_outputs(12414) <= (layer0_outputs(2680)) or (layer0_outputs(7448));
    layer1_outputs(12415) <= not(layer0_outputs(12170));
    layer1_outputs(12416) <= not(layer0_outputs(10251));
    layer1_outputs(12417) <= not((layer0_outputs(5116)) and (layer0_outputs(12139)));
    layer1_outputs(12418) <= '1';
    layer1_outputs(12419) <= not(layer0_outputs(11869));
    layer1_outputs(12420) <= not(layer0_outputs(8098));
    layer1_outputs(12421) <= '0';
    layer1_outputs(12422) <= (layer0_outputs(8589)) and not (layer0_outputs(3985));
    layer1_outputs(12423) <= (layer0_outputs(3416)) and (layer0_outputs(3217));
    layer1_outputs(12424) <= layer0_outputs(8349);
    layer1_outputs(12425) <= not(layer0_outputs(4764));
    layer1_outputs(12426) <= not(layer0_outputs(10956)) or (layer0_outputs(4190));
    layer1_outputs(12427) <= (layer0_outputs(3302)) and not (layer0_outputs(10521));
    layer1_outputs(12428) <= layer0_outputs(12645);
    layer1_outputs(12429) <= (layer0_outputs(8534)) and not (layer0_outputs(3160));
    layer1_outputs(12430) <= (layer0_outputs(6037)) and not (layer0_outputs(10966));
    layer1_outputs(12431) <= not((layer0_outputs(1837)) and (layer0_outputs(602)));
    layer1_outputs(12432) <= not(layer0_outputs(965));
    layer1_outputs(12433) <= (layer0_outputs(8139)) xor (layer0_outputs(2451));
    layer1_outputs(12434) <= (layer0_outputs(3587)) and not (layer0_outputs(2047));
    layer1_outputs(12435) <= layer0_outputs(662);
    layer1_outputs(12436) <= not(layer0_outputs(712));
    layer1_outputs(12437) <= not(layer0_outputs(2732)) or (layer0_outputs(11818));
    layer1_outputs(12438) <= (layer0_outputs(2954)) and (layer0_outputs(5314));
    layer1_outputs(12439) <= layer0_outputs(11152);
    layer1_outputs(12440) <= layer0_outputs(12113);
    layer1_outputs(12441) <= not(layer0_outputs(8858)) or (layer0_outputs(2849));
    layer1_outputs(12442) <= not((layer0_outputs(4072)) xor (layer0_outputs(2750)));
    layer1_outputs(12443) <= (layer0_outputs(5041)) and (layer0_outputs(2037));
    layer1_outputs(12444) <= (layer0_outputs(9208)) xor (layer0_outputs(1769));
    layer1_outputs(12445) <= layer0_outputs(3195);
    layer1_outputs(12446) <= (layer0_outputs(3709)) xor (layer0_outputs(5650));
    layer1_outputs(12447) <= not(layer0_outputs(7293)) or (layer0_outputs(11383));
    layer1_outputs(12448) <= (layer0_outputs(10067)) and (layer0_outputs(12219));
    layer1_outputs(12449) <= not((layer0_outputs(4175)) and (layer0_outputs(7554)));
    layer1_outputs(12450) <= not(layer0_outputs(9327));
    layer1_outputs(12451) <= layer0_outputs(598);
    layer1_outputs(12452) <= layer0_outputs(2865);
    layer1_outputs(12453) <= (layer0_outputs(12081)) and not (layer0_outputs(9201));
    layer1_outputs(12454) <= (layer0_outputs(302)) or (layer0_outputs(106));
    layer1_outputs(12455) <= (layer0_outputs(12104)) and (layer0_outputs(6374));
    layer1_outputs(12456) <= not(layer0_outputs(1872));
    layer1_outputs(12457) <= layer0_outputs(11108);
    layer1_outputs(12458) <= layer0_outputs(4097);
    layer1_outputs(12459) <= layer0_outputs(10893);
    layer1_outputs(12460) <= layer0_outputs(2196);
    layer1_outputs(12461) <= (layer0_outputs(8208)) and not (layer0_outputs(2974));
    layer1_outputs(12462) <= layer0_outputs(1437);
    layer1_outputs(12463) <= layer0_outputs(5889);
    layer1_outputs(12464) <= (layer0_outputs(7747)) and not (layer0_outputs(2353));
    layer1_outputs(12465) <= not((layer0_outputs(12167)) or (layer0_outputs(9343)));
    layer1_outputs(12466) <= not(layer0_outputs(5213));
    layer1_outputs(12467) <= not(layer0_outputs(415));
    layer1_outputs(12468) <= (layer0_outputs(629)) and (layer0_outputs(4929));
    layer1_outputs(12469) <= not(layer0_outputs(9139)) or (layer0_outputs(6797));
    layer1_outputs(12470) <= layer0_outputs(5824);
    layer1_outputs(12471) <= not((layer0_outputs(12351)) xor (layer0_outputs(12755)));
    layer1_outputs(12472) <= (layer0_outputs(3487)) and not (layer0_outputs(2170));
    layer1_outputs(12473) <= layer0_outputs(3030);
    layer1_outputs(12474) <= (layer0_outputs(9365)) and not (layer0_outputs(6855));
    layer1_outputs(12475) <= layer0_outputs(3132);
    layer1_outputs(12476) <= layer0_outputs(6112);
    layer1_outputs(12477) <= not(layer0_outputs(1108));
    layer1_outputs(12478) <= not((layer0_outputs(4887)) or (layer0_outputs(1093)));
    layer1_outputs(12479) <= layer0_outputs(440);
    layer1_outputs(12480) <= not(layer0_outputs(8442)) or (layer0_outputs(2584));
    layer1_outputs(12481) <= layer0_outputs(7542);
    layer1_outputs(12482) <= not(layer0_outputs(12042));
    layer1_outputs(12483) <= (layer0_outputs(210)) and not (layer0_outputs(11900));
    layer1_outputs(12484) <= (layer0_outputs(11696)) or (layer0_outputs(9461));
    layer1_outputs(12485) <= not(layer0_outputs(11475));
    layer1_outputs(12486) <= (layer0_outputs(6487)) xor (layer0_outputs(8324));
    layer1_outputs(12487) <= (layer0_outputs(5189)) and not (layer0_outputs(8143));
    layer1_outputs(12488) <= (layer0_outputs(1891)) and not (layer0_outputs(4203));
    layer1_outputs(12489) <= (layer0_outputs(4748)) xor (layer0_outputs(10914));
    layer1_outputs(12490) <= layer0_outputs(4331);
    layer1_outputs(12491) <= not((layer0_outputs(7000)) and (layer0_outputs(12188)));
    layer1_outputs(12492) <= layer0_outputs(6559);
    layer1_outputs(12493) <= (layer0_outputs(7983)) or (layer0_outputs(11391));
    layer1_outputs(12494) <= not(layer0_outputs(8724));
    layer1_outputs(12495) <= not(layer0_outputs(11005));
    layer1_outputs(12496) <= '1';
    layer1_outputs(12497) <= not(layer0_outputs(4040));
    layer1_outputs(12498) <= layer0_outputs(3309);
    layer1_outputs(12499) <= (layer0_outputs(4473)) and not (layer0_outputs(3374));
    layer1_outputs(12500) <= (layer0_outputs(10269)) and not (layer0_outputs(8782));
    layer1_outputs(12501) <= layer0_outputs(8107);
    layer1_outputs(12502) <= not((layer0_outputs(3604)) and (layer0_outputs(11554)));
    layer1_outputs(12503) <= not(layer0_outputs(4212));
    layer1_outputs(12504) <= (layer0_outputs(12574)) xor (layer0_outputs(8550));
    layer1_outputs(12505) <= not((layer0_outputs(11065)) and (layer0_outputs(2444)));
    layer1_outputs(12506) <= (layer0_outputs(9714)) and not (layer0_outputs(4792));
    layer1_outputs(12507) <= not(layer0_outputs(11791));
    layer1_outputs(12508) <= (layer0_outputs(9399)) and not (layer0_outputs(2231));
    layer1_outputs(12509) <= not(layer0_outputs(10062));
    layer1_outputs(12510) <= not((layer0_outputs(6775)) or (layer0_outputs(2367)));
    layer1_outputs(12511) <= (layer0_outputs(2509)) xor (layer0_outputs(3877));
    layer1_outputs(12512) <= not((layer0_outputs(12263)) and (layer0_outputs(9338)));
    layer1_outputs(12513) <= not(layer0_outputs(2074)) or (layer0_outputs(11941));
    layer1_outputs(12514) <= (layer0_outputs(6574)) and (layer0_outputs(9773));
    layer1_outputs(12515) <= (layer0_outputs(8701)) or (layer0_outputs(10096));
    layer1_outputs(12516) <= (layer0_outputs(7186)) xor (layer0_outputs(11701));
    layer1_outputs(12517) <= not((layer0_outputs(2898)) xor (layer0_outputs(8901)));
    layer1_outputs(12518) <= not(layer0_outputs(3612));
    layer1_outputs(12519) <= not(layer0_outputs(6605));
    layer1_outputs(12520) <= not((layer0_outputs(2825)) or (layer0_outputs(9729)));
    layer1_outputs(12521) <= (layer0_outputs(816)) and (layer0_outputs(3719));
    layer1_outputs(12522) <= not(layer0_outputs(5105));
    layer1_outputs(12523) <= not(layer0_outputs(9813));
    layer1_outputs(12524) <= layer0_outputs(12460);
    layer1_outputs(12525) <= not((layer0_outputs(10585)) xor (layer0_outputs(2063)));
    layer1_outputs(12526) <= not(layer0_outputs(5226));
    layer1_outputs(12527) <= not(layer0_outputs(10540));
    layer1_outputs(12528) <= not(layer0_outputs(9061)) or (layer0_outputs(8237));
    layer1_outputs(12529) <= not((layer0_outputs(7527)) and (layer0_outputs(1904)));
    layer1_outputs(12530) <= not(layer0_outputs(12638));
    layer1_outputs(12531) <= not((layer0_outputs(7915)) xor (layer0_outputs(7248)));
    layer1_outputs(12532) <= not((layer0_outputs(10627)) and (layer0_outputs(6060)));
    layer1_outputs(12533) <= layer0_outputs(8323);
    layer1_outputs(12534) <= layer0_outputs(3359);
    layer1_outputs(12535) <= not(layer0_outputs(3045)) or (layer0_outputs(3185));
    layer1_outputs(12536) <= layer0_outputs(10212);
    layer1_outputs(12537) <= not(layer0_outputs(5444)) or (layer0_outputs(11437));
    layer1_outputs(12538) <= (layer0_outputs(11557)) xor (layer0_outputs(6476));
    layer1_outputs(12539) <= not((layer0_outputs(2719)) and (layer0_outputs(10970)));
    layer1_outputs(12540) <= (layer0_outputs(9609)) and not (layer0_outputs(12156));
    layer1_outputs(12541) <= not(layer0_outputs(12030)) or (layer0_outputs(12305));
    layer1_outputs(12542) <= (layer0_outputs(12348)) xor (layer0_outputs(1328));
    layer1_outputs(12543) <= layer0_outputs(9397);
    layer1_outputs(12544) <= not((layer0_outputs(4687)) and (layer0_outputs(8522)));
    layer1_outputs(12545) <= not(layer0_outputs(2181)) or (layer0_outputs(6107));
    layer1_outputs(12546) <= not(layer0_outputs(12443));
    layer1_outputs(12547) <= layer0_outputs(9555);
    layer1_outputs(12548) <= not((layer0_outputs(7548)) and (layer0_outputs(3970)));
    layer1_outputs(12549) <= layer0_outputs(895);
    layer1_outputs(12550) <= not((layer0_outputs(3458)) xor (layer0_outputs(9278)));
    layer1_outputs(12551) <= layer0_outputs(7341);
    layer1_outputs(12552) <= not((layer0_outputs(7267)) or (layer0_outputs(808)));
    layer1_outputs(12553) <= not(layer0_outputs(8790)) or (layer0_outputs(809));
    layer1_outputs(12554) <= (layer0_outputs(3771)) xor (layer0_outputs(12278));
    layer1_outputs(12555) <= (layer0_outputs(3734)) and (layer0_outputs(3671));
    layer1_outputs(12556) <= layer0_outputs(6751);
    layer1_outputs(12557) <= (layer0_outputs(11788)) xor (layer0_outputs(12493));
    layer1_outputs(12558) <= (layer0_outputs(12233)) and not (layer0_outputs(5857));
    layer1_outputs(12559) <= not(layer0_outputs(4558)) or (layer0_outputs(44));
    layer1_outputs(12560) <= '0';
    layer1_outputs(12561) <= layer0_outputs(12262);
    layer1_outputs(12562) <= not(layer0_outputs(11981));
    layer1_outputs(12563) <= '0';
    layer1_outputs(12564) <= not(layer0_outputs(11427)) or (layer0_outputs(10952));
    layer1_outputs(12565) <= not(layer0_outputs(3499)) or (layer0_outputs(7310));
    layer1_outputs(12566) <= (layer0_outputs(34)) and not (layer0_outputs(8317));
    layer1_outputs(12567) <= not((layer0_outputs(8027)) xor (layer0_outputs(8857)));
    layer1_outputs(12568) <= layer0_outputs(111);
    layer1_outputs(12569) <= (layer0_outputs(100)) and not (layer0_outputs(6390));
    layer1_outputs(12570) <= not(layer0_outputs(12283));
    layer1_outputs(12571) <= (layer0_outputs(12316)) or (layer0_outputs(2385));
    layer1_outputs(12572) <= not((layer0_outputs(3489)) and (layer0_outputs(8674)));
    layer1_outputs(12573) <= (layer0_outputs(6980)) and not (layer0_outputs(4684));
    layer1_outputs(12574) <= not(layer0_outputs(11643));
    layer1_outputs(12575) <= layer0_outputs(8564);
    layer1_outputs(12576) <= not(layer0_outputs(10982));
    layer1_outputs(12577) <= not(layer0_outputs(4019));
    layer1_outputs(12578) <= not((layer0_outputs(8988)) and (layer0_outputs(5908)));
    layer1_outputs(12579) <= (layer0_outputs(8452)) xor (layer0_outputs(2747));
    layer1_outputs(12580) <= (layer0_outputs(1460)) and (layer0_outputs(1495));
    layer1_outputs(12581) <= not(layer0_outputs(8688));
    layer1_outputs(12582) <= (layer0_outputs(4386)) and not (layer0_outputs(6741));
    layer1_outputs(12583) <= not((layer0_outputs(7322)) or (layer0_outputs(8910)));
    layer1_outputs(12584) <= layer0_outputs(12721);
    layer1_outputs(12585) <= (layer0_outputs(5410)) or (layer0_outputs(357));
    layer1_outputs(12586) <= not(layer0_outputs(12190));
    layer1_outputs(12587) <= not(layer0_outputs(5076)) or (layer0_outputs(6542));
    layer1_outputs(12588) <= (layer0_outputs(3950)) and not (layer0_outputs(3800));
    layer1_outputs(12589) <= not((layer0_outputs(7905)) xor (layer0_outputs(3722)));
    layer1_outputs(12590) <= (layer0_outputs(9293)) and not (layer0_outputs(9695));
    layer1_outputs(12591) <= (layer0_outputs(1657)) xor (layer0_outputs(2622));
    layer1_outputs(12592) <= (layer0_outputs(9767)) and (layer0_outputs(9493));
    layer1_outputs(12593) <= not((layer0_outputs(5560)) and (layer0_outputs(10566)));
    layer1_outputs(12594) <= not(layer0_outputs(7858));
    layer1_outputs(12595) <= (layer0_outputs(6873)) and not (layer0_outputs(8972));
    layer1_outputs(12596) <= (layer0_outputs(1027)) or (layer0_outputs(6923));
    layer1_outputs(12597) <= not(layer0_outputs(8315)) or (layer0_outputs(6863));
    layer1_outputs(12598) <= not((layer0_outputs(1496)) or (layer0_outputs(5575)));
    layer1_outputs(12599) <= not(layer0_outputs(6300));
    layer1_outputs(12600) <= not(layer0_outputs(4585)) or (layer0_outputs(9273));
    layer1_outputs(12601) <= not((layer0_outputs(6426)) and (layer0_outputs(11009)));
    layer1_outputs(12602) <= (layer0_outputs(11238)) or (layer0_outputs(5992));
    layer1_outputs(12603) <= not(layer0_outputs(3695)) or (layer0_outputs(11651));
    layer1_outputs(12604) <= layer0_outputs(877);
    layer1_outputs(12605) <= not(layer0_outputs(10546));
    layer1_outputs(12606) <= (layer0_outputs(11164)) or (layer0_outputs(177));
    layer1_outputs(12607) <= (layer0_outputs(7081)) xor (layer0_outputs(5704));
    layer1_outputs(12608) <= layer0_outputs(8275);
    layer1_outputs(12609) <= not(layer0_outputs(4785)) or (layer0_outputs(5067));
    layer1_outputs(12610) <= not((layer0_outputs(9200)) and (layer0_outputs(4039)));
    layer1_outputs(12611) <= (layer0_outputs(1988)) xor (layer0_outputs(7769));
    layer1_outputs(12612) <= (layer0_outputs(7285)) and not (layer0_outputs(8813));
    layer1_outputs(12613) <= not((layer0_outputs(1264)) or (layer0_outputs(2610)));
    layer1_outputs(12614) <= not((layer0_outputs(11875)) or (layer0_outputs(11431)));
    layer1_outputs(12615) <= not(layer0_outputs(2521));
    layer1_outputs(12616) <= (layer0_outputs(10441)) xor (layer0_outputs(3512));
    layer1_outputs(12617) <= (layer0_outputs(5909)) and not (layer0_outputs(6337));
    layer1_outputs(12618) <= not((layer0_outputs(780)) and (layer0_outputs(1364)));
    layer1_outputs(12619) <= layer0_outputs(5737);
    layer1_outputs(12620) <= not(layer0_outputs(10245));
    layer1_outputs(12621) <= (layer0_outputs(7430)) and not (layer0_outputs(579));
    layer1_outputs(12622) <= (layer0_outputs(7707)) and not (layer0_outputs(11186));
    layer1_outputs(12623) <= not((layer0_outputs(8788)) and (layer0_outputs(1718)));
    layer1_outputs(12624) <= layer0_outputs(7027);
    layer1_outputs(12625) <= (layer0_outputs(8145)) and not (layer0_outputs(11664));
    layer1_outputs(12626) <= not(layer0_outputs(3568));
    layer1_outputs(12627) <= not(layer0_outputs(12325)) or (layer0_outputs(4047));
    layer1_outputs(12628) <= not(layer0_outputs(8206));
    layer1_outputs(12629) <= layer0_outputs(3355);
    layer1_outputs(12630) <= (layer0_outputs(9923)) and not (layer0_outputs(10259));
    layer1_outputs(12631) <= not(layer0_outputs(8940)) or (layer0_outputs(7666));
    layer1_outputs(12632) <= not(layer0_outputs(8995)) or (layer0_outputs(9362));
    layer1_outputs(12633) <= not(layer0_outputs(9670));
    layer1_outputs(12634) <= (layer0_outputs(1341)) or (layer0_outputs(8560));
    layer1_outputs(12635) <= layer0_outputs(9520);
    layer1_outputs(12636) <= layer0_outputs(1638);
    layer1_outputs(12637) <= (layer0_outputs(5839)) and not (layer0_outputs(3487));
    layer1_outputs(12638) <= not(layer0_outputs(1053));
    layer1_outputs(12639) <= not(layer0_outputs(8189));
    layer1_outputs(12640) <= not(layer0_outputs(6504));
    layer1_outputs(12641) <= not(layer0_outputs(9983)) or (layer0_outputs(11528));
    layer1_outputs(12642) <= not((layer0_outputs(1823)) and (layer0_outputs(7321)));
    layer1_outputs(12643) <= (layer0_outputs(8369)) xor (layer0_outputs(3931));
    layer1_outputs(12644) <= not(layer0_outputs(12561));
    layer1_outputs(12645) <= not(layer0_outputs(10831)) or (layer0_outputs(4276));
    layer1_outputs(12646) <= not(layer0_outputs(11540)) or (layer0_outputs(8064));
    layer1_outputs(12647) <= not((layer0_outputs(11059)) and (layer0_outputs(4888)));
    layer1_outputs(12648) <= (layer0_outputs(872)) and not (layer0_outputs(5291));
    layer1_outputs(12649) <= layer0_outputs(4431);
    layer1_outputs(12650) <= not((layer0_outputs(7578)) and (layer0_outputs(5616)));
    layer1_outputs(12651) <= layer0_outputs(11096);
    layer1_outputs(12652) <= not(layer0_outputs(2790));
    layer1_outputs(12653) <= not((layer0_outputs(12686)) xor (layer0_outputs(5349)));
    layer1_outputs(12654) <= not(layer0_outputs(5531));
    layer1_outputs(12655) <= not(layer0_outputs(8656)) or (layer0_outputs(10319));
    layer1_outputs(12656) <= not(layer0_outputs(5870));
    layer1_outputs(12657) <= not((layer0_outputs(10028)) xor (layer0_outputs(12455)));
    layer1_outputs(12658) <= layer0_outputs(7739);
    layer1_outputs(12659) <= not(layer0_outputs(170));
    layer1_outputs(12660) <= layer0_outputs(6422);
    layer1_outputs(12661) <= not((layer0_outputs(2458)) and (layer0_outputs(4518)));
    layer1_outputs(12662) <= layer0_outputs(5453);
    layer1_outputs(12663) <= not(layer0_outputs(1066)) or (layer0_outputs(4439));
    layer1_outputs(12664) <= (layer0_outputs(10783)) and not (layer0_outputs(2398));
    layer1_outputs(12665) <= not(layer0_outputs(6981));
    layer1_outputs(12666) <= not((layer0_outputs(7381)) and (layer0_outputs(12550)));
    layer1_outputs(12667) <= (layer0_outputs(12644)) and not (layer0_outputs(10012));
    layer1_outputs(12668) <= not(layer0_outputs(5755));
    layer1_outputs(12669) <= (layer0_outputs(6937)) and (layer0_outputs(11234));
    layer1_outputs(12670) <= not((layer0_outputs(9763)) or (layer0_outputs(10737)));
    layer1_outputs(12671) <= not((layer0_outputs(1707)) and (layer0_outputs(7119)));
    layer1_outputs(12672) <= not(layer0_outputs(10963));
    layer1_outputs(12673) <= not(layer0_outputs(3953)) or (layer0_outputs(3906));
    layer1_outputs(12674) <= (layer0_outputs(10733)) xor (layer0_outputs(5316));
    layer1_outputs(12675) <= not(layer0_outputs(12121));
    layer1_outputs(12676) <= layer0_outputs(4837);
    layer1_outputs(12677) <= layer0_outputs(7959);
    layer1_outputs(12678) <= layer0_outputs(10131);
    layer1_outputs(12679) <= (layer0_outputs(3721)) and not (layer0_outputs(9528));
    layer1_outputs(12680) <= layer0_outputs(2851);
    layer1_outputs(12681) <= layer0_outputs(4071);
    layer1_outputs(12682) <= not(layer0_outputs(12500));
    layer1_outputs(12683) <= layer0_outputs(2028);
    layer1_outputs(12684) <= not(layer0_outputs(10827)) or (layer0_outputs(4151));
    layer1_outputs(12685) <= (layer0_outputs(11499)) and not (layer0_outputs(1126));
    layer1_outputs(12686) <= (layer0_outputs(8786)) xor (layer0_outputs(8836));
    layer1_outputs(12687) <= not((layer0_outputs(7838)) or (layer0_outputs(8636)));
    layer1_outputs(12688) <= layer0_outputs(9896);
    layer1_outputs(12689) <= not(layer0_outputs(4092));
    layer1_outputs(12690) <= layer0_outputs(174);
    layer1_outputs(12691) <= not(layer0_outputs(5879));
    layer1_outputs(12692) <= layer0_outputs(11764);
    layer1_outputs(12693) <= not((layer0_outputs(280)) xor (layer0_outputs(9558)));
    layer1_outputs(12694) <= not((layer0_outputs(9279)) or (layer0_outputs(6682)));
    layer1_outputs(12695) <= not(layer0_outputs(10736)) or (layer0_outputs(2121));
    layer1_outputs(12696) <= (layer0_outputs(1486)) and (layer0_outputs(1772));
    layer1_outputs(12697) <= not((layer0_outputs(7246)) and (layer0_outputs(11850)));
    layer1_outputs(12698) <= (layer0_outputs(2033)) or (layer0_outputs(11795));
    layer1_outputs(12699) <= not((layer0_outputs(5581)) and (layer0_outputs(11738)));
    layer1_outputs(12700) <= layer0_outputs(4808);
    layer1_outputs(12701) <= (layer0_outputs(49)) and (layer0_outputs(11920));
    layer1_outputs(12702) <= '0';
    layer1_outputs(12703) <= layer0_outputs(4851);
    layer1_outputs(12704) <= not(layer0_outputs(479));
    layer1_outputs(12705) <= not((layer0_outputs(5651)) xor (layer0_outputs(10983)));
    layer1_outputs(12706) <= not(layer0_outputs(4611));
    layer1_outputs(12707) <= layer0_outputs(12413);
    layer1_outputs(12708) <= not(layer0_outputs(8673));
    layer1_outputs(12709) <= not(layer0_outputs(6475)) or (layer0_outputs(3182));
    layer1_outputs(12710) <= not((layer0_outputs(1691)) or (layer0_outputs(7821)));
    layer1_outputs(12711) <= not(layer0_outputs(5788)) or (layer0_outputs(6213));
    layer1_outputs(12712) <= (layer0_outputs(2002)) and (layer0_outputs(10855));
    layer1_outputs(12713) <= (layer0_outputs(11591)) and (layer0_outputs(4300));
    layer1_outputs(12714) <= not(layer0_outputs(3653));
    layer1_outputs(12715) <= not((layer0_outputs(11368)) and (layer0_outputs(11022)));
    layer1_outputs(12716) <= layer0_outputs(10236);
    layer1_outputs(12717) <= not(layer0_outputs(542)) or (layer0_outputs(6501));
    layer1_outputs(12718) <= (layer0_outputs(1349)) and not (layer0_outputs(4784));
    layer1_outputs(12719) <= layer0_outputs(2130);
    layer1_outputs(12720) <= not((layer0_outputs(11150)) and (layer0_outputs(2677)));
    layer1_outputs(12721) <= not((layer0_outputs(7173)) and (layer0_outputs(9737)));
    layer1_outputs(12722) <= not(layer0_outputs(7250));
    layer1_outputs(12723) <= (layer0_outputs(7251)) and not (layer0_outputs(9759));
    layer1_outputs(12724) <= not((layer0_outputs(11294)) and (layer0_outputs(4143)));
    layer1_outputs(12725) <= (layer0_outputs(10837)) and not (layer0_outputs(11862));
    layer1_outputs(12726) <= (layer0_outputs(10762)) and not (layer0_outputs(7389));
    layer1_outputs(12727) <= layer0_outputs(12493);
    layer1_outputs(12728) <= not((layer0_outputs(2474)) and (layer0_outputs(1265)));
    layer1_outputs(12729) <= '1';
    layer1_outputs(12730) <= not(layer0_outputs(10457)) or (layer0_outputs(3316));
    layer1_outputs(12731) <= '0';
    layer1_outputs(12732) <= not((layer0_outputs(6361)) or (layer0_outputs(8939)));
    layer1_outputs(12733) <= layer0_outputs(5697);
    layer1_outputs(12734) <= (layer0_outputs(6721)) xor (layer0_outputs(187));
    layer1_outputs(12735) <= layer0_outputs(578);
    layer1_outputs(12736) <= (layer0_outputs(9328)) and not (layer0_outputs(11505));
    layer1_outputs(12737) <= layer0_outputs(8190);
    layer1_outputs(12738) <= (layer0_outputs(5428)) and (layer0_outputs(10593));
    layer1_outputs(12739) <= not((layer0_outputs(4578)) and (layer0_outputs(1254)));
    layer1_outputs(12740) <= layer0_outputs(9025);
    layer1_outputs(12741) <= not((layer0_outputs(205)) and (layer0_outputs(4680)));
    layer1_outputs(12742) <= layer0_outputs(5626);
    layer1_outputs(12743) <= '0';
    layer1_outputs(12744) <= (layer0_outputs(12187)) and (layer0_outputs(4647));
    layer1_outputs(12745) <= (layer0_outputs(2096)) and not (layer0_outputs(3949));
    layer1_outputs(12746) <= layer0_outputs(1135);
    layer1_outputs(12747) <= not((layer0_outputs(10060)) and (layer0_outputs(7845)));
    layer1_outputs(12748) <= not(layer0_outputs(7253));
    layer1_outputs(12749) <= (layer0_outputs(12277)) xor (layer0_outputs(9971));
    layer1_outputs(12750) <= (layer0_outputs(4991)) and not (layer0_outputs(10947));
    layer1_outputs(12751) <= '1';
    layer1_outputs(12752) <= not(layer0_outputs(9426)) or (layer0_outputs(12321));
    layer1_outputs(12753) <= layer0_outputs(2955);
    layer1_outputs(12754) <= (layer0_outputs(6670)) and not (layer0_outputs(6302));
    layer1_outputs(12755) <= not(layer0_outputs(8823));
    layer1_outputs(12756) <= not(layer0_outputs(3263)) or (layer0_outputs(943));
    layer1_outputs(12757) <= (layer0_outputs(4693)) xor (layer0_outputs(257));
    layer1_outputs(12758) <= (layer0_outputs(539)) and not (layer0_outputs(2645));
    layer1_outputs(12759) <= (layer0_outputs(2361)) and (layer0_outputs(10091));
    layer1_outputs(12760) <= not(layer0_outputs(10416));
    layer1_outputs(12761) <= (layer0_outputs(855)) and not (layer0_outputs(7264));
    layer1_outputs(12762) <= (layer0_outputs(9198)) and not (layer0_outputs(2048));
    layer1_outputs(12763) <= (layer0_outputs(2360)) and not (layer0_outputs(11873));
    layer1_outputs(12764) <= not((layer0_outputs(6454)) xor (layer0_outputs(11228)));
    layer1_outputs(12765) <= not((layer0_outputs(8341)) or (layer0_outputs(2060)));
    layer1_outputs(12766) <= not(layer0_outputs(10283));
    layer1_outputs(12767) <= not((layer0_outputs(9662)) xor (layer0_outputs(5733)));
    layer1_outputs(12768) <= layer0_outputs(11515);
    layer1_outputs(12769) <= not(layer0_outputs(7277));
    layer1_outputs(12770) <= (layer0_outputs(47)) and not (layer0_outputs(8810));
    layer1_outputs(12771) <= (layer0_outputs(937)) and not (layer0_outputs(6007));
    layer1_outputs(12772) <= (layer0_outputs(4970)) and not (layer0_outputs(8726));
    layer1_outputs(12773) <= (layer0_outputs(10499)) or (layer0_outputs(12434));
    layer1_outputs(12774) <= not(layer0_outputs(7914)) or (layer0_outputs(11862));
    layer1_outputs(12775) <= not((layer0_outputs(10136)) and (layer0_outputs(258)));
    layer1_outputs(12776) <= not(layer0_outputs(11553)) or (layer0_outputs(9023));
    layer1_outputs(12777) <= layer0_outputs(7984);
    layer1_outputs(12778) <= not(layer0_outputs(5066));
    layer1_outputs(12779) <= layer0_outputs(3252);
    layer1_outputs(12780) <= not(layer0_outputs(11309));
    layer1_outputs(12781) <= (layer0_outputs(5408)) or (layer0_outputs(3271));
    layer1_outputs(12782) <= (layer0_outputs(12111)) and (layer0_outputs(3934));
    layer1_outputs(12783) <= not(layer0_outputs(2120));
    layer1_outputs(12784) <= not(layer0_outputs(2638));
    layer1_outputs(12785) <= not(layer0_outputs(8205));
    layer1_outputs(12786) <= not(layer0_outputs(10234));
    layer1_outputs(12787) <= (layer0_outputs(554)) and not (layer0_outputs(9366));
    layer1_outputs(12788) <= not(layer0_outputs(5016));
    layer1_outputs(12789) <= layer0_outputs(5770);
    layer1_outputs(12790) <= not((layer0_outputs(3768)) or (layer0_outputs(8586)));
    layer1_outputs(12791) <= not((layer0_outputs(11340)) or (layer0_outputs(1034)));
    layer1_outputs(12792) <= not(layer0_outputs(5310));
    layer1_outputs(12793) <= not(layer0_outputs(1490)) or (layer0_outputs(3625));
    layer1_outputs(12794) <= not(layer0_outputs(9211));
    layer1_outputs(12795) <= not(layer0_outputs(257));
    layer1_outputs(12796) <= (layer0_outputs(6331)) and not (layer0_outputs(1827));
    layer1_outputs(12797) <= layer0_outputs(10215);
    layer1_outputs(12798) <= not(layer0_outputs(1767)) or (layer0_outputs(7127));
    layer1_outputs(12799) <= not(layer0_outputs(12524));
    layer2_outputs(0) <= layer1_outputs(5610);
    layer2_outputs(1) <= not((layer1_outputs(6367)) and (layer1_outputs(8112)));
    layer2_outputs(2) <= layer1_outputs(2629);
    layer2_outputs(3) <= layer1_outputs(4634);
    layer2_outputs(4) <= not(layer1_outputs(723));
    layer2_outputs(5) <= not(layer1_outputs(3399));
    layer2_outputs(6) <= (layer1_outputs(8317)) and not (layer1_outputs(7366));
    layer2_outputs(7) <= not(layer1_outputs(3896));
    layer2_outputs(8) <= (layer1_outputs(3767)) and not (layer1_outputs(2774));
    layer2_outputs(9) <= not(layer1_outputs(12121));
    layer2_outputs(10) <= not((layer1_outputs(3344)) or (layer1_outputs(8473)));
    layer2_outputs(11) <= layer1_outputs(451);
    layer2_outputs(12) <= layer1_outputs(1371);
    layer2_outputs(13) <= not((layer1_outputs(8428)) xor (layer1_outputs(9939)));
    layer2_outputs(14) <= not(layer1_outputs(3952));
    layer2_outputs(15) <= layer1_outputs(5963);
    layer2_outputs(16) <= not(layer1_outputs(8704));
    layer2_outputs(17) <= not((layer1_outputs(4949)) xor (layer1_outputs(10257)));
    layer2_outputs(18) <= (layer1_outputs(8497)) and (layer1_outputs(4733));
    layer2_outputs(19) <= not((layer1_outputs(2730)) and (layer1_outputs(1542)));
    layer2_outputs(20) <= (layer1_outputs(4342)) and not (layer1_outputs(6110));
    layer2_outputs(21) <= layer1_outputs(6504);
    layer2_outputs(22) <= not(layer1_outputs(3606));
    layer2_outputs(23) <= not(layer1_outputs(4936));
    layer2_outputs(24) <= not(layer1_outputs(6315)) or (layer1_outputs(7331));
    layer2_outputs(25) <= not(layer1_outputs(9918));
    layer2_outputs(26) <= layer1_outputs(6206);
    layer2_outputs(27) <= not((layer1_outputs(257)) xor (layer1_outputs(12126)));
    layer2_outputs(28) <= layer1_outputs(181);
    layer2_outputs(29) <= layer1_outputs(7604);
    layer2_outputs(30) <= not(layer1_outputs(1409));
    layer2_outputs(31) <= not(layer1_outputs(8576));
    layer2_outputs(32) <= layer1_outputs(6177);
    layer2_outputs(33) <= layer1_outputs(1632);
    layer2_outputs(34) <= layer1_outputs(221);
    layer2_outputs(35) <= not(layer1_outputs(11843));
    layer2_outputs(36) <= (layer1_outputs(5418)) and not (layer1_outputs(10480));
    layer2_outputs(37) <= not(layer1_outputs(10531));
    layer2_outputs(38) <= (layer1_outputs(8550)) xor (layer1_outputs(5982));
    layer2_outputs(39) <= not(layer1_outputs(11333)) or (layer1_outputs(7826));
    layer2_outputs(40) <= layer1_outputs(10407);
    layer2_outputs(41) <= not((layer1_outputs(4961)) xor (layer1_outputs(3056)));
    layer2_outputs(42) <= not(layer1_outputs(10796));
    layer2_outputs(43) <= not(layer1_outputs(2538));
    layer2_outputs(44) <= not((layer1_outputs(5492)) or (layer1_outputs(4718)));
    layer2_outputs(45) <= layer1_outputs(4305);
    layer2_outputs(46) <= not(layer1_outputs(12014));
    layer2_outputs(47) <= (layer1_outputs(9920)) or (layer1_outputs(4331));
    layer2_outputs(48) <= not(layer1_outputs(4857));
    layer2_outputs(49) <= not((layer1_outputs(2856)) and (layer1_outputs(10446)));
    layer2_outputs(50) <= (layer1_outputs(12591)) and (layer1_outputs(8933));
    layer2_outputs(51) <= layer1_outputs(3506);
    layer2_outputs(52) <= layer1_outputs(8440);
    layer2_outputs(53) <= (layer1_outputs(1724)) xor (layer1_outputs(8664));
    layer2_outputs(54) <= not(layer1_outputs(476));
    layer2_outputs(55) <= not(layer1_outputs(11468)) or (layer1_outputs(2203));
    layer2_outputs(56) <= layer1_outputs(8432);
    layer2_outputs(57) <= layer1_outputs(10703);
    layer2_outputs(58) <= not(layer1_outputs(4870)) or (layer1_outputs(4894));
    layer2_outputs(59) <= layer1_outputs(7237);
    layer2_outputs(60) <= (layer1_outputs(9579)) xor (layer1_outputs(12155));
    layer2_outputs(61) <= not(layer1_outputs(8347));
    layer2_outputs(62) <= not(layer1_outputs(4974));
    layer2_outputs(63) <= (layer1_outputs(12306)) and (layer1_outputs(10069));
    layer2_outputs(64) <= (layer1_outputs(5810)) and not (layer1_outputs(5795));
    layer2_outputs(65) <= layer1_outputs(11013);
    layer2_outputs(66) <= layer1_outputs(12480);
    layer2_outputs(67) <= not(layer1_outputs(4008));
    layer2_outputs(68) <= not(layer1_outputs(1482));
    layer2_outputs(69) <= not(layer1_outputs(7308));
    layer2_outputs(70) <= not((layer1_outputs(7502)) xor (layer1_outputs(6941)));
    layer2_outputs(71) <= not((layer1_outputs(9242)) and (layer1_outputs(5398)));
    layer2_outputs(72) <= layer1_outputs(1379);
    layer2_outputs(73) <= layer1_outputs(7412);
    layer2_outputs(74) <= layer1_outputs(1016);
    layer2_outputs(75) <= layer1_outputs(6561);
    layer2_outputs(76) <= (layer1_outputs(2846)) and not (layer1_outputs(9105));
    layer2_outputs(77) <= not(layer1_outputs(5417));
    layer2_outputs(78) <= (layer1_outputs(9820)) and (layer1_outputs(12729));
    layer2_outputs(79) <= (layer1_outputs(3071)) and not (layer1_outputs(11888));
    layer2_outputs(80) <= (layer1_outputs(4735)) or (layer1_outputs(10739));
    layer2_outputs(81) <= not((layer1_outputs(10866)) xor (layer1_outputs(8041)));
    layer2_outputs(82) <= not(layer1_outputs(3111));
    layer2_outputs(83) <= not((layer1_outputs(1860)) or (layer1_outputs(12558)));
    layer2_outputs(84) <= (layer1_outputs(8007)) and not (layer1_outputs(9099));
    layer2_outputs(85) <= not(layer1_outputs(5386));
    layer2_outputs(86) <= '1';
    layer2_outputs(87) <= not((layer1_outputs(10462)) xor (layer1_outputs(2095)));
    layer2_outputs(88) <= not((layer1_outputs(10147)) xor (layer1_outputs(9515)));
    layer2_outputs(89) <= not((layer1_outputs(11632)) xor (layer1_outputs(0)));
    layer2_outputs(90) <= (layer1_outputs(5848)) xor (layer1_outputs(9677));
    layer2_outputs(91) <= not(layer1_outputs(1807));
    layer2_outputs(92) <= (layer1_outputs(2932)) and (layer1_outputs(12716));
    layer2_outputs(93) <= layer1_outputs(4432);
    layer2_outputs(94) <= not(layer1_outputs(5301));
    layer2_outputs(95) <= (layer1_outputs(2849)) or (layer1_outputs(7745));
    layer2_outputs(96) <= layer1_outputs(2034);
    layer2_outputs(97) <= not(layer1_outputs(12291)) or (layer1_outputs(10882));
    layer2_outputs(98) <= (layer1_outputs(3243)) and not (layer1_outputs(12700));
    layer2_outputs(99) <= not(layer1_outputs(7212));
    layer2_outputs(100) <= (layer1_outputs(2669)) or (layer1_outputs(875));
    layer2_outputs(101) <= (layer1_outputs(6695)) or (layer1_outputs(6401));
    layer2_outputs(102) <= (layer1_outputs(6564)) xor (layer1_outputs(11673));
    layer2_outputs(103) <= not((layer1_outputs(12775)) or (layer1_outputs(2918)));
    layer2_outputs(104) <= (layer1_outputs(9414)) and not (layer1_outputs(8274));
    layer2_outputs(105) <= not((layer1_outputs(2423)) or (layer1_outputs(6733)));
    layer2_outputs(106) <= not(layer1_outputs(12652));
    layer2_outputs(107) <= layer1_outputs(10492);
    layer2_outputs(108) <= layer1_outputs(5412);
    layer2_outputs(109) <= (layer1_outputs(6459)) or (layer1_outputs(7526));
    layer2_outputs(110) <= (layer1_outputs(3368)) xor (layer1_outputs(3345));
    layer2_outputs(111) <= not((layer1_outputs(6106)) xor (layer1_outputs(173)));
    layer2_outputs(112) <= layer1_outputs(762);
    layer2_outputs(113) <= not(layer1_outputs(1745)) or (layer1_outputs(9651));
    layer2_outputs(114) <= (layer1_outputs(3802)) and not (layer1_outputs(3800));
    layer2_outputs(115) <= (layer1_outputs(1118)) and not (layer1_outputs(12721));
    layer2_outputs(116) <= layer1_outputs(8645);
    layer2_outputs(117) <= (layer1_outputs(8731)) and not (layer1_outputs(4135));
    layer2_outputs(118) <= (layer1_outputs(11456)) and (layer1_outputs(18));
    layer2_outputs(119) <= not(layer1_outputs(1771));
    layer2_outputs(120) <= not(layer1_outputs(3239));
    layer2_outputs(121) <= layer1_outputs(10856);
    layer2_outputs(122) <= not((layer1_outputs(11235)) and (layer1_outputs(11993)));
    layer2_outputs(123) <= not(layer1_outputs(2942));
    layer2_outputs(124) <= (layer1_outputs(2154)) and not (layer1_outputs(1760));
    layer2_outputs(125) <= not(layer1_outputs(11778)) or (layer1_outputs(2448));
    layer2_outputs(126) <= layer1_outputs(2078);
    layer2_outputs(127) <= not((layer1_outputs(11825)) or (layer1_outputs(4267)));
    layer2_outputs(128) <= not(layer1_outputs(8325)) or (layer1_outputs(1013));
    layer2_outputs(129) <= (layer1_outputs(8489)) and not (layer1_outputs(529));
    layer2_outputs(130) <= (layer1_outputs(6834)) or (layer1_outputs(4653));
    layer2_outputs(131) <= layer1_outputs(8737);
    layer2_outputs(132) <= not(layer1_outputs(10337));
    layer2_outputs(133) <= not(layer1_outputs(4618));
    layer2_outputs(134) <= not(layer1_outputs(10490));
    layer2_outputs(135) <= layer1_outputs(1668);
    layer2_outputs(136) <= not((layer1_outputs(1987)) and (layer1_outputs(10625)));
    layer2_outputs(137) <= layer1_outputs(11850);
    layer2_outputs(138) <= (layer1_outputs(1743)) or (layer1_outputs(4885));
    layer2_outputs(139) <= not(layer1_outputs(10997));
    layer2_outputs(140) <= not(layer1_outputs(788)) or (layer1_outputs(2350));
    layer2_outputs(141) <= (layer1_outputs(12252)) and (layer1_outputs(12616));
    layer2_outputs(142) <= (layer1_outputs(11757)) xor (layer1_outputs(4696));
    layer2_outputs(143) <= layer1_outputs(7533);
    layer2_outputs(144) <= layer1_outputs(5047);
    layer2_outputs(145) <= layer1_outputs(8617);
    layer2_outputs(146) <= not(layer1_outputs(12686));
    layer2_outputs(147) <= not((layer1_outputs(4803)) xor (layer1_outputs(4770)));
    layer2_outputs(148) <= (layer1_outputs(4284)) and not (layer1_outputs(8164));
    layer2_outputs(149) <= not(layer1_outputs(2931));
    layer2_outputs(150) <= layer1_outputs(3066);
    layer2_outputs(151) <= not(layer1_outputs(1183));
    layer2_outputs(152) <= layer1_outputs(12296);
    layer2_outputs(153) <= layer1_outputs(8310);
    layer2_outputs(154) <= layer1_outputs(8028);
    layer2_outputs(155) <= not(layer1_outputs(6698));
    layer2_outputs(156) <= not(layer1_outputs(6400));
    layer2_outputs(157) <= not(layer1_outputs(10976));
    layer2_outputs(158) <= not((layer1_outputs(12519)) xor (layer1_outputs(9527)));
    layer2_outputs(159) <= not(layer1_outputs(6922));
    layer2_outputs(160) <= (layer1_outputs(3957)) xor (layer1_outputs(11907));
    layer2_outputs(161) <= '0';
    layer2_outputs(162) <= layer1_outputs(3387);
    layer2_outputs(163) <= not(layer1_outputs(8214));
    layer2_outputs(164) <= not((layer1_outputs(693)) xor (layer1_outputs(2534)));
    layer2_outputs(165) <= (layer1_outputs(4079)) and not (layer1_outputs(1820));
    layer2_outputs(166) <= (layer1_outputs(3470)) and not (layer1_outputs(10289));
    layer2_outputs(167) <= layer1_outputs(5426);
    layer2_outputs(168) <= layer1_outputs(1400);
    layer2_outputs(169) <= (layer1_outputs(7134)) or (layer1_outputs(5555));
    layer2_outputs(170) <= not(layer1_outputs(3648));
    layer2_outputs(171) <= not(layer1_outputs(10343)) or (layer1_outputs(4676));
    layer2_outputs(172) <= (layer1_outputs(10339)) and (layer1_outputs(3915));
    layer2_outputs(173) <= (layer1_outputs(10829)) or (layer1_outputs(7176));
    layer2_outputs(174) <= not(layer1_outputs(5370));
    layer2_outputs(175) <= not(layer1_outputs(11798));
    layer2_outputs(176) <= not((layer1_outputs(6391)) and (layer1_outputs(12771)));
    layer2_outputs(177) <= not(layer1_outputs(7217));
    layer2_outputs(178) <= not(layer1_outputs(12188)) or (layer1_outputs(495));
    layer2_outputs(179) <= not(layer1_outputs(10342)) or (layer1_outputs(9448));
    layer2_outputs(180) <= layer1_outputs(9410);
    layer2_outputs(181) <= not(layer1_outputs(2542));
    layer2_outputs(182) <= not((layer1_outputs(9700)) and (layer1_outputs(4363)));
    layer2_outputs(183) <= not(layer1_outputs(11232));
    layer2_outputs(184) <= not(layer1_outputs(2522)) or (layer1_outputs(5374));
    layer2_outputs(185) <= layer1_outputs(12508);
    layer2_outputs(186) <= not(layer1_outputs(7148)) or (layer1_outputs(2123));
    layer2_outputs(187) <= not((layer1_outputs(8242)) or (layer1_outputs(1283)));
    layer2_outputs(188) <= not(layer1_outputs(6452)) or (layer1_outputs(8725));
    layer2_outputs(189) <= not(layer1_outputs(10160));
    layer2_outputs(190) <= (layer1_outputs(2021)) and not (layer1_outputs(6175));
    layer2_outputs(191) <= not(layer1_outputs(7164));
    layer2_outputs(192) <= layer1_outputs(1930);
    layer2_outputs(193) <= layer1_outputs(7260);
    layer2_outputs(194) <= not(layer1_outputs(9271));
    layer2_outputs(195) <= (layer1_outputs(71)) xor (layer1_outputs(3466));
    layer2_outputs(196) <= layer1_outputs(4539);
    layer2_outputs(197) <= layer1_outputs(7285);
    layer2_outputs(198) <= (layer1_outputs(605)) and not (layer1_outputs(6226));
    layer2_outputs(199) <= layer1_outputs(3313);
    layer2_outputs(200) <= not(layer1_outputs(10915));
    layer2_outputs(201) <= layer1_outputs(6156);
    layer2_outputs(202) <= layer1_outputs(8585);
    layer2_outputs(203) <= (layer1_outputs(2824)) or (layer1_outputs(4225));
    layer2_outputs(204) <= layer1_outputs(390);
    layer2_outputs(205) <= layer1_outputs(5988);
    layer2_outputs(206) <= layer1_outputs(2694);
    layer2_outputs(207) <= not(layer1_outputs(2725));
    layer2_outputs(208) <= layer1_outputs(8453);
    layer2_outputs(209) <= not(layer1_outputs(5412));
    layer2_outputs(210) <= not((layer1_outputs(1619)) and (layer1_outputs(6741)));
    layer2_outputs(211) <= not(layer1_outputs(10500)) or (layer1_outputs(8635));
    layer2_outputs(212) <= not((layer1_outputs(8299)) xor (layer1_outputs(5922)));
    layer2_outputs(213) <= (layer1_outputs(10053)) and not (layer1_outputs(6859));
    layer2_outputs(214) <= not(layer1_outputs(9252));
    layer2_outputs(215) <= not((layer1_outputs(9394)) xor (layer1_outputs(4593)));
    layer2_outputs(216) <= layer1_outputs(11972);
    layer2_outputs(217) <= (layer1_outputs(4968)) or (layer1_outputs(11270));
    layer2_outputs(218) <= not(layer1_outputs(12445));
    layer2_outputs(219) <= not(layer1_outputs(3914));
    layer2_outputs(220) <= not(layer1_outputs(361));
    layer2_outputs(221) <= (layer1_outputs(2557)) and not (layer1_outputs(7005));
    layer2_outputs(222) <= layer1_outputs(4812);
    layer2_outputs(223) <= not(layer1_outputs(11243));
    layer2_outputs(224) <= (layer1_outputs(5153)) or (layer1_outputs(5293));
    layer2_outputs(225) <= not(layer1_outputs(8494)) or (layer1_outputs(6899));
    layer2_outputs(226) <= '1';
    layer2_outputs(227) <= layer1_outputs(1064);
    layer2_outputs(228) <= layer1_outputs(3827);
    layer2_outputs(229) <= layer1_outputs(97);
    layer2_outputs(230) <= (layer1_outputs(607)) xor (layer1_outputs(1933));
    layer2_outputs(231) <= not(layer1_outputs(9991));
    layer2_outputs(232) <= not((layer1_outputs(7291)) and (layer1_outputs(9567)));
    layer2_outputs(233) <= not((layer1_outputs(3098)) or (layer1_outputs(8548)));
    layer2_outputs(234) <= not(layer1_outputs(7274)) or (layer1_outputs(10986));
    layer2_outputs(235) <= layer1_outputs(6664);
    layer2_outputs(236) <= not(layer1_outputs(2274));
    layer2_outputs(237) <= not(layer1_outputs(6080));
    layer2_outputs(238) <= not(layer1_outputs(4185)) or (layer1_outputs(11221));
    layer2_outputs(239) <= (layer1_outputs(8160)) xor (layer1_outputs(9248));
    layer2_outputs(240) <= not(layer1_outputs(3361));
    layer2_outputs(241) <= not((layer1_outputs(12345)) or (layer1_outputs(9152)));
    layer2_outputs(242) <= not(layer1_outputs(8193));
    layer2_outputs(243) <= not((layer1_outputs(5727)) xor (layer1_outputs(11261)));
    layer2_outputs(244) <= (layer1_outputs(8919)) and not (layer1_outputs(2131));
    layer2_outputs(245) <= layer1_outputs(4564);
    layer2_outputs(246) <= not((layer1_outputs(3705)) and (layer1_outputs(9784)));
    layer2_outputs(247) <= not(layer1_outputs(5724));
    layer2_outputs(248) <= not(layer1_outputs(9906));
    layer2_outputs(249) <= layer1_outputs(10733);
    layer2_outputs(250) <= (layer1_outputs(2986)) and (layer1_outputs(7425));
    layer2_outputs(251) <= (layer1_outputs(5564)) and not (layer1_outputs(8619));
    layer2_outputs(252) <= (layer1_outputs(11757)) and not (layer1_outputs(2863));
    layer2_outputs(253) <= not(layer1_outputs(10073));
    layer2_outputs(254) <= not(layer1_outputs(8541));
    layer2_outputs(255) <= layer1_outputs(2324);
    layer2_outputs(256) <= (layer1_outputs(8988)) and (layer1_outputs(7));
    layer2_outputs(257) <= (layer1_outputs(6891)) and (layer1_outputs(4498));
    layer2_outputs(258) <= (layer1_outputs(8382)) and not (layer1_outputs(4405));
    layer2_outputs(259) <= layer1_outputs(3021);
    layer2_outputs(260) <= (layer1_outputs(1740)) and not (layer1_outputs(3437));
    layer2_outputs(261) <= layer1_outputs(7417);
    layer2_outputs(262) <= layer1_outputs(10785);
    layer2_outputs(263) <= layer1_outputs(11809);
    layer2_outputs(264) <= not(layer1_outputs(12368));
    layer2_outputs(265) <= layer1_outputs(2941);
    layer2_outputs(266) <= (layer1_outputs(9233)) xor (layer1_outputs(80));
    layer2_outputs(267) <= not(layer1_outputs(7991)) or (layer1_outputs(1686));
    layer2_outputs(268) <= layer1_outputs(10357);
    layer2_outputs(269) <= '0';
    layer2_outputs(270) <= (layer1_outputs(2457)) xor (layer1_outputs(1121));
    layer2_outputs(271) <= not((layer1_outputs(642)) and (layer1_outputs(10830)));
    layer2_outputs(272) <= '0';
    layer2_outputs(273) <= layer1_outputs(8803);
    layer2_outputs(274) <= layer1_outputs(2949);
    layer2_outputs(275) <= (layer1_outputs(7125)) xor (layer1_outputs(5268));
    layer2_outputs(276) <= not(layer1_outputs(2705));
    layer2_outputs(277) <= layer1_outputs(5435);
    layer2_outputs(278) <= layer1_outputs(12626);
    layer2_outputs(279) <= layer1_outputs(3183);
    layer2_outputs(280) <= not((layer1_outputs(8615)) xor (layer1_outputs(11856)));
    layer2_outputs(281) <= (layer1_outputs(2292)) or (layer1_outputs(485));
    layer2_outputs(282) <= not((layer1_outputs(1736)) xor (layer1_outputs(4479)));
    layer2_outputs(283) <= not(layer1_outputs(7882)) or (layer1_outputs(12263));
    layer2_outputs(284) <= layer1_outputs(3223);
    layer2_outputs(285) <= not(layer1_outputs(2412));
    layer2_outputs(286) <= (layer1_outputs(4222)) and not (layer1_outputs(9678));
    layer2_outputs(287) <= (layer1_outputs(12128)) or (layer1_outputs(1681));
    layer2_outputs(288) <= not((layer1_outputs(11021)) xor (layer1_outputs(11290)));
    layer2_outputs(289) <= layer1_outputs(3123);
    layer2_outputs(290) <= not((layer1_outputs(7334)) xor (layer1_outputs(4615)));
    layer2_outputs(291) <= layer1_outputs(12591);
    layer2_outputs(292) <= (layer1_outputs(5424)) and (layer1_outputs(4173));
    layer2_outputs(293) <= not(layer1_outputs(6902));
    layer2_outputs(294) <= not((layer1_outputs(8289)) xor (layer1_outputs(7907)));
    layer2_outputs(295) <= layer1_outputs(7460);
    layer2_outputs(296) <= (layer1_outputs(2744)) and not (layer1_outputs(3727));
    layer2_outputs(297) <= not(layer1_outputs(10444));
    layer2_outputs(298) <= not(layer1_outputs(3445));
    layer2_outputs(299) <= not(layer1_outputs(3391));
    layer2_outputs(300) <= not(layer1_outputs(5871));
    layer2_outputs(301) <= layer1_outputs(2783);
    layer2_outputs(302) <= not((layer1_outputs(1030)) xor (layer1_outputs(10278)));
    layer2_outputs(303) <= not(layer1_outputs(3102)) or (layer1_outputs(27));
    layer2_outputs(304) <= not(layer1_outputs(3115));
    layer2_outputs(305) <= not(layer1_outputs(11245));
    layer2_outputs(306) <= not(layer1_outputs(5691)) or (layer1_outputs(4851));
    layer2_outputs(307) <= not(layer1_outputs(2754));
    layer2_outputs(308) <= not((layer1_outputs(9833)) or (layer1_outputs(2)));
    layer2_outputs(309) <= not(layer1_outputs(7424));
    layer2_outputs(310) <= (layer1_outputs(10527)) or (layer1_outputs(11941));
    layer2_outputs(311) <= not(layer1_outputs(3330));
    layer2_outputs(312) <= not(layer1_outputs(7624));
    layer2_outputs(313) <= layer1_outputs(8322);
    layer2_outputs(314) <= not(layer1_outputs(8532));
    layer2_outputs(315) <= layer1_outputs(1390);
    layer2_outputs(316) <= (layer1_outputs(8857)) and (layer1_outputs(5726));
    layer2_outputs(317) <= not((layer1_outputs(3481)) and (layer1_outputs(10119)));
    layer2_outputs(318) <= (layer1_outputs(8831)) xor (layer1_outputs(7219));
    layer2_outputs(319) <= (layer1_outputs(10944)) and not (layer1_outputs(11429));
    layer2_outputs(320) <= layer1_outputs(6969);
    layer2_outputs(321) <= not(layer1_outputs(6735));
    layer2_outputs(322) <= (layer1_outputs(2944)) or (layer1_outputs(4632));
    layer2_outputs(323) <= not(layer1_outputs(3675));
    layer2_outputs(324) <= layer1_outputs(6514);
    layer2_outputs(325) <= not(layer1_outputs(1367));
    layer2_outputs(326) <= layer1_outputs(8727);
    layer2_outputs(327) <= not((layer1_outputs(1092)) and (layer1_outputs(10522)));
    layer2_outputs(328) <= not(layer1_outputs(1026));
    layer2_outputs(329) <= (layer1_outputs(6961)) xor (layer1_outputs(2217));
    layer2_outputs(330) <= (layer1_outputs(10641)) and not (layer1_outputs(2022));
    layer2_outputs(331) <= (layer1_outputs(6455)) and (layer1_outputs(10734));
    layer2_outputs(332) <= (layer1_outputs(9086)) and not (layer1_outputs(1296));
    layer2_outputs(333) <= not(layer1_outputs(8801));
    layer2_outputs(334) <= (layer1_outputs(4645)) and not (layer1_outputs(10674));
    layer2_outputs(335) <= not((layer1_outputs(9769)) xor (layer1_outputs(11820)));
    layer2_outputs(336) <= not(layer1_outputs(5392)) or (layer1_outputs(5999));
    layer2_outputs(337) <= not(layer1_outputs(10623)) or (layer1_outputs(11024));
    layer2_outputs(338) <= not(layer1_outputs(280)) or (layer1_outputs(3785));
    layer2_outputs(339) <= not(layer1_outputs(794)) or (layer1_outputs(7185));
    layer2_outputs(340) <= (layer1_outputs(1588)) xor (layer1_outputs(8597));
    layer2_outputs(341) <= not(layer1_outputs(10678));
    layer2_outputs(342) <= not(layer1_outputs(6772));
    layer2_outputs(343) <= (layer1_outputs(5601)) and not (layer1_outputs(8435));
    layer2_outputs(344) <= not(layer1_outputs(10832));
    layer2_outputs(345) <= not(layer1_outputs(4137));
    layer2_outputs(346) <= layer1_outputs(12690);
    layer2_outputs(347) <= not(layer1_outputs(7663)) or (layer1_outputs(11239));
    layer2_outputs(348) <= not(layer1_outputs(12263));
    layer2_outputs(349) <= (layer1_outputs(11587)) and not (layer1_outputs(3045));
    layer2_outputs(350) <= not(layer1_outputs(3253)) or (layer1_outputs(7875));
    layer2_outputs(351) <= (layer1_outputs(10313)) xor (layer1_outputs(7754));
    layer2_outputs(352) <= not((layer1_outputs(6593)) xor (layer1_outputs(1701)));
    layer2_outputs(353) <= layer1_outputs(9066);
    layer2_outputs(354) <= not(layer1_outputs(8725));
    layer2_outputs(355) <= not(layer1_outputs(5777));
    layer2_outputs(356) <= layer1_outputs(7771);
    layer2_outputs(357) <= (layer1_outputs(11285)) and not (layer1_outputs(7065));
    layer2_outputs(358) <= (layer1_outputs(11223)) xor (layer1_outputs(11833));
    layer2_outputs(359) <= layer1_outputs(6039);
    layer2_outputs(360) <= layer1_outputs(8451);
    layer2_outputs(361) <= (layer1_outputs(6110)) or (layer1_outputs(4327));
    layer2_outputs(362) <= layer1_outputs(2451);
    layer2_outputs(363) <= layer1_outputs(473);
    layer2_outputs(364) <= layer1_outputs(6298);
    layer2_outputs(365) <= layer1_outputs(5433);
    layer2_outputs(366) <= not((layer1_outputs(3882)) xor (layer1_outputs(10539)));
    layer2_outputs(367) <= layer1_outputs(5297);
    layer2_outputs(368) <= layer1_outputs(2170);
    layer2_outputs(369) <= (layer1_outputs(12460)) or (layer1_outputs(7840));
    layer2_outputs(370) <= (layer1_outputs(3603)) and not (layer1_outputs(603));
    layer2_outputs(371) <= layer1_outputs(6359);
    layer2_outputs(372) <= not(layer1_outputs(12099)) or (layer1_outputs(8533));
    layer2_outputs(373) <= layer1_outputs(4677);
    layer2_outputs(374) <= not((layer1_outputs(2732)) or (layer1_outputs(10321)));
    layer2_outputs(375) <= layer1_outputs(4319);
    layer2_outputs(376) <= (layer1_outputs(2995)) or (layer1_outputs(3673));
    layer2_outputs(377) <= not((layer1_outputs(6123)) or (layer1_outputs(5307)));
    layer2_outputs(378) <= (layer1_outputs(4076)) and not (layer1_outputs(1245));
    layer2_outputs(379) <= not((layer1_outputs(9811)) xor (layer1_outputs(8008)));
    layer2_outputs(380) <= layer1_outputs(8314);
    layer2_outputs(381) <= not((layer1_outputs(6877)) or (layer1_outputs(2287)));
    layer2_outputs(382) <= not(layer1_outputs(11226)) or (layer1_outputs(1486));
    layer2_outputs(383) <= layer1_outputs(1463);
    layer2_outputs(384) <= (layer1_outputs(11803)) or (layer1_outputs(1166));
    layer2_outputs(385) <= not(layer1_outputs(12603)) or (layer1_outputs(6527));
    layer2_outputs(386) <= not(layer1_outputs(6861));
    layer2_outputs(387) <= not((layer1_outputs(10181)) xor (layer1_outputs(9169)));
    layer2_outputs(388) <= (layer1_outputs(11256)) xor (layer1_outputs(4860));
    layer2_outputs(389) <= layer1_outputs(4911);
    layer2_outputs(390) <= layer1_outputs(10400);
    layer2_outputs(391) <= not(layer1_outputs(8364));
    layer2_outputs(392) <= not(layer1_outputs(11451));
    layer2_outputs(393) <= not(layer1_outputs(9458)) or (layer1_outputs(6511));
    layer2_outputs(394) <= not(layer1_outputs(5851));
    layer2_outputs(395) <= layer1_outputs(12283);
    layer2_outputs(396) <= (layer1_outputs(5371)) or (layer1_outputs(5036));
    layer2_outputs(397) <= not((layer1_outputs(922)) xor (layer1_outputs(288)));
    layer2_outputs(398) <= not(layer1_outputs(5136)) or (layer1_outputs(1286));
    layer2_outputs(399) <= layer1_outputs(3203);
    layer2_outputs(400) <= layer1_outputs(3543);
    layer2_outputs(401) <= not((layer1_outputs(2481)) and (layer1_outputs(6893)));
    layer2_outputs(402) <= not(layer1_outputs(10529));
    layer2_outputs(403) <= not((layer1_outputs(2495)) and (layer1_outputs(1366)));
    layer2_outputs(404) <= (layer1_outputs(7429)) and not (layer1_outputs(7923));
    layer2_outputs(405) <= '0';
    layer2_outputs(406) <= layer1_outputs(3305);
    layer2_outputs(407) <= (layer1_outputs(4666)) and (layer1_outputs(8413));
    layer2_outputs(408) <= (layer1_outputs(1426)) or (layer1_outputs(11549));
    layer2_outputs(409) <= (layer1_outputs(6512)) and not (layer1_outputs(6546));
    layer2_outputs(410) <= (layer1_outputs(11471)) and (layer1_outputs(5567));
    layer2_outputs(411) <= layer1_outputs(9649);
    layer2_outputs(412) <= (layer1_outputs(9063)) or (layer1_outputs(91));
    layer2_outputs(413) <= (layer1_outputs(2274)) or (layer1_outputs(7493));
    layer2_outputs(414) <= (layer1_outputs(3256)) or (layer1_outputs(5175));
    layer2_outputs(415) <= not(layer1_outputs(745));
    layer2_outputs(416) <= (layer1_outputs(10850)) and not (layer1_outputs(3));
    layer2_outputs(417) <= layer1_outputs(6191);
    layer2_outputs(418) <= not(layer1_outputs(3537));
    layer2_outputs(419) <= not((layer1_outputs(9272)) and (layer1_outputs(9522)));
    layer2_outputs(420) <= not((layer1_outputs(3614)) and (layer1_outputs(4775)));
    layer2_outputs(421) <= not(layer1_outputs(8309));
    layer2_outputs(422) <= (layer1_outputs(9284)) and (layer1_outputs(4165));
    layer2_outputs(423) <= (layer1_outputs(10531)) and (layer1_outputs(6224));
    layer2_outputs(424) <= layer1_outputs(9939);
    layer2_outputs(425) <= layer1_outputs(6160);
    layer2_outputs(426) <= layer1_outputs(7047);
    layer2_outputs(427) <= (layer1_outputs(3506)) xor (layer1_outputs(4212));
    layer2_outputs(428) <= not((layer1_outputs(4491)) or (layer1_outputs(5397)));
    layer2_outputs(429) <= layer1_outputs(1373);
    layer2_outputs(430) <= (layer1_outputs(1658)) xor (layer1_outputs(10123));
    layer2_outputs(431) <= layer1_outputs(7223);
    layer2_outputs(432) <= layer1_outputs(11627);
    layer2_outputs(433) <= not(layer1_outputs(2919)) or (layer1_outputs(6426));
    layer2_outputs(434) <= layer1_outputs(3854);
    layer2_outputs(435) <= layer1_outputs(6757);
    layer2_outputs(436) <= not(layer1_outputs(12047));
    layer2_outputs(437) <= layer1_outputs(8139);
    layer2_outputs(438) <= layer1_outputs(4319);
    layer2_outputs(439) <= layer1_outputs(8569);
    layer2_outputs(440) <= not(layer1_outputs(7757));
    layer2_outputs(441) <= '1';
    layer2_outputs(442) <= (layer1_outputs(5715)) and not (layer1_outputs(11250));
    layer2_outputs(443) <= not(layer1_outputs(3763)) or (layer1_outputs(10569));
    layer2_outputs(444) <= (layer1_outputs(4665)) and not (layer1_outputs(1528));
    layer2_outputs(445) <= (layer1_outputs(7488)) and not (layer1_outputs(376));
    layer2_outputs(446) <= not((layer1_outputs(4793)) or (layer1_outputs(4416)));
    layer2_outputs(447) <= layer1_outputs(11677);
    layer2_outputs(448) <= (layer1_outputs(7815)) and not (layer1_outputs(7774));
    layer2_outputs(449) <= not((layer1_outputs(5473)) and (layer1_outputs(11383)));
    layer2_outputs(450) <= not(layer1_outputs(11512));
    layer2_outputs(451) <= (layer1_outputs(10285)) and (layer1_outputs(4848));
    layer2_outputs(452) <= layer1_outputs(9052);
    layer2_outputs(453) <= not((layer1_outputs(8060)) xor (layer1_outputs(5257)));
    layer2_outputs(454) <= not(layer1_outputs(10978));
    layer2_outputs(455) <= not(layer1_outputs(10463));
    layer2_outputs(456) <= not(layer1_outputs(6167)) or (layer1_outputs(7027));
    layer2_outputs(457) <= not((layer1_outputs(903)) xor (layer1_outputs(5932)));
    layer2_outputs(458) <= not((layer1_outputs(10048)) xor (layer1_outputs(5672)));
    layer2_outputs(459) <= (layer1_outputs(6558)) and not (layer1_outputs(9847));
    layer2_outputs(460) <= not(layer1_outputs(7453));
    layer2_outputs(461) <= not(layer1_outputs(12391));
    layer2_outputs(462) <= layer1_outputs(2745);
    layer2_outputs(463) <= (layer1_outputs(10901)) and not (layer1_outputs(10445));
    layer2_outputs(464) <= layer1_outputs(10638);
    layer2_outputs(465) <= not(layer1_outputs(3576)) or (layer1_outputs(12138));
    layer2_outputs(466) <= not(layer1_outputs(11681));
    layer2_outputs(467) <= not((layer1_outputs(12433)) xor (layer1_outputs(4579)));
    layer2_outputs(468) <= not((layer1_outputs(6257)) or (layer1_outputs(7912)));
    layer2_outputs(469) <= not((layer1_outputs(10187)) and (layer1_outputs(4810)));
    layer2_outputs(470) <= not(layer1_outputs(8763)) or (layer1_outputs(10635));
    layer2_outputs(471) <= not((layer1_outputs(233)) xor (layer1_outputs(382)));
    layer2_outputs(472) <= not(layer1_outputs(3961));
    layer2_outputs(473) <= not(layer1_outputs(10437));
    layer2_outputs(474) <= not(layer1_outputs(2256));
    layer2_outputs(475) <= not(layer1_outputs(473));
    layer2_outputs(476) <= layer1_outputs(1379);
    layer2_outputs(477) <= not(layer1_outputs(9350)) or (layer1_outputs(4489));
    layer2_outputs(478) <= (layer1_outputs(6287)) and not (layer1_outputs(9876));
    layer2_outputs(479) <= '0';
    layer2_outputs(480) <= not(layer1_outputs(11362));
    layer2_outputs(481) <= layer1_outputs(4847);
    layer2_outputs(482) <= (layer1_outputs(7484)) xor (layer1_outputs(8534));
    layer2_outputs(483) <= layer1_outputs(9562);
    layer2_outputs(484) <= not((layer1_outputs(9513)) xor (layer1_outputs(728)));
    layer2_outputs(485) <= layer1_outputs(3352);
    layer2_outputs(486) <= not(layer1_outputs(3757));
    layer2_outputs(487) <= not(layer1_outputs(7976));
    layer2_outputs(488) <= not((layer1_outputs(4120)) or (layer1_outputs(10768)));
    layer2_outputs(489) <= not(layer1_outputs(2476)) or (layer1_outputs(1538));
    layer2_outputs(490) <= not((layer1_outputs(1431)) or (layer1_outputs(7721)));
    layer2_outputs(491) <= (layer1_outputs(7143)) and (layer1_outputs(996));
    layer2_outputs(492) <= not((layer1_outputs(9625)) and (layer1_outputs(5611)));
    layer2_outputs(493) <= not(layer1_outputs(11533));
    layer2_outputs(494) <= not(layer1_outputs(10984)) or (layer1_outputs(3508));
    layer2_outputs(495) <= not(layer1_outputs(3981));
    layer2_outputs(496) <= not(layer1_outputs(8387));
    layer2_outputs(497) <= not(layer1_outputs(4774)) or (layer1_outputs(10792));
    layer2_outputs(498) <= '1';
    layer2_outputs(499) <= not((layer1_outputs(3831)) xor (layer1_outputs(7805)));
    layer2_outputs(500) <= (layer1_outputs(8108)) and not (layer1_outputs(1816));
    layer2_outputs(501) <= layer1_outputs(10962);
    layer2_outputs(502) <= (layer1_outputs(9192)) and not (layer1_outputs(6089));
    layer2_outputs(503) <= layer1_outputs(12303);
    layer2_outputs(504) <= (layer1_outputs(4332)) and (layer1_outputs(8952));
    layer2_outputs(505) <= layer1_outputs(10961);
    layer2_outputs(506) <= (layer1_outputs(2510)) and not (layer1_outputs(1679));
    layer2_outputs(507) <= not((layer1_outputs(3925)) xor (layer1_outputs(100)));
    layer2_outputs(508) <= not((layer1_outputs(730)) or (layer1_outputs(9572)));
    layer2_outputs(509) <= not(layer1_outputs(91));
    layer2_outputs(510) <= (layer1_outputs(11482)) xor (layer1_outputs(9709));
    layer2_outputs(511) <= not((layer1_outputs(987)) and (layer1_outputs(12330)));
    layer2_outputs(512) <= (layer1_outputs(9073)) xor (layer1_outputs(8189));
    layer2_outputs(513) <= (layer1_outputs(12603)) and (layer1_outputs(11930));
    layer2_outputs(514) <= not((layer1_outputs(10627)) xor (layer1_outputs(2707)));
    layer2_outputs(515) <= '0';
    layer2_outputs(516) <= not(layer1_outputs(2677)) or (layer1_outputs(7294));
    layer2_outputs(517) <= layer1_outputs(12762);
    layer2_outputs(518) <= layer1_outputs(6998);
    layer2_outputs(519) <= (layer1_outputs(4182)) and not (layer1_outputs(10089));
    layer2_outputs(520) <= layer1_outputs(11140);
    layer2_outputs(521) <= (layer1_outputs(7261)) xor (layer1_outputs(1573));
    layer2_outputs(522) <= (layer1_outputs(6078)) xor (layer1_outputs(8799));
    layer2_outputs(523) <= not((layer1_outputs(4924)) and (layer1_outputs(11673)));
    layer2_outputs(524) <= not(layer1_outputs(8222));
    layer2_outputs(525) <= not(layer1_outputs(7502));
    layer2_outputs(526) <= not((layer1_outputs(4275)) xor (layer1_outputs(2822)));
    layer2_outputs(527) <= layer1_outputs(9622);
    layer2_outputs(528) <= (layer1_outputs(10717)) or (layer1_outputs(5148));
    layer2_outputs(529) <= not(layer1_outputs(5007)) or (layer1_outputs(5476));
    layer2_outputs(530) <= not(layer1_outputs(4024));
    layer2_outputs(531) <= not(layer1_outputs(12298)) or (layer1_outputs(1560));
    layer2_outputs(532) <= layer1_outputs(9328);
    layer2_outputs(533) <= layer1_outputs(10320);
    layer2_outputs(534) <= (layer1_outputs(12609)) or (layer1_outputs(8665));
    layer2_outputs(535) <= not(layer1_outputs(9834));
    layer2_outputs(536) <= (layer1_outputs(5009)) xor (layer1_outputs(876));
    layer2_outputs(537) <= not((layer1_outputs(10059)) and (layer1_outputs(933)));
    layer2_outputs(538) <= layer1_outputs(2440);
    layer2_outputs(539) <= (layer1_outputs(10348)) or (layer1_outputs(9260));
    layer2_outputs(540) <= layer1_outputs(1667);
    layer2_outputs(541) <= (layer1_outputs(11008)) and not (layer1_outputs(947));
    layer2_outputs(542) <= layer1_outputs(9259);
    layer2_outputs(543) <= (layer1_outputs(8867)) or (layer1_outputs(12310));
    layer2_outputs(544) <= not((layer1_outputs(10775)) or (layer1_outputs(1270)));
    layer2_outputs(545) <= (layer1_outputs(10513)) and (layer1_outputs(11918));
    layer2_outputs(546) <= layer1_outputs(7377);
    layer2_outputs(547) <= (layer1_outputs(3306)) and not (layer1_outputs(8808));
    layer2_outputs(548) <= not(layer1_outputs(1962));
    layer2_outputs(549) <= (layer1_outputs(7642)) xor (layer1_outputs(5539));
    layer2_outputs(550) <= not((layer1_outputs(10518)) xor (layer1_outputs(6156)));
    layer2_outputs(551) <= not(layer1_outputs(7004));
    layer2_outputs(552) <= not(layer1_outputs(2992));
    layer2_outputs(553) <= not(layer1_outputs(10322));
    layer2_outputs(554) <= (layer1_outputs(9843)) and (layer1_outputs(12090));
    layer2_outputs(555) <= not(layer1_outputs(12158));
    layer2_outputs(556) <= not(layer1_outputs(5974));
    layer2_outputs(557) <= (layer1_outputs(7470)) and (layer1_outputs(8411));
    layer2_outputs(558) <= not(layer1_outputs(4139));
    layer2_outputs(559) <= not((layer1_outputs(12375)) xor (layer1_outputs(6747)));
    layer2_outputs(560) <= layer1_outputs(5261);
    layer2_outputs(561) <= not(layer1_outputs(8930));
    layer2_outputs(562) <= not((layer1_outputs(8279)) or (layer1_outputs(2865)));
    layer2_outputs(563) <= layer1_outputs(7594);
    layer2_outputs(564) <= (layer1_outputs(11933)) and (layer1_outputs(9679));
    layer2_outputs(565) <= not(layer1_outputs(11660));
    layer2_outputs(566) <= layer1_outputs(12365);
    layer2_outputs(567) <= not(layer1_outputs(4772));
    layer2_outputs(568) <= layer1_outputs(5409);
    layer2_outputs(569) <= (layer1_outputs(10102)) xor (layer1_outputs(9583));
    layer2_outputs(570) <= (layer1_outputs(5773)) or (layer1_outputs(8506));
    layer2_outputs(571) <= not((layer1_outputs(7521)) xor (layer1_outputs(5511)));
    layer2_outputs(572) <= layer1_outputs(4090);
    layer2_outputs(573) <= not(layer1_outputs(8462));
    layer2_outputs(574) <= not(layer1_outputs(665));
    layer2_outputs(575) <= not((layer1_outputs(3547)) or (layer1_outputs(7288)));
    layer2_outputs(576) <= (layer1_outputs(8040)) or (layer1_outputs(12505));
    layer2_outputs(577) <= not(layer1_outputs(2864));
    layer2_outputs(578) <= not(layer1_outputs(347));
    layer2_outputs(579) <= layer1_outputs(6491);
    layer2_outputs(580) <= not((layer1_outputs(2712)) or (layer1_outputs(2626)));
    layer2_outputs(581) <= (layer1_outputs(12547)) xor (layer1_outputs(2209));
    layer2_outputs(582) <= layer1_outputs(9756);
    layer2_outputs(583) <= (layer1_outputs(5991)) and not (layer1_outputs(6799));
    layer2_outputs(584) <= (layer1_outputs(3451)) or (layer1_outputs(11434));
    layer2_outputs(585) <= layer1_outputs(5684);
    layer2_outputs(586) <= layer1_outputs(7889);
    layer2_outputs(587) <= not(layer1_outputs(1908));
    layer2_outputs(588) <= not(layer1_outputs(10492)) or (layer1_outputs(527));
    layer2_outputs(589) <= not(layer1_outputs(5990));
    layer2_outputs(590) <= not(layer1_outputs(5456));
    layer2_outputs(591) <= (layer1_outputs(472)) xor (layer1_outputs(2784));
    layer2_outputs(592) <= (layer1_outputs(1469)) and (layer1_outputs(3993));
    layer2_outputs(593) <= (layer1_outputs(8957)) and (layer1_outputs(1640));
    layer2_outputs(594) <= not(layer1_outputs(10280));
    layer2_outputs(595) <= not(layer1_outputs(5234));
    layer2_outputs(596) <= layer1_outputs(2998);
    layer2_outputs(597) <= layer1_outputs(3332);
    layer2_outputs(598) <= layer1_outputs(10967);
    layer2_outputs(599) <= layer1_outputs(10267);
    layer2_outputs(600) <= layer1_outputs(1089);
    layer2_outputs(601) <= layer1_outputs(4637);
    layer2_outputs(602) <= (layer1_outputs(12739)) xor (layer1_outputs(2413));
    layer2_outputs(603) <= (layer1_outputs(6130)) and not (layer1_outputs(4180));
    layer2_outputs(604) <= layer1_outputs(6896);
    layer2_outputs(605) <= layer1_outputs(530);
    layer2_outputs(606) <= not(layer1_outputs(3840));
    layer2_outputs(607) <= not(layer1_outputs(4250));
    layer2_outputs(608) <= not(layer1_outputs(6196));
    layer2_outputs(609) <= (layer1_outputs(3606)) or (layer1_outputs(6625));
    layer2_outputs(610) <= (layer1_outputs(9373)) xor (layer1_outputs(4904));
    layer2_outputs(611) <= (layer1_outputs(9699)) and not (layer1_outputs(1947));
    layer2_outputs(612) <= not(layer1_outputs(5573)) or (layer1_outputs(10504));
    layer2_outputs(613) <= not(layer1_outputs(12779)) or (layer1_outputs(1225));
    layer2_outputs(614) <= layer1_outputs(6714);
    layer2_outputs(615) <= layer1_outputs(481);
    layer2_outputs(616) <= (layer1_outputs(11989)) xor (layer1_outputs(11771));
    layer2_outputs(617) <= layer1_outputs(10776);
    layer2_outputs(618) <= not(layer1_outputs(2397));
    layer2_outputs(619) <= (layer1_outputs(4057)) or (layer1_outputs(11102));
    layer2_outputs(620) <= (layer1_outputs(2363)) xor (layer1_outputs(3385));
    layer2_outputs(621) <= (layer1_outputs(4357)) xor (layer1_outputs(9275));
    layer2_outputs(622) <= not(layer1_outputs(6541)) or (layer1_outputs(11233));
    layer2_outputs(623) <= not((layer1_outputs(6813)) or (layer1_outputs(12754)));
    layer2_outputs(624) <= not(layer1_outputs(12718));
    layer2_outputs(625) <= not(layer1_outputs(10704)) or (layer1_outputs(11216));
    layer2_outputs(626) <= (layer1_outputs(2706)) and (layer1_outputs(10126));
    layer2_outputs(627) <= layer1_outputs(2039);
    layer2_outputs(628) <= not(layer1_outputs(3500));
    layer2_outputs(629) <= not(layer1_outputs(1173));
    layer2_outputs(630) <= not(layer1_outputs(10688));
    layer2_outputs(631) <= (layer1_outputs(3918)) xor (layer1_outputs(11278));
    layer2_outputs(632) <= '1';
    layer2_outputs(633) <= not(layer1_outputs(2077));
    layer2_outputs(634) <= not(layer1_outputs(1708));
    layer2_outputs(635) <= not(layer1_outputs(4148));
    layer2_outputs(636) <= layer1_outputs(5606);
    layer2_outputs(637) <= not(layer1_outputs(12328)) or (layer1_outputs(8137));
    layer2_outputs(638) <= layer1_outputs(5396);
    layer2_outputs(639) <= (layer1_outputs(11110)) and not (layer1_outputs(3668));
    layer2_outputs(640) <= layer1_outputs(4510);
    layer2_outputs(641) <= not((layer1_outputs(861)) or (layer1_outputs(10904)));
    layer2_outputs(642) <= layer1_outputs(6737);
    layer2_outputs(643) <= layer1_outputs(4680);
    layer2_outputs(644) <= not(layer1_outputs(4433));
    layer2_outputs(645) <= not((layer1_outputs(10049)) xor (layer1_outputs(11444)));
    layer2_outputs(646) <= not(layer1_outputs(5127));
    layer2_outputs(647) <= not(layer1_outputs(12314)) or (layer1_outputs(2592));
    layer2_outputs(648) <= (layer1_outputs(5809)) and (layer1_outputs(9316));
    layer2_outputs(649) <= not(layer1_outputs(12778));
    layer2_outputs(650) <= not(layer1_outputs(4405));
    layer2_outputs(651) <= layer1_outputs(8329);
    layer2_outputs(652) <= (layer1_outputs(5523)) and (layer1_outputs(9877));
    layer2_outputs(653) <= (layer1_outputs(3106)) and not (layer1_outputs(9452));
    layer2_outputs(654) <= not(layer1_outputs(7977)) or (layer1_outputs(2400));
    layer2_outputs(655) <= layer1_outputs(11583);
    layer2_outputs(656) <= not(layer1_outputs(4011));
    layer2_outputs(657) <= not(layer1_outputs(6952));
    layer2_outputs(658) <= (layer1_outputs(7315)) and (layer1_outputs(5254));
    layer2_outputs(659) <= not((layer1_outputs(9069)) and (layer1_outputs(5254)));
    layer2_outputs(660) <= not(layer1_outputs(3059));
    layer2_outputs(661) <= (layer1_outputs(10940)) and not (layer1_outputs(4402));
    layer2_outputs(662) <= not(layer1_outputs(11469)) or (layer1_outputs(3850));
    layer2_outputs(663) <= layer1_outputs(4516);
    layer2_outputs(664) <= not(layer1_outputs(9154));
    layer2_outputs(665) <= not(layer1_outputs(2279));
    layer2_outputs(666) <= not((layer1_outputs(4440)) xor (layer1_outputs(5954)));
    layer2_outputs(667) <= layer1_outputs(748);
    layer2_outputs(668) <= (layer1_outputs(3442)) or (layer1_outputs(3188));
    layer2_outputs(669) <= (layer1_outputs(6181)) and not (layer1_outputs(7968));
    layer2_outputs(670) <= not((layer1_outputs(4884)) or (layer1_outputs(6904)));
    layer2_outputs(671) <= not((layer1_outputs(8709)) xor (layer1_outputs(42)));
    layer2_outputs(672) <= (layer1_outputs(10158)) and (layer1_outputs(667));
    layer2_outputs(673) <= layer1_outputs(6850);
    layer2_outputs(674) <= not((layer1_outputs(12495)) or (layer1_outputs(4473)));
    layer2_outputs(675) <= layer1_outputs(11643);
    layer2_outputs(676) <= not(layer1_outputs(10433));
    layer2_outputs(677) <= (layer1_outputs(11810)) and not (layer1_outputs(8165));
    layer2_outputs(678) <= not((layer1_outputs(4158)) and (layer1_outputs(12510)));
    layer2_outputs(679) <= not(layer1_outputs(4604)) or (layer1_outputs(2161));
    layer2_outputs(680) <= not((layer1_outputs(9981)) and (layer1_outputs(8637)));
    layer2_outputs(681) <= not(layer1_outputs(2175)) or (layer1_outputs(11957));
    layer2_outputs(682) <= layer1_outputs(6872);
    layer2_outputs(683) <= not((layer1_outputs(1682)) or (layer1_outputs(3650)));
    layer2_outputs(684) <= (layer1_outputs(5745)) and not (layer1_outputs(4597));
    layer2_outputs(685) <= not(layer1_outputs(10095));
    layer2_outputs(686) <= not(layer1_outputs(8945));
    layer2_outputs(687) <= layer1_outputs(4226);
    layer2_outputs(688) <= (layer1_outputs(5496)) or (layer1_outputs(3727));
    layer2_outputs(689) <= not(layer1_outputs(7616)) or (layer1_outputs(668));
    layer2_outputs(690) <= not(layer1_outputs(4516));
    layer2_outputs(691) <= (layer1_outputs(11558)) and not (layer1_outputs(11003));
    layer2_outputs(692) <= not((layer1_outputs(948)) and (layer1_outputs(6233)));
    layer2_outputs(693) <= not(layer1_outputs(9724));
    layer2_outputs(694) <= layer1_outputs(2332);
    layer2_outputs(695) <= layer1_outputs(5575);
    layer2_outputs(696) <= layer1_outputs(4123);
    layer2_outputs(697) <= not(layer1_outputs(6449)) or (layer1_outputs(3894));
    layer2_outputs(698) <= not((layer1_outputs(12193)) xor (layer1_outputs(4871)));
    layer2_outputs(699) <= not(layer1_outputs(6341));
    layer2_outputs(700) <= layer1_outputs(6251);
    layer2_outputs(701) <= not((layer1_outputs(7657)) or (layer1_outputs(1076)));
    layer2_outputs(702) <= not(layer1_outputs(9772)) or (layer1_outputs(6666));
    layer2_outputs(703) <= (layer1_outputs(1282)) xor (layer1_outputs(6727));
    layer2_outputs(704) <= layer1_outputs(9474);
    layer2_outputs(705) <= (layer1_outputs(10315)) xor (layer1_outputs(8505));
    layer2_outputs(706) <= not((layer1_outputs(3760)) xor (layer1_outputs(9567)));
    layer2_outputs(707) <= '0';
    layer2_outputs(708) <= layer1_outputs(1074);
    layer2_outputs(709) <= not(layer1_outputs(12600));
    layer2_outputs(710) <= not(layer1_outputs(11575));
    layer2_outputs(711) <= not(layer1_outputs(771));
    layer2_outputs(712) <= layer1_outputs(4865);
    layer2_outputs(713) <= (layer1_outputs(7974)) xor (layer1_outputs(9345));
    layer2_outputs(714) <= (layer1_outputs(9932)) or (layer1_outputs(7398));
    layer2_outputs(715) <= layer1_outputs(8859);
    layer2_outputs(716) <= not((layer1_outputs(3826)) and (layer1_outputs(5674)));
    layer2_outputs(717) <= (layer1_outputs(12095)) and (layer1_outputs(3052));
    layer2_outputs(718) <= not((layer1_outputs(11881)) and (layer1_outputs(7791)));
    layer2_outputs(719) <= (layer1_outputs(5902)) and (layer1_outputs(5010));
    layer2_outputs(720) <= (layer1_outputs(9013)) or (layer1_outputs(11664));
    layer2_outputs(721) <= layer1_outputs(9158);
    layer2_outputs(722) <= layer1_outputs(1146);
    layer2_outputs(723) <= layer1_outputs(6366);
    layer2_outputs(724) <= (layer1_outputs(6595)) xor (layer1_outputs(2093));
    layer2_outputs(725) <= (layer1_outputs(3929)) and not (layer1_outputs(7882));
    layer2_outputs(726) <= (layer1_outputs(8623)) and (layer1_outputs(8093));
    layer2_outputs(727) <= layer1_outputs(6915);
    layer2_outputs(728) <= not(layer1_outputs(11590));
    layer2_outputs(729) <= '0';
    layer2_outputs(730) <= (layer1_outputs(2491)) and (layer1_outputs(477));
    layer2_outputs(731) <= not(layer1_outputs(2717)) or (layer1_outputs(1014));
    layer2_outputs(732) <= not(layer1_outputs(1764)) or (layer1_outputs(232));
    layer2_outputs(733) <= not(layer1_outputs(3878));
    layer2_outputs(734) <= not(layer1_outputs(2399));
    layer2_outputs(735) <= (layer1_outputs(1142)) xor (layer1_outputs(7750));
    layer2_outputs(736) <= (layer1_outputs(1763)) xor (layer1_outputs(8949));
    layer2_outputs(737) <= not(layer1_outputs(3903));
    layer2_outputs(738) <= (layer1_outputs(1828)) and not (layer1_outputs(12731));
    layer2_outputs(739) <= layer1_outputs(7999);
    layer2_outputs(740) <= (layer1_outputs(2465)) and (layer1_outputs(5420));
    layer2_outputs(741) <= layer1_outputs(3050);
    layer2_outputs(742) <= not((layer1_outputs(5351)) and (layer1_outputs(2572)));
    layer2_outputs(743) <= not(layer1_outputs(3533));
    layer2_outputs(744) <= layer1_outputs(1782);
    layer2_outputs(745) <= layer1_outputs(6949);
    layer2_outputs(746) <= not(layer1_outputs(1182)) or (layer1_outputs(6494));
    layer2_outputs(747) <= not((layer1_outputs(37)) xor (layer1_outputs(7287)));
    layer2_outputs(748) <= not(layer1_outputs(8367)) or (layer1_outputs(6203));
    layer2_outputs(749) <= not((layer1_outputs(11867)) and (layer1_outputs(3844)));
    layer2_outputs(750) <= (layer1_outputs(6346)) or (layer1_outputs(8547));
    layer2_outputs(751) <= not(layer1_outputs(1996));
    layer2_outputs(752) <= not(layer1_outputs(9449));
    layer2_outputs(753) <= (layer1_outputs(12675)) or (layer1_outputs(4916));
    layer2_outputs(754) <= not(layer1_outputs(1287)) or (layer1_outputs(703));
    layer2_outputs(755) <= not(layer1_outputs(566)) or (layer1_outputs(8452));
    layer2_outputs(756) <= layer1_outputs(488);
    layer2_outputs(757) <= not(layer1_outputs(12615)) or (layer1_outputs(10816));
    layer2_outputs(758) <= (layer1_outputs(9753)) xor (layer1_outputs(9049));
    layer2_outputs(759) <= layer1_outputs(487);
    layer2_outputs(760) <= not((layer1_outputs(8051)) or (layer1_outputs(10824)));
    layer2_outputs(761) <= not((layer1_outputs(6863)) xor (layer1_outputs(4650)));
    layer2_outputs(762) <= layer1_outputs(1866);
    layer2_outputs(763) <= not((layer1_outputs(5055)) or (layer1_outputs(3755)));
    layer2_outputs(764) <= not(layer1_outputs(757));
    layer2_outputs(765) <= not(layer1_outputs(2330)) or (layer1_outputs(12098));
    layer2_outputs(766) <= (layer1_outputs(6031)) or (layer1_outputs(11758));
    layer2_outputs(767) <= not((layer1_outputs(10722)) and (layer1_outputs(10985)));
    layer2_outputs(768) <= layer1_outputs(1249);
    layer2_outputs(769) <= not((layer1_outputs(124)) and (layer1_outputs(3181)));
    layer2_outputs(770) <= not(layer1_outputs(2641)) or (layer1_outputs(1846));
    layer2_outputs(771) <= '0';
    layer2_outputs(772) <= layer1_outputs(7918);
    layer2_outputs(773) <= not(layer1_outputs(413));
    layer2_outputs(774) <= not((layer1_outputs(3697)) or (layer1_outputs(365)));
    layer2_outputs(775) <= not(layer1_outputs(4497));
    layer2_outputs(776) <= (layer1_outputs(2543)) xor (layer1_outputs(7894));
    layer2_outputs(777) <= layer1_outputs(10726);
    layer2_outputs(778) <= layer1_outputs(1900);
    layer2_outputs(779) <= (layer1_outputs(2532)) xor (layer1_outputs(110));
    layer2_outputs(780) <= not((layer1_outputs(2838)) and (layer1_outputs(2873)));
    layer2_outputs(781) <= not(layer1_outputs(46)) or (layer1_outputs(4331));
    layer2_outputs(782) <= (layer1_outputs(10532)) and not (layer1_outputs(8994));
    layer2_outputs(783) <= layer1_outputs(2253);
    layer2_outputs(784) <= not(layer1_outputs(9633));
    layer2_outputs(785) <= (layer1_outputs(5073)) and (layer1_outputs(12273));
    layer2_outputs(786) <= layer1_outputs(9620);
    layer2_outputs(787) <= layer1_outputs(4972);
    layer2_outputs(788) <= layer1_outputs(8814);
    layer2_outputs(789) <= not(layer1_outputs(2530)) or (layer1_outputs(1049));
    layer2_outputs(790) <= layer1_outputs(303);
    layer2_outputs(791) <= not(layer1_outputs(11643));
    layer2_outputs(792) <= (layer1_outputs(9807)) and not (layer1_outputs(2321));
    layer2_outputs(793) <= (layer1_outputs(11266)) xor (layer1_outputs(958));
    layer2_outputs(794) <= not((layer1_outputs(7970)) and (layer1_outputs(1296)));
    layer2_outputs(795) <= layer1_outputs(11001);
    layer2_outputs(796) <= (layer1_outputs(4262)) and not (layer1_outputs(11650));
    layer2_outputs(797) <= not((layer1_outputs(11766)) xor (layer1_outputs(145)));
    layer2_outputs(798) <= not((layer1_outputs(5978)) xor (layer1_outputs(10926)));
    layer2_outputs(799) <= (layer1_outputs(9882)) xor (layer1_outputs(6510));
    layer2_outputs(800) <= not(layer1_outputs(8075));
    layer2_outputs(801) <= not(layer1_outputs(8645));
    layer2_outputs(802) <= '1';
    layer2_outputs(803) <= not((layer1_outputs(9642)) and (layer1_outputs(4131)));
    layer2_outputs(804) <= layer1_outputs(10638);
    layer2_outputs(805) <= not((layer1_outputs(12796)) xor (layer1_outputs(8980)));
    layer2_outputs(806) <= not((layer1_outputs(5377)) xor (layer1_outputs(10869)));
    layer2_outputs(807) <= not((layer1_outputs(6974)) and (layer1_outputs(760)));
    layer2_outputs(808) <= not(layer1_outputs(3568));
    layer2_outputs(809) <= layer1_outputs(11031);
    layer2_outputs(810) <= not(layer1_outputs(3685));
    layer2_outputs(811) <= (layer1_outputs(9320)) or (layer1_outputs(3340));
    layer2_outputs(812) <= layer1_outputs(6051);
    layer2_outputs(813) <= not(layer1_outputs(9161)) or (layer1_outputs(6623));
    layer2_outputs(814) <= (layer1_outputs(1688)) and not (layer1_outputs(1764));
    layer2_outputs(815) <= not((layer1_outputs(2634)) xor (layer1_outputs(7197)));
    layer2_outputs(816) <= layer1_outputs(5790);
    layer2_outputs(817) <= not(layer1_outputs(8991));
    layer2_outputs(818) <= not((layer1_outputs(1246)) xor (layer1_outputs(4077)));
    layer2_outputs(819) <= not((layer1_outputs(10992)) or (layer1_outputs(12518)));
    layer2_outputs(820) <= (layer1_outputs(6241)) and not (layer1_outputs(1317));
    layer2_outputs(821) <= not((layer1_outputs(8931)) xor (layer1_outputs(11900)));
    layer2_outputs(822) <= layer1_outputs(784);
    layer2_outputs(823) <= not(layer1_outputs(7265)) or (layer1_outputs(3257));
    layer2_outputs(824) <= layer1_outputs(1699);
    layer2_outputs(825) <= not(layer1_outputs(2580)) or (layer1_outputs(3014));
    layer2_outputs(826) <= (layer1_outputs(3274)) xor (layer1_outputs(2281));
    layer2_outputs(827) <= not(layer1_outputs(11366)) or (layer1_outputs(8029));
    layer2_outputs(828) <= layer1_outputs(7554);
    layer2_outputs(829) <= layer1_outputs(7680);
    layer2_outputs(830) <= (layer1_outputs(10566)) and not (layer1_outputs(4055));
    layer2_outputs(831) <= not(layer1_outputs(4632)) or (layer1_outputs(1632));
    layer2_outputs(832) <= (layer1_outputs(1050)) and not (layer1_outputs(8389));
    layer2_outputs(833) <= not((layer1_outputs(2541)) or (layer1_outputs(6047)));
    layer2_outputs(834) <= '1';
    layer2_outputs(835) <= layer1_outputs(7011);
    layer2_outputs(836) <= not(layer1_outputs(1061));
    layer2_outputs(837) <= layer1_outputs(11730);
    layer2_outputs(838) <= layer1_outputs(2883);
    layer2_outputs(839) <= layer1_outputs(8186);
    layer2_outputs(840) <= layer1_outputs(7733);
    layer2_outputs(841) <= not(layer1_outputs(10912));
    layer2_outputs(842) <= layer1_outputs(7639);
    layer2_outputs(843) <= layer1_outputs(2458);
    layer2_outputs(844) <= layer1_outputs(5289);
    layer2_outputs(845) <= not((layer1_outputs(9332)) xor (layer1_outputs(12191)));
    layer2_outputs(846) <= (layer1_outputs(4665)) and not (layer1_outputs(3000));
    layer2_outputs(847) <= not((layer1_outputs(8917)) xor (layer1_outputs(9259)));
    layer2_outputs(848) <= not((layer1_outputs(5568)) or (layer1_outputs(402)));
    layer2_outputs(849) <= not(layer1_outputs(3990));
    layer2_outputs(850) <= not(layer1_outputs(12127));
    layer2_outputs(851) <= not((layer1_outputs(12411)) and (layer1_outputs(9296)));
    layer2_outputs(852) <= layer1_outputs(10705);
    layer2_outputs(853) <= layer1_outputs(8413);
    layer2_outputs(854) <= layer1_outputs(2561);
    layer2_outputs(855) <= not(layer1_outputs(1947));
    layer2_outputs(856) <= layer1_outputs(1124);
    layer2_outputs(857) <= (layer1_outputs(10252)) or (layer1_outputs(2771));
    layer2_outputs(858) <= (layer1_outputs(10067)) and not (layer1_outputs(7226));
    layer2_outputs(859) <= not(layer1_outputs(12281));
    layer2_outputs(860) <= not(layer1_outputs(9747));
    layer2_outputs(861) <= '0';
    layer2_outputs(862) <= not((layer1_outputs(2613)) or (layer1_outputs(3160)));
    layer2_outputs(863) <= layer1_outputs(8555);
    layer2_outputs(864) <= not(layer1_outputs(5441));
    layer2_outputs(865) <= layer1_outputs(1498);
    layer2_outputs(866) <= (layer1_outputs(4647)) xor (layer1_outputs(8741));
    layer2_outputs(867) <= layer1_outputs(12406);
    layer2_outputs(868) <= not(layer1_outputs(6777));
    layer2_outputs(869) <= not((layer1_outputs(9735)) or (layer1_outputs(5915)));
    layer2_outputs(870) <= not(layer1_outputs(11172));
    layer2_outputs(871) <= not(layer1_outputs(9056));
    layer2_outputs(872) <= not(layer1_outputs(6741));
    layer2_outputs(873) <= (layer1_outputs(12079)) and not (layer1_outputs(4051));
    layer2_outputs(874) <= (layer1_outputs(1943)) and not (layer1_outputs(11432));
    layer2_outputs(875) <= not((layer1_outputs(9730)) or (layer1_outputs(6999)));
    layer2_outputs(876) <= (layer1_outputs(9274)) and (layer1_outputs(9956));
    layer2_outputs(877) <= not((layer1_outputs(5622)) or (layer1_outputs(8351)));
    layer2_outputs(878) <= not((layer1_outputs(6413)) xor (layer1_outputs(25)));
    layer2_outputs(879) <= not(layer1_outputs(7560));
    layer2_outputs(880) <= not(layer1_outputs(5083));
    layer2_outputs(881) <= layer1_outputs(6340);
    layer2_outputs(882) <= not((layer1_outputs(812)) and (layer1_outputs(5849)));
    layer2_outputs(883) <= not((layer1_outputs(2403)) xor (layer1_outputs(7281)));
    layer2_outputs(884) <= not(layer1_outputs(1797)) or (layer1_outputs(3198));
    layer2_outputs(885) <= layer1_outputs(64);
    layer2_outputs(886) <= layer1_outputs(4914);
    layer2_outputs(887) <= (layer1_outputs(8431)) and (layer1_outputs(11488));
    layer2_outputs(888) <= (layer1_outputs(11826)) and (layer1_outputs(6683));
    layer2_outputs(889) <= layer1_outputs(7906);
    layer2_outputs(890) <= (layer1_outputs(3913)) and not (layer1_outputs(546));
    layer2_outputs(891) <= not((layer1_outputs(3793)) xor (layer1_outputs(9860)));
    layer2_outputs(892) <= layer1_outputs(2875);
    layer2_outputs(893) <= (layer1_outputs(10955)) and not (layer1_outputs(3080));
    layer2_outputs(894) <= (layer1_outputs(12324)) and not (layer1_outputs(7036));
    layer2_outputs(895) <= not(layer1_outputs(1514));
    layer2_outputs(896) <= not(layer1_outputs(8759));
    layer2_outputs(897) <= not(layer1_outputs(5280));
    layer2_outputs(898) <= layer1_outputs(985);
    layer2_outputs(899) <= not((layer1_outputs(6505)) and (layer1_outputs(5193)));
    layer2_outputs(900) <= not((layer1_outputs(2381)) xor (layer1_outputs(810)));
    layer2_outputs(901) <= (layer1_outputs(11780)) and not (layer1_outputs(5091));
    layer2_outputs(902) <= not(layer1_outputs(2212));
    layer2_outputs(903) <= (layer1_outputs(5808)) and not (layer1_outputs(4817));
    layer2_outputs(904) <= layer1_outputs(12562);
    layer2_outputs(905) <= layer1_outputs(8026);
    layer2_outputs(906) <= (layer1_outputs(1192)) and not (layer1_outputs(6903));
    layer2_outputs(907) <= not(layer1_outputs(3042));
    layer2_outputs(908) <= (layer1_outputs(5223)) and (layer1_outputs(8774));
    layer2_outputs(909) <= not(layer1_outputs(11454)) or (layer1_outputs(3485));
    layer2_outputs(910) <= (layer1_outputs(11817)) xor (layer1_outputs(9733));
    layer2_outputs(911) <= (layer1_outputs(8553)) and not (layer1_outputs(10301));
    layer2_outputs(912) <= not(layer1_outputs(8283));
    layer2_outputs(913) <= layer1_outputs(11430);
    layer2_outputs(914) <= (layer1_outputs(4562)) xor (layer1_outputs(3524));
    layer2_outputs(915) <= not(layer1_outputs(4407));
    layer2_outputs(916) <= not((layer1_outputs(1719)) and (layer1_outputs(6588)));
    layer2_outputs(917) <= not(layer1_outputs(1702)) or (layer1_outputs(11577));
    layer2_outputs(918) <= layer1_outputs(8915);
    layer2_outputs(919) <= not((layer1_outputs(5992)) or (layer1_outputs(6396)));
    layer2_outputs(920) <= not(layer1_outputs(6584));
    layer2_outputs(921) <= not(layer1_outputs(4915));
    layer2_outputs(922) <= (layer1_outputs(4030)) or (layer1_outputs(11371));
    layer2_outputs(923) <= (layer1_outputs(888)) xor (layer1_outputs(2686));
    layer2_outputs(924) <= not(layer1_outputs(8066));
    layer2_outputs(925) <= (layer1_outputs(5649)) and not (layer1_outputs(12486));
    layer2_outputs(926) <= not((layer1_outputs(3743)) xor (layer1_outputs(12227)));
    layer2_outputs(927) <= (layer1_outputs(5703)) and not (layer1_outputs(7324));
    layer2_outputs(928) <= not(layer1_outputs(1991)) or (layer1_outputs(7772));
    layer2_outputs(929) <= not(layer1_outputs(7547));
    layer2_outputs(930) <= not(layer1_outputs(2576));
    layer2_outputs(931) <= layer1_outputs(10412);
    layer2_outputs(932) <= not(layer1_outputs(763)) or (layer1_outputs(12075));
    layer2_outputs(933) <= not((layer1_outputs(7790)) xor (layer1_outputs(1524)));
    layer2_outputs(934) <= layer1_outputs(10829);
    layer2_outputs(935) <= '0';
    layer2_outputs(936) <= (layer1_outputs(4743)) and (layer1_outputs(10057));
    layer2_outputs(937) <= not(layer1_outputs(136)) or (layer1_outputs(9135));
    layer2_outputs(938) <= layer1_outputs(6665);
    layer2_outputs(939) <= not(layer1_outputs(1158));
    layer2_outputs(940) <= not(layer1_outputs(7016));
    layer2_outputs(941) <= (layer1_outputs(12276)) or (layer1_outputs(8001));
    layer2_outputs(942) <= (layer1_outputs(6817)) xor (layer1_outputs(550));
    layer2_outputs(943) <= (layer1_outputs(3848)) and not (layer1_outputs(2074));
    layer2_outputs(944) <= not(layer1_outputs(669));
    layer2_outputs(945) <= layer1_outputs(6831);
    layer2_outputs(946) <= not(layer1_outputs(8315));
    layer2_outputs(947) <= (layer1_outputs(5355)) and not (layer1_outputs(4704));
    layer2_outputs(948) <= layer1_outputs(2188);
    layer2_outputs(949) <= '0';
    layer2_outputs(950) <= (layer1_outputs(294)) or (layer1_outputs(12759));
    layer2_outputs(951) <= not(layer1_outputs(8813));
    layer2_outputs(952) <= not(layer1_outputs(10063)) or (layer1_outputs(6070));
    layer2_outputs(953) <= not((layer1_outputs(337)) xor (layer1_outputs(6084)));
    layer2_outputs(954) <= not(layer1_outputs(8132));
    layer2_outputs(955) <= (layer1_outputs(2749)) and (layer1_outputs(5520));
    layer2_outputs(956) <= layer1_outputs(646);
    layer2_outputs(957) <= layer1_outputs(482);
    layer2_outputs(958) <= layer1_outputs(10366);
    layer2_outputs(959) <= not((layer1_outputs(6477)) xor (layer1_outputs(5393)));
    layer2_outputs(960) <= layer1_outputs(11280);
    layer2_outputs(961) <= (layer1_outputs(11291)) and not (layer1_outputs(2271));
    layer2_outputs(962) <= not(layer1_outputs(8519));
    layer2_outputs(963) <= (layer1_outputs(9466)) and not (layer1_outputs(7227));
    layer2_outputs(964) <= layer1_outputs(11370);
    layer2_outputs(965) <= not((layer1_outputs(7723)) xor (layer1_outputs(4004)));
    layer2_outputs(966) <= not((layer1_outputs(3170)) and (layer1_outputs(12088)));
    layer2_outputs(967) <= layer1_outputs(7857);
    layer2_outputs(968) <= (layer1_outputs(4942)) and (layer1_outputs(3005));
    layer2_outputs(969) <= (layer1_outputs(2967)) and not (layer1_outputs(5367));
    layer2_outputs(970) <= (layer1_outputs(7900)) xor (layer1_outputs(4550));
    layer2_outputs(971) <= not(layer1_outputs(10766));
    layer2_outputs(972) <= layer1_outputs(12284);
    layer2_outputs(973) <= (layer1_outputs(4998)) and not (layer1_outputs(10794));
    layer2_outputs(974) <= not((layer1_outputs(10255)) xor (layer1_outputs(582)));
    layer2_outputs(975) <= layer1_outputs(713);
    layer2_outputs(976) <= not((layer1_outputs(5444)) xor (layer1_outputs(5901)));
    layer2_outputs(977) <= not(layer1_outputs(241));
    layer2_outputs(978) <= layer1_outputs(9104);
    layer2_outputs(979) <= not(layer1_outputs(11283)) or (layer1_outputs(4058));
    layer2_outputs(980) <= '0';
    layer2_outputs(981) <= layer1_outputs(6041);
    layer2_outputs(982) <= not(layer1_outputs(11969));
    layer2_outputs(983) <= (layer1_outputs(7031)) xor (layer1_outputs(2968));
    layer2_outputs(984) <= (layer1_outputs(10136)) xor (layer1_outputs(7597));
    layer2_outputs(985) <= layer1_outputs(2076);
    layer2_outputs(986) <= not(layer1_outputs(9961)) or (layer1_outputs(4773));
    layer2_outputs(987) <= (layer1_outputs(1313)) xor (layer1_outputs(610));
    layer2_outputs(988) <= not((layer1_outputs(6130)) or (layer1_outputs(3483)));
    layer2_outputs(989) <= (layer1_outputs(2074)) xor (layer1_outputs(11830));
    layer2_outputs(990) <= not(layer1_outputs(9342));
    layer2_outputs(991) <= not(layer1_outputs(4434)) or (layer1_outputs(1946));
    layer2_outputs(992) <= (layer1_outputs(7487)) and not (layer1_outputs(5898));
    layer2_outputs(993) <= layer1_outputs(9646);
    layer2_outputs(994) <= layer1_outputs(7481);
    layer2_outputs(995) <= (layer1_outputs(3224)) xor (layer1_outputs(8711));
    layer2_outputs(996) <= (layer1_outputs(11710)) xor (layer1_outputs(10085));
    layer2_outputs(997) <= layer1_outputs(10787);
    layer2_outputs(998) <= not(layer1_outputs(3665)) or (layer1_outputs(7171));
    layer2_outputs(999) <= layer1_outputs(3710);
    layer2_outputs(1000) <= not(layer1_outputs(4608));
    layer2_outputs(1001) <= not(layer1_outputs(10543));
    layer2_outputs(1002) <= (layer1_outputs(6868)) xor (layer1_outputs(2369));
    layer2_outputs(1003) <= (layer1_outputs(12443)) or (layer1_outputs(10293));
    layer2_outputs(1004) <= not((layer1_outputs(10735)) or (layer1_outputs(9770)));
    layer2_outputs(1005) <= not((layer1_outputs(1062)) or (layer1_outputs(10413)));
    layer2_outputs(1006) <= not(layer1_outputs(3196));
    layer2_outputs(1007) <= not(layer1_outputs(11334)) or (layer1_outputs(3146));
    layer2_outputs(1008) <= (layer1_outputs(11737)) xor (layer1_outputs(3001));
    layer2_outputs(1009) <= layer1_outputs(5947);
    layer2_outputs(1010) <= not(layer1_outputs(2791));
    layer2_outputs(1011) <= (layer1_outputs(3857)) and not (layer1_outputs(5473));
    layer2_outputs(1012) <= not(layer1_outputs(11350));
    layer2_outputs(1013) <= layer1_outputs(11806);
    layer2_outputs(1014) <= layer1_outputs(9741);
    layer2_outputs(1015) <= (layer1_outputs(8575)) xor (layer1_outputs(10786));
    layer2_outputs(1016) <= layer1_outputs(9930);
    layer2_outputs(1017) <= layer1_outputs(11222);
    layer2_outputs(1018) <= not(layer1_outputs(5467));
    layer2_outputs(1019) <= layer1_outputs(9837);
    layer2_outputs(1020) <= not(layer1_outputs(5179));
    layer2_outputs(1021) <= not(layer1_outputs(3703));
    layer2_outputs(1022) <= (layer1_outputs(10221)) and not (layer1_outputs(10034));
    layer2_outputs(1023) <= layer1_outputs(1583);
    layer2_outputs(1024) <= not(layer1_outputs(12082));
    layer2_outputs(1025) <= not(layer1_outputs(1417));
    layer2_outputs(1026) <= layer1_outputs(8053);
    layer2_outputs(1027) <= not(layer1_outputs(3300));
    layer2_outputs(1028) <= not(layer1_outputs(4856)) or (layer1_outputs(12049));
    layer2_outputs(1029) <= not(layer1_outputs(8074));
    layer2_outputs(1030) <= layer1_outputs(11987);
    layer2_outputs(1031) <= layer1_outputs(250);
    layer2_outputs(1032) <= (layer1_outputs(12574)) and not (layer1_outputs(7397));
    layer2_outputs(1033) <= not(layer1_outputs(9106));
    layer2_outputs(1034) <= (layer1_outputs(6006)) or (layer1_outputs(1246));
    layer2_outputs(1035) <= not(layer1_outputs(5070)) or (layer1_outputs(12195));
    layer2_outputs(1036) <= (layer1_outputs(3749)) or (layer1_outputs(4660));
    layer2_outputs(1037) <= (layer1_outputs(5981)) or (layer1_outputs(2102));
    layer2_outputs(1038) <= (layer1_outputs(3803)) xor (layer1_outputs(8492));
    layer2_outputs(1039) <= (layer1_outputs(7403)) or (layer1_outputs(204));
    layer2_outputs(1040) <= layer1_outputs(1695);
    layer2_outputs(1041) <= (layer1_outputs(617)) and not (layer1_outputs(5510));
    layer2_outputs(1042) <= not((layer1_outputs(10403)) or (layer1_outputs(9812)));
    layer2_outputs(1043) <= (layer1_outputs(144)) and (layer1_outputs(7580));
    layer2_outputs(1044) <= not((layer1_outputs(10935)) or (layer1_outputs(1289)));
    layer2_outputs(1045) <= not((layer1_outputs(10671)) xor (layer1_outputs(5932)));
    layer2_outputs(1046) <= not((layer1_outputs(7885)) xor (layer1_outputs(412)));
    layer2_outputs(1047) <= (layer1_outputs(4941)) or (layer1_outputs(6580));
    layer2_outputs(1048) <= not((layer1_outputs(12327)) and (layer1_outputs(4207)));
    layer2_outputs(1049) <= not(layer1_outputs(10606));
    layer2_outputs(1050) <= not(layer1_outputs(4404));
    layer2_outputs(1051) <= not(layer1_outputs(4766));
    layer2_outputs(1052) <= layer1_outputs(10330);
    layer2_outputs(1053) <= not((layer1_outputs(8533)) or (layer1_outputs(1229)));
    layer2_outputs(1054) <= not(layer1_outputs(10282)) or (layer1_outputs(5489));
    layer2_outputs(1055) <= layer1_outputs(2593);
    layer2_outputs(1056) <= not(layer1_outputs(790));
    layer2_outputs(1057) <= not(layer1_outputs(10980));
    layer2_outputs(1058) <= not(layer1_outputs(913));
    layer2_outputs(1059) <= (layer1_outputs(166)) and not (layer1_outputs(5829));
    layer2_outputs(1060) <= not(layer1_outputs(1388));
    layer2_outputs(1061) <= not(layer1_outputs(11940));
    layer2_outputs(1062) <= not((layer1_outputs(6542)) and (layer1_outputs(12659)));
    layer2_outputs(1063) <= layer1_outputs(9273);
    layer2_outputs(1064) <= not(layer1_outputs(121));
    layer2_outputs(1065) <= (layer1_outputs(3019)) and not (layer1_outputs(2137));
    layer2_outputs(1066) <= layer1_outputs(10876);
    layer2_outputs(1067) <= not(layer1_outputs(6907));
    layer2_outputs(1068) <= not(layer1_outputs(11842)) or (layer1_outputs(3870));
    layer2_outputs(1069) <= (layer1_outputs(10540)) and not (layer1_outputs(7365));
    layer2_outputs(1070) <= not(layer1_outputs(5140)) or (layer1_outputs(11761));
    layer2_outputs(1071) <= not(layer1_outputs(2667));
    layer2_outputs(1072) <= (layer1_outputs(5451)) and not (layer1_outputs(3398));
    layer2_outputs(1073) <= layer1_outputs(102);
    layer2_outputs(1074) <= (layer1_outputs(9163)) and (layer1_outputs(9706));
    layer2_outputs(1075) <= (layer1_outputs(11314)) and not (layer1_outputs(8241));
    layer2_outputs(1076) <= not(layer1_outputs(7603));
    layer2_outputs(1077) <= layer1_outputs(1188);
    layer2_outputs(1078) <= layer1_outputs(6200);
    layer2_outputs(1079) <= not((layer1_outputs(61)) and (layer1_outputs(598)));
    layer2_outputs(1080) <= layer1_outputs(5846);
    layer2_outputs(1081) <= not(layer1_outputs(9536));
    layer2_outputs(1082) <= not(layer1_outputs(6501));
    layer2_outputs(1083) <= '1';
    layer2_outputs(1084) <= not(layer1_outputs(8762)) or (layer1_outputs(8101));
    layer2_outputs(1085) <= not(layer1_outputs(6418));
    layer2_outputs(1086) <= not(layer1_outputs(7454));
    layer2_outputs(1087) <= not(layer1_outputs(6819));
    layer2_outputs(1088) <= not(layer1_outputs(8581));
    layer2_outputs(1089) <= not(layer1_outputs(2098));
    layer2_outputs(1090) <= layer1_outputs(2027);
    layer2_outputs(1091) <= (layer1_outputs(8828)) or (layer1_outputs(7784));
    layer2_outputs(1092) <= layer1_outputs(2006);
    layer2_outputs(1093) <= (layer1_outputs(10971)) xor (layer1_outputs(7560));
    layer2_outputs(1094) <= not(layer1_outputs(1826));
    layer2_outputs(1095) <= (layer1_outputs(9554)) xor (layer1_outputs(11601));
    layer2_outputs(1096) <= not(layer1_outputs(11571));
    layer2_outputs(1097) <= not((layer1_outputs(6149)) xor (layer1_outputs(9759)));
    layer2_outputs(1098) <= (layer1_outputs(7490)) xor (layer1_outputs(11706));
    layer2_outputs(1099) <= '1';
    layer2_outputs(1100) <= not((layer1_outputs(12648)) xor (layer1_outputs(7114)));
    layer2_outputs(1101) <= not(layer1_outputs(8733)) or (layer1_outputs(8749));
    layer2_outputs(1102) <= layer1_outputs(10236);
    layer2_outputs(1103) <= not(layer1_outputs(1215));
    layer2_outputs(1104) <= not(layer1_outputs(946));
    layer2_outputs(1105) <= layer1_outputs(11984);
    layer2_outputs(1106) <= (layer1_outputs(7267)) xor (layer1_outputs(10369));
    layer2_outputs(1107) <= not(layer1_outputs(11416));
    layer2_outputs(1108) <= not((layer1_outputs(10515)) xor (layer1_outputs(2191)));
    layer2_outputs(1109) <= (layer1_outputs(3280)) or (layer1_outputs(2142));
    layer2_outputs(1110) <= (layer1_outputs(1302)) and not (layer1_outputs(7070));
    layer2_outputs(1111) <= (layer1_outputs(2055)) and not (layer1_outputs(8434));
    layer2_outputs(1112) <= layer1_outputs(10805);
    layer2_outputs(1113) <= not((layer1_outputs(956)) xor (layer1_outputs(10141)));
    layer2_outputs(1114) <= (layer1_outputs(2403)) and (layer1_outputs(1230));
    layer2_outputs(1115) <= not((layer1_outputs(2388)) xor (layer1_outputs(11181)));
    layer2_outputs(1116) <= not((layer1_outputs(1193)) and (layer1_outputs(4834)));
    layer2_outputs(1117) <= not(layer1_outputs(10396));
    layer2_outputs(1118) <= not(layer1_outputs(7175));
    layer2_outputs(1119) <= not(layer1_outputs(309));
    layer2_outputs(1120) <= not(layer1_outputs(4468));
    layer2_outputs(1121) <= layer1_outputs(1484);
    layer2_outputs(1122) <= (layer1_outputs(2987)) and (layer1_outputs(10055));
    layer2_outputs(1123) <= (layer1_outputs(7008)) and (layer1_outputs(8273));
    layer2_outputs(1124) <= not(layer1_outputs(4966));
    layer2_outputs(1125) <= (layer1_outputs(6712)) and (layer1_outputs(6824));
    layer2_outputs(1126) <= layer1_outputs(165);
    layer2_outputs(1127) <= not(layer1_outputs(4277));
    layer2_outputs(1128) <= not(layer1_outputs(1159));
    layer2_outputs(1129) <= (layer1_outputs(6872)) or (layer1_outputs(8032));
    layer2_outputs(1130) <= not(layer1_outputs(12017));
    layer2_outputs(1131) <= not(layer1_outputs(773));
    layer2_outputs(1132) <= (layer1_outputs(6195)) xor (layer1_outputs(8769));
    layer2_outputs(1133) <= not(layer1_outputs(9730));
    layer2_outputs(1134) <= not(layer1_outputs(5840));
    layer2_outputs(1135) <= not(layer1_outputs(6081));
    layer2_outputs(1136) <= not(layer1_outputs(6597)) or (layer1_outputs(11132));
    layer2_outputs(1137) <= not((layer1_outputs(11878)) and (layer1_outputs(9897)));
    layer2_outputs(1138) <= (layer1_outputs(8120)) and (layer1_outputs(497));
    layer2_outputs(1139) <= layer1_outputs(9577);
    layer2_outputs(1140) <= not(layer1_outputs(12469));
    layer2_outputs(1141) <= not(layer1_outputs(7907)) or (layer1_outputs(10125));
    layer2_outputs(1142) <= not(layer1_outputs(11158));
    layer2_outputs(1143) <= (layer1_outputs(8349)) and not (layer1_outputs(1872));
    layer2_outputs(1144) <= (layer1_outputs(8722)) and not (layer1_outputs(3718));
    layer2_outputs(1145) <= not((layer1_outputs(6029)) and (layer1_outputs(4866)));
    layer2_outputs(1146) <= not((layer1_outputs(1295)) and (layer1_outputs(4365)));
    layer2_outputs(1147) <= not(layer1_outputs(11550)) or (layer1_outputs(9390));
    layer2_outputs(1148) <= not(layer1_outputs(489));
    layer2_outputs(1149) <= not(layer1_outputs(9676));
    layer2_outputs(1150) <= not((layer1_outputs(1647)) or (layer1_outputs(7324)));
    layer2_outputs(1151) <= not((layer1_outputs(4421)) xor (layer1_outputs(10906)));
    layer2_outputs(1152) <= not(layer1_outputs(5));
    layer2_outputs(1153) <= not(layer1_outputs(159)) or (layer1_outputs(8827));
    layer2_outputs(1154) <= not((layer1_outputs(10605)) xor (layer1_outputs(3472)));
    layer2_outputs(1155) <= (layer1_outputs(6119)) and not (layer1_outputs(671));
    layer2_outputs(1156) <= (layer1_outputs(11800)) or (layer1_outputs(1564));
    layer2_outputs(1157) <= not(layer1_outputs(8085));
    layer2_outputs(1158) <= (layer1_outputs(1515)) xor (layer1_outputs(2805));
    layer2_outputs(1159) <= not(layer1_outputs(5872));
    layer2_outputs(1160) <= not((layer1_outputs(10412)) and (layer1_outputs(10567)));
    layer2_outputs(1161) <= (layer1_outputs(4996)) or (layer1_outputs(6723));
    layer2_outputs(1162) <= not(layer1_outputs(5973));
    layer2_outputs(1163) <= (layer1_outputs(4834)) xor (layer1_outputs(4663));
    layer2_outputs(1164) <= layer1_outputs(11029);
    layer2_outputs(1165) <= (layer1_outputs(12398)) or (layer1_outputs(6995));
    layer2_outputs(1166) <= (layer1_outputs(7651)) and (layer1_outputs(4195));
    layer2_outputs(1167) <= layer1_outputs(2588);
    layer2_outputs(1168) <= layer1_outputs(10976);
    layer2_outputs(1169) <= (layer1_outputs(9507)) xor (layer1_outputs(3380));
    layer2_outputs(1170) <= not((layer1_outputs(7167)) or (layer1_outputs(8158)));
    layer2_outputs(1171) <= (layer1_outputs(12312)) xor (layer1_outputs(5353));
    layer2_outputs(1172) <= not(layer1_outputs(2657));
    layer2_outputs(1173) <= not((layer1_outputs(7642)) xor (layer1_outputs(11075)));
    layer2_outputs(1174) <= not(layer1_outputs(7545));
    layer2_outputs(1175) <= (layer1_outputs(7798)) xor (layer1_outputs(5088));
    layer2_outputs(1176) <= (layer1_outputs(8846)) xor (layer1_outputs(5199));
    layer2_outputs(1177) <= not((layer1_outputs(9234)) xor (layer1_outputs(8017)));
    layer2_outputs(1178) <= layer1_outputs(6773);
    layer2_outputs(1179) <= not(layer1_outputs(4755)) or (layer1_outputs(2340));
    layer2_outputs(1180) <= not(layer1_outputs(10631)) or (layer1_outputs(6215));
    layer2_outputs(1181) <= layer1_outputs(7835);
    layer2_outputs(1182) <= not(layer1_outputs(8952));
    layer2_outputs(1183) <= not((layer1_outputs(9674)) or (layer1_outputs(12250)));
    layer2_outputs(1184) <= not((layer1_outputs(6190)) or (layer1_outputs(918)));
    layer2_outputs(1185) <= not(layer1_outputs(6954));
    layer2_outputs(1186) <= not(layer1_outputs(8149));
    layer2_outputs(1187) <= layer1_outputs(10269);
    layer2_outputs(1188) <= (layer1_outputs(7801)) or (layer1_outputs(6990));
    layer2_outputs(1189) <= layer1_outputs(3745);
    layer2_outputs(1190) <= not((layer1_outputs(2454)) or (layer1_outputs(1531)));
    layer2_outputs(1191) <= not((layer1_outputs(1232)) or (layer1_outputs(10510)));
    layer2_outputs(1192) <= not(layer1_outputs(967));
    layer2_outputs(1193) <= not(layer1_outputs(1698));
    layer2_outputs(1194) <= not(layer1_outputs(1907));
    layer2_outputs(1195) <= not(layer1_outputs(12317));
    layer2_outputs(1196) <= layer1_outputs(11271);
    layer2_outputs(1197) <= not(layer1_outputs(2823));
    layer2_outputs(1198) <= (layer1_outputs(11388)) and not (layer1_outputs(2901));
    layer2_outputs(1199) <= (layer1_outputs(10345)) xor (layer1_outputs(6192));
    layer2_outputs(1200) <= (layer1_outputs(1544)) and not (layer1_outputs(8014));
    layer2_outputs(1201) <= (layer1_outputs(11035)) and not (layer1_outputs(1553));
    layer2_outputs(1202) <= (layer1_outputs(11897)) xor (layer1_outputs(2656));
    layer2_outputs(1203) <= (layer1_outputs(6634)) and (layer1_outputs(7621));
    layer2_outputs(1204) <= layer1_outputs(7499);
    layer2_outputs(1205) <= not(layer1_outputs(9734));
    layer2_outputs(1206) <= layer1_outputs(7654);
    layer2_outputs(1207) <= layer1_outputs(10177);
    layer2_outputs(1208) <= (layer1_outputs(1125)) and not (layer1_outputs(7111));
    layer2_outputs(1209) <= layer1_outputs(3463);
    layer2_outputs(1210) <= not(layer1_outputs(9964)) or (layer1_outputs(2073));
    layer2_outputs(1211) <= not((layer1_outputs(8926)) or (layer1_outputs(6675)));
    layer2_outputs(1212) <= not(layer1_outputs(7034)) or (layer1_outputs(9341));
    layer2_outputs(1213) <= not(layer1_outputs(10951));
    layer2_outputs(1214) <= (layer1_outputs(5969)) and not (layer1_outputs(8873));
    layer2_outputs(1215) <= (layer1_outputs(823)) xor (layer1_outputs(2534));
    layer2_outputs(1216) <= layer1_outputs(2934);
    layer2_outputs(1217) <= not(layer1_outputs(766));
    layer2_outputs(1218) <= layer1_outputs(2101);
    layer2_outputs(1219) <= not(layer1_outputs(9780)) or (layer1_outputs(4352));
    layer2_outputs(1220) <= not(layer1_outputs(10089));
    layer2_outputs(1221) <= layer1_outputs(10841);
    layer2_outputs(1222) <= (layer1_outputs(6831)) and not (layer1_outputs(4172));
    layer2_outputs(1223) <= not(layer1_outputs(8383));
    layer2_outputs(1224) <= layer1_outputs(3658);
    layer2_outputs(1225) <= not((layer1_outputs(3205)) and (layer1_outputs(12754)));
    layer2_outputs(1226) <= '0';
    layer2_outputs(1227) <= not(layer1_outputs(6988));
    layer2_outputs(1228) <= (layer1_outputs(8291)) and (layer1_outputs(281));
    layer2_outputs(1229) <= (layer1_outputs(2925)) or (layer1_outputs(11363));
    layer2_outputs(1230) <= (layer1_outputs(11533)) or (layer1_outputs(8372));
    layer2_outputs(1231) <= layer1_outputs(7127);
    layer2_outputs(1232) <= layer1_outputs(12285);
    layer2_outputs(1233) <= (layer1_outputs(81)) xor (layer1_outputs(12576));
    layer2_outputs(1234) <= (layer1_outputs(5059)) xor (layer1_outputs(8312));
    layer2_outputs(1235) <= layer1_outputs(10265);
    layer2_outputs(1236) <= not(layer1_outputs(2179)) or (layer1_outputs(7576));
    layer2_outputs(1237) <= layer1_outputs(5243);
    layer2_outputs(1238) <= layer1_outputs(7621);
    layer2_outputs(1239) <= (layer1_outputs(8652)) and (layer1_outputs(2836));
    layer2_outputs(1240) <= not(layer1_outputs(5255));
    layer2_outputs(1241) <= (layer1_outputs(27)) and not (layer1_outputs(10582));
    layer2_outputs(1242) <= (layer1_outputs(4256)) xor (layer1_outputs(3022));
    layer2_outputs(1243) <= not(layer1_outputs(10687));
    layer2_outputs(1244) <= (layer1_outputs(11985)) xor (layer1_outputs(9476));
    layer2_outputs(1245) <= not(layer1_outputs(395));
    layer2_outputs(1246) <= layer1_outputs(7168);
    layer2_outputs(1247) <= not((layer1_outputs(3013)) xor (layer1_outputs(8220)));
    layer2_outputs(1248) <= layer1_outputs(8777);
    layer2_outputs(1249) <= not((layer1_outputs(2819)) and (layer1_outputs(1815)));
    layer2_outputs(1250) <= not(layer1_outputs(1604));
    layer2_outputs(1251) <= not((layer1_outputs(6508)) or (layer1_outputs(7312)));
    layer2_outputs(1252) <= (layer1_outputs(11313)) xor (layer1_outputs(7678));
    layer2_outputs(1253) <= (layer1_outputs(12383)) and not (layer1_outputs(1065));
    layer2_outputs(1254) <= (layer1_outputs(10344)) xor (layer1_outputs(7693));
    layer2_outputs(1255) <= not(layer1_outputs(12043));
    layer2_outputs(1256) <= not((layer1_outputs(8278)) xor (layer1_outputs(3101)));
    layer2_outputs(1257) <= layer1_outputs(8259);
    layer2_outputs(1258) <= not(layer1_outputs(9096)) or (layer1_outputs(2430));
    layer2_outputs(1259) <= (layer1_outputs(8791)) and (layer1_outputs(11923));
    layer2_outputs(1260) <= layer1_outputs(940);
    layer2_outputs(1261) <= (layer1_outputs(8921)) and (layer1_outputs(1595));
    layer2_outputs(1262) <= (layer1_outputs(2375)) or (layer1_outputs(18));
    layer2_outputs(1263) <= not((layer1_outputs(6135)) or (layer1_outputs(11922)));
    layer2_outputs(1264) <= (layer1_outputs(2485)) xor (layer1_outputs(9200));
    layer2_outputs(1265) <= not(layer1_outputs(2279)) or (layer1_outputs(1006));
    layer2_outputs(1266) <= (layer1_outputs(2540)) and (layer1_outputs(4674));
    layer2_outputs(1267) <= (layer1_outputs(10008)) xor (layer1_outputs(10127));
    layer2_outputs(1268) <= layer1_outputs(3294);
    layer2_outputs(1269) <= '1';
    layer2_outputs(1270) <= not(layer1_outputs(9125)) or (layer1_outputs(11497));
    layer2_outputs(1271) <= not(layer1_outputs(6062));
    layer2_outputs(1272) <= not((layer1_outputs(6022)) and (layer1_outputs(12234)));
    layer2_outputs(1273) <= (layer1_outputs(5278)) and (layer1_outputs(4517));
    layer2_outputs(1274) <= layer1_outputs(5752);
    layer2_outputs(1275) <= (layer1_outputs(330)) and not (layer1_outputs(1986));
    layer2_outputs(1276) <= not((layer1_outputs(10364)) xor (layer1_outputs(1168)));
    layer2_outputs(1277) <= not(layer1_outputs(5847)) or (layer1_outputs(9141));
    layer2_outputs(1278) <= layer1_outputs(7608);
    layer2_outputs(1279) <= layer1_outputs(1159);
    layer2_outputs(1280) <= not(layer1_outputs(5167)) or (layer1_outputs(10114));
    layer2_outputs(1281) <= not(layer1_outputs(11326));
    layer2_outputs(1282) <= layer1_outputs(8233);
    layer2_outputs(1283) <= not(layer1_outputs(7220));
    layer2_outputs(1284) <= not(layer1_outputs(9791));
    layer2_outputs(1285) <= (layer1_outputs(10459)) and (layer1_outputs(12266));
    layer2_outputs(1286) <= (layer1_outputs(9944)) and not (layer1_outputs(3070));
    layer2_outputs(1287) <= (layer1_outputs(11290)) or (layer1_outputs(12758));
    layer2_outputs(1288) <= layer1_outputs(12068);
    layer2_outputs(1289) <= not((layer1_outputs(12210)) or (layer1_outputs(10088)));
    layer2_outputs(1290) <= (layer1_outputs(3946)) and (layer1_outputs(6889));
    layer2_outputs(1291) <= not(layer1_outputs(6749));
    layer2_outputs(1292) <= not((layer1_outputs(3779)) xor (layer1_outputs(3377)));
    layer2_outputs(1293) <= not((layer1_outputs(7957)) or (layer1_outputs(584)));
    layer2_outputs(1294) <= layer1_outputs(826);
    layer2_outputs(1295) <= layer1_outputs(5111);
    layer2_outputs(1296) <= not(layer1_outputs(7349));
    layer2_outputs(1297) <= not(layer1_outputs(3151)) or (layer1_outputs(10460));
    layer2_outputs(1298) <= layer1_outputs(3545);
    layer2_outputs(1299) <= not(layer1_outputs(10484));
    layer2_outputs(1300) <= (layer1_outputs(2800)) xor (layer1_outputs(2704));
    layer2_outputs(1301) <= layer1_outputs(8834);
    layer2_outputs(1302) <= (layer1_outputs(11508)) and not (layer1_outputs(4655));
    layer2_outputs(1303) <= not(layer1_outputs(5549));
    layer2_outputs(1304) <= (layer1_outputs(2818)) xor (layer1_outputs(4640));
    layer2_outputs(1305) <= not((layer1_outputs(2749)) and (layer1_outputs(9630)));
    layer2_outputs(1306) <= layer1_outputs(4369);
    layer2_outputs(1307) <= (layer1_outputs(4316)) xor (layer1_outputs(10246));
    layer2_outputs(1308) <= not(layer1_outputs(3079));
    layer2_outputs(1309) <= layer1_outputs(10830);
    layer2_outputs(1310) <= not((layer1_outputs(6232)) and (layer1_outputs(3752)));
    layer2_outputs(1311) <= not(layer1_outputs(5891));
    layer2_outputs(1312) <= not(layer1_outputs(10678));
    layer2_outputs(1313) <= layer1_outputs(5627);
    layer2_outputs(1314) <= layer1_outputs(3676);
    layer2_outputs(1315) <= layer1_outputs(10148);
    layer2_outputs(1316) <= not(layer1_outputs(9384));
    layer2_outputs(1317) <= not(layer1_outputs(8854));
    layer2_outputs(1318) <= layer1_outputs(4485);
    layer2_outputs(1319) <= not(layer1_outputs(9868)) or (layer1_outputs(5381));
    layer2_outputs(1320) <= not(layer1_outputs(3166));
    layer2_outputs(1321) <= not(layer1_outputs(8476)) or (layer1_outputs(8734));
    layer2_outputs(1322) <= (layer1_outputs(8656)) and (layer1_outputs(724));
    layer2_outputs(1323) <= layer1_outputs(5045);
    layer2_outputs(1324) <= not(layer1_outputs(3697));
    layer2_outputs(1325) <= not(layer1_outputs(2027)) or (layer1_outputs(10848));
    layer2_outputs(1326) <= not(layer1_outputs(7707)) or (layer1_outputs(1515));
    layer2_outputs(1327) <= not(layer1_outputs(10663));
    layer2_outputs(1328) <= layer1_outputs(2394);
    layer2_outputs(1329) <= layer1_outputs(4490);
    layer2_outputs(1330) <= (layer1_outputs(9585)) and not (layer1_outputs(1214));
    layer2_outputs(1331) <= not((layer1_outputs(5798)) or (layer1_outputs(9955)));
    layer2_outputs(1332) <= not(layer1_outputs(8003)) or (layer1_outputs(21));
    layer2_outputs(1333) <= (layer1_outputs(5753)) xor (layer1_outputs(9493));
    layer2_outputs(1334) <= (layer1_outputs(5125)) and not (layer1_outputs(10619));
    layer2_outputs(1335) <= not(layer1_outputs(9501));
    layer2_outputs(1336) <= layer1_outputs(4536);
    layer2_outputs(1337) <= layer1_outputs(11085);
    layer2_outputs(1338) <= not((layer1_outputs(6540)) or (layer1_outputs(1620)));
    layer2_outputs(1339) <= not(layer1_outputs(1082));
    layer2_outputs(1340) <= (layer1_outputs(6274)) xor (layer1_outputs(8157));
    layer2_outputs(1341) <= layer1_outputs(2974);
    layer2_outputs(1342) <= (layer1_outputs(9782)) and (layer1_outputs(5839));
    layer2_outputs(1343) <= '0';
    layer2_outputs(1344) <= not((layer1_outputs(3780)) or (layer1_outputs(12020)));
    layer2_outputs(1345) <= not((layer1_outputs(1248)) or (layer1_outputs(10102)));
    layer2_outputs(1346) <= layer1_outputs(3003);
    layer2_outputs(1347) <= not(layer1_outputs(9738)) or (layer1_outputs(8806));
    layer2_outputs(1348) <= '1';
    layer2_outputs(1349) <= layer1_outputs(9042);
    layer2_outputs(1350) <= not(layer1_outputs(10802)) or (layer1_outputs(11262));
    layer2_outputs(1351) <= layer1_outputs(10894);
    layer2_outputs(1352) <= (layer1_outputs(7971)) xor (layer1_outputs(8603));
    layer2_outputs(1353) <= layer1_outputs(9651);
    layer2_outputs(1354) <= not(layer1_outputs(3234));
    layer2_outputs(1355) <= layer1_outputs(1992);
    layer2_outputs(1356) <= '1';
    layer2_outputs(1357) <= (layer1_outputs(5514)) or (layer1_outputs(12062));
    layer2_outputs(1358) <= not(layer1_outputs(12252));
    layer2_outputs(1359) <= not(layer1_outputs(7773));
    layer2_outputs(1360) <= not(layer1_outputs(11764));
    layer2_outputs(1361) <= not((layer1_outputs(6205)) xor (layer1_outputs(4430)));
    layer2_outputs(1362) <= layer1_outputs(1067);
    layer2_outputs(1363) <= (layer1_outputs(571)) and not (layer1_outputs(2744));
    layer2_outputs(1364) <= not(layer1_outputs(11853)) or (layer1_outputs(8425));
    layer2_outputs(1365) <= (layer1_outputs(12703)) and not (layer1_outputs(10138));
    layer2_outputs(1366) <= (layer1_outputs(10950)) or (layer1_outputs(8136));
    layer2_outputs(1367) <= layer1_outputs(3861);
    layer2_outputs(1368) <= not((layer1_outputs(1346)) xor (layer1_outputs(496)));
    layer2_outputs(1369) <= layer1_outputs(1978);
    layer2_outputs(1370) <= not(layer1_outputs(11905));
    layer2_outputs(1371) <= not((layer1_outputs(12492)) xor (layer1_outputs(2058)));
    layer2_outputs(1372) <= not((layer1_outputs(1572)) xor (layer1_outputs(9995)));
    layer2_outputs(1373) <= (layer1_outputs(4039)) and not (layer1_outputs(2468));
    layer2_outputs(1374) <= not((layer1_outputs(639)) or (layer1_outputs(1570)));
    layer2_outputs(1375) <= not(layer1_outputs(8642));
    layer2_outputs(1376) <= not(layer1_outputs(6332)) or (layer1_outputs(8679));
    layer2_outputs(1377) <= not((layer1_outputs(3605)) or (layer1_outputs(6969)));
    layer2_outputs(1378) <= not((layer1_outputs(5782)) xor (layer1_outputs(100)));
    layer2_outputs(1379) <= not(layer1_outputs(1502));
    layer2_outputs(1380) <= layer1_outputs(3525);
    layer2_outputs(1381) <= not((layer1_outputs(8520)) xor (layer1_outputs(3865)));
    layer2_outputs(1382) <= (layer1_outputs(4600)) xor (layer1_outputs(1459));
    layer2_outputs(1383) <= not(layer1_outputs(11974));
    layer2_outputs(1384) <= (layer1_outputs(2987)) xor (layer1_outputs(8465));
    layer2_outputs(1385) <= not(layer1_outputs(4049));
    layer2_outputs(1386) <= (layer1_outputs(9510)) and (layer1_outputs(3372));
    layer2_outputs(1387) <= not(layer1_outputs(7133)) or (layer1_outputs(1793));
    layer2_outputs(1388) <= (layer1_outputs(9975)) or (layer1_outputs(9692));
    layer2_outputs(1389) <= layer1_outputs(11605);
    layer2_outputs(1390) <= not((layer1_outputs(784)) xor (layer1_outputs(7643)));
    layer2_outputs(1391) <= layer1_outputs(6756);
    layer2_outputs(1392) <= not((layer1_outputs(7017)) and (layer1_outputs(11268)));
    layer2_outputs(1393) <= (layer1_outputs(7018)) and (layer1_outputs(5203));
    layer2_outputs(1394) <= not((layer1_outputs(6719)) and (layer1_outputs(1184)));
    layer2_outputs(1395) <= (layer1_outputs(8621)) or (layer1_outputs(10845));
    layer2_outputs(1396) <= not((layer1_outputs(3947)) and (layer1_outputs(1517)));
    layer2_outputs(1397) <= (layer1_outputs(595)) and (layer1_outputs(938));
    layer2_outputs(1398) <= not((layer1_outputs(9185)) xor (layer1_outputs(3484)));
    layer2_outputs(1399) <= layer1_outputs(10063);
    layer2_outputs(1400) <= layer1_outputs(2185);
    layer2_outputs(1401) <= not(layer1_outputs(11756));
    layer2_outputs(1402) <= layer1_outputs(11067);
    layer2_outputs(1403) <= (layer1_outputs(5769)) or (layer1_outputs(9733));
    layer2_outputs(1404) <= not(layer1_outputs(5228));
    layer2_outputs(1405) <= (layer1_outputs(7194)) or (layer1_outputs(5013));
    layer2_outputs(1406) <= not(layer1_outputs(6651)) or (layer1_outputs(7121));
    layer2_outputs(1407) <= (layer1_outputs(9860)) xor (layer1_outputs(1382));
    layer2_outputs(1408) <= not(layer1_outputs(12430));
    layer2_outputs(1409) <= (layer1_outputs(11115)) xor (layer1_outputs(11820));
    layer2_outputs(1410) <= (layer1_outputs(6906)) or (layer1_outputs(4527));
    layer2_outputs(1411) <= (layer1_outputs(9383)) xor (layer1_outputs(5664));
    layer2_outputs(1412) <= (layer1_outputs(10519)) and not (layer1_outputs(7866));
    layer2_outputs(1413) <= not(layer1_outputs(4777));
    layer2_outputs(1414) <= not((layer1_outputs(8435)) xor (layer1_outputs(6072)));
    layer2_outputs(1415) <= (layer1_outputs(724)) and not (layer1_outputs(9879));
    layer2_outputs(1416) <= layer1_outputs(2761);
    layer2_outputs(1417) <= not(layer1_outputs(1841));
    layer2_outputs(1418) <= not(layer1_outputs(11770));
    layer2_outputs(1419) <= not((layer1_outputs(6060)) xor (layer1_outputs(3842)));
    layer2_outputs(1420) <= not(layer1_outputs(2012)) or (layer1_outputs(6524));
    layer2_outputs(1421) <= not(layer1_outputs(4126));
    layer2_outputs(1422) <= not(layer1_outputs(1858));
    layer2_outputs(1423) <= (layer1_outputs(8768)) and not (layer1_outputs(10394));
    layer2_outputs(1424) <= not(layer1_outputs(273));
    layer2_outputs(1425) <= (layer1_outputs(7744)) and not (layer1_outputs(7174));
    layer2_outputs(1426) <= not((layer1_outputs(8625)) or (layer1_outputs(6194)));
    layer2_outputs(1427) <= (layer1_outputs(12154)) and not (layer1_outputs(8744));
    layer2_outputs(1428) <= not((layer1_outputs(7023)) and (layer1_outputs(5617)));
    layer2_outputs(1429) <= (layer1_outputs(2096)) or (layer1_outputs(1639));
    layer2_outputs(1430) <= (layer1_outputs(6701)) and not (layer1_outputs(3347));
    layer2_outputs(1431) <= (layer1_outputs(7665)) xor (layer1_outputs(5501));
    layer2_outputs(1432) <= layer1_outputs(5908);
    layer2_outputs(1433) <= layer1_outputs(8464);
    layer2_outputs(1434) <= layer1_outputs(4638);
    layer2_outputs(1435) <= layer1_outputs(10194);
    layer2_outputs(1436) <= not(layer1_outputs(1032));
    layer2_outputs(1437) <= not((layer1_outputs(4228)) xor (layer1_outputs(11016)));
    layer2_outputs(1438) <= layer1_outputs(11338);
    layer2_outputs(1439) <= (layer1_outputs(7327)) and (layer1_outputs(102));
    layer2_outputs(1440) <= not(layer1_outputs(4287));
    layer2_outputs(1441) <= (layer1_outputs(2779)) and not (layer1_outputs(11958));
    layer2_outputs(1442) <= not(layer1_outputs(8836));
    layer2_outputs(1443) <= layer1_outputs(12417);
    layer2_outputs(1444) <= not(layer1_outputs(1794));
    layer2_outputs(1445) <= not(layer1_outputs(9835));
    layer2_outputs(1446) <= (layer1_outputs(10285)) xor (layer1_outputs(11999));
    layer2_outputs(1447) <= layer1_outputs(5625);
    layer2_outputs(1448) <= (layer1_outputs(3992)) or (layer1_outputs(441));
    layer2_outputs(1449) <= not((layer1_outputs(4026)) and (layer1_outputs(11138)));
    layer2_outputs(1450) <= (layer1_outputs(3111)) xor (layer1_outputs(10069));
    layer2_outputs(1451) <= layer1_outputs(3891);
    layer2_outputs(1452) <= not(layer1_outputs(4125));
    layer2_outputs(1453) <= (layer1_outputs(64)) and not (layer1_outputs(7083));
    layer2_outputs(1454) <= not(layer1_outputs(6116)) or (layer1_outputs(6920));
    layer2_outputs(1455) <= layer1_outputs(8338);
    layer2_outputs(1456) <= layer1_outputs(253);
    layer2_outputs(1457) <= not(layer1_outputs(3097));
    layer2_outputs(1458) <= not(layer1_outputs(125));
    layer2_outputs(1459) <= (layer1_outputs(1137)) or (layer1_outputs(956));
    layer2_outputs(1460) <= not(layer1_outputs(2416));
    layer2_outputs(1461) <= not((layer1_outputs(9611)) and (layer1_outputs(345)));
    layer2_outputs(1462) <= not((layer1_outputs(9954)) xor (layer1_outputs(3031)));
    layer2_outputs(1463) <= not((layer1_outputs(8558)) and (layer1_outputs(6222)));
    layer2_outputs(1464) <= (layer1_outputs(85)) and (layer1_outputs(6888));
    layer2_outputs(1465) <= (layer1_outputs(8339)) and not (layer1_outputs(12675));
    layer2_outputs(1466) <= (layer1_outputs(4073)) and not (layer1_outputs(5340));
    layer2_outputs(1467) <= not((layer1_outputs(142)) xor (layer1_outputs(11440)));
    layer2_outputs(1468) <= layer1_outputs(5476);
    layer2_outputs(1469) <= not((layer1_outputs(4211)) or (layer1_outputs(3144)));
    layer2_outputs(1470) <= not(layer1_outputs(9298));
    layer2_outputs(1471) <= not((layer1_outputs(3731)) xor (layer1_outputs(1094)));
    layer2_outputs(1472) <= (layer1_outputs(8539)) or (layer1_outputs(12327));
    layer2_outputs(1473) <= (layer1_outputs(10811)) and not (layer1_outputs(5150));
    layer2_outputs(1474) <= layer1_outputs(8945);
    layer2_outputs(1475) <= not(layer1_outputs(11112));
    layer2_outputs(1476) <= not(layer1_outputs(835)) or (layer1_outputs(40));
    layer2_outputs(1477) <= layer1_outputs(524);
    layer2_outputs(1478) <= (layer1_outputs(12477)) and not (layer1_outputs(9508));
    layer2_outputs(1479) <= (layer1_outputs(2742)) and not (layer1_outputs(5207));
    layer2_outputs(1480) <= not(layer1_outputs(2395));
    layer2_outputs(1481) <= (layer1_outputs(8383)) and (layer1_outputs(12544));
    layer2_outputs(1482) <= layer1_outputs(3652);
    layer2_outputs(1483) <= layer1_outputs(10410);
    layer2_outputs(1484) <= layer1_outputs(5493);
    layer2_outputs(1485) <= (layer1_outputs(3103)) xor (layer1_outputs(7234));
    layer2_outputs(1486) <= (layer1_outputs(10635)) and (layer1_outputs(2225));
    layer2_outputs(1487) <= (layer1_outputs(11805)) and (layer1_outputs(10273));
    layer2_outputs(1488) <= not(layer1_outputs(3302));
    layer2_outputs(1489) <= layer1_outputs(10153);
    layer2_outputs(1490) <= (layer1_outputs(3886)) and not (layer1_outputs(6038));
    layer2_outputs(1491) <= (layer1_outputs(12696)) and not (layer1_outputs(7268));
    layer2_outputs(1492) <= not((layer1_outputs(4480)) xor (layer1_outputs(7422)));
    layer2_outputs(1493) <= not((layer1_outputs(11495)) xor (layer1_outputs(7320)));
    layer2_outputs(1494) <= (layer1_outputs(8273)) or (layer1_outputs(6567));
    layer2_outputs(1495) <= layer1_outputs(289);
    layer2_outputs(1496) <= '0';
    layer2_outputs(1497) <= not((layer1_outputs(6608)) and (layer1_outputs(8355)));
    layer2_outputs(1498) <= not((layer1_outputs(4369)) or (layer1_outputs(8238)));
    layer2_outputs(1499) <= not((layer1_outputs(11839)) xor (layer1_outputs(1195)));
    layer2_outputs(1500) <= layer1_outputs(6740);
    layer2_outputs(1501) <= (layer1_outputs(9788)) xor (layer1_outputs(5046));
    layer2_outputs(1502) <= (layer1_outputs(3439)) and not (layer1_outputs(9494));
    layer2_outputs(1503) <= (layer1_outputs(5690)) and not (layer1_outputs(2907));
    layer2_outputs(1504) <= (layer1_outputs(12506)) and not (layer1_outputs(3668));
    layer2_outputs(1505) <= (layer1_outputs(9312)) xor (layer1_outputs(10222));
    layer2_outputs(1506) <= not((layer1_outputs(9720)) xor (layer1_outputs(9813)));
    layer2_outputs(1507) <= layer1_outputs(11358);
    layer2_outputs(1508) <= not(layer1_outputs(2477));
    layer2_outputs(1509) <= not(layer1_outputs(4006));
    layer2_outputs(1510) <= not(layer1_outputs(605)) or (layer1_outputs(645));
    layer2_outputs(1511) <= not((layer1_outputs(1691)) or (layer1_outputs(4997)));
    layer2_outputs(1512) <= not(layer1_outputs(12018));
    layer2_outputs(1513) <= (layer1_outputs(5432)) and not (layer1_outputs(1518));
    layer2_outputs(1514) <= layer1_outputs(10415);
    layer2_outputs(1515) <= not((layer1_outputs(6564)) xor (layer1_outputs(5195)));
    layer2_outputs(1516) <= not(layer1_outputs(6403));
    layer2_outputs(1517) <= layer1_outputs(4926);
    layer2_outputs(1518) <= not(layer1_outputs(301));
    layer2_outputs(1519) <= (layer1_outputs(6197)) and not (layer1_outputs(9336));
    layer2_outputs(1520) <= (layer1_outputs(3099)) xor (layer1_outputs(12044));
    layer2_outputs(1521) <= not(layer1_outputs(3837));
    layer2_outputs(1522) <= not(layer1_outputs(5363));
    layer2_outputs(1523) <= layer1_outputs(3522);
    layer2_outputs(1524) <= not(layer1_outputs(3422));
    layer2_outputs(1525) <= (layer1_outputs(1209)) and not (layer1_outputs(11720));
    layer2_outputs(1526) <= (layer1_outputs(11772)) and (layer1_outputs(4098));
    layer2_outputs(1527) <= not(layer1_outputs(7897));
    layer2_outputs(1528) <= not(layer1_outputs(7992)) or (layer1_outputs(5260));
    layer2_outputs(1529) <= (layer1_outputs(11589)) xor (layer1_outputs(8666));
    layer2_outputs(1530) <= not(layer1_outputs(10681));
    layer2_outputs(1531) <= not(layer1_outputs(969)) or (layer1_outputs(9149));
    layer2_outputs(1532) <= (layer1_outputs(8479)) xor (layer1_outputs(2386));
    layer2_outputs(1533) <= (layer1_outputs(12171)) xor (layer1_outputs(11225));
    layer2_outputs(1534) <= layer1_outputs(3671);
    layer2_outputs(1535) <= not(layer1_outputs(2678)) or (layer1_outputs(1699));
    layer2_outputs(1536) <= (layer1_outputs(2280)) or (layer1_outputs(7233));
    layer2_outputs(1537) <= not(layer1_outputs(10871));
    layer2_outputs(1538) <= not((layer1_outputs(887)) xor (layer1_outputs(4738)));
    layer2_outputs(1539) <= not(layer1_outputs(7212));
    layer2_outputs(1540) <= not(layer1_outputs(1103));
    layer2_outputs(1541) <= not(layer1_outputs(5022)) or (layer1_outputs(7536));
    layer2_outputs(1542) <= not((layer1_outputs(6015)) xor (layer1_outputs(12294)));
    layer2_outputs(1543) <= layer1_outputs(2924);
    layer2_outputs(1544) <= layer1_outputs(7458);
    layer2_outputs(1545) <= (layer1_outputs(1519)) or (layer1_outputs(9809));
    layer2_outputs(1546) <= not(layer1_outputs(9044));
    layer2_outputs(1547) <= (layer1_outputs(12136)) xor (layer1_outputs(12216));
    layer2_outputs(1548) <= not(layer1_outputs(4455));
    layer2_outputs(1549) <= not(layer1_outputs(9788));
    layer2_outputs(1550) <= (layer1_outputs(6490)) xor (layer1_outputs(8226));
    layer2_outputs(1551) <= not((layer1_outputs(10103)) xor (layer1_outputs(7536)));
    layer2_outputs(1552) <= layer1_outputs(7153);
    layer2_outputs(1553) <= not(layer1_outputs(11460)) or (layer1_outputs(11153));
    layer2_outputs(1554) <= layer1_outputs(9909);
    layer2_outputs(1555) <= layer1_outputs(1467);
    layer2_outputs(1556) <= (layer1_outputs(2387)) or (layer1_outputs(6995));
    layer2_outputs(1557) <= not(layer1_outputs(8460)) or (layer1_outputs(10518));
    layer2_outputs(1558) <= (layer1_outputs(12783)) and not (layer1_outputs(10653));
    layer2_outputs(1559) <= layer1_outputs(2157);
    layer2_outputs(1560) <= layer1_outputs(5715);
    layer2_outputs(1561) <= not(layer1_outputs(9017));
    layer2_outputs(1562) <= not(layer1_outputs(3572)) or (layer1_outputs(6006));
    layer2_outputs(1563) <= not((layer1_outputs(1221)) xor (layer1_outputs(9927)));
    layer2_outputs(1564) <= layer1_outputs(5506);
    layer2_outputs(1565) <= (layer1_outputs(3711)) and not (layer1_outputs(1097));
    layer2_outputs(1566) <= (layer1_outputs(3)) or (layer1_outputs(9219));
    layer2_outputs(1567) <= layer1_outputs(7902);
    layer2_outputs(1568) <= not(layer1_outputs(8237)) or (layer1_outputs(8143));
    layer2_outputs(1569) <= not(layer1_outputs(2255));
    layer2_outputs(1570) <= not(layer1_outputs(2637));
    layer2_outputs(1571) <= not((layer1_outputs(842)) and (layer1_outputs(1575)));
    layer2_outputs(1572) <= layer1_outputs(5544);
    layer2_outputs(1573) <= not(layer1_outputs(11458));
    layer2_outputs(1574) <= not((layer1_outputs(5700)) or (layer1_outputs(7803)));
    layer2_outputs(1575) <= (layer1_outputs(3973)) xor (layer1_outputs(3557));
    layer2_outputs(1576) <= not(layer1_outputs(4620));
    layer2_outputs(1577) <= (layer1_outputs(2437)) or (layer1_outputs(5182));
    layer2_outputs(1578) <= layer1_outputs(8791);
    layer2_outputs(1579) <= not((layer1_outputs(12651)) xor (layer1_outputs(521)));
    layer2_outputs(1580) <= not(layer1_outputs(630));
    layer2_outputs(1581) <= layer1_outputs(4255);
    layer2_outputs(1582) <= layer1_outputs(909);
    layer2_outputs(1583) <= layer1_outputs(10828);
    layer2_outputs(1584) <= layer1_outputs(1311);
    layer2_outputs(1585) <= not(layer1_outputs(2152)) or (layer1_outputs(1261));
    layer2_outputs(1586) <= (layer1_outputs(11306)) xor (layer1_outputs(1173));
    layer2_outputs(1587) <= not(layer1_outputs(10728)) or (layer1_outputs(4031));
    layer2_outputs(1588) <= (layer1_outputs(5274)) or (layer1_outputs(2233));
    layer2_outputs(1589) <= not(layer1_outputs(4675)) or (layer1_outputs(6076));
    layer2_outputs(1590) <= not((layer1_outputs(3624)) xor (layer1_outputs(3588)));
    layer2_outputs(1591) <= layer1_outputs(7269);
    layer2_outputs(1592) <= layer1_outputs(2840);
    layer2_outputs(1593) <= layer1_outputs(1665);
    layer2_outputs(1594) <= (layer1_outputs(7235)) and not (layer1_outputs(4355));
    layer2_outputs(1595) <= layer1_outputs(4681);
    layer2_outputs(1596) <= (layer1_outputs(10280)) xor (layer1_outputs(96));
    layer2_outputs(1597) <= layer1_outputs(1549);
    layer2_outputs(1598) <= not(layer1_outputs(6162));
    layer2_outputs(1599) <= not(layer1_outputs(4617));
    layer2_outputs(1600) <= not(layer1_outputs(10652)) or (layer1_outputs(10948));
    layer2_outputs(1601) <= (layer1_outputs(7961)) and not (layer1_outputs(4146));
    layer2_outputs(1602) <= not(layer1_outputs(3084));
    layer2_outputs(1603) <= not(layer1_outputs(5707));
    layer2_outputs(1604) <= not((layer1_outputs(2943)) xor (layer1_outputs(4475)));
    layer2_outputs(1605) <= not(layer1_outputs(4220));
    layer2_outputs(1606) <= (layer1_outputs(8312)) and not (layer1_outputs(4983));
    layer2_outputs(1607) <= layer1_outputs(12377);
    layer2_outputs(1608) <= not(layer1_outputs(4037));
    layer2_outputs(1609) <= (layer1_outputs(2083)) xor (layer1_outputs(8597));
    layer2_outputs(1610) <= (layer1_outputs(2603)) and (layer1_outputs(3255));
    layer2_outputs(1611) <= not((layer1_outputs(12119)) or (layer1_outputs(8946)));
    layer2_outputs(1612) <= (layer1_outputs(9869)) or (layer1_outputs(7176));
    layer2_outputs(1613) <= not(layer1_outputs(2721));
    layer2_outputs(1614) <= layer1_outputs(4184);
    layer2_outputs(1615) <= (layer1_outputs(5259)) xor (layer1_outputs(6430));
    layer2_outputs(1616) <= not(layer1_outputs(7434));
    layer2_outputs(1617) <= layer1_outputs(3742);
    layer2_outputs(1618) <= not(layer1_outputs(8717));
    layer2_outputs(1619) <= layer1_outputs(5187);
    layer2_outputs(1620) <= (layer1_outputs(1074)) and not (layer1_outputs(4904));
    layer2_outputs(1621) <= (layer1_outputs(11686)) or (layer1_outputs(5135));
    layer2_outputs(1622) <= not(layer1_outputs(11319)) or (layer1_outputs(6276));
    layer2_outputs(1623) <= layer1_outputs(3417);
    layer2_outputs(1624) <= layer1_outputs(10942);
    layer2_outputs(1625) <= not((layer1_outputs(2035)) and (layer1_outputs(4317)));
    layer2_outputs(1626) <= (layer1_outputs(8315)) and not (layer1_outputs(9549));
    layer2_outputs(1627) <= not(layer1_outputs(9148));
    layer2_outputs(1628) <= layer1_outputs(12338);
    layer2_outputs(1629) <= not(layer1_outputs(2856)) or (layer1_outputs(12010));
    layer2_outputs(1630) <= not(layer1_outputs(5003));
    layer2_outputs(1631) <= not(layer1_outputs(3478));
    layer2_outputs(1632) <= layer1_outputs(1119);
    layer2_outputs(1633) <= not(layer1_outputs(270));
    layer2_outputs(1634) <= not((layer1_outputs(3968)) xor (layer1_outputs(11721)));
    layer2_outputs(1635) <= not(layer1_outputs(7474));
    layer2_outputs(1636) <= not(layer1_outputs(768));
    layer2_outputs(1637) <= not(layer1_outputs(5105));
    layer2_outputs(1638) <= layer1_outputs(4574);
    layer2_outputs(1639) <= not((layer1_outputs(9451)) or (layer1_outputs(11595)));
    layer2_outputs(1640) <= layer1_outputs(12222);
    layer2_outputs(1641) <= layer1_outputs(1120);
    layer2_outputs(1642) <= (layer1_outputs(11378)) xor (layer1_outputs(7169));
    layer2_outputs(1643) <= (layer1_outputs(5408)) and not (layer1_outputs(5461));
    layer2_outputs(1644) <= layer1_outputs(747);
    layer2_outputs(1645) <= (layer1_outputs(9314)) and not (layer1_outputs(6365));
    layer2_outputs(1646) <= '1';
    layer2_outputs(1647) <= (layer1_outputs(5907)) and not (layer1_outputs(297));
    layer2_outputs(1648) <= layer1_outputs(6196);
    layer2_outputs(1649) <= not(layer1_outputs(132));
    layer2_outputs(1650) <= layer1_outputs(803);
    layer2_outputs(1651) <= not((layer1_outputs(6330)) and (layer1_outputs(697)));
    layer2_outputs(1652) <= layer1_outputs(9353);
    layer2_outputs(1653) <= not(layer1_outputs(3193));
    layer2_outputs(1654) <= not(layer1_outputs(2845));
    layer2_outputs(1655) <= layer1_outputs(4417);
    layer2_outputs(1656) <= (layer1_outputs(1536)) and not (layer1_outputs(6589));
    layer2_outputs(1657) <= not((layer1_outputs(3930)) xor (layer1_outputs(115)));
    layer2_outputs(1658) <= (layer1_outputs(8667)) and (layer1_outputs(5889));
    layer2_outputs(1659) <= not(layer1_outputs(12307));
    layer2_outputs(1660) <= not(layer1_outputs(7100));
    layer2_outputs(1661) <= layer1_outputs(2695);
    layer2_outputs(1662) <= not((layer1_outputs(7144)) or (layer1_outputs(5944)));
    layer2_outputs(1663) <= (layer1_outputs(8426)) or (layer1_outputs(2615));
    layer2_outputs(1664) <= (layer1_outputs(12672)) xor (layer1_outputs(9130));
    layer2_outputs(1665) <= layer1_outputs(2516);
    layer2_outputs(1666) <= not(layer1_outputs(11089)) or (layer1_outputs(5444));
    layer2_outputs(1667) <= not(layer1_outputs(11521)) or (layer1_outputs(10478));
    layer2_outputs(1668) <= layer1_outputs(9617);
    layer2_outputs(1669) <= (layer1_outputs(12517)) or (layer1_outputs(5983));
    layer2_outputs(1670) <= layer1_outputs(11562);
    layer2_outputs(1671) <= layer1_outputs(4565);
    layer2_outputs(1672) <= not(layer1_outputs(10547));
    layer2_outputs(1673) <= layer1_outputs(8993);
    layer2_outputs(1674) <= (layer1_outputs(7347)) xor (layer1_outputs(8876));
    layer2_outputs(1675) <= (layer1_outputs(3681)) or (layer1_outputs(8480));
    layer2_outputs(1676) <= (layer1_outputs(9121)) or (layer1_outputs(11825));
    layer2_outputs(1677) <= (layer1_outputs(5575)) or (layer1_outputs(11263));
    layer2_outputs(1678) <= (layer1_outputs(12139)) or (layer1_outputs(1903));
    layer2_outputs(1679) <= not(layer1_outputs(159));
    layer2_outputs(1680) <= layer1_outputs(8069);
    layer2_outputs(1681) <= layer1_outputs(12305);
    layer2_outputs(1682) <= layer1_outputs(10505);
    layer2_outputs(1683) <= not((layer1_outputs(6589)) xor (layer1_outputs(8928)));
    layer2_outputs(1684) <= not(layer1_outputs(9935));
    layer2_outputs(1685) <= not((layer1_outputs(3536)) xor (layer1_outputs(10530)));
    layer2_outputs(1686) <= not((layer1_outputs(3578)) or (layer1_outputs(119)));
    layer2_outputs(1687) <= not((layer1_outputs(12225)) xor (layer1_outputs(4392)));
    layer2_outputs(1688) <= layer1_outputs(1899);
    layer2_outputs(1689) <= (layer1_outputs(6884)) xor (layer1_outputs(12315));
    layer2_outputs(1690) <= layer1_outputs(7820);
    layer2_outputs(1691) <= layer1_outputs(6220);
    layer2_outputs(1692) <= not(layer1_outputs(11147));
    layer2_outputs(1693) <= '0';
    layer2_outputs(1694) <= (layer1_outputs(4387)) and (layer1_outputs(4377));
    layer2_outputs(1695) <= not(layer1_outputs(6161));
    layer2_outputs(1696) <= (layer1_outputs(11033)) xor (layer1_outputs(671));
    layer2_outputs(1697) <= not(layer1_outputs(12269));
    layer2_outputs(1698) <= (layer1_outputs(49)) and not (layer1_outputs(6708));
    layer2_outputs(1699) <= layer1_outputs(5533);
    layer2_outputs(1700) <= not((layer1_outputs(116)) and (layer1_outputs(3709)));
    layer2_outputs(1701) <= not((layer1_outputs(3590)) or (layer1_outputs(33)));
    layer2_outputs(1702) <= not(layer1_outputs(2899));
    layer2_outputs(1703) <= (layer1_outputs(12411)) and not (layer1_outputs(8659));
    layer2_outputs(1704) <= layer1_outputs(323);
    layer2_outputs(1705) <= not((layer1_outputs(2880)) or (layer1_outputs(9195)));
    layer2_outputs(1706) <= (layer1_outputs(12481)) xor (layer1_outputs(4360));
    layer2_outputs(1707) <= layer1_outputs(2514);
    layer2_outputs(1708) <= (layer1_outputs(9262)) xor (layer1_outputs(11173));
    layer2_outputs(1709) <= not((layer1_outputs(5552)) xor (layer1_outputs(7726)));
    layer2_outputs(1710) <= not(layer1_outputs(11725)) or (layer1_outputs(571));
    layer2_outputs(1711) <= not(layer1_outputs(11185));
    layer2_outputs(1712) <= layer1_outputs(9906);
    layer2_outputs(1713) <= layer1_outputs(10242);
    layer2_outputs(1714) <= (layer1_outputs(4999)) and not (layer1_outputs(5466));
    layer2_outputs(1715) <= not(layer1_outputs(4979)) or (layer1_outputs(12202));
    layer2_outputs(1716) <= not(layer1_outputs(5052));
    layer2_outputs(1717) <= (layer1_outputs(1734)) or (layer1_outputs(4494));
    layer2_outputs(1718) <= not((layer1_outputs(11443)) xor (layer1_outputs(7115)));
    layer2_outputs(1719) <= layer1_outputs(9095);
    layer2_outputs(1720) <= not(layer1_outputs(11040));
    layer2_outputs(1721) <= layer1_outputs(7092);
    layer2_outputs(1722) <= (layer1_outputs(5862)) or (layer1_outputs(5906));
    layer2_outputs(1723) <= layer1_outputs(1512);
    layer2_outputs(1724) <= not(layer1_outputs(3460));
    layer2_outputs(1725) <= layer1_outputs(4351);
    layer2_outputs(1726) <= not(layer1_outputs(4721));
    layer2_outputs(1727) <= not(layer1_outputs(8508));
    layer2_outputs(1728) <= layer1_outputs(11563);
    layer2_outputs(1729) <= layer1_outputs(5069);
    layer2_outputs(1730) <= layer1_outputs(7667);
    layer2_outputs(1731) <= not((layer1_outputs(4094)) xor (layer1_outputs(4928)));
    layer2_outputs(1732) <= not(layer1_outputs(8698));
    layer2_outputs(1733) <= (layer1_outputs(8654)) xor (layer1_outputs(5738));
    layer2_outputs(1734) <= not(layer1_outputs(12690));
    layer2_outputs(1735) <= not(layer1_outputs(9620));
    layer2_outputs(1736) <= '0';
    layer2_outputs(1737) <= not(layer1_outputs(1454)) or (layer1_outputs(3825));
    layer2_outputs(1738) <= layer1_outputs(3556);
    layer2_outputs(1739) <= not(layer1_outputs(9071)) or (layer1_outputs(6266));
    layer2_outputs(1740) <= not(layer1_outputs(12069)) or (layer1_outputs(7437));
    layer2_outputs(1741) <= not((layer1_outputs(1873)) and (layer1_outputs(5012)));
    layer2_outputs(1742) <= layer1_outputs(5263);
    layer2_outputs(1743) <= not((layer1_outputs(10114)) xor (layer1_outputs(12152)));
    layer2_outputs(1744) <= '1';
    layer2_outputs(1745) <= not(layer1_outputs(4377));
    layer2_outputs(1746) <= layer1_outputs(8866);
    layer2_outputs(1747) <= not(layer1_outputs(5736));
    layer2_outputs(1748) <= not((layer1_outputs(9525)) or (layer1_outputs(11938)));
    layer2_outputs(1749) <= not((layer1_outputs(12047)) xor (layer1_outputs(3024)));
    layer2_outputs(1750) <= layer1_outputs(8792);
    layer2_outputs(1751) <= not(layer1_outputs(4056)) or (layer1_outputs(328));
    layer2_outputs(1752) <= layer1_outputs(9474);
    layer2_outputs(1753) <= layer1_outputs(4964);
    layer2_outputs(1754) <= not(layer1_outputs(10135)) or (layer1_outputs(2176));
    layer2_outputs(1755) <= not(layer1_outputs(4448));
    layer2_outputs(1756) <= (layer1_outputs(2410)) and not (layer1_outputs(3398));
    layer2_outputs(1757) <= not(layer1_outputs(1495));
    layer2_outputs(1758) <= not((layer1_outputs(7318)) and (layer1_outputs(8887)));
    layer2_outputs(1759) <= not(layer1_outputs(1802));
    layer2_outputs(1760) <= layer1_outputs(7468);
    layer2_outputs(1761) <= not((layer1_outputs(11879)) xor (layer1_outputs(6769)));
    layer2_outputs(1762) <= not((layer1_outputs(4075)) or (layer1_outputs(10527)));
    layer2_outputs(1763) <= (layer1_outputs(5092)) and (layer1_outputs(9656));
    layer2_outputs(1764) <= (layer1_outputs(5865)) or (layer1_outputs(409));
    layer2_outputs(1765) <= layer1_outputs(5625);
    layer2_outputs(1766) <= layer1_outputs(2813);
    layer2_outputs(1767) <= not(layer1_outputs(3775));
    layer2_outputs(1768) <= not(layer1_outputs(9952));
    layer2_outputs(1769) <= not(layer1_outputs(9685));
    layer2_outputs(1770) <= layer1_outputs(313);
    layer2_outputs(1771) <= not((layer1_outputs(11069)) xor (layer1_outputs(10956)));
    layer2_outputs(1772) <= not((layer1_outputs(11687)) xor (layer1_outputs(11774)));
    layer2_outputs(1773) <= layer1_outputs(7025);
    layer2_outputs(1774) <= (layer1_outputs(427)) and (layer1_outputs(11527));
    layer2_outputs(1775) <= (layer1_outputs(4576)) or (layer1_outputs(6082));
    layer2_outputs(1776) <= not(layer1_outputs(8200)) or (layer1_outputs(9968));
    layer2_outputs(1777) <= not(layer1_outputs(7472));
    layer2_outputs(1778) <= not(layer1_outputs(10070));
    layer2_outputs(1779) <= not(layer1_outputs(7142));
    layer2_outputs(1780) <= not((layer1_outputs(2786)) xor (layer1_outputs(2361)));
    layer2_outputs(1781) <= layer1_outputs(9090);
    layer2_outputs(1782) <= layer1_outputs(2862);
    layer2_outputs(1783) <= not(layer1_outputs(9644));
    layer2_outputs(1784) <= not((layer1_outputs(5126)) xor (layer1_outputs(836)));
    layer2_outputs(1785) <= not(layer1_outputs(6766));
    layer2_outputs(1786) <= (layer1_outputs(10848)) and not (layer1_outputs(9480));
    layer2_outputs(1787) <= not(layer1_outputs(8977));
    layer2_outputs(1788) <= not((layer1_outputs(9756)) and (layer1_outputs(6909)));
    layer2_outputs(1789) <= not(layer1_outputs(1436));
    layer2_outputs(1790) <= layer1_outputs(7102);
    layer2_outputs(1791) <= not((layer1_outputs(8275)) or (layer1_outputs(1304)));
    layer2_outputs(1792) <= not(layer1_outputs(4310)) or (layer1_outputs(3078));
    layer2_outputs(1793) <= not((layer1_outputs(1789)) or (layer1_outputs(5024)));
    layer2_outputs(1794) <= not((layer1_outputs(11402)) xor (layer1_outputs(6081)));
    layer2_outputs(1795) <= not((layer1_outputs(2442)) xor (layer1_outputs(2663)));
    layer2_outputs(1796) <= (layer1_outputs(7082)) and not (layer1_outputs(10738));
    layer2_outputs(1797) <= layer1_outputs(10762);
    layer2_outputs(1798) <= not(layer1_outputs(11546)) or (layer1_outputs(8648));
    layer2_outputs(1799) <= not((layer1_outputs(12686)) and (layer1_outputs(11716)));
    layer2_outputs(1800) <= not((layer1_outputs(4980)) xor (layer1_outputs(9636)));
    layer2_outputs(1801) <= not(layer1_outputs(4934));
    layer2_outputs(1802) <= not(layer1_outputs(3846));
    layer2_outputs(1803) <= not((layer1_outputs(10760)) xor (layer1_outputs(9377)));
    layer2_outputs(1804) <= (layer1_outputs(6594)) and (layer1_outputs(7208));
    layer2_outputs(1805) <= layer1_outputs(1469);
    layer2_outputs(1806) <= (layer1_outputs(113)) and (layer1_outputs(2952));
    layer2_outputs(1807) <= (layer1_outputs(3450)) xor (layer1_outputs(8936));
    layer2_outputs(1808) <= layer1_outputs(7123);
    layer2_outputs(1809) <= not((layer1_outputs(499)) xor (layer1_outputs(10043)));
    layer2_outputs(1810) <= (layer1_outputs(4788)) xor (layer1_outputs(7238));
    layer2_outputs(1811) <= not(layer1_outputs(12371)) or (layer1_outputs(3286));
    layer2_outputs(1812) <= (layer1_outputs(3538)) and (layer1_outputs(8681));
    layer2_outputs(1813) <= layer1_outputs(3745);
    layer2_outputs(1814) <= layer1_outputs(5143);
    layer2_outputs(1815) <= layer1_outputs(6172);
    layer2_outputs(1816) <= (layer1_outputs(1525)) xor (layer1_outputs(5032));
    layer2_outputs(1817) <= layer1_outputs(10193);
    layer2_outputs(1818) <= not((layer1_outputs(1364)) and (layer1_outputs(643)));
    layer2_outputs(1819) <= not(layer1_outputs(11153));
    layer2_outputs(1820) <= '0';
    layer2_outputs(1821) <= layer1_outputs(11561);
    layer2_outputs(1822) <= (layer1_outputs(9007)) and not (layer1_outputs(4763));
    layer2_outputs(1823) <= not(layer1_outputs(7629));
    layer2_outputs(1824) <= (layer1_outputs(10870)) and not (layer1_outputs(7485));
    layer2_outputs(1825) <= (layer1_outputs(7690)) and (layer1_outputs(3302));
    layer2_outputs(1826) <= not(layer1_outputs(10251));
    layer2_outputs(1827) <= (layer1_outputs(7258)) and (layer1_outputs(8564));
    layer2_outputs(1828) <= not(layer1_outputs(4217));
    layer2_outputs(1829) <= (layer1_outputs(1530)) and not (layer1_outputs(7224));
    layer2_outputs(1830) <= not((layer1_outputs(3295)) xor (layer1_outputs(6271)));
    layer2_outputs(1831) <= layer1_outputs(8737);
    layer2_outputs(1832) <= not((layer1_outputs(3356)) and (layer1_outputs(7321)));
    layer2_outputs(1833) <= '1';
    layer2_outputs(1834) <= not(layer1_outputs(11159));
    layer2_outputs(1835) <= not(layer1_outputs(7222)) or (layer1_outputs(9727));
    layer2_outputs(1836) <= not(layer1_outputs(6443)) or (layer1_outputs(4129));
    layer2_outputs(1837) <= not(layer1_outputs(3182)) or (layer1_outputs(5490));
    layer2_outputs(1838) <= not(layer1_outputs(242));
    layer2_outputs(1839) <= not((layer1_outputs(2060)) and (layer1_outputs(4661)));
    layer2_outputs(1840) <= not(layer1_outputs(410));
    layer2_outputs(1841) <= layer1_outputs(6894);
    layer2_outputs(1842) <= layer1_outputs(8849);
    layer2_outputs(1843) <= (layer1_outputs(11971)) and (layer1_outputs(8938));
    layer2_outputs(1844) <= layer1_outputs(6294);
    layer2_outputs(1845) <= layer1_outputs(3892);
    layer2_outputs(1846) <= not(layer1_outputs(4215));
    layer2_outputs(1847) <= (layer1_outputs(11512)) and not (layer1_outputs(11965));
    layer2_outputs(1848) <= (layer1_outputs(11262)) and not (layer1_outputs(678));
    layer2_outputs(1849) <= not((layer1_outputs(11327)) xor (layer1_outputs(7035)));
    layer2_outputs(1850) <= not((layer1_outputs(4631)) xor (layer1_outputs(5093)));
    layer2_outputs(1851) <= not((layer1_outputs(10734)) and (layer1_outputs(3567)));
    layer2_outputs(1852) <= not(layer1_outputs(12051)) or (layer1_outputs(3736));
    layer2_outputs(1853) <= layer1_outputs(6769);
    layer2_outputs(1854) <= (layer1_outputs(11591)) and (layer1_outputs(2579));
    layer2_outputs(1855) <= not(layer1_outputs(620));
    layer2_outputs(1856) <= (layer1_outputs(9072)) xor (layer1_outputs(10788));
    layer2_outputs(1857) <= not(layer1_outputs(12483));
    layer2_outputs(1858) <= '1';
    layer2_outputs(1859) <= not((layer1_outputs(12336)) xor (layer1_outputs(10099)));
    layer2_outputs(1860) <= not(layer1_outputs(6218)) or (layer1_outputs(11335));
    layer2_outputs(1861) <= layer1_outputs(217);
    layer2_outputs(1862) <= not((layer1_outputs(12617)) or (layer1_outputs(9781)));
    layer2_outputs(1863) <= layer1_outputs(4783);
    layer2_outputs(1864) <= layer1_outputs(8501);
    layer2_outputs(1865) <= (layer1_outputs(1243)) and not (layer1_outputs(9166));
    layer2_outputs(1866) <= (layer1_outputs(4740)) xor (layer1_outputs(447));
    layer2_outputs(1867) <= not(layer1_outputs(6514)) or (layer1_outputs(7205));
    layer2_outputs(1868) <= layer1_outputs(1829);
    layer2_outputs(1869) <= not(layer1_outputs(12688));
    layer2_outputs(1870) <= not(layer1_outputs(5589));
    layer2_outputs(1871) <= layer1_outputs(2134);
    layer2_outputs(1872) <= not(layer1_outputs(9439));
    layer2_outputs(1873) <= layer1_outputs(10555);
    layer2_outputs(1874) <= (layer1_outputs(7856)) xor (layer1_outputs(1172));
    layer2_outputs(1875) <= not(layer1_outputs(7435)) or (layer1_outputs(4417));
    layer2_outputs(1876) <= not((layer1_outputs(4406)) or (layer1_outputs(380)));
    layer2_outputs(1877) <= (layer1_outputs(1844)) and not (layer1_outputs(4547));
    layer2_outputs(1878) <= layer1_outputs(11679);
    layer2_outputs(1879) <= not((layer1_outputs(3252)) and (layer1_outputs(3589)));
    layer2_outputs(1880) <= (layer1_outputs(9232)) and not (layer1_outputs(6561));
    layer2_outputs(1881) <= layer1_outputs(6395);
    layer2_outputs(1882) <= (layer1_outputs(10909)) or (layer1_outputs(12676));
    layer2_outputs(1883) <= (layer1_outputs(9164)) and not (layer1_outputs(10597));
    layer2_outputs(1884) <= (layer1_outputs(5615)) xor (layer1_outputs(1619));
    layer2_outputs(1885) <= not(layer1_outputs(1332));
    layer2_outputs(1886) <= layer1_outputs(3694);
    layer2_outputs(1887) <= (layer1_outputs(3983)) and not (layer1_outputs(2332));
    layer2_outputs(1888) <= (layer1_outputs(3114)) xor (layer1_outputs(9039));
    layer2_outputs(1889) <= not(layer1_outputs(3684));
    layer2_outputs(1890) <= layer1_outputs(12158);
    layer2_outputs(1891) <= not(layer1_outputs(6614));
    layer2_outputs(1892) <= not(layer1_outputs(8186)) or (layer1_outputs(4192));
    layer2_outputs(1893) <= not((layer1_outputs(7921)) or (layer1_outputs(3129)));
    layer2_outputs(1894) <= not((layer1_outputs(9367)) xor (layer1_outputs(9272)));
    layer2_outputs(1895) <= not(layer1_outputs(7751));
    layer2_outputs(1896) <= layer1_outputs(3577);
    layer2_outputs(1897) <= layer1_outputs(3258);
    layer2_outputs(1898) <= not((layer1_outputs(7058)) xor (layer1_outputs(3241)));
    layer2_outputs(1899) <= not(layer1_outputs(1408)) or (layer1_outputs(11656));
    layer2_outputs(1900) <= (layer1_outputs(9972)) and not (layer1_outputs(10858));
    layer2_outputs(1901) <= (layer1_outputs(6131)) xor (layer1_outputs(4770));
    layer2_outputs(1902) <= not(layer1_outputs(11519));
    layer2_outputs(1903) <= not(layer1_outputs(11551));
    layer2_outputs(1904) <= layer1_outputs(12261);
    layer2_outputs(1905) <= (layer1_outputs(9590)) and not (layer1_outputs(2319));
    layer2_outputs(1906) <= (layer1_outputs(5393)) xor (layer1_outputs(8892));
    layer2_outputs(1907) <= layer1_outputs(7270);
    layer2_outputs(1908) <= layer1_outputs(8897);
    layer2_outputs(1909) <= not((layer1_outputs(487)) or (layer1_outputs(1800)));
    layer2_outputs(1910) <= not((layer1_outputs(11453)) and (layer1_outputs(10573)));
    layer2_outputs(1911) <= not(layer1_outputs(4622));
    layer2_outputs(1912) <= not(layer1_outputs(6918));
    layer2_outputs(1913) <= layer1_outputs(2164);
    layer2_outputs(1914) <= layer1_outputs(5669);
    layer2_outputs(1915) <= not(layer1_outputs(9161));
    layer2_outputs(1916) <= '1';
    layer2_outputs(1917) <= (layer1_outputs(10020)) and not (layer1_outputs(2231));
    layer2_outputs(1918) <= not(layer1_outputs(10278));
    layer2_outputs(1919) <= not(layer1_outputs(267));
    layer2_outputs(1920) <= not(layer1_outputs(11114)) or (layer1_outputs(6898));
    layer2_outputs(1921) <= layer1_outputs(4174);
    layer2_outputs(1922) <= layer1_outputs(6862);
    layer2_outputs(1923) <= layer1_outputs(559);
    layer2_outputs(1924) <= (layer1_outputs(2616)) xor (layer1_outputs(354));
    layer2_outputs(1925) <= layer1_outputs(1053);
    layer2_outputs(1926) <= not((layer1_outputs(9299)) and (layer1_outputs(3206)));
    layer2_outputs(1927) <= layer1_outputs(2037);
    layer2_outputs(1928) <= layer1_outputs(10894);
    layer2_outputs(1929) <= layer1_outputs(12241);
    layer2_outputs(1930) <= not((layer1_outputs(5927)) or (layer1_outputs(2018)));
    layer2_outputs(1931) <= (layer1_outputs(6276)) and (layer1_outputs(3502));
    layer2_outputs(1932) <= (layer1_outputs(8448)) and not (layer1_outputs(7404));
    layer2_outputs(1933) <= (layer1_outputs(2134)) and not (layer1_outputs(8118));
    layer2_outputs(1934) <= not(layer1_outputs(1004));
    layer2_outputs(1935) <= not(layer1_outputs(3270));
    layer2_outputs(1936) <= (layer1_outputs(6038)) and not (layer1_outputs(4564));
    layer2_outputs(1937) <= layer1_outputs(1101);
    layer2_outputs(1938) <= (layer1_outputs(3083)) and not (layer1_outputs(4941));
    layer2_outputs(1939) <= not(layer1_outputs(4220));
    layer2_outputs(1940) <= not(layer1_outputs(6469));
    layer2_outputs(1941) <= layer1_outputs(2596);
    layer2_outputs(1942) <= layer1_outputs(5942);
    layer2_outputs(1943) <= (layer1_outputs(871)) and not (layer1_outputs(10997));
    layer2_outputs(1944) <= not(layer1_outputs(2305)) or (layer1_outputs(11788));
    layer2_outputs(1945) <= layer1_outputs(1255);
    layer2_outputs(1946) <= not(layer1_outputs(11215)) or (layer1_outputs(8177));
    layer2_outputs(1947) <= (layer1_outputs(4002)) or (layer1_outputs(8378));
    layer2_outputs(1948) <= not((layer1_outputs(9222)) xor (layer1_outputs(720)));
    layer2_outputs(1949) <= layer1_outputs(8036);
    layer2_outputs(1950) <= (layer1_outputs(8483)) and not (layer1_outputs(3662));
    layer2_outputs(1951) <= not(layer1_outputs(4165));
    layer2_outputs(1952) <= not((layer1_outputs(3808)) xor (layer1_outputs(2460)));
    layer2_outputs(1953) <= not((layer1_outputs(3048)) or (layer1_outputs(5453)));
    layer2_outputs(1954) <= (layer1_outputs(5292)) and not (layer1_outputs(3762));
    layer2_outputs(1955) <= not(layer1_outputs(10577));
    layer2_outputs(1956) <= layer1_outputs(2116);
    layer2_outputs(1957) <= not(layer1_outputs(8761));
    layer2_outputs(1958) <= not(layer1_outputs(4382)) or (layer1_outputs(12357));
    layer2_outputs(1959) <= (layer1_outputs(2890)) and (layer1_outputs(2527));
    layer2_outputs(1960) <= (layer1_outputs(8604)) and not (layer1_outputs(2591));
    layer2_outputs(1961) <= not(layer1_outputs(10216));
    layer2_outputs(1962) <= not(layer1_outputs(4947));
    layer2_outputs(1963) <= not(layer1_outputs(12345));
    layer2_outputs(1964) <= layer1_outputs(2895);
    layer2_outputs(1965) <= not(layer1_outputs(8579));
    layer2_outputs(1966) <= not(layer1_outputs(2254));
    layer2_outputs(1967) <= (layer1_outputs(3810)) and not (layer1_outputs(5110));
    layer2_outputs(1968) <= layer1_outputs(106);
    layer2_outputs(1969) <= not(layer1_outputs(4359));
    layer2_outputs(1970) <= not((layer1_outputs(4818)) or (layer1_outputs(11069)));
    layer2_outputs(1971) <= layer1_outputs(9538);
    layer2_outputs(1972) <= (layer1_outputs(1280)) and not (layer1_outputs(4549));
    layer2_outputs(1973) <= not(layer1_outputs(7751));
    layer2_outputs(1974) <= not(layer1_outputs(4759)) or (layer1_outputs(6451));
    layer2_outputs(1975) <= (layer1_outputs(731)) and (layer1_outputs(12767));
    layer2_outputs(1976) <= layer1_outputs(11682);
    layer2_outputs(1977) <= not(layer1_outputs(3214));
    layer2_outputs(1978) <= not(layer1_outputs(6289));
    layer2_outputs(1979) <= not((layer1_outputs(270)) and (layer1_outputs(8360)));
    layer2_outputs(1980) <= not(layer1_outputs(3900));
    layer2_outputs(1981) <= layer1_outputs(4337);
    layer2_outputs(1982) <= layer1_outputs(8347);
    layer2_outputs(1983) <= not(layer1_outputs(7719));
    layer2_outputs(1984) <= not((layer1_outputs(2183)) or (layer1_outputs(5264)));
    layer2_outputs(1985) <= not(layer1_outputs(1313));
    layer2_outputs(1986) <= not(layer1_outputs(12177));
    layer2_outputs(1987) <= layer1_outputs(9395);
    layer2_outputs(1988) <= layer1_outputs(7162);
    layer2_outputs(1989) <= layer1_outputs(5106);
    layer2_outputs(1990) <= layer1_outputs(9369);
    layer2_outputs(1991) <= (layer1_outputs(4392)) or (layer1_outputs(2449));
    layer2_outputs(1992) <= not((layer1_outputs(3839)) and (layer1_outputs(12785)));
    layer2_outputs(1993) <= not(layer1_outputs(12130));
    layer2_outputs(1994) <= layer1_outputs(5962);
    layer2_outputs(1995) <= layer1_outputs(1558);
    layer2_outputs(1996) <= not((layer1_outputs(5331)) or (layer1_outputs(2959)));
    layer2_outputs(1997) <= not((layer1_outputs(2383)) and (layer1_outputs(8348)));
    layer2_outputs(1998) <= (layer1_outputs(1856)) and not (layer1_outputs(9920));
    layer2_outputs(1999) <= not(layer1_outputs(6643));
    layer2_outputs(2000) <= (layer1_outputs(3972)) or (layer1_outputs(12405));
    layer2_outputs(2001) <= not((layer1_outputs(7330)) xor (layer1_outputs(8851)));
    layer2_outputs(2002) <= not(layer1_outputs(8049));
    layer2_outputs(2003) <= not((layer1_outputs(7477)) xor (layer1_outputs(2396)));
    layer2_outputs(2004) <= (layer1_outputs(5695)) xor (layer1_outputs(5422));
    layer2_outputs(2005) <= layer1_outputs(10998);
    layer2_outputs(2006) <= not((layer1_outputs(11041)) or (layer1_outputs(187)));
    layer2_outputs(2007) <= not((layer1_outputs(4122)) xor (layer1_outputs(7819)));
    layer2_outputs(2008) <= (layer1_outputs(9080)) xor (layer1_outputs(3145));
    layer2_outputs(2009) <= layer1_outputs(2457);
    layer2_outputs(2010) <= layer1_outputs(107);
    layer2_outputs(2011) <= (layer1_outputs(4824)) xor (layer1_outputs(7142));
    layer2_outputs(2012) <= (layer1_outputs(9904)) or (layer1_outputs(6973));
    layer2_outputs(2013) <= not(layer1_outputs(4294)) or (layer1_outputs(2689));
    layer2_outputs(2014) <= not((layer1_outputs(7606)) or (layer1_outputs(7634)));
    layer2_outputs(2015) <= (layer1_outputs(5637)) and not (layer1_outputs(161));
    layer2_outputs(2016) <= not((layer1_outputs(3459)) xor (layer1_outputs(11057)));
    layer2_outputs(2017) <= not((layer1_outputs(2049)) xor (layer1_outputs(7851)));
    layer2_outputs(2018) <= '1';
    layer2_outputs(2019) <= not(layer1_outputs(548));
    layer2_outputs(2020) <= (layer1_outputs(4881)) xor (layer1_outputs(333));
    layer2_outputs(2021) <= not(layer1_outputs(6940));
    layer2_outputs(2022) <= not(layer1_outputs(1051));
    layer2_outputs(2023) <= not((layer1_outputs(3316)) or (layer1_outputs(4401)));
    layer2_outputs(2024) <= not((layer1_outputs(555)) or (layer1_outputs(209)));
    layer2_outputs(2025) <= layer1_outputs(6024);
    layer2_outputs(2026) <= layer1_outputs(1920);
    layer2_outputs(2027) <= (layer1_outputs(3523)) xor (layer1_outputs(258));
    layer2_outputs(2028) <= not(layer1_outputs(4020));
    layer2_outputs(2029) <= (layer1_outputs(8116)) and not (layer1_outputs(5654));
    layer2_outputs(2030) <= (layer1_outputs(5701)) and not (layer1_outputs(9147));
    layer2_outputs(2031) <= not(layer1_outputs(350));
    layer2_outputs(2032) <= not(layer1_outputs(6951));
    layer2_outputs(2033) <= layer1_outputs(5073);
    layer2_outputs(2034) <= not(layer1_outputs(10378)) or (layer1_outputs(1959));
    layer2_outputs(2035) <= layer1_outputs(1046);
    layer2_outputs(2036) <= layer1_outputs(3586);
    layer2_outputs(2037) <= layer1_outputs(94);
    layer2_outputs(2038) <= not((layer1_outputs(2178)) and (layer1_outputs(2292)));
    layer2_outputs(2039) <= layer1_outputs(8915);
    layer2_outputs(2040) <= not(layer1_outputs(9439));
    layer2_outputs(2041) <= (layer1_outputs(5690)) and not (layer1_outputs(9176));
    layer2_outputs(2042) <= (layer1_outputs(3024)) xor (layer1_outputs(10006));
    layer2_outputs(2043) <= not(layer1_outputs(12409));
    layer2_outputs(2044) <= not(layer1_outputs(5881)) or (layer1_outputs(3600));
    layer2_outputs(2045) <= (layer1_outputs(1175)) and not (layer1_outputs(4290));
    layer2_outputs(2046) <= layer1_outputs(6310);
    layer2_outputs(2047) <= not(layer1_outputs(8480)) or (layer1_outputs(10250));
    layer2_outputs(2048) <= layer1_outputs(12685);
    layer2_outputs(2049) <= layer1_outputs(3552);
    layer2_outputs(2050) <= layer1_outputs(4599);
    layer2_outputs(2051) <= not(layer1_outputs(12194));
    layer2_outputs(2052) <= layer1_outputs(7281);
    layer2_outputs(2053) <= (layer1_outputs(10712)) and not (layer1_outputs(442));
    layer2_outputs(2054) <= not(layer1_outputs(8071));
    layer2_outputs(2055) <= (layer1_outputs(7057)) xor (layer1_outputs(2548));
    layer2_outputs(2056) <= layer1_outputs(5987);
    layer2_outputs(2057) <= not(layer1_outputs(3291));
    layer2_outputs(2058) <= (layer1_outputs(12280)) or (layer1_outputs(10961));
    layer2_outputs(2059) <= not(layer1_outputs(11121));
    layer2_outputs(2060) <= (layer1_outputs(3947)) and not (layer1_outputs(3260));
    layer2_outputs(2061) <= layer1_outputs(10698);
    layer2_outputs(2062) <= not(layer1_outputs(6708));
    layer2_outputs(2063) <= not(layer1_outputs(11614));
    layer2_outputs(2064) <= not(layer1_outputs(5680));
    layer2_outputs(2065) <= not(layer1_outputs(6221));
    layer2_outputs(2066) <= (layer1_outputs(6945)) or (layer1_outputs(5707));
    layer2_outputs(2067) <= (layer1_outputs(6978)) xor (layer1_outputs(6604));
    layer2_outputs(2068) <= layer1_outputs(3910);
    layer2_outputs(2069) <= not(layer1_outputs(2758));
    layer2_outputs(2070) <= not((layer1_outputs(1464)) xor (layer1_outputs(2533)));
    layer2_outputs(2071) <= (layer1_outputs(6198)) xor (layer1_outputs(8540));
    layer2_outputs(2072) <= not(layer1_outputs(8462));
    layer2_outputs(2073) <= layer1_outputs(11356);
    layer2_outputs(2074) <= not(layer1_outputs(3144));
    layer2_outputs(2075) <= layer1_outputs(11850);
    layer2_outputs(2076) <= layer1_outputs(7656);
    layer2_outputs(2077) <= layer1_outputs(12341);
    layer2_outputs(2078) <= not((layer1_outputs(9790)) and (layer1_outputs(875)));
    layer2_outputs(2079) <= (layer1_outputs(7819)) and not (layer1_outputs(916));
    layer2_outputs(2080) <= layer1_outputs(9101);
    layer2_outputs(2081) <= layer1_outputs(8918);
    layer2_outputs(2082) <= not(layer1_outputs(4858));
    layer2_outputs(2083) <= layer1_outputs(2182);
    layer2_outputs(2084) <= (layer1_outputs(5385)) or (layer1_outputs(652));
    layer2_outputs(2085) <= layer1_outputs(3288);
    layer2_outputs(2086) <= (layer1_outputs(5032)) and not (layer1_outputs(7762));
    layer2_outputs(2087) <= not(layer1_outputs(3772));
    layer2_outputs(2088) <= not(layer1_outputs(902));
    layer2_outputs(2089) <= not((layer1_outputs(10108)) and (layer1_outputs(11277)));
    layer2_outputs(2090) <= not(layer1_outputs(5418));
    layer2_outputs(2091) <= not((layer1_outputs(2743)) xor (layer1_outputs(10474)));
    layer2_outputs(2092) <= not(layer1_outputs(9515)) or (layer1_outputs(6543));
    layer2_outputs(2093) <= not(layer1_outputs(3130));
    layer2_outputs(2094) <= not((layer1_outputs(4141)) and (layer1_outputs(231)));
    layer2_outputs(2095) <= '1';
    layer2_outputs(2096) <= layer1_outputs(1339);
    layer2_outputs(2097) <= not((layer1_outputs(8946)) xor (layer1_outputs(6209)));
    layer2_outputs(2098) <= (layer1_outputs(12221)) and not (layer1_outputs(10507));
    layer2_outputs(2099) <= (layer1_outputs(2221)) xor (layer1_outputs(6573));
    layer2_outputs(2100) <= not((layer1_outputs(8221)) xor (layer1_outputs(3527)));
    layer2_outputs(2101) <= not(layer1_outputs(5047));
    layer2_outputs(2102) <= not((layer1_outputs(4766)) xor (layer1_outputs(1671)));
    layer2_outputs(2103) <= layer1_outputs(6356);
    layer2_outputs(2104) <= not((layer1_outputs(9278)) and (layer1_outputs(6811)));
    layer2_outputs(2105) <= not(layer1_outputs(5313)) or (layer1_outputs(3924));
    layer2_outputs(2106) <= layer1_outputs(2318);
    layer2_outputs(2107) <= layer1_outputs(1385);
    layer2_outputs(2108) <= (layer1_outputs(4624)) and (layer1_outputs(9739));
    layer2_outputs(2109) <= layer1_outputs(11177);
    layer2_outputs(2110) <= (layer1_outputs(10464)) and not (layer1_outputs(6009));
    layer2_outputs(2111) <= not(layer1_outputs(5498)) or (layer1_outputs(2625));
    layer2_outputs(2112) <= layer1_outputs(6744);
    layer2_outputs(2113) <= not(layer1_outputs(4301));
    layer2_outputs(2114) <= not(layer1_outputs(12691)) or (layer1_outputs(10991));
    layer2_outputs(2115) <= (layer1_outputs(1443)) and not (layer1_outputs(5366));
    layer2_outputs(2116) <= not((layer1_outputs(9717)) xor (layer1_outputs(7965)));
    layer2_outputs(2117) <= layer1_outputs(11399);
    layer2_outputs(2118) <= not(layer1_outputs(8913)) or (layer1_outputs(4933));
    layer2_outputs(2119) <= not((layer1_outputs(7879)) or (layer1_outputs(1722)));
    layer2_outputs(2120) <= layer1_outputs(241);
    layer2_outputs(2121) <= layer1_outputs(464);
    layer2_outputs(2122) <= layer1_outputs(4005);
    layer2_outputs(2123) <= '1';
    layer2_outputs(2124) <= not(layer1_outputs(10319));
    layer2_outputs(2125) <= not((layer1_outputs(10896)) or (layer1_outputs(456)));
    layer2_outputs(2126) <= not((layer1_outputs(4198)) xor (layer1_outputs(6219)));
    layer2_outputs(2127) <= (layer1_outputs(6542)) or (layer1_outputs(7953));
    layer2_outputs(2128) <= (layer1_outputs(9794)) and (layer1_outputs(5832));
    layer2_outputs(2129) <= not(layer1_outputs(2555));
    layer2_outputs(2130) <= layer1_outputs(12124);
    layer2_outputs(2131) <= not((layer1_outputs(1684)) xor (layer1_outputs(998)));
    layer2_outputs(2132) <= not((layer1_outputs(9366)) or (layer1_outputs(12530)));
    layer2_outputs(2133) <= (layer1_outputs(10831)) and not (layer1_outputs(10496));
    layer2_outputs(2134) <= not((layer1_outputs(9657)) and (layer1_outputs(4843)));
    layer2_outputs(2135) <= (layer1_outputs(5454)) and not (layer1_outputs(5579));
    layer2_outputs(2136) <= layer1_outputs(8074);
    layer2_outputs(2137) <= layer1_outputs(8970);
    layer2_outputs(2138) <= not(layer1_outputs(9885));
    layer2_outputs(2139) <= layer1_outputs(2737);
    layer2_outputs(2140) <= (layer1_outputs(6913)) and not (layer1_outputs(8872));
    layer2_outputs(2141) <= not(layer1_outputs(5164)) or (layer1_outputs(8349));
    layer2_outputs(2142) <= not((layer1_outputs(10899)) and (layer1_outputs(4816)));
    layer2_outputs(2143) <= not((layer1_outputs(6305)) xor (layer1_outputs(9205)));
    layer2_outputs(2144) <= not((layer1_outputs(5513)) and (layer1_outputs(384)));
    layer2_outputs(2145) <= not(layer1_outputs(10996));
    layer2_outputs(2146) <= not((layer1_outputs(9776)) xor (layer1_outputs(3734)));
    layer2_outputs(2147) <= (layer1_outputs(6028)) xor (layer1_outputs(10364));
    layer2_outputs(2148) <= (layer1_outputs(8262)) or (layer1_outputs(7768));
    layer2_outputs(2149) <= layer1_outputs(12635);
    layer2_outputs(2150) <= not(layer1_outputs(7525));
    layer2_outputs(2151) <= layer1_outputs(11124);
    layer2_outputs(2152) <= not(layer1_outputs(8035));
    layer2_outputs(2153) <= not(layer1_outputs(3500)) or (layer1_outputs(4128));
    layer2_outputs(2154) <= not(layer1_outputs(12579));
    layer2_outputs(2155) <= not((layer1_outputs(2936)) xor (layer1_outputs(7371)));
    layer2_outputs(2156) <= (layer1_outputs(8154)) xor (layer1_outputs(9962));
    layer2_outputs(2157) <= not(layer1_outputs(11082));
    layer2_outputs(2158) <= not(layer1_outputs(8172));
    layer2_outputs(2159) <= not(layer1_outputs(10662)) or (layer1_outputs(2490));
    layer2_outputs(2160) <= layer1_outputs(11593);
    layer2_outputs(2161) <= not((layer1_outputs(5563)) xor (layer1_outputs(1216)));
    layer2_outputs(2162) <= not(layer1_outputs(4986));
    layer2_outputs(2163) <= layer1_outputs(9360);
    layer2_outputs(2164) <= not(layer1_outputs(1487));
    layer2_outputs(2165) <= (layer1_outputs(11531)) xor (layer1_outputs(5137));
    layer2_outputs(2166) <= not(layer1_outputs(1206));
    layer2_outputs(2167) <= not((layer1_outputs(2384)) or (layer1_outputs(3883)));
    layer2_outputs(2168) <= layer1_outputs(11652);
    layer2_outputs(2169) <= layer1_outputs(7972);
    layer2_outputs(2170) <= (layer1_outputs(10780)) and not (layer1_outputs(151));
    layer2_outputs(2171) <= (layer1_outputs(445)) and (layer1_outputs(4833));
    layer2_outputs(2172) <= layer1_outputs(1865);
    layer2_outputs(2173) <= layer1_outputs(12795);
    layer2_outputs(2174) <= not(layer1_outputs(5325)) or (layer1_outputs(4427));
    layer2_outputs(2175) <= not(layer1_outputs(7019)) or (layer1_outputs(9958));
    layer2_outputs(2176) <= not((layer1_outputs(12381)) or (layer1_outputs(4508)));
    layer2_outputs(2177) <= (layer1_outputs(579)) and not (layer1_outputs(672));
    layer2_outputs(2178) <= not(layer1_outputs(1372));
    layer2_outputs(2179) <= not((layer1_outputs(9048)) and (layer1_outputs(2668)));
    layer2_outputs(2180) <= (layer1_outputs(2301)) and not (layer1_outputs(5828));
    layer2_outputs(2181) <= not((layer1_outputs(7576)) xor (layer1_outputs(8687)));
    layer2_outputs(2182) <= not(layer1_outputs(12544));
    layer2_outputs(2183) <= not(layer1_outputs(6048)) or (layer1_outputs(10196));
    layer2_outputs(2184) <= not(layer1_outputs(11396));
    layer2_outputs(2185) <= (layer1_outputs(2110)) xor (layer1_outputs(10528));
    layer2_outputs(2186) <= not(layer1_outputs(2195)) or (layer1_outputs(8166));
    layer2_outputs(2187) <= (layer1_outputs(8587)) xor (layer1_outputs(9372));
    layer2_outputs(2188) <= layer1_outputs(5864);
    layer2_outputs(2189) <= not((layer1_outputs(8730)) and (layer1_outputs(624)));
    layer2_outputs(2190) <= not(layer1_outputs(9680));
    layer2_outputs(2191) <= (layer1_outputs(2265)) or (layer1_outputs(1132));
    layer2_outputs(2192) <= not(layer1_outputs(12375));
    layer2_outputs(2193) <= (layer1_outputs(1331)) xor (layer1_outputs(10811));
    layer2_outputs(2194) <= (layer1_outputs(12077)) and not (layer1_outputs(7818));
    layer2_outputs(2195) <= layer1_outputs(9819);
    layer2_outputs(2196) <= layer1_outputs(12084);
    layer2_outputs(2197) <= (layer1_outputs(4189)) and not (layer1_outputs(12589));
    layer2_outputs(2198) <= not(layer1_outputs(2032));
    layer2_outputs(2199) <= (layer1_outputs(5326)) xor (layer1_outputs(10807));
    layer2_outputs(2200) <= not(layer1_outputs(7997));
    layer2_outputs(2201) <= (layer1_outputs(7780)) xor (layer1_outputs(635));
    layer2_outputs(2202) <= not((layer1_outputs(6104)) xor (layer1_outputs(9420)));
    layer2_outputs(2203) <= not(layer1_outputs(4657));
    layer2_outputs(2204) <= not(layer1_outputs(1890));
    layer2_outputs(2205) <= (layer1_outputs(1753)) and not (layer1_outputs(6303));
    layer2_outputs(2206) <= (layer1_outputs(6490)) xor (layer1_outputs(7436));
    layer2_outputs(2207) <= layer1_outputs(4936);
    layer2_outputs(2208) <= (layer1_outputs(7619)) and (layer1_outputs(1718));
    layer2_outputs(2209) <= not(layer1_outputs(6599));
    layer2_outputs(2210) <= layer1_outputs(7475);
    layer2_outputs(2211) <= not(layer1_outputs(4382)) or (layer1_outputs(8011));
    layer2_outputs(2212) <= not(layer1_outputs(6341));
    layer2_outputs(2213) <= not(layer1_outputs(2933));
    layer2_outputs(2214) <= not(layer1_outputs(6164));
    layer2_outputs(2215) <= (layer1_outputs(10402)) xor (layer1_outputs(4619));
    layer2_outputs(2216) <= (layer1_outputs(7077)) xor (layer1_outputs(3521));
    layer2_outputs(2217) <= layer1_outputs(10858);
    layer2_outputs(2218) <= not((layer1_outputs(5739)) or (layer1_outputs(8877)));
    layer2_outputs(2219) <= not(layer1_outputs(5087));
    layer2_outputs(2220) <= layer1_outputs(6441);
    layer2_outputs(2221) <= layer1_outputs(7420);
    layer2_outputs(2222) <= layer1_outputs(8779);
    layer2_outputs(2223) <= layer1_outputs(452);
    layer2_outputs(2224) <= layer1_outputs(12135);
    layer2_outputs(2225) <= not(layer1_outputs(10479));
    layer2_outputs(2226) <= (layer1_outputs(5589)) xor (layer1_outputs(3304));
    layer2_outputs(2227) <= layer1_outputs(2851);
    layer2_outputs(2228) <= (layer1_outputs(8292)) xor (layer1_outputs(11118));
    layer2_outputs(2229) <= not(layer1_outputs(2205));
    layer2_outputs(2230) <= layer1_outputs(3635);
    layer2_outputs(2231) <= not((layer1_outputs(8350)) or (layer1_outputs(5861)));
    layer2_outputs(2232) <= not(layer1_outputs(1181));
    layer2_outputs(2233) <= layer1_outputs(10397);
    layer2_outputs(2234) <= layer1_outputs(5324);
    layer2_outputs(2235) <= (layer1_outputs(52)) and not (layer1_outputs(1648));
    layer2_outputs(2236) <= layer1_outputs(1264);
    layer2_outputs(2237) <= not(layer1_outputs(7177));
    layer2_outputs(2238) <= not(layer1_outputs(7590));
    layer2_outputs(2239) <= not(layer1_outputs(7392)) or (layer1_outputs(1220));
    layer2_outputs(2240) <= (layer1_outputs(5373)) and (layer1_outputs(6173));
    layer2_outputs(2241) <= (layer1_outputs(11693)) and not (layer1_outputs(11807));
    layer2_outputs(2242) <= not(layer1_outputs(9967));
    layer2_outputs(2243) <= '0';
    layer2_outputs(2244) <= (layer1_outputs(4103)) or (layer1_outputs(9748));
    layer2_outputs(2245) <= not(layer1_outputs(8257));
    layer2_outputs(2246) <= not(layer1_outputs(960));
    layer2_outputs(2247) <= not((layer1_outputs(9352)) or (layer1_outputs(10897)));
    layer2_outputs(2248) <= layer1_outputs(3926);
    layer2_outputs(2249) <= layer1_outputs(11170);
    layer2_outputs(2250) <= layer1_outputs(11550);
    layer2_outputs(2251) <= not((layer1_outputs(8581)) and (layer1_outputs(8157)));
    layer2_outputs(2252) <= layer1_outputs(12356);
    layer2_outputs(2253) <= layer1_outputs(10546);
    layer2_outputs(2254) <= layer1_outputs(1239);
    layer2_outputs(2255) <= not(layer1_outputs(6610));
    layer2_outputs(2256) <= (layer1_outputs(4411)) and not (layer1_outputs(7630));
    layer2_outputs(2257) <= '1';
    layer2_outputs(2258) <= layer1_outputs(5925);
    layer2_outputs(2259) <= (layer1_outputs(5936)) and (layer1_outputs(5878));
    layer2_outputs(2260) <= (layer1_outputs(3541)) and not (layer1_outputs(11390));
    layer2_outputs(2261) <= not(layer1_outputs(6441));
    layer2_outputs(2262) <= layer1_outputs(4451);
    layer2_outputs(2263) <= layer1_outputs(4586);
    layer2_outputs(2264) <= not((layer1_outputs(519)) xor (layer1_outputs(12097)));
    layer2_outputs(2265) <= (layer1_outputs(6713)) or (layer1_outputs(2141));
    layer2_outputs(2266) <= not(layer1_outputs(9896));
    layer2_outputs(2267) <= not((layer1_outputs(6684)) xor (layer1_outputs(9775)));
    layer2_outputs(2268) <= not(layer1_outputs(5812)) or (layer1_outputs(4101));
    layer2_outputs(2269) <= layer1_outputs(7013);
    layer2_outputs(2270) <= (layer1_outputs(4310)) and (layer1_outputs(8269));
    layer2_outputs(2271) <= (layer1_outputs(3828)) and not (layer1_outputs(3416));
    layer2_outputs(2272) <= layer1_outputs(1153);
    layer2_outputs(2273) <= not(layer1_outputs(6558));
    layer2_outputs(2274) <= layer1_outputs(248);
    layer2_outputs(2275) <= not(layer1_outputs(3168)) or (layer1_outputs(6600));
    layer2_outputs(2276) <= not(layer1_outputs(11017)) or (layer1_outputs(3855));
    layer2_outputs(2277) <= not((layer1_outputs(3698)) or (layer1_outputs(9188)));
    layer2_outputs(2278) <= not(layer1_outputs(5731)) or (layer1_outputs(3764));
    layer2_outputs(2279) <= layer1_outputs(9893);
    layer2_outputs(2280) <= not(layer1_outputs(10551));
    layer2_outputs(2281) <= layer1_outputs(4238);
    layer2_outputs(2282) <= layer1_outputs(11699);
    layer2_outputs(2283) <= layer1_outputs(9189);
    layer2_outputs(2284) <= not((layer1_outputs(8755)) xor (layer1_outputs(4493)));
    layer2_outputs(2285) <= (layer1_outputs(6670)) xor (layer1_outputs(11777));
    layer2_outputs(2286) <= layer1_outputs(7557);
    layer2_outputs(2287) <= not(layer1_outputs(8690));
    layer2_outputs(2288) <= not(layer1_outputs(9767)) or (layer1_outputs(2287));
    layer2_outputs(2289) <= not((layer1_outputs(4780)) and (layer1_outputs(4254)));
    layer2_outputs(2290) <= not(layer1_outputs(5184));
    layer2_outputs(2291) <= not(layer1_outputs(10711));
    layer2_outputs(2292) <= not(layer1_outputs(5077));
    layer2_outputs(2293) <= not((layer1_outputs(6671)) xor (layer1_outputs(12253)));
    layer2_outputs(2294) <= (layer1_outputs(11555)) and (layer1_outputs(8388));
    layer2_outputs(2295) <= layer1_outputs(8128);
    layer2_outputs(2296) <= not(layer1_outputs(6853));
    layer2_outputs(2297) <= (layer1_outputs(3860)) or (layer1_outputs(3709));
    layer2_outputs(2298) <= layer1_outputs(12297);
    layer2_outputs(2299) <= not((layer1_outputs(1187)) and (layer1_outputs(2687)));
    layer2_outputs(2300) <= (layer1_outputs(9433)) or (layer1_outputs(10776));
    layer2_outputs(2301) <= (layer1_outputs(3215)) and (layer1_outputs(3377));
    layer2_outputs(2302) <= not(layer1_outputs(10491));
    layer2_outputs(2303) <= (layer1_outputs(4658)) or (layer1_outputs(1212));
    layer2_outputs(2304) <= not(layer1_outputs(564));
    layer2_outputs(2305) <= not(layer1_outputs(3409));
    layer2_outputs(2306) <= not((layer1_outputs(3453)) or (layer1_outputs(11322)));
    layer2_outputs(2307) <= (layer1_outputs(3507)) and not (layer1_outputs(2380));
    layer2_outputs(2308) <= not((layer1_outputs(4707)) xor (layer1_outputs(5019)));
    layer2_outputs(2309) <= layer1_outputs(1554);
    layer2_outputs(2310) <= not(layer1_outputs(7994));
    layer2_outputs(2311) <= not(layer1_outputs(7575));
    layer2_outputs(2312) <= not(layer1_outputs(184)) or (layer1_outputs(8406));
    layer2_outputs(2313) <= not((layer1_outputs(226)) and (layer1_outputs(2327)));
    layer2_outputs(2314) <= layer1_outputs(912);
    layer2_outputs(2315) <= not(layer1_outputs(1427));
    layer2_outputs(2316) <= layer1_outputs(10696);
    layer2_outputs(2317) <= (layer1_outputs(399)) or (layer1_outputs(9037));
    layer2_outputs(2318) <= not((layer1_outputs(10170)) xor (layer1_outputs(12789)));
    layer2_outputs(2319) <= not((layer1_outputs(9138)) and (layer1_outputs(398)));
    layer2_outputs(2320) <= layer1_outputs(11966);
    layer2_outputs(2321) <= layer1_outputs(5456);
    layer2_outputs(2322) <= '1';
    layer2_outputs(2323) <= (layer1_outputs(1596)) and not (layer1_outputs(10509));
    layer2_outputs(2324) <= (layer1_outputs(3766)) and (layer1_outputs(11061));
    layer2_outputs(2325) <= layer1_outputs(580);
    layer2_outputs(2326) <= (layer1_outputs(1502)) and (layer1_outputs(6565));
    layer2_outputs(2327) <= layer1_outputs(10884);
    layer2_outputs(2328) <= not(layer1_outputs(4761));
    layer2_outputs(2329) <= (layer1_outputs(3582)) and not (layer1_outputs(12149));
    layer2_outputs(2330) <= not(layer1_outputs(3534)) or (layer1_outputs(9551));
    layer2_outputs(2331) <= not(layer1_outputs(3532));
    layer2_outputs(2332) <= layer1_outputs(1659);
    layer2_outputs(2333) <= not(layer1_outputs(422));
    layer2_outputs(2334) <= layer1_outputs(10477);
    layer2_outputs(2335) <= (layer1_outputs(12735)) and not (layer1_outputs(9213));
    layer2_outputs(2336) <= not(layer1_outputs(2098));
    layer2_outputs(2337) <= (layer1_outputs(6055)) or (layer1_outputs(508));
    layer2_outputs(2338) <= not(layer1_outputs(10077));
    layer2_outputs(2339) <= not(layer1_outputs(11984)) or (layer1_outputs(8844));
    layer2_outputs(2340) <= (layer1_outputs(8344)) and (layer1_outputs(4375));
    layer2_outputs(2341) <= (layer1_outputs(7154)) and (layer1_outputs(5622));
    layer2_outputs(2342) <= not(layer1_outputs(8960)) or (layer1_outputs(4689));
    layer2_outputs(2343) <= (layer1_outputs(6296)) xor (layer1_outputs(6445));
    layer2_outputs(2344) <= not(layer1_outputs(1836));
    layer2_outputs(2345) <= not(layer1_outputs(11774));
    layer2_outputs(2346) <= not((layer1_outputs(12414)) or (layer1_outputs(12379)));
    layer2_outputs(2347) <= not(layer1_outputs(10033));
    layer2_outputs(2348) <= not((layer1_outputs(5795)) and (layer1_outputs(5156)));
    layer2_outputs(2349) <= layer1_outputs(1561);
    layer2_outputs(2350) <= not((layer1_outputs(9249)) and (layer1_outputs(675)));
    layer2_outputs(2351) <= layer1_outputs(5153);
    layer2_outputs(2352) <= layer1_outputs(4757);
    layer2_outputs(2353) <= (layer1_outputs(5450)) and (layer1_outputs(2762));
    layer2_outputs(2354) <= (layer1_outputs(824)) xor (layer1_outputs(6582));
    layer2_outputs(2355) <= layer1_outputs(9573);
    layer2_outputs(2356) <= layer1_outputs(9039);
    layer2_outputs(2357) <= not(layer1_outputs(2739)) or (layer1_outputs(1126));
    layer2_outputs(2358) <= not(layer1_outputs(3879)) or (layer1_outputs(5362));
    layer2_outputs(2359) <= layer1_outputs(7550);
    layer2_outputs(2360) <= (layer1_outputs(8018)) or (layer1_outputs(9190));
    layer2_outputs(2361) <= not(layer1_outputs(1170));
    layer2_outputs(2362) <= not((layer1_outputs(1129)) and (layer1_outputs(4726)));
    layer2_outputs(2363) <= not((layer1_outputs(5870)) or (layer1_outputs(5762)));
    layer2_outputs(2364) <= not((layer1_outputs(9476)) and (layer1_outputs(10944)));
    layer2_outputs(2365) <= layer1_outputs(1762);
    layer2_outputs(2366) <= layer1_outputs(7518);
    layer2_outputs(2367) <= layer1_outputs(11098);
    layer2_outputs(2368) <= (layer1_outputs(10684)) xor (layer1_outputs(11548));
    layer2_outputs(2369) <= '1';
    layer2_outputs(2370) <= not(layer1_outputs(839));
    layer2_outputs(2371) <= (layer1_outputs(12503)) or (layer1_outputs(9346));
    layer2_outputs(2372) <= not((layer1_outputs(389)) xor (layer1_outputs(9356)));
    layer2_outputs(2373) <= not(layer1_outputs(8956)) or (layer1_outputs(11414));
    layer2_outputs(2374) <= (layer1_outputs(5376)) xor (layer1_outputs(8543));
    layer2_outputs(2375) <= layer1_outputs(1869);
    layer2_outputs(2376) <= layer1_outputs(7089);
    layer2_outputs(2377) <= not((layer1_outputs(12159)) and (layer1_outputs(4298)));
    layer2_outputs(2378) <= (layer1_outputs(12641)) and not (layer1_outputs(4113));
    layer2_outputs(2379) <= layer1_outputs(1078);
    layer2_outputs(2380) <= layer1_outputs(12692);
    layer2_outputs(2381) <= not((layer1_outputs(174)) or (layer1_outputs(5178)));
    layer2_outputs(2382) <= (layer1_outputs(268)) xor (layer1_outputs(7595));
    layer2_outputs(2383) <= layer1_outputs(9874);
    layer2_outputs(2384) <= layer1_outputs(12320);
    layer2_outputs(2385) <= not(layer1_outputs(11753));
    layer2_outputs(2386) <= (layer1_outputs(10087)) xor (layer1_outputs(4558));
    layer2_outputs(2387) <= (layer1_outputs(3770)) and (layer1_outputs(11962));
    layer2_outputs(2388) <= (layer1_outputs(12029)) or (layer1_outputs(6730));
    layer2_outputs(2389) <= not((layer1_outputs(3806)) xor (layer1_outputs(2390)));
    layer2_outputs(2390) <= not(layer1_outputs(1603)) or (layer1_outputs(2822));
    layer2_outputs(2391) <= not((layer1_outputs(5048)) xor (layer1_outputs(8998)));
    layer2_outputs(2392) <= not(layer1_outputs(10881));
    layer2_outputs(2393) <= (layer1_outputs(6460)) and (layer1_outputs(5789));
    layer2_outputs(2394) <= layer1_outputs(6379);
    layer2_outputs(2395) <= not(layer1_outputs(8286)) or (layer1_outputs(10764));
    layer2_outputs(2396) <= not((layer1_outputs(3915)) xor (layer1_outputs(795)));
    layer2_outputs(2397) <= not((layer1_outputs(11354)) and (layer1_outputs(5599)));
    layer2_outputs(2398) <= (layer1_outputs(5280)) and (layer1_outputs(3539));
    layer2_outputs(2399) <= not(layer1_outputs(3863)) or (layer1_outputs(6742));
    layer2_outputs(2400) <= not((layer1_outputs(11808)) and (layer1_outputs(10927)));
    layer2_outputs(2401) <= not(layer1_outputs(2440));
    layer2_outputs(2402) <= not((layer1_outputs(6386)) or (layer1_outputs(9993)));
    layer2_outputs(2403) <= layer1_outputs(11866);
    layer2_outputs(2404) <= not(layer1_outputs(11907));
    layer2_outputs(2405) <= (layer1_outputs(7859)) and not (layer1_outputs(5878));
    layer2_outputs(2406) <= layer1_outputs(3219);
    layer2_outputs(2407) <= layer1_outputs(10899);
    layer2_outputs(2408) <= not(layer1_outputs(9689));
    layer2_outputs(2409) <= not((layer1_outputs(6506)) or (layer1_outputs(3876)));
    layer2_outputs(2410) <= layer1_outputs(12363);
    layer2_outputs(2411) <= layer1_outputs(788);
    layer2_outputs(2412) <= not((layer1_outputs(1170)) and (layer1_outputs(7224)));
    layer2_outputs(2413) <= (layer1_outputs(759)) or (layer1_outputs(6027));
    layer2_outputs(2414) <= not((layer1_outputs(188)) xor (layer1_outputs(3804)));
    layer2_outputs(2415) <= (layer1_outputs(4184)) or (layer1_outputs(9612));
    layer2_outputs(2416) <= layer1_outputs(11267);
    layer2_outputs(2417) <= not(layer1_outputs(2267));
    layer2_outputs(2418) <= layer1_outputs(1935);
    layer2_outputs(2419) <= not(layer1_outputs(2223));
    layer2_outputs(2420) <= not(layer1_outputs(2109));
    layer2_outputs(2421) <= layer1_outputs(3100);
    layer2_outputs(2422) <= not((layer1_outputs(6830)) xor (layer1_outputs(4018)));
    layer2_outputs(2423) <= not((layer1_outputs(10173)) xor (layer1_outputs(8140)));
    layer2_outputs(2424) <= not(layer1_outputs(596));
    layer2_outputs(2425) <= layer1_outputs(5504);
    layer2_outputs(2426) <= not(layer1_outputs(8551));
    layer2_outputs(2427) <= layer1_outputs(431);
    layer2_outputs(2428) <= not(layer1_outputs(8180));
    layer2_outputs(2429) <= layer1_outputs(11455);
    layer2_outputs(2430) <= not(layer1_outputs(11886)) or (layer1_outputs(7955));
    layer2_outputs(2431) <= not(layer1_outputs(8969));
    layer2_outputs(2432) <= not((layer1_outputs(12203)) xor (layer1_outputs(1197)));
    layer2_outputs(2433) <= not(layer1_outputs(8484));
    layer2_outputs(2434) <= (layer1_outputs(4897)) or (layer1_outputs(4623));
    layer2_outputs(2435) <= layer1_outputs(2631);
    layer2_outputs(2436) <= not(layer1_outputs(10772)) or (layer1_outputs(3339));
    layer2_outputs(2437) <= (layer1_outputs(6636)) xor (layer1_outputs(8794));
    layer2_outputs(2438) <= not(layer1_outputs(5191));
    layer2_outputs(2439) <= not(layer1_outputs(4149));
    layer2_outputs(2440) <= not(layer1_outputs(1850));
    layer2_outputs(2441) <= (layer1_outputs(2299)) and not (layer1_outputs(4446));
    layer2_outputs(2442) <= (layer1_outputs(1418)) xor (layer1_outputs(10682));
    layer2_outputs(2443) <= (layer1_outputs(7117)) and (layer1_outputs(1042));
    layer2_outputs(2444) <= (layer1_outputs(7306)) or (layer1_outputs(5081));
    layer2_outputs(2445) <= layer1_outputs(3515);
    layer2_outputs(2446) <= not(layer1_outputs(3903));
    layer2_outputs(2447) <= not(layer1_outputs(2312)) or (layer1_outputs(12108));
    layer2_outputs(2448) <= not((layer1_outputs(3837)) or (layer1_outputs(3477)));
    layer2_outputs(2449) <= (layer1_outputs(1912)) xor (layer1_outputs(11616));
    layer2_outputs(2450) <= layer1_outputs(11294);
    layer2_outputs(2451) <= (layer1_outputs(469)) and not (layer1_outputs(12174));
    layer2_outputs(2452) <= layer1_outputs(3616);
    layer2_outputs(2453) <= not(layer1_outputs(901));
    layer2_outputs(2454) <= not(layer1_outputs(2341));
    layer2_outputs(2455) <= not(layer1_outputs(7951)) or (layer1_outputs(3753));
    layer2_outputs(2456) <= (layer1_outputs(9662)) xor (layer1_outputs(3284));
    layer2_outputs(2457) <= not(layer1_outputs(3125));
    layer2_outputs(2458) <= (layer1_outputs(4078)) xor (layer1_outputs(508));
    layer2_outputs(2459) <= not(layer1_outputs(9428));
    layer2_outputs(2460) <= layer1_outputs(6523);
    layer2_outputs(2461) <= layer1_outputs(3153);
    layer2_outputs(2462) <= not(layer1_outputs(498));
    layer2_outputs(2463) <= (layer1_outputs(5582)) and not (layer1_outputs(6353));
    layer2_outputs(2464) <= not((layer1_outputs(5964)) or (layer1_outputs(10949)));
    layer2_outputs(2465) <= (layer1_outputs(2692)) and not (layer1_outputs(9006));
    layer2_outputs(2466) <= layer1_outputs(6608);
    layer2_outputs(2467) <= not(layer1_outputs(3461));
    layer2_outputs(2468) <= not(layer1_outputs(6371));
    layer2_outputs(2469) <= not(layer1_outputs(4913));
    layer2_outputs(2470) <= not((layer1_outputs(6122)) and (layer1_outputs(8091)));
    layer2_outputs(2471) <= not(layer1_outputs(9012)) or (layer1_outputs(6008));
    layer2_outputs(2472) <= not((layer1_outputs(10179)) and (layer1_outputs(6467)));
    layer2_outputs(2473) <= not(layer1_outputs(8396)) or (layer1_outputs(3358));
    layer2_outputs(2474) <= layer1_outputs(1592);
    layer2_outputs(2475) <= (layer1_outputs(12525)) and (layer1_outputs(5916));
    layer2_outputs(2476) <= layer1_outputs(2183);
    layer2_outputs(2477) <= (layer1_outputs(4060)) and (layer1_outputs(5480));
    layer2_outputs(2478) <= not((layer1_outputs(11960)) and (layer1_outputs(7172)));
    layer2_outputs(2479) <= not((layer1_outputs(4391)) xor (layer1_outputs(10661)));
    layer2_outputs(2480) <= (layer1_outputs(105)) and (layer1_outputs(2046));
    layer2_outputs(2481) <= not(layer1_outputs(2769));
    layer2_outputs(2482) <= not(layer1_outputs(6376));
    layer2_outputs(2483) <= layer1_outputs(5348);
    layer2_outputs(2484) <= not((layer1_outputs(2247)) and (layer1_outputs(123)));
    layer2_outputs(2485) <= layer1_outputs(3751);
    layer2_outputs(2486) <= (layer1_outputs(11591)) and (layer1_outputs(11623));
    layer2_outputs(2487) <= not(layer1_outputs(2455));
    layer2_outputs(2488) <= not((layer1_outputs(1520)) and (layer1_outputs(10741)));
    layer2_outputs(2489) <= layer1_outputs(2792);
    layer2_outputs(2490) <= not(layer1_outputs(8266)) or (layer1_outputs(56));
    layer2_outputs(2491) <= (layer1_outputs(5720)) or (layer1_outputs(9320));
    layer2_outputs(2492) <= (layer1_outputs(11777)) or (layer1_outputs(11814));
    layer2_outputs(2493) <= not(layer1_outputs(5340));
    layer2_outputs(2494) <= not((layer1_outputs(8359)) and (layer1_outputs(9565)));
    layer2_outputs(2495) <= not(layer1_outputs(3436));
    layer2_outputs(2496) <= layer1_outputs(2503);
    layer2_outputs(2497) <= not(layer1_outputs(3701));
    layer2_outputs(2498) <= not(layer1_outputs(12364));
    layer2_outputs(2499) <= not(layer1_outputs(5913));
    layer2_outputs(2500) <= not(layer1_outputs(4378));
    layer2_outputs(2501) <= not(layer1_outputs(8765)) or (layer1_outputs(72));
    layer2_outputs(2502) <= (layer1_outputs(12693)) or (layer1_outputs(8925));
    layer2_outputs(2503) <= (layer1_outputs(6679)) and not (layer1_outputs(1344));
    layer2_outputs(2504) <= (layer1_outputs(10259)) xor (layer1_outputs(3494));
    layer2_outputs(2505) <= (layer1_outputs(3677)) and (layer1_outputs(5411));
    layer2_outputs(2506) <= not(layer1_outputs(12130)) or (layer1_outputs(10504));
    layer2_outputs(2507) <= not(layer1_outputs(191));
    layer2_outputs(2508) <= (layer1_outputs(12070)) and (layer1_outputs(7146));
    layer2_outputs(2509) <= layer1_outputs(2171);
    layer2_outputs(2510) <= layer1_outputs(4902);
    layer2_outputs(2511) <= layer1_outputs(5467);
    layer2_outputs(2512) <= (layer1_outputs(3672)) xor (layer1_outputs(6431));
    layer2_outputs(2513) <= not(layer1_outputs(2536)) or (layer1_outputs(5892));
    layer2_outputs(2514) <= not(layer1_outputs(2828));
    layer2_outputs(2515) <= layer1_outputs(945);
    layer2_outputs(2516) <= not(layer1_outputs(11649));
    layer2_outputs(2517) <= layer1_outputs(6270);
    layer2_outputs(2518) <= (layer1_outputs(3853)) and not (layer1_outputs(9381));
    layer2_outputs(2519) <= not(layer1_outputs(8826)) or (layer1_outputs(3054));
    layer2_outputs(2520) <= not((layer1_outputs(1569)) xor (layer1_outputs(9913)));
    layer2_outputs(2521) <= not(layer1_outputs(5315)) or (layer1_outputs(12709));
    layer2_outputs(2522) <= not(layer1_outputs(7381)) or (layer1_outputs(9583));
    layer2_outputs(2523) <= layer1_outputs(10207);
    layer2_outputs(2524) <= layer1_outputs(10181);
    layer2_outputs(2525) <= not((layer1_outputs(3540)) xor (layer1_outputs(7191)));
    layer2_outputs(2526) <= not(layer1_outputs(5484));
    layer2_outputs(2527) <= layer1_outputs(7);
    layer2_outputs(2528) <= not((layer1_outputs(8669)) and (layer1_outputs(1063)));
    layer2_outputs(2529) <= layer1_outputs(9946);
    layer2_outputs(2530) <= not(layer1_outputs(8948));
    layer2_outputs(2531) <= not((layer1_outputs(6221)) and (layer1_outputs(6327)));
    layer2_outputs(2532) <= (layer1_outputs(3058)) and not (layer1_outputs(2037));
    layer2_outputs(2533) <= not(layer1_outputs(910));
    layer2_outputs(2534) <= (layer1_outputs(10284)) and not (layer1_outputs(4950));
    layer2_outputs(2535) <= layer1_outputs(12409);
    layer2_outputs(2536) <= not(layer1_outputs(8255)) or (layer1_outputs(11487));
    layer2_outputs(2537) <= (layer1_outputs(9307)) and (layer1_outputs(8539));
    layer2_outputs(2538) <= (layer1_outputs(11959)) or (layer1_outputs(8099));
    layer2_outputs(2539) <= layer1_outputs(6246);
    layer2_outputs(2540) <= not(layer1_outputs(7345));
    layer2_outputs(2541) <= layer1_outputs(7371);
    layer2_outputs(2542) <= (layer1_outputs(5763)) and (layer1_outputs(10615));
    layer2_outputs(2543) <= layer1_outputs(7228);
    layer2_outputs(2544) <= (layer1_outputs(1433)) or (layer1_outputs(10622));
    layer2_outputs(2545) <= not((layer1_outputs(2229)) xor (layer1_outputs(8096)));
    layer2_outputs(2546) <= not(layer1_outputs(12176)) or (layer1_outputs(10549));
    layer2_outputs(2547) <= (layer1_outputs(824)) xor (layer1_outputs(5702));
    layer2_outputs(2548) <= layer1_outputs(2912);
    layer2_outputs(2549) <= not((layer1_outputs(294)) xor (layer1_outputs(3425)));
    layer2_outputs(2550) <= not(layer1_outputs(6260)) or (layer1_outputs(3325));
    layer2_outputs(2551) <= (layer1_outputs(9790)) and (layer1_outputs(4813));
    layer2_outputs(2552) <= not(layer1_outputs(5322));
    layer2_outputs(2553) <= (layer1_outputs(11222)) xor (layer1_outputs(8796));
    layer2_outputs(2554) <= not(layer1_outputs(5893));
    layer2_outputs(2555) <= not(layer1_outputs(12144));
    layer2_outputs(2556) <= (layer1_outputs(7650)) and not (layer1_outputs(195));
    layer2_outputs(2557) <= not((layer1_outputs(1114)) xor (layer1_outputs(11728)));
    layer2_outputs(2558) <= not(layer1_outputs(10740));
    layer2_outputs(2559) <= '1';
    layer2_outputs(2560) <= (layer1_outputs(6555)) xor (layer1_outputs(82));
    layer2_outputs(2561) <= (layer1_outputs(2990)) and not (layer1_outputs(11648));
    layer2_outputs(2562) <= (layer1_outputs(4597)) or (layer1_outputs(12251));
    layer2_outputs(2563) <= not(layer1_outputs(8460));
    layer2_outputs(2564) <= layer1_outputs(12392);
    layer2_outputs(2565) <= layer1_outputs(12516);
    layer2_outputs(2566) <= (layer1_outputs(10647)) and not (layer1_outputs(7967));
    layer2_outputs(2567) <= (layer1_outputs(945)) or (layer1_outputs(8210));
    layer2_outputs(2568) <= (layer1_outputs(4636)) and not (layer1_outputs(9631));
    layer2_outputs(2569) <= not((layer1_outputs(7787)) or (layer1_outputs(8647)));
    layer2_outputs(2570) <= layer1_outputs(9490);
    layer2_outputs(2571) <= not(layer1_outputs(7409));
    layer2_outputs(2572) <= layer1_outputs(9613);
    layer2_outputs(2573) <= not(layer1_outputs(7682));
    layer2_outputs(2574) <= layer1_outputs(8543);
    layer2_outputs(2575) <= not(layer1_outputs(9919));
    layer2_outputs(2576) <= not((layer1_outputs(6356)) or (layer1_outputs(5106)));
    layer2_outputs(2577) <= layer1_outputs(10990);
    layer2_outputs(2578) <= (layer1_outputs(3604)) and not (layer1_outputs(4701));
    layer2_outputs(2579) <= not((layer1_outputs(11132)) and (layer1_outputs(6936)));
    layer2_outputs(2580) <= layer1_outputs(9804);
    layer2_outputs(2581) <= (layer1_outputs(2257)) and not (layer1_outputs(11368));
    layer2_outputs(2582) <= layer1_outputs(9261);
    layer2_outputs(2583) <= not((layer1_outputs(1152)) and (layer1_outputs(3176)));
    layer2_outputs(2584) <= (layer1_outputs(1116)) and not (layer1_outputs(656));
    layer2_outputs(2585) <= not(layer1_outputs(6642)) or (layer1_outputs(11961));
    layer2_outputs(2586) <= layer1_outputs(1994);
    layer2_outputs(2587) <= layer1_outputs(4328);
    layer2_outputs(2588) <= (layer1_outputs(10093)) and not (layer1_outputs(4204));
    layer2_outputs(2589) <= not((layer1_outputs(12172)) and (layer1_outputs(7086)));
    layer2_outputs(2590) <= not((layer1_outputs(8572)) and (layer1_outputs(9961)));
    layer2_outputs(2591) <= not((layer1_outputs(2587)) or (layer1_outputs(9023)));
    layer2_outputs(2592) <= layer1_outputs(11745);
    layer2_outputs(2593) <= (layer1_outputs(5837)) and (layer1_outputs(10214));
    layer2_outputs(2594) <= layer1_outputs(4792);
    layer2_outputs(2595) <= (layer1_outputs(11159)) xor (layer1_outputs(9499));
    layer2_outputs(2596) <= not(layer1_outputs(5391));
    layer2_outputs(2597) <= layer1_outputs(4556);
    layer2_outputs(2598) <= (layer1_outputs(9548)) and not (layer1_outputs(368));
    layer2_outputs(2599) <= (layer1_outputs(10096)) xor (layer1_outputs(3859));
    layer2_outputs(2600) <= not(layer1_outputs(12561)) or (layer1_outputs(10142));
    layer2_outputs(2601) <= layer1_outputs(8275);
    layer2_outputs(2602) <= not(layer1_outputs(1382));
    layer2_outputs(2603) <= not(layer1_outputs(117)) or (layer1_outputs(1233));
    layer2_outputs(2604) <= not(layer1_outputs(5137));
    layer2_outputs(2605) <= not((layer1_outputs(1300)) and (layer1_outputs(11343)));
    layer2_outputs(2606) <= not(layer1_outputs(11678));
    layer2_outputs(2607) <= layer1_outputs(10584);
    layer2_outputs(2608) <= layer1_outputs(7243);
    layer2_outputs(2609) <= (layer1_outputs(9938)) xor (layer1_outputs(2754));
    layer2_outputs(2610) <= not(layer1_outputs(10403)) or (layer1_outputs(9680));
    layer2_outputs(2611) <= not(layer1_outputs(2281)) or (layer1_outputs(3303));
    layer2_outputs(2612) <= layer1_outputs(12077);
    layer2_outputs(2613) <= not(layer1_outputs(8082));
    layer2_outputs(2614) <= not(layer1_outputs(9109));
    layer2_outputs(2615) <= not(layer1_outputs(12404)) or (layer1_outputs(9062));
    layer2_outputs(2616) <= not((layer1_outputs(748)) or (layer1_outputs(3746)));
    layer2_outputs(2617) <= layer1_outputs(11322);
    layer2_outputs(2618) <= layer1_outputs(4368);
    layer2_outputs(2619) <= (layer1_outputs(7073)) xor (layer1_outputs(4824));
    layer2_outputs(2620) <= (layer1_outputs(11452)) and not (layer1_outputs(10790));
    layer2_outputs(2621) <= layer1_outputs(7203);
    layer2_outputs(2622) <= (layer1_outputs(1766)) xor (layer1_outputs(12432));
    layer2_outputs(2623) <= not(layer1_outputs(12336));
    layer2_outputs(2624) <= not(layer1_outputs(2723));
    layer2_outputs(2625) <= not(layer1_outputs(8517));
    layer2_outputs(2626) <= not(layer1_outputs(6457));
    layer2_outputs(2627) <= not(layer1_outputs(1090));
    layer2_outputs(2628) <= not((layer1_outputs(2216)) or (layer1_outputs(69)));
    layer2_outputs(2629) <= not(layer1_outputs(32));
    layer2_outputs(2630) <= (layer1_outputs(9045)) or (layer1_outputs(4486));
    layer2_outputs(2631) <= not(layer1_outputs(6382));
    layer2_outputs(2632) <= layer1_outputs(1588);
    layer2_outputs(2633) <= (layer1_outputs(6533)) and not (layer1_outputs(11449));
    layer2_outputs(2634) <= layer1_outputs(214);
    layer2_outputs(2635) <= not(layer1_outputs(9590)) or (layer1_outputs(7460));
    layer2_outputs(2636) <= not(layer1_outputs(12032));
    layer2_outputs(2637) <= layer1_outputs(5900);
    layer2_outputs(2638) <= (layer1_outputs(693)) or (layer1_outputs(11168));
    layer2_outputs(2639) <= not((layer1_outputs(2989)) xor (layer1_outputs(4612)));
    layer2_outputs(2640) <= layer1_outputs(1541);
    layer2_outputs(2641) <= (layer1_outputs(7498)) xor (layer1_outputs(12329));
    layer2_outputs(2642) <= layer1_outputs(3916);
    layer2_outputs(2643) <= not((layer1_outputs(5415)) xor (layer1_outputs(10569)));
    layer2_outputs(2644) <= (layer1_outputs(6867)) and (layer1_outputs(4020));
    layer2_outputs(2645) <= not((layer1_outputs(11012)) or (layer1_outputs(7121)));
    layer2_outputs(2646) <= (layer1_outputs(6516)) and not (layer1_outputs(5095));
    layer2_outputs(2647) <= layer1_outputs(10279);
    layer2_outputs(2648) <= not(layer1_outputs(11784)) or (layer1_outputs(6743));
    layer2_outputs(2649) <= not(layer1_outputs(2950)) or (layer1_outputs(3654));
    layer2_outputs(2650) <= (layer1_outputs(1261)) xor (layer1_outputs(7359));
    layer2_outputs(2651) <= (layer1_outputs(2570)) and not (layer1_outputs(11697));
    layer2_outputs(2652) <= not(layer1_outputs(6099));
    layer2_outputs(2653) <= not(layer1_outputs(11500)) or (layer1_outputs(5236));
    layer2_outputs(2654) <= not((layer1_outputs(3712)) or (layer1_outputs(1247)));
    layer2_outputs(2655) <= not(layer1_outputs(8333));
    layer2_outputs(2656) <= not(layer1_outputs(6191)) or (layer1_outputs(8369));
    layer2_outputs(2657) <= (layer1_outputs(502)) and not (layer1_outputs(2331));
    layer2_outputs(2658) <= not((layer1_outputs(4140)) xor (layer1_outputs(7786)));
    layer2_outputs(2659) <= not(layer1_outputs(304));
    layer2_outputs(2660) <= not(layer1_outputs(1477));
    layer2_outputs(2661) <= not(layer1_outputs(1694));
    layer2_outputs(2662) <= not(layer1_outputs(1924));
    layer2_outputs(2663) <= not(layer1_outputs(1713));
    layer2_outputs(2664) <= layer1_outputs(1946);
    layer2_outputs(2665) <= not(layer1_outputs(8878));
    layer2_outputs(2666) <= layer1_outputs(397);
    layer2_outputs(2667) <= (layer1_outputs(11755)) and not (layer1_outputs(5535));
    layer2_outputs(2668) <= not(layer1_outputs(1018));
    layer2_outputs(2669) <= not(layer1_outputs(6428));
    layer2_outputs(2670) <= not((layer1_outputs(9975)) xor (layer1_outputs(12243)));
    layer2_outputs(2671) <= (layer1_outputs(2112)) or (layer1_outputs(6135));
    layer2_outputs(2672) <= not((layer1_outputs(5399)) xor (layer1_outputs(420)));
    layer2_outputs(2673) <= (layer1_outputs(9879)) and (layer1_outputs(9978));
    layer2_outputs(2674) <= layer1_outputs(8938);
    layer2_outputs(2675) <= layer1_outputs(505);
    layer2_outputs(2676) <= layer1_outputs(1845);
    layer2_outputs(2677) <= layer1_outputs(8271);
    layer2_outputs(2678) <= not((layer1_outputs(6362)) or (layer1_outputs(602)));
    layer2_outputs(2679) <= not(layer1_outputs(12173)) or (layer1_outputs(5486));
    layer2_outputs(2680) <= (layer1_outputs(4442)) or (layer1_outputs(9672));
    layer2_outputs(2681) <= not(layer1_outputs(3729));
    layer2_outputs(2682) <= not(layer1_outputs(1389));
    layer2_outputs(2683) <= (layer1_outputs(10519)) and not (layer1_outputs(8105));
    layer2_outputs(2684) <= not(layer1_outputs(3287));
    layer2_outputs(2685) <= (layer1_outputs(2372)) and not (layer1_outputs(10250));
    layer2_outputs(2686) <= (layer1_outputs(7651)) and (layer1_outputs(8728));
    layer2_outputs(2687) <= layer1_outputs(8839);
    layer2_outputs(2688) <= (layer1_outputs(10971)) and not (layer1_outputs(12284));
    layer2_outputs(2689) <= not((layer1_outputs(4898)) xor (layer1_outputs(3904)));
    layer2_outputs(2690) <= not(layer1_outputs(1439));
    layer2_outputs(2691) <= (layer1_outputs(12704)) xor (layer1_outputs(9581));
    layer2_outputs(2692) <= (layer1_outputs(4937)) or (layer1_outputs(2389));
    layer2_outputs(2693) <= (layer1_outputs(8023)) and not (layer1_outputs(2801));
    layer2_outputs(2694) <= not(layer1_outputs(10691));
    layer2_outputs(2695) <= not(layer1_outputs(1999));
    layer2_outputs(2696) <= not((layer1_outputs(9690)) xor (layer1_outputs(9276)));
    layer2_outputs(2697) <= layer1_outputs(4567);
    layer2_outputs(2698) <= not((layer1_outputs(1735)) and (layer1_outputs(4010)));
    layer2_outputs(2699) <= not((layer1_outputs(10384)) or (layer1_outputs(10448)));
    layer2_outputs(2700) <= not(layer1_outputs(1802));
    layer2_outputs(2701) <= (layer1_outputs(11249)) or (layer1_outputs(3184));
    layer2_outputs(2702) <= layer1_outputs(2888);
    layer2_outputs(2703) <= layer1_outputs(8334);
    layer2_outputs(2704) <= (layer1_outputs(11994)) xor (layer1_outputs(1254));
    layer2_outputs(2705) <= not(layer1_outputs(11844));
    layer2_outputs(2706) <= not((layer1_outputs(2651)) and (layer1_outputs(9060)));
    layer2_outputs(2707) <= not(layer1_outputs(7746));
    layer2_outputs(2708) <= not(layer1_outputs(6113));
    layer2_outputs(2709) <= layer1_outputs(2266);
    layer2_outputs(2710) <= not((layer1_outputs(7296)) xor (layer1_outputs(7913)));
    layer2_outputs(2711) <= (layer1_outputs(7077)) and not (layer1_outputs(11631));
    layer2_outputs(2712) <= not(layer1_outputs(8067));
    layer2_outputs(2713) <= not((layer1_outputs(661)) xor (layer1_outputs(9413)));
    layer2_outputs(2714) <= (layer1_outputs(1892)) and (layer1_outputs(12184));
    layer2_outputs(2715) <= layer1_outputs(3560);
    layer2_outputs(2716) <= layer1_outputs(10769);
    layer2_outputs(2717) <= not((layer1_outputs(4686)) xor (layer1_outputs(10171)));
    layer2_outputs(2718) <= (layer1_outputs(10710)) xor (layer1_outputs(7517));
    layer2_outputs(2719) <= not(layer1_outputs(4082));
    layer2_outputs(2720) <= (layer1_outputs(7504)) and not (layer1_outputs(2793));
    layer2_outputs(2721) <= not(layer1_outputs(9492));
    layer2_outputs(2722) <= (layer1_outputs(10435)) and (layer1_outputs(10079));
    layer2_outputs(2723) <= layer1_outputs(11156);
    layer2_outputs(2724) <= not((layer1_outputs(10483)) and (layer1_outputs(10697)));
    layer2_outputs(2725) <= (layer1_outputs(3637)) and not (layer1_outputs(1500));
    layer2_outputs(2726) <= not(layer1_outputs(7736));
    layer2_outputs(2727) <= not(layer1_outputs(243)) or (layer1_outputs(6940));
    layer2_outputs(2728) <= not(layer1_outputs(12040));
    layer2_outputs(2729) <= not(layer1_outputs(5979)) or (layer1_outputs(8863));
    layer2_outputs(2730) <= (layer1_outputs(12656)) and not (layer1_outputs(7699));
    layer2_outputs(2731) <= (layer1_outputs(10959)) xor (layer1_outputs(10274));
    layer2_outputs(2732) <= layer1_outputs(7173);
    layer2_outputs(2733) <= layer1_outputs(10937);
    layer2_outputs(2734) <= not((layer1_outputs(6057)) or (layer1_outputs(12321)));
    layer2_outputs(2735) <= layer1_outputs(3444);
    layer2_outputs(2736) <= layer1_outputs(7369);
    layer2_outputs(2737) <= layer1_outputs(8393);
    layer2_outputs(2738) <= not(layer1_outputs(12190));
    layer2_outputs(2739) <= (layer1_outputs(11319)) and (layer1_outputs(7149));
    layer2_outputs(2740) <= not((layer1_outputs(8115)) or (layer1_outputs(408)));
    layer2_outputs(2741) <= layer1_outputs(2025);
    layer2_outputs(2742) <= layer1_outputs(3520);
    layer2_outputs(2743) <= layer1_outputs(6435);
    layer2_outputs(2744) <= '1';
    layer2_outputs(2745) <= layer1_outputs(12512);
    layer2_outputs(2746) <= not(layer1_outputs(1369));
    layer2_outputs(2747) <= layer1_outputs(2972);
    layer2_outputs(2748) <= not(layer1_outputs(3293));
    layer2_outputs(2749) <= (layer1_outputs(6745)) and not (layer1_outputs(5465));
    layer2_outputs(2750) <= layer1_outputs(6323);
    layer2_outputs(2751) <= (layer1_outputs(8064)) xor (layer1_outputs(1135));
    layer2_outputs(2752) <= layer1_outputs(7070);
    layer2_outputs(2753) <= not((layer1_outputs(3912)) and (layer1_outputs(4858)));
    layer2_outputs(2754) <= layer1_outputs(9045);
    layer2_outputs(2755) <= layer1_outputs(5547);
    layer2_outputs(2756) <= not((layer1_outputs(60)) and (layer1_outputs(274)));
    layer2_outputs(2757) <= layer1_outputs(6220);
    layer2_outputs(2758) <= not(layer1_outputs(10914)) or (layer1_outputs(2854));
    layer2_outputs(2759) <= layer1_outputs(2601);
    layer2_outputs(2760) <= (layer1_outputs(7857)) and not (layer1_outputs(10896));
    layer2_outputs(2761) <= not(layer1_outputs(1590)) or (layer1_outputs(6476));
    layer2_outputs(2762) <= not(layer1_outputs(4240)) or (layer1_outputs(674));
    layer2_outputs(2763) <= not(layer1_outputs(10535));
    layer2_outputs(2764) <= not(layer1_outputs(11600)) or (layer1_outputs(1979));
    layer2_outputs(2765) <= '0';
    layer2_outputs(2766) <= layer1_outputs(10892);
    layer2_outputs(2767) <= not((layer1_outputs(7861)) and (layer1_outputs(5157)));
    layer2_outputs(2768) <= layer1_outputs(3595);
    layer2_outputs(2769) <= not(layer1_outputs(10928));
    layer2_outputs(2770) <= not(layer1_outputs(8691)) or (layer1_outputs(1529));
    layer2_outputs(2771) <= layer1_outputs(2825);
    layer2_outputs(2772) <= not((layer1_outputs(2478)) xor (layer1_outputs(9891)));
    layer2_outputs(2773) <= not(layer1_outputs(289));
    layer2_outputs(2774) <= (layer1_outputs(1552)) and not (layer1_outputs(66));
    layer2_outputs(2775) <= not(layer1_outputs(8044)) or (layer1_outputs(9682));
    layer2_outputs(2776) <= layer1_outputs(8298);
    layer2_outputs(2777) <= not(layer1_outputs(11408));
    layer2_outputs(2778) <= layer1_outputs(12466);
    layer2_outputs(2779) <= (layer1_outputs(11045)) or (layer1_outputs(3732));
    layer2_outputs(2780) <= (layer1_outputs(2523)) xor (layer1_outputs(1524));
    layer2_outputs(2781) <= not(layer1_outputs(2054));
    layer2_outputs(2782) <= layer1_outputs(9726);
    layer2_outputs(2783) <= not((layer1_outputs(11738)) xor (layer1_outputs(8296)));
    layer2_outputs(2784) <= not((layer1_outputs(11085)) xor (layer1_outputs(3623)));
    layer2_outputs(2785) <= not(layer1_outputs(353));
    layer2_outputs(2786) <= not(layer1_outputs(9209)) or (layer1_outputs(707));
    layer2_outputs(2787) <= not((layer1_outputs(9533)) or (layer1_outputs(9011)));
    layer2_outputs(2788) <= (layer1_outputs(9401)) or (layer1_outputs(1972));
    layer2_outputs(2789) <= layer1_outputs(3895);
    layer2_outputs(2790) <= not((layer1_outputs(9296)) xor (layer1_outputs(2670)));
    layer2_outputs(2791) <= not((layer1_outputs(1984)) xor (layer1_outputs(5398)));
    layer2_outputs(2792) <= (layer1_outputs(11298)) and (layer1_outputs(12620));
    layer2_outputs(2793) <= not((layer1_outputs(3841)) and (layer1_outputs(9800)));
    layer2_outputs(2794) <= not(layer1_outputs(4841));
    layer2_outputs(2795) <= layer1_outputs(8613);
    layer2_outputs(2796) <= not(layer1_outputs(8975));
    layer2_outputs(2797) <= not(layer1_outputs(105));
    layer2_outputs(2798) <= (layer1_outputs(4296)) or (layer1_outputs(11926));
    layer2_outputs(2799) <= (layer1_outputs(8439)) and not (layer1_outputs(9009));
    layer2_outputs(2800) <= layer1_outputs(4512);
    layer2_outputs(2801) <= layer1_outputs(1653);
    layer2_outputs(2802) <= not((layer1_outputs(5305)) and (layer1_outputs(11578)));
    layer2_outputs(2803) <= (layer1_outputs(1995)) xor (layer1_outputs(10664));
    layer2_outputs(2804) <= layer1_outputs(8813);
    layer2_outputs(2805) <= (layer1_outputs(317)) and not (layer1_outputs(9726));
    layer2_outputs(2806) <= not(layer1_outputs(9631)) or (layer1_outputs(10904));
    layer2_outputs(2807) <= not(layer1_outputs(8775));
    layer2_outputs(2808) <= not(layer1_outputs(5166));
    layer2_outputs(2809) <= layer1_outputs(7523);
    layer2_outputs(2810) <= layer1_outputs(9351);
    layer2_outputs(2811) <= (layer1_outputs(3430)) and not (layer1_outputs(8280));
    layer2_outputs(2812) <= not(layer1_outputs(3609)) or (layer1_outputs(10003));
    layer2_outputs(2813) <= (layer1_outputs(8947)) and (layer1_outputs(9901));
    layer2_outputs(2814) <= not(layer1_outputs(5068));
    layer2_outputs(2815) <= not(layer1_outputs(6888));
    layer2_outputs(2816) <= (layer1_outputs(11357)) or (layer1_outputs(8222));
    layer2_outputs(2817) <= (layer1_outputs(6847)) xor (layer1_outputs(6389));
    layer2_outputs(2818) <= not((layer1_outputs(2803)) or (layer1_outputs(10184)));
    layer2_outputs(2819) <= layer1_outputs(3613);
    layer2_outputs(2820) <= not((layer1_outputs(3204)) and (layer1_outputs(8874)));
    layer2_outputs(2821) <= layer1_outputs(1662);
    layer2_outputs(2822) <= layer1_outputs(3028);
    layer2_outputs(2823) <= not(layer1_outputs(1015));
    layer2_outputs(2824) <= not(layer1_outputs(341));
    layer2_outputs(2825) <= (layer1_outputs(3967)) and not (layer1_outputs(967));
    layer2_outputs(2826) <= (layer1_outputs(11145)) and not (layer1_outputs(4426));
    layer2_outputs(2827) <= not((layer1_outputs(1205)) xor (layer1_outputs(1881)));
    layer2_outputs(2828) <= layer1_outputs(5910);
    layer2_outputs(2829) <= not(layer1_outputs(10572));
    layer2_outputs(2830) <= not((layer1_outputs(181)) xor (layer1_outputs(11635)));
    layer2_outputs(2831) <= layer1_outputs(4047);
    layer2_outputs(2832) <= not(layer1_outputs(1673));
    layer2_outputs(2833) <= not((layer1_outputs(8899)) and (layer1_outputs(6767)));
    layer2_outputs(2834) <= not((layer1_outputs(8326)) xor (layer1_outputs(10130)));
    layer2_outputs(2835) <= layer1_outputs(4748);
    layer2_outputs(2836) <= (layer1_outputs(8552)) and (layer1_outputs(9663));
    layer2_outputs(2837) <= (layer1_outputs(7605)) and not (layer1_outputs(3138));
    layer2_outputs(2838) <= layer1_outputs(8149);
    layer2_outputs(2839) <= not((layer1_outputs(9252)) and (layer1_outputs(9308)));
    layer2_outputs(2840) <= layer1_outputs(5539);
    layer2_outputs(2841) <= layer1_outputs(5440);
    layer2_outputs(2842) <= not(layer1_outputs(11358));
    layer2_outputs(2843) <= layer1_outputs(3182);
    layer2_outputs(2844) <= not(layer1_outputs(10190));
    layer2_outputs(2845) <= (layer1_outputs(1489)) and not (layer1_outputs(8430));
    layer2_outputs(2846) <= not(layer1_outputs(2808));
    layer2_outputs(2847) <= not(layer1_outputs(4445));
    layer2_outputs(2848) <= (layer1_outputs(4402)) and not (layer1_outputs(7210));
    layer2_outputs(2849) <= layer1_outputs(1191);
    layer2_outputs(2850) <= not((layer1_outputs(6487)) xor (layer1_outputs(12205)));
    layer2_outputs(2851) <= layer1_outputs(12589);
    layer2_outputs(2852) <= not(layer1_outputs(381)) or (layer1_outputs(6688));
    layer2_outputs(2853) <= layer1_outputs(11079);
    layer2_outputs(2854) <= layer1_outputs(11394);
    layer2_outputs(2855) <= not(layer1_outputs(1623)) or (layer1_outputs(779));
    layer2_outputs(2856) <= not((layer1_outputs(10939)) or (layer1_outputs(8212)));
    layer2_outputs(2857) <= '0';
    layer2_outputs(2858) <= not(layer1_outputs(1010));
    layer2_outputs(2859) <= not(layer1_outputs(3796));
    layer2_outputs(2860) <= not((layer1_outputs(12318)) or (layer1_outputs(12289)));
    layer2_outputs(2861) <= not(layer1_outputs(2233)) or (layer1_outputs(1760));
    layer2_outputs(2862) <= layer1_outputs(12663);
    layer2_outputs(2863) <= layer1_outputs(6066);
    layer2_outputs(2864) <= layer1_outputs(11371);
    layer2_outputs(2865) <= layer1_outputs(7055);
    layer2_outputs(2866) <= not(layer1_outputs(507));
    layer2_outputs(2867) <= layer1_outputs(1030);
    layer2_outputs(2868) <= not(layer1_outputs(9462)) or (layer1_outputs(11827));
    layer2_outputs(2869) <= not(layer1_outputs(1705)) or (layer1_outputs(2283));
    layer2_outputs(2870) <= not(layer1_outputs(11139)) or (layer1_outputs(2994));
    layer2_outputs(2871) <= not(layer1_outputs(756));
    layer2_outputs(2872) <= not(layer1_outputs(11328)) or (layer1_outputs(1681));
    layer2_outputs(2873) <= not(layer1_outputs(3379));
    layer2_outputs(2874) <= layer1_outputs(1101);
    layer2_outputs(2875) <= layer1_outputs(4183);
    layer2_outputs(2876) <= layer1_outputs(5154);
    layer2_outputs(2877) <= layer1_outputs(3544);
    layer2_outputs(2878) <= layer1_outputs(9097);
    layer2_outputs(2879) <= not(layer1_outputs(5705));
    layer2_outputs(2880) <= not(layer1_outputs(7676));
    layer2_outputs(2881) <= layer1_outputs(5855);
    layer2_outputs(2882) <= (layer1_outputs(10623)) xor (layer1_outputs(4239));
    layer2_outputs(2883) <= not(layer1_outputs(2015));
    layer2_outputs(2884) <= (layer1_outputs(1203)) and not (layer1_outputs(4812));
    layer2_outputs(2885) <= (layer1_outputs(9774)) or (layer1_outputs(6000));
    layer2_outputs(2886) <= not(layer1_outputs(10234));
    layer2_outputs(2887) <= not(layer1_outputs(12008));
    layer2_outputs(2888) <= layer1_outputs(6697);
    layer2_outputs(2889) <= not(layer1_outputs(5634));
    layer2_outputs(2890) <= (layer1_outputs(8724)) or (layer1_outputs(1405));
    layer2_outputs(2891) <= layer1_outputs(2501);
    layer2_outputs(2892) <= (layer1_outputs(3803)) xor (layer1_outputs(4182));
    layer2_outputs(2893) <= (layer1_outputs(2270)) and not (layer1_outputs(12033));
    layer2_outputs(2894) <= layer1_outputs(10449);
    layer2_outputs(2895) <= not(layer1_outputs(6655));
    layer2_outputs(2896) <= layer1_outputs(3870);
    layer2_outputs(2897) <= not((layer1_outputs(238)) or (layer1_outputs(6685)));
    layer2_outputs(2898) <= not(layer1_outputs(12328));
    layer2_outputs(2899) <= (layer1_outputs(3423)) or (layer1_outputs(5925));
    layer2_outputs(2900) <= (layer1_outputs(6615)) or (layer1_outputs(7984));
    layer2_outputs(2901) <= '1';
    layer2_outputs(2902) <= (layer1_outputs(5769)) xor (layer1_outputs(6920));
    layer2_outputs(2903) <= not(layer1_outputs(5996));
    layer2_outputs(2904) <= not((layer1_outputs(7315)) xor (layer1_outputs(11128)));
    layer2_outputs(2905) <= layer1_outputs(1786);
    layer2_outputs(2906) <= layer1_outputs(12147);
    layer2_outputs(2907) <= not(layer1_outputs(10002));
    layer2_outputs(2908) <= (layer1_outputs(5214)) and not (layer1_outputs(3965));
    layer2_outputs(2909) <= (layer1_outputs(3511)) and not (layer1_outputs(9645));
    layer2_outputs(2910) <= (layer1_outputs(2629)) xor (layer1_outputs(9062));
    layer2_outputs(2911) <= layer1_outputs(3579);
    layer2_outputs(2912) <= (layer1_outputs(3807)) or (layer1_outputs(3165));
    layer2_outputs(2913) <= not(layer1_outputs(2213)) or (layer1_outputs(12456));
    layer2_outputs(2914) <= (layer1_outputs(5343)) xor (layer1_outputs(2997));
    layer2_outputs(2915) <= layer1_outputs(9531);
    layer2_outputs(2916) <= not(layer1_outputs(3890));
    layer2_outputs(2917) <= layer1_outputs(11205);
    layer2_outputs(2918) <= (layer1_outputs(6453)) and (layer1_outputs(1434));
    layer2_outputs(2919) <= not((layer1_outputs(5176)) xor (layer1_outputs(3610)));
    layer2_outputs(2920) <= not(layer1_outputs(4162));
    layer2_outputs(2921) <= layer1_outputs(303);
    layer2_outputs(2922) <= not((layer1_outputs(6802)) or (layer1_outputs(6304)));
    layer2_outputs(2923) <= (layer1_outputs(2147)) or (layer1_outputs(23));
    layer2_outputs(2924) <= not((layer1_outputs(2714)) or (layer1_outputs(2196)));
    layer2_outputs(2925) <= (layer1_outputs(5375)) or (layer1_outputs(7883));
    layer2_outputs(2926) <= layer1_outputs(9300);
    layer2_outputs(2927) <= not(layer1_outputs(2193)) or (layer1_outputs(5160));
    layer2_outputs(2928) <= not(layer1_outputs(11105));
    layer2_outputs(2929) <= layer1_outputs(12156);
    layer2_outputs(2930) <= not((layer1_outputs(10735)) xor (layer1_outputs(4160)));
    layer2_outputs(2931) <= layer1_outputs(5300);
    layer2_outputs(2932) <= layer1_outputs(11880);
    layer2_outputs(2933) <= (layer1_outputs(2944)) or (layer1_outputs(7289));
    layer2_outputs(2934) <= not(layer1_outputs(9638));
    layer2_outputs(2935) <= not(layer1_outputs(9817));
    layer2_outputs(2936) <= not(layer1_outputs(2863));
    layer2_outputs(2937) <= layer1_outputs(7036);
    layer2_outputs(2938) <= not((layer1_outputs(7286)) and (layer1_outputs(9640)));
    layer2_outputs(2939) <= layer1_outputs(6582);
    layer2_outputs(2940) <= (layer1_outputs(6079)) or (layer1_outputs(1395));
    layer2_outputs(2941) <= not((layer1_outputs(10892)) xor (layer1_outputs(716)));
    layer2_outputs(2942) <= not(layer1_outputs(3756));
    layer2_outputs(2943) <= layer1_outputs(2443);
    layer2_outputs(2944) <= (layer1_outputs(8823)) xor (layer1_outputs(7538));
    layer2_outputs(2945) <= layer1_outputs(8374);
    layer2_outputs(2946) <= not(layer1_outputs(9925));
    layer2_outputs(2947) <= layer1_outputs(7972);
    layer2_outputs(2948) <= layer1_outputs(5497);
    layer2_outputs(2949) <= (layer1_outputs(4910)) or (layer1_outputs(2644));
    layer2_outputs(2950) <= not(layer1_outputs(10142));
    layer2_outputs(2951) <= not(layer1_outputs(11219)) or (layer1_outputs(943));
    layer2_outputs(2952) <= not((layer1_outputs(10083)) or (layer1_outputs(7647)));
    layer2_outputs(2953) <= layer1_outputs(8653);
    layer2_outputs(2954) <= not(layer1_outputs(5591));
    layer2_outputs(2955) <= (layer1_outputs(6507)) xor (layer1_outputs(5372));
    layer2_outputs(2956) <= not((layer1_outputs(6985)) or (layer1_outputs(5076)));
    layer2_outputs(2957) <= not(layer1_outputs(4029)) or (layer1_outputs(11540));
    layer2_outputs(2958) <= '0';
    layer2_outputs(2959) <= not((layer1_outputs(4348)) xor (layer1_outputs(867)));
    layer2_outputs(2960) <= layer1_outputs(5727);
    layer2_outputs(2961) <= not(layer1_outputs(7046)) or (layer1_outputs(7807));
    layer2_outputs(2962) <= layer1_outputs(6696);
    layer2_outputs(2963) <= (layer1_outputs(9885)) or (layer1_outputs(11426));
    layer2_outputs(2964) <= (layer1_outputs(12192)) and not (layer1_outputs(11510));
    layer2_outputs(2965) <= (layer1_outputs(12382)) and (layer1_outputs(5823));
    layer2_outputs(2966) <= layer1_outputs(11696);
    layer2_outputs(2967) <= not(layer1_outputs(9535));
    layer2_outputs(2968) <= not(layer1_outputs(7804)) or (layer1_outputs(11187));
    layer2_outputs(2969) <= layer1_outputs(11640);
    layer2_outputs(2970) <= (layer1_outputs(4320)) or (layer1_outputs(1867));
    layer2_outputs(2971) <= layer1_outputs(2072);
    layer2_outputs(2972) <= not((layer1_outputs(4424)) and (layer1_outputs(6493)));
    layer2_outputs(2973) <= layer1_outputs(2167);
    layer2_outputs(2974) <= layer1_outputs(8090);
    layer2_outputs(2975) <= not(layer1_outputs(9199)) or (layer1_outputs(4841));
    layer2_outputs(2976) <= not((layer1_outputs(4560)) or (layer1_outputs(10781)));
    layer2_outputs(2977) <= not(layer1_outputs(5687)) or (layer1_outputs(5879));
    layer2_outputs(2978) <= not(layer1_outputs(2886));
    layer2_outputs(2979) <= layer1_outputs(4040);
    layer2_outputs(2980) <= not((layer1_outputs(2422)) xor (layer1_outputs(1818)));
    layer2_outputs(2981) <= not((layer1_outputs(9882)) or (layer1_outputs(3460)));
    layer2_outputs(2982) <= layer1_outputs(1597);
    layer2_outputs(2983) <= (layer1_outputs(2024)) and not (layer1_outputs(8016));
    layer2_outputs(2984) <= (layer1_outputs(3767)) and not (layer1_outputs(10624));
    layer2_outputs(2985) <= (layer1_outputs(7110)) or (layer1_outputs(662));
    layer2_outputs(2986) <= not(layer1_outputs(11822));
    layer2_outputs(2987) <= (layer1_outputs(4581)) xor (layer1_outputs(3331));
    layer2_outputs(2988) <= not(layer1_outputs(6689));
    layer2_outputs(2989) <= (layer1_outputs(2334)) and not (layer1_outputs(10113));
    layer2_outputs(2990) <= not(layer1_outputs(8245));
    layer2_outputs(2991) <= layer1_outputs(7520);
    layer2_outputs(2992) <= not(layer1_outputs(10455)) or (layer1_outputs(4618));
    layer2_outputs(2993) <= not(layer1_outputs(8973)) or (layer1_outputs(6211));
    layer2_outputs(2994) <= not(layer1_outputs(732));
    layer2_outputs(2995) <= not(layer1_outputs(4419));
    layer2_outputs(2996) <= not(layer1_outputs(7136));
    layer2_outputs(2997) <= layer1_outputs(4778);
    layer2_outputs(2998) <= (layer1_outputs(10593)) xor (layer1_outputs(4554));
    layer2_outputs(2999) <= not(layer1_outputs(5128));
    layer2_outputs(3000) <= not((layer1_outputs(6682)) xor (layer1_outputs(6887)));
    layer2_outputs(3001) <= not(layer1_outputs(6311));
    layer2_outputs(3002) <= not((layer1_outputs(11230)) or (layer1_outputs(6930)));
    layer2_outputs(3003) <= (layer1_outputs(10426)) and not (layer1_outputs(3354));
    layer2_outputs(3004) <= not((layer1_outputs(3561)) and (layer1_outputs(11939)));
    layer2_outputs(3005) <= not(layer1_outputs(3936));
    layer2_outputs(3006) <= (layer1_outputs(8864)) xor (layer1_outputs(733));
    layer2_outputs(3007) <= (layer1_outputs(2456)) or (layer1_outputs(11994));
    layer2_outputs(3008) <= not(layer1_outputs(11149));
    layer2_outputs(3009) <= not(layer1_outputs(10178));
    layer2_outputs(3010) <= not((layer1_outputs(3029)) and (layer1_outputs(11278)));
    layer2_outputs(3011) <= not(layer1_outputs(9870)) or (layer1_outputs(3725));
    layer2_outputs(3012) <= not((layer1_outputs(4298)) and (layer1_outputs(6538)));
    layer2_outputs(3013) <= not(layer1_outputs(8257));
    layer2_outputs(3014) <= (layer1_outputs(568)) and not (layer1_outputs(7442));
    layer2_outputs(3015) <= layer1_outputs(10256);
    layer2_outputs(3016) <= not((layer1_outputs(6201)) xor (layer1_outputs(8039)));
    layer2_outputs(3017) <= not((layer1_outputs(1581)) xor (layer1_outputs(9254)));
    layer2_outputs(3018) <= not(layer1_outputs(10930));
    layer2_outputs(3019) <= (layer1_outputs(7638)) and (layer1_outputs(8258));
    layer2_outputs(3020) <= (layer1_outputs(9945)) and not (layer1_outputs(11641));
    layer2_outputs(3021) <= not(layer1_outputs(1587));
    layer2_outputs(3022) <= layer1_outputs(6098);
    layer2_outputs(3023) <= layer1_outputs(1109);
    layer2_outputs(3024) <= not(layer1_outputs(4994));
    layer2_outputs(3025) <= not(layer1_outputs(3003));
    layer2_outputs(3026) <= (layer1_outputs(8621)) xor (layer1_outputs(2473));
    layer2_outputs(3027) <= not(layer1_outputs(11499));
    layer2_outputs(3028) <= not(layer1_outputs(12070));
    layer2_outputs(3029) <= layer1_outputs(4479);
    layer2_outputs(3030) <= not(layer1_outputs(3465));
    layer2_outputs(3031) <= not(layer1_outputs(1326));
    layer2_outputs(3032) <= (layer1_outputs(7026)) and not (layer1_outputs(4635));
    layer2_outputs(3033) <= not((layer1_outputs(5225)) and (layer1_outputs(2303)));
    layer2_outputs(3034) <= layer1_outputs(2067);
    layer2_outputs(3035) <= '1';
    layer2_outputs(3036) <= (layer1_outputs(8194)) xor (layer1_outputs(7130));
    layer2_outputs(3037) <= layer1_outputs(3577);
    layer2_outputs(3038) <= layer1_outputs(8225);
    layer2_outputs(3039) <= not(layer1_outputs(9324));
    layer2_outputs(3040) <= not(layer1_outputs(9949));
    layer2_outputs(3041) <= (layer1_outputs(563)) and (layer1_outputs(7649));
    layer2_outputs(3042) <= (layer1_outputs(7939)) or (layer1_outputs(10401));
    layer2_outputs(3043) <= (layer1_outputs(6990)) xor (layer1_outputs(8170));
    layer2_outputs(3044) <= (layer1_outputs(5317)) and not (layer1_outputs(11743));
    layer2_outputs(3045) <= not((layer1_outputs(10021)) and (layer1_outputs(1832)));
    layer2_outputs(3046) <= not(layer1_outputs(1970));
    layer2_outputs(3047) <= (layer1_outputs(1228)) or (layer1_outputs(7032));
    layer2_outputs(3048) <= not((layer1_outputs(517)) and (layer1_outputs(11741)));
    layer2_outputs(3049) <= layer1_outputs(1835);
    layer2_outputs(3050) <= layer1_outputs(2925);
    layer2_outputs(3051) <= (layer1_outputs(3770)) and not (layer1_outputs(12275));
    layer2_outputs(3052) <= layer1_outputs(9840);
    layer2_outputs(3053) <= (layer1_outputs(5267)) and not (layer1_outputs(11768));
    layer2_outputs(3054) <= (layer1_outputs(8449)) or (layer1_outputs(2234));
    layer2_outputs(3055) <= not((layer1_outputs(3113)) xor (layer1_outputs(2455)));
    layer2_outputs(3056) <= (layer1_outputs(1128)) or (layer1_outputs(10462));
    layer2_outputs(3057) <= (layer1_outputs(8311)) or (layer1_outputs(5529));
    layer2_outputs(3058) <= not((layer1_outputs(4038)) and (layer1_outputs(2229)));
    layer2_outputs(3059) <= not(layer1_outputs(9694));
    layer2_outputs(3060) <= not((layer1_outputs(10603)) or (layer1_outputs(67)));
    layer2_outputs(3061) <= not((layer1_outputs(526)) and (layer1_outputs(1742)));
    layer2_outputs(3062) <= not((layer1_outputs(10336)) xor (layer1_outputs(7551)));
    layer2_outputs(3063) <= not(layer1_outputs(7107));
    layer2_outputs(3064) <= layer1_outputs(8162);
    layer2_outputs(3065) <= (layer1_outputs(4219)) and not (layer1_outputs(12140));
    layer2_outputs(3066) <= '1';
    layer2_outputs(3067) <= (layer1_outputs(9547)) xor (layer1_outputs(11421));
    layer2_outputs(3068) <= not((layer1_outputs(821)) or (layer1_outputs(2336)));
    layer2_outputs(3069) <= not((layer1_outputs(1509)) xor (layer1_outputs(10335)));
    layer2_outputs(3070) <= not((layer1_outputs(7045)) xor (layer1_outputs(5930)));
    layer2_outputs(3071) <= layer1_outputs(4276);
    layer2_outputs(3072) <= not((layer1_outputs(49)) and (layer1_outputs(6405)));
    layer2_outputs(3073) <= not(layer1_outputs(3456));
    layer2_outputs(3074) <= not(layer1_outputs(205));
    layer2_outputs(3075) <= not(layer1_outputs(9265));
    layer2_outputs(3076) <= (layer1_outputs(7610)) or (layer1_outputs(10475));
    layer2_outputs(3077) <= not(layer1_outputs(3504));
    layer2_outputs(3078) <= layer1_outputs(9278);
    layer2_outputs(3079) <= (layer1_outputs(8126)) and (layer1_outputs(8344));
    layer2_outputs(3080) <= not(layer1_outputs(10929));
    layer2_outputs(3081) <= (layer1_outputs(3066)) xor (layer1_outputs(2127));
    layer2_outputs(3082) <= not(layer1_outputs(4054));
    layer2_outputs(3083) <= not((layer1_outputs(911)) or (layer1_outputs(9970)));
    layer2_outputs(3084) <= not(layer1_outputs(710));
    layer2_outputs(3085) <= not(layer1_outputs(10215));
    layer2_outputs(3086) <= not(layer1_outputs(9184));
    layer2_outputs(3087) <= (layer1_outputs(4294)) and (layer1_outputs(2715));
    layer2_outputs(3088) <= layer1_outputs(9679);
    layer2_outputs(3089) <= layer1_outputs(6911);
    layer2_outputs(3090) <= not(layer1_outputs(6816));
    layer2_outputs(3091) <= layer1_outputs(1747);
    layer2_outputs(3092) <= not(layer1_outputs(10991));
    layer2_outputs(3093) <= not(layer1_outputs(11951)) or (layer1_outputs(10497));
    layer2_outputs(3094) <= not(layer1_outputs(3874)) or (layer1_outputs(2836));
    layer2_outputs(3095) <= not((layer1_outputs(9347)) xor (layer1_outputs(11385)));
    layer2_outputs(3096) <= not(layer1_outputs(6459));
    layer2_outputs(3097) <= layer1_outputs(11499);
    layer2_outputs(3098) <= not(layer1_outputs(5480));
    layer2_outputs(3099) <= layer1_outputs(10132);
    layer2_outputs(3100) <= (layer1_outputs(3064)) and (layer1_outputs(6058));
    layer2_outputs(3101) <= not(layer1_outputs(2590));
    layer2_outputs(3102) <= (layer1_outputs(3643)) xor (layer1_outputs(6828));
    layer2_outputs(3103) <= not((layer1_outputs(9118)) xor (layer1_outputs(9545)));
    layer2_outputs(3104) <= (layer1_outputs(11584)) xor (layer1_outputs(7119));
    layer2_outputs(3105) <= not(layer1_outputs(1184));
    layer2_outputs(3106) <= (layer1_outputs(6463)) or (layer1_outputs(7310));
    layer2_outputs(3107) <= (layer1_outputs(7908)) and (layer1_outputs(225));
    layer2_outputs(3108) <= not(layer1_outputs(1732));
    layer2_outputs(3109) <= layer1_outputs(786);
    layer2_outputs(3110) <= (layer1_outputs(1831)) or (layer1_outputs(12385));
    layer2_outputs(3111) <= not((layer1_outputs(6439)) xor (layer1_outputs(7414)));
    layer2_outputs(3112) <= layer1_outputs(3554);
    layer2_outputs(3113) <= (layer1_outputs(6394)) and not (layer1_outputs(630));
    layer2_outputs(3114) <= not(layer1_outputs(1089));
    layer2_outputs(3115) <= (layer1_outputs(1021)) and not (layer1_outputs(14));
    layer2_outputs(3116) <= not(layer1_outputs(2062));
    layer2_outputs(3117) <= layer1_outputs(9297);
    layer2_outputs(3118) <= not(layer1_outputs(5085));
    layer2_outputs(3119) <= not((layer1_outputs(7753)) xor (layer1_outputs(11903)));
    layer2_outputs(3120) <= layer1_outputs(198);
    layer2_outputs(3121) <= not((layer1_outputs(5919)) or (layer1_outputs(4075)));
    layer2_outputs(3122) <= layer1_outputs(5144);
    layer2_outputs(3123) <= (layer1_outputs(11062)) and (layer1_outputs(5595));
    layer2_outputs(3124) <= not((layer1_outputs(4364)) xor (layer1_outputs(10653)));
    layer2_outputs(3125) <= not((layer1_outputs(10817)) xor (layer1_outputs(11877)));
    layer2_outputs(3126) <= (layer1_outputs(158)) xor (layer1_outputs(9621));
    layer2_outputs(3127) <= layer1_outputs(4649);
    layer2_outputs(3128) <= not(layer1_outputs(10781));
    layer2_outputs(3129) <= layer1_outputs(7490);
    layer2_outputs(3130) <= layer1_outputs(8147);
    layer2_outputs(3131) <= not(layer1_outputs(4203));
    layer2_outputs(3132) <= (layer1_outputs(1141)) and not (layer1_outputs(3009));
    layer2_outputs(3133) <= not(layer1_outputs(3997));
    layer2_outputs(3134) <= (layer1_outputs(11466)) or (layer1_outputs(1808));
    layer2_outputs(3135) <= layer1_outputs(8790);
    layer2_outputs(3136) <= layer1_outputs(9129);
    layer2_outputs(3137) <= not((layer1_outputs(7700)) xor (layer1_outputs(4694)));
    layer2_outputs(3138) <= not((layer1_outputs(2703)) and (layer1_outputs(9859)));
    layer2_outputs(3139) <= layer1_outputs(12039);
    layer2_outputs(3140) <= (layer1_outputs(12021)) and not (layer1_outputs(10968));
    layer2_outputs(3141) <= layer1_outputs(7858);
    layer2_outputs(3142) <= not(layer1_outputs(8075)) or (layer1_outputs(4697));
    layer2_outputs(3143) <= (layer1_outputs(11017)) and not (layer1_outputs(3471));
    layer2_outputs(3144) <= not(layer1_outputs(3715)) or (layer1_outputs(10155));
    layer2_outputs(3145) <= not(layer1_outputs(6539));
    layer2_outputs(3146) <= not((layer1_outputs(10466)) xor (layer1_outputs(4514)));
    layer2_outputs(3147) <= (layer1_outputs(4257)) and not (layer1_outputs(5843));
    layer2_outputs(3148) <= layer1_outputs(5367);
    layer2_outputs(3149) <= layer1_outputs(2677);
    layer2_outputs(3150) <= not(layer1_outputs(12727));
    layer2_outputs(3151) <= (layer1_outputs(5820)) and not (layer1_outputs(2401));
    layer2_outputs(3152) <= layer1_outputs(8107);
    layer2_outputs(3153) <= not((layer1_outputs(1630)) xor (layer1_outputs(12757)));
    layer2_outputs(3154) <= '1';
    layer2_outputs(3155) <= not(layer1_outputs(2884));
    layer2_outputs(3156) <= layer1_outputs(12064);
    layer2_outputs(3157) <= not((layer1_outputs(2224)) xor (layer1_outputs(4731)));
    layer2_outputs(3158) <= not((layer1_outputs(9536)) and (layer1_outputs(4989)));
    layer2_outputs(3159) <= not(layer1_outputs(6301));
    layer2_outputs(3160) <= layer1_outputs(1277);
    layer2_outputs(3161) <= not(layer1_outputs(6828)) or (layer1_outputs(889));
    layer2_outputs(3162) <= not(layer1_outputs(5271));
    layer2_outputs(3163) <= not(layer1_outputs(36));
    layer2_outputs(3164) <= (layer1_outputs(12293)) xor (layer1_outputs(5748));
    layer2_outputs(3165) <= not(layer1_outputs(10795)) or (layer1_outputs(2273));
    layer2_outputs(3166) <= not((layer1_outputs(12712)) xor (layer1_outputs(542)));
    layer2_outputs(3167) <= (layer1_outputs(7654)) and not (layer1_outputs(5129));
    layer2_outputs(3168) <= not((layer1_outputs(8316)) or (layer1_outputs(806)));
    layer2_outputs(3169) <= not((layer1_outputs(12403)) xor (layer1_outputs(1917)));
    layer2_outputs(3170) <= (layer1_outputs(3575)) or (layer1_outputs(9089));
    layer2_outputs(3171) <= layer1_outputs(2657);
    layer2_outputs(3172) <= layer1_outputs(1247);
    layer2_outputs(3173) <= (layer1_outputs(129)) or (layer1_outputs(5835));
    layer2_outputs(3174) <= (layer1_outputs(4115)) or (layer1_outputs(8113));
    layer2_outputs(3175) <= not(layer1_outputs(8241));
    layer2_outputs(3176) <= not(layer1_outputs(5760)) or (layer1_outputs(11978));
    layer2_outputs(3177) <= not(layer1_outputs(5883));
    layer2_outputs(3178) <= (layer1_outputs(239)) or (layer1_outputs(1488));
    layer2_outputs(3179) <= not(layer1_outputs(9454));
    layer2_outputs(3180) <= (layer1_outputs(7727)) or (layer1_outputs(1231));
    layer2_outputs(3181) <= not((layer1_outputs(7740)) and (layer1_outputs(10172)));
    layer2_outputs(3182) <= not((layer1_outputs(11303)) xor (layer1_outputs(10405)));
    layer2_outputs(3183) <= not(layer1_outputs(476));
    layer2_outputs(3184) <= (layer1_outputs(4337)) and (layer1_outputs(6676));
    layer2_outputs(3185) <= not(layer1_outputs(5869));
    layer2_outputs(3186) <= (layer1_outputs(9354)) and not (layer1_outputs(6380));
    layer2_outputs(3187) <= not(layer1_outputs(4116));
    layer2_outputs(3188) <= not(layer1_outputs(6357)) or (layer1_outputs(11634));
    layer2_outputs(3189) <= not((layer1_outputs(11250)) or (layer1_outputs(12246)));
    layer2_outputs(3190) <= not(layer1_outputs(8622));
    layer2_outputs(3191) <= layer1_outputs(11435);
    layer2_outputs(3192) <= not((layer1_outputs(4720)) or (layer1_outputs(5405)));
    layer2_outputs(3193) <= not(layer1_outputs(8139));
    layer2_outputs(3194) <= (layer1_outputs(9240)) xor (layer1_outputs(6446));
    layer2_outputs(3195) <= not(layer1_outputs(5834));
    layer2_outputs(3196) <= not((layer1_outputs(2605)) xor (layer1_outputs(4080)));
    layer2_outputs(3197) <= (layer1_outputs(6155)) and not (layer1_outputs(8375));
    layer2_outputs(3198) <= (layer1_outputs(4260)) and not (layer1_outputs(8346));
    layer2_outputs(3199) <= not((layer1_outputs(2238)) xor (layer1_outputs(6740)));
    layer2_outputs(3200) <= not(layer1_outputs(2411));
    layer2_outputs(3201) <= not((layer1_outputs(2910)) or (layer1_outputs(9417)));
    layer2_outputs(3202) <= not(layer1_outputs(3847)) or (layer1_outputs(8950));
    layer2_outputs(3203) <= not(layer1_outputs(3126));
    layer2_outputs(3204) <= not(layer1_outputs(2954)) or (layer1_outputs(1523));
    layer2_outputs(3205) <= layer1_outputs(462);
    layer2_outputs(3206) <= not((layer1_outputs(4076)) or (layer1_outputs(3622)));
    layer2_outputs(3207) <= not((layer1_outputs(5260)) and (layer1_outputs(2963)));
    layer2_outputs(3208) <= layer1_outputs(3384);
    layer2_outputs(3209) <= not(layer1_outputs(9542));
    layer2_outputs(3210) <= not(layer1_outputs(12474)) or (layer1_outputs(5039));
    layer2_outputs(3211) <= not((layer1_outputs(11916)) and (layer1_outputs(7928)));
    layer2_outputs(3212) <= not(layer1_outputs(6288));
    layer2_outputs(3213) <= layer1_outputs(3789);
    layer2_outputs(3214) <= not(layer1_outputs(1536));
    layer2_outputs(3215) <= not(layer1_outputs(1349));
    layer2_outputs(3216) <= not(layer1_outputs(10509));
    layer2_outputs(3217) <= not(layer1_outputs(12055));
    layer2_outputs(3218) <= (layer1_outputs(2802)) xor (layer1_outputs(7302));
    layer2_outputs(3219) <= (layer1_outputs(2406)) and (layer1_outputs(10225));
    layer2_outputs(3220) <= '1';
    layer2_outputs(3221) <= not(layer1_outputs(8885));
    layer2_outputs(3222) <= not((layer1_outputs(8579)) and (layer1_outputs(10062)));
    layer2_outputs(3223) <= not(layer1_outputs(9142));
    layer2_outputs(3224) <= '0';
    layer2_outputs(3225) <= not(layer1_outputs(649));
    layer2_outputs(3226) <= (layer1_outputs(5115)) and not (layer1_outputs(6218));
    layer2_outputs(3227) <= not(layer1_outputs(3049)) or (layer1_outputs(7855));
    layer2_outputs(3228) <= not((layer1_outputs(1559)) and (layer1_outputs(2737)));
    layer2_outputs(3229) <= layer1_outputs(9494);
    layer2_outputs(3230) <= not((layer1_outputs(4728)) xor (layer1_outputs(11119)));
    layer2_outputs(3231) <= layer1_outputs(10129);
    layer2_outputs(3232) <= not(layer1_outputs(2695));
    layer2_outputs(3233) <= layer1_outputs(12514);
    layer2_outputs(3234) <= (layer1_outputs(5696)) and not (layer1_outputs(494));
    layer2_outputs(3235) <= not(layer1_outputs(1741)) or (layer1_outputs(2980));
    layer2_outputs(3236) <= not(layer1_outputs(12749));
    layer2_outputs(3237) <= layer1_outputs(11404);
    layer2_outputs(3238) <= layer1_outputs(616);
    layer2_outputs(3239) <= not((layer1_outputs(5821)) or (layer1_outputs(9217)));
    layer2_outputs(3240) <= not(layer1_outputs(7245));
    layer2_outputs(3241) <= not(layer1_outputs(8819));
    layer2_outputs(3242) <= (layer1_outputs(804)) and not (layer1_outputs(426));
    layer2_outputs(3243) <= (layer1_outputs(3376)) or (layer1_outputs(11473));
    layer2_outputs(3244) <= layer1_outputs(2346);
    layer2_outputs(3245) <= not(layer1_outputs(11670));
    layer2_outputs(3246) <= not((layer1_outputs(10442)) xor (layer1_outputs(2950)));
    layer2_outputs(3247) <= not((layer1_outputs(9080)) or (layer1_outputs(6529)));
    layer2_outputs(3248) <= (layer1_outputs(8914)) xor (layer1_outputs(3419));
    layer2_outputs(3249) <= layer1_outputs(4159);
    layer2_outputs(3250) <= (layer1_outputs(4953)) xor (layer1_outputs(10419));
    layer2_outputs(3251) <= not((layer1_outputs(2064)) xor (layer1_outputs(9565)));
    layer2_outputs(3252) <= not(layer1_outputs(8216));
    layer2_outputs(3253) <= (layer1_outputs(921)) and not (layer1_outputs(6351));
    layer2_outputs(3254) <= not(layer1_outputs(7265)) or (layer1_outputs(10658));
    layer2_outputs(3255) <= not(layer1_outputs(9840));
    layer2_outputs(3256) <= layer1_outputs(11399);
    layer2_outputs(3257) <= (layer1_outputs(189)) and not (layer1_outputs(9830));
    layer2_outputs(3258) <= not((layer1_outputs(8663)) or (layer1_outputs(9588)));
    layer2_outputs(3259) <= layer1_outputs(158);
    layer2_outputs(3260) <= not(layer1_outputs(3876));
    layer2_outputs(3261) <= not((layer1_outputs(11400)) or (layer1_outputs(6258)));
    layer2_outputs(3262) <= not(layer1_outputs(10277));
    layer2_outputs(3263) <= layer1_outputs(11662);
    layer2_outputs(3264) <= layer1_outputs(5618);
    layer2_outputs(3265) <= (layer1_outputs(11559)) and not (layer1_outputs(11254));
    layer2_outputs(3266) <= not(layer1_outputs(5431));
    layer2_outputs(3267) <= layer1_outputs(1398);
    layer2_outputs(3268) <= not((layer1_outputs(4063)) and (layer1_outputs(11588)));
    layer2_outputs(3269) <= (layer1_outputs(1607)) or (layer1_outputs(10296));
    layer2_outputs(3270) <= not(layer1_outputs(1939));
    layer2_outputs(3271) <= (layer1_outputs(6729)) and (layer1_outputs(5677));
    layer2_outputs(3272) <= (layer1_outputs(10502)) and not (layer1_outputs(5054));
    layer2_outputs(3273) <= layer1_outputs(10245);
    layer2_outputs(3274) <= layer1_outputs(8058);
    layer2_outputs(3275) <= not((layer1_outputs(2807)) or (layer1_outputs(2624)));
    layer2_outputs(3276) <= not(layer1_outputs(12655));
    layer2_outputs(3277) <= layer1_outputs(9422);
    layer2_outputs(3278) <= not((layer1_outputs(10511)) xor (layer1_outputs(9495)));
    layer2_outputs(3279) <= not((layer1_outputs(9817)) and (layer1_outputs(3773)));
    layer2_outputs(3280) <= (layer1_outputs(12389)) or (layer1_outputs(3540));
    layer2_outputs(3281) <= not((layer1_outputs(11021)) xor (layer1_outputs(7801)));
    layer2_outputs(3282) <= (layer1_outputs(2023)) xor (layer1_outputs(10331));
    layer2_outputs(3283) <= layer1_outputs(4521);
    layer2_outputs(3284) <= layer1_outputs(6344);
    layer2_outputs(3285) <= (layer1_outputs(6630)) xor (layer1_outputs(8602));
    layer2_outputs(3286) <= (layer1_outputs(1367)) or (layer1_outputs(7778));
    layer2_outputs(3287) <= not(layer1_outputs(4878));
    layer2_outputs(3288) <= layer1_outputs(873);
    layer2_outputs(3289) <= not((layer1_outputs(179)) xor (layer1_outputs(4318)));
    layer2_outputs(3290) <= (layer1_outputs(7909)) and not (layer1_outputs(7668));
    layer2_outputs(3291) <= layer1_outputs(2841);
    layer2_outputs(3292) <= not(layer1_outputs(2316)) or (layer1_outputs(9752));
    layer2_outputs(3293) <= layer1_outputs(5093);
    layer2_outputs(3294) <= not((layer1_outputs(12785)) and (layer1_outputs(3907)));
    layer2_outputs(3295) <= layer1_outputs(10027);
    layer2_outputs(3296) <= not(layer1_outputs(9721));
    layer2_outputs(3297) <= not(layer1_outputs(8470));
    layer2_outputs(3298) <= not(layer1_outputs(7454)) or (layer1_outputs(11440));
    layer2_outputs(3299) <= layer1_outputs(8827);
    layer2_outputs(3300) <= not((layer1_outputs(5095)) xor (layer1_outputs(10756)));
    layer2_outputs(3301) <= layer1_outputs(11146);
    layer2_outputs(3302) <= not(layer1_outputs(11791));
    layer2_outputs(3303) <= (layer1_outputs(8366)) or (layer1_outputs(7744));
    layer2_outputs(3304) <= not(layer1_outputs(12467));
    layer2_outputs(3305) <= not(layer1_outputs(12621));
    layer2_outputs(3306) <= (layer1_outputs(10442)) xor (layer1_outputs(9966));
    layer2_outputs(3307) <= not(layer1_outputs(12763));
    layer2_outputs(3308) <= layer1_outputs(9134);
    layer2_outputs(3309) <= not(layer1_outputs(9677));
    layer2_outputs(3310) <= not(layer1_outputs(8109));
    layer2_outputs(3311) <= layer1_outputs(9934);
    layer2_outputs(3312) <= (layer1_outputs(10308)) and (layer1_outputs(11137));
    layer2_outputs(3313) <= not(layer1_outputs(8235));
    layer2_outputs(3314) <= (layer1_outputs(5197)) and not (layer1_outputs(3361));
    layer2_outputs(3315) <= not(layer1_outputs(4603)) or (layer1_outputs(12558));
    layer2_outputs(3316) <= not(layer1_outputs(6406));
    layer2_outputs(3317) <= layer1_outputs(1900);
    layer2_outputs(3318) <= (layer1_outputs(11626)) and not (layer1_outputs(7161));
    layer2_outputs(3319) <= layer1_outputs(6999);
    layer2_outputs(3320) <= layer1_outputs(9953);
    layer2_outputs(3321) <= (layer1_outputs(8384)) and not (layer1_outputs(12114));
    layer2_outputs(3322) <= layer1_outputs(6738);
    layer2_outputs(3323) <= not(layer1_outputs(2125));
    layer2_outputs(3324) <= (layer1_outputs(3277)) xor (layer1_outputs(10350));
    layer2_outputs(3325) <= not(layer1_outputs(10297));
    layer2_outputs(3326) <= layer1_outputs(4642);
    layer2_outputs(3327) <= (layer1_outputs(5232)) xor (layer1_outputs(2113));
    layer2_outputs(3328) <= not(layer1_outputs(1054)) or (layer1_outputs(1161));
    layer2_outputs(3329) <= not((layer1_outputs(9446)) or (layer1_outputs(11716)));
    layer2_outputs(3330) <= (layer1_outputs(7332)) xor (layer1_outputs(12655));
    layer2_outputs(3331) <= (layer1_outputs(2805)) and not (layer1_outputs(10616));
    layer2_outputs(3332) <= (layer1_outputs(1451)) and (layer1_outputs(9501));
    layer2_outputs(3333) <= not(layer1_outputs(5230)) or (layer1_outputs(7065));
    layer2_outputs(3334) <= not(layer1_outputs(7507));
    layer2_outputs(3335) <= layer1_outputs(11067);
    layer2_outputs(3336) <= layer1_outputs(5952);
    layer2_outputs(3337) <= not(layer1_outputs(6645));
    layer2_outputs(3338) <= not((layer1_outputs(11981)) or (layer1_outputs(1201)));
    layer2_outputs(3339) <= (layer1_outputs(6592)) xor (layer1_outputs(11648));
    layer2_outputs(3340) <= not((layer1_outputs(360)) and (layer1_outputs(5936)));
    layer2_outputs(3341) <= (layer1_outputs(9319)) or (layer1_outputs(8683));
    layer2_outputs(3342) <= not(layer1_outputs(6516));
    layer2_outputs(3343) <= not(layer1_outputs(1000)) or (layer1_outputs(1965));
    layer2_outputs(3344) <= (layer1_outputs(7343)) and not (layer1_outputs(4804));
    layer2_outputs(3345) <= not(layer1_outputs(9047));
    layer2_outputs(3346) <= layer1_outputs(5502);
    layer2_outputs(3347) <= (layer1_outputs(3557)) and not (layer1_outputs(4264));
    layer2_outputs(3348) <= not(layer1_outputs(5318)) or (layer1_outputs(7516));
    layer2_outputs(3349) <= (layer1_outputs(2756)) or (layer1_outputs(4549));
    layer2_outputs(3350) <= layer1_outputs(4509);
    layer2_outputs(3351) <= layer1_outputs(2969);
    layer2_outputs(3352) <= layer1_outputs(6147);
    layer2_outputs(3353) <= not((layer1_outputs(3655)) xor (layer1_outputs(839)));
    layer2_outputs(3354) <= layer1_outputs(3678);
    layer2_outputs(3355) <= layer1_outputs(101);
    layer2_outputs(3356) <= not((layer1_outputs(7704)) xor (layer1_outputs(11840)));
    layer2_outputs(3357) <= not(layer1_outputs(9028));
    layer2_outputs(3358) <= layer1_outputs(12628);
    layer2_outputs(3359) <= not((layer1_outputs(7747)) xor (layer1_outputs(364)));
    layer2_outputs(3360) <= layer1_outputs(6528);
    layer2_outputs(3361) <= not(layer1_outputs(1437));
    layer2_outputs(3362) <= not(layer1_outputs(93)) or (layer1_outputs(5205));
    layer2_outputs(3363) <= layer1_outputs(6137);
    layer2_outputs(3364) <= (layer1_outputs(8025)) or (layer1_outputs(6570));
    layer2_outputs(3365) <= (layer1_outputs(11197)) and not (layer1_outputs(2180));
    layer2_outputs(3366) <= (layer1_outputs(2575)) and not (layer1_outputs(4112));
    layer2_outputs(3367) <= layer1_outputs(2760);
    layer2_outputs(3368) <= layer1_outputs(5896);
    layer2_outputs(3369) <= layer1_outputs(7895);
    layer2_outputs(3370) <= not(layer1_outputs(2663));
    layer2_outputs(3371) <= not(layer1_outputs(5037));
    layer2_outputs(3372) <= not(layer1_outputs(4531));
    layer2_outputs(3373) <= layer1_outputs(7354);
    layer2_outputs(3374) <= not(layer1_outputs(388));
    layer2_outputs(3375) <= (layer1_outputs(11308)) and not (layer1_outputs(8605));
    layer2_outputs(3376) <= layer1_outputs(1710);
    layer2_outputs(3377) <= layer1_outputs(247);
    layer2_outputs(3378) <= '0';
    layer2_outputs(3379) <= not(layer1_outputs(5840));
    layer2_outputs(3380) <= not((layer1_outputs(6918)) and (layer1_outputs(10030)));
    layer2_outputs(3381) <= (layer1_outputs(10979)) and not (layer1_outputs(5805));
    layer2_outputs(3382) <= layer1_outputs(2482);
    layer2_outputs(3383) <= not(layer1_outputs(4463)) or (layer1_outputs(7852));
    layer2_outputs(3384) <= not(layer1_outputs(2586));
    layer2_outputs(3385) <= not((layer1_outputs(1781)) xor (layer1_outputs(9795)));
    layer2_outputs(3386) <= (layer1_outputs(1667)) and (layer1_outputs(3705));
    layer2_outputs(3387) <= not(layer1_outputs(3462));
    layer2_outputs(3388) <= not(layer1_outputs(5124));
    layer2_outputs(3389) <= layer1_outputs(11333);
    layer2_outputs(3390) <= (layer1_outputs(9219)) xor (layer1_outputs(5545));
    layer2_outputs(3391) <= (layer1_outputs(10547)) or (layer1_outputs(4875));
    layer2_outputs(3392) <= layer1_outputs(9004);
    layer2_outputs(3393) <= layer1_outputs(7570);
    layer2_outputs(3394) <= (layer1_outputs(4990)) and (layer1_outputs(5907));
    layer2_outputs(3395) <= not((layer1_outputs(6132)) and (layer1_outputs(7540)));
    layer2_outputs(3396) <= layer1_outputs(10163);
    layer2_outputs(3397) <= not(layer1_outputs(1806));
    layer2_outputs(3398) <= layer1_outputs(7128);
    layer2_outputs(3399) <= not(layer1_outputs(11932));
    layer2_outputs(3400) <= not((layer1_outputs(4206)) or (layer1_outputs(9698)));
    layer2_outputs(3401) <= not((layer1_outputs(8668)) xor (layer1_outputs(2673)));
    layer2_outputs(3402) <= not(layer1_outputs(4685)) or (layer1_outputs(11226));
    layer2_outputs(3403) <= layer1_outputs(5429);
    layer2_outputs(3404) <= layer1_outputs(1521);
    layer2_outputs(3405) <= not(layer1_outputs(6734));
    layer2_outputs(3406) <= not(layer1_outputs(2350));
    layer2_outputs(3407) <= not(layer1_outputs(12784)) or (layer1_outputs(10263));
    layer2_outputs(3408) <= not((layer1_outputs(7904)) and (layer1_outputs(1366)));
    layer2_outputs(3409) <= layer1_outputs(9523);
    layer2_outputs(3410) <= not(layer1_outputs(2433)) or (layer1_outputs(2622));
    layer2_outputs(3411) <= not(layer1_outputs(1094)) or (layer1_outputs(930));
    layer2_outputs(3412) <= layer1_outputs(9302);
    layer2_outputs(3413) <= layer1_outputs(10468);
    layer2_outputs(3414) <= layer1_outputs(3012);
    layer2_outputs(3415) <= layer1_outputs(10064);
    layer2_outputs(3416) <= layer1_outputs(2899);
    layer2_outputs(3417) <= (layer1_outputs(532)) or (layer1_outputs(9223));
    layer2_outputs(3418) <= not(layer1_outputs(8373)) or (layer1_outputs(2525));
    layer2_outputs(3419) <= (layer1_outputs(10167)) and not (layer1_outputs(5911));
    layer2_outputs(3420) <= layer1_outputs(1971);
    layer2_outputs(3421) <= (layer1_outputs(8772)) xor (layer1_outputs(1775));
    layer2_outputs(3422) <= not((layer1_outputs(8130)) and (layer1_outputs(8656)));
    layer2_outputs(3423) <= layer1_outputs(4694);
    layer2_outputs(3424) <= (layer1_outputs(6434)) xor (layer1_outputs(10774));
    layer2_outputs(3425) <= not(layer1_outputs(11238));
    layer2_outputs(3426) <= (layer1_outputs(9001)) xor (layer1_outputs(4700));
    layer2_outputs(3427) <= not(layer1_outputs(8343)) or (layer1_outputs(3355));
    layer2_outputs(3428) <= not(layer1_outputs(1974));
    layer2_outputs(3429) <= not((layer1_outputs(9569)) xor (layer1_outputs(11179)));
    layer2_outputs(3430) <= (layer1_outputs(802)) and not (layer1_outputs(7334));
    layer2_outputs(3431) <= (layer1_outputs(9739)) and not (layer1_outputs(11486));
    layer2_outputs(3432) <= not(layer1_outputs(4291)) or (layer1_outputs(767));
    layer2_outputs(3433) <= not(layer1_outputs(11594));
    layer2_outputs(3434) <= not((layer1_outputs(5891)) or (layer1_outputs(6693)));
    layer2_outputs(3435) <= not(layer1_outputs(9507));
    layer2_outputs(3436) <= layer1_outputs(11880);
    layer2_outputs(3437) <= (layer1_outputs(7892)) xor (layer1_outputs(11859));
    layer2_outputs(3438) <= layer1_outputs(5039);
    layer2_outputs(3439) <= layer1_outputs(10177);
    layer2_outputs(3440) <= not((layer1_outputs(4533)) xor (layer1_outputs(10880)));
    layer2_outputs(3441) <= (layer1_outputs(5388)) and (layer1_outputs(5169));
    layer2_outputs(3442) <= layer1_outputs(10047);
    layer2_outputs(3443) <= not(layer1_outputs(7838)) or (layer1_outputs(9216));
    layer2_outputs(3444) <= not(layer1_outputs(3271)) or (layer1_outputs(11202));
    layer2_outputs(3445) <= not(layer1_outputs(8374));
    layer2_outputs(3446) <= (layer1_outputs(8644)) and not (layer1_outputs(6143));
    layer2_outputs(3447) <= layer1_outputs(1720);
    layer2_outputs(3448) <= not(layer1_outputs(11332)) or (layer1_outputs(718));
    layer2_outputs(3449) <= not((layer1_outputs(1951)) and (layer1_outputs(7064)));
    layer2_outputs(3450) <= (layer1_outputs(3656)) and not (layer1_outputs(12595));
    layer2_outputs(3451) <= layer1_outputs(1687);
    layer2_outputs(3452) <= (layer1_outputs(2390)) xor (layer1_outputs(12488));
    layer2_outputs(3453) <= not(layer1_outputs(4155));
    layer2_outputs(3454) <= not((layer1_outputs(5605)) or (layer1_outputs(12710)));
    layer2_outputs(3455) <= not((layer1_outputs(8747)) and (layer1_outputs(12204)));
    layer2_outputs(3456) <= (layer1_outputs(3863)) or (layer1_outputs(3438));
    layer2_outputs(3457) <= not(layer1_outputs(7809));
    layer2_outputs(3458) <= not(layer1_outputs(9002));
    layer2_outputs(3459) <= not(layer1_outputs(9520));
    layer2_outputs(3460) <= (layer1_outputs(6502)) xor (layer1_outputs(1941));
    layer2_outputs(3461) <= not(layer1_outputs(261)) or (layer1_outputs(8407));
    layer2_outputs(3462) <= layer1_outputs(589);
    layer2_outputs(3463) <= not(layer1_outputs(10241));
    layer2_outputs(3464) <= (layer1_outputs(10889)) and not (layer1_outputs(10540));
    layer2_outputs(3465) <= not(layer1_outputs(10745));
    layer2_outputs(3466) <= layer1_outputs(6772);
    layer2_outputs(3467) <= layer1_outputs(1811);
    layer2_outputs(3468) <= not((layer1_outputs(2814)) and (layer1_outputs(8868)));
    layer2_outputs(3469) <= not((layer1_outputs(8420)) or (layer1_outputs(3678)));
    layer2_outputs(3470) <= not(layer1_outputs(2857));
    layer2_outputs(3471) <= layer1_outputs(2724);
    layer2_outputs(3472) <= not(layer1_outputs(12493));
    layer2_outputs(3473) <= layer1_outputs(10970);
    layer2_outputs(3474) <= layer1_outputs(845);
    layer2_outputs(3475) <= not(layer1_outputs(9082));
    layer2_outputs(3476) <= not(layer1_outputs(261));
    layer2_outputs(3477) <= not(layer1_outputs(10587)) or (layer1_outputs(5029));
    layer2_outputs(3478) <= not(layer1_outputs(4334));
    layer2_outputs(3479) <= not(layer1_outputs(8750)) or (layer1_outputs(12514));
    layer2_outputs(3480) <= (layer1_outputs(9714)) or (layer1_outputs(3447));
    layer2_outputs(3481) <= (layer1_outputs(8368)) and not (layer1_outputs(9598));
    layer2_outputs(3482) <= layer1_outputs(3387);
    layer2_outputs(3483) <= (layer1_outputs(29)) xor (layer1_outputs(9073));
    layer2_outputs(3484) <= not(layer1_outputs(10855));
    layer2_outputs(3485) <= layer1_outputs(3026);
    layer2_outputs(3486) <= (layer1_outputs(10286)) and not (layer1_outputs(12177));
    layer2_outputs(3487) <= '0';
    layer2_outputs(3488) <= layer1_outputs(4579);
    layer2_outputs(3489) <= not(layer1_outputs(6060));
    layer2_outputs(3490) <= not(layer1_outputs(10576));
    layer2_outputs(3491) <= layer1_outputs(8635);
    layer2_outputs(3492) <= not(layer1_outputs(8507));
    layer2_outputs(3493) <= not(layer1_outputs(10404));
    layer2_outputs(3494) <= not(layer1_outputs(12541));
    layer2_outputs(3495) <= layer1_outputs(12627);
    layer2_outputs(3496) <= not(layer1_outputs(3882));
    layer2_outputs(3497) <= not(layer1_outputs(8451));
    layer2_outputs(3498) <= not(layer1_outputs(5321));
    layer2_outputs(3499) <= not(layer1_outputs(4339));
    layer2_outputs(3500) <= not(layer1_outputs(10618));
    layer2_outputs(3501) <= not((layer1_outputs(7299)) and (layer1_outputs(11536)));
    layer2_outputs(3502) <= layer1_outputs(7491);
    layer2_outputs(3503) <= (layer1_outputs(9516)) or (layer1_outputs(9124));
    layer2_outputs(3504) <= not(layer1_outputs(2165)) or (layer1_outputs(11198));
    layer2_outputs(3505) <= layer1_outputs(979);
    layer2_outputs(3506) <= not((layer1_outputs(11736)) xor (layer1_outputs(3674)));
    layer2_outputs(3507) <= not(layer1_outputs(9115)) or (layer1_outputs(7441));
    layer2_outputs(3508) <= not(layer1_outputs(596));
    layer2_outputs(3509) <= not(layer1_outputs(10342));
    layer2_outputs(3510) <= layer1_outputs(7157);
    layer2_outputs(3511) <= not(layer1_outputs(2707));
    layer2_outputs(3512) <= layer1_outputs(6363);
    layer2_outputs(3513) <= not(layer1_outputs(6063));
    layer2_outputs(3514) <= not(layer1_outputs(4054));
    layer2_outputs(3515) <= not(layer1_outputs(7319));
    layer2_outputs(3516) <= layer1_outputs(5221);
    layer2_outputs(3517) <= layer1_outputs(2227);
    layer2_outputs(3518) <= not(layer1_outputs(7124));
    layer2_outputs(3519) <= not(layer1_outputs(8692)) or (layer1_outputs(7627));
    layer2_outputs(3520) <= layer1_outputs(12781);
    layer2_outputs(3521) <= not((layer1_outputs(8243)) and (layer1_outputs(12634)));
    layer2_outputs(3522) <= layer1_outputs(7332);
    layer2_outputs(3523) <= layer1_outputs(7558);
    layer2_outputs(3524) <= not(layer1_outputs(2709)) or (layer1_outputs(12399));
    layer2_outputs(3525) <= not(layer1_outputs(12596));
    layer2_outputs(3526) <= not((layer1_outputs(1559)) xor (layer1_outputs(12163)));
    layer2_outputs(3527) <= not((layer1_outputs(8524)) or (layer1_outputs(12797)));
    layer2_outputs(3528) <= not(layer1_outputs(9329));
    layer2_outputs(3529) <= layer1_outputs(6900);
    layer2_outputs(3530) <= not((layer1_outputs(6267)) xor (layer1_outputs(6331)));
    layer2_outputs(3531) <= layer1_outputs(4613);
    layer2_outputs(3532) <= not(layer1_outputs(10847));
    layer2_outputs(3533) <= not(layer1_outputs(7322));
    layer2_outputs(3534) <= layer1_outputs(9477);
    layer2_outputs(3535) <= not(layer1_outputs(7132)) or (layer1_outputs(1683));
    layer2_outputs(3536) <= (layer1_outputs(898)) and not (layer1_outputs(5926));
    layer2_outputs(3537) <= not((layer1_outputs(11167)) xor (layer1_outputs(12755)));
    layer2_outputs(3538) <= not(layer1_outputs(461)) or (layer1_outputs(11723));
    layer2_outputs(3539) <= not(layer1_outputs(781));
    layer2_outputs(3540) <= not(layer1_outputs(6656));
    layer2_outputs(3541) <= not(layer1_outputs(4889)) or (layer1_outputs(7940));
    layer2_outputs(3542) <= (layer1_outputs(7463)) and not (layer1_outputs(2607));
    layer2_outputs(3543) <= layer1_outputs(1909);
    layer2_outputs(3544) <= '0';
    layer2_outputs(3545) <= (layer1_outputs(3919)) and (layer1_outputs(2650));
    layer2_outputs(3546) <= not((layer1_outputs(4162)) or (layer1_outputs(11046)));
    layer2_outputs(3547) <= '0';
    layer2_outputs(3548) <= not(layer1_outputs(2136)) or (layer1_outputs(7652));
    layer2_outputs(3549) <= not(layer1_outputs(377)) or (layer1_outputs(4938));
    layer2_outputs(3550) <= not(layer1_outputs(3447));
    layer2_outputs(3551) <= layer1_outputs(244);
    layer2_outputs(3552) <= layer1_outputs(8843);
    layer2_outputs(3553) <= not(layer1_outputs(6323));
    layer2_outputs(3554) <= not(layer1_outputs(2619));
    layer2_outputs(3555) <= layer1_outputs(8528);
    layer2_outputs(3556) <= layer1_outputs(6576);
    layer2_outputs(3557) <= (layer1_outputs(838)) or (layer1_outputs(6164));
    layer2_outputs(3558) <= layer1_outputs(11469);
    layer2_outputs(3559) <= not(layer1_outputs(5520));
    layer2_outputs(3560) <= (layer1_outputs(830)) or (layer1_outputs(2515));
    layer2_outputs(3561) <= (layer1_outputs(7743)) or (layer1_outputs(4536));
    layer2_outputs(3562) <= not(layer1_outputs(11320));
    layer2_outputs(3563) <= layer1_outputs(2740);
    layer2_outputs(3564) <= layer1_outputs(11514);
    layer2_outputs(3565) <= not(layer1_outputs(6059));
    layer2_outputs(3566) <= not(layer1_outputs(5004));
    layer2_outputs(3567) <= layer1_outputs(1651);
    layer2_outputs(3568) <= layer1_outputs(5186);
    layer2_outputs(3569) <= not(layer1_outputs(7562));
    layer2_outputs(3570) <= layer1_outputs(5765);
    layer2_outputs(3571) <= (layer1_outputs(10893)) xor (layer1_outputs(1546));
    layer2_outputs(3572) <= not(layer1_outputs(167));
    layer2_outputs(3573) <= not(layer1_outputs(8465));
    layer2_outputs(3574) <= not(layer1_outputs(8521));
    layer2_outputs(3575) <= not(layer1_outputs(3565));
    layer2_outputs(3576) <= layer1_outputs(12147);
    layer2_outputs(3577) <= (layer1_outputs(74)) and (layer1_outputs(11424));
    layer2_outputs(3578) <= layer1_outputs(8442);
    layer2_outputs(3579) <= (layer1_outputs(6752)) and (layer1_outputs(1165));
    layer2_outputs(3580) <= (layer1_outputs(7509)) or (layer1_outputs(5617));
    layer2_outputs(3581) <= not(layer1_outputs(2487));
    layer2_outputs(3582) <= layer1_outputs(8671);
    layer2_outputs(3583) <= not((layer1_outputs(1422)) and (layer1_outputs(5519)));
    layer2_outputs(3584) <= not((layer1_outputs(7302)) or (layer1_outputs(391)));
    layer2_outputs(3585) <= not((layer1_outputs(129)) xor (layer1_outputs(1351)));
    layer2_outputs(3586) <= not(layer1_outputs(7736));
    layer2_outputs(3587) <= layer1_outputs(3136);
    layer2_outputs(3588) <= not((layer1_outputs(12232)) and (layer1_outputs(6244)));
    layer2_outputs(3589) <= not(layer1_outputs(6537)) or (layer1_outputs(2711));
    layer2_outputs(3590) <= (layer1_outputs(6630)) and (layer1_outputs(10963));
    layer2_outputs(3591) <= layer1_outputs(2595);
    layer2_outputs(3592) <= not(layer1_outputs(7241));
    layer2_outputs(3593) <= not(layer1_outputs(6320));
    layer2_outputs(3594) <= layer1_outputs(10297);
    layer2_outputs(3595) <= (layer1_outputs(9464)) and not (layer1_outputs(410));
    layer2_outputs(3596) <= layer1_outputs(12507);
    layer2_outputs(3597) <= not(layer1_outputs(9971));
    layer2_outputs(3598) <= layer1_outputs(8511);
    layer2_outputs(3599) <= not(layer1_outputs(4692)) or (layer1_outputs(7230));
    layer2_outputs(3600) <= not(layer1_outputs(701)) or (layer1_outputs(9854));
    layer2_outputs(3601) <= (layer1_outputs(9456)) and not (layer1_outputs(2788));
    layer2_outputs(3602) <= (layer1_outputs(4515)) or (layer1_outputs(2910));
    layer2_outputs(3603) <= not(layer1_outputs(4634));
    layer2_outputs(3604) <= not(layer1_outputs(9962));
    layer2_outputs(3605) <= not(layer1_outputs(9684));
    layer2_outputs(3606) <= layer1_outputs(11338);
    layer2_outputs(3607) <= not((layer1_outputs(1047)) xor (layer1_outputs(218)));
    layer2_outputs(3608) <= not((layer1_outputs(331)) or (layer1_outputs(5155)));
    layer2_outputs(3609) <= (layer1_outputs(8681)) and (layer1_outputs(10414));
    layer2_outputs(3610) <= (layer1_outputs(8456)) and not (layer1_outputs(5395));
    layer2_outputs(3611) <= (layer1_outputs(5071)) and not (layer1_outputs(10785));
    layer2_outputs(3612) <= (layer1_outputs(4658)) and not (layer1_outputs(11627));
    layer2_outputs(3613) <= not(layer1_outputs(2343));
    layer2_outputs(3614) <= layer1_outputs(1210);
    layer2_outputs(3615) <= (layer1_outputs(10846)) and not (layer1_outputs(7025));
    layer2_outputs(3616) <= (layer1_outputs(3210)) or (layer1_outputs(4897));
    layer2_outputs(3617) <= (layer1_outputs(10686)) and not (layer1_outputs(10150));
    layer2_outputs(3618) <= layer1_outputs(5233);
    layer2_outputs(3619) <= (layer1_outputs(8570)) or (layer1_outputs(11592));
    layer2_outputs(3620) <= not(layer1_outputs(982));
    layer2_outputs(3621) <= not((layer1_outputs(11018)) xor (layer1_outputs(5329)));
    layer2_outputs(3622) <= layer1_outputs(5166);
    layer2_outputs(3623) <= not((layer1_outputs(12371)) or (layer1_outputs(5211)));
    layer2_outputs(3624) <= (layer1_outputs(966)) and (layer1_outputs(1351));
    layer2_outputs(3625) <= (layer1_outputs(7673)) and (layer1_outputs(5062));
    layer2_outputs(3626) <= (layer1_outputs(11493)) xor (layer1_outputs(8117));
    layer2_outputs(3627) <= not(layer1_outputs(5983));
    layer2_outputs(3628) <= not((layer1_outputs(4385)) xor (layer1_outputs(10333)));
    layer2_outputs(3629) <= not(layer1_outputs(12215));
    layer2_outputs(3630) <= layer1_outputs(6055);
    layer2_outputs(3631) <= not(layer1_outputs(9492));
    layer2_outputs(3632) <= not((layer1_outputs(7854)) and (layer1_outputs(5424)));
    layer2_outputs(3633) <= layer1_outputs(5018);
    layer2_outputs(3634) <= (layer1_outputs(12056)) or (layer1_outputs(8591));
    layer2_outputs(3635) <= layer1_outputs(8986);
    layer2_outputs(3636) <= not(layer1_outputs(11253));
    layer2_outputs(3637) <= not((layer1_outputs(8657)) or (layer1_outputs(7622)));
    layer2_outputs(3638) <= layer1_outputs(5149);
    layer2_outputs(3639) <= layer1_outputs(2249);
    layer2_outputs(3640) <= not((layer1_outputs(4918)) and (layer1_outputs(10083)));
    layer2_outputs(3641) <= (layer1_outputs(10261)) and (layer1_outputs(10878));
    layer2_outputs(3642) <= layer1_outputs(392);
    layer2_outputs(3643) <= not(layer1_outputs(7501));
    layer2_outputs(3644) <= not((layer1_outputs(3360)) and (layer1_outputs(5569)));
    layer2_outputs(3645) <= not(layer1_outputs(4828));
    layer2_outputs(3646) <= not(layer1_outputs(1114)) or (layer1_outputs(6883));
    layer2_outputs(3647) <= layer1_outputs(4326);
    layer2_outputs(3648) <= layer1_outputs(10836);
    layer2_outputs(3649) <= not(layer1_outputs(4526));
    layer2_outputs(3650) <= layer1_outputs(1503);
    layer2_outputs(3651) <= not(layer1_outputs(8610));
    layer2_outputs(3652) <= layer1_outputs(9407);
    layer2_outputs(3653) <= (layer1_outputs(11199)) xor (layer1_outputs(10925));
    layer2_outputs(3654) <= layer1_outputs(44);
    layer2_outputs(3655) <= not(layer1_outputs(960));
    layer2_outputs(3656) <= not(layer1_outputs(10398));
    layer2_outputs(3657) <= not(layer1_outputs(255));
    layer2_outputs(3658) <= not(layer1_outputs(5299));
    layer2_outputs(3659) <= layer1_outputs(48);
    layer2_outputs(3660) <= (layer1_outputs(7540)) and not (layer1_outputs(8265));
    layer2_outputs(3661) <= not(layer1_outputs(12025));
    layer2_outputs(3662) <= (layer1_outputs(3967)) and not (layer1_outputs(192));
    layer2_outputs(3663) <= not((layer1_outputs(5698)) and (layer1_outputs(5161)));
    layer2_outputs(3664) <= not((layer1_outputs(1825)) or (layer1_outputs(8523)));
    layer2_outputs(3665) <= (layer1_outputs(9430)) and not (layer1_outputs(1793));
    layer2_outputs(3666) <= (layer1_outputs(3412)) or (layer1_outputs(7340));
    layer2_outputs(3667) <= layer1_outputs(7346);
    layer2_outputs(3668) <= not((layer1_outputs(8307)) xor (layer1_outputs(5227)));
    layer2_outputs(3669) <= layer1_outputs(10884);
    layer2_outputs(3670) <= not((layer1_outputs(5601)) and (layer1_outputs(5860)));
    layer2_outputs(3671) <= not((layer1_outputs(9487)) xor (layer1_outputs(10974)));
    layer2_outputs(3672) <= not((layer1_outputs(11748)) or (layer1_outputs(4957)));
    layer2_outputs(3673) <= layer1_outputs(9867);
    layer2_outputs(3674) <= not(layer1_outputs(4797)) or (layer1_outputs(891));
    layer2_outputs(3675) <= not(layer1_outputs(8376)) or (layer1_outputs(5614));
    layer2_outputs(3676) <= not((layer1_outputs(10554)) and (layer1_outputs(8237)));
    layer2_outputs(3677) <= '0';
    layer2_outputs(3678) <= layer1_outputs(10441);
    layer2_outputs(3679) <= (layer1_outputs(10514)) and not (layer1_outputs(506));
    layer2_outputs(3680) <= layer1_outputs(7273);
    layer2_outputs(3681) <= layer1_outputs(5955);
    layer2_outputs(3682) <= (layer1_outputs(12311)) and (layer1_outputs(11056));
    layer2_outputs(3683) <= (layer1_outputs(3766)) xor (layer1_outputs(4251));
    layer2_outputs(3684) <= layer1_outputs(3432);
    layer2_outputs(3685) <= (layer1_outputs(10254)) and (layer1_outputs(1938));
    layer2_outputs(3686) <= not(layer1_outputs(6268));
    layer2_outputs(3687) <= not(layer1_outputs(10727));
    layer2_outputs(3688) <= not(layer1_outputs(6287));
    layer2_outputs(3689) <= (layer1_outputs(10863)) or (layer1_outputs(12772));
    layer2_outputs(3690) <= not(layer1_outputs(10696)) or (layer1_outputs(2879));
    layer2_outputs(3691) <= not(layer1_outputs(1925));
    layer2_outputs(3692) <= not(layer1_outputs(3431));
    layer2_outputs(3693) <= not(layer1_outputs(3687));
    layer2_outputs(3694) <= not(layer1_outputs(6547));
    layer2_outputs(3695) <= layer1_outputs(4773);
    layer2_outputs(3696) <= layer1_outputs(11913);
    layer2_outputs(3697) <= layer1_outputs(8511);
    layer2_outputs(3698) <= not(layer1_outputs(12206));
    layer2_outputs(3699) <= not(layer1_outputs(484));
    layer2_outputs(3700) <= layer1_outputs(2902);
    layer2_outputs(3701) <= not((layer1_outputs(11885)) xor (layer1_outputs(1242)));
    layer2_outputs(3702) <= (layer1_outputs(692)) or (layer1_outputs(4710));
    layer2_outputs(3703) <= (layer1_outputs(11356)) and not (layer1_outputs(1913));
    layer2_outputs(3704) <= layer1_outputs(5926);
    layer2_outputs(3705) <= not(layer1_outputs(4964));
    layer2_outputs(3706) <= not((layer1_outputs(470)) or (layer1_outputs(3181)));
    layer2_outputs(3707) <= layer1_outputs(9315);
    layer2_outputs(3708) <= not(layer1_outputs(10544));
    layer2_outputs(3709) <= layer1_outputs(4601);
    layer2_outputs(3710) <= (layer1_outputs(6308)) and not (layer1_outputs(3137));
    layer2_outputs(3711) <= not(layer1_outputs(425)) or (layer1_outputs(3692));
    layer2_outputs(3712) <= not((layer1_outputs(1526)) or (layer1_outputs(7084)));
    layer2_outputs(3713) <= layer1_outputs(9405);
    layer2_outputs(3714) <= not((layer1_outputs(7588)) or (layer1_outputs(12784)));
    layer2_outputs(3715) <= not(layer1_outputs(1821));
    layer2_outputs(3716) <= (layer1_outputs(5455)) xor (layer1_outputs(12668));
    layer2_outputs(3717) <= (layer1_outputs(6043)) xor (layer1_outputs(259));
    layer2_outputs(3718) <= (layer1_outputs(4754)) and (layer1_outputs(7844));
    layer2_outputs(3719) <= (layer1_outputs(4850)) or (layer1_outputs(7655));
    layer2_outputs(3720) <= not((layer1_outputs(5201)) xor (layer1_outputs(6027)));
    layer2_outputs(3721) <= not((layer1_outputs(8684)) and (layer1_outputs(5957)));
    layer2_outputs(3722) <= not(layer1_outputs(2030));
    layer2_outputs(3723) <= layer1_outputs(4739);
    layer2_outputs(3724) <= not(layer1_outputs(7079));
    layer2_outputs(3725) <= (layer1_outputs(275)) and not (layer1_outputs(8385));
    layer2_outputs(3726) <= (layer1_outputs(10158)) xor (layer1_outputs(11403));
    layer2_outputs(3727) <= not(layer1_outputs(10013));
    layer2_outputs(3728) <= not(layer1_outputs(4808));
    layer2_outputs(3729) <= layer1_outputs(2559);
    layer2_outputs(3730) <= not((layer1_outputs(10375)) xor (layer1_outputs(9156)));
    layer2_outputs(3731) <= layer1_outputs(4033);
    layer2_outputs(3732) <= layer1_outputs(8414);
    layer2_outputs(3733) <= (layer1_outputs(646)) and not (layer1_outputs(5287));
    layer2_outputs(3734) <= not((layer1_outputs(12200)) xor (layer1_outputs(5297)));
    layer2_outputs(3735) <= (layer1_outputs(3443)) and (layer1_outputs(1948));
    layer2_outputs(3736) <= (layer1_outputs(2155)) and not (layer1_outputs(4795));
    layer2_outputs(3737) <= not((layer1_outputs(7959)) or (layer1_outputs(3027)));
    layer2_outputs(3738) <= not(layer1_outputs(3832));
    layer2_outputs(3739) <= (layer1_outputs(10477)) xor (layer1_outputs(7193));
    layer2_outputs(3740) <= not(layer1_outputs(3554));
    layer2_outputs(3741) <= not((layer1_outputs(10337)) and (layer1_outputs(11446)));
    layer2_outputs(3742) <= layer1_outputs(7532);
    layer2_outputs(3743) <= layer1_outputs(3119);
    layer2_outputs(3744) <= (layer1_outputs(11874)) or (layer1_outputs(916));
    layer2_outputs(3745) <= not(layer1_outputs(2364));
    layer2_outputs(3746) <= (layer1_outputs(2347)) and not (layer1_outputs(137));
    layer2_outputs(3747) <= not(layer1_outputs(2566));
    layer2_outputs(3748) <= not((layer1_outputs(9000)) xor (layer1_outputs(6694)));
    layer2_outputs(3749) <= (layer1_outputs(2915)) and not (layer1_outputs(10629));
    layer2_outputs(3750) <= layer1_outputs(6254);
    layer2_outputs(3751) <= not(layer1_outputs(7802)) or (layer1_outputs(6057));
    layer2_outputs(3752) <= (layer1_outputs(3838)) xor (layer1_outputs(4955));
    layer2_outputs(3753) <= (layer1_outputs(1814)) or (layer1_outputs(11050));
    layer2_outputs(3754) <= not(layer1_outputs(1024));
    layer2_outputs(3755) <= (layer1_outputs(5796)) and not (layer1_outputs(9973));
    layer2_outputs(3756) <= not((layer1_outputs(814)) or (layer1_outputs(11686)));
    layer2_outputs(3757) <= (layer1_outputs(5627)) and not (layer1_outputs(1761));
    layer2_outputs(3758) <= layer1_outputs(10755);
    layer2_outputs(3759) <= (layer1_outputs(3983)) xor (layer1_outputs(2269));
    layer2_outputs(3760) <= not(layer1_outputs(1924));
    layer2_outputs(3761) <= not(layer1_outputs(11131)) or (layer1_outputs(11388));
    layer2_outputs(3762) <= (layer1_outputs(4870)) and (layer1_outputs(5824));
    layer2_outputs(3763) <= not(layer1_outputs(8693));
    layer2_outputs(3764) <= (layer1_outputs(8702)) or (layer1_outputs(3848));
    layer2_outputs(3765) <= not(layer1_outputs(6748));
    layer2_outputs(3766) <= (layer1_outputs(534)) and not (layer1_outputs(5468));
    layer2_outputs(3767) <= layer1_outputs(8589);
    layer2_outputs(3768) <= not((layer1_outputs(7081)) xor (layer1_outputs(10239)));
    layer2_outputs(3769) <= not(layer1_outputs(5146)) or (layer1_outputs(2624));
    layer2_outputs(3770) <= layer1_outputs(6981);
    layer2_outputs(3771) <= layer1_outputs(10821);
    layer2_outputs(3772) <= (layer1_outputs(5295)) xor (layer1_outputs(11813));
    layer2_outputs(3773) <= layer1_outputs(10176);
    layer2_outputs(3774) <= layer1_outputs(1085);
    layer2_outputs(3775) <= (layer1_outputs(8148)) and (layer1_outputs(12480));
    layer2_outputs(3776) <= (layer1_outputs(9098)) xor (layer1_outputs(5811));
    layer2_outputs(3777) <= layer1_outputs(7386);
    layer2_outputs(3778) <= (layer1_outputs(1652)) and not (layer1_outputs(6471));
    layer2_outputs(3779) <= not(layer1_outputs(11382)) or (layer1_outputs(8345));
    layer2_outputs(3780) <= not((layer1_outputs(9534)) or (layer1_outputs(3579)));
    layer2_outputs(3781) <= layer1_outputs(6659);
    layer2_outputs(3782) <= layer1_outputs(1140);
    layer2_outputs(3783) <= not(layer1_outputs(8884));
    layer2_outputs(3784) <= (layer1_outputs(7451)) and (layer1_outputs(1744));
    layer2_outputs(3785) <= not(layer1_outputs(6830));
    layer2_outputs(3786) <= layer1_outputs(9331);
    layer2_outputs(3787) <= layer1_outputs(4876);
    layer2_outputs(3788) <= not(layer1_outputs(11256));
    layer2_outputs(3789) <= (layer1_outputs(3127)) and not (layer1_outputs(5089));
    layer2_outputs(3790) <= (layer1_outputs(6431)) xor (layer1_outputs(7541));
    layer2_outputs(3791) <= (layer1_outputs(3777)) and (layer1_outputs(9750));
    layer2_outputs(3792) <= not((layer1_outputs(8228)) xor (layer1_outputs(11949)));
    layer2_outputs(3793) <= not(layer1_outputs(10679)) or (layer1_outputs(9952));
    layer2_outputs(3794) <= not(layer1_outputs(12613));
    layer2_outputs(3795) <= not((layer1_outputs(5938)) and (layer1_outputs(3807)));
    layer2_outputs(3796) <= not(layer1_outputs(10549));
    layer2_outputs(3797) <= not(layer1_outputs(2547));
    layer2_outputs(3798) <= not(layer1_outputs(7555));
    layer2_outputs(3799) <= layer1_outputs(4570);
    layer2_outputs(3800) <= layer1_outputs(10431);
    layer2_outputs(3801) <= layer1_outputs(11808);
    layer2_outputs(3802) <= layer1_outputs(6572);
    layer2_outputs(3803) <= not(layer1_outputs(3040));
    layer2_outputs(3804) <= layer1_outputs(10038);
    layer2_outputs(3805) <= not((layer1_outputs(3818)) xor (layer1_outputs(10130)));
    layer2_outputs(3806) <= not((layer1_outputs(1582)) or (layer1_outputs(5103)));
    layer2_outputs(3807) <= not(layer1_outputs(4575)) or (layer1_outputs(5970));
    layer2_outputs(3808) <= (layer1_outputs(2163)) and (layer1_outputs(7815));
    layer2_outputs(3809) <= (layer1_outputs(3541)) xor (layer1_outputs(10510));
    layer2_outputs(3810) <= not(layer1_outputs(10538));
    layer2_outputs(3811) <= not((layer1_outputs(9368)) or (layer1_outputs(466)));
    layer2_outputs(3812) <= not(layer1_outputs(1044)) or (layer1_outputs(6069));
    layer2_outputs(3813) <= not((layer1_outputs(12170)) and (layer1_outputs(7269)));
    layer2_outputs(3814) <= not(layer1_outputs(85));
    layer2_outputs(3815) <= (layer1_outputs(2118)) and not (layer1_outputs(8188));
    layer2_outputs(3816) <= (layer1_outputs(6217)) and not (layer1_outputs(11529));
    layer2_outputs(3817) <= layer1_outputs(3864);
    layer2_outputs(3818) <= layer1_outputs(7086);
    layer2_outputs(3819) <= layer1_outputs(8673);
    layer2_outputs(3820) <= not((layer1_outputs(11037)) xor (layer1_outputs(2625)));
    layer2_outputs(3821) <= layer1_outputs(3937);
    layer2_outputs(3822) <= layer1_outputs(12532);
    layer2_outputs(3823) <= (layer1_outputs(10709)) and not (layer1_outputs(2909));
    layer2_outputs(3824) <= not(layer1_outputs(6437)) or (layer1_outputs(7200));
    layer2_outputs(3825) <= not(layer1_outputs(586));
    layer2_outputs(3826) <= not(layer1_outputs(2710)) or (layer1_outputs(6591));
    layer2_outputs(3827) <= not(layer1_outputs(1040)) or (layer1_outputs(9412));
    layer2_outputs(3828) <= not((layer1_outputs(11769)) or (layer1_outputs(9848)));
    layer2_outputs(3829) <= not(layer1_outputs(4525)) or (layer1_outputs(11883));
    layer2_outputs(3830) <= (layer1_outputs(11734)) xor (layer1_outputs(4079));
    layer2_outputs(3831) <= '0';
    layer2_outputs(3832) <= (layer1_outputs(2445)) and (layer1_outputs(9661));
    layer2_outputs(3833) <= not(layer1_outputs(6793));
    layer2_outputs(3834) <= not(layer1_outputs(10290));
    layer2_outputs(3835) <= layer1_outputs(1031);
    layer2_outputs(3836) <= not(layer1_outputs(11341));
    layer2_outputs(3837) <= not((layer1_outputs(2344)) and (layer1_outputs(2613)));
    layer2_outputs(3838) <= not(layer1_outputs(11441));
    layer2_outputs(3839) <= layer1_outputs(10715);
    layer2_outputs(3840) <= (layer1_outputs(2352)) and not (layer1_outputs(4066));
    layer2_outputs(3841) <= (layer1_outputs(5427)) xor (layer1_outputs(7387));
    layer2_outputs(3842) <= not(layer1_outputs(8246));
    layer2_outputs(3843) <= not(layer1_outputs(3644));
    layer2_outputs(3844) <= layer1_outputs(12000);
    layer2_outputs(3845) <= (layer1_outputs(5754)) xor (layer1_outputs(5968));
    layer2_outputs(3846) <= not(layer1_outputs(9826));
    layer2_outputs(3847) <= '1';
    layer2_outputs(3848) <= (layer1_outputs(4132)) xor (layer1_outputs(10145));
    layer2_outputs(3849) <= not(layer1_outputs(920));
    layer2_outputs(3850) <= (layer1_outputs(4198)) and (layer1_outputs(7057));
    layer2_outputs(3851) <= not(layer1_outputs(7873)) or (layer1_outputs(1737));
    layer2_outputs(3852) <= not(layer1_outputs(10911));
    layer2_outputs(3853) <= not((layer1_outputs(8736)) or (layer1_outputs(11987)));
    layer2_outputs(3854) <= not((layer1_outputs(2832)) xor (layer1_outputs(4803)));
    layer2_outputs(3855) <= (layer1_outputs(1799)) or (layer1_outputs(10307));
    layer2_outputs(3856) <= not(layer1_outputs(2531));
    layer2_outputs(3857) <= layer1_outputs(10762);
    layer2_outputs(3858) <= not(layer1_outputs(7952));
    layer2_outputs(3859) <= not(layer1_outputs(6489));
    layer2_outputs(3860) <= not(layer1_outputs(1456));
    layer2_outputs(3861) <= not((layer1_outputs(5827)) and (layer1_outputs(12398)));
    layer2_outputs(3862) <= not(layer1_outputs(10760));
    layer2_outputs(3863) <= layer1_outputs(5214);
    layer2_outputs(3864) <= layer1_outputs(9306);
    layer2_outputs(3865) <= layer1_outputs(9613);
    layer2_outputs(3866) <= (layer1_outputs(12458)) or (layer1_outputs(6825));
    layer2_outputs(3867) <= layer1_outputs(4289);
    layer2_outputs(3868) <= not(layer1_outputs(3700));
    layer2_outputs(3869) <= not(layer1_outputs(12680));
    layer2_outputs(3870) <= not((layer1_outputs(6032)) xor (layer1_outputs(11248)));
    layer2_outputs(3871) <= not((layer1_outputs(3263)) xor (layer1_outputs(7167)));
    layer2_outputs(3872) <= not(layer1_outputs(11));
    layer2_outputs(3873) <= not(layer1_outputs(9284));
    layer2_outputs(3874) <= not(layer1_outputs(9036));
    layer2_outputs(3875) <= not((layer1_outputs(8819)) or (layer1_outputs(6526)));
    layer2_outputs(3876) <= (layer1_outputs(6971)) xor (layer1_outputs(3683));
    layer2_outputs(3877) <= (layer1_outputs(3433)) xor (layer1_outputs(2266));
    layer2_outputs(3878) <= not(layer1_outputs(973));
    layer2_outputs(3879) <= (layer1_outputs(1117)) or (layer1_outputs(1125));
    layer2_outputs(3880) <= not((layer1_outputs(3383)) xor (layer1_outputs(5924)));
    layer2_outputs(3881) <= (layer1_outputs(4940)) and not (layer1_outputs(4303));
    layer2_outputs(3882) <= layer1_outputs(10088);
    layer2_outputs(3883) <= layer1_outputs(155);
    layer2_outputs(3884) <= not((layer1_outputs(4292)) and (layer1_outputs(8614)));
    layer2_outputs(3885) <= not((layer1_outputs(4862)) and (layer1_outputs(4526)));
    layer2_outputs(3886) <= not(layer1_outputs(7847));
    layer2_outputs(3887) <= not((layer1_outputs(7641)) or (layer1_outputs(3569)));
    layer2_outputs(3888) <= (layer1_outputs(5355)) xor (layer1_outputs(5027));
    layer2_outputs(3889) <= not(layer1_outputs(7566)) or (layer1_outputs(1263));
    layer2_outputs(3890) <= layer1_outputs(5721);
    layer2_outputs(3891) <= not((layer1_outputs(4734)) or (layer1_outputs(3667)));
    layer2_outputs(3892) <= not(layer1_outputs(2316));
    layer2_outputs(3893) <= (layer1_outputs(5057)) and not (layer1_outputs(4806));
    layer2_outputs(3894) <= layer1_outputs(7043);
    layer2_outputs(3895) <= layer1_outputs(10266);
    layer2_outputs(3896) <= (layer1_outputs(9969)) xor (layer1_outputs(2853));
    layer2_outputs(3897) <= not(layer1_outputs(3649));
    layer2_outputs(3898) <= not(layer1_outputs(768));
    layer2_outputs(3899) <= not((layer1_outputs(11545)) xor (layer1_outputs(9856)));
    layer2_outputs(3900) <= (layer1_outputs(9250)) or (layer1_outputs(947));
    layer2_outputs(3901) <= not(layer1_outputs(4531));
    layer2_outputs(3902) <= not((layer1_outputs(4193)) xor (layer1_outputs(6105)));
    layer2_outputs(3903) <= not(layer1_outputs(4414));
    layer2_outputs(3904) <= not(layer1_outputs(9378));
    layer2_outputs(3905) <= not((layer1_outputs(9610)) xor (layer1_outputs(2979)));
    layer2_outputs(3906) <= not(layer1_outputs(12453));
    layer2_outputs(3907) <= not((layer1_outputs(3655)) xor (layer1_outputs(10229)));
    layer2_outputs(3908) <= not(layer1_outputs(8421)) or (layer1_outputs(5802));
    layer2_outputs(3909) <= (layer1_outputs(4017)) or (layer1_outputs(11524));
    layer2_outputs(3910) <= not((layer1_outputs(5842)) xor (layer1_outputs(4264)));
    layer2_outputs(3911) <= not(layer1_outputs(397));
    layer2_outputs(3912) <= '1';
    layer2_outputs(3913) <= (layer1_outputs(8436)) xor (layer1_outputs(532));
    layer2_outputs(3914) <= layer1_outputs(10591);
    layer2_outputs(3915) <= not(layer1_outputs(9842));
    layer2_outputs(3916) <= layer1_outputs(9532);
    layer2_outputs(3917) <= not(layer1_outputs(1735));
    layer2_outputs(3918) <= not(layer1_outputs(4308)) or (layer1_outputs(5065));
    layer2_outputs(3919) <= not(layer1_outputs(541)) or (layer1_outputs(10476));
    layer2_outputs(3920) <= layer1_outputs(682);
    layer2_outputs(3921) <= (layer1_outputs(8133)) and (layer1_outputs(4472));
    layer2_outputs(3922) <= not(layer1_outputs(12207));
    layer2_outputs(3923) <= not(layer1_outputs(9653));
    layer2_outputs(3924) <= not(layer1_outputs(7509));
    layer2_outputs(3925) <= not(layer1_outputs(12715));
    layer2_outputs(3926) <= not((layer1_outputs(12725)) or (layer1_outputs(9376)));
    layer2_outputs(3927) <= not(layer1_outputs(12641));
    layer2_outputs(3928) <= layer1_outputs(5050);
    layer2_outputs(3929) <= (layer1_outputs(8051)) or (layer1_outputs(7790));
    layer2_outputs(3930) <= not((layer1_outputs(930)) xor (layer1_outputs(12076)));
    layer2_outputs(3931) <= not((layer1_outputs(10019)) or (layer1_outputs(4678)));
    layer2_outputs(3932) <= not(layer1_outputs(9078));
    layer2_outputs(3933) <= layer1_outputs(4003);
    layer2_outputs(3934) <= not(layer1_outputs(2963)) or (layer1_outputs(11337));
    layer2_outputs(3935) <= (layer1_outputs(2391)) and not (layer1_outputs(5272));
    layer2_outputs(3936) <= layer1_outputs(983);
    layer2_outputs(3937) <= (layer1_outputs(6205)) and not (layer1_outputs(3707));
    layer2_outputs(3938) <= not((layer1_outputs(3510)) or (layer1_outputs(7287)));
    layer2_outputs(3939) <= layer1_outputs(199);
    layer2_outputs(3940) <= not((layer1_outputs(5374)) and (layer1_outputs(152)));
    layer2_outputs(3941) <= not(layer1_outputs(2482));
    layer2_outputs(3942) <= not((layer1_outputs(2587)) xor (layer1_outputs(3784)));
    layer2_outputs(3943) <= not(layer1_outputs(2919));
    layer2_outputs(3944) <= not(layer1_outputs(1576));
    layer2_outputs(3945) <= layer1_outputs(4206);
    layer2_outputs(3946) <= not(layer1_outputs(10103));
    layer2_outputs(3947) <= layer1_outputs(927);
    layer2_outputs(3948) <= not(layer1_outputs(2405));
    layer2_outputs(3949) <= not(layer1_outputs(2324)) or (layer1_outputs(638));
    layer2_outputs(3950) <= '1';
    layer2_outputs(3951) <= '0';
    layer2_outputs(3952) <= not(layer1_outputs(4682));
    layer2_outputs(3953) <= not(layer1_outputs(5025)) or (layer1_outputs(5584));
    layer2_outputs(3954) <= not(layer1_outputs(4459)) or (layer1_outputs(5438));
    layer2_outputs(3955) <= not((layer1_outputs(8000)) or (layer1_outputs(9500)));
    layer2_outputs(3956) <= not((layer1_outputs(98)) xor (layer1_outputs(10198)));
    layer2_outputs(3957) <= not(layer1_outputs(1203));
    layer2_outputs(3958) <= not(layer1_outputs(8829));
    layer2_outputs(3959) <= not(layer1_outputs(10427)) or (layer1_outputs(5211));
    layer2_outputs(3960) <= not((layer1_outputs(322)) or (layer1_outputs(9795)));
    layer2_outputs(3961) <= (layer1_outputs(1887)) xor (layer1_outputs(11567));
    layer2_outputs(3962) <= not(layer1_outputs(362)) or (layer1_outputs(3275));
    layer2_outputs(3963) <= (layer1_outputs(3107)) and not (layer1_outputs(886));
    layer2_outputs(3964) <= (layer1_outputs(11810)) and not (layer1_outputs(2143));
    layer2_outputs(3965) <= not((layer1_outputs(10624)) xor (layer1_outputs(6833)));
    layer2_outputs(3966) <= not((layer1_outputs(11117)) xor (layer1_outputs(11238)));
    layer2_outputs(3967) <= not(layer1_outputs(5581)) or (layer1_outputs(7753));
    layer2_outputs(3968) <= (layer1_outputs(1748)) or (layer1_outputs(4450));
    layer2_outputs(3969) <= not(layer1_outputs(4409));
    layer2_outputs(3970) <= (layer1_outputs(2119)) and (layer1_outputs(1813));
    layer2_outputs(3971) <= (layer1_outputs(202)) and not (layer1_outputs(9067));
    layer2_outputs(3972) <= not(layer1_outputs(12044));
    layer2_outputs(3973) <= layer1_outputs(7124);
    layer2_outputs(3974) <= (layer1_outputs(7979)) and not (layer1_outputs(1488));
    layer2_outputs(3975) <= not(layer1_outputs(10336));
    layer2_outputs(3976) <= not(layer1_outputs(8130));
    layer2_outputs(3977) <= layer1_outputs(5644);
    layer2_outputs(3978) <= not(layer1_outputs(3754)) or (layer1_outputs(822));
    layer2_outputs(3979) <= not(layer1_outputs(10416));
    layer2_outputs(3980) <= not((layer1_outputs(12376)) and (layer1_outputs(5559)));
    layer2_outputs(3981) <= layer1_outputs(293);
    layer2_outputs(3982) <= layer1_outputs(8807);
    layer2_outputs(3983) <= layer1_outputs(6214);
    layer2_outputs(3984) <= layer1_outputs(5656);
    layer2_outputs(3985) <= not((layer1_outputs(3627)) xor (layer1_outputs(2865)));
    layer2_outputs(3986) <= layer1_outputs(7443);
    layer2_outputs(3987) <= not((layer1_outputs(6942)) xor (layer1_outputs(12734)));
    layer2_outputs(3988) <= (layer1_outputs(5266)) xor (layer1_outputs(6260));
    layer2_outputs(3989) <= not(layer1_outputs(10487));
    layer2_outputs(3990) <= (layer1_outputs(8544)) or (layer1_outputs(2149));
    layer2_outputs(3991) <= not(layer1_outputs(10467));
    layer2_outputs(3992) <= layer1_outputs(5967);
    layer2_outputs(3993) <= (layer1_outputs(1886)) xor (layer1_outputs(5880));
    layer2_outputs(3994) <= not(layer1_outputs(263));
    layer2_outputs(3995) <= (layer1_outputs(10012)) xor (layer1_outputs(1599));
    layer2_outputs(3996) <= not(layer1_outputs(1375)) or (layer1_outputs(3131));
    layer2_outputs(3997) <= layer1_outputs(2891);
    layer2_outputs(3998) <= not(layer1_outputs(10574));
    layer2_outputs(3999) <= layer1_outputs(6841);
    layer2_outputs(4000) <= not(layer1_outputs(1387)) or (layer1_outputs(5107));
    layer2_outputs(4001) <= not(layer1_outputs(808));
    layer2_outputs(4002) <= layer1_outputs(8920);
    layer2_outputs(4003) <= (layer1_outputs(1570)) or (layer1_outputs(7677));
    layer2_outputs(4004) <= layer1_outputs(3382);
    layer2_outputs(4005) <= not(layer1_outputs(2468));
    layer2_outputs(4006) <= not((layer1_outputs(9477)) and (layer1_outputs(2878)));
    layer2_outputs(4007) <= not(layer1_outputs(8745));
    layer2_outputs(4008) <= layer1_outputs(8356);
    layer2_outputs(4009) <= layer1_outputs(2546);
    layer2_outputs(4010) <= layer1_outputs(1036);
    layer2_outputs(4011) <= not(layer1_outputs(3899));
    layer2_outputs(4012) <= not(layer1_outputs(764));
    layer2_outputs(4013) <= (layer1_outputs(7915)) xor (layer1_outputs(2079));
    layer2_outputs(4014) <= not(layer1_outputs(5656)) or (layer1_outputs(6183));
    layer2_outputs(4015) <= not(layer1_outputs(6757)) or (layer1_outputs(4998));
    layer2_outputs(4016) <= not((layer1_outputs(10875)) xor (layer1_outputs(1077)));
    layer2_outputs(4017) <= not((layer1_outputs(1369)) and (layer1_outputs(8616)));
    layer2_outputs(4018) <= not(layer1_outputs(9370));
    layer2_outputs(4019) <= (layer1_outputs(10018)) and (layer1_outputs(511));
    layer2_outputs(4020) <= not(layer1_outputs(3671));
    layer2_outputs(4021) <= not(layer1_outputs(2385));
    layer2_outputs(4022) <= not(layer1_outputs(6866));
    layer2_outputs(4023) <= not((layer1_outputs(4197)) xor (layer1_outputs(5792)));
    layer2_outputs(4024) <= layer1_outputs(6648);
    layer2_outputs(4025) <= not((layer1_outputs(738)) and (layer1_outputs(12339)));
    layer2_outputs(4026) <= layer1_outputs(3278);
    layer2_outputs(4027) <= not(layer1_outputs(1630));
    layer2_outputs(4028) <= layer1_outputs(892);
    layer2_outputs(4029) <= layer1_outputs(10033);
    layer2_outputs(4030) <= not(layer1_outputs(1569));
    layer2_outputs(4031) <= (layer1_outputs(5903)) or (layer1_outputs(1025));
    layer2_outputs(4032) <= (layer1_outputs(9442)) and not (layer1_outputs(12554));
    layer2_outputs(4033) <= not(layer1_outputs(4872));
    layer2_outputs(4034) <= not(layer1_outputs(1822));
    layer2_outputs(4035) <= layer1_outputs(722);
    layer2_outputs(4036) <= (layer1_outputs(795)) and (layer1_outputs(8571));
    layer2_outputs(4037) <= layer1_outputs(435);
    layer2_outputs(4038) <= not(layer1_outputs(11031)) or (layer1_outputs(1381));
    layer2_outputs(4039) <= not(layer1_outputs(10328));
    layer2_outputs(4040) <= (layer1_outputs(1292)) xor (layer1_outputs(2083));
    layer2_outputs(4041) <= not(layer1_outputs(4730));
    layer2_outputs(4042) <= not((layer1_outputs(11999)) and (layer1_outputs(7821)));
    layer2_outputs(4043) <= not(layer1_outputs(9693)) or (layer1_outputs(11911));
    layer2_outputs(4044) <= layer1_outputs(4695);
    layer2_outputs(4045) <= (layer1_outputs(9414)) xor (layer1_outputs(3110));
    layer2_outputs(4046) <= (layer1_outputs(6178)) or (layer1_outputs(1819));
    layer2_outputs(4047) <= (layer1_outputs(6125)) xor (layer1_outputs(9844));
    layer2_outputs(4048) <= not((layer1_outputs(428)) and (layer1_outputs(9623)));
    layer2_outputs(4049) <= not(layer1_outputs(3115));
    layer2_outputs(4050) <= not(layer1_outputs(4532));
    layer2_outputs(4051) <= (layer1_outputs(11006)) and not (layer1_outputs(4681));
    layer2_outputs(4052) <= not(layer1_outputs(10857));
    layer2_outputs(4053) <= (layer1_outputs(12247)) or (layer1_outputs(9114));
    layer2_outputs(4054) <= not(layer1_outputs(8458));
    layer2_outputs(4055) <= not((layer1_outputs(3353)) or (layer1_outputs(11331)));
    layer2_outputs(4056) <= not(layer1_outputs(12619)) or (layer1_outputs(6413));
    layer2_outputs(4057) <= layer1_outputs(1451);
    layer2_outputs(4058) <= not(layer1_outputs(10578));
    layer2_outputs(4059) <= not(layer1_outputs(9175));
    layer2_outputs(4060) <= not(layer1_outputs(2660));
    layer2_outputs(4061) <= not((layer1_outputs(9615)) xor (layer1_outputs(11225)));
    layer2_outputs(4062) <= not(layer1_outputs(5570));
    layer2_outputs(4063) <= not(layer1_outputs(11572));
    layer2_outputs(4064) <= not(layer1_outputs(7639)) or (layer1_outputs(8450));
    layer2_outputs(4065) <= (layer1_outputs(7507)) and not (layer1_outputs(1755));
    layer2_outputs(4066) <= not((layer1_outputs(9298)) or (layer1_outputs(12713)));
    layer2_outputs(4067) <= (layer1_outputs(9132)) xor (layer1_outputs(11717));
    layer2_outputs(4068) <= (layer1_outputs(1059)) or (layer1_outputs(6087));
    layer2_outputs(4069) <= layer1_outputs(8481);
    layer2_outputs(4070) <= layer1_outputs(229);
    layer2_outputs(4071) <= not((layer1_outputs(974)) or (layer1_outputs(10007)));
    layer2_outputs(4072) <= not(layer1_outputs(8118));
    layer2_outputs(4073) <= not(layer1_outputs(5580));
    layer2_outputs(4074) <= not((layer1_outputs(12380)) xor (layer1_outputs(12227)));
    layer2_outputs(4075) <= (layer1_outputs(5788)) or (layer1_outputs(8301));
    layer2_outputs(4076) <= layer1_outputs(2775);
    layer2_outputs(4077) <= layer1_outputs(840);
    layer2_outputs(4078) <= (layer1_outputs(6127)) and (layer1_outputs(2033));
    layer2_outputs(4079) <= (layer1_outputs(1155)) xor (layer1_outputs(12143));
    layer2_outputs(4080) <= not((layer1_outputs(1316)) xor (layer1_outputs(1468)));
    layer2_outputs(4081) <= (layer1_outputs(8213)) and (layer1_outputs(3725));
    layer2_outputs(4082) <= not((layer1_outputs(47)) and (layer1_outputs(3200)));
    layer2_outputs(4083) <= (layer1_outputs(2921)) and not (layer1_outputs(7763));
    layer2_outputs(4084) <= not(layer1_outputs(5780)) or (layer1_outputs(9361));
    layer2_outputs(4085) <= not((layer1_outputs(11)) or (layer1_outputs(8283)));
    layer2_outputs(4086) <= (layer1_outputs(8438)) xor (layer1_outputs(10744));
    layer2_outputs(4087) <= not(layer1_outputs(8682));
    layer2_outputs(4088) <= layer1_outputs(1011);
    layer2_outputs(4089) <= layer1_outputs(5204);
    layer2_outputs(4090) <= not((layer1_outputs(2003)) xor (layer1_outputs(3758)));
    layer2_outputs(4091) <= not((layer1_outputs(9300)) and (layer1_outputs(11839)));
    layer2_outputs(4092) <= not(layer1_outputs(4275));
    layer2_outputs(4093) <= '0';
    layer2_outputs(4094) <= not(layer1_outputs(6211));
    layer2_outputs(4095) <= layer1_outputs(3519);
    layer2_outputs(4096) <= not(layer1_outputs(11265)) or (layer1_outputs(4508));
    layer2_outputs(4097) <= not(layer1_outputs(8850));
    layer2_outputs(4098) <= layer1_outputs(4673);
    layer2_outputs(4099) <= not((layer1_outputs(1016)) and (layer1_outputs(12295)));
    layer2_outputs(4100) <= (layer1_outputs(2376)) and not (layer1_outputs(8577));
    layer2_outputs(4101) <= not((layer1_outputs(7231)) xor (layer1_outputs(4193)));
    layer2_outputs(4102) <= not(layer1_outputs(7277));
    layer2_outputs(4103) <= (layer1_outputs(3064)) and not (layer1_outputs(3718));
    layer2_outputs(4104) <= (layer1_outputs(2833)) xor (layer1_outputs(1862));
    layer2_outputs(4105) <= layer1_outputs(6786);
    layer2_outputs(4106) <= not(layer1_outputs(4170));
    layer2_outputs(4107) <= not(layer1_outputs(8340));
    layer2_outputs(4108) <= layer1_outputs(8324);
    layer2_outputs(4109) <= not((layer1_outputs(9615)) or (layer1_outputs(1834)));
    layer2_outputs(4110) <= not((layer1_outputs(12460)) and (layer1_outputs(2102)));
    layer2_outputs(4111) <= layer1_outputs(1333);
    layer2_outputs(4112) <= not(layer1_outputs(334)) or (layer1_outputs(512));
    layer2_outputs(4113) <= not((layer1_outputs(4862)) and (layer1_outputs(53)));
    layer2_outputs(4114) <= layer1_outputs(3717);
    layer2_outputs(4115) <= layer1_outputs(6732);
    layer2_outputs(4116) <= layer1_outputs(5172);
    layer2_outputs(4117) <= not(layer1_outputs(12744)) or (layer1_outputs(5940));
    layer2_outputs(4118) <= layer1_outputs(4323);
    layer2_outputs(4119) <= (layer1_outputs(5671)) xor (layer1_outputs(2814));
    layer2_outputs(4120) <= layer1_outputs(8096);
    layer2_outputs(4121) <= not(layer1_outputs(1019)) or (layer1_outputs(7966));
    layer2_outputs(4122) <= (layer1_outputs(11794)) and not (layer1_outputs(5361));
    layer2_outputs(4123) <= not((layer1_outputs(6534)) or (layer1_outputs(5359)));
    layer2_outputs(4124) <= '0';
    layer2_outputs(4125) <= (layer1_outputs(7056)) xor (layer1_outputs(1145));
    layer2_outputs(4126) <= not(layer1_outputs(470));
    layer2_outputs(4127) <= layer1_outputs(7880);
    layer2_outputs(4128) <= layer1_outputs(6402);
    layer2_outputs(4129) <= not(layer1_outputs(9697));
    layer2_outputs(4130) <= not(layer1_outputs(5291));
    layer2_outputs(4131) <= not(layer1_outputs(8018));
    layer2_outputs(4132) <= not((layer1_outputs(327)) xor (layer1_outputs(4835)));
    layer2_outputs(4133) <= layer1_outputs(2031);
    layer2_outputs(4134) <= layer1_outputs(3764);
    layer2_outputs(4135) <= not(layer1_outputs(3216));
    layer2_outputs(4136) <= not((layer1_outputs(114)) and (layer1_outputs(10810)));
    layer2_outputs(4137) <= not(layer1_outputs(50));
    layer2_outputs(4138) <= (layer1_outputs(4826)) xor (layer1_outputs(764));
    layer2_outputs(4139) <= (layer1_outputs(3558)) or (layer1_outputs(2688));
    layer2_outputs(4140) <= not(layer1_outputs(5854)) or (layer1_outputs(11980));
    layer2_outputs(4141) <= not((layer1_outputs(6704)) or (layer1_outputs(1400)));
    layer2_outputs(4142) <= not(layer1_outputs(2308)) or (layer1_outputs(3666));
    layer2_outputs(4143) <= not((layer1_outputs(1703)) and (layer1_outputs(2977)));
    layer2_outputs(4144) <= not((layer1_outputs(12681)) or (layer1_outputs(7770)));
    layer2_outputs(4145) <= (layer1_outputs(893)) or (layer1_outputs(234));
    layer2_outputs(4146) <= not((layer1_outputs(3143)) or (layer1_outputs(4993)));
    layer2_outputs(4147) <= not(layer1_outputs(8542)) or (layer1_outputs(1663));
    layer2_outputs(4148) <= (layer1_outputs(8745)) and (layer1_outputs(9888));
    layer2_outputs(4149) <= (layer1_outputs(1323)) or (layer1_outputs(7160));
    layer2_outputs(4150) <= layer1_outputs(10840);
    layer2_outputs(4151) <= layer1_outputs(208);
    layer2_outputs(4152) <= not(layer1_outputs(10367));
    layer2_outputs(4153) <= (layer1_outputs(10115)) or (layer1_outputs(1617));
    layer2_outputs(4154) <= not(layer1_outputs(9006));
    layer2_outputs(4155) <= layer1_outputs(1340);
    layer2_outputs(4156) <= not(layer1_outputs(10929));
    layer2_outputs(4157) <= layer1_outputs(2116);
    layer2_outputs(4158) <= not(layer1_outputs(12076));
    layer2_outputs(4159) <= not(layer1_outputs(1243)) or (layer1_outputs(5980));
    layer2_outputs(4160) <= not(layer1_outputs(9464));
    layer2_outputs(4161) <= not((layer1_outputs(11969)) or (layer1_outputs(4884)));
    layer2_outputs(4162) <= not(layer1_outputs(11315));
    layer2_outputs(4163) <= not(layer1_outputs(12026));
    layer2_outputs(4164) <= not(layer1_outputs(9854)) or (layer1_outputs(9024));
    layer2_outputs(4165) <= not(layer1_outputs(1007));
    layer2_outputs(4166) <= layer1_outputs(414);
    layer2_outputs(4167) <= (layer1_outputs(7023)) xor (layer1_outputs(265));
    layer2_outputs(4168) <= not(layer1_outputs(3065));
    layer2_outputs(4169) <= (layer1_outputs(1859)) and not (layer1_outputs(4671));
    layer2_outputs(4170) <= not((layer1_outputs(5574)) or (layer1_outputs(6633)));
    layer2_outputs(4171) <= not((layer1_outputs(9951)) or (layer1_outputs(6926)));
    layer2_outputs(4172) <= (layer1_outputs(28)) xor (layer1_outputs(5847));
    layer2_outputs(4173) <= layer1_outputs(11646);
    layer2_outputs(4174) <= not((layer1_outputs(3543)) xor (layer1_outputs(8713)));
    layer2_outputs(4175) <= not((layer1_outputs(3177)) xor (layer1_outputs(11228)));
    layer2_outputs(4176) <= (layer1_outputs(10367)) or (layer1_outputs(7005));
    layer2_outputs(4177) <= not(layer1_outputs(6465));
    layer2_outputs(4178) <= not(layer1_outputs(11786));
    layer2_outputs(4179) <= layer1_outputs(3830);
    layer2_outputs(4180) <= layer1_outputs(10804);
    layer2_outputs(4181) <= not((layer1_outputs(6611)) and (layer1_outputs(5076)));
    layer2_outputs(4182) <= (layer1_outputs(9815)) and (layer1_outputs(11848));
    layer2_outputs(4183) <= not(layer1_outputs(12211));
    layer2_outputs(4184) <= layer1_outputs(5984);
    layer2_outputs(4185) <= layer1_outputs(11633);
    layer2_outputs(4186) <= not(layer1_outputs(8602));
    layer2_outputs(4187) <= layer1_outputs(12384);
    layer2_outputs(4188) <= not(layer1_outputs(2404));
    layer2_outputs(4189) <= not(layer1_outputs(7545));
    layer2_outputs(4190) <= (layer1_outputs(4668)) xor (layer1_outputs(1845));
    layer2_outputs(4191) <= not(layer1_outputs(73));
    layer2_outputs(4192) <= (layer1_outputs(6753)) and (layer1_outputs(3503));
    layer2_outputs(4193) <= (layer1_outputs(3670)) and (layer1_outputs(11522));
    layer2_outputs(4194) <= not((layer1_outputs(7581)) and (layer1_outputs(8190)));
    layer2_outputs(4195) <= (layer1_outputs(4227)) and (layer1_outputs(10050));
    layer2_outputs(4196) <= (layer1_outputs(10302)) and (layer1_outputs(7081));
    layer2_outputs(4197) <= not(layer1_outputs(1412)) or (layer1_outputs(9859));
    layer2_outputs(4198) <= not(layer1_outputs(4336)) or (layer1_outputs(4896));
    layer2_outputs(4199) <= (layer1_outputs(8288)) and not (layer1_outputs(5409));
    layer2_outputs(4200) <= not(layer1_outputs(10494));
    layer2_outputs(4201) <= not(layer1_outputs(876)) or (layer1_outputs(11300));
    layer2_outputs(4202) <= not(layer1_outputs(5917));
    layer2_outputs(4203) <= layer1_outputs(11702);
    layer2_outputs(4204) <= layer1_outputs(2381);
    layer2_outputs(4205) <= layer1_outputs(1874);
    layer2_outputs(4206) <= layer1_outputs(12094);
    layer2_outputs(4207) <= not(layer1_outputs(2474));
    layer2_outputs(4208) <= (layer1_outputs(2653)) xor (layer1_outputs(8943));
    layer2_outputs(4209) <= (layer1_outputs(11367)) and not (layer1_outputs(4898));
    layer2_outputs(4210) <= layer1_outputs(306);
    layer2_outputs(4211) <= layer1_outputs(9383);
    layer2_outputs(4212) <= (layer1_outputs(4566)) and (layer1_outputs(4015));
    layer2_outputs(4213) <= not(layer1_outputs(11015)) or (layer1_outputs(9759));
    layer2_outputs(4214) <= layer1_outputs(9301);
    layer2_outputs(4215) <= (layer1_outputs(11210)) and (layer1_outputs(6031));
    layer2_outputs(4216) <= layer1_outputs(7985);
    layer2_outputs(4217) <= (layer1_outputs(11554)) and (layer1_outputs(658));
    layer2_outputs(4218) <= not(layer1_outputs(11321));
    layer2_outputs(4219) <= layer1_outputs(1029);
    layer2_outputs(4220) <= (layer1_outputs(7905)) or (layer1_outputs(9213));
    layer2_outputs(4221) <= layer1_outputs(6116);
    layer2_outputs(4222) <= not((layer1_outputs(8675)) xor (layer1_outputs(8904)));
    layer2_outputs(4223) <= not(layer1_outputs(8935));
    layer2_outputs(4224) <= layer1_outputs(12190);
    layer2_outputs(4225) <= not(layer1_outputs(12773)) or (layer1_outputs(5964));
    layer2_outputs(4226) <= (layer1_outputs(12106)) and not (layer1_outputs(12658));
    layer2_outputs(4227) <= layer1_outputs(6470);
    layer2_outputs(4228) <= not((layer1_outputs(10006)) xor (layer1_outputs(7164)));
    layer2_outputs(4229) <= layer1_outputs(9100);
    layer2_outputs(4230) <= not(layer1_outputs(11677));
    layer2_outputs(4231) <= (layer1_outputs(374)) or (layer1_outputs(6605));
    layer2_outputs(4232) <= layer1_outputs(7059);
    layer2_outputs(4233) <= layer1_outputs(1419);
    layer2_outputs(4234) <= not(layer1_outputs(3644));
    layer2_outputs(4235) <= (layer1_outputs(10397)) and not (layer1_outputs(6312));
    layer2_outputs(4236) <= layer1_outputs(5704);
    layer2_outputs(4237) <= not(layer1_outputs(9475)) or (layer1_outputs(6548));
    layer2_outputs(4238) <= not((layer1_outputs(11896)) xor (layer1_outputs(9051)));
    layer2_outputs(4239) <= not((layer1_outputs(7172)) xor (layer1_outputs(4429)));
    layer2_outputs(4240) <= (layer1_outputs(12166)) and (layer1_outputs(11690));
    layer2_outputs(4241) <= not(layer1_outputs(1127)) or (layer1_outputs(7162));
    layer2_outputs(4242) <= not(layer1_outputs(11730));
    layer2_outputs(4243) <= not(layer1_outputs(10116)) or (layer1_outputs(12346));
    layer2_outputs(4244) <= (layer1_outputs(11532)) xor (layer1_outputs(12134));
    layer2_outputs(4245) <= (layer1_outputs(4948)) or (layer1_outputs(12350));
    layer2_outputs(4246) <= (layer1_outputs(2159)) or (layer1_outputs(12191));
    layer2_outputs(4247) <= not(layer1_outputs(312)) or (layer1_outputs(8239));
    layer2_outputs(4248) <= not(layer1_outputs(3780));
    layer2_outputs(4249) <= (layer1_outputs(10726)) and (layer1_outputs(2068));
    layer2_outputs(4250) <= not(layer1_outputs(407)) or (layer1_outputs(10864));
    layer2_outputs(4251) <= not(layer1_outputs(5726)) or (layer1_outputs(4444));
    layer2_outputs(4252) <= (layer1_outputs(7980)) xor (layer1_outputs(1238));
    layer2_outputs(4253) <= not((layer1_outputs(3357)) and (layer1_outputs(12733)));
    layer2_outputs(4254) <= not((layer1_outputs(12706)) xor (layer1_outputs(828)));
    layer2_outputs(4255) <= not(layer1_outputs(12456));
    layer2_outputs(4256) <= not(layer1_outputs(8526));
    layer2_outputs(4257) <= (layer1_outputs(8643)) and not (layer1_outputs(11195));
    layer2_outputs(4258) <= not(layer1_outputs(6355)) or (layer1_outputs(6283));
    layer2_outputs(4259) <= (layer1_outputs(984)) and not (layer1_outputs(7800));
    layer2_outputs(4260) <= not((layer1_outputs(4083)) and (layer1_outputs(12713)));
    layer2_outputs(4261) <= (layer1_outputs(3203)) or (layer1_outputs(9578));
    layer2_outputs(4262) <= not(layer1_outputs(10030));
    layer2_outputs(4263) <= layer1_outputs(8473);
    layer2_outputs(4264) <= not((layer1_outputs(8377)) or (layer1_outputs(4081)));
    layer2_outputs(4265) <= layer1_outputs(10701);
    layer2_outputs(4266) <= not((layer1_outputs(6215)) or (layer1_outputs(8573)));
    layer2_outputs(4267) <= not((layer1_outputs(6662)) and (layer1_outputs(868)));
    layer2_outputs(4268) <= (layer1_outputs(7105)) and (layer1_outputs(10855));
    layer2_outputs(4269) <= not((layer1_outputs(7342)) xor (layer1_outputs(8651)));
    layer2_outputs(4270) <= layer1_outputs(436);
    layer2_outputs(4271) <= layer1_outputs(4538);
    layer2_outputs(4272) <= layer1_outputs(6876);
    layer2_outputs(4273) <= not(layer1_outputs(8743)) or (layer1_outputs(4576));
    layer2_outputs(4274) <= not((layer1_outputs(10533)) xor (layer1_outputs(2793)));
    layer2_outputs(4275) <= layer1_outputs(6954);
    layer2_outputs(4276) <= not((layer1_outputs(5912)) xor (layer1_outputs(5177)));
    layer2_outputs(4277) <= layer1_outputs(10);
    layer2_outputs(4278) <= (layer1_outputs(12305)) and not (layer1_outputs(2835));
    layer2_outputs(4279) <= layer1_outputs(6633);
    layer2_outputs(4280) <= layer1_outputs(1585);
    layer2_outputs(4281) <= not(layer1_outputs(4416));
    layer2_outputs(4282) <= layer1_outputs(8365);
    layer2_outputs(4283) <= not(layer1_outputs(11051));
    layer2_outputs(4284) <= not(layer1_outputs(1918));
    layer2_outputs(4285) <= (layer1_outputs(12612)) and not (layer1_outputs(5987));
    layer2_outputs(4286) <= (layer1_outputs(4373)) xor (layer1_outputs(1095));
    layer2_outputs(4287) <= not(layer1_outputs(9589));
    layer2_outputs(4288) <= layer1_outputs(3750);
    layer2_outputs(4289) <= layer1_outputs(2201);
    layer2_outputs(4290) <= (layer1_outputs(8160)) or (layer1_outputs(7030));
    layer2_outputs(4291) <= (layer1_outputs(1356)) or (layer1_outputs(9030));
    layer2_outputs(4292) <= not(layer1_outputs(6854)) or (layer1_outputs(6371));
    layer2_outputs(4293) <= not((layer1_outputs(6236)) or (layer1_outputs(6794)));
    layer2_outputs(4294) <= not((layer1_outputs(8985)) or (layer1_outputs(6924)));
    layer2_outputs(4295) <= layer1_outputs(6825);
    layer2_outputs(4296) <= not(layer1_outputs(12467)) or (layer1_outputs(12428));
    layer2_outputs(4297) <= not(layer1_outputs(3368)) or (layer1_outputs(357));
    layer2_outputs(4298) <= (layer1_outputs(12698)) xor (layer1_outputs(6455));
    layer2_outputs(4299) <= layer1_outputs(433);
    layer2_outputs(4300) <= not(layer1_outputs(10608));
    layer2_outputs(4301) <= not(layer1_outputs(1343));
    layer2_outputs(4302) <= (layer1_outputs(4023)) and not (layer1_outputs(7627));
    layer2_outputs(4303) <= not(layer1_outputs(1784)) or (layer1_outputs(7346));
    layer2_outputs(4304) <= not(layer1_outputs(9089)) or (layer1_outputs(9563));
    layer2_outputs(4305) <= layer1_outputs(825);
    layer2_outputs(4306) <= layer1_outputs(1891);
    layer2_outputs(4307) <= (layer1_outputs(6826)) and not (layer1_outputs(9029));
    layer2_outputs(4308) <= (layer1_outputs(3771)) and (layer1_outputs(11217));
    layer2_outputs(4309) <= not((layer1_outputs(8299)) and (layer1_outputs(9015)));
    layer2_outputs(4310) <= not((layer1_outputs(4714)) and (layer1_outputs(1391)));
    layer2_outputs(4311) <= not(layer1_outputs(440));
    layer2_outputs(4312) <= not(layer1_outputs(3680));
    layer2_outputs(4313) <= not(layer1_outputs(11537));
    layer2_outputs(4314) <= not((layer1_outputs(388)) xor (layer1_outputs(1882)));
    layer2_outputs(4315) <= layer1_outputs(7750);
    layer2_outputs(4316) <= not(layer1_outputs(12504));
    layer2_outputs(4317) <= layer1_outputs(7527);
    layer2_outputs(4318) <= layer1_outputs(11655);
    layer2_outputs(4319) <= not(layer1_outputs(10538)) or (layer1_outputs(2309));
    layer2_outputs(4320) <= not((layer1_outputs(12552)) xor (layer1_outputs(7198)));
    layer2_outputs(4321) <= (layer1_outputs(3948)) xor (layer1_outputs(4648));
    layer2_outputs(4322) <= not((layer1_outputs(4188)) and (layer1_outputs(11846)));
    layer2_outputs(4323) <= (layer1_outputs(5512)) and (layer1_outputs(10298));
    layer2_outputs(4324) <= not((layer1_outputs(4873)) or (layer1_outputs(1894)));
    layer2_outputs(4325) <= (layer1_outputs(6472)) or (layer1_outputs(3951));
    layer2_outputs(4326) <= not(layer1_outputs(11000));
    layer2_outputs(4327) <= not(layer1_outputs(12761));
    layer2_outputs(4328) <= not(layer1_outputs(6796));
    layer2_outputs(4329) <= not((layer1_outputs(9595)) and (layer1_outputs(6286)));
    layer2_outputs(4330) <= not(layer1_outputs(8366));
    layer2_outputs(4331) <= not(layer1_outputs(10582));
    layer2_outputs(4332) <= (layer1_outputs(9635)) or (layer1_outputs(9841));
    layer2_outputs(4333) <= not((layer1_outputs(570)) and (layer1_outputs(5750)));
    layer2_outputs(4334) <= not(layer1_outputs(5314)) or (layer1_outputs(7891));
    layer2_outputs(4335) <= (layer1_outputs(7481)) and (layer1_outputs(9864));
    layer2_outputs(4336) <= not(layer1_outputs(63));
    layer2_outputs(4337) <= not((layer1_outputs(8818)) or (layer1_outputs(10190)));
    layer2_outputs(4338) <= not(layer1_outputs(9612));
    layer2_outputs(4339) <= layer1_outputs(7831);
    layer2_outputs(4340) <= (layer1_outputs(2196)) and not (layer1_outputs(2799));
    layer2_outputs(4341) <= (layer1_outputs(1356)) and (layer1_outputs(12330));
    layer2_outputs(4342) <= (layer1_outputs(1952)) xor (layer1_outputs(7189));
    layer2_outputs(4343) <= (layer1_outputs(1557)) or (layer1_outputs(1210));
    layer2_outputs(4344) <= (layer1_outputs(153)) and not (layer1_outputs(11763));
    layer2_outputs(4345) <= (layer1_outputs(11164)) xor (layer1_outputs(1466));
    layer2_outputs(4346) <= (layer1_outputs(4169)) and (layer1_outputs(5198));
    layer2_outputs(4347) <= not(layer1_outputs(11472));
    layer2_outputs(4348) <= not((layer1_outputs(12116)) and (layer1_outputs(4362)));
    layer2_outputs(4349) <= layer1_outputs(7500);
    layer2_outputs(4350) <= layer1_outputs(1782);
    layer2_outputs(4351) <= (layer1_outputs(266)) xor (layer1_outputs(12423));
    layer2_outputs(4352) <= not(layer1_outputs(6747));
    layer2_outputs(4353) <= not(layer1_outputs(5091));
    layer2_outputs(4354) <= not(layer1_outputs(6397)) or (layer1_outputs(1723));
    layer2_outputs(4355) <= not((layer1_outputs(10598)) xor (layer1_outputs(10996)));
    layer2_outputs(4356) <= not((layer1_outputs(8787)) or (layer1_outputs(296)));
    layer2_outputs(4357) <= layer1_outputs(11911);
    layer2_outputs(4358) <= layer1_outputs(11864);
    layer2_outputs(4359) <= not(layer1_outputs(8562));
    layer2_outputs(4360) <= layer1_outputs(4519);
    layer2_outputs(4361) <= not((layer1_outputs(10391)) or (layer1_outputs(7591)));
    layer2_outputs(4362) <= not((layer1_outputs(12016)) xor (layer1_outputs(11309)));
    layer2_outputs(4363) <= not((layer1_outputs(5391)) xor (layer1_outputs(399)));
    layer2_outputs(4364) <= not(layer1_outputs(10694)) or (layer1_outputs(11887));
    layer2_outputs(4365) <= layer1_outputs(8069);
    layer2_outputs(4366) <= not(layer1_outputs(11894));
    layer2_outputs(4367) <= not((layer1_outputs(10373)) or (layer1_outputs(3805)));
    layer2_outputs(4368) <= (layer1_outputs(794)) xor (layer1_outputs(8606));
    layer2_outputs(4369) <= (layer1_outputs(4393)) and not (layer1_outputs(11184));
    layer2_outputs(4370) <= not(layer1_outputs(9303));
    layer2_outputs(4371) <= (layer1_outputs(8869)) or (layer1_outputs(7118));
    layer2_outputs(4372) <= not(layer1_outputs(2130));
    layer2_outputs(4373) <= not((layer1_outputs(1527)) xor (layer1_outputs(1302)));
    layer2_outputs(4374) <= layer1_outputs(9732);
    layer2_outputs(4375) <= not(layer1_outputs(2796)) or (layer1_outputs(12079));
    layer2_outputs(4376) <= layer1_outputs(9283);
    layer2_outputs(4377) <= (layer1_outputs(10599)) or (layer1_outputs(8471));
    layer2_outputs(4378) <= layer1_outputs(7782);
    layer2_outputs(4379) <= not(layer1_outputs(9970));
    layer2_outputs(4380) <= (layer1_outputs(886)) or (layer1_outputs(9327));
    layer2_outputs(4381) <= layer1_outputs(483);
    layer2_outputs(4382) <= not(layer1_outputs(5537));
    layer2_outputs(4383) <= layer1_outputs(2355);
    layer2_outputs(4384) <= (layer1_outputs(11683)) and (layer1_outputs(11128));
    layer2_outputs(4385) <= layer1_outputs(8198);
    layer2_outputs(4386) <= not(layer1_outputs(3830)) or (layer1_outputs(1563));
    layer2_outputs(4387) <= (layer1_outputs(6066)) or (layer1_outputs(8280));
    layer2_outputs(4388) <= not(layer1_outputs(10204));
    layer2_outputs(4389) <= layer1_outputs(7674);
    layer2_outputs(4390) <= not(layer1_outputs(1134));
    layer2_outputs(4391) <= layer1_outputs(539);
    layer2_outputs(4392) <= (layer1_outputs(926)) and not (layer1_outputs(7067));
    layer2_outputs(4393) <= not(layer1_outputs(3257)) or (layer1_outputs(7024));
    layer2_outputs(4394) <= layer1_outputs(6106);
    layer2_outputs(4395) <= not((layer1_outputs(12472)) or (layer1_outputs(4555)));
    layer2_outputs(4396) <= (layer1_outputs(576)) and not (layer1_outputs(11306));
    layer2_outputs(4397) <= not(layer1_outputs(9865));
    layer2_outputs(4398) <= not(layer1_outputs(325));
    layer2_outputs(4399) <= layer1_outputs(7389);
    layer2_outputs(4400) <= not(layer1_outputs(6766));
    layer2_outputs(4401) <= layer1_outputs(5213);
    layer2_outputs(4402) <= not(layer1_outputs(1916)) or (layer1_outputs(5326));
    layer2_outputs(4403) <= not(layer1_outputs(10987));
    layer2_outputs(4404) <= '1';
    layer2_outputs(4405) <= layer1_outputs(6092);
    layer2_outputs(4406) <= not(layer1_outputs(8914)) or (layer1_outputs(10072));
    layer2_outputs(4407) <= not(layer1_outputs(9781));
    layer2_outputs(4408) <= (layer1_outputs(12719)) and not (layer1_outputs(1642));
    layer2_outputs(4409) <= (layer1_outputs(12236)) xor (layer1_outputs(6128));
    layer2_outputs(4410) <= not(layer1_outputs(1263));
    layer2_outputs(4411) <= layer1_outputs(6095);
    layer2_outputs(4412) <= layer1_outputs(6136);
    layer2_outputs(4413) <= '1';
    layer2_outputs(4414) <= '1';
    layer2_outputs(4415) <= not(layer1_outputs(5923)) or (layer1_outputs(12771));
    layer2_outputs(4416) <= (layer1_outputs(3435)) and not (layer1_outputs(7117));
    layer2_outputs(4417) <= layer1_outputs(10380);
    layer2_outputs(4418) <= layer1_outputs(5281);
    layer2_outputs(4419) <= (layer1_outputs(2150)) xor (layer1_outputs(216));
    layer2_outputs(4420) <= layer1_outputs(2872);
    layer2_outputs(4421) <= not(layer1_outputs(1429));
    layer2_outputs(4422) <= not(layer1_outputs(2676));
    layer2_outputs(4423) <= (layer1_outputs(10911)) xor (layer1_outputs(3744));
    layer2_outputs(4424) <= (layer1_outputs(1441)) and not (layer1_outputs(5222));
    layer2_outputs(4425) <= not(layer1_outputs(11329));
    layer2_outputs(4426) <= not(layer1_outputs(10640)) or (layer1_outputs(55));
    layer2_outputs(4427) <= layer1_outputs(5213);
    layer2_outputs(4428) <= layer1_outputs(547);
    layer2_outputs(4429) <= not(layer1_outputs(3809));
    layer2_outputs(4430) <= (layer1_outputs(8866)) and (layer1_outputs(4346));
    layer2_outputs(4431) <= not((layer1_outputs(9864)) xor (layer1_outputs(12072)));
    layer2_outputs(4432) <= layer1_outputs(2288);
    layer2_outputs(4433) <= (layer1_outputs(4469)) and not (layer1_outputs(1107));
    layer2_outputs(4434) <= not((layer1_outputs(5533)) xor (layer1_outputs(12153)));
    layer2_outputs(4435) <= (layer1_outputs(10838)) xor (layer1_outputs(690));
    layer2_outputs(4436) <= layer1_outputs(2608);
    layer2_outputs(4437) <= (layer1_outputs(10393)) and not (layer1_outputs(12436));
    layer2_outputs(4438) <= (layer1_outputs(1499)) and (layer1_outputs(3756));
    layer2_outputs(4439) <= layer1_outputs(516);
    layer2_outputs(4440) <= not(layer1_outputs(12266));
    layer2_outputs(4441) <= layer1_outputs(6511);
    layer2_outputs(4442) <= not(layer1_outputs(5818)) or (layer1_outputs(4034));
    layer2_outputs(4443) <= not((layer1_outputs(2905)) xor (layer1_outputs(2580)));
    layer2_outputs(4444) <= not(layer1_outputs(6390));
    layer2_outputs(4445) <= (layer1_outputs(1969)) or (layer1_outputs(6559));
    layer2_outputs(4446) <= layer1_outputs(9361);
    layer2_outputs(4447) <= '0';
    layer2_outputs(4448) <= (layer1_outputs(1589)) xor (layer1_outputs(5131));
    layer2_outputs(4449) <= layer1_outputs(1621);
    layer2_outputs(4450) <= not(layer1_outputs(2908)) or (layer1_outputs(10244));
    layer2_outputs(4451) <= not((layer1_outputs(6979)) and (layer1_outputs(8411)));
    layer2_outputs(4452) <= (layer1_outputs(10024)) xor (layer1_outputs(11628));
    layer2_outputs(4453) <= layer1_outputs(8373);
    layer2_outputs(4454) <= (layer1_outputs(12288)) and not (layer1_outputs(8608));
    layer2_outputs(4455) <= (layer1_outputs(1691)) xor (layer1_outputs(9862));
    layer2_outputs(4456) <= not(layer1_outputs(8263));
    layer2_outputs(4457) <= layer1_outputs(552);
    layer2_outputs(4458) <= layer1_outputs(631);
    layer2_outputs(4459) <= not(layer1_outputs(9340));
    layer2_outputs(4460) <= layer1_outputs(5527);
    layer2_outputs(4461) <= layer1_outputs(3324);
    layer2_outputs(4462) <= not((layer1_outputs(9446)) and (layer1_outputs(3397)));
    layer2_outputs(4463) <= (layer1_outputs(8386)) and not (layer1_outputs(6326));
    layer2_outputs(4464) <= not((layer1_outputs(2831)) xor (layer1_outputs(2947)));
    layer2_outputs(4465) <= not((layer1_outputs(1143)) xor (layer1_outputs(2564)));
    layer2_outputs(4466) <= (layer1_outputs(6576)) xor (layer1_outputs(9444));
    layer2_outputs(4467) <= layer1_outputs(10068);
    layer2_outputs(4468) <= not(layer1_outputs(7949));
    layer2_outputs(4469) <= not(layer1_outputs(5383));
    layer2_outputs(4470) <= not(layer1_outputs(11161));
    layer2_outputs(4471) <= (layer1_outputs(2879)) xor (layer1_outputs(308));
    layer2_outputs(4472) <= layer1_outputs(7931);
    layer2_outputs(4473) <= layer1_outputs(386);
    layer2_outputs(4474) <= (layer1_outputs(12277)) xor (layer1_outputs(8206));
    layer2_outputs(4475) <= (layer1_outputs(2276)) and not (layer1_outputs(2024));
    layer2_outputs(4476) <= layer1_outputs(6602);
    layer2_outputs(4477) <= layer1_outputs(2219);
    layer2_outputs(4478) <= not((layer1_outputs(8902)) xor (layer1_outputs(12709)));
    layer2_outputs(4479) <= layer1_outputs(8712);
    layer2_outputs(4480) <= not(layer1_outputs(5371));
    layer2_outputs(4481) <= not((layer1_outputs(2359)) xor (layer1_outputs(565)));
    layer2_outputs(4482) <= not(layer1_outputs(12640)) or (layer1_outputs(9734));
    layer2_outputs(4483) <= (layer1_outputs(11110)) and not (layer1_outputs(7061));
    layer2_outputs(4484) <= not((layer1_outputs(8996)) xor (layer1_outputs(4522)));
    layer2_outputs(4485) <= not(layer1_outputs(2661)) or (layer1_outputs(1580));
    layer2_outputs(4486) <= not(layer1_outputs(8136));
    layer2_outputs(4487) <= not(layer1_outputs(4032));
    layer2_outputs(4488) <= not((layer1_outputs(9148)) xor (layer1_outputs(10788)));
    layer2_outputs(4489) <= (layer1_outputs(567)) and not (layer1_outputs(3968));
    layer2_outputs(4490) <= not(layer1_outputs(4917));
    layer2_outputs(4491) <= (layer1_outputs(919)) or (layer1_outputs(7565));
    layer2_outputs(4492) <= not((layer1_outputs(4329)) and (layer1_outputs(12004)));
    layer2_outputs(4493) <= (layer1_outputs(3860)) or (layer1_outputs(10255));
    layer2_outputs(4494) <= not((layer1_outputs(4257)) or (layer1_outputs(6)));
    layer2_outputs(4495) <= layer1_outputs(9277);
    layer2_outputs(4496) <= not(layer1_outputs(5382));
    layer2_outputs(4497) <= not(layer1_outputs(9472)) or (layer1_outputs(4743));
    layer2_outputs(4498) <= not((layer1_outputs(6404)) xor (layer1_outputs(12781)));
    layer2_outputs(4499) <= not(layer1_outputs(12060));
    layer2_outputs(4500) <= not((layer1_outputs(197)) or (layer1_outputs(2535)));
    layer2_outputs(4501) <= (layer1_outputs(8026)) or (layer1_outputs(1012));
    layer2_outputs(4502) <= (layer1_outputs(4104)) or (layer1_outputs(10672));
    layer2_outputs(4503) <= (layer1_outputs(7466)) and not (layer1_outputs(2506));
    layer2_outputs(4504) <= not((layer1_outputs(7139)) xor (layer1_outputs(6724)));
    layer2_outputs(4505) <= layer1_outputs(3462);
    layer2_outputs(4506) <= (layer1_outputs(3232)) and (layer1_outputs(6864));
    layer2_outputs(4507) <= (layer1_outputs(502)) xor (layer1_outputs(1777));
    layer2_outputs(4508) <= not(layer1_outputs(6498));
    layer2_outputs(4509) <= not(layer1_outputs(4293));
    layer2_outputs(4510) <= layer1_outputs(4199);
    layer2_outputs(4511) <= layer1_outputs(2088);
    layer2_outputs(4512) <= not(layer1_outputs(10211)) or (layer1_outputs(904));
    layer2_outputs(4513) <= layer1_outputs(5748);
    layer2_outputs(4514) <= layer1_outputs(9210);
    layer2_outputs(4515) <= not(layer1_outputs(10723));
    layer2_outputs(4516) <= not(layer1_outputs(8880));
    layer2_outputs(4517) <= layer1_outputs(3552);
    layer2_outputs(4518) <= not(layer1_outputs(9862)) or (layer1_outputs(2511));
    layer2_outputs(4519) <= not((layer1_outputs(7437)) or (layer1_outputs(8084)));
    layer2_outputs(4520) <= layer1_outputs(7755);
    layer2_outputs(4521) <= (layer1_outputs(1279)) and (layer1_outputs(6189));
    layer2_outputs(4522) <= not((layer1_outputs(4381)) xor (layer1_outputs(1716)));
    layer2_outputs(4523) <= layer1_outputs(8589);
    layer2_outputs(4524) <= (layer1_outputs(7644)) and not (layer1_outputs(2620));
    layer2_outputs(4525) <= layer1_outputs(12487);
    layer2_outputs(4526) <= (layer1_outputs(5590)) xor (layer1_outputs(6646));
    layer2_outputs(4527) <= not(layer1_outputs(11525));
    layer2_outputs(4528) <= not((layer1_outputs(8304)) or (layer1_outputs(1634)));
    layer2_outputs(4529) <= not(layer1_outputs(513));
    layer2_outputs(4530) <= (layer1_outputs(3418)) and (layer1_outputs(8331));
    layer2_outputs(4531) <= (layer1_outputs(12599)) or (layer1_outputs(4302));
    layer2_outputs(4532) <= (layer1_outputs(1186)) or (layer1_outputs(4372));
    layer2_outputs(4533) <= not(layer1_outputs(7079));
    layer2_outputs(4534) <= not(layer1_outputs(2479));
    layer2_outputs(4535) <= not(layer1_outputs(7841));
    layer2_outputs(4536) <= layer1_outputs(1674);
    layer2_outputs(4537) <= layer1_outputs(2606);
    layer2_outputs(4538) <= layer1_outputs(9218);
    layer2_outputs(4539) <= not((layer1_outputs(5730)) xor (layer1_outputs(2142)));
    layer2_outputs(4540) <= (layer1_outputs(3289)) and not (layer1_outputs(3748));
    layer2_outputs(4541) <= not((layer1_outputs(4347)) xor (layer1_outputs(9534)));
    layer2_outputs(4542) <= (layer1_outputs(10685)) xor (layer1_outputs(12344));
    layer2_outputs(4543) <= not((layer1_outputs(4094)) xor (layer1_outputs(3206)));
    layer2_outputs(4544) <= not((layer1_outputs(6499)) xor (layer1_outputs(3071)));
    layer2_outputs(4545) <= not((layer1_outputs(10165)) or (layer1_outputs(3806)));
    layer2_outputs(4546) <= layer1_outputs(4156);
    layer2_outputs(4547) <= not(layer1_outputs(11847));
    layer2_outputs(4548) <= not(layer1_outputs(12074));
    layer2_outputs(4549) <= (layer1_outputs(1436)) xor (layer1_outputs(8134));
    layer2_outputs(4550) <= not(layer1_outputs(3220)) or (layer1_outputs(12435));
    layer2_outputs(4551) <= not(layer1_outputs(2635)) or (layer1_outputs(2631));
    layer2_outputs(4552) <= not(layer1_outputs(11381));
    layer2_outputs(4553) <= layer1_outputs(1622);
    layer2_outputs(4554) <= (layer1_outputs(7214)) and (layer1_outputs(2549));
    layer2_outputs(4555) <= layer1_outputs(10157);
    layer2_outputs(4556) <= not(layer1_outputs(12708));
    layer2_outputs(4557) <= not(layer1_outputs(3427)) or (layer1_outputs(11214));
    layer2_outputs(4558) <= not(layer1_outputs(3384)) or (layer1_outputs(3262));
    layer2_outputs(4559) <= layer1_outputs(316);
    layer2_outputs(4560) <= not(layer1_outputs(2514));
    layer2_outputs(4561) <= (layer1_outputs(9573)) or (layer1_outputs(422));
    layer2_outputs(4562) <= (layer1_outputs(968)) and not (layer1_outputs(1293));
    layer2_outputs(4563) <= (layer1_outputs(1846)) and not (layer1_outputs(1728));
    layer2_outputs(4564) <= layer1_outputs(1939);
    layer2_outputs(4565) <= not(layer1_outputs(2060));
    layer2_outputs(4566) <= not((layer1_outputs(10554)) and (layer1_outputs(750)));
    layer2_outputs(4567) <= layer1_outputs(8293);
    layer2_outputs(4568) <= layer1_outputs(2194);
    layer2_outputs(4569) <= not(layer1_outputs(4183));
    layer2_outputs(4570) <= not((layer1_outputs(8135)) or (layer1_outputs(6764)));
    layer2_outputs(4571) <= (layer1_outputs(11704)) and not (layer1_outputs(5319));
    layer2_outputs(4572) <= not(layer1_outputs(6815));
    layer2_outputs(4573) <= layer1_outputs(5109);
    layer2_outputs(4574) <= not(layer1_outputs(10498));
    layer2_outputs(4575) <= layer1_outputs(4008);
    layer2_outputs(4576) <= not((layer1_outputs(10173)) xor (layer1_outputs(8786)));
    layer2_outputs(4577) <= not(layer1_outputs(7690));
    layer2_outputs(4578) <= not(layer1_outputs(5825)) or (layer1_outputs(5777));
    layer2_outputs(4579) <= (layer1_outputs(3478)) xor (layer1_outputs(4888));
    layer2_outputs(4580) <= layer1_outputs(10392);
    layer2_outputs(4581) <= (layer1_outputs(5750)) xor (layer1_outputs(1479));
    layer2_outputs(4582) <= not(layer1_outputs(6706));
    layer2_outputs(4583) <= not(layer1_outputs(10632));
    layer2_outputs(4584) <= layer1_outputs(7089);
    layer2_outputs(4585) <= layer1_outputs(11615);
    layer2_outputs(4586) <= not(layer1_outputs(5302));
    layer2_outputs(4587) <= not((layer1_outputs(6440)) xor (layer1_outputs(10877)));
    layer2_outputs(4588) <= (layer1_outputs(9668)) and not (layer1_outputs(12304));
    layer2_outputs(4589) <= layer1_outputs(3407);
    layer2_outputs(4590) <= not((layer1_outputs(8837)) xor (layer1_outputs(6470)));
    layer2_outputs(4591) <= not((layer1_outputs(5414)) xor (layer1_outputs(12013)));
    layer2_outputs(4592) <= not(layer1_outputs(10986));
    layer2_outputs(4593) <= not(layer1_outputs(4633));
    layer2_outputs(4594) <= not(layer1_outputs(4266));
    layer2_outputs(4595) <= layer1_outputs(5053);
    layer2_outputs(4596) <= not(layer1_outputs(11266)) or (layer1_outputs(11315));
    layer2_outputs(4597) <= not(layer1_outputs(7943));
    layer2_outputs(4598) <= layer1_outputs(7619);
    layer2_outputs(4599) <= (layer1_outputs(8030)) and (layer1_outputs(11232));
    layer2_outputs(4600) <= not(layer1_outputs(12105));
    layer2_outputs(4601) <= (layer1_outputs(5104)) and not (layer1_outputs(791));
    layer2_outputs(4602) <= not(layer1_outputs(1108));
    layer2_outputs(4603) <= not(layer1_outputs(5521));
    layer2_outputs(4604) <= not(layer1_outputs(2829));
    layer2_outputs(4605) <= (layer1_outputs(3227)) xor (layer1_outputs(11023));
    layer2_outputs(4606) <= layer1_outputs(7926);
    layer2_outputs(4607) <= (layer1_outputs(6758)) and (layer1_outputs(6306));
    layer2_outputs(4608) <= not(layer1_outputs(276));
    layer2_outputs(4609) <= (layer1_outputs(4269)) and not (layer1_outputs(2792));
    layer2_outputs(4610) <= (layer1_outputs(12775)) and not (layer1_outputs(5234));
    layer2_outputs(4611) <= layer1_outputs(10702);
    layer2_outputs(4612) <= not(layer1_outputs(11630));
    layer2_outputs(4613) <= not(layer1_outputs(5172));
    layer2_outputs(4614) <= layer1_outputs(127);
    layer2_outputs(4615) <= (layer1_outputs(8932)) and not (layer1_outputs(4446));
    layer2_outputs(4616) <= (layer1_outputs(10010)) and not (layer1_outputs(335));
    layer2_outputs(4617) <= not(layer1_outputs(1934));
    layer2_outputs(4618) <= (layer1_outputs(5239)) and not (layer1_outputs(8248));
    layer2_outputs(4619) <= layer1_outputs(3075);
    layer2_outputs(4620) <= not((layer1_outputs(6175)) xor (layer1_outputs(7473)));
    layer2_outputs(4621) <= layer1_outputs(7339);
    layer2_outputs(4622) <= not((layer1_outputs(10819)) or (layer1_outputs(8984)));
    layer2_outputs(4623) <= layer1_outputs(7313);
    layer2_outputs(4624) <= layer1_outputs(2907);
    layer2_outputs(4625) <= not(layer1_outputs(409)) or (layer1_outputs(11892));
    layer2_outputs(4626) <= not((layer1_outputs(1689)) xor (layer1_outputs(222)));
    layer2_outputs(4627) <= not((layer1_outputs(8895)) and (layer1_outputs(2084)));
    layer2_outputs(4628) <= layer1_outputs(7166);
    layer2_outputs(4629) <= not(layer1_outputs(5800));
    layer2_outputs(4630) <= not(layer1_outputs(3498));
    layer2_outputs(4631) <= layer1_outputs(9641);
    layer2_outputs(4632) <= not(layer1_outputs(5791));
    layer2_outputs(4633) <= layer1_outputs(9326);
    layer2_outputs(4634) <= layer1_outputs(8821);
    layer2_outputs(4635) <= not(layer1_outputs(3495));
    layer2_outputs(4636) <= (layer1_outputs(2422)) and not (layer1_outputs(4081));
    layer2_outputs(4637) <= layer1_outputs(3124);
    layer2_outputs(4638) <= layer1_outputs(6318);
    layer2_outputs(4639) <= not(layer1_outputs(6911));
    layer2_outputs(4640) <= not((layer1_outputs(10319)) or (layer1_outputs(6552)));
    layer2_outputs(4641) <= not(layer1_outputs(353));
    layer2_outputs(4642) <= (layer1_outputs(10330)) and not (layer1_outputs(3970));
    layer2_outputs(4643) <= not(layer1_outputs(7196));
    layer2_outputs(4644) <= not((layer1_outputs(4127)) and (layer1_outputs(1040)));
    layer2_outputs(4645) <= (layer1_outputs(3292)) or (layer1_outputs(9452));
    layer2_outputs(4646) <= (layer1_outputs(549)) or (layer1_outputs(2293));
    layer2_outputs(4647) <= not(layer1_outputs(264));
    layer2_outputs(4648) <= (layer1_outputs(9334)) or (layer1_outputs(4606));
    layer2_outputs(4649) <= layer1_outputs(9146);
    layer2_outputs(4650) <= not(layer1_outputs(6635));
    layer2_outputs(4651) <= layer1_outputs(11530);
    layer2_outputs(4652) <= (layer1_outputs(12098)) xor (layer1_outputs(12430));
    layer2_outputs(4653) <= (layer1_outputs(659)) and not (layer1_outputs(9204));
    layer2_outputs(4654) <= layer1_outputs(243);
    layer2_outputs(4655) <= not(layer1_outputs(5342)) or (layer1_outputs(889));
    layer2_outputs(4656) <= (layer1_outputs(5028)) or (layer1_outputs(1798));
    layer2_outputs(4657) <= layer1_outputs(9081);
    layer2_outputs(4658) <= (layer1_outputs(5956)) xor (layer1_outputs(3651));
    layer2_outputs(4659) <= not(layer1_outputs(11690)) or (layer1_outputs(9773));
    layer2_outputs(4660) <= not(layer1_outputs(8703));
    layer2_outputs(4661) <= not(layer1_outputs(4982));
    layer2_outputs(4662) <= layer1_outputs(9564);
    layer2_outputs(4663) <= not((layer1_outputs(2353)) or (layer1_outputs(5179)));
    layer2_outputs(4664) <= layer1_outputs(131);
    layer2_outputs(4665) <= not(layer1_outputs(10704)) or (layer1_outputs(26));
    layer2_outputs(4666) <= not(layer1_outputs(2650));
    layer2_outputs(4667) <= layer1_outputs(357);
    layer2_outputs(4668) <= not(layer1_outputs(4709));
    layer2_outputs(4669) <= not(layer1_outputs(2526));
    layer2_outputs(4670) <= (layer1_outputs(9289)) and not (layer1_outputs(10825));
    layer2_outputs(4671) <= (layer1_outputs(12484)) and not (layer1_outputs(12029));
    layer2_outputs(4672) <= layer1_outputs(7893);
    layer2_outputs(4673) <= not(layer1_outputs(9827));
    layer2_outputs(4674) <= '0';
    layer2_outputs(4675) <= layer1_outputs(6506);
    layer2_outputs(4676) <= (layer1_outputs(11603)) or (layer1_outputs(4141));
    layer2_outputs(4677) <= (layer1_outputs(7888)) and not (layer1_outputs(4130));
    layer2_outputs(4678) <= not(layer1_outputs(8776));
    layer2_outputs(4679) <= (layer1_outputs(9025)) xor (layer1_outputs(1746));
    layer2_outputs(4680) <= not(layer1_outputs(12182));
    layer2_outputs(4681) <= not((layer1_outputs(10985)) or (layer1_outputs(9600)));
    layer2_outputs(4682) <= (layer1_outputs(4218)) and not (layer1_outputs(9765));
    layer2_outputs(4683) <= not((layer1_outputs(3180)) xor (layer1_outputs(12015)));
    layer2_outputs(4684) <= not(layer1_outputs(5134));
    layer2_outputs(4685) <= layer1_outputs(12794);
    layer2_outputs(4686) <= layer1_outputs(854);
    layer2_outputs(4687) <= (layer1_outputs(12490)) and (layer1_outputs(1147));
    layer2_outputs(4688) <= (layer1_outputs(7076)) xor (layer1_outputs(3400));
    layer2_outputs(4689) <= (layer1_outputs(10448)) and (layer1_outputs(10827));
    layer2_outputs(4690) <= layer1_outputs(4374);
    layer2_outputs(4691) <= not(layer1_outputs(7766));
    layer2_outputs(4692) <= not(layer1_outputs(602));
    layer2_outputs(4693) <= (layer1_outputs(1812)) and not (layer1_outputs(1131));
    layer2_outputs(4694) <= layer1_outputs(7432);
    layer2_outputs(4695) <= not(layer1_outputs(2286));
    layer2_outputs(4696) <= not((layer1_outputs(2812)) or (layer1_outputs(8325)));
    layer2_outputs(4697) <= not(layer1_outputs(3740));
    layer2_outputs(4698) <= not(layer1_outputs(9317));
    layer2_outputs(4699) <= not(layer1_outputs(12243));
    layer2_outputs(4700) <= (layer1_outputs(4122)) and (layer1_outputs(10565));
    layer2_outputs(4701) <= not(layer1_outputs(11072));
    layer2_outputs(4702) <= not(layer1_outputs(6987));
    layer2_outputs(4703) <= not(layer1_outputs(10793));
    layer2_outputs(4704) <= not((layer1_outputs(9132)) or (layer1_outputs(4074)));
    layer2_outputs(4705) <= layer1_outputs(4745);
    layer2_outputs(4706) <= not(layer1_outputs(10017));
    layer2_outputs(4707) <= layer1_outputs(7589);
    layer2_outputs(4708) <= not((layer1_outputs(2417)) and (layer1_outputs(1678)));
    layer2_outputs(4709) <= not((layer1_outputs(2582)) xor (layer1_outputs(9664)));
    layer2_outputs(4710) <= layer1_outputs(2132);
    layer2_outputs(4711) <= (layer1_outputs(594)) and (layer1_outputs(291));
    layer2_outputs(4712) <= (layer1_outputs(7152)) xor (layer1_outputs(6640));
    layer2_outputs(4713) <= '1';
    layer2_outputs(4714) <= not((layer1_outputs(3633)) xor (layer1_outputs(3060)));
    layer2_outputs(4715) <= not((layer1_outputs(4815)) xor (layer1_outputs(9050)));
    layer2_outputs(4716) <= not(layer1_outputs(4739));
    layer2_outputs(4717) <= not(layer1_outputs(1543));
    layer2_outputs(4718) <= (layer1_outputs(12273)) and not (layer1_outputs(7194));
    layer2_outputs(4719) <= not(layer1_outputs(2427));
    layer2_outputs(4720) <= not(layer1_outputs(12235));
    layer2_outputs(4721) <= (layer1_outputs(8778)) and not (layer1_outputs(2300));
    layer2_outputs(4722) <= not(layer1_outputs(10104)) or (layer1_outputs(10372));
    layer2_outputs(4723) <= layer1_outputs(8913);
    layer2_outputs(4724) <= not(layer1_outputs(7683)) or (layer1_outputs(8959));
    layer2_outputs(4725) <= not((layer1_outputs(3945)) xor (layer1_outputs(11656)));
    layer2_outputs(4726) <= (layer1_outputs(12148)) and not (layer1_outputs(3962));
    layer2_outputs(4727) <= not(layer1_outputs(7841)) or (layer1_outputs(7444));
    layer2_outputs(4728) <= not(layer1_outputs(6645));
    layer2_outputs(4729) <= not(layer1_outputs(10650));
    layer2_outputs(4730) <= (layer1_outputs(9101)) xor (layer1_outputs(3509));
    layer2_outputs(4731) <= layer1_outputs(5210);
    layer2_outputs(4732) <= (layer1_outputs(12516)) and not (layer1_outputs(7860));
    layer2_outputs(4733) <= (layer1_outputs(1338)) and (layer1_outputs(10086));
    layer2_outputs(4734) <= not((layer1_outputs(3319)) xor (layer1_outputs(11991)));
    layer2_outputs(4735) <= not((layer1_outputs(6684)) or (layer1_outputs(593)));
    layer2_outputs(4736) <= not((layer1_outputs(9721)) xor (layer1_outputs(11386)));
    layer2_outputs(4737) <= not((layer1_outputs(10905)) xor (layer1_outputs(3231)));
    layer2_outputs(4738) <= not(layer1_outputs(9987));
    layer2_outputs(4739) <= not(layer1_outputs(11246)) or (layer1_outputs(11928));
    layer2_outputs(4740) <= layer1_outputs(4730);
    layer2_outputs(4741) <= (layer1_outputs(4666)) and not (layer1_outputs(3245));
    layer2_outputs(4742) <= not(layer1_outputs(12111));
    layer2_outputs(4743) <= layer1_outputs(8502);
    layer2_outputs(4744) <= not(layer1_outputs(8100)) or (layer1_outputs(8165));
    layer2_outputs(4745) <= layer1_outputs(3842);
    layer2_outputs(4746) <= (layer1_outputs(8142)) xor (layer1_outputs(1461));
    layer2_outputs(4747) <= layer1_outputs(4299);
    layer2_outputs(4748) <= not(layer1_outputs(7931));
    layer2_outputs(4749) <= (layer1_outputs(5806)) or (layer1_outputs(11028));
    layer2_outputs(4750) <= (layer1_outputs(12559)) or (layer1_outputs(4143));
    layer2_outputs(4751) <= (layer1_outputs(5011)) and (layer1_outputs(5697));
    layer2_outputs(4752) <= not(layer1_outputs(5789));
    layer2_outputs(4753) <= not(layer1_outputs(589));
    layer2_outputs(4754) <= not(layer1_outputs(9892));
    layer2_outputs(4755) <= (layer1_outputs(2782)) and not (layer1_outputs(9825));
    layer2_outputs(4756) <= layer1_outputs(9752);
    layer2_outputs(4757) <= not(layer1_outputs(8553)) or (layer1_outputs(12037));
    layer2_outputs(4758) <= layer1_outputs(5710);
    layer2_outputs(4759) <= not((layer1_outputs(329)) xor (layer1_outputs(8068)));
    layer2_outputs(4760) <= layer1_outputs(953);
    layer2_outputs(4761) <= not(layer1_outputs(1967)) or (layer1_outputs(10939));
    layer2_outputs(4762) <= layer1_outputs(7829);
    layer2_outputs(4763) <= not((layer1_outputs(11206)) or (layer1_outputs(8210)));
    layer2_outputs(4764) <= layer1_outputs(2684);
    layer2_outputs(4765) <= layer1_outputs(1294);
    layer2_outputs(4766) <= layer1_outputs(8086);
    layer2_outputs(4767) <= (layer1_outputs(6641)) or (layer1_outputs(1894));
    layer2_outputs(4768) <= not(layer1_outputs(8837));
    layer2_outputs(4769) <= (layer1_outputs(312)) and (layer1_outputs(4520));
    layer2_outputs(4770) <= layer1_outputs(10238);
    layer2_outputs(4771) <= not(layer1_outputs(11558));
    layer2_outputs(4772) <= not(layer1_outputs(5688));
    layer2_outputs(4773) <= (layer1_outputs(3268)) xor (layer1_outputs(6115));
    layer2_outputs(4774) <= (layer1_outputs(3748)) or (layer1_outputs(6626));
    layer2_outputs(4775) <= layer1_outputs(3103);
    layer2_outputs(4776) <= not((layer1_outputs(11210)) xor (layer1_outputs(7542)));
    layer2_outputs(4777) <= layer1_outputs(6021);
    layer2_outputs(4778) <= not(layer1_outputs(2602));
    layer2_outputs(4779) <= not(layer1_outputs(3449)) or (layer1_outputs(1083));
    layer2_outputs(4780) <= not(layer1_outputs(8817));
    layer2_outputs(4781) <= not(layer1_outputs(10377));
    layer2_outputs(4782) <= not(layer1_outputs(10423));
    layer2_outputs(4783) <= (layer1_outputs(12740)) and not (layer1_outputs(2949));
    layer2_outputs(4784) <= not(layer1_outputs(3893));
    layer2_outputs(4785) <= not(layer1_outputs(8119));
    layer2_outputs(4786) <= not(layer1_outputs(1865));
    layer2_outputs(4787) <= (layer1_outputs(6261)) and (layer1_outputs(6612));
    layer2_outputs(4788) <= layer1_outputs(10466);
    layer2_outputs(4789) <= layer1_outputs(6100);
    layer2_outputs(4790) <= layer1_outputs(11126);
    layer2_outputs(4791) <= not(layer1_outputs(1359));
    layer2_outputs(4792) <= not((layer1_outputs(3834)) xor (layer1_outputs(12135)));
    layer2_outputs(4793) <= (layer1_outputs(648)) and (layer1_outputs(5368));
    layer2_outputs(4794) <= layer1_outputs(4490);
    layer2_outputs(4795) <= (layer1_outputs(2590)) xor (layer1_outputs(9289));
    layer2_outputs(4796) <= not((layer1_outputs(175)) xor (layer1_outputs(3030)));
    layer2_outputs(4797) <= not((layer1_outputs(9965)) or (layer1_outputs(163)));
    layer2_outputs(4798) <= layer1_outputs(8699);
    layer2_outputs(4799) <= not(layer1_outputs(11549));
    layer2_outputs(4800) <= (layer1_outputs(6090)) and not (layer1_outputs(7054));
    layer2_outputs(4801) <= not((layer1_outputs(3135)) xor (layer1_outputs(11748)));
    layer2_outputs(4802) <= not(layer1_outputs(9437));
    layer2_outputs(4803) <= not(layer1_outputs(10265));
    layer2_outputs(4804) <= not((layer1_outputs(6476)) or (layer1_outputs(11072)));
    layer2_outputs(4805) <= not(layer1_outputs(657));
    layer2_outputs(4806) <= not(layer1_outputs(1578));
    layer2_outputs(4807) <= not(layer1_outputs(10268));
    layer2_outputs(4808) <= layer1_outputs(168);
    layer2_outputs(4809) <= layer1_outputs(6832);
    layer2_outputs(4810) <= not((layer1_outputs(7417)) and (layer1_outputs(11629)));
    layer2_outputs(4811) <= (layer1_outputs(12614)) and not (layer1_outputs(5084));
    layer2_outputs(4812) <= (layer1_outputs(7602)) or (layer1_outputs(10842));
    layer2_outputs(4813) <= not((layer1_outputs(7940)) xor (layer1_outputs(1273)));
    layer2_outputs(4814) <= (layer1_outputs(6406)) and (layer1_outputs(2530));
    layer2_outputs(4815) <= (layer1_outputs(8828)) and not (layer1_outputs(3601));
    layer2_outputs(4816) <= layer1_outputs(7242);
    layer2_outputs(4817) <= layer1_outputs(7684);
    layer2_outputs(4818) <= (layer1_outputs(9192)) xor (layer1_outputs(5078));
    layer2_outputs(4819) <= not((layer1_outputs(6834)) xor (layer1_outputs(9513)));
    layer2_outputs(4820) <= not(layer1_outputs(6357));
    layer2_outputs(4821) <= layer1_outputs(12058);
    layer2_outputs(4822) <= not(layer1_outputs(7694));
    layer2_outputs(4823) <= (layer1_outputs(7867)) xor (layer1_outputs(8907));
    layer2_outputs(4824) <= not((layer1_outputs(4387)) xor (layer1_outputs(8518)));
    layer2_outputs(4825) <= layer1_outputs(6965);
    layer2_outputs(4826) <= not(layer1_outputs(1688));
    layer2_outputs(4827) <= not(layer1_outputs(10951)) or (layer1_outputs(1113));
    layer2_outputs(4828) <= layer1_outputs(3814);
    layer2_outputs(4829) <= not(layer1_outputs(9872)) or (layer1_outputs(11546));
    layer2_outputs(4830) <= not((layer1_outputs(1310)) xor (layer1_outputs(9302)));
    layer2_outputs(4831) <= (layer1_outputs(2569)) and not (layer1_outputs(5471));
    layer2_outputs(4832) <= not(layer1_outputs(7692));
    layer2_outputs(4833) <= layer1_outputs(10684);
    layer2_outputs(4834) <= not(layer1_outputs(4938));
    layer2_outputs(4835) <= (layer1_outputs(3979)) xor (layer1_outputs(8448));
    layer2_outputs(4836) <= (layer1_outputs(1756)) or (layer1_outputs(1530));
    layer2_outputs(4837) <= layer1_outputs(4342);
    layer2_outputs(4838) <= layer1_outputs(12103);
    layer2_outputs(4839) <= (layer1_outputs(8510)) xor (layer1_outputs(1303));
    layer2_outputs(4840) <= not((layer1_outputs(343)) xor (layer1_outputs(1454)));
    layer2_outputs(4841) <= layer1_outputs(12520);
    layer2_outputs(4842) <= not(layer1_outputs(12270));
    layer2_outputs(4843) <= (layer1_outputs(7022)) or (layer1_outputs(12707));
    layer2_outputs(4844) <= (layer1_outputs(8469)) xor (layer1_outputs(2246));
    layer2_outputs(4845) <= not((layer1_outputs(12105)) xor (layer1_outputs(441)));
    layer2_outputs(4846) <= not(layer1_outputs(561));
    layer2_outputs(4847) <= (layer1_outputs(5136)) and (layer1_outputs(9270));
    layer2_outputs(4848) <= not((layer1_outputs(6145)) xor (layer1_outputs(2190)));
    layer2_outputs(4849) <= not(layer1_outputs(10008)) or (layer1_outputs(12332));
    layer2_outputs(4850) <= not((layer1_outputs(8197)) and (layer1_outputs(1392)));
    layer2_outputs(4851) <= not(layer1_outputs(8463));
    layer2_outputs(4852) <= not(layer1_outputs(9684));
    layer2_outputs(4853) <= (layer1_outputs(3521)) and not (layer1_outputs(7040));
    layer2_outputs(4854) <= layer1_outputs(7485);
    layer2_outputs(4855) <= not((layer1_outputs(3132)) and (layer1_outputs(4155)));
    layer2_outputs(4856) <= layer1_outputs(1014);
    layer2_outputs(4857) <= (layer1_outputs(3503)) and not (layer1_outputs(10613));
    layer2_outputs(4858) <= layer1_outputs(2844);
    layer2_outputs(4859) <= not(layer1_outputs(7729));
    layer2_outputs(4860) <= not((layer1_outputs(1463)) or (layer1_outputs(5612)));
    layer2_outputs(4861) <= not(layer1_outputs(4211));
    layer2_outputs(4862) <= (layer1_outputs(10359)) and not (layer1_outputs(7236));
    layer2_outputs(4863) <= (layer1_outputs(9145)) xor (layer1_outputs(11990));
    layer2_outputs(4864) <= not((layer1_outputs(6254)) xor (layer1_outputs(5378)));
    layer2_outputs(4865) <= layer1_outputs(827);
    layer2_outputs(4866) <= (layer1_outputs(12432)) xor (layer1_outputs(318));
    layer2_outputs(4867) <= (layer1_outputs(3597)) and (layer1_outputs(10349));
    layer2_outputs(4868) <= layer1_outputs(3737);
    layer2_outputs(4869) <= not(layer1_outputs(542));
    layer2_outputs(4870) <= layer1_outputs(12260);
    layer2_outputs(4871) <= (layer1_outputs(8434)) and (layer1_outputs(6715));
    layer2_outputs(4872) <= (layer1_outputs(7403)) and not (layer1_outputs(7278));
    layer2_outputs(4873) <= not(layer1_outputs(10920));
    layer2_outputs(4874) <= not(layer1_outputs(9033)) or (layer1_outputs(5903));
    layer2_outputs(4875) <= (layer1_outputs(588)) xor (layer1_outputs(10707));
    layer2_outputs(4876) <= not(layer1_outputs(10134)) or (layer1_outputs(3608));
    layer2_outputs(4877) <= layer1_outputs(2241);
    layer2_outputs(4878) <= layer1_outputs(8463);
    layer2_outputs(4879) <= layer1_outputs(11410);
    layer2_outputs(4880) <= not((layer1_outputs(6366)) xor (layer1_outputs(2646)));
    layer2_outputs(4881) <= layer1_outputs(12766);
    layer2_outputs(4882) <= not(layer1_outputs(9375));
    layer2_outputs(4883) <= not((layer1_outputs(5813)) or (layer1_outputs(946)));
    layer2_outputs(4884) <= not(layer1_outputs(8103));
    layer2_outputs(4885) <= layer1_outputs(9900);
    layer2_outputs(4886) <= not(layer1_outputs(581));
    layer2_outputs(4887) <= (layer1_outputs(4664)) and not (layer1_outputs(7811));
    layer2_outputs(4888) <= not(layer1_outputs(3364));
    layer2_outputs(4889) <= not(layer1_outputs(9982));
    layer2_outputs(4890) <= (layer1_outputs(5079)) and not (layer1_outputs(914));
    layer2_outputs(4891) <= layer1_outputs(2165);
    layer2_outputs(4892) <= (layer1_outputs(3941)) and (layer1_outputs(12419));
    layer2_outputs(4893) <= (layer1_outputs(6396)) and not (layer1_outputs(10754));
    layer2_outputs(4894) <= (layer1_outputs(1396)) xor (layer1_outputs(8094));
    layer2_outputs(4895) <= not((layer1_outputs(3180)) and (layer1_outputs(9591)));
    layer2_outputs(4896) <= layer1_outputs(3528);
    layer2_outputs(4897) <= not((layer1_outputs(8429)) and (layer1_outputs(10465)));
    layer2_outputs(4898) <= (layer1_outputs(6777)) xor (layer1_outputs(11049));
    layer2_outputs(4899) <= not(layer1_outputs(6053)) or (layer1_outputs(5363));
    layer2_outputs(4900) <= layer1_outputs(8857);
    layer2_outputs(4901) <= layer1_outputs(9443);
    layer2_outputs(4902) <= (layer1_outputs(7723)) and not (layer1_outputs(12620));
    layer2_outputs(4903) <= not(layer1_outputs(7659));
    layer2_outputs(4904) <= (layer1_outputs(5071)) or (layer1_outputs(1839));
    layer2_outputs(4905) <= (layer1_outputs(7094)) and not (layer1_outputs(11505));
    layer2_outputs(4906) <= layer1_outputs(9704);
    layer2_outputs(4907) <= layer1_outputs(10315);
    layer2_outputs(4908) <= (layer1_outputs(9809)) xor (layer1_outputs(1686));
    layer2_outputs(4909) <= (layer1_outputs(2331)) or (layer1_outputs(8057));
    layer2_outputs(4910) <= (layer1_outputs(3928)) and (layer1_outputs(3039));
    layer2_outputs(4911) <= layer1_outputs(1621);
    layer2_outputs(4912) <= (layer1_outputs(9937)) xor (layer1_outputs(2493));
    layer2_outputs(4913) <= not(layer1_outputs(3483));
    layer2_outputs(4914) <= layer1_outputs(3831);
    layer2_outputs(4915) <= not((layer1_outputs(4404)) xor (layer1_outputs(8410)));
    layer2_outputs(4916) <= layer1_outputs(11750);
    layer2_outputs(4917) <= not(layer1_outputs(11642));
    layer2_outputs(4918) <= layer1_outputs(9074);
    layer2_outputs(4919) <= not(layer1_outputs(12102));
    layer2_outputs(4920) <= (layer1_outputs(11167)) and (layer1_outputs(5528));
    layer2_outputs(4921) <= not((layer1_outputs(11556)) or (layer1_outputs(2780)));
    layer2_outputs(4922) <= not((layer1_outputs(5385)) xor (layer1_outputs(1683)));
    layer2_outputs(4923) <= not(layer1_outputs(3647));
    layer2_outputs(4924) <= not(layer1_outputs(4057));
    layer2_outputs(4925) <= layer1_outputs(2355);
    layer2_outputs(4926) <= not(layer1_outputs(4097));
    layer2_outputs(4927) <= not((layer1_outputs(5636)) or (layer1_outputs(6486)));
    layer2_outputs(4928) <= not(layer1_outputs(1690));
    layer2_outputs(4929) <= not(layer1_outputs(11948));
    layer2_outputs(4930) <= not((layer1_outputs(1715)) xor (layer1_outputs(6373)));
    layer2_outputs(4931) <= not(layer1_outputs(7445));
    layer2_outputs(4932) <= (layer1_outputs(2089)) and not (layer1_outputs(6790));
    layer2_outputs(4933) <= not(layer1_outputs(4956)) or (layer1_outputs(7648));
    layer2_outputs(4934) <= not((layer1_outputs(3564)) xor (layer1_outputs(5406)));
    layer2_outputs(4935) <= layer1_outputs(9398);
    layer2_outputs(4936) <= (layer1_outputs(1611)) and not (layer1_outputs(894));
    layer2_outputs(4937) <= not(layer1_outputs(5689));
    layer2_outputs(4938) <= layer1_outputs(7885);
    layer2_outputs(4939) <= layer1_outputs(9072);
    layer2_outputs(4940) <= not(layer1_outputs(10595));
    layer2_outputs(4941) <= not((layer1_outputs(5477)) xor (layer1_outputs(1734)));
    layer2_outputs(4942) <= (layer1_outputs(6871)) xor (layer1_outputs(9820));
    layer2_outputs(4943) <= layer1_outputs(7235);
    layer2_outputs(4944) <= (layer1_outputs(9750)) xor (layer1_outputs(3049));
    layer2_outputs(4945) <= layer1_outputs(36);
    layer2_outputs(4946) <= layer1_outputs(11462);
    layer2_outputs(4947) <= (layer1_outputs(774)) or (layer1_outputs(5257));
    layer2_outputs(4948) <= not(layer1_outputs(11882));
    layer2_outputs(4949) <= (layer1_outputs(4843)) or (layer1_outputs(10467));
    layer2_outputs(4950) <= not(layer1_outputs(6273));
    layer2_outputs(4951) <= not(layer1_outputs(6846));
    layer2_outputs(4952) <= layer1_outputs(5359);
    layer2_outputs(4953) <= (layer1_outputs(5242)) xor (layer1_outputs(2009));
    layer2_outputs(4954) <= (layer1_outputs(5270)) xor (layer1_outputs(10833));
    layer2_outputs(4955) <= (layer1_outputs(5346)) and not (layer1_outputs(2529));
    layer2_outputs(4956) <= layer1_outputs(2633);
    layer2_outputs(4957) <= not((layer1_outputs(2641)) or (layer1_outputs(10878)));
    layer2_outputs(4958) <= (layer1_outputs(7631)) and (layer1_outputs(7537));
    layer2_outputs(4959) <= layer1_outputs(1258);
    layer2_outputs(4960) <= (layer1_outputs(1720)) and not (layer1_outputs(6071));
    layer2_outputs(4961) <= not((layer1_outputs(11474)) or (layer1_outputs(2002)));
    layer2_outputs(4962) <= layer1_outputs(11921);
    layer2_outputs(4963) <= not(layer1_outputs(2139));
    layer2_outputs(4964) <= (layer1_outputs(10092)) and not (layer1_outputs(12644));
    layer2_outputs(4965) <= (layer1_outputs(2311)) and (layer1_outputs(3110));
    layer2_outputs(4966) <= not(layer1_outputs(12565));
    layer2_outputs(4967) <= not((layer1_outputs(5556)) or (layer1_outputs(4500)));
    layer2_outputs(4968) <= not(layer1_outputs(8574)) or (layer1_outputs(11412));
    layer2_outputs(4969) <= (layer1_outputs(5820)) or (layer1_outputs(7165));
    layer2_outputs(4970) <= layer1_outputs(10575);
    layer2_outputs(4971) <= layer1_outputs(12513);
    layer2_outputs(4972) <= not(layer1_outputs(7948)) or (layer1_outputs(5327));
    layer2_outputs(4973) <= not((layer1_outputs(11576)) xor (layer1_outputs(9622)));
    layer2_outputs(4974) <= not(layer1_outputs(6034));
    layer2_outputs(4975) <= layer1_outputs(6801);
    layer2_outputs(4976) <= not(layer1_outputs(12324));
    layer2_outputs(4977) <= (layer1_outputs(3791)) and not (layer1_outputs(7760));
    layer2_outputs(4978) <= not(layer1_outputs(12797));
    layer2_outputs(4979) <= not(layer1_outputs(6931));
    layer2_outputs(4980) <= not(layer1_outputs(2701));
    layer2_outputs(4981) <= layer1_outputs(3219);
    layer2_outputs(4982) <= (layer1_outputs(3359)) and not (layer1_outputs(1233));
    layer2_outputs(4983) <= (layer1_outputs(5644)) and (layer1_outputs(11345));
    layer2_outputs(4984) <= not(layer1_outputs(1501)) or (layer1_outputs(3486));
    layer2_outputs(4985) <= not(layer1_outputs(11942));
    layer2_outputs(4986) <= not((layer1_outputs(12208)) and (layer1_outputs(5250)));
    layer2_outputs(4987) <= layer1_outputs(4478);
    layer2_outputs(4988) <= not(layer1_outputs(9787));
    layer2_outputs(4989) <= not(layer1_outputs(11468));
    layer2_outputs(4990) <= layer1_outputs(12096);
    layer2_outputs(4991) <= (layer1_outputs(12530)) or (layer1_outputs(11651));
    layer2_outputs(4992) <= (layer1_outputs(6783)) or (layer1_outputs(2630));
    layer2_outputs(4993) <= not(layer1_outputs(12639)) or (layer1_outputs(7539));
    layer2_outputs(4994) <= not(layer1_outputs(2399)) or (layer1_outputs(10101));
    layer2_outputs(4995) <= (layer1_outputs(636)) or (layer1_outputs(11160));
    layer2_outputs(4996) <= (layer1_outputs(3835)) and not (layer1_outputs(7122));
    layer2_outputs(4997) <= layer1_outputs(5050);
    layer2_outputs(4998) <= not((layer1_outputs(5129)) and (layer1_outputs(7122)));
    layer2_outputs(4999) <= layer1_outputs(5863);
    layer2_outputs(5000) <= layer1_outputs(1015);
    layer2_outputs(5001) <= (layer1_outputs(7373)) and not (layer1_outputs(8131));
    layer2_outputs(5002) <= not(layer1_outputs(2007));
    layer2_outputs(5003) <= not(layer1_outputs(7410));
    layer2_outputs(5004) <= not((layer1_outputs(6050)) and (layer1_outputs(12051)));
    layer2_outputs(5005) <= not(layer1_outputs(3369)) or (layer1_outputs(6508));
    layer2_outputs(5006) <= not((layer1_outputs(11480)) and (layer1_outputs(2522)));
    layer2_outputs(5007) <= layer1_outputs(5180);
    layer2_outputs(5008) <= layer1_outputs(12038);
    layer2_outputs(5009) <= not(layer1_outputs(9102));
    layer2_outputs(5010) <= layer1_outputs(7123);
    layer2_outputs(5011) <= not(layer1_outputs(12181));
    layer2_outputs(5012) <= (layer1_outputs(8004)) xor (layer1_outputs(912));
    layer2_outputs(5013) <= not(layer1_outputs(2694));
    layer2_outputs(5014) <= not(layer1_outputs(10808));
    layer2_outputs(5015) <= (layer1_outputs(11780)) and not (layer1_outputs(12723));
    layer2_outputs(5016) <= (layer1_outputs(2585)) and not (layer1_outputs(7225));
    layer2_outputs(5017) <= (layer1_outputs(11188)) and not (layer1_outputs(4495));
    layer2_outputs(5018) <= not(layer1_outputs(7119));
    layer2_outputs(5019) <= not((layer1_outputs(406)) and (layer1_outputs(8578)));
    layer2_outputs(5020) <= not(layer1_outputs(11372)) or (layer1_outputs(10473));
    layer2_outputs(5021) <= layer1_outputs(3706);
    layer2_outputs(5022) <= (layer1_outputs(12001)) and (layer1_outputs(2011));
    layer2_outputs(5023) <= layer1_outputs(11345);
    layer2_outputs(5024) <= (layer1_outputs(11617)) xor (layer1_outputs(4714));
    layer2_outputs(5025) <= not((layer1_outputs(12080)) xor (layer1_outputs(4188)));
    layer2_outputs(5026) <= (layer1_outputs(9541)) xor (layer1_outputs(7047));
    layer2_outputs(5027) <= not((layer1_outputs(10950)) or (layer1_outputs(7704)));
    layer2_outputs(5028) <= not((layer1_outputs(10605)) or (layer1_outputs(8187)));
    layer2_outputs(5029) <= not(layer1_outputs(7359));
    layer2_outputs(5030) <= layer1_outputs(11312);
    layer2_outputs(5031) <= not((layer1_outputs(8595)) or (layer1_outputs(12287)));
    layer2_outputs(5032) <= not((layer1_outputs(3954)) and (layer1_outputs(10275)));
    layer2_outputs(5033) <= layer1_outputs(7091);
    layer2_outputs(5034) <= (layer1_outputs(7411)) xor (layer1_outputs(500));
    layer2_outputs(5035) <= layer1_outputs(4197);
    layer2_outputs(5036) <= (layer1_outputs(9164)) xor (layer1_outputs(182));
    layer2_outputs(5037) <= not(layer1_outputs(2541));
    layer2_outputs(5038) <= not(layer1_outputs(3477));
    layer2_outputs(5039) <= layer1_outputs(8040);
    layer2_outputs(5040) <= (layer1_outputs(8964)) xor (layer1_outputs(11271));
    layer2_outputs(5041) <= layer1_outputs(12533);
    layer2_outputs(5042) <= not((layer1_outputs(9327)) or (layer1_outputs(704)));
    layer2_outputs(5043) <= not(layer1_outputs(4146));
    layer2_outputs(5044) <= layer1_outputs(10487);
    layer2_outputs(5045) <= not((layer1_outputs(403)) xor (layer1_outputs(3958)));
    layer2_outputs(5046) <= not(layer1_outputs(3392)) or (layer1_outputs(7945));
    layer2_outputs(5047) <= not(layer1_outputs(4602));
    layer2_outputs(5048) <= layer1_outputs(8313);
    layer2_outputs(5049) <= (layer1_outputs(6697)) and (layer1_outputs(12749));
    layer2_outputs(5050) <= (layer1_outputs(456)) and not (layer1_outputs(2582));
    layer2_outputs(5051) <= not(layer1_outputs(2660));
    layer2_outputs(5052) <= not(layer1_outputs(4656));
    layer2_outputs(5053) <= layer1_outputs(1599);
    layer2_outputs(5054) <= layer1_outputs(12034);
    layer2_outputs(5055) <= (layer1_outputs(379)) and not (layer1_outputs(3015));
    layer2_outputs(5056) <= layer1_outputs(10140);
    layer2_outputs(5057) <= not(layer1_outputs(9305));
    layer2_outputs(5058) <= not(layer1_outputs(12419));
    layer2_outputs(5059) <= not(layer1_outputs(12445));
    layer2_outputs(5060) <= not(layer1_outputs(6583));
    layer2_outputs(5061) <= not(layer1_outputs(10562));
    layer2_outputs(5062) <= (layer1_outputs(1604)) and not (layer1_outputs(10524));
    layer2_outputs(5063) <= (layer1_outputs(9692)) and (layer1_outputs(6079));
    layer2_outputs(5064) <= not((layer1_outputs(11938)) or (layer1_outputs(798)));
    layer2_outputs(5065) <= (layer1_outputs(4334)) and not (layer1_outputs(12038));
    layer2_outputs(5066) <= not(layer1_outputs(10675));
    layer2_outputs(5067) <= layer1_outputs(1440);
    layer2_outputs(5068) <= not((layer1_outputs(3465)) or (layer1_outputs(10656)));
    layer2_outputs(5069) <= layer1_outputs(7932);
    layer2_outputs(5070) <= not((layer1_outputs(9489)) or (layer1_outputs(4269)));
    layer2_outputs(5071) <= (layer1_outputs(3898)) and (layer1_outputs(4789));
    layer2_outputs(5072) <= layer1_outputs(6158);
    layer2_outputs(5073) <= (layer1_outputs(9716)) and not (layer1_outputs(11411));
    layer2_outputs(5074) <= '0';
    layer2_outputs(5075) <= (layer1_outputs(2272)) or (layer1_outputs(6806));
    layer2_outputs(5076) <= not(layer1_outputs(3228));
    layer2_outputs(5077) <= not(layer1_outputs(2451));
    layer2_outputs(5078) <= not((layer1_outputs(6524)) and (layer1_outputs(6788)));
    layer2_outputs(5079) <= not(layer1_outputs(10862)) or (layer1_outputs(5255));
    layer2_outputs(5080) <= (layer1_outputs(4367)) xor (layer1_outputs(10245));
    layer2_outputs(5081) <= layer1_outputs(3735);
    layer2_outputs(5082) <= layer1_outputs(3984);
    layer2_outputs(5083) <= not(layer1_outputs(4825));
    layer2_outputs(5084) <= (layer1_outputs(10052)) xor (layer1_outputs(8281));
    layer2_outputs(5085) <= not(layer1_outputs(1552));
    layer2_outputs(5086) <= (layer1_outputs(4499)) and not (layer1_outputs(9198));
    layer2_outputs(5087) <= not(layer1_outputs(7503));
    layer2_outputs(5088) <= not(layer1_outputs(3247)) or (layer1_outputs(6518));
    layer2_outputs(5089) <= layer1_outputs(2133);
    layer2_outputs(5090) <= not(layer1_outputs(1922)) or (layer1_outputs(4403));
    layer2_outputs(5091) <= layer1_outputs(2354);
    layer2_outputs(5092) <= not((layer1_outputs(8113)) xor (layer1_outputs(12241)));
    layer2_outputs(5093) <= (layer1_outputs(6532)) or (layer1_outputs(9895));
    layer2_outputs(5094) <= layer1_outputs(4434);
    layer2_outputs(5095) <= layer1_outputs(9285);
    layer2_outputs(5096) <= (layer1_outputs(9011)) xor (layer1_outputs(10592));
    layer2_outputs(5097) <= (layer1_outputs(6380)) and not (layer1_outputs(8337));
    layer2_outputs(5098) <= not(layer1_outputs(333)) or (layer1_outputs(5171));
    layer2_outputs(5099) <= not(layer1_outputs(6437)) or (layer1_outputs(7546));
    layer2_outputs(5100) <= layer1_outputs(11129);
    layer2_outputs(5101) <= not(layer1_outputs(7837)) or (layer1_outputs(7138));
    layer2_outputs(5102) <= (layer1_outputs(4352)) or (layer1_outputs(1174));
    layer2_outputs(5103) <= (layer1_outputs(3891)) and not (layer1_outputs(10118));
    layer2_outputs(5104) <= layer1_outputs(4943);
    layer2_outputs(5105) <= (layer1_outputs(5332)) xor (layer1_outputs(2424));
    layer2_outputs(5106) <= not(layer1_outputs(8825)) or (layer1_outputs(10199));
    layer2_outputs(5107) <= (layer1_outputs(2052)) xor (layer1_outputs(8891));
    layer2_outputs(5108) <= layer1_outputs(8192);
    layer2_outputs(5109) <= not(layer1_outputs(11925));
    layer2_outputs(5110) <= not((layer1_outputs(1262)) xor (layer1_outputs(478)));
    layer2_outputs(5111) <= layer1_outputs(6702);
    layer2_outputs(5112) <= (layer1_outputs(10927)) and not (layer1_outputs(9797));
    layer2_outputs(5113) <= not(layer1_outputs(2759));
    layer2_outputs(5114) <= (layer1_outputs(8754)) xor (layer1_outputs(7478));
    layer2_outputs(5115) <= (layer1_outputs(5683)) or (layer1_outputs(4762));
    layer2_outputs(5116) <= not(layer1_outputs(9908));
    layer2_outputs(5117) <= not(layer1_outputs(5673));
    layer2_outputs(5118) <= layer1_outputs(10070);
    layer2_outputs(5119) <= not(layer1_outputs(11665));
    layer2_outputs(5120) <= not(layer1_outputs(10532)) or (layer1_outputs(9423));
    layer2_outputs(5121) <= (layer1_outputs(9155)) xor (layer1_outputs(6848));
    layer2_outputs(5122) <= layer1_outputs(12228);
    layer2_outputs(5123) <= not((layer1_outputs(4663)) xor (layer1_outputs(4353)));
    layer2_outputs(5124) <= not(layer1_outputs(10451));
    layer2_outputs(5125) <= not(layer1_outputs(11841)) or (layer1_outputs(12219));
    layer2_outputs(5126) <= not(layer1_outputs(7768));
    layer2_outputs(5127) <= (layer1_outputs(10347)) and not (layer1_outputs(2211));
    layer2_outputs(5128) <= layer1_outputs(12410);
    layer2_outputs(5129) <= not(layer1_outputs(298));
    layer2_outputs(5130) <= '0';
    layer2_outputs(5131) <= layer1_outputs(5838);
    layer2_outputs(5132) <= (layer1_outputs(6320)) xor (layer1_outputs(11231));
    layer2_outputs(5133) <= layer1_outputs(12741);
    layer2_outputs(5134) <= layer1_outputs(12760);
    layer2_outputs(5135) <= layer1_outputs(11307);
    layer2_outputs(5136) <= layer1_outputs(6718);
    layer2_outputs(5137) <= layer1_outputs(2726);
    layer2_outputs(5138) <= not(layer1_outputs(10926));
    layer2_outputs(5139) <= not(layer1_outputs(2220));
    layer2_outputs(5140) <= layer1_outputs(3211);
    layer2_outputs(5141) <= (layer1_outputs(3289)) and not (layer1_outputs(1911));
    layer2_outputs(5142) <= not(layer1_outputs(3404));
    layer2_outputs(5143) <= (layer1_outputs(10303)) xor (layer1_outputs(7703));
    layer2_outputs(5144) <= not((layer1_outputs(2523)) xor (layer1_outputs(1840)));
    layer2_outputs(5145) <= not(layer1_outputs(6688)) or (layer1_outputs(1377));
    layer2_outputs(5146) <= not(layer1_outputs(7645));
    layer2_outputs(5147) <= not((layer1_outputs(9956)) xor (layer1_outputs(3390)));
    layer2_outputs(5148) <= layer1_outputs(7003);
    layer2_outputs(5149) <= (layer1_outputs(3015)) and not (layer1_outputs(10489));
    layer2_outputs(5150) <= not(layer1_outputs(5963)) or (layer1_outputs(12089));
    layer2_outputs(5151) <= layer1_outputs(4271);
    layer2_outputs(5152) <= not((layer1_outputs(2784)) xor (layer1_outputs(5218)));
    layer2_outputs(5153) <= layer1_outputs(11545);
    layer2_outputs(5154) <= (layer1_outputs(10981)) xor (layer1_outputs(7537));
    layer2_outputs(5155) <= not((layer1_outputs(12600)) xor (layer1_outputs(917)));
    layer2_outputs(5156) <= not(layer1_outputs(8634));
    layer2_outputs(5157) <= layer1_outputs(1198);
    layer2_outputs(5158) <= not(layer1_outputs(11806));
    layer2_outputs(5159) <= layer1_outputs(6704);
    layer2_outputs(5160) <= (layer1_outputs(12337)) xor (layer1_outputs(6482));
    layer2_outputs(5161) <= (layer1_outputs(9358)) xor (layer1_outputs(5764));
    layer2_outputs(5162) <= (layer1_outputs(10331)) and (layer1_outputs(10484));
    layer2_outputs(5163) <= layer1_outputs(8327);
    layer2_outputs(5164) <= not((layer1_outputs(12647)) xor (layer1_outputs(10916)));
    layer2_outputs(5165) <= layer1_outputs(6483);
    layer2_outputs(5166) <= not(layer1_outputs(11074)) or (layer1_outputs(7345));
    layer2_outputs(5167) <= (layer1_outputs(2914)) xor (layer1_outputs(447));
    layer2_outputs(5168) <= not((layer1_outputs(7754)) and (layer1_outputs(8094)));
    layer2_outputs(5169) <= layer1_outputs(1655);
    layer2_outputs(5170) <= not(layer1_outputs(4330));
    layer2_outputs(5171) <= not(layer1_outputs(7572));
    layer2_outputs(5172) <= layer1_outputs(6932);
    layer2_outputs(5173) <= layer1_outputs(4593);
    layer2_outputs(5174) <= not((layer1_outputs(382)) xor (layer1_outputs(11794)));
    layer2_outputs(5175) <= not(layer1_outputs(5722));
    layer2_outputs(5176) <= layer1_outputs(326);
    layer2_outputs(5177) <= not((layer1_outputs(9393)) or (layer1_outputs(5596)));
    layer2_outputs(5178) <= not(layer1_outputs(2900)) or (layer1_outputs(11380));
    layer2_outputs(5179) <= layer1_outputs(1180);
    layer2_outputs(5180) <= not(layer1_outputs(301));
    layer2_outputs(5181) <= not(layer1_outputs(8254)) or (layer1_outputs(3528));
    layer2_outputs(5182) <= (layer1_outputs(336)) xor (layer1_outputs(10843));
    layer2_outputs(5183) <= (layer1_outputs(2113)) xor (layer1_outputs(9029));
    layer2_outputs(5184) <= not(layer1_outputs(5496));
    layer2_outputs(5185) <= layer1_outputs(12788);
    layer2_outputs(5186) <= not(layer1_outputs(931)) or (layer1_outputs(10536));
    layer2_outputs(5187) <= not((layer1_outputs(7685)) or (layer1_outputs(3551)));
    layer2_outputs(5188) <= (layer1_outputs(5021)) xor (layer1_outputs(3364));
    layer2_outputs(5189) <= not(layer1_outputs(4927)) or (layer1_outputs(4815));
    layer2_outputs(5190) <= not((layer1_outputs(3673)) xor (layer1_outputs(4216)));
    layer2_outputs(5191) <= layer1_outputs(8145);
    layer2_outputs(5192) <= not(layer1_outputs(6082));
    layer2_outputs(5193) <= layer1_outputs(5892);
    layer2_outputs(5194) <= not(layer1_outputs(2126)) or (layer1_outputs(10761));
    layer2_outputs(5195) <= not(layer1_outputs(11600));
    layer2_outputs(5196) <= (layer1_outputs(11943)) xor (layer1_outputs(72));
    layer2_outputs(5197) <= not((layer1_outputs(395)) xor (layer1_outputs(5174)));
    layer2_outputs(5198) <= (layer1_outputs(2028)) and (layer1_outputs(367));
    layer2_outputs(5199) <= not(layer1_outputs(12677));
    layer2_outputs(5200) <= layer1_outputs(10123);
    layer2_outputs(5201) <= layer1_outputs(5311);
    layer2_outputs(5202) <= not(layer1_outputs(3178)) or (layer1_outputs(7232));
    layer2_outputs(5203) <= not(layer1_outputs(8705));
    layer2_outputs(5204) <= not(layer1_outputs(10568)) or (layer1_outputs(7084));
    layer2_outputs(5205) <= not(layer1_outputs(6279));
    layer2_outputs(5206) <= layer1_outputs(10713);
    layer2_outputs(5207) <= not(layer1_outputs(1058));
    layer2_outputs(5208) <= not(layer1_outputs(1882));
    layer2_outputs(5209) <= not((layer1_outputs(11461)) and (layer1_outputs(5006)));
    layer2_outputs(5210) <= not((layer1_outputs(267)) and (layer1_outputs(3119)));
    layer2_outputs(5211) <= layer1_outputs(5794);
    layer2_outputs(5212) <= (layer1_outputs(8554)) xor (layer1_outputs(3724));
    layer2_outputs(5213) <= (layer1_outputs(11107)) and (layer1_outputs(8560));
    layer2_outputs(5214) <= not(layer1_outputs(3034));
    layer2_outputs(5215) <= layer1_outputs(7189);
    layer2_outputs(5216) <= not((layer1_outputs(2976)) or (layer1_outputs(1414)));
    layer2_outputs(5217) <= layer1_outputs(210);
    layer2_outputs(5218) <= (layer1_outputs(7793)) and not (layer1_outputs(8410));
    layer2_outputs(5219) <= (layer1_outputs(10053)) and not (layer1_outputs(9040));
    layer2_outputs(5220) <= not(layer1_outputs(3026));
    layer2_outputs(5221) <= (layer1_outputs(7682)) xor (layer1_outputs(9078));
    layer2_outputs(5222) <= not(layer1_outputs(5475)) or (layer1_outputs(6682));
    layer2_outputs(5223) <= not(layer1_outputs(7456)) or (layer1_outputs(6420));
    layer2_outputs(5224) <= layer1_outputs(311);
    layer2_outputs(5225) <= (layer1_outputs(6591)) or (layer1_outputs(8156));
    layer2_outputs(5226) <= not(layer1_outputs(2701));
    layer2_outputs(5227) <= not(layer1_outputs(4117));
    layer2_outputs(5228) <= layer1_outputs(12525);
    layer2_outputs(5229) <= not(layer1_outputs(1872));
    layer2_outputs(5230) <= not((layer1_outputs(7504)) and (layer1_outputs(11463)));
    layer2_outputs(5231) <= not((layer1_outputs(12014)) and (layer1_outputs(5904)));
    layer2_outputs(5232) <= (layer1_outputs(1772)) and (layer1_outputs(7209));
    layer2_outputs(5233) <= not(layer1_outputs(12635));
    layer2_outputs(5234) <= layer1_outputs(6124);
    layer2_outputs(5235) <= (layer1_outputs(12009)) or (layer1_outputs(6997));
    layer2_outputs(5236) <= not((layer1_outputs(9717)) or (layer1_outputs(3359)));
    layer2_outputs(5237) <= layer1_outputs(682);
    layer2_outputs(5238) <= (layer1_outputs(11206)) or (layer1_outputs(2690));
    layer2_outputs(5239) <= not(layer1_outputs(12292)) or (layer1_outputs(1383));
    layer2_outputs(5240) <= layer1_outputs(387);
    layer2_outputs(5241) <= (layer1_outputs(12662)) or (layer1_outputs(5636));
    layer2_outputs(5242) <= not(layer1_outputs(7933));
    layer2_outputs(5243) <= not((layer1_outputs(10411)) or (layer1_outputs(12066)));
    layer2_outputs(5244) <= not(layer1_outputs(9496)) or (layer1_outputs(5744));
    layer2_outputs(5245) <= not(layer1_outputs(11264));
    layer2_outputs(5246) <= layer1_outputs(11144);
    layer2_outputs(5247) <= not((layer1_outputs(321)) or (layer1_outputs(10113)));
    layer2_outputs(5248) <= not(layer1_outputs(10244));
    layer2_outputs(5249) <= layer1_outputs(172);
    layer2_outputs(5250) <= not((layer1_outputs(10680)) xor (layer1_outputs(5287)));
    layer2_outputs(5251) <= layer1_outputs(12124);
    layer2_outputs(5252) <= not(layer1_outputs(12707)) or (layer1_outputs(4620));
    layer2_outputs(5253) <= layer1_outputs(5684);
    layer2_outputs(5254) <= not(layer1_outputs(7154));
    layer2_outputs(5255) <= (layer1_outputs(1704)) and not (layer1_outputs(3942));
    layer2_outputs(5256) <= not(layer1_outputs(531));
    layer2_outputs(5257) <= layer1_outputs(3781);
    layer2_outputs(5258) <= (layer1_outputs(4512)) and not (layer1_outputs(3031));
    layer2_outputs(5259) <= (layer1_outputs(8379)) or (layer1_outputs(3041));
    layer2_outputs(5260) <= not(layer1_outputs(12592));
    layer2_outputs(5261) <= not((layer1_outputs(12450)) xor (layer1_outputs(5219)));
    layer2_outputs(5262) <= not((layer1_outputs(8409)) and (layer1_outputs(12783)));
    layer2_outputs(5263) <= (layer1_outputs(8878)) and not (layer1_outputs(12067));
    layer2_outputs(5264) <= not(layer1_outputs(11589));
    layer2_outputs(5265) <= not(layer1_outputs(9486));
    layer2_outputs(5266) <= not((layer1_outputs(10530)) and (layer1_outputs(10189)));
    layer2_outputs(5267) <= not((layer1_outputs(8806)) or (layer1_outputs(8772)));
    layer2_outputs(5268) <= '0';
    layer2_outputs(5269) <= layer1_outputs(4224);
    layer2_outputs(5270) <= not(layer1_outputs(8797));
    layer2_outputs(5271) <= not(layer1_outputs(2436));
    layer2_outputs(5272) <= not(layer1_outputs(9517));
    layer2_outputs(5273) <= layer1_outputs(9279);
    layer2_outputs(5274) <= not(layer1_outputs(4629)) or (layer1_outputs(11331));
    layer2_outputs(5275) <= not((layer1_outputs(10556)) and (layer1_outputs(5919)));
    layer2_outputs(5276) <= (layer1_outputs(7901)) xor (layer1_outputs(1596));
    layer2_outputs(5277) <= layer1_outputs(7998);
    layer2_outputs(5278) <= not(layer1_outputs(20));
    layer2_outputs(5279) <= (layer1_outputs(4899)) and not (layer1_outputs(8663));
    layer2_outputs(5280) <= not((layer1_outputs(12329)) and (layer1_outputs(417)));
    layer2_outputs(5281) <= layer1_outputs(965);
    layer2_outputs(5282) <= not(layer1_outputs(833));
    layer2_outputs(5283) <= (layer1_outputs(10529)) and not (layer1_outputs(4151));
    layer2_outputs(5284) <= layer1_outputs(12141);
    layer2_outputs(5285) <= not((layer1_outputs(6780)) and (layer1_outputs(1784)));
    layer2_outputs(5286) <= (layer1_outputs(3324)) and not (layer1_outputs(6424));
    layer2_outputs(5287) <= layer1_outputs(1230);
    layer2_outputs(5288) <= not(layer1_outputs(6700));
    layer2_outputs(5289) <= not(layer1_outputs(6721));
    layer2_outputs(5290) <= not(layer1_outputs(10622));
    layer2_outputs(5291) <= not(layer1_outputs(12229)) or (layer1_outputs(5261));
    layer2_outputs(5292) <= not(layer1_outputs(5997));
    layer2_outputs(5293) <= layer1_outputs(6043);
    layer2_outputs(5294) <= not(layer1_outputs(11363));
    layer2_outputs(5295) <= not(layer1_outputs(9212)) or (layer1_outputs(3965));
    layer2_outputs(5296) <= layer1_outputs(1730);
    layer2_outputs(5297) <= layer1_outputs(7199);
    layer2_outputs(5298) <= (layer1_outputs(11804)) and not (layer1_outputs(8500));
    layer2_outputs(5299) <= not((layer1_outputs(1061)) and (layer1_outputs(3414)));
    layer2_outputs(5300) <= not((layer1_outputs(10410)) xor (layer1_outputs(8726)));
    layer2_outputs(5301) <= layer1_outputs(1444);
    layer2_outputs(5302) <= layer1_outputs(5177);
    layer2_outputs(5303) <= layer1_outputs(7300);
    layer2_outputs(5304) <= not((layer1_outputs(7017)) and (layer1_outputs(3322)));
    layer2_outputs(5305) <= not(layer1_outputs(5446)) or (layer1_outputs(9059));
    layer2_outputs(5306) <= not(layer1_outputs(8820));
    layer2_outputs(5307) <= layer1_outputs(1353);
    layer2_outputs(5308) <= not((layer1_outputs(9791)) xor (layer1_outputs(9363)));
    layer2_outputs(5309) <= layer1_outputs(7469);
    layer2_outputs(5310) <= (layer1_outputs(6293)) and (layer1_outputs(3204));
    layer2_outputs(5311) <= not(layer1_outputs(10779));
    layer2_outputs(5312) <= (layer1_outputs(1035)) and (layer1_outputs(1993));
    layer2_outputs(5313) <= not(layer1_outputs(11762));
    layer2_outputs(5314) <= (layer1_outputs(2250)) xor (layer1_outputs(8902));
    layer2_outputs(5315) <= not((layer1_outputs(11065)) and (layer1_outputs(10358)));
    layer2_outputs(5316) <= layer1_outputs(219);
    layer2_outputs(5317) <= not(layer1_outputs(12732));
    layer2_outputs(5318) <= (layer1_outputs(10643)) xor (layer1_outputs(902));
    layer2_outputs(5319) <= layer1_outputs(6190);
    layer2_outputs(5320) <= (layer1_outputs(4470)) xor (layer1_outputs(1156));
    layer2_outputs(5321) <= layer1_outputs(5874);
    layer2_outputs(5322) <= not(layer1_outputs(1453));
    layer2_outputs(5323) <= (layer1_outputs(9546)) xor (layer1_outputs(412));
    layer2_outputs(5324) <= (layer1_outputs(1424)) or (layer1_outputs(4757));
    layer2_outputs(5325) <= not(layer1_outputs(10550));
    layer2_outputs(5326) <= not((layer1_outputs(8842)) xor (layer1_outputs(12440)));
    layer2_outputs(5327) <= not(layer1_outputs(8354));
    layer2_outputs(5328) <= (layer1_outputs(38)) and (layer1_outputs(3263));
    layer2_outputs(5329) <= (layer1_outputs(11927)) xor (layer1_outputs(7326));
    layer2_outputs(5330) <= not(layer1_outputs(7072));
    layer2_outputs(5331) <= (layer1_outputs(4024)) and (layer1_outputs(1425));
    layer2_outputs(5332) <= layer1_outputs(4655);
    layer2_outputs(5333) <= not(layer1_outputs(8146)) or (layer1_outputs(6739));
    layer2_outputs(5334) <= not((layer1_outputs(1792)) and (layer1_outputs(11108)));
    layer2_outputs(5335) <= not(layer1_outputs(5229));
    layer2_outputs(5336) <= not(layer1_outputs(8531)) or (layer1_outputs(11816));
    layer2_outputs(5337) <= (layer1_outputs(2933)) and not (layer1_outputs(12278));
    layer2_outputs(5338) <= not(layer1_outputs(1803)) or (layer1_outputs(736));
    layer2_outputs(5339) <= not(layer1_outputs(11163));
    layer2_outputs(5340) <= (layer1_outputs(8673)) and (layer1_outputs(61));
    layer2_outputs(5341) <= not((layer1_outputs(9447)) xor (layer1_outputs(1494)));
    layer2_outputs(5342) <= not(layer1_outputs(7728));
    layer2_outputs(5343) <= not(layer1_outputs(6811));
    layer2_outputs(5344) <= not(layer1_outputs(8036));
    layer2_outputs(5345) <= (layer1_outputs(11797)) xor (layer1_outputs(4551));
    layer2_outputs(5346) <= not(layer1_outputs(1656));
    layer2_outputs(5347) <= not(layer1_outputs(5170));
    layer2_outputs(5348) <= (layer1_outputs(5774)) and (layer1_outputs(8513));
    layer2_outputs(5349) <= not((layer1_outputs(9910)) and (layer1_outputs(1360)));
    layer2_outputs(5350) <= (layer1_outputs(2296)) xor (layer1_outputs(2768));
    layer2_outputs(5351) <= (layer1_outputs(5007)) and not (layer1_outputs(11434));
    layer2_outputs(5352) <= layer1_outputs(6382);
    layer2_outputs(5353) <= (layer1_outputs(3395)) or (layer1_outputs(2337));
    layer2_outputs(5354) <= (layer1_outputs(3143)) xor (layer1_outputs(12075));
    layer2_outputs(5355) <= layer1_outputs(10170);
    layer2_outputs(5356) <= layer1_outputs(2199);
    layer2_outputs(5357) <= layer1_outputs(12680);
    layer2_outputs(5358) <= (layer1_outputs(2136)) and not (layer1_outputs(12770));
    layer2_outputs(5359) <= (layer1_outputs(998)) and not (layer1_outputs(3627));
    layer2_outputs(5360) <= layer1_outputs(4227);
    layer2_outputs(5361) <= (layer1_outputs(12524)) and not (layer1_outputs(11547));
    layer2_outputs(5362) <= not(layer1_outputs(11735));
    layer2_outputs(5363) <= not(layer1_outputs(9201));
    layer2_outputs(5364) <= not(layer1_outputs(4174));
    layer2_outputs(5365) <= (layer1_outputs(3442)) and (layer1_outputs(9121));
    layer2_outputs(5366) <= not(layer1_outputs(7934));
    layer2_outputs(5367) <= (layer1_outputs(2545)) or (layer1_outputs(6447));
    layer2_outputs(5368) <= layer1_outputs(8808);
    layer2_outputs(5369) <= not(layer1_outputs(10915));
    layer2_outputs(5370) <= not((layer1_outputs(9174)) xor (layer1_outputs(9317)));
    layer2_outputs(5371) <= (layer1_outputs(4385)) and not (layer1_outputs(2681));
    layer2_outputs(5372) <= (layer1_outputs(1150)) and not (layer1_outputs(2343));
    layer2_outputs(5373) <= (layer1_outputs(8111)) or (layer1_outputs(134));
    layer2_outputs(5374) <= not((layer1_outputs(5119)) or (layer1_outputs(4425)));
    layer2_outputs(5375) <= not(layer1_outputs(3429));
    layer2_outputs(5376) <= layer1_outputs(11776);
    layer2_outputs(5377) <= layer1_outputs(2);
    layer2_outputs(5378) <= layer1_outputs(11714);
    layer2_outputs(5379) <= not((layer1_outputs(1116)) and (layer1_outputs(5929)));
    layer2_outputs(5380) <= layer1_outputs(10326);
    layer2_outputs(5381) <= not(layer1_outputs(1767)) or (layer1_outputs(1407));
    layer2_outputs(5382) <= (layer1_outputs(7769)) xor (layer1_outputs(6631));
    layer2_outputs(5383) <= not(layer1_outputs(7897));
    layer2_outputs(5384) <= layer1_outputs(5152);
    layer2_outputs(5385) <= (layer1_outputs(6307)) xor (layer1_outputs(401));
    layer2_outputs(5386) <= (layer1_outputs(4846)) or (layer1_outputs(10312));
    layer2_outputs(5387) <= layer1_outputs(10262);
    layer2_outputs(5388) <= layer1_outputs(5514);
    layer2_outputs(5389) <= not(layer1_outputs(9886));
    layer2_outputs(5390) <= not(layer1_outputs(12463));
    layer2_outputs(5391) <= not(layer1_outputs(1628));
    layer2_outputs(5392) <= (layer1_outputs(1788)) and (layer1_outputs(11902));
    layer2_outputs(5393) <= not(layer1_outputs(2148));
    layer2_outputs(5394) <= layer1_outputs(5841);
    layer2_outputs(5395) <= not(layer1_outputs(12585));
    layer2_outputs(5396) <= layer1_outputs(2198);
    layer2_outputs(5397) <= (layer1_outputs(6716)) or (layer1_outputs(3501));
    layer2_outputs(5398) <= not((layer1_outputs(7256)) and (layer1_outputs(2478)));
    layer2_outputs(5399) <= (layer1_outputs(5943)) xor (layer1_outputs(7248));
    layer2_outputs(5400) <= not(layer1_outputs(7922));
    layer2_outputs(5401) <= (layer1_outputs(5689)) or (layer1_outputs(444));
    layer2_outputs(5402) <= not(layer1_outputs(5199));
    layer2_outputs(5403) <= not(layer1_outputs(5632));
    layer2_outputs(5404) <= (layer1_outputs(10937)) and not (layer1_outputs(4028));
    layer2_outputs(5405) <= not((layer1_outputs(10609)) and (layer1_outputs(3010)));
    layer2_outputs(5406) <= not((layer1_outputs(8250)) and (layer1_outputs(8)));
    layer2_outputs(5407) <= not(layer1_outputs(4445)) or (layer1_outputs(78));
    layer2_outputs(5408) <= (layer1_outputs(9972)) xor (layer1_outputs(10634));
    layer2_outputs(5409) <= layer1_outputs(9990);
    layer2_outputs(5410) <= layer1_outputs(19);
    layer2_outputs(5411) <= not(layer1_outputs(12373)) or (layer1_outputs(3167));
    layer2_outputs(5412) <= not(layer1_outputs(1319)) or (layer1_outputs(9131));
    layer2_outputs(5413) <= layer1_outputs(8022);
    layer2_outputs(5414) <= layer1_outputs(2159);
    layer2_outputs(5415) <= not(layer1_outputs(6726));
    layer2_outputs(5416) <= not((layer1_outputs(6475)) and (layer1_outputs(7040)));
    layer2_outputs(5417) <= layer1_outputs(11472);
    layer2_outputs(5418) <= not(layer1_outputs(10917));
    layer2_outputs(5419) <= not(layer1_outputs(6001));
    layer2_outputs(5420) <= (layer1_outputs(7231)) or (layer1_outputs(12217));
    layer2_outputs(5421) <= (layer1_outputs(12482)) and not (layer1_outputs(11267));
    layer2_outputs(5422) <= layer1_outputs(9949);
    layer2_outputs(5423) <= layer1_outputs(504);
    layer2_outputs(5424) <= not(layer1_outputs(1669));
    layer2_outputs(5425) <= layer1_outputs(3045);
    layer2_outputs(5426) <= not((layer1_outputs(1565)) or (layer1_outputs(3095)));
    layer2_outputs(5427) <= layer1_outputs(2380);
    layer2_outputs(5428) <= layer1_outputs(1019);
    layer2_outputs(5429) <= (layer1_outputs(10062)) and not (layer1_outputs(3169));
    layer2_outputs(5430) <= not(layer1_outputs(2563));
    layer2_outputs(5431) <= layer1_outputs(10286);
    layer2_outputs(5432) <= layer1_outputs(4186);
    layer2_outputs(5433) <= not(layer1_outputs(9904));
    layer2_outputs(5434) <= not(layer1_outputs(2305));
    layer2_outputs(5435) <= not(layer1_outputs(6167));
    layer2_outputs(5436) <= not(layer1_outputs(6873)) or (layer1_outputs(1962));
    layer2_outputs(5437) <= not(layer1_outputs(3667));
    layer2_outputs(5438) <= (layer1_outputs(6049)) and not (layer1_outputs(6101));
    layer2_outputs(5439) <= (layer1_outputs(5123)) and not (layer1_outputs(12102));
    layer2_outputs(5440) <= not((layer1_outputs(806)) xor (layer1_outputs(2465)));
    layer2_outputs(5441) <= layer1_outputs(10710);
    layer2_outputs(5442) <= not((layer1_outputs(287)) or (layer1_outputs(4948)));
    layer2_outputs(5443) <= layer1_outputs(7180);
    layer2_outputs(5444) <= layer1_outputs(5183);
    layer2_outputs(5445) <= not(layer1_outputs(6473));
    layer2_outputs(5446) <= (layer1_outputs(12133)) and not (layer1_outputs(1944));
    layer2_outputs(5447) <= not(layer1_outputs(2099)) or (layer1_outputs(8335));
    layer2_outputs(5448) <= not(layer1_outputs(8600));
    layer2_outputs(5449) <= (layer1_outputs(5158)) and not (layer1_outputs(7659));
    layer2_outputs(5450) <= layer1_outputs(9084);
    layer2_outputs(5451) <= (layer1_outputs(153)) and not (layer1_outputs(3942));
    layer2_outputs(5452) <= not(layer1_outputs(4482));
    layer2_outputs(5453) <= layer1_outputs(2852);
    layer2_outputs(5454) <= not(layer1_outputs(7745));
    layer2_outputs(5455) <= layer1_outputs(4895);
    layer2_outputs(5456) <= not(layer1_outputs(4010)) or (layer1_outputs(5945));
    layer2_outputs(5457) <= (layer1_outputs(8620)) or (layer1_outputs(11437));
    layer2_outputs(5458) <= layer1_outputs(285);
    layer2_outputs(5459) <= not(layer1_outputs(1873));
    layer2_outputs(5460) <= layer1_outputs(6922);
    layer2_outputs(5461) <= not(layer1_outputs(5651)) or (layer1_outputs(11101));
    layer2_outputs(5462) <= not(layer1_outputs(12248));
    layer2_outputs(5463) <= not(layer1_outputs(1207));
    layer2_outputs(5464) <= (layer1_outputs(5159)) and (layer1_outputs(6245));
    layer2_outputs(5465) <= layer1_outputs(6865);
    layer2_outputs(5466) <= layer1_outputs(11504);
    layer2_outputs(5467) <= not(layer1_outputs(11921)) or (layer1_outputs(12296));
    layer2_outputs(5468) <= not((layer1_outputs(1244)) or (layer1_outputs(9718)));
    layer2_outputs(5469) <= not(layer1_outputs(9343));
    layer2_outputs(5470) <= layer1_outputs(4702);
    layer2_outputs(5471) <= (layer1_outputs(2654)) xor (layer1_outputs(8685));
    layer2_outputs(5472) <= layer1_outputs(4427);
    layer2_outputs(5473) <= '0';
    layer2_outputs(5474) <= (layer1_outputs(12689)) and not (layer1_outputs(11498));
    layer2_outputs(5475) <= not(layer1_outputs(1769));
    layer2_outputs(5476) <= layer1_outputs(1119);
    layer2_outputs(5477) <= layer1_outputs(9997);
    layer2_outputs(5478) <= layer1_outputs(6492);
    layer2_outputs(5479) <= not((layer1_outputs(9629)) xor (layer1_outputs(962)));
    layer2_outputs(5480) <= not(layer1_outputs(11700)) or (layer1_outputs(7752));
    layer2_outputs(5481) <= (layer1_outputs(5965)) or (layer1_outputs(5551));
    layer2_outputs(5482) <= layer1_outputs(11834);
    layer2_outputs(5483) <= not((layer1_outputs(8918)) and (layer1_outputs(12381)));
    layer2_outputs(5484) <= not(layer1_outputs(4710)) or (layer1_outputs(482));
    layer2_outputs(5485) <= (layer1_outputs(11249)) or (layer1_outputs(10918));
    layer2_outputs(5486) <= not(layer1_outputs(10974));
    layer2_outputs(5487) <= not(layer1_outputs(12285)) or (layer1_outputs(3608));
    layer2_outputs(5488) <= not(layer1_outputs(8757)) or (layer1_outputs(6064));
    layer2_outputs(5489) <= not((layer1_outputs(6185)) xor (layer1_outputs(12793)));
    layer2_outputs(5490) <= layer1_outputs(9421);
    layer2_outputs(5491) <= (layer1_outputs(11505)) xor (layer1_outputs(8271));
    layer2_outputs(5492) <= (layer1_outputs(1472)) and not (layer1_outputs(7112));
    layer2_outputs(5493) <= not(layer1_outputs(11791));
    layer2_outputs(5494) <= layer1_outputs(2999);
    layer2_outputs(5495) <= layer1_outputs(11276);
    layer2_outputs(5496) <= (layer1_outputs(4409)) xor (layer1_outputs(5457));
    layer2_outputs(5497) <= layer1_outputs(2499);
    layer2_outputs(5498) <= layer1_outputs(11081);
    layer2_outputs(5499) <= (layer1_outputs(3023)) or (layer1_outputs(2700));
    layer2_outputs(5500) <= layer1_outputs(1056);
    layer2_outputs(5501) <= not(layer1_outputs(11575));
    layer2_outputs(5502) <= (layer1_outputs(2781)) or (layer1_outputs(633));
    layer2_outputs(5503) <= layer1_outputs(4823);
    layer2_outputs(5504) <= (layer1_outputs(11086)) and not (layer1_outputs(2621));
    layer2_outputs(5505) <= not((layer1_outputs(8824)) xor (layer1_outputs(4575)));
    layer2_outputs(5506) <= not((layer1_outputs(3254)) and (layer1_outputs(869)));
    layer2_outputs(5507) <= (layer1_outputs(4449)) and (layer1_outputs(828));
    layer2_outputs(5508) <= (layer1_outputs(10525)) and (layer1_outputs(5535));
    layer2_outputs(5509) <= not(layer1_outputs(9936)) or (layer1_outputs(5087));
    layer2_outputs(5510) <= not((layer1_outputs(8921)) xor (layer1_outputs(8629)));
    layer2_outputs(5511) <= (layer1_outputs(6478)) and (layer1_outputs(6282));
    layer2_outputs(5512) <= (layer1_outputs(7797)) and not (layer1_outputs(4176));
    layer2_outputs(5513) <= (layer1_outputs(8731)) xor (layer1_outputs(10091));
    layer2_outputs(5514) <= (layer1_outputs(12604)) xor (layer1_outputs(10972));
    layer2_outputs(5515) <= layer1_outputs(8823);
    layer2_outputs(5516) <= not(layer1_outputs(5459));
    layer2_outputs(5517) <= not(layer1_outputs(1458));
    layer2_outputs(5518) <= layer1_outputs(5126);
    layer2_outputs(5519) <= not((layer1_outputs(9695)) or (layer1_outputs(11272)));
    layer2_outputs(5520) <= layer1_outputs(9491);
    layer2_outputs(5521) <= (layer1_outputs(11275)) xor (layer1_outputs(1696));
    layer2_outputs(5522) <= not((layer1_outputs(6193)) xor (layer1_outputs(12362)));
    layer2_outputs(5523) <= not((layer1_outputs(12573)) or (layer1_outputs(12319)));
    layer2_outputs(5524) <= not((layer1_outputs(2600)) xor (layer1_outputs(4222)));
    layer2_outputs(5525) <= not((layer1_outputs(5146)) xor (layer1_outputs(10713)));
    layer2_outputs(5526) <= (layer1_outputs(4688)) and (layer1_outputs(7556));
    layer2_outputs(5527) <= not(layer1_outputs(311));
    layer2_outputs(5528) <= not(layer1_outputs(6845));
    layer2_outputs(5529) <= layer1_outputs(10982);
    layer2_outputs(5530) <= not(layer1_outputs(4453));
    layer2_outputs(5531) <= not((layer1_outputs(634)) and (layer1_outputs(11042)));
    layer2_outputs(5532) <= layer1_outputs(785);
    layer2_outputs(5533) <= (layer1_outputs(5624)) or (layer1_outputs(8477));
    layer2_outputs(5534) <= not(layer1_outputs(9467));
    layer2_outputs(5535) <= (layer1_outputs(6827)) or (layer1_outputs(180));
    layer2_outputs(5536) <= layer1_outputs(9486);
    layer2_outputs(5537) <= not((layer1_outputs(207)) or (layer1_outputs(7383)));
    layer2_outputs(5538) <= not((layer1_outputs(10044)) or (layer1_outputs(10061)));
    layer2_outputs(5539) <= layer1_outputs(10456);
    layer2_outputs(5540) <= not(layer1_outputs(11928));
    layer2_outputs(5541) <= (layer1_outputs(3279)) and not (layer1_outputs(5905));
    layer2_outputs(5542) <= (layer1_outputs(9783)) and not (layer1_outputs(3114));
    layer2_outputs(5543) <= (layer1_outputs(5695)) or (layer1_outputs(3385));
    layer2_outputs(5544) <= not(layer1_outputs(9364));
    layer2_outputs(5545) <= not(layer1_outputs(9960));
    layer2_outputs(5546) <= not(layer1_outputs(5599));
    layer2_outputs(5547) <= not(layer1_outputs(10901));
    layer2_outputs(5548) <= not((layer1_outputs(2956)) xor (layer1_outputs(4855)));
    layer2_outputs(5549) <= not((layer1_outputs(8785)) or (layer1_outputs(11717)));
    layer2_outputs(5550) <= not((layer1_outputs(9593)) and (layer1_outputs(8135)));
    layer2_outputs(5551) <= not(layer1_outputs(6268));
    layer2_outputs(5552) <= layer1_outputs(8319);
    layer2_outputs(5553) <= (layer1_outputs(2326)) xor (layer1_outputs(12208));
    layer2_outputs(5554) <= not(layer1_outputs(9855));
    layer2_outputs(5555) <= not(layer1_outputs(2167));
    layer2_outputs(5556) <= layer1_outputs(5460);
    layer2_outputs(5557) <= not(layer1_outputs(7075));
    layer2_outputs(5558) <= layer1_outputs(6562);
    layer2_outputs(5559) <= not((layer1_outputs(6657)) xor (layer1_outputs(4354)));
    layer2_outputs(5560) <= (layer1_outputs(6158)) and (layer1_outputs(4698));
    layer2_outputs(5561) <= (layer1_outputs(192)) or (layer1_outputs(3229));
    layer2_outputs(5562) <= layer1_outputs(10675);
    layer2_outputs(5563) <= layer1_outputs(292);
    layer2_outputs(5564) <= layer1_outputs(11953);
    layer2_outputs(5565) <= layer1_outputs(11640);
    layer2_outputs(5566) <= (layer1_outputs(1649)) xor (layer1_outputs(10668));
    layer2_outputs(5567) <= (layer1_outputs(12786)) and not (layer1_outputs(12755));
    layer2_outputs(5568) <= not(layer1_outputs(4848));
    layer2_outputs(5569) <= not(layer1_outputs(10092));
    layer2_outputs(5570) <= not(layer1_outputs(6168));
    layer2_outputs(5571) <= layer1_outputs(1256);
    layer2_outputs(5572) <= (layer1_outputs(3369)) xor (layer1_outputs(1345));
    layer2_outputs(5573) <= layer1_outputs(8879);
    layer2_outputs(5574) <= layer1_outputs(12203);
    layer2_outputs(5575) <= layer1_outputs(1208);
    layer2_outputs(5576) <= not(layer1_outputs(5570));
    layer2_outputs(5577) <= layer1_outputs(5884);
    layer2_outputs(5578) <= not(layer1_outputs(3963));
    layer2_outputs(5579) <= not(layer1_outputs(3923)) or (layer1_outputs(8290));
    layer2_outputs(5580) <= not((layer1_outputs(6687)) and (layer1_outputs(1849)));
    layer2_outputs(5581) <= layer1_outputs(5540);
    layer2_outputs(5582) <= layer1_outputs(3712);
    layer2_outputs(5583) <= layer1_outputs(7685);
    layer2_outputs(5584) <= (layer1_outputs(11093)) xor (layer1_outputs(3246));
    layer2_outputs(5585) <= not(layer1_outputs(11569));
    layer2_outputs(5586) <= layer1_outputs(263);
    layer2_outputs(5587) <= not((layer1_outputs(3194)) xor (layer1_outputs(7675)));
    layer2_outputs(5588) <= (layer1_outputs(10845)) xor (layer1_outputs(515));
    layer2_outputs(5589) <= not(layer1_outputs(10791));
    layer2_outputs(5590) <= (layer1_outputs(10168)) and not (layer1_outputs(11009));
    layer2_outputs(5591) <= (layer1_outputs(10886)) xor (layer1_outputs(1730));
    layer2_outputs(5592) <= not((layer1_outputs(1751)) xor (layer1_outputs(9503)));
    layer2_outputs(5593) <= not(layer1_outputs(717));
    layer2_outputs(5594) <= not((layer1_outputs(5020)) and (layer1_outputs(5833)));
    layer2_outputs(5595) <= (layer1_outputs(10305)) or (layer1_outputs(6782));
    layer2_outputs(5596) <= not(layer1_outputs(2843));
    layer2_outputs(5597) <= not(layer1_outputs(11241));
    layer2_outputs(5598) <= not(layer1_outputs(6790)) or (layer1_outputs(31));
    layer2_outputs(5599) <= not(layer1_outputs(4614));
    layer2_outputs(5600) <= layer1_outputs(9258);
    layer2_outputs(5601) <= not(layer1_outputs(1207));
    layer2_outputs(5602) <= layer1_outputs(12667);
    layer2_outputs(5603) <= not(layer1_outputs(533));
    layer2_outputs(5604) <= layer1_outputs(12757);
    layer2_outputs(5605) <= not(layer1_outputs(6840));
    layer2_outputs(5606) <= not(layer1_outputs(8089));
    layer2_outputs(5607) <= (layer1_outputs(103)) and not (layer1_outputs(5988));
    layer2_outputs(5608) <= layer1_outputs(9160);
    layer2_outputs(5609) <= (layer1_outputs(5866)) xor (layer1_outputs(7755));
    layer2_outputs(5610) <= layer1_outputs(2938);
    layer2_outputs(5611) <= (layer1_outputs(8290)) and not (layer1_outputs(228));
    layer2_outputs(5612) <= not(layer1_outputs(2841));
    layer2_outputs(5613) <= not(layer1_outputs(4000));
    layer2_outputs(5614) <= layer1_outputs(12041);
    layer2_outputs(5615) <= (layer1_outputs(5822)) or (layer1_outputs(2153));
    layer2_outputs(5616) <= not((layer1_outputs(12242)) xor (layer1_outputs(10773)));
    layer2_outputs(5617) <= not(layer1_outputs(11269));
    layer2_outputs(5618) <= not(layer1_outputs(8618));
    layer2_outputs(5619) <= (layer1_outputs(11446)) and not (layer1_outputs(8967));
    layer2_outputs(5620) <= not((layer1_outputs(3498)) or (layer1_outputs(5033)));
    layer2_outputs(5621) <= not(layer1_outputs(2756));
    layer2_outputs(5622) <= not(layer1_outputs(5119));
    layer2_outputs(5623) <= not((layer1_outputs(4013)) and (layer1_outputs(6992)));
    layer2_outputs(5624) <= layer1_outputs(11805);
    layer2_outputs(5625) <= not(layer1_outputs(10782));
    layer2_outputs(5626) <= not(layer1_outputs(11800));
    layer2_outputs(5627) <= (layer1_outputs(6019)) and not (layer1_outputs(1183));
    layer2_outputs(5628) <= not(layer1_outputs(866));
    layer2_outputs(5629) <= not(layer1_outputs(9825)) or (layer1_outputs(4171));
    layer2_outputs(5630) <= (layer1_outputs(10143)) and not (layer1_outputs(2249));
    layer2_outputs(5631) <= not(layer1_outputs(10023));
    layer2_outputs(5632) <= layer1_outputs(10732);
    layer2_outputs(5633) <= layer1_outputs(8676);
    layer2_outputs(5634) <= (layer1_outputs(7980)) and not (layer1_outputs(12194));
    layer2_outputs(5635) <= not((layer1_outputs(6925)) and (layer1_outputs(319)));
    layer2_outputs(5636) <= layer1_outputs(8903);
    layer2_outputs(5637) <= (layer1_outputs(4478)) or (layer1_outputs(8384));
    layer2_outputs(5638) <= not(layer1_outputs(10393));
    layer2_outputs(5639) <= not(layer1_outputs(3233));
    layer2_outputs(5640) <= not(layer1_outputs(7896));
    layer2_outputs(5641) <= not(layer1_outputs(5487));
    layer2_outputs(5642) <= not(layer1_outputs(1759));
    layer2_outputs(5643) <= not(layer1_outputs(8352));
    layer2_outputs(5644) <= (layer1_outputs(7364)) xor (layer1_outputs(7826));
    layer2_outputs(5645) <= not(layer1_outputs(9225));
    layer2_outputs(5646) <= not(layer1_outputs(5678));
    layer2_outputs(5647) <= not(layer1_outputs(2067));
    layer2_outputs(5648) <= not(layer1_outputs(2939));
    layer2_outputs(5649) <= layer1_outputs(11904);
    layer2_outputs(5650) <= not((layer1_outputs(5282)) and (layer1_outputs(8342)));
    layer2_outputs(5651) <= not((layer1_outputs(10241)) or (layer1_outputs(3801)));
    layer2_outputs(5652) <= not(layer1_outputs(7646));
    layer2_outputs(5653) <= (layer1_outputs(6876)) or (layer1_outputs(11416));
    layer2_outputs(5654) <= (layer1_outputs(3945)) xor (layer1_outputs(8932));
    layer2_outputs(5655) <= layer1_outputs(3008);
    layer2_outputs(5656) <= not((layer1_outputs(7253)) xor (layer1_outputs(8416)));
    layer2_outputs(5657) <= (layer1_outputs(9647)) xor (layer1_outputs(3397));
    layer2_outputs(5658) <= not(layer1_outputs(1497));
    layer2_outputs(5659) <= layer1_outputs(10046);
    layer2_outputs(5660) <= not(layer1_outputs(3630));
    layer2_outputs(5661) <= (layer1_outputs(2425)) and (layer1_outputs(3240));
    layer2_outputs(5662) <= not((layer1_outputs(1676)) or (layer1_outputs(284)));
    layer2_outputs(5663) <= not(layer1_outputs(6795));
    layer2_outputs(5664) <= not((layer1_outputs(9632)) and (layer1_outputs(4447)));
    layer2_outputs(5665) <= layer1_outputs(4378);
    layer2_outputs(5666) <= not(layer1_outputs(3170));
    layer2_outputs(5667) <= (layer1_outputs(1271)) and (layer1_outputs(3774));
    layer2_outputs(5668) <= layer1_outputs(3988);
    layer2_outputs(5669) <= (layer1_outputs(5417)) and not (layer1_outputs(3813));
    layer2_outputs(5670) <= layer1_outputs(7729);
    layer2_outputs(5671) <= not(layer1_outputs(7716));
    layer2_outputs(5672) <= not((layer1_outputs(11801)) xor (layer1_outputs(899)));
    layer2_outputs(5673) <= (layer1_outputs(8805)) and not (layer1_outputs(1020));
    layer2_outputs(5674) <= layer1_outputs(11864);
    layer2_outputs(5675) <= not((layer1_outputs(1585)) xor (layer1_outputs(2004)));
    layer2_outputs(5676) <= not(layer1_outputs(39)) or (layer1_outputs(4080));
    layer2_outputs(5677) <= (layer1_outputs(4230)) or (layer1_outputs(1631));
    layer2_outputs(5678) <= layer1_outputs(8080);
    layer2_outputs(5679) <= not(layer1_outputs(12179));
    layer2_outputs(5680) <= layer1_outputs(4868);
    layer2_outputs(5681) <= layer1_outputs(8142);
    layer2_outputs(5682) <= not((layer1_outputs(7358)) xor (layer1_outputs(8091)));
    layer2_outputs(5683) <= not((layer1_outputs(10227)) xor (layer1_outputs(350)));
    layer2_outputs(5684) <= not(layer1_outputs(5757));
    layer2_outputs(5685) <= not(layer1_outputs(12431)) or (layer1_outputs(7889));
    layer2_outputs(5686) <= not(layer1_outputs(7618));
    layer2_outputs(5687) <= not((layer1_outputs(862)) and (layer1_outputs(7201)));
    layer2_outputs(5688) <= (layer1_outputs(9530)) and not (layer1_outputs(8282));
    layer2_outputs(5689) <= (layer1_outputs(7954)) and not (layer1_outputs(12622));
    layer2_outputs(5690) <= not(layer1_outputs(10327));
    layer2_outputs(5691) <= layer1_outputs(11346);
    layer2_outputs(5692) <= not(layer1_outputs(3972));
    layer2_outputs(5693) <= (layer1_outputs(9311)) xor (layer1_outputs(8083));
    layer2_outputs(5694) <= layer1_outputs(11667);
    layer2_outputs(5695) <= not(layer1_outputs(8259));
    layer2_outputs(5696) <= not(layer1_outputs(4585));
    layer2_outputs(5697) <= (layer1_outputs(9922)) or (layer1_outputs(3632));
    layer2_outputs(5698) <= (layer1_outputs(11379)) or (layer1_outputs(8994));
    layer2_outputs(5699) <= not(layer1_outputs(6690));
    layer2_outputs(5700) <= not((layer1_outputs(8487)) or (layer1_outputs(7015)));
    layer2_outputs(5701) <= not(layer1_outputs(8378));
    layer2_outputs(5702) <= (layer1_outputs(12046)) and not (layer1_outputs(1636));
    layer2_outputs(5703) <= not(layer1_outputs(9027));
    layer2_outputs(5704) <= not(layer1_outputs(9814));
    layer2_outputs(5705) <= not((layer1_outputs(8585)) xor (layer1_outputs(9364)));
    layer2_outputs(5706) <= layer1_outputs(358);
    layer2_outputs(5707) <= not((layer1_outputs(486)) and (layer1_outputs(3091)));
    layer2_outputs(5708) <= not(layer1_outputs(9197));
    layer2_outputs(5709) <= layer1_outputs(7681);
    layer2_outputs(5710) <= (layer1_outputs(700)) xor (layer1_outputs(9408));
    layer2_outputs(5711) <= (layer1_outputs(12262)) and (layer1_outputs(12281));
    layer2_outputs(5712) <= layer1_outputs(183);
    layer2_outputs(5713) <= (layer1_outputs(8440)) and (layer1_outputs(8468));
    layer2_outputs(5714) <= (layer1_outputs(2414)) and not (layer1_outputs(8207));
    layer2_outputs(5715) <= (layer1_outputs(3371)) xor (layer1_outputs(7796));
    layer2_outputs(5716) <= (layer1_outputs(9055)) and not (layer1_outputs(6850));
    layer2_outputs(5717) <= not(layer1_outputs(1545)) or (layer1_outputs(4686));
    layer2_outputs(5718) <= not(layer1_outputs(2140));
    layer2_outputs(5719) <= layer1_outputs(8030);
    layer2_outputs(5720) <= not(layer1_outputs(2091));
    layer2_outputs(5721) <= (layer1_outputs(8456)) and not (layer1_outputs(1151));
    layer2_outputs(5722) <= not(layer1_outputs(4179));
    layer2_outputs(5723) <= not((layer1_outputs(4176)) and (layer1_outputs(3809)));
    layer2_outputs(5724) <= layer1_outputs(11833);
    layer2_outputs(5725) <= not((layer1_outputs(8233)) and (layer1_outputs(6784)));
    layer2_outputs(5726) <= not((layer1_outputs(7240)) and (layer1_outputs(3007)));
    layer2_outputs(5727) <= not((layer1_outputs(3382)) xor (layer1_outputs(6720)));
    layer2_outputs(5728) <= layer1_outputs(6819);
    layer2_outputs(5729) <= (layer1_outputs(5532)) or (layer1_outputs(8140));
    layer2_outputs(5730) <= layer1_outputs(2811);
    layer2_outputs(5731) <= (layer1_outputs(6109)) xor (layer1_outputs(9898));
    layer2_outputs(5732) <= not(layer1_outputs(10841));
    layer2_outputs(5733) <= (layer1_outputs(164)) or (layer1_outputs(11187));
    layer2_outputs(5734) <= not((layer1_outputs(7159)) or (layer1_outputs(7201)));
    layer2_outputs(5735) <= layer1_outputs(7971);
    layer2_outputs(5736) <= not(layer1_outputs(7288));
    layer2_outputs(5737) <= not(layer1_outputs(8483)) or (layer1_outputs(2020));
    layer2_outputs(5738) <= layer1_outputs(6942);
    layer2_outputs(5739) <= not(layer1_outputs(3440));
    layer2_outputs(5740) <= not(layer1_outputs(10677)) or (layer1_outputs(1909));
    layer2_outputs(5741) <= not(layer1_outputs(6803));
    layer2_outputs(5742) <= not(layer1_outputs(1105));
    layer2_outputs(5743) <= not(layer1_outputs(11095)) or (layer1_outputs(7531));
    layer2_outputs(5744) <= layer1_outputs(9853);
    layer2_outputs(5745) <= not(layer1_outputs(3122));
    layer2_outputs(5746) <= not(layer1_outputs(8662));
    layer2_outputs(5747) <= not((layer1_outputs(4216)) and (layer1_outputs(329)));
    layer2_outputs(5748) <= not(layer1_outputs(10716)) or (layer1_outputs(12257));
    layer2_outputs(5749) <= not((layer1_outputs(10156)) or (layer1_outputs(7703)));
    layer2_outputs(5750) <= (layer1_outputs(3298)) and (layer1_outputs(5770));
    layer2_outputs(5751) <= layer1_outputs(3304);
    layer2_outputs(5752) <= not((layer1_outputs(2736)) and (layer1_outputs(2149)));
    layer2_outputs(5753) <= layer1_outputs(11624);
    layer2_outputs(5754) <= layer1_outputs(4809);
    layer2_outputs(5755) <= not(layer1_outputs(1951)) or (layer1_outputs(10670));
    layer2_outputs(5756) <= layer1_outputs(5122);
    layer2_outputs(5757) <= layer1_outputs(10236);
    layer2_outputs(5758) <= not(layer1_outputs(3017));
    layer2_outputs(5759) <= layer1_outputs(4464);
    layer2_outputs(5760) <= not((layer1_outputs(8123)) or (layer1_outputs(9384)));
    layer2_outputs(5761) <= (layer1_outputs(9491)) xor (layer1_outputs(10334));
    layer2_outputs(5762) <= layer1_outputs(8323);
    layer2_outputs(5763) <= (layer1_outputs(6624)) and not (layer1_outputs(6281));
    layer2_outputs(5764) <= not(layer1_outputs(541));
    layer2_outputs(5765) <= not(layer1_outputs(4335));
    layer2_outputs(5766) <= (layer1_outputs(4215)) xor (layer1_outputs(2507));
    layer2_outputs(5767) <= layer1_outputs(239);
    layer2_outputs(5768) <= not((layer1_outputs(6534)) xor (layer1_outputs(10144)));
    layer2_outputs(5769) <= (layer1_outputs(7912)) xor (layer1_outputs(5977));
    layer2_outputs(5770) <= (layer1_outputs(2549)) and not (layer1_outputs(11020));
    layer2_outputs(5771) <= not(layer1_outputs(3328));
    layer2_outputs(5772) <= not(layer1_outputs(7614));
    layer2_outputs(5773) <= layer1_outputs(11403);
    layer2_outputs(5774) <= (layer1_outputs(7605)) or (layer1_outputs(2276));
    layer2_outputs(5775) <= not(layer1_outputs(20));
    layer2_outputs(5776) <= not(layer1_outputs(9397));
    layer2_outputs(5777) <= layer1_outputs(4708);
    layer2_outputs(5778) <= not(layer1_outputs(2578));
    layer2_outputs(5779) <= not(layer1_outputs(9776));
    layer2_outputs(5780) <= not((layer1_outputs(1022)) and (layer1_outputs(5782)));
    layer2_outputs(5781) <= layer1_outputs(8830);
    layer2_outputs(5782) <= not((layer1_outputs(4194)) xor (layer1_outputs(1130)));
    layer2_outputs(5783) <= not(layer1_outputs(8790));
    layer2_outputs(5784) <= not(layer1_outputs(4796));
    layer2_outputs(5785) <= layer1_outputs(8774);
    layer2_outputs(5786) <= '0';
    layer2_outputs(5787) <= not((layer1_outputs(4030)) xor (layer1_outputs(1057)));
    layer2_outputs(5788) <= (layer1_outputs(679)) and (layer1_outputs(8816));
    layer2_outputs(5789) <= (layer1_outputs(613)) and (layer1_outputs(9385));
    layer2_outputs(5790) <= not(layer1_outputs(3582));
    layer2_outputs(5791) <= layer1_outputs(8601);
    layer2_outputs(5792) <= (layer1_outputs(2662)) and (layer1_outputs(11989));
    layer2_outputs(5793) <= (layer1_outputs(6980)) and (layer1_outputs(975));
    layer2_outputs(5794) <= (layer1_outputs(9159)) xor (layer1_outputs(1633));
    layer2_outputs(5795) <= not((layer1_outputs(11568)) xor (layer1_outputs(11158)));
    layer2_outputs(5796) <= layer1_outputs(12410);
    layer2_outputs(5797) <= not((layer1_outputs(11344)) and (layer1_outputs(11352)));
    layer2_outputs(5798) <= layer1_outputs(2982);
    layer2_outputs(5799) <= not(layer1_outputs(10983)) or (layer1_outputs(6300));
    layer2_outputs(5800) <= (layer1_outputs(3276)) and not (layer1_outputs(8350));
    layer2_outputs(5801) <= not(layer1_outputs(5534));
    layer2_outputs(5802) <= layer1_outputs(12564);
    layer2_outputs(5803) <= not(layer1_outputs(10124)) or (layer1_outputs(10320));
    layer2_outputs(5804) <= not(layer1_outputs(4819));
    layer2_outputs(5805) <= not((layer1_outputs(7356)) xor (layer1_outputs(4379)));
    layer2_outputs(5806) <= not(layer1_outputs(2139));
    layer2_outputs(5807) <= not(layer1_outputs(4340));
    layer2_outputs(5808) <= layer1_outputs(7448);
    layer2_outputs(5809) <= not(layer1_outputs(9655));
    layer2_outputs(5810) <= not(layer1_outputs(5542));
    layer2_outputs(5811) <= (layer1_outputs(5971)) xor (layer1_outputs(6744));
    layer2_outputs(5812) <= not((layer1_outputs(7412)) and (layer1_outputs(8098)));
    layer2_outputs(5813) <= not(layer1_outputs(10473)) or (layer1_outputs(3795));
    layer2_outputs(5814) <= not(layer1_outputs(2137));
    layer2_outputs(5815) <= layer1_outputs(4315);
    layer2_outputs(5816) <= not(layer1_outputs(1641));
    layer2_outputs(5817) <= (layer1_outputs(12528)) xor (layer1_outputs(4131));
    layer2_outputs(5818) <= (layer1_outputs(2513)) and (layer1_outputs(1384));
    layer2_outputs(5819) <= (layer1_outputs(7406)) xor (layer1_outputs(11353));
    layer2_outputs(5820) <= not(layer1_outputs(11097)) or (layer1_outputs(10343));
    layer2_outputs(5821) <= (layer1_outputs(2187)) and not (layer1_outputs(1120));
    layer2_outputs(5822) <= (layer1_outputs(4557)) or (layer1_outputs(11538));
    layer2_outputs(5823) <= (layer1_outputs(5868)) and not (layer1_outputs(3841));
    layer2_outputs(5824) <= not((layer1_outputs(11920)) or (layer1_outputs(2932)));
    layer2_outputs(5825) <= layer1_outputs(5468);
    layer2_outputs(5826) <= not(layer1_outputs(11767)) or (layer1_outputs(6559));
    layer2_outputs(5827) <= not(layer1_outputs(3794)) or (layer1_outputs(4654));
    layer2_outputs(5828) <= not(layer1_outputs(7304)) or (layer1_outputs(9451));
    layer2_outputs(5829) <= layer1_outputs(10982);
    layer2_outputs(5830) <= (layer1_outputs(7990)) and not (layer1_outputs(5273));
    layer2_outputs(5831) <= (layer1_outputs(12224)) xor (layer1_outputs(5645));
    layer2_outputs(5832) <= (layer1_outputs(1108)) xor (layer1_outputs(7471));
    layer2_outputs(5833) <= layer1_outputs(12722);
    layer2_outputs(5834) <= not(layer1_outputs(7617));
    layer2_outputs(5835) <= layer1_outputs(12321);
    layer2_outputs(5836) <= not(layer1_outputs(4837));
    layer2_outputs(5837) <= (layer1_outputs(5593)) and not (layer1_outputs(3202));
    layer2_outputs(5838) <= not(layer1_outputs(4567));
    layer2_outputs(5839) <= not(layer1_outputs(11557));
    layer2_outputs(5840) <= not(layer1_outputs(8046));
    layer2_outputs(5841) <= (layer1_outputs(8371)) xor (layer1_outputs(3536));
    layer2_outputs(5842) <= (layer1_outputs(2063)) and not (layer1_outputs(8504));
    layer2_outputs(5843) <= not(layer1_outputs(12538));
    layer2_outputs(5844) <= layer1_outputs(6427);
    layer2_outputs(5845) <= layer1_outputs(480);
    layer2_outputs(5846) <= not((layer1_outputs(5184)) and (layer1_outputs(10890)));
    layer2_outputs(5847) <= not(layer1_outputs(2367));
    layer2_outputs(5848) <= layer1_outputs(3207);
    layer2_outputs(5849) <= not(layer1_outputs(10795));
    layer2_outputs(5850) <= layer1_outputs(10443);
    layer2_outputs(5851) <= not((layer1_outputs(11983)) xor (layer1_outputs(1200)));
    layer2_outputs(5852) <= layer1_outputs(1291);
    layer2_outputs(5853) <= layer1_outputs(7208);
    layer2_outputs(5854) <= (layer1_outputs(7376)) and (layer1_outputs(1547));
    layer2_outputs(5855) <= not(layer1_outputs(6809)) or (layer1_outputs(4107));
    layer2_outputs(5856) <= (layer1_outputs(1950)) and not (layer1_outputs(921));
    layer2_outputs(5857) <= not((layer1_outputs(10674)) and (layer1_outputs(12157)));
    layer2_outputs(5858) <= (layer1_outputs(7071)) and not (layer1_outputs(7311));
    layer2_outputs(5859) <= (layer1_outputs(10749)) xor (layer1_outputs(4013));
    layer2_outputs(5860) <= not(layer1_outputs(5682)) or (layer1_outputs(3216));
    layer2_outputs(5861) <= (layer1_outputs(2738)) or (layer1_outputs(5574));
    layer2_outputs(5862) <= not((layer1_outputs(3434)) xor (layer1_outputs(4906)));
    layer2_outputs(5863) <= layer1_outputs(2059);
    layer2_outputs(5864) <= layer1_outputs(2648);
    layer2_outputs(5865) <= (layer1_outputs(1091)) or (layer1_outputs(2166));
    layer2_outputs(5866) <= not((layer1_outputs(12684)) xor (layer1_outputs(2573)));
    layer2_outputs(5867) <= not(layer1_outputs(12739)) or (layer1_outputs(4307));
    layer2_outputs(5868) <= not((layer1_outputs(1767)) or (layer1_outputs(4623)));
    layer2_outputs(5869) <= not((layer1_outputs(4595)) xor (layer1_outputs(12452)));
    layer2_outputs(5870) <= layer1_outputs(3157);
    layer2_outputs(5871) <= not(layer1_outputs(5380));
    layer2_outputs(5872) <= not((layer1_outputs(10517)) and (layer1_outputs(12003)));
    layer2_outputs(5873) <= not(layer1_outputs(5350));
    layer2_outputs(5874) <= not(layer1_outputs(9245));
    layer2_outputs(5875) <= not(layer1_outputs(4583));
    layer2_outputs(5876) <= not(layer1_outputs(7098));
    layer2_outputs(5877) <= not(layer1_outputs(9166)) or (layer1_outputs(1884));
    layer2_outputs(5878) <= not(layer1_outputs(11011));
    layer2_outputs(5879) <= not((layer1_outputs(6925)) or (layer1_outputs(6474)));
    layer2_outputs(5880) <= layer1_outputs(8973);
    layer2_outputs(5881) <= layer1_outputs(1076);
    layer2_outputs(5882) <= not(layer1_outputs(3402));
    layer2_outputs(5883) <= layer1_outputs(2383);
    layer2_outputs(5884) <= layer1_outputs(1727);
    layer2_outputs(5885) <= not((layer1_outputs(10345)) xor (layer1_outputs(6824)));
    layer2_outputs(5886) <= layer1_outputs(12551);
    layer2_outputs(5887) <= (layer1_outputs(8307)) and not (layer1_outputs(1837));
    layer2_outputs(5888) <= (layer1_outputs(5324)) xor (layer1_outputs(68));
    layer2_outputs(5889) <= layer1_outputs(8464);
    layer2_outputs(5890) <= not((layer1_outputs(7109)) xor (layer1_outputs(4058)));
    layer2_outputs(5891) <= (layer1_outputs(10105)) or (layer1_outputs(3047));
    layer2_outputs(5892) <= not(layer1_outputs(8792));
    layer2_outputs(5893) <= layer1_outputs(354);
    layer2_outputs(5894) <= not(layer1_outputs(7738)) or (layer1_outputs(11700));
    layer2_outputs(5895) <= layer1_outputs(2356);
    layer2_outputs(5896) <= not((layer1_outputs(3981)) xor (layer1_outputs(3929)));
    layer2_outputs(5897) <= (layer1_outputs(10589)) xor (layer1_outputs(6537));
    layer2_outputs(5898) <= layer1_outputs(6858);
    layer2_outputs(5899) <= (layer1_outputs(338)) xor (layer1_outputs(3930));
    layer2_outputs(5900) <= not(layer1_outputs(7680));
    layer2_outputs(5901) <= layer1_outputs(4140);
    layer2_outputs(5902) <= not(layer1_outputs(1856));
    layer2_outputs(5903) <= layer1_outputs(11233);
    layer2_outputs(5904) <= layer1_outputs(11027);
    layer2_outputs(5905) <= not(layer1_outputs(5231));
    layer2_outputs(5906) <= '1';
    layer2_outputs(5907) <= layer1_outputs(11478);
    layer2_outputs(5908) <= not(layer1_outputs(4251));
    layer2_outputs(5909) <= not((layer1_outputs(1386)) xor (layer1_outputs(5387)));
    layer2_outputs(5910) <= not(layer1_outputs(987)) or (layer1_outputs(5152));
    layer2_outputs(5911) <= layer1_outputs(8496);
    layer2_outputs(5912) <= layer1_outputs(6806);
    layer2_outputs(5913) <= not(layer1_outputs(4469));
    layer2_outputs(5914) <= not(layer1_outputs(9484));
    layer2_outputs(5915) <= (layer1_outputs(4859)) and (layer1_outputs(11086));
    layer2_outputs(5916) <= not(layer1_outputs(1322)) or (layer1_outputs(7613));
    layer2_outputs(5917) <= not((layer1_outputs(522)) and (layer1_outputs(2033)));
    layer2_outputs(5918) <= layer1_outputs(9497);
    layer2_outputs(5919) <= layer1_outputs(11214);
    layer2_outputs(5920) <= (layer1_outputs(7147)) or (layer1_outputs(9297));
    layer2_outputs(5921) <= not(layer1_outputs(9051));
    layer2_outputs(5922) <= not(layer1_outputs(7069));
    layer2_outputs(5923) <= (layer1_outputs(10273)) xor (layer1_outputs(12438));
    layer2_outputs(5924) <= (layer1_outputs(952)) xor (layer1_outputs(7875));
    layer2_outputs(5925) <= layer1_outputs(11807);
    layer2_outputs(5926) <= not(layer1_outputs(1438));
    layer2_outputs(5927) <= layer1_outputs(6195);
    layer2_outputs(5928) <= not(layer1_outputs(228));
    layer2_outputs(5929) <= not((layer1_outputs(8862)) xor (layer1_outputs(2220)));
    layer2_outputs(5930) <= layer1_outputs(11816);
    layer2_outputs(5931) <= not((layer1_outputs(7421)) xor (layer1_outputs(2711)));
    layer2_outputs(5932) <= layer1_outputs(2789);
    layer2_outputs(5933) <= not((layer1_outputs(4045)) xor (layer1_outputs(10147)));
    layer2_outputs(5934) <= layer1_outputs(485);
    layer2_outputs(5935) <= layer1_outputs(12719);
    layer2_outputs(5936) <= not((layer1_outputs(7671)) xor (layer1_outputs(9821)));
    layer2_outputs(5937) <= not((layer1_outputs(11773)) or (layer1_outputs(120)));
    layer2_outputs(5938) <= (layer1_outputs(11398)) and not (layer1_outputs(8549));
    layer2_outputs(5939) <= layer1_outputs(11882);
    layer2_outputs(5940) <= not(layer1_outputs(11827)) or (layer1_outputs(2088));
    layer2_outputs(5941) <= not(layer1_outputs(11317));
    layer2_outputs(5942) <= (layer1_outputs(6166)) xor (layer1_outputs(3626));
    layer2_outputs(5943) <= layer1_outputs(6659);
    layer2_outputs(5944) <= not(layer1_outputs(4312));
    layer2_outputs(5945) <= layer1_outputs(885);
    layer2_outputs(5946) <= layer1_outputs(825);
    layer2_outputs(5947) <= not((layer1_outputs(12729)) xor (layer1_outputs(1636)));
    layer2_outputs(5948) <= not((layer1_outputs(695)) or (layer1_outputs(8488)));
    layer2_outputs(5949) <= layer1_outputs(3686);
    layer2_outputs(5950) <= not((layer1_outputs(1534)) or (layer1_outputs(11584)));
    layer2_outputs(5951) <= layer1_outputs(3342);
    layer2_outputs(5952) <= (layer1_outputs(11895)) and (layer1_outputs(9666));
    layer2_outputs(5953) <= not(layer1_outputs(12239));
    layer2_outputs(5954) <= (layer1_outputs(427)) and not (layer1_outputs(7318));
    layer2_outputs(5955) <= not(layer1_outputs(3341));
    layer2_outputs(5956) <= not(layer1_outputs(3683)) or (layer1_outputs(12731));
    layer2_outputs(5957) <= not(layer1_outputs(9238)) or (layer1_outputs(3140));
    layer2_outputs(5958) <= layer1_outputs(38);
    layer2_outputs(5959) <= layer1_outputs(2604);
    layer2_outputs(5960) <= not(layer1_outputs(8292));
    layer2_outputs(5961) <= not(layer1_outputs(12405));
    layer2_outputs(5962) <= not(layer1_outputs(3301)) or (layer1_outputs(4133));
    layer2_outputs(5963) <= not(layer1_outputs(9100));
    layer2_outputs(5964) <= not(layer1_outputs(6172)) or (layer1_outputs(8152));
    layer2_outputs(5965) <= not((layer1_outputs(3141)) xor (layer1_outputs(628)));
    layer2_outputs(5966) <= not(layer1_outputs(12023)) or (layer1_outputs(8217));
    layer2_outputs(5967) <= layer1_outputs(7769);
    layer2_outputs(5968) <= (layer1_outputs(7156)) and not (layer1_outputs(10806));
    layer2_outputs(5969) <= (layer1_outputs(11669)) and (layer1_outputs(2990));
    layer2_outputs(5970) <= not(layer1_outputs(11696));
    layer2_outputs(5971) <= layer1_outputs(2190);
    layer2_outputs(5972) <= not(layer1_outputs(1505));
    layer2_outputs(5973) <= layer1_outputs(1770);
    layer2_outputs(5974) <= layer1_outputs(9754);
    layer2_outputs(5975) <= (layer1_outputs(6105)) and (layer1_outputs(12673));
    layer2_outputs(5976) <= not(layer1_outputs(8974));
    layer2_outputs(5977) <= not(layer1_outputs(3824));
    layer2_outputs(5978) <= not(layer1_outputs(9798));
    layer2_outputs(5979) <= not(layer1_outputs(11713)) or (layer1_outputs(11895));
    layer2_outputs(5980) <= not((layer1_outputs(3525)) and (layer1_outputs(10810)));
    layer2_outputs(5981) <= (layer1_outputs(3765)) and not (layer1_outputs(5221));
    layer2_outputs(5982) <= not(layer1_outputs(799));
    layer2_outputs(5983) <= not((layer1_outputs(11169)) or (layer1_outputs(607)));
    layer2_outputs(5984) <= not(layer1_outputs(9091));
    layer2_outputs(5985) <= (layer1_outputs(2881)) and (layer1_outputs(2736));
    layer2_outputs(5986) <= (layer1_outputs(2362)) and not (layer1_outputs(7071));
    layer2_outputs(5987) <= layer1_outputs(4221);
    layer2_outputs(5988) <= not(layer1_outputs(6679));
    layer2_outputs(5989) <= not((layer1_outputs(11779)) xor (layer1_outputs(10602)));
    layer2_outputs(5990) <= not(layer1_outputs(4684));
    layer2_outputs(5991) <= not(layer1_outputs(11968));
    layer2_outputs(5992) <= not(layer1_outputs(9411));
    layer2_outputs(5993) <= (layer1_outputs(3887)) and (layer1_outputs(5587));
    layer2_outputs(5994) <= (layer1_outputs(7518)) and (layer1_outputs(12521));
    layer2_outputs(5995) <= not(layer1_outputs(11653)) or (layer1_outputs(11580));
    layer2_outputs(5996) <= not(layer1_outputs(7213));
    layer2_outputs(5997) <= not((layer1_outputs(3242)) or (layer1_outputs(24)));
    layer2_outputs(5998) <= not(layer1_outputs(11659));
    layer2_outputs(5999) <= not(layer1_outputs(7599));
    layer2_outputs(6000) <= layer1_outputs(10552);
    layer2_outputs(6001) <= not(layer1_outputs(8510)) or (layer1_outputs(1268));
    layer2_outputs(6002) <= (layer1_outputs(12601)) xor (layer1_outputs(10562));
    layer2_outputs(6003) <= not(layer1_outputs(4428));
    layer2_outputs(6004) <= (layer1_outputs(2470)) and not (layer1_outputs(6751));
    layer2_outputs(6005) <= layer1_outputs(6374);
    layer2_outputs(6006) <= not(layer1_outputs(9357));
    layer2_outputs(6007) <= layer1_outputs(8628);
    layer2_outputs(6008) <= layer1_outputs(7647);
    layer2_outputs(6009) <= (layer1_outputs(12717)) and (layer1_outputs(7264));
    layer2_outputs(6010) <= layer1_outputs(5772);
    layer2_outputs(6011) <= layer1_outputs(10456);
    layer2_outputs(6012) <= layer1_outputs(7442);
    layer2_outputs(6013) <= not(layer1_outputs(7817));
    layer2_outputs(6014) <= not(layer1_outputs(8079));
    layer2_outputs(6015) <= not(layer1_outputs(2685));
    layer2_outputs(6016) <= (layer1_outputs(10381)) and not (layer1_outputs(6007));
    layer2_outputs(6017) <= not(layer1_outputs(527)) or (layer1_outputs(3290));
    layer2_outputs(6018) <= not(layer1_outputs(725)) or (layer1_outputs(6617));
    layer2_outputs(6019) <= not(layer1_outputs(8883));
    layer2_outputs(6020) <= not(layer1_outputs(10887));
    layer2_outputs(6021) <= not((layer1_outputs(4167)) or (layer1_outputs(11104)));
    layer2_outputs(6022) <= not(layer1_outputs(10317));
    layer2_outputs(6023) <= (layer1_outputs(1355)) xor (layer1_outputs(1341));
    layer2_outputs(6024) <= not((layer1_outputs(2238)) or (layer1_outputs(6729)));
    layer2_outputs(6025) <= not(layer1_outputs(1157));
    layer2_outputs(6026) <= not((layer1_outputs(6228)) and (layer1_outputs(8080)));
    layer2_outputs(6027) <= layer1_outputs(2682);
    layer2_outputs(6028) <= not((layer1_outputs(3213)) xor (layer1_outputs(5740)));
    layer2_outputs(6029) <= not(layer1_outputs(5720));
    layer2_outputs(6030) <= (layer1_outputs(6989)) and (layer1_outputs(11427));
    layer2_outputs(6031) <= not(layer1_outputs(10719)) or (layer1_outputs(8146));
    layer2_outputs(6032) <= layer1_outputs(9374);
    layer2_outputs(6033) <= layer1_outputs(11405);
    layer2_outputs(6034) <= not(layer1_outputs(8900));
    layer2_outputs(6035) <= (layer1_outputs(10186)) and not (layer1_outputs(8106));
    layer2_outputs(6036) <= (layer1_outputs(11295)) xor (layer1_outputs(9557));
    layer2_outputs(6037) <= layer1_outputs(3458);
    layer2_outputs(6038) <= not(layer1_outputs(12564));
    layer2_outputs(6039) <= not(layer1_outputs(12145)) or (layer1_outputs(9917));
    layer2_outputs(6040) <= layer1_outputs(3954);
    layer2_outputs(6041) <= (layer1_outputs(11727)) and not (layer1_outputs(310));
    layer2_outputs(6042) <= layer1_outputs(12536);
    layer2_outputs(6043) <= not(layer1_outputs(4973));
    layer2_outputs(6044) <= layer1_outputs(2057);
    layer2_outputs(6045) <= (layer1_outputs(5655)) and not (layer1_outputs(5906));
    layer2_outputs(6046) <= not(layer1_outputs(8940));
    layer2_outputs(6047) <= not(layer1_outputs(11414)) or (layer1_outputs(2019));
    layer2_outputs(6048) <= not(layer1_outputs(1139)) or (layer1_outputs(6812));
    layer2_outputs(6049) <= layer1_outputs(10913);
    layer2_outputs(6050) <= (layer1_outputs(9915)) and not (layer1_outputs(1168));
    layer2_outputs(6051) <= (layer1_outputs(810)) and (layer1_outputs(4636));
    layer2_outputs(6052) <= not(layer1_outputs(9520));
    layer2_outputs(6053) <= not(layer1_outputs(1970)) or (layer1_outputs(12168));
    layer2_outputs(6054) <= not((layer1_outputs(3759)) and (layer1_outputs(10361)));
    layer2_outputs(6055) <= not((layer1_outputs(3585)) and (layer1_outputs(187)));
    layer2_outputs(6056) <= not(layer1_outputs(8509));
    layer2_outputs(6057) <= not(layer1_outputs(3309));
    layer2_outputs(6058) <= layer1_outputs(10543);
    layer2_outputs(6059) <= not(layer1_outputs(11205));
    layer2_outputs(6060) <= layer1_outputs(6842);
    layer2_outputs(6061) <= not((layer1_outputs(7505)) xor (layer1_outputs(9110)));
    layer2_outputs(6062) <= '1';
    layer2_outputs(6063) <= not(layer1_outputs(9743));
    layer2_outputs(6064) <= layer1_outputs(9896);
    layer2_outputs(6065) <= (layer1_outputs(6123)) and (layer1_outputs(3099));
    layer2_outputs(6066) <= not(layer1_outputs(9316));
    layer2_outputs(6067) <= (layer1_outputs(10402)) and not (layer1_outputs(728));
    layer2_outputs(6068) <= layer1_outputs(9744);
    layer2_outputs(6069) <= not(layer1_outputs(275)) or (layer1_outputs(11813));
    layer2_outputs(6070) <= not(layer1_outputs(1387));
    layer2_outputs(6071) <= not(layer1_outputs(6279)) or (layer1_outputs(1276));
    layer2_outputs(6072) <= (layer1_outputs(2439)) and (layer1_outputs(775));
    layer2_outputs(6073) <= not(layer1_outputs(4258)) or (layer1_outputs(5939));
    layer2_outputs(6074) <= not(layer1_outputs(119));
    layer2_outputs(6075) <= (layer1_outputs(8592)) and not (layer1_outputs(11728));
    layer2_outputs(6076) <= (layer1_outputs(5396)) xor (layer1_outputs(9871));
    layer2_outputs(6077) <= (layer1_outputs(1773)) xor (layer1_outputs(3414));
    layer2_outputs(6078) <= (layer1_outputs(7250)) and not (layer1_outputs(2319));
    layer2_outputs(6079) <= not(layer1_outputs(8390)) or (layer1_outputs(8906));
    layer2_outputs(6080) <= layer1_outputs(3254);
    layer2_outputs(6081) <= layer1_outputs(3341);
    layer2_outputs(6082) <= (layer1_outputs(8651)) and not (layer1_outputs(11892));
    layer2_outputs(6083) <= not(layer1_outputs(10618)) or (layer1_outputs(11495));
    layer2_outputs(6084) <= not((layer1_outputs(11924)) or (layer1_outputs(9987)));
    layer2_outputs(6085) <= layer1_outputs(5469);
    layer2_outputs(6086) <= layer1_outputs(8560);
    layer2_outputs(6087) <= not((layer1_outputs(1187)) xor (layer1_outputs(12488)));
    layer2_outputs(6088) <= (layer1_outputs(2602)) and not (layer1_outputs(4414));
    layer2_outputs(6089) <= not((layer1_outputs(7418)) xor (layer1_outputs(8163)));
    layer2_outputs(6090) <= (layer1_outputs(8763)) or (layer1_outputs(7413));
    layer2_outputs(6091) <= layer1_outputs(8481);
    layer2_outputs(6092) <= layer1_outputs(6061);
    layer2_outputs(6093) <= not(layer1_outputs(8108)) or (layer1_outputs(12524));
    layer2_outputs(6094) <= (layer1_outputs(9818)) xor (layer1_outputs(8317));
    layer2_outputs(6095) <= not((layer1_outputs(1453)) or (layer1_outputs(7317)));
    layer2_outputs(6096) <= (layer1_outputs(9703)) and not (layer1_outputs(1963));
    layer2_outputs(6097) <= not((layer1_outputs(8561)) and (layer1_outputs(4762)));
    layer2_outputs(6098) <= layer1_outputs(5462);
    layer2_outputs(6099) <= layer1_outputs(7033);
    layer2_outputs(6100) <= not(layer1_outputs(3510));
    layer2_outputs(6101) <= layer1_outputs(8909);
    layer2_outputs(6102) <= layer1_outputs(2777);
    layer2_outputs(6103) <= layer1_outputs(87);
    layer2_outputs(6104) <= not((layer1_outputs(10186)) xor (layer1_outputs(2158)));
    layer2_outputs(6105) <= (layer1_outputs(7963)) and not (layer1_outputs(12486));
    layer2_outputs(6106) <= (layer1_outputs(2217)) and (layer1_outputs(425));
    layer2_outputs(6107) <= layer1_outputs(12325);
    layer2_outputs(6108) <= layer1_outputs(9980);
    layer2_outputs(6109) <= (layer1_outputs(11186)) xor (layer1_outputs(3980));
    layer2_outputs(6110) <= not((layer1_outputs(5937)) and (layer1_outputs(11329)));
    layer2_outputs(6111) <= not((layer1_outputs(1327)) xor (layer1_outputs(8922)));
    layer2_outputs(6112) <= not((layer1_outputs(6124)) or (layer1_outputs(5785)));
    layer2_outputs(6113) <= not((layer1_outputs(8332)) and (layer1_outputs(8264)));
    layer2_outputs(6114) <= (layer1_outputs(9940)) xor (layer1_outputs(2550));
    layer2_outputs(6115) <= not((layer1_outputs(9887)) and (layer1_outputs(6897)));
    layer2_outputs(6116) <= layer1_outputs(5650);
    layer2_outputs(6117) <= (layer1_outputs(10184)) and not (layer1_outputs(7764));
    layer2_outputs(6118) <= (layer1_outputs(4202)) and not (layer1_outputs(10990));
    layer2_outputs(6119) <= not(layer1_outputs(1474));
    layer2_outputs(6120) <= not(layer1_outputs(10323));
    layer2_outputs(6121) <= not((layer1_outputs(4854)) and (layer1_outputs(3381)));
    layer2_outputs(6122) <= (layer1_outputs(8954)) xor (layer1_outputs(6343));
    layer2_outputs(6123) <= not(layer1_outputs(12662));
    layer2_outputs(6124) <= (layer1_outputs(10197)) and not (layer1_outputs(3176));
    layer2_outputs(6125) <= not(layer1_outputs(5663)) or (layer1_outputs(9321));
    layer2_outputs(6126) <= (layer1_outputs(6605)) and not (layer1_outputs(9443));
    layer2_outputs(6127) <= layer1_outputs(3133);
    layer2_outputs(6128) <= not((layer1_outputs(938)) and (layer1_outputs(12354)));
    layer2_outputs(6129) <= not(layer1_outputs(2679));
    layer2_outputs(6130) <= layer1_outputs(1603);
    layer2_outputs(6131) <= layer1_outputs(10924);
    layer2_outputs(6132) <= not(layer1_outputs(4888));
    layer2_outputs(6133) <= layer1_outputs(12760);
    layer2_outputs(6134) <= not(layer1_outputs(5163)) or (layer1_outputs(2020));
    layer2_outputs(6135) <= not(layer1_outputs(12720));
    layer2_outputs(6136) <= not((layer1_outputs(134)) or (layer1_outputs(9948)));
    layer2_outputs(6137) <= layer1_outputs(2554);
    layer2_outputs(6138) <= not(layer1_outputs(3513)) or (layer1_outputs(5189));
    layer2_outputs(6139) <= (layer1_outputs(1259)) and not (layer1_outputs(9460));
    layer2_outputs(6140) <= layer1_outputs(9003);
    layer2_outputs(6141) <= not(layer1_outputs(9255)) or (layer1_outputs(4764));
    layer2_outputs(6142) <= not(layer1_outputs(4237));
    layer2_outputs(6143) <= not(layer1_outputs(8852)) or (layer1_outputs(4727));
    layer2_outputs(6144) <= layer1_outputs(880);
    layer2_outputs(6145) <= not(layer1_outputs(4462));
    layer2_outputs(6146) <= not((layer1_outputs(8122)) xor (layer1_outputs(8236)));
    layer2_outputs(6147) <= layer1_outputs(5056);
    layer2_outputs(6148) <= (layer1_outputs(194)) xor (layer1_outputs(4095));
    layer2_outputs(6149) <= (layer1_outputs(691)) and (layer1_outputs(12752));
    layer2_outputs(6150) <= (layer1_outputs(1149)) or (layer1_outputs(12459));
    layer2_outputs(6151) <= not(layer1_outputs(8302));
    layer2_outputs(6152) <= layer1_outputs(3629);
    layer2_outputs(6153) <= layer1_outputs(4937);
    layer2_outputs(6154) <= not(layer1_outputs(7886));
    layer2_outputs(6155) <= layer1_outputs(7988);
    layer2_outputs(6156) <= not((layer1_outputs(2951)) and (layer1_outputs(7832)));
    layer2_outputs(6157) <= not((layer1_outputs(8358)) and (layer1_outputs(6062)));
    layer2_outputs(6158) <= layer1_outputs(5083);
    layer2_outputs(6159) <= not(layer1_outputs(6515)) or (layer1_outputs(8337));
    layer2_outputs(6160) <= not((layer1_outputs(9016)) or (layer1_outputs(2253)));
    layer2_outputs(6161) <= layer1_outputs(6604);
    layer2_outputs(6162) <= not(layer1_outputs(8960));
    layer2_outputs(6163) <= not(layer1_outputs(9226));
    layer2_outputs(6164) <= not(layer1_outputs(10457));
    layer2_outputs(6165) <= not(layer1_outputs(1680)) or (layer1_outputs(9295));
    layer2_outputs(6166) <= not(layer1_outputs(3618));
    layer2_outputs(6167) <= not(layer1_outputs(10817));
    layer2_outputs(6168) <= not(layer1_outputs(5381));
    layer2_outputs(6169) <= not(layer1_outputs(5941));
    layer2_outputs(6170) <= layer1_outputs(3421);
    layer2_outputs(6171) <= layer1_outputs(11364);
    layer2_outputs(6172) <= (layer1_outputs(9754)) xor (layer1_outputs(1154));
    layer2_outputs(6173) <= not(layer1_outputs(3468));
    layer2_outputs(6174) <= layer1_outputs(1467);
    layer2_outputs(6175) <= layer1_outputs(7547);
    layer2_outputs(6176) <= '1';
    layer2_outputs(6177) <= (layer1_outputs(5122)) or (layer1_outputs(10630));
    layer2_outputs(6178) <= not(layer1_outputs(3283));
    layer2_outputs(6179) <= layer1_outputs(10311);
    layer2_outputs(6180) <= (layer1_outputs(5306)) and not (layer1_outputs(6134));
    layer2_outputs(6181) <= '1';
    layer2_outputs(6182) <= layer1_outputs(2051);
    layer2_outputs(6183) <= not((layer1_outputs(844)) or (layer1_outputs(12629)));
    layer2_outputs(6184) <= '1';
    layer2_outputs(6185) <= (layer1_outputs(1511)) or (layer1_outputs(8503));
    layer2_outputs(6186) <= (layer1_outputs(5130)) or (layer1_outputs(2262));
    layer2_outputs(6187) <= not(layer1_outputs(9181));
    layer2_outputs(6188) <= not(layer1_outputs(11782)) or (layer1_outputs(4900));
    layer2_outputs(6189) <= (layer1_outputs(2035)) xor (layer1_outputs(12725));
    layer2_outputs(6190) <= not(layer1_outputs(4354));
    layer2_outputs(6191) <= not(layer1_outputs(8110));
    layer2_outputs(6192) <= (layer1_outputs(10651)) xor (layer1_outputs(12698));
    layer2_outputs(6193) <= not(layer1_outputs(10744));
    layer2_outputs(6194) <= not(layer1_outputs(8817));
    layer2_outputs(6195) <= layer1_outputs(7559);
    layer2_outputs(6196) <= layer1_outputs(1829);
    layer2_outputs(6197) <= (layer1_outputs(11246)) and not (layer1_outputs(7447));
    layer2_outputs(6198) <= not((layer1_outputs(11535)) and (layer1_outputs(10784)));
    layer2_outputs(6199) <= (layer1_outputs(2519)) xor (layer1_outputs(52));
    layer2_outputs(6200) <= not(layer1_outputs(8485)) or (layer1_outputs(8353));
    layer2_outputs(6201) <= not((layer1_outputs(1774)) and (layer1_outputs(9841)));
    layer2_outputs(6202) <= '0';
    layer2_outputs(6203) <= not((layer1_outputs(12682)) and (layer1_outputs(7970)));
    layer2_outputs(6204) <= not(layer1_outputs(9043));
    layer2_outputs(6205) <= not(layer1_outputs(237)) or (layer1_outputs(4248));
    layer2_outputs(6206) <= layer1_outputs(11893);
    layer2_outputs(6207) <= (layer1_outputs(2005)) and not (layer1_outputs(1038));
    layer2_outputs(6208) <= not(layer1_outputs(3611)) or (layer1_outputs(11450));
    layer2_outputs(6209) <= not(layer1_outputs(9743));
    layer2_outputs(6210) <= not(layer1_outputs(11670));
    layer2_outputs(6211) <= not(layer1_outputs(8804));
    layer2_outputs(6212) <= not((layer1_outputs(338)) xor (layer1_outputs(7712)));
    layer2_outputs(6213) <= (layer1_outputs(7469)) and not (layer1_outputs(681));
    layer2_outputs(6214) <= layer1_outputs(10156);
    layer2_outputs(6215) <= not(layer1_outputs(614));
    layer2_outputs(6216) <= not(layer1_outputs(2115));
    layer2_outputs(6217) <= (layer1_outputs(2435)) and (layer1_outputs(8565));
    layer2_outputs(6218) <= not(layer1_outputs(1071));
    layer2_outputs(6219) <= not(layer1_outputs(2315)) or (layer1_outputs(10288));
    layer2_outputs(6220) <= not(layer1_outputs(4787));
    layer2_outputs(6221) <= (layer1_outputs(9521)) xor (layer1_outputs(9116));
    layer2_outputs(6222) <= not(layer1_outputs(11369));
    layer2_outputs(6223) <= not(layer1_outputs(5600));
    layer2_outputs(6224) <= not(layer1_outputs(6207));
    layer2_outputs(6225) <= (layer1_outputs(4115)) and not (layer1_outputs(5062));
    layer2_outputs(6226) <= not((layer1_outputs(11588)) xor (layer1_outputs(665)));
    layer2_outputs(6227) <= (layer1_outputs(6891)) xor (layer1_outputs(12572));
    layer2_outputs(6228) <= (layer1_outputs(9050)) or (layer1_outputs(8881));
    layer2_outputs(6229) <= (layer1_outputs(4817)) xor (layer1_outputs(12378));
    layer2_outputs(6230) <= not((layer1_outputs(7844)) and (layer1_outputs(7434)));
    layer2_outputs(6231) <= layer1_outputs(8319);
    layer2_outputs(6232) <= not((layer1_outputs(2285)) xor (layer1_outputs(4324)));
    layer2_outputs(6233) <= not(layer1_outputs(7858));
    layer2_outputs(6234) <= (layer1_outputs(1884)) xor (layer1_outputs(8208));
    layer2_outputs(6235) <= not(layer1_outputs(3832)) or (layer1_outputs(4676));
    layer2_outputs(6236) <= layer1_outputs(6250);
    layer2_outputs(6237) <= (layer1_outputs(12210)) and not (layer1_outputs(11213));
    layer2_outputs(6238) <= not(layer1_outputs(2335)) or (layer1_outputs(7229));
    layer2_outputs(6239) <= (layer1_outputs(5115)) and (layer1_outputs(12003));
    layer2_outputs(6240) <= layer1_outputs(2314);
    layer2_outputs(6241) <= layer1_outputs(432);
    layer2_outputs(6242) <= (layer1_outputs(10481)) or (layer1_outputs(3088));
    layer2_outputs(6243) <= layer1_outputs(8976);
    layer2_outputs(6244) <= layer1_outputs(712);
    layer2_outputs(6245) <= not(layer1_outputs(3825)) or (layer1_outputs(7830));
    layer2_outputs(6246) <= not(layer1_outputs(12559));
    layer2_outputs(6247) <= layer1_outputs(709);
    layer2_outputs(6248) <= not(layer1_outputs(8322));
    layer2_outputs(6249) <= not(layer1_outputs(429));
    layer2_outputs(6250) <= not(layer1_outputs(5870)) or (layer1_outputs(11829));
    layer2_outputs(6251) <= (layer1_outputs(2034)) or (layer1_outputs(11303));
    layer2_outputs(6252) <= layer1_outputs(10700);
    layer2_outputs(6253) <= not(layer1_outputs(8035));
    layer2_outputs(6254) <= not(layer1_outputs(2466));
    layer2_outputs(6255) <= layer1_outputs(12359);
    layer2_outputs(6256) <= (layer1_outputs(2858)) and not (layer1_outputs(8491));
    layer2_outputs(6257) <= layer1_outputs(4603);
    layer2_outputs(6258) <= layer1_outputs(1381);
    layer2_outputs(6259) <= not(layer1_outputs(12661));
    layer2_outputs(6260) <= (layer1_outputs(1088)) xor (layer1_outputs(9968));
    layer2_outputs(6261) <= not(layer1_outputs(8472));
    layer2_outputs(6262) <= (layer1_outputs(5285)) or (layer1_outputs(1728));
    layer2_outputs(6263) <= not(layer1_outputs(2870)) or (layer1_outputs(9550));
    layer2_outputs(6264) <= layer1_outputs(4208);
    layer2_outputs(6265) <= not(layer1_outputs(5815));
    layer2_outputs(6266) <= (layer1_outputs(9010)) and not (layer1_outputs(9201));
    layer2_outputs(6267) <= (layer1_outputs(11916)) and not (layer1_outputs(6644));
    layer2_outputs(6268) <= (layer1_outputs(9729)) or (layer1_outputs(7198));
    layer2_outputs(6269) <= not(layer1_outputs(4839));
    layer2_outputs(6270) <= not(layer1_outputs(7488));
    layer2_outputs(6271) <= layer1_outputs(81);
    layer2_outputs(6272) <= layer1_outputs(12136);
    layer2_outputs(6273) <= not((layer1_outputs(10756)) and (layer1_outputs(963)));
    layer2_outputs(6274) <= (layer1_outputs(3061)) xor (layer1_outputs(8739));
    layer2_outputs(6275) <= (layer1_outputs(9206)) or (layer1_outputs(1903));
    layer2_outputs(6276) <= not(layer1_outputs(9911));
    layer2_outputs(6277) <= not((layer1_outputs(7132)) xor (layer1_outputs(126)));
    layer2_outputs(6278) <= not(layer1_outputs(7816));
    layer2_outputs(6279) <= not(layer1_outputs(12611));
    layer2_outputs(6280) <= not(layer1_outputs(8598));
    layer2_outputs(6281) <= not(layer1_outputs(6133));
    layer2_outputs(6282) <= layer1_outputs(4644);
    layer2_outputs(6283) <= not(layer1_outputs(3513));
    layer2_outputs(6284) <= layer1_outputs(536);
    layer2_outputs(6285) <= not((layer1_outputs(3795)) or (layer1_outputs(439)));
    layer2_outputs(6286) <= layer1_outputs(3394);
    layer2_outputs(6287) <= layer1_outputs(4566);
    layer2_outputs(6288) <= layer1_outputs(4932);
    layer2_outputs(6289) <= (layer1_outputs(2280)) and not (layer1_outputs(7990));
    layer2_outputs(6290) <= (layer1_outputs(416)) and (layer1_outputs(11858));
    layer2_outputs(6291) <= not(layer1_outputs(2179));
    layer2_outputs(6292) <= '1';
    layer2_outputs(6293) <= not(layer1_outputs(1736));
    layer2_outputs(6294) <= not(layer1_outputs(3463));
    layer2_outputs(6295) <= (layer1_outputs(11038)) and not (layer1_outputs(744));
    layer2_outputs(6296) <= (layer1_outputs(1450)) and (layer1_outputs(5147));
    layer2_outputs(6297) <= layer1_outputs(8867);
    layer2_outputs(6298) <= not(layer1_outputs(9390));
    layer2_outputs(6299) <= not((layer1_outputs(2317)) xor (layer1_outputs(10747)));
    layer2_outputs(6300) <= not((layer1_outputs(3346)) xor (layer1_outputs(5181)));
    layer2_outputs(6301) <= layer1_outputs(317);
    layer2_outputs(6302) <= (layer1_outputs(10258)) xor (layer1_outputs(12494));
    layer2_outputs(6303) <= not(layer1_outputs(8013));
    layer2_outputs(6304) <= not(layer1_outputs(9065));
    layer2_outputs(6305) <= not((layer1_outputs(11943)) xor (layer1_outputs(10493)));
    layer2_outputs(6306) <= not(layer1_outputs(11109));
    layer2_outputs(6307) <= not(layer1_outputs(1750));
    layer2_outputs(6308) <= not((layer1_outputs(3046)) or (layer1_outputs(6976)));
    layer2_outputs(6309) <= not(layer1_outputs(6581));
    layer2_outputs(6310) <= not(layer1_outputs(10118));
    layer2_outputs(6311) <= not(layer1_outputs(5572));
    layer2_outputs(6312) <= not(layer1_outputs(9301));
    layer2_outputs(6313) <= not((layer1_outputs(8706)) or (layer1_outputs(9010)));
    layer2_outputs(6314) <= (layer1_outputs(5484)) and not (layer1_outputs(3081));
    layer2_outputs(6315) <= layer1_outputs(6169);
    layer2_outputs(6316) <= not(layer1_outputs(1916));
    layer2_outputs(6317) <= (layer1_outputs(1755)) or (layer1_outputs(12421));
    layer2_outputs(6318) <= not((layer1_outputs(4935)) and (layer1_outputs(869)));
    layer2_outputs(6319) <= layer1_outputs(8611);
    layer2_outputs(6320) <= not((layer1_outputs(2974)) or (layer1_outputs(10770)));
    layer2_outputs(6321) <= layer1_outputs(10358);
    layer2_outputs(6322) <= layer1_outputs(414);
    layer2_outputs(6323) <= not((layer1_outputs(1799)) and (layer1_outputs(501)));
    layer2_outputs(6324) <= layer1_outputs(8285);
    layer2_outputs(6325) <= not(layer1_outputs(1360));
    layer2_outputs(6326) <= not(layer1_outputs(7188));
    layer2_outputs(6327) <= not(layer1_outputs(9021));
    layer2_outputs(6328) <= (layer1_outputs(5701)) and (layer1_outputs(4304));
    layer2_outputs(6329) <= not(layer1_outputs(8522));
    layer2_outputs(6330) <= not(layer1_outputs(5218));
    layer2_outputs(6331) <= layer1_outputs(6610);
    layer2_outputs(6332) <= not((layer1_outputs(8935)) and (layer1_outputs(8252)));
    layer2_outputs(6333) <= (layer1_outputs(1697)) and not (layer1_outputs(6152));
    layer2_outputs(6334) <= layer1_outputs(8289);
    layer2_outputs(6335) <= not((layer1_outputs(2261)) xor (layer1_outputs(3958)));
    layer2_outputs(6336) <= not(layer1_outputs(160)) or (layer1_outputs(5989));
    layer2_outputs(6337) <= layer1_outputs(10695);
    layer2_outputs(6338) <= not(layer1_outputs(4296));
    layer2_outputs(6339) <= layer1_outputs(6851);
    layer2_outputs(6340) <= layer1_outputs(10233);
    layer2_outputs(6341) <= not(layer1_outputs(9463));
    layer2_outputs(6342) <= not((layer1_outputs(8184)) or (layer1_outputs(7210)));
    layer2_outputs(6343) <= (layer1_outputs(3783)) xor (layer1_outputs(12272));
    layer2_outputs(6344) <= (layer1_outputs(10871)) and not (layer1_outputs(12560));
    layer2_outputs(6345) <= (layer1_outputs(3197)) and (layer1_outputs(877));
    layer2_outputs(6346) <= not(layer1_outputs(3530));
    layer2_outputs(6347) <= (layer1_outputs(4552)) xor (layer1_outputs(11733));
    layer2_outputs(6348) <= (layer1_outputs(7874)) and (layer1_outputs(10596));
    layer2_outputs(6349) <= not(layer1_outputs(10870)) or (layer1_outputs(2722));
    layer2_outputs(6350) <= not(layer1_outputs(9020));
    layer2_outputs(6351) <= not((layer1_outputs(9828)) xor (layer1_outputs(1608)));
    layer2_outputs(6352) <= not(layer1_outputs(2177)) or (layer1_outputs(2344));
    layer2_outputs(6353) <= not((layer1_outputs(205)) xor (layer1_outputs(6549)));
    layer2_outputs(6354) <= layer1_outputs(359);
    layer2_outputs(6355) <= layer1_outputs(5110);
    layer2_outputs(6356) <= (layer1_outputs(11215)) xor (layer1_outputs(2615));
    layer2_outputs(6357) <= layer1_outputs(76);
    layer2_outputs(6358) <= not((layer1_outputs(4340)) and (layer1_outputs(8314)));
    layer2_outputs(6359) <= not((layer1_outputs(5657)) and (layer1_outputs(7546)));
    layer2_outputs(6360) <= (layer1_outputs(6733)) or (layer1_outputs(11175));
    layer2_outputs(6361) <= (layer1_outputs(6882)) and not (layer1_outputs(7405));
    layer2_outputs(6362) <= (layer1_outputs(8557)) or (layer1_outputs(11674));
    layer2_outputs(6363) <= (layer1_outputs(5724)) xor (layer1_outputs(2928));
    layer2_outputs(6364) <= not(layer1_outputs(12776)) or (layer1_outputs(11498));
    layer2_outputs(6365) <= not(layer1_outputs(6159));
    layer2_outputs(6366) <= not((layer1_outputs(9829)) xor (layer1_outputs(4825)));
    layer2_outputs(6367) <= layer1_outputs(820);
    layer2_outputs(6368) <= (layer1_outputs(854)) and (layer1_outputs(11497));
    layer2_outputs(6369) <= layer1_outputs(6108);
    layer2_outputs(6370) <= (layer1_outputs(7528)) or (layer1_outputs(12002));
    layer2_outputs(6371) <= not(layer1_outputs(10587));
    layer2_outputs(6372) <= not(layer1_outputs(1257));
    layer2_outputs(6373) <= not(layer1_outputs(5171));
    layer2_outputs(6374) <= not(layer1_outputs(1163));
    layer2_outputs(6375) <= not(layer1_outputs(12309));
    layer2_outputs(6376) <= not(layer1_outputs(4210));
    layer2_outputs(6377) <= layer1_outputs(7842);
    layer2_outputs(6378) <= (layer1_outputs(6275)) and not (layer1_outputs(2659));
    layer2_outputs(6379) <= not(layer1_outputs(363)) or (layer1_outputs(11170));
    layer2_outputs(6380) <= not((layer1_outputs(2753)) xor (layer1_outputs(9394)));
    layer2_outputs(6381) <= (layer1_outputs(5787)) xor (layer1_outputs(3975));
    layer2_outputs(6382) <= not((layer1_outputs(6193)) xor (layer1_outputs(6004)));
    layer2_outputs(6383) <= not(layer1_outputs(9749));
    layer2_outputs(6384) <= not(layer1_outputs(4125));
    layer2_outputs(6385) <= layer1_outputs(3215);
    layer2_outputs(6386) <= not(layer1_outputs(10271));
    layer2_outputs(6387) <= not(layer1_outputs(6728));
    layer2_outputs(6388) <= (layer1_outputs(965)) and not (layer1_outputs(7513));
    layer2_outputs(6389) <= layer1_outputs(7090);
    layer2_outputs(6390) <= (layer1_outputs(1812)) and not (layer1_outputs(9698));
    layer2_outputs(6391) <= not(layer1_outputs(983)) or (layer1_outputs(12342));
    layer2_outputs(6392) <= not((layer1_outputs(12019)) xor (layer1_outputs(1190)));
    layer2_outputs(6393) <= (layer1_outputs(6435)) and (layer1_outputs(4037));
    layer2_outputs(6394) <= not(layer1_outputs(4511)) or (layer1_outputs(10505));
    layer2_outputs(6395) <= (layer1_outputs(4748)) xor (layer1_outputs(865));
    layer2_outputs(6396) <= layer1_outputs(7891);
    layer2_outputs(6397) <= not(layer1_outputs(5019)) or (layer1_outputs(2237));
    layer2_outputs(6398) <= not(layer1_outputs(11645)) or (layer1_outputs(2090));
    layer2_outputs(6399) <= not(layer1_outputs(4048));
    layer2_outputs(6400) <= not(layer1_outputs(3994)) or (layer1_outputs(2511));
    layer2_outputs(6401) <= (layer1_outputs(9122)) and (layer1_outputs(12395));
    layer2_outputs(6402) <= not(layer1_outputs(5850));
    layer2_outputs(6403) <= not(layer1_outputs(7222)) or (layer1_outputs(8562));
    layer2_outputs(6404) <= not(layer1_outputs(5117));
    layer2_outputs(6405) <= not(layer1_outputs(927));
    layer2_outputs(6406) <= (layer1_outputs(2764)) and not (layer1_outputs(7623));
    layer2_outputs(6407) <= (layer1_outputs(9512)) xor (layer1_outputs(4840));
    layer2_outputs(6408) <= (layer1_outputs(11304)) and (layer1_outputs(2156));
    layer2_outputs(6409) <= layer1_outputs(3299);
    layer2_outputs(6410) <= not(layer1_outputs(2564));
    layer2_outputs(6411) <= (layer1_outputs(6804)) xor (layer1_outputs(11357));
    layer2_outputs(6412) <= layer1_outputs(4502);
    layer2_outputs(6413) <= (layer1_outputs(9502)) or (layer1_outputs(7711));
    layer2_outputs(6414) <= not((layer1_outputs(1852)) or (layer1_outputs(3937)));
    layer2_outputs(6415) <= layer1_outputs(7932);
    layer2_outputs(6416) <= not((layer1_outputs(1943)) or (layer1_outputs(5251)));
    layer2_outputs(6417) <= (layer1_outputs(6960)) xor (layer1_outputs(12518));
    layer2_outputs(6418) <= layer1_outputs(9548);
    layer2_outputs(6419) <= not(layer1_outputs(2309));
    layer2_outputs(6420) <= (layer1_outputs(4977)) or (layer1_outputs(5259));
    layer2_outputs(6421) <= not(layer1_outputs(755));
    layer2_outputs(6422) <= not(layer1_outputs(2351));
    layer2_outputs(6423) <= (layer1_outputs(5266)) and not (layer1_outputs(10773));
    layer2_outputs(6424) <= (layer1_outputs(11840)) xor (layer1_outputs(6515));
    layer2_outputs(6425) <= (layer1_outputs(6500)) or (layer1_outputs(9147));
    layer2_outputs(6426) <= not(layer1_outputs(11199));
    layer2_outputs(6427) <= layer1_outputs(11926);
    layer2_outputs(6428) <= (layer1_outputs(12214)) or (layer1_outputs(8361));
    layer2_outputs(6429) <= layer1_outputs(6075);
    layer2_outputs(6430) <= not(layer1_outputs(1231));
    layer2_outputs(6431) <= not(layer1_outputs(11841));
    layer2_outputs(6432) <= layer1_outputs(2542);
    layer2_outputs(6433) <= not(layer1_outputs(7400));
    layer2_outputs(6434) <= (layer1_outputs(2041)) and (layer1_outputs(2533));
    layer2_outputs(6435) <= not(layer1_outputs(41)) or (layer1_outputs(1974));
    layer2_outputs(6436) <= not(layer1_outputs(10275));
    layer2_outputs(6437) <= layer1_outputs(8490);
    layer2_outputs(6438) <= layer1_outputs(1333);
    layer2_outputs(6439) <= not((layer1_outputs(12068)) xor (layer1_outputs(5895)));
    layer2_outputs(6440) <= not((layer1_outputs(1393)) or (layer1_outputs(5000)));
    layer2_outputs(6441) <= not(layer1_outputs(1717)) or (layer1_outputs(7945));
    layer2_outputs(6442) <= not(layer1_outputs(3075)) or (layer1_outputs(10231));
    layer2_outputs(6443) <= (layer1_outputs(9655)) or (layer1_outputs(12251));
    layer2_outputs(6444) <= not(layer1_outputs(4988));
    layer2_outputs(6445) <= not((layer1_outputs(3444)) and (layer1_outputs(3233)));
    layer2_outputs(6446) <= not(layer1_outputs(6845));
    layer2_outputs(6447) <= not((layer1_outputs(1996)) and (layer1_outputs(6802)));
    layer2_outputs(6448) <= (layer1_outputs(10837)) and (layer1_outputs(1672));
    layer2_outputs(6449) <= layer1_outputs(6668);
    layer2_outputs(6450) <= not(layer1_outputs(2418));
    layer2_outputs(6451) <= not(layer1_outputs(9053));
    layer2_outputs(6452) <= not(layer1_outputs(1226)) or (layer1_outputs(11667));
    layer2_outputs(6453) <= not(layer1_outputs(9371));
    layer2_outputs(6454) <= not((layer1_outputs(5725)) or (layer1_outputs(3820)));
    layer2_outputs(6455) <= layer1_outputs(5621);
    layer2_outputs(6456) <= not(layer1_outputs(1507));
    layer2_outputs(6457) <= not((layer1_outputs(3459)) and (layer1_outputs(7104)));
    layer2_outputs(6458) <= (layer1_outputs(11101)) and (layer1_outputs(1503));
    layer2_outputs(6459) <= layer1_outputs(2824);
    layer2_outputs(6460) <= (layer1_outputs(5085)) and (layer1_outputs(6640));
    layer2_outputs(6461) <= layer1_outputs(11785);
    layer2_outputs(6462) <= not(layer1_outputs(9519));
    layer2_outputs(6463) <= (layer1_outputs(8002)) xor (layer1_outputs(9977));
    layer2_outputs(6464) <= (layer1_outputs(11577)) or (layer1_outputs(440));
    layer2_outputs(6465) <= layer1_outputs(9836);
    layer2_outputs(6466) <= not((layer1_outputs(5859)) xor (layer1_outputs(546)));
    layer2_outputs(6467) <= not((layer1_outputs(9409)) and (layer1_outputs(5392)));
    layer2_outputs(6468) <= not(layer1_outputs(2377));
    layer2_outputs(6469) <= layer1_outputs(2884);
    layer2_outputs(6470) <= layer1_outputs(8454);
    layer2_outputs(6471) <= not((layer1_outputs(4161)) or (layer1_outputs(8159)));
    layer2_outputs(6472) <= layer1_outputs(11407);
    layer2_outputs(6473) <= (layer1_outputs(9334)) or (layer1_outputs(7393));
    layer2_outputs(6474) <= not((layer1_outputs(7279)) xor (layer1_outputs(7045)));
    layer2_outputs(6475) <= not(layer1_outputs(5947));
    layer2_outputs(6476) <= not(layer1_outputs(10059));
    layer2_outputs(6477) <= (layer1_outputs(2410)) and not (layer1_outputs(1123));
    layer2_outputs(6478) <= not(layer1_outputs(2869));
    layer2_outputs(6479) <= not(layer1_outputs(1320));
    layer2_outputs(6480) <= not(layer1_outputs(1264)) or (layer1_outputs(10074));
    layer2_outputs(6481) <= (layer1_outputs(2474)) and not (layer1_outputs(898));
    layer2_outputs(6482) <= (layer1_outputs(7459)) and not (layer1_outputs(6058));
    layer2_outputs(6483) <= layer1_outputs(10324);
    layer2_outputs(6484) <= not(layer1_outputs(4154)) or (layer1_outputs(7737));
    layer2_outputs(6485) <= layer1_outputs(10041);
    layer2_outputs(6486) <= not(layer1_outputs(11480));
    layer2_outputs(6487) <= layer1_outputs(9202);
    layer2_outputs(6488) <= not(layer1_outputs(8722));
    layer2_outputs(6489) <= not(layer1_outputs(9946));
    layer2_outputs(6490) <= not(layer1_outputs(5164));
    layer2_outputs(6491) <= layer1_outputs(2566);
    layer2_outputs(6492) <= layer1_outputs(11946);
    layer2_outputs(6493) <= layer1_outputs(3365);
    layer2_outputs(6494) <= not(layer1_outputs(12074)) or (layer1_outputs(5247));
    layer2_outputs(6495) <= not(layer1_outputs(5616)) or (layer1_outputs(1325));
    layer2_outputs(6496) <= layer1_outputs(807);
    layer2_outputs(6497) <= '1';
    layer2_outputs(6498) <= layer1_outputs(1192);
    layer2_outputs(6499) <= layer1_outputs(8887);
    layer2_outputs(6500) <= not((layer1_outputs(2235)) and (layer1_outputs(5604)));
    layer2_outputs(6501) <= (layer1_outputs(8983)) and (layer1_outputs(776));
    layer2_outputs(6502) <= not((layer1_outputs(999)) xor (layer1_outputs(3820)));
    layer2_outputs(6503) <= layer1_outputs(2479);
    layer2_outputs(6504) <= not(layer1_outputs(8576));
    layer2_outputs(6505) <= layer1_outputs(11489);
    layer2_outputs(6506) <= (layer1_outputs(11258)) xor (layer1_outputs(6555));
    layer2_outputs(6507) <= layer1_outputs(9764);
    layer2_outputs(6508) <= layer1_outputs(796);
    layer2_outputs(6509) <= (layer1_outputs(9387)) or (layer1_outputs(11828));
    layer2_outputs(6510) <= layer1_outputs(5133);
    layer2_outputs(6511) <= (layer1_outputs(7355)) or (layer1_outputs(10616));
    layer2_outputs(6512) <= layer1_outputs(10563);
    layer2_outputs(6513) <= not(layer1_outputs(1097));
    layer2_outputs(6514) <= layer1_outputs(9504);
    layer2_outputs(6515) <= not((layer1_outputs(10869)) xor (layer1_outputs(3195)));
    layer2_outputs(6516) <= layer1_outputs(4285);
    layer2_outputs(6517) <= not(layer1_outputs(10469));
    layer2_outputs(6518) <= not(layer1_outputs(9328));
    layer2_outputs(6519) <= not((layer1_outputs(8188)) xor (layer1_outputs(695)));
    layer2_outputs(6520) <= not(layer1_outputs(7317));
    layer2_outputs(6521) <= layer1_outputs(2444);
    layer2_outputs(6522) <= not((layer1_outputs(4983)) and (layer1_outputs(118)));
    layer2_outputs(6523) <= not(layer1_outputs(296));
    layer2_outputs(6524) <= not(layer1_outputs(23));
    layer2_outputs(6525) <= (layer1_outputs(5022)) xor (layer1_outputs(10078));
    layer2_outputs(6526) <= layer1_outputs(11869);
    layer2_outputs(6527) <= layer1_outputs(4317);
    layer2_outputs(6528) <= not(layer1_outputs(7960));
    layer2_outputs(6529) <= '0';
    layer2_outputs(6530) <= layer1_outputs(6753);
    layer2_outputs(6531) <= not(layer1_outputs(11867));
    layer2_outputs(6532) <= '1';
    layer2_outputs(6533) <= not(layer1_outputs(7310));
    layer2_outputs(6534) <= layer1_outputs(4313);
    layer2_outputs(6535) <= (layer1_outputs(5630)) and not (layer1_outputs(4437));
    layer2_outputs(6536) <= (layer1_outputs(6209)) xor (layer1_outputs(9821));
    layer2_outputs(6537) <= not(layer1_outputs(2722));
    layer2_outputs(6538) <= not(layer1_outputs(76));
    layer2_outputs(6539) <= not(layer1_outputs(9208));
    layer2_outputs(6540) <= not((layer1_outputs(4235)) or (layer1_outputs(1868)));
    layer2_outputs(6541) <= not(layer1_outputs(4014));
    layer2_outputs(6542) <= not(layer1_outputs(10299));
    layer2_outputs(6543) <= (layer1_outputs(860)) xor (layer1_outputs(12586));
    layer2_outputs(6544) <= (layer1_outputs(4484)) xor (layer1_outputs(6433));
    layer2_outputs(6545) <= not(layer1_outputs(4097));
    layer2_outputs(6546) <= not((layer1_outputs(11650)) xor (layer1_outputs(12765)));
    layer2_outputs(6547) <= (layer1_outputs(2174)) or (layer1_outputs(6968));
    layer2_outputs(6548) <= not(layer1_outputs(11456));
    layer2_outputs(6549) <= not((layer1_outputs(2438)) and (layer1_outputs(9322)));
    layer2_outputs(6550) <= not(layer1_outputs(7825)) or (layer1_outputs(3264));
    layer2_outputs(6551) <= (layer1_outputs(7581)) and (layer1_outputs(6095));
    layer2_outputs(6552) <= (layer1_outputs(11874)) and not (layer1_outputs(1344));
    layer2_outputs(6553) <= not(layer1_outputs(9487));
    layer2_outputs(6554) <= not(layer1_outputs(3595)) or (layer1_outputs(5843));
    layer2_outputs(6555) <= not(layer1_outputs(11010));
    layer2_outputs(6556) <= not((layer1_outputs(1644)) xor (layer1_outputs(4533)));
    layer2_outputs(6557) <= not((layer1_outputs(4435)) or (layer1_outputs(4963)));
    layer2_outputs(6558) <= not(layer1_outputs(5369));
    layer2_outputs(6559) <= layer1_outputs(4814);
    layer2_outputs(6560) <= (layer1_outputs(10360)) and not (layer1_outputs(604));
    layer2_outputs(6561) <= layer1_outputs(7161);
    layer2_outputs(6562) <= (layer1_outputs(1204)) and (layer1_outputs(5669));
    layer2_outputs(6563) <= not((layer1_outputs(5316)) and (layer1_outputs(1801)));
    layer2_outputs(6564) <= not(layer1_outputs(293)) or (layer1_outputs(1180));
    layer2_outputs(6565) <= not(layer1_outputs(2904));
    layer2_outputs(6566) <= not((layer1_outputs(11729)) or (layer1_outputs(557)));
    layer2_outputs(6567) <= (layer1_outputs(8899)) and not (layer1_outputs(537));
    layer2_outputs(6568) <= not((layer1_outputs(5578)) and (layer1_outputs(8674)));
    layer2_outputs(6569) <= not((layer1_outputs(8215)) and (layer1_outputs(2780)));
    layer2_outputs(6570) <= (layer1_outputs(890)) and not (layer1_outputs(12425));
    layer2_outputs(6571) <= layer1_outputs(991);
    layer2_outputs(6572) <= not(layer1_outputs(9436));
    layer2_outputs(6573) <= layer1_outputs(4273);
    layer2_outputs(6574) <= not(layer1_outputs(10992));
    layer2_outputs(6575) <= not(layer1_outputs(10511)) or (layer1_outputs(6838));
    layer2_outputs(6576) <= not(layer1_outputs(7090));
    layer2_outputs(6577) <= not((layer1_outputs(2389)) xor (layer1_outputs(1717)));
    layer2_outputs(6578) <= layer1_outputs(9371);
    layer2_outputs(6579) <= layer1_outputs(10849);
    layer2_outputs(6580) <= (layer1_outputs(7603)) xor (layer1_outputs(3482));
    layer2_outputs(6581) <= not(layer1_outputs(1863));
    layer2_outputs(6582) <= layer1_outputs(719);
    layer2_outputs(6583) <= (layer1_outputs(12091)) and not (layer1_outputs(1215));
    layer2_outputs(6584) <= not(layer1_outputs(10514));
    layer2_outputs(6585) <= (layer1_outputs(2581)) and not (layer1_outputs(7425));
    layer2_outputs(6586) <= not(layer1_outputs(8888)) or (layer1_outputs(10914));
    layer2_outputs(6587) <= layer1_outputs(10866);
    layer2_outputs(6588) <= not(layer1_outputs(8196));
    layer2_outputs(6589) <= not((layer1_outputs(11936)) xor (layer1_outputs(6182)));
    layer2_outputs(6590) <= '1';
    layer2_outputs(6591) <= not(layer1_outputs(9116));
    layer2_outputs(6592) <= layer1_outputs(5070);
    layer2_outputs(6593) <= layer1_outputs(2861);
    layer2_outputs(6594) <= (layer1_outputs(9428)) and not (layer1_outputs(9470));
    layer2_outputs(6595) <= not(layer1_outputs(8606));
    layer2_outputs(6596) <= layer1_outputs(6730);
    layer2_outputs(6597) <= not(layer1_outputs(3455));
    layer2_outputs(6598) <= (layer1_outputs(9466)) and (layer1_outputs(426));
    layer2_outputs(6599) <= layer1_outputs(9823);
    layer2_outputs(6600) <= not((layer1_outputs(2168)) xor (layer1_outputs(9895)));
    layer2_outputs(6601) <= (layer1_outputs(5606)) and not (layer1_outputs(6907));
    layer2_outputs(6602) <= (layer1_outputs(11674)) xor (layer1_outputs(7722));
    layer2_outputs(6603) <= layer1_outputs(22);
    layer2_outputs(6604) <= (layer1_outputs(8034)) or (layer1_outputs(10499));
    layer2_outputs(6605) <= (layer1_outputs(6823)) or (layer1_outputs(10783));
    layer2_outputs(6606) <= layer1_outputs(11137);
    layer2_outputs(6607) <= (layer1_outputs(9095)) and not (layer1_outputs(7792));
    layer2_outputs(6608) <= not((layer1_outputs(3808)) xor (layer1_outputs(10718)));
    layer2_outputs(6609) <= layer1_outputs(12293);
    layer2_outputs(6610) <= not((layer1_outputs(8622)) xor (layer1_outputs(2823)));
    layer2_outputs(6611) <= not((layer1_outputs(5308)) and (layer1_outputs(2172)));
    layer2_outputs(6612) <= (layer1_outputs(11393)) xor (layer1_outputs(9757));
    layer2_outputs(6613) <= not((layer1_outputs(7952)) or (layer1_outputs(11387)));
    layer2_outputs(6614) <= layer1_outputs(6210);
    layer2_outputs(6615) <= not(layer1_outputs(1357));
    layer2_outputs(6616) <= not(layer1_outputs(3792));
    layer2_outputs(6617) <= layer1_outputs(4033);
    layer2_outputs(6618) <= (layer1_outputs(1113)) and (layer1_outputs(7773));
    layer2_outputs(6619) <= layer1_outputs(7180);
    layer2_outputs(6620) <= (layer1_outputs(10064)) and not (layer1_outputs(8238));
    layer2_outputs(6621) <= (layer1_outputs(10580)) xor (layer1_outputs(7670));
    layer2_outputs(6622) <= (layer1_outputs(4100)) and (layer1_outputs(7973));
    layer2_outputs(6623) <= not(layer1_outputs(8764));
    layer2_outputs(6624) <= layer1_outputs(11000);
    layer2_outputs(6625) <= not(layer1_outputs(142));
    layer2_outputs(6626) <= layer1_outputs(6866);
    layer2_outputs(6627) <= (layer1_outputs(4209)) xor (layer1_outputs(5799));
    layer2_outputs(6628) <= not(layer1_outputs(994));
    layer2_outputs(6629) <= not((layer1_outputs(5562)) xor (layer1_outputs(139)));
    layer2_outputs(6630) <= layer1_outputs(8765);
    layer2_outputs(6631) <= layer1_outputs(3642);
    layer2_outputs(6632) <= not(layer1_outputs(2460));
    layer2_outputs(6633) <= (layer1_outputs(11908)) or (layer1_outputs(10193));
    layer2_outputs(6634) <= layer1_outputs(8967);
    layer2_outputs(6635) <= layer1_outputs(77);
    layer2_outputs(6636) <= layer1_outputs(2243);
    layer2_outputs(6637) <= layer1_outputs(5966);
    layer2_outputs(6638) <= not(layer1_outputs(6910));
    layer2_outputs(6639) <= not((layer1_outputs(2476)) and (layer1_outputs(9450)));
    layer2_outputs(6640) <= not(layer1_outputs(8939));
    layer2_outputs(6641) <= (layer1_outputs(6560)) xor (layer1_outputs(12519));
    layer2_outputs(6642) <= (layer1_outputs(1919)) and not (layer1_outputs(8454));
    layer2_outputs(6643) <= layer1_outputs(9237);
    layer2_outputs(6644) <= (layer1_outputs(3752)) and not (layer1_outputs(7073));
    layer2_outputs(6645) <= layer1_outputs(11837);
    layer2_outputs(6646) <= not(layer1_outputs(4744));
    layer2_outputs(6647) <= not(layer1_outputs(8989)) or (layer1_outputs(1223));
    layer2_outputs(6648) <= (layer1_outputs(6140)) or (layer1_outputs(9905));
    layer2_outputs(6649) <= not((layer1_outputs(6227)) or (layer1_outputs(11988)));
    layer2_outputs(6650) <= layer1_outputs(3022);
    layer2_outputs(6651) <= layer1_outputs(4120);
    layer2_outputs(6652) <= (layer1_outputs(6668)) or (layer1_outputs(6975));
    layer2_outputs(6653) <= (layer1_outputs(6574)) and (layer1_outputs(9982));
    layer2_outputs(6654) <= not((layer1_outputs(643)) xor (layer1_outputs(10612)));
    layer2_outputs(6655) <= (layer1_outputs(10178)) and not (layer1_outputs(8390));
    layer2_outputs(6656) <= not(layer1_outputs(11973));
    layer2_outputs(6657) <= layer1_outputs(1942);
    layer2_outputs(6658) <= layer1_outputs(8407);
    layer2_outputs(6659) <= not(layer1_outputs(4358));
    layer2_outputs(6660) <= not((layer1_outputs(6807)) xor (layer1_outputs(1251)));
    layer2_outputs(6661) <= layer1_outputs(12211);
    layer2_outputs(6662) <= not(layer1_outputs(9628));
    layer2_outputs(6663) <= (layer1_outputs(11312)) and not (layer1_outputs(9238));
    layer2_outputs(6664) <= not(layer1_outputs(8037));
    layer2_outputs(6665) <= layer1_outputs(4864);
    layer2_outputs(6666) <= (layer1_outputs(6953)) xor (layer1_outputs(4901));
    layer2_outputs(6667) <= layer1_outputs(6019);
    layer2_outputs(6668) <= not(layer1_outputs(773));
    layer2_outputs(6669) <= (layer1_outputs(10471)) or (layer1_outputs(429));
    layer2_outputs(6670) <= not(layer1_outputs(12704));
    layer2_outputs(6671) <= not((layer1_outputs(10097)) or (layer1_outputs(9558)));
    layer2_outputs(6672) <= layer1_outputs(2765);
    layer2_outputs(6673) <= not(layer1_outputs(4703));
    layer2_outputs(6674) <= (layer1_outputs(8081)) and not (layer1_outputs(6448));
    layer2_outputs(6675) <= not(layer1_outputs(3159)) or (layer1_outputs(4347));
    layer2_outputs(6676) <= layer1_outputs(3849);
    layer2_outputs(6677) <= not((layer1_outputs(5286)) xor (layer1_outputs(2086)));
    layer2_outputs(6678) <= layer1_outputs(4368);
    layer2_outputs(6679) <= not((layer1_outputs(2568)) xor (layer1_outputs(8971)));
    layer2_outputs(6680) <= not(layer1_outputs(11531)) or (layer1_outputs(7843));
    layer2_outputs(6681) <= layer1_outputs(2406);
    layer2_outputs(6682) <= not(layer1_outputs(2157));
    layer2_outputs(6683) <= not(layer1_outputs(5711));
    layer2_outputs(6684) <= not(layer1_outputs(10856));
    layer2_outputs(6685) <= layer1_outputs(7983);
    layer2_outputs(6686) <= layer1_outputs(419);
    layer2_outputs(6687) <= not(layer1_outputs(6798));
    layer2_outputs(6688) <= not(layer1_outputs(12471));
    layer2_outputs(6689) <= layer1_outputs(11626);
    layer2_outputs(6690) <= layer1_outputs(4454);
    layer2_outputs(6691) <= layer1_outputs(1322);
    layer2_outputs(6692) <= not(layer1_outputs(8461)) or (layer1_outputs(11992));
    layer2_outputs(6693) <= not((layer1_outputs(5005)) or (layer1_outputs(1823)));
    layer2_outputs(6694) <= not(layer1_outputs(8388)) or (layer1_outputs(7964));
    layer2_outputs(6695) <= (layer1_outputs(5108)) xor (layer1_outputs(12618));
    layer2_outputs(6696) <= not((layer1_outputs(4071)) and (layer1_outputs(6863)));
    layer2_outputs(6697) <= not((layer1_outputs(12026)) xor (layer1_outputs(10434)));
    layer2_outputs(6698) <= not(layer1_outputs(12050));
    layer2_outputs(6699) <= not(layer1_outputs(6154));
    layer2_outputs(6700) <= not(layer1_outputs(12495));
    layer2_outputs(6701) <= '1';
    layer2_outputs(6702) <= layer1_outputs(345);
    layer2_outputs(6703) <= not((layer1_outputs(6461)) or (layer1_outputs(2871)));
    layer2_outputs(6704) <= not(layer1_outputs(4511));
    layer2_outputs(6705) <= (layer1_outputs(601)) and not (layer1_outputs(11220));
    layer2_outputs(6706) <= layer1_outputs(1409);
    layer2_outputs(6707) <= '0';
    layer2_outputs(6708) <= layer1_outputs(8245);
    layer2_outputs(6709) <= (layer1_outputs(8636)) and (layer1_outputs(10714));
    layer2_outputs(6710) <= not(layer1_outputs(2585)) or (layer1_outputs(12728));
    layer2_outputs(6711) <= layer1_outputs(11325);
    layer2_outputs(6712) <= (layer1_outputs(3187)) and (layer1_outputs(2811));
    layer2_outputs(6713) <= layer1_outputs(3058);
    layer2_outputs(6714) <= not(layer1_outputs(1955));
    layer2_outputs(6715) <= not(layer1_outputs(11608));
    layer2_outputs(6716) <= not((layer1_outputs(5753)) xor (layer1_outputs(166)));
    layer2_outputs(6717) <= layer1_outputs(7847);
    layer2_outputs(6718) <= not((layer1_outputs(3050)) and (layer1_outputs(9036)));
    layer2_outputs(6719) <= not(layer1_outputs(2298));
    layer2_outputs(6720) <= not((layer1_outputs(6597)) xor (layer1_outputs(8995)));
    layer2_outputs(6721) <= '0';
    layer2_outputs(6722) <= layer1_outputs(9318);
    layer2_outputs(6723) <= layer1_outputs(5361);
    layer2_outputs(6724) <= not(layer1_outputs(1223));
    layer2_outputs(6725) <= layer1_outputs(8611);
    layer2_outputs(6726) <= layer1_outputs(250);
    layer2_outputs(6727) <= '1';
    layer2_outputs(6728) <= not(layer1_outputs(9768));
    layer2_outputs(6729) <= (layer1_outputs(8632)) and not (layer1_outputs(5320));
    layer2_outputs(6730) <= (layer1_outputs(7262)) xor (layer1_outputs(11564));
    layer2_outputs(6731) <= layer1_outputs(1677);
    layer2_outputs(6732) <= not(layer1_outputs(8232));
    layer2_outputs(6733) <= not(layer1_outputs(6792));
    layer2_outputs(6734) <= layer1_outputs(991);
    layer2_outputs(6735) <= layer1_outputs(12533);
    layer2_outputs(6736) <= layer1_outputs(10836);
    layer2_outputs(6737) <= not((layer1_outputs(2011)) or (layer1_outputs(11513)));
    layer2_outputs(6738) <= not((layer1_outputs(9418)) xor (layer1_outputs(6617)));
    layer2_outputs(6739) <= (layer1_outputs(2321)) and not (layer1_outputs(6056));
    layer2_outputs(6740) <= not((layer1_outputs(11740)) and (layer1_outputs(525)));
    layer2_outputs(6741) <= not((layer1_outputs(8710)) and (layer1_outputs(5646)));
    layer2_outputs(6742) <= layer1_outputs(8159);
    layer2_outputs(6743) <= not((layer1_outputs(10671)) and (layer1_outputs(12706)));
    layer2_outputs(6744) <= layer1_outputs(9712);
    layer2_outputs(6745) <= not((layer1_outputs(12730)) xor (layer1_outputs(2452)));
    layer2_outputs(6746) <= (layer1_outputs(4476)) or (layer1_outputs(9611));
    layer2_outputs(6747) <= layer1_outputs(12571);
    layer2_outputs(6748) <= not((layer1_outputs(10131)) xor (layer1_outputs(4102)));
    layer2_outputs(6749) <= not(layer1_outputs(5436)) or (layer1_outputs(6216));
    layer2_outputs(6750) <= not(layer1_outputs(5967));
    layer2_outputs(6751) <= layer1_outputs(10217);
    layer2_outputs(6752) <= not(layer1_outputs(220));
    layer2_outputs(6753) <= not(layer1_outputs(9081));
    layer2_outputs(6754) <= not(layer1_outputs(851)) or (layer1_outputs(3669));
    layer2_outputs(6755) <= not((layer1_outputs(8219)) or (layer1_outputs(12423)));
    layer2_outputs(6756) <= (layer1_outputs(8598)) and not (layer1_outputs(6302));
    layer2_outputs(6757) <= (layer1_outputs(12002)) or (layer1_outputs(276));
    layer2_outputs(6758) <= layer1_outputs(6536);
    layer2_outputs(6759) <= (layer1_outputs(5759)) xor (layer1_outputs(9848));
    layer2_outputs(6760) <= layer1_outputs(3275);
    layer2_outputs(6761) <= not((layer1_outputs(9412)) xor (layer1_outputs(5512)));
    layer2_outputs(6762) <= layer1_outputs(10128);
    layer2_outputs(6763) <= not(layer1_outputs(752));
    layer2_outputs(6764) <= layer1_outputs(7021);
    layer2_outputs(6765) <= not(layer1_outputs(4005));
    layer2_outputs(6766) <= not(layer1_outputs(791));
    layer2_outputs(6767) <= not((layer1_outputs(1948)) and (layer1_outputs(2868)));
    layer2_outputs(6768) <= layer1_outputs(9472);
    layer2_outputs(6769) <= (layer1_outputs(7855)) and (layer1_outputs(5446));
    layer2_outputs(6770) <= not((layer1_outputs(3196)) xor (layer1_outputs(4901)));
    layer2_outputs(6771) <= (layer1_outputs(484)) xor (layer1_outputs(6336));
    layer2_outputs(6772) <= layer1_outputs(11873);
    layer2_outputs(6773) <= not((layer1_outputs(10648)) xor (layer1_outputs(1342)));
    layer2_outputs(6774) <= not(layer1_outputs(1762));
    layer2_outputs(6775) <= (layer1_outputs(6748)) and (layer1_outputs(12774));
    layer2_outputs(6776) <= not(layer1_outputs(722));
    layer2_outputs(6777) <= (layer1_outputs(5696)) and (layer1_outputs(10791));
    layer2_outputs(6778) <= layer1_outputs(12556);
    layer2_outputs(6779) <= layer1_outputs(4978);
    layer2_outputs(6780) <= (layer1_outputs(8328)) and (layer1_outputs(9228));
    layer2_outputs(6781) <= not(layer1_outputs(111));
    layer2_outputs(6782) <= not(layer1_outputs(11330));
    layer2_outputs(6783) <= not((layer1_outputs(10636)) xor (layer1_outputs(7266)));
    layer2_outputs(6784) <= not(layer1_outputs(7392));
    layer2_outputs(6785) <= layer1_outputs(10405);
    layer2_outputs(6786) <= not(layer1_outputs(7440));
    layer2_outputs(6787) <= not((layer1_outputs(11076)) or (layer1_outputs(10310)));
    layer2_outputs(6788) <= (layer1_outputs(6619)) and not (layer1_outputs(10117));
    layer2_outputs(6789) <= not(layer1_outputs(5253)) or (layer1_outputs(5252));
    layer2_outputs(6790) <= layer1_outputs(10736);
    layer2_outputs(6791) <= layer1_outputs(8566);
    layer2_outputs(6792) <= (layer1_outputs(5485)) or (layer1_outputs(3073));
    layer2_outputs(6793) <= (layer1_outputs(398)) and (layer1_outputs(2991));
    layer2_outputs(6794) <= not(layer1_outputs(986));
    layer2_outputs(6795) <= (layer1_outputs(3096)) and not (layer1_outputs(5245));
    layer2_outputs(6796) <= layer1_outputs(1982);
    layer2_outputs(6797) <= layer1_outputs(7975);
    layer2_outputs(6798) <= not((layer1_outputs(1731)) and (layer1_outputs(12730)));
    layer2_outputs(6799) <= (layer1_outputs(2512)) or (layer1_outputs(1489));
    layer2_outputs(6800) <= not(layer1_outputs(3162)) or (layer1_outputs(9974));
    layer2_outputs(6801) <= (layer1_outputs(12569)) or (layer1_outputs(11819));
    layer2_outputs(6802) <= not(layer1_outputs(8892)) or (layer1_outputs(9780));
    layer2_outputs(6803) <= layer1_outputs(7640);
    layer2_outputs(6804) <= not(layer1_outputs(10482));
    layer2_outputs(6805) <= (layer1_outputs(4089)) xor (layer1_outputs(8488));
    layer2_outputs(6806) <= layer1_outputs(1481);
    layer2_outputs(6807) <= layer1_outputs(5835);
    layer2_outputs(6808) <= not(layer1_outputs(6340));
    layer2_outputs(6809) <= not(layer1_outputs(6231));
    layer2_outputs(6810) <= not((layer1_outputs(4542)) xor (layer1_outputs(6348)));
    layer2_outputs(6811) <= not(layer1_outputs(2409));
    layer2_outputs(6812) <= not(layer1_outputs(12644));
    layer2_outputs(6813) <= not(layer1_outputs(83));
    layer2_outputs(6814) <= not((layer1_outputs(8901)) xor (layer1_outputs(5874)));
    layer2_outputs(6815) <= not((layer1_outputs(12493)) or (layer1_outputs(2156)));
    layer2_outputs(6816) <= (layer1_outputs(118)) and not (layer1_outputs(3239));
    layer2_outputs(6817) <= (layer1_outputs(765)) xor (layer1_outputs(7993));
    layer2_outputs(6818) <= layer1_outputs(6539);
    layer2_outputs(6819) <= not(layer1_outputs(9381));
    layer2_outputs(6820) <= layer1_outputs(271);
    layer2_outputs(6821) <= not((layer1_outputs(5668)) xor (layer1_outputs(7446)));
    layer2_outputs(6822) <= not(layer1_outputs(7696));
    layer2_outputs(6823) <= not((layer1_outputs(9396)) and (layer1_outputs(10934)));
    layer2_outputs(6824) <= not(layer1_outputs(10703));
    layer2_outputs(6825) <= not((layer1_outputs(5595)) or (layer1_outputs(8045)));
    layer2_outputs(6826) <= layer1_outputs(8068);
    layer2_outputs(6827) <= (layer1_outputs(683)) xor (layer1_outputs(9024));
    layer2_outputs(6828) <= layer1_outputs(11402);
    layer2_outputs(6829) <= not(layer1_outputs(6650));
    layer2_outputs(6830) <= (layer1_outputs(2446)) and (layer1_outputs(455));
    layer2_outputs(6831) <= not((layer1_outputs(4050)) and (layer1_outputs(8311)));
    layer2_outputs(6832) <= not(layer1_outputs(11625));
    layer2_outputs(6833) <= not((layer1_outputs(4844)) xor (layer1_outputs(12303)));
    layer2_outputs(6834) <= not(layer1_outputs(4505));
    layer2_outputs(6835) <= layer1_outputs(5472);
    layer2_outputs(6836) <= not((layer1_outputs(9571)) xor (layer1_outputs(8206)));
    layer2_outputs(6837) <= not(layer1_outputs(1118));
    layer2_outputs(6838) <= not(layer1_outputs(10807));
    layer2_outputs(6839) <= not(layer1_outputs(5051));
    layer2_outputs(6840) <= not(layer1_outputs(8755));
    layer2_outputs(6841) <= (layer1_outputs(4021)) xor (layer1_outputs(6595));
    layer2_outputs(6842) <= (layer1_outputs(9375)) or (layer1_outputs(6347));
    layer2_outputs(6843) <= layer1_outputs(9925);
    layer2_outputs(6844) <= not((layer1_outputs(1628)) and (layer1_outputs(7681)));
    layer2_outputs(6845) <= not(layer1_outputs(9137));
    layer2_outputs(6846) <= not((layer1_outputs(1926)) and (layer1_outputs(9800)));
    layer2_outputs(6847) <= layer1_outputs(7673);
    layer2_outputs(6848) <= layer1_outputs(9442);
    layer2_outputs(6849) <= not(layer1_outputs(5075));
    layer2_outputs(6850) <= (layer1_outputs(9483)) xor (layer1_outputs(11286));
    layer2_outputs(6851) <= layer1_outputs(9715);
    layer2_outputs(6852) <= (layer1_outputs(5464)) and (layer1_outputs(9391));
    layer2_outputs(6853) <= not(layer1_outputs(4472)) or (layer1_outputs(8840));
    layer2_outputs(6854) <= not(layer1_outputs(3851));
    layer2_outputs(6855) <= layer1_outputs(11451);
    layer2_outputs(6856) <= (layer1_outputs(7522)) or (layer1_outputs(3177));
    layer2_outputs(6857) <= layer1_outputs(5734);
    layer2_outputs(6858) <= not(layer1_outputs(618));
    layer2_outputs(6859) <= not(layer1_outputs(5443));
    layer2_outputs(6860) <= not(layer1_outputs(4515));
    layer2_outputs(6861) <= not((layer1_outputs(9094)) and (layer1_outputs(12471)));
    layer2_outputs(6862) <= layer1_outputs(6148);
    layer2_outputs(6863) <= layer1_outputs(1445);
    layer2_outputs(6864) <= not(layer1_outputs(12521));
    layer2_outputs(6865) <= (layer1_outputs(8092)) or (layer1_outputs(458));
    layer2_outputs(6866) <= not(layer1_outputs(184));
    layer2_outputs(6867) <= (layer1_outputs(8610)) and not (layer1_outputs(4942));
    layer2_outputs(6868) <= (layer1_outputs(7296)) and not (layer1_outputs(4312));
    layer2_outputs(6869) <= (layer1_outputs(12111)) or (layer1_outputs(8894));
    layer2_outputs(6870) <= not(layer1_outputs(2328)) or (layer1_outputs(5914));
    layer2_outputs(6871) <= layer1_outputs(10783);
    layer2_outputs(6872) <= not(layer1_outputs(10699)) or (layer1_outputs(6653));
    layer2_outputs(6873) <= not(layer1_outputs(5850));
    layer2_outputs(6874) <= not((layer1_outputs(5958)) and (layer1_outputs(1396)));
    layer2_outputs(6875) <= not(layer1_outputs(11786)) or (layer1_outputs(6504));
    layer2_outputs(6876) <= layer1_outputs(11819);
    layer2_outputs(6877) <= not(layer1_outputs(1163)) or (layer1_outputs(1871));
    layer2_outputs(6878) <= (layer1_outputs(4253)) and (layer1_outputs(12322));
    layer2_outputs(6879) <= not(layer1_outputs(9488));
    layer2_outputs(6880) <= not(layer1_outputs(5935));
    layer2_outputs(6881) <= layer1_outputs(2787);
    layer2_outputs(6882) <= not(layer1_outputs(8515));
    layer2_outputs(6883) <= not(layer1_outputs(6240)) or (layer1_outputs(11348));
    layer2_outputs(6884) <= not(layer1_outputs(8015)) or (layer1_outputs(12073));
    layer2_outputs(6885) <= not(layer1_outputs(2126)) or (layer1_outputs(3192));
    layer2_outputs(6886) <= layer1_outputs(10815);
    layer2_outputs(6887) <= not(layer1_outputs(10786));
    layer2_outputs(6888) <= not(layer1_outputs(5659)) or (layer1_outputs(3399));
    layer2_outputs(6889) <= not((layer1_outputs(5042)) and (layer1_outputs(7700)));
    layer2_outputs(6890) <= not((layer1_outputs(5356)) xor (layer1_outputs(553)));
    layer2_outputs(6891) <= not(layer1_outputs(1093));
    layer2_outputs(6892) <= (layer1_outputs(6952)) xor (layer1_outputs(4583));
    layer2_outputs(6893) <= (layer1_outputs(692)) or (layer1_outputs(8961));
    layer2_outputs(6894) <= not(layer1_outputs(6959));
    layer2_outputs(6895) <= layer1_outputs(2748);
    layer2_outputs(6896) <= (layer1_outputs(7886)) xor (layer1_outputs(8934));
    layer2_outputs(6897) <= (layer1_outputs(12125)) and not (layer1_outputs(3698));
    layer2_outputs(6898) <= layer1_outputs(6002);
    layer2_outputs(6899) <= not(layer1_outputs(10464));
    layer2_outputs(6900) <= (layer1_outputs(6398)) and not (layer1_outputs(3918));
    layer2_outputs(6901) <= layer1_outputs(9941);
    layer2_outputs(6902) <= not((layer1_outputs(6899)) and (layer1_outputs(9109)));
    layer2_outputs(6903) <= layer1_outputs(4230);
    layer2_outputs(6904) <= not((layer1_outputs(5590)) xor (layer1_outputs(7426)));
    layer2_outputs(6905) <= not(layer1_outputs(4153));
    layer2_outputs(6906) <= (layer1_outputs(10499)) and not (layer1_outputs(7843));
    layer2_outputs(6907) <= layer1_outputs(3238);
    layer2_outputs(6908) <= (layer1_outputs(3739)) or (layer1_outputs(9777));
    layer2_outputs(6909) <= not(layer1_outputs(7223));
    layer2_outputs(6910) <= layer1_outputs(2948);
    layer2_outputs(6911) <= not(layer1_outputs(6660));
    layer2_outputs(6912) <= not((layer1_outputs(7846)) xor (layer1_outputs(4249)));
    layer2_outputs(6913) <= not((layer1_outputs(11234)) and (layer1_outputs(1705)));
    layer2_outputs(6914) <= layer1_outputs(1439);
    layer2_outputs(6915) <= layer1_outputs(3195);
    layer2_outputs(6916) <= not(layer1_outputs(5483));
    layer2_outputs(6917) <= not(layer1_outputs(5267));
    layer2_outputs(6918) <= layer1_outputs(7544);
    layer2_outputs(6919) <= layer1_outputs(751);
    layer2_outputs(6920) <= not(layer1_outputs(6189));
    layer2_outputs(6921) <= not(layer1_outputs(6103)) or (layer1_outputs(12308));
    layer2_outputs(6922) <= not(layer1_outputs(7166)) or (layer1_outputs(1561));
    layer2_outputs(6923) <= (layer1_outputs(3348)) or (layer1_outputs(4143));
    layer2_outputs(6924) <= layer1_outputs(9999);
    layer2_outputs(6925) <= layer1_outputs(4221);
    layer2_outputs(6926) <= layer1_outputs(12221);
    layer2_outputs(6927) <= not(layer1_outputs(8006));
    layer2_outputs(6928) <= not(layer1_outputs(2888));
    layer2_outputs(6929) <= (layer1_outputs(6839)) and (layer1_outputs(4025));
    layer2_outputs(6930) <= not(layer1_outputs(12531));
    layer2_outputs(6931) <= (layer1_outputs(11297)) or (layer1_outputs(9599));
    layer2_outputs(6932) <= (layer1_outputs(10917)) and not (layer1_outputs(8535));
    layer2_outputs(6933) <= not(layer1_outputs(9008));
    layer2_outputs(6934) <= (layer1_outputs(7293)) and (layer1_outputs(70));
    layer2_outputs(6935) <= not(layer1_outputs(11886));
    layer2_outputs(6936) <= not((layer1_outputs(2611)) and (layer1_outputs(2480)));
    layer2_outputs(6937) <= not(layer1_outputs(7543)) or (layer1_outputs(11186));
    layer2_outputs(6938) <= not(layer1_outputs(2894));
    layer2_outputs(6939) <= not((layer1_outputs(8580)) or (layer1_outputs(6330)));
    layer2_outputs(6940) <= layer1_outputs(3682);
    layer2_outputs(6941) <= layer1_outputs(9641);
    layer2_outputs(6942) <= layer1_outputs(7399);
    layer2_outputs(6943) <= (layer1_outputs(7741)) and not (layer1_outputs(9978));
    layer2_outputs(6944) <= not((layer1_outputs(7743)) or (layer1_outputs(4626)));
    layer2_outputs(6945) <= not(layer1_outputs(11711)) or (layer1_outputs(10197));
    layer2_outputs(6946) <= not(layer1_outputs(11408));
    layer2_outputs(6947) <= (layer1_outputs(9212)) and (layer1_outputs(11180));
    layer2_outputs(6948) <= layer1_outputs(9918);
    layer2_outputs(6949) <= layer1_outputs(12413);
    layer2_outputs(6950) <= (layer1_outputs(11162)) or (layer1_outputs(11956));
    layer2_outputs(6951) <= not(layer1_outputs(9088));
    layer2_outputs(6952) <= not(layer1_outputs(9591));
    layer2_outputs(6953) <= not((layer1_outputs(6755)) or (layer1_outputs(5813)));
    layer2_outputs(6954) <= not(layer1_outputs(555));
    layer2_outputs(6955) <= not(layer1_outputs(4295));
    layer2_outputs(6956) <= (layer1_outputs(7297)) and not (layer1_outputs(5648));
    layer2_outputs(6957) <= not(layer1_outputs(7393)) or (layer1_outputs(7467));
    layer2_outputs(6958) <= not(layer1_outputs(7881)) or (layer1_outputs(11930));
    layer2_outputs(6959) <= not(layer1_outputs(7612));
    layer2_outputs(6960) <= layer1_outputs(1880);
    layer2_outputs(6961) <= not(layer1_outputs(8033));
    layer2_outputs(6962) <= not(layer1_outputs(9202));
    layer2_outputs(6963) <= (layer1_outputs(1712)) and not (layer1_outputs(11481));
    layer2_outputs(6964) <= not(layer1_outputs(2048));
    layer2_outputs(6965) <= layer1_outputs(1084);
    layer2_outputs(6966) <= not((layer1_outputs(2138)) and (layer1_outputs(10408)));
    layer2_outputs(6967) <= not(layer1_outputs(8127));
    layer2_outputs(6968) <= (layer1_outputs(11623)) and (layer1_outputs(11022));
    layer2_outputs(6969) <= not(layer1_outputs(10551)) or (layer1_outputs(12777));
    layer2_outputs(6970) <= not(layer1_outputs(10743)) or (layer1_outputs(1650));
    layer2_outputs(6971) <= layer1_outputs(1838);
    layer2_outputs(6972) <= (layer1_outputs(4976)) and not (layer1_outputs(7241));
    layer2_outputs(6973) <= not(layer1_outputs(11071)) or (layer1_outputs(3546));
    layer2_outputs(6974) <= not(layer1_outputs(9523));
    layer2_outputs(6975) <= (layer1_outputs(3186)) or (layer1_outputs(8875));
    layer2_outputs(6976) <= layer1_outputs(10648);
    layer2_outputs(6977) <= layer1_outputs(4277);
    layer2_outputs(6978) <= (layer1_outputs(7839)) xor (layer1_outputs(3468));
    layer2_outputs(6979) <= not(layer1_outputs(1269));
    layer2_outputs(6980) <= not((layer1_outputs(8369)) xor (layer1_outputs(2713)));
    layer2_outputs(6981) <= (layer1_outputs(10009)) and (layer1_outputs(1277));
    layer2_outputs(6982) <= not((layer1_outputs(12434)) or (layer1_outputs(5960)));
    layer2_outputs(6983) <= (layer1_outputs(4451)) and (layer1_outputs(2448));
    layer2_outputs(6984) <= (layer1_outputs(452)) and not (layer1_outputs(9624));
    layer2_outputs(6985) <= not((layer1_outputs(8815)) and (layer1_outputs(4584)));
    layer2_outputs(6986) <= layer1_outputs(1054);
    layer2_outputs(6987) <= not(layer1_outputs(10789));
    layer2_outputs(6988) <= not((layer1_outputs(8038)) and (layer1_outputs(632)));
    layer2_outputs(6989) <= layer1_outputs(2916);
    layer2_outputs(6990) <= not(layer1_outputs(8399));
    layer2_outputs(6991) <= (layer1_outputs(3875)) and (layer1_outputs(6035));
    layer2_outputs(6992) <= layer1_outputs(3775);
    layer2_outputs(6993) <= layer1_outputs(11032);
    layer2_outputs(6994) <= layer1_outputs(6881);
    layer2_outputs(6995) <= not(layer1_outputs(3432));
    layer2_outputs(6996) <= (layer1_outputs(1692)) and (layer1_outputs(3922));
    layer2_outputs(6997) <= layer1_outputs(2725);
    layer2_outputs(6998) <= layer1_outputs(4236);
    layer2_outputs(6999) <= not(layer1_outputs(10378));
    layer2_outputs(7000) <= not(layer1_outputs(3792));
    layer2_outputs(7001) <= (layer1_outputs(7513)) and (layer1_outputs(1493));
    layer2_outputs(7002) <= layer1_outputs(950);
    layer2_outputs(7003) <= (layer1_outputs(963)) xor (layer1_outputs(8740));
    layer2_outputs(7004) <= (layer1_outputs(1529)) and not (layer1_outputs(12080));
    layer2_outputs(7005) <= layer1_outputs(9191);
    layer2_outputs(7006) <= layer1_outputs(8115);
    layer2_outputs(7007) <= (layer1_outputs(11590)) or (layer1_outputs(12333));
    layer2_outputs(7008) <= not(layer1_outputs(815));
    layer2_outputs(7009) <= layer1_outputs(12258);
    layer2_outputs(7010) <= (layer1_outputs(5801)) and not (layer1_outputs(4563));
    layer2_outputs(7011) <= (layer1_outputs(6332)) and (layer1_outputs(8208));
    layer2_outputs(7012) <= (layer1_outputs(12301)) and (layer1_outputs(4877));
    layer2_outputs(7013) <= (layer1_outputs(995)) and not (layer1_outputs(4077));
    layer2_outputs(7014) <= layer1_outputs(10334);
    layer2_outputs(7015) <= (layer1_outputs(7254)) and not (layer1_outputs(4152));
    layer2_outputs(7016) <= not(layer1_outputs(6163));
    layer2_outputs(7017) <= (layer1_outputs(2693)) and (layer1_outputs(6629));
    layer2_outputs(7018) <= layer1_outputs(3663);
    layer2_outputs(7019) <= not(layer1_outputs(2561));
    layer2_outputs(7020) <= (layer1_outputs(5524)) and (layer1_outputs(7668));
    layer2_outputs(7021) <= not((layer1_outputs(12420)) and (layer1_outputs(8397)));
    layer2_outputs(7022) <= not(layer1_outputs(6624));
    layer2_outputs(7023) <= not(layer1_outputs(3221)) or (layer1_outputs(9688));
    layer2_outputs(7024) <= not((layer1_outputs(5778)) xor (layer1_outputs(2647)));
    layer2_outputs(7025) <= layer1_outputs(9220);
    layer2_outputs(7026) <= not((layer1_outputs(11875)) and (layer1_outputs(9585)));
    layer2_outputs(7027) <= (layer1_outputs(3174)) and not (layer1_outputs(4));
    layer2_outputs(7028) <= layer1_outputs(1073);
    layer2_outputs(7029) <= (layer1_outputs(11661)) and not (layer1_outputs(12566));
    layer2_outputs(7030) <= layer1_outputs(9489);
    layer2_outputs(7031) <= not((layer1_outputs(8230)) xor (layer1_outputs(12474)));
    layer2_outputs(7032) <= layer1_outputs(8191);
    layer2_outputs(7033) <= (layer1_outputs(8940)) and (layer1_outputs(2714));
    layer2_outputs(7034) <= (layer1_outputs(7538)) or (layer1_outputs(9293));
    layer2_outputs(7035) <= not((layer1_outputs(7374)) or (layer1_outputs(5803)));
    layer2_outputs(7036) <= not(layer1_outputs(3989)) or (layer1_outputs(7848));
    layer2_outputs(7037) <= layer1_outputs(811);
    layer2_outputs(7038) <= not(layer1_outputs(6061));
    layer2_outputs(7039) <= not(layer1_outputs(9669));
    layer2_outputs(7040) <= (layer1_outputs(7845)) xor (layer1_outputs(12389));
    layer2_outputs(7041) <= not((layer1_outputs(2726)) and (layer1_outputs(3722)));
    layer2_outputs(7042) <= not(layer1_outputs(4744));
    layer2_outputs(7043) <= (layer1_outputs(3896)) and (layer1_outputs(1687));
    layer2_outputs(7044) <= layer1_outputs(9735);
    layer2_outputs(7045) <= layer1_outputs(9715);
    layer2_outputs(7046) <= not((layer1_outputs(961)) and (layer1_outputs(4985)));
    layer2_outputs(7047) <= not((layer1_outputs(1640)) and (layer1_outputs(11412)));
    layer2_outputs(7048) <= '0';
    layer2_outputs(7049) <= not((layer1_outputs(7979)) or (layer1_outputs(1670)));
    layer2_outputs(7050) <= not(layer1_outputs(3106));
    layer2_outputs(7051) <= layer1_outputs(10164);
    layer2_outputs(7052) <= not(layer1_outputs(7411));
    layer2_outputs(7053) <= (layer1_outputs(9703)) and not (layer1_outputs(9673));
    layer2_outputs(7054) <= (layer1_outputs(4399)) or (layer1_outputs(3342));
    layer2_outputs(7055) <= (layer1_outputs(9724)) xor (layer1_outputs(9810));
    layer2_outputs(7056) <= layer1_outputs(10546);
    layer2_outputs(7057) <= not(layer1_outputs(9898));
    layer2_outputs(7058) <= not(layer1_outputs(1235));
    layer2_outputs(7059) <= not((layer1_outputs(3308)) xor (layer1_outputs(11709)));
    layer2_outputs(7060) <= not(layer1_outputs(2576));
    layer2_outputs(7061) <= layer1_outputs(11054);
    layer2_outputs(7062) <= layer1_outputs(8423);
    layer2_outputs(7063) <= not((layer1_outputs(4322)) xor (layer1_outputs(8527)));
    layer2_outputs(7064) <= not((layer1_outputs(10000)) xor (layer1_outputs(2985)));
    layer2_outputs(7065) <= layer1_outputs(4586);
    layer2_outputs(7066) <= not((layer1_outputs(622)) xor (layer1_outputs(6033)));
    layer2_outputs(7067) <= (layer1_outputs(9415)) and not (layer1_outputs(6556));
    layer2_outputs(7068) <= layer1_outputs(10260);
    layer2_outputs(7069) <= not((layer1_outputs(12174)) and (layer1_outputs(402)));
    layer2_outputs(7070) <= layer1_outputs(8145);
    layer2_outputs(7071) <= not(layer1_outputs(6285));
    layer2_outputs(7072) <= not(layer1_outputs(453));
    layer2_outputs(7073) <= (layer1_outputs(5238)) or (layer1_outputs(9816));
    layer2_outputs(7074) <= layer1_outputs(2268);
    layer2_outputs(7075) <= layer1_outputs(743);
    layer2_outputs(7076) <= (layer1_outputs(8022)) or (layer1_outputs(5737));
    layer2_outputs(7077) <= not((layer1_outputs(8855)) or (layer1_outputs(7333)));
    layer2_outputs(7078) <= layer1_outputs(3810);
    layer2_outputs(7079) <= not(layer1_outputs(3160));
    layer2_outputs(7080) <= (layer1_outputs(6421)) and (layer1_outputs(7551));
    layer2_outputs(7081) <= layer1_outputs(7996);
    layer2_outputs(7082) <= not(layer1_outputs(9199)) or (layer1_outputs(6939));
    layer2_outputs(7083) <= layer1_outputs(9208);
    layer2_outputs(7084) <= (layer1_outputs(11373)) and (layer1_outputs(387));
    layer2_outputs(7085) <= (layer1_outputs(5216)) xor (layer1_outputs(12537));
    layer2_outputs(7086) <= (layer1_outputs(6232)) xor (layer1_outputs(1759));
    layer2_outputs(7087) <= (layer1_outputs(11638)) xor (layer1_outputs(8427));
    layer2_outputs(7088) <= not((layer1_outputs(7674)) or (layer1_outputs(12796)));
    layer2_outputs(7089) <= (layer1_outputs(2219)) and not (layer1_outputs(4164));
    layer2_outputs(7090) <= not((layer1_outputs(11783)) or (layer1_outputs(9856)));
    layer2_outputs(7091) <= layer1_outputs(11447);
    layer2_outputs(7092) <= layer1_outputs(3824);
    layer2_outputs(7093) <= not((layer1_outputs(9687)) and (layer1_outputs(7572)));
    layer2_outputs(7094) <= not(layer1_outputs(3389));
    layer2_outputs(7095) <= not((layer1_outputs(4724)) xor (layer1_outputs(950)));
    layer2_outputs(7096) <= (layer1_outputs(2765)) and not (layer1_outputs(3433));
    layer2_outputs(7097) <= not(layer1_outputs(5770)) or (layer1_outputs(1044));
    layer2_outputs(7098) <= not(layer1_outputs(7782)) or (layer1_outputs(5608));
    layer2_outputs(7099) <= (layer1_outputs(6596)) and not (layer1_outputs(10801));
    layer2_outputs(7100) <= layer1_outputs(8591);
    layer2_outputs(7101) <= (layer1_outputs(11832)) or (layer1_outputs(7573));
    layer2_outputs(7102) <= layer1_outputs(10084);
    layer2_outputs(7103) <= not(layer1_outputs(11293));
    layer2_outputs(7104) <= layer1_outputs(7285);
    layer2_outputs(7105) <= layer1_outputs(4735);
    layer2_outputs(7106) <= not(layer1_outputs(7155));
    layer2_outputs(7107) <= not((layer1_outputs(12294)) or (layer1_outputs(1904)));
    layer2_outputs(7108) <= not((layer1_outputs(10131)) and (layer1_outputs(7964)));
    layer2_outputs(7109) <= not(layer1_outputs(12104));
    layer2_outputs(7110) <= not(layer1_outputs(2906));
    layer2_outputs(7111) <= not((layer1_outputs(10436)) xor (layer1_outputs(10627)));
    layer2_outputs(7112) <= layer1_outputs(46);
    layer2_outputs(7113) <= layer1_outputs(10908);
    layer2_outputs(7114) <= layer1_outputs(2356);
    layer2_outputs(7115) <= layer1_outputs(8928);
    layer2_outputs(7116) <= layer1_outputs(7336);
    layer2_outputs(7117) <= not(layer1_outputs(3265)) or (layer1_outputs(3951));
    layer2_outputs(7118) <= layer1_outputs(4758);
    layer2_outputs(7119) <= not(layer1_outputs(1581));
    layer2_outputs(7120) <= not(layer1_outputs(10325));
    layer2_outputs(7121) <= not(layer1_outputs(9916)) or (layer1_outputs(10874));
    layer2_outputs(7122) <= layer1_outputs(4804);
    layer2_outputs(7123) <= (layer1_outputs(2365)) and not (layer1_outputs(4987));
    layer2_outputs(7124) <= not((layer1_outputs(10407)) xor (layer1_outputs(766)));
    layer2_outputs(7125) <= layer1_outputs(6978);
    layer2_outputs(7126) <= not(layer1_outputs(4535));
    layer2_outputs(7127) <= not((layer1_outputs(9076)) or (layer1_outputs(8223)));
    layer2_outputs(7128) <= (layer1_outputs(2154)) and not (layer1_outputs(6429));
    layer2_outputs(7129) <= not((layer1_outputs(9005)) and (layer1_outputs(11467)));
    layer2_outputs(7130) <= not(layer1_outputs(12199));
    layer2_outputs(7131) <= (layer1_outputs(11019)) and not (layer1_outputs(11765));
    layer2_outputs(7132) <= (layer1_outputs(5316)) and not (layer1_outputs(12695));
    layer2_outputs(7133) <= layer1_outputs(9469);
    layer2_outputs(7134) <= not(layer1_outputs(10433));
    layer2_outputs(7135) <= layer1_outputs(7063);
    layer2_outputs(7136) <= not(layer1_outputs(6454));
    layer2_outputs(7137) <= not((layer1_outputs(223)) or (layer1_outputs(5698)));
    layer2_outputs(7138) <= (layer1_outputs(3173)) xor (layer1_outputs(2304));
    layer2_outputs(7139) <= not(layer1_outputs(667));
    layer2_outputs(7140) <= layer1_outputs(10893);
    layer2_outputs(7141) <= not((layer1_outputs(11950)) xor (layer1_outputs(9913)));
    layer2_outputs(7142) <= (layer1_outputs(650)) xor (layer1_outputs(8258));
    layer2_outputs(7143) <= not(layer1_outputs(2450));
    layer2_outputs(7144) <= not((layer1_outputs(12466)) or (layer1_outputs(8010)));
    layer2_outputs(7145) <= not((layer1_outputs(1650)) xor (layer1_outputs(11860)));
    layer2_outputs(7146) <= layer1_outputs(12714);
    layer2_outputs(7147) <= (layer1_outputs(9349)) and not (layer1_outputs(5247));
    layer2_outputs(7148) <= layer1_outputs(7008);
    layer2_outputs(7149) <= (layer1_outputs(6852)) and (layer1_outputs(7327));
    layer2_outputs(7150) <= layer1_outputs(2317);
    layer2_outputs(7151) <= not(layer1_outputs(852));
    layer2_outputs(7152) <= (layer1_outputs(5797)) or (layer1_outputs(11520));
    layer2_outputs(7153) <= layer1_outputs(1485);
    layer2_outputs(7154) <= (layer1_outputs(8779)) and not (layer1_outputs(1220));
    layer2_outputs(7155) <= not(layer1_outputs(2497));
    layer2_outputs(7156) <= not((layer1_outputs(1413)) or (layer1_outputs(7910)));
    layer2_outputs(7157) <= not(layer1_outputs(714));
    layer2_outputs(7158) <= not(layer1_outputs(3406));
    layer2_outputs(7159) <= '1';
    layer2_outputs(7160) <= not(layer1_outputs(11977));
    layer2_outputs(7161) <= not(layer1_outputs(680)) or (layer1_outputs(7695));
    layer2_outputs(7162) <= not(layer1_outputs(7930));
    layer2_outputs(7163) <= (layer1_outputs(10202)) or (layer1_outputs(5678));
    layer2_outputs(7164) <= (layer1_outputs(3437)) xor (layer1_outputs(10291));
    layer2_outputs(7165) <= (layer1_outputs(5358)) xor (layer1_outputs(1196));
    layer2_outputs(7166) <= not((layer1_outputs(2889)) or (layer1_outputs(5994)));
    layer2_outputs(7167) <= not((layer1_outputs(915)) or (layer1_outputs(10952)));
    layer2_outputs(7168) <= not((layer1_outputs(11878)) xor (layer1_outputs(10612)));
    layer2_outputs(7169) <= not(layer1_outputs(8306)) or (layer1_outputs(4821));
    layer2_outputs(7170) <= layer1_outputs(9382);
    layer2_outputs(7171) <= (layer1_outputs(10943)) and not (layer1_outputs(10745));
    layer2_outputs(7172) <= not((layer1_outputs(8688)) or (layer1_outputs(1485)));
    layer2_outputs(7173) <= layer1_outputs(6902);
    layer2_outputs(7174) <= (layer1_outputs(10240)) xor (layer1_outputs(12224));
    layer2_outputs(7175) <= layer1_outputs(5743);
    layer2_outputs(7176) <= not((layer1_outputs(3333)) xor (layer1_outputs(730)));
    layer2_outputs(7177) <= layer1_outputs(10399);
    layer2_outputs(7178) <= not((layer1_outputs(2434)) or (layer1_outputs(608)));
    layer2_outputs(7179) <= '1';
    layer2_outputs(7180) <= layer1_outputs(746);
    layer2_outputs(7181) <= not(layer1_outputs(9082));
    layer2_outputs(7182) <= not((layer1_outputs(5556)) or (layer1_outputs(9250)));
    layer2_outputs(7183) <= layer1_outputs(837);
    layer2_outputs(7184) <= not(layer1_outputs(4823));
    layer2_outputs(7185) <= layer1_outputs(3118);
    layer2_outputs(7186) <= not((layer1_outputs(5747)) xor (layer1_outputs(2799)));
    layer2_outputs(7187) <= not(layer1_outputs(8263));
    layer2_outputs(7188) <= not(layer1_outputs(9897));
    layer2_outputs(7189) <= not(layer1_outputs(10409));
    layer2_outputs(7190) <= layer1_outputs(316);
    layer2_outputs(7191) <= not(layer1_outputs(8358));
    layer2_outputs(7192) <= not((layer1_outputs(1535)) and (layer1_outputs(10169)));
    layer2_outputs(7193) <= (layer1_outputs(3638)) and (layer1_outputs(4279));
    layer2_outputs(7194) <= (layer1_outputs(9338)) and not (layer1_outputs(1920));
    layer2_outputs(7195) <= layer1_outputs(10691);
    layer2_outputs(7196) <= (layer1_outputs(11118)) and not (layer1_outputs(11351));
    layer2_outputs(7197) <= not(layer1_outputs(120));
    layer2_outputs(7198) <= not(layer1_outputs(985)) or (layer1_outputs(2206));
    layer2_outputs(7199) <= not(layer1_outputs(12304));
    layer2_outputs(7200) <= not((layer1_outputs(2866)) xor (layer1_outputs(9853)));
    layer2_outputs(7201) <= layer1_outputs(586);
    layer2_outputs(7202) <= not(layer1_outputs(6317));
    layer2_outputs(7203) <= not(layer1_outputs(3245));
    layer2_outputs(7204) <= not(layer1_outputs(8962));
    layer2_outputs(7205) <= not(layer1_outputs(4242)) or (layer1_outputs(1104));
    layer2_outputs(7206) <= not((layer1_outputs(11829)) and (layer1_outputs(11793)));
    layer2_outputs(7207) <= not(layer1_outputs(12534));
    layer2_outputs(7208) <= not((layer1_outputs(2471)) and (layer1_outputs(5327)));
    layer2_outputs(7209) <= (layer1_outputs(10066)) and not (layer1_outputs(878));
    layer2_outputs(7210) <= not((layer1_outputs(3020)) or (layer1_outputs(12015)));
    layer2_outputs(7211) <= layer1_outputs(7420);
    layer2_outputs(7212) <= not(layer1_outputs(2089));
    layer2_outputs(7213) <= not((layer1_outputs(8955)) or (layer1_outputs(5505)));
    layer2_outputs(7214) <= (layer1_outputs(10757)) and (layer1_outputs(8550));
    layer2_outputs(7215) <= layer1_outputs(5900);
    layer2_outputs(7216) <= layer1_outputs(11311);
    layer2_outputs(7217) <= not(layer1_outputs(7758)) or (layer1_outputs(8106));
    layer2_outputs(7218) <= not((layer1_outputs(8710)) xor (layer1_outputs(4786)));
    layer2_outputs(7219) <= not((layer1_outputs(9917)) and (layer1_outputs(562)));
    layer2_outputs(7220) <= not(layer1_outputs(5097));
    layer2_outputs(7221) <= layer1_outputs(3208);
    layer2_outputs(7222) <= not(layer1_outputs(1457));
    layer2_outputs(7223) <= not(layer1_outputs(9203));
    layer2_outputs(7224) <= '1';
    layer2_outputs(7225) <= (layer1_outputs(8559)) xor (layer1_outputs(11884));
    layer2_outputs(7226) <= not(layer1_outputs(11212));
    layer2_outputs(7227) <= not((layer1_outputs(3701)) or (layer1_outputs(9725)));
    layer2_outputs(7228) <= (layer1_outputs(12740)) and not (layer1_outputs(2124));
    layer2_outputs(7229) <= not(layer1_outputs(3141)) or (layer1_outputs(3935));
    layer2_outputs(7230) <= layer1_outputs(2121);
    layer2_outputs(7231) <= layer1_outputs(5365);
    layer2_outputs(7232) <= not((layer1_outputs(1448)) xor (layer1_outputs(255)));
    layer2_outputs(7233) <= not((layer1_outputs(5336)) xor (layer1_outputs(1519)));
    layer2_outputs(7234) <= not(layer1_outputs(4835));
    layer2_outputs(7235) <= not(layer1_outputs(4659));
    layer2_outputs(7236) <= not(layer1_outputs(7407)) or (layer1_outputs(9362));
    layer2_outputs(7237) <= (layer1_outputs(2809)) xor (layer1_outputs(9877));
    layer2_outputs(7238) <= not((layer1_outputs(1238)) xor (layer1_outputs(10548)));
    layer2_outputs(7239) <= not(layer1_outputs(4082));
    layer2_outputs(7240) <= not(layer1_outputs(12437));
    layer2_outputs(7241) <= not(layer1_outputs(8552));
    layer2_outputs(7242) <= layer1_outputs(7492);
    layer2_outputs(7243) <= not(layer1_outputs(2858)) or (layer1_outputs(6171));
    layer2_outputs(7244) <= not(layer1_outputs(4772)) or (layer1_outputs(6180));
    layer2_outputs(7245) <= (layer1_outputs(5868)) and not (layer1_outputs(10134));
    layer2_outputs(7246) <= not(layer1_outputs(2480));
    layer2_outputs(7247) <= not(layer1_outputs(8977)) or (layer1_outputs(7096));
    layer2_outputs(7248) <= (layer1_outputs(11718)) and (layer1_outputs(7200));
    layer2_outputs(7249) <= not((layer1_outputs(8569)) or (layer1_outputs(5913)));
    layer2_outputs(7250) <= (layer1_outputs(3269)) and not (layer1_outputs(6955));
    layer2_outputs(7251) <= not((layer1_outputs(5003)) xor (layer1_outputs(417)));
    layer2_outputs(7252) <= not(layer1_outputs(11978)) or (layer1_outputs(12299));
    layer2_outputs(7253) <= not(layer1_outputs(6338));
    layer2_outputs(7254) <= not(layer1_outputs(1471));
    layer2_outputs(7255) <= layer1_outputs(7732);
    layer2_outputs(7256) <= not(layer1_outputs(1306));
    layer2_outputs(7257) <= not((layer1_outputs(2759)) xor (layer1_outputs(1477)));
    layer2_outputs(7258) <= not((layer1_outputs(2114)) and (layer1_outputs(9796)));
    layer2_outputs(7259) <= layer1_outputs(7514);
    layer2_outputs(7260) <= layer1_outputs(7244);
    layer2_outputs(7261) <= not(layer1_outputs(11134));
    layer2_outputs(7262) <= layer1_outputs(9468);
    layer2_outputs(7263) <= layer1_outputs(9184);
    layer2_outputs(7264) <= layer1_outputs(882);
    layer2_outputs(7265) <= layer1_outputs(8236);
    layer2_outputs(7266) <= not((layer1_outputs(2379)) xor (layer1_outputs(4683)));
    layer2_outputs(7267) <= not(layer1_outputs(4071));
    layer2_outputs(7268) <= (layer1_outputs(2398)) xor (layer1_outputs(505));
    layer2_outputs(7269) <= (layer1_outputs(3200)) or (layer1_outputs(12615));
    layer2_outputs(7270) <= not((layer1_outputs(2353)) xor (layer1_outputs(2000)));
    layer2_outputs(7271) <= (layer1_outputs(5723)) and (layer1_outputs(2577));
    layer2_outputs(7272) <= not((layer1_outputs(1462)) xor (layer1_outputs(5034)));
    layer2_outputs(7273) <= layer1_outputs(245);
    layer2_outputs(7274) <= layer1_outputs(8097);
    layer2_outputs(7275) <= (layer1_outputs(832)) xor (layer1_outputs(609));
    layer2_outputs(7276) <= not(layer1_outputs(8964)) or (layer1_outputs(2708));
    layer2_outputs(7277) <= (layer1_outputs(3664)) and not (layer1_outputs(2433));
    layer2_outputs(7278) <= layer1_outputs(7929);
    layer2_outputs(7279) <= not(layer1_outputs(3645));
    layer2_outputs(7280) <= layer1_outputs(6950);
    layer2_outputs(7281) <= layer1_outputs(10555);
    layer2_outputs(7282) <= not(layer1_outputs(12767));
    layer2_outputs(7283) <= not(layer1_outputs(6249)) or (layer1_outputs(7406));
    layer2_outputs(7284) <= (layer1_outputs(6349)) and not (layer1_outputs(8810));
    layer2_outputs(7285) <= not(layer1_outputs(3393));
    layer2_outputs(7286) <= not(layer1_outputs(4715));
    layer2_outputs(7287) <= (layer1_outputs(2348)) xor (layer1_outputs(12422));
    layer2_outputs(7288) <= not((layer1_outputs(12265)) xor (layer1_outputs(9387)));
    layer2_outputs(7289) <= not((layer1_outputs(11494)) or (layer1_outputs(6407)));
    layer2_outputs(7290) <= (layer1_outputs(9044)) and not (layer1_outputs(8773));
    layer2_outputs(7291) <= not(layer1_outputs(7061));
    layer2_outputs(7292) <= not((layer1_outputs(12071)) xor (layer1_outputs(11231)));
    layer2_outputs(7293) <= not(layer1_outputs(1792));
    layer2_outputs(7294) <= not(layer1_outputs(6791));
    layer2_outputs(7295) <= (layer1_outputs(3040)) and not (layer1_outputs(8527));
    layer2_outputs(7296) <= layer1_outputs(861);
    layer2_outputs(7297) <= not(layer1_outputs(9988));
    layer2_outputs(7298) <= (layer1_outputs(11707)) and (layer1_outputs(11688));
    layer2_outputs(7299) <= (layer1_outputs(10396)) and not (layer1_outputs(6579));
    layer2_outputs(7300) <= not(layer1_outputs(3307));
    layer2_outputs(7301) <= not(layer1_outputs(9459));
    layer2_outputs(7302) <= layer1_outputs(4100);
    layer2_outputs(7303) <= (layer1_outputs(10685)) and not (layer1_outputs(2006));
    layer2_outputs(7304) <= (layer1_outputs(7491)) or (layer1_outputs(4476));
    layer2_outputs(7305) <= layer1_outputs(4691);
    layer2_outputs(7306) <= (layer1_outputs(6522)) xor (layer1_outputs(11783));
    layer2_outputs(7307) <= layer1_outputs(6717);
    layer2_outputs(7308) <= not(layer1_outputs(3812));
    layer2_outputs(7309) <= not(layer1_outputs(8615));
    layer2_outputs(7310) <= (layer1_outputs(4395)) or (layer1_outputs(11848));
    layer2_outputs(7311) <= '0';
    layer2_outputs(7312) <= '0';
    layer2_outputs(7313) <= not(layer1_outputs(12759));
    layer2_outputs(7314) <= layer1_outputs(4999);
    layer2_outputs(7315) <= (layer1_outputs(3871)) or (layer1_outputs(10191));
    layer2_outputs(7316) <= not(layer1_outputs(9207));
    layer2_outputs(7317) <= layer1_outputs(4517);
    layer2_outputs(7318) <= not(layer1_outputs(11133)) or (layer1_outputs(9814));
    layer2_outputs(7319) <= layer1_outputs(12575);
    layer2_outputs(7320) <= (layer1_outputs(2445)) and (layer1_outputs(11756));
    layer2_outputs(7321) <= (layer1_outputs(12638)) or (layer1_outputs(466));
    layer2_outputs(7322) <= '0';
    layer2_outputs(7323) <= not(layer1_outputs(1976));
    layer2_outputs(7324) <= (layer1_outputs(12684)) xor (layer1_outputs(11235));
    layer2_outputs(7325) <= not(layer1_outputs(4291));
    layer2_outputs(7326) <= not((layer1_outputs(5504)) or (layer1_outputs(10344)));
    layer2_outputs(7327) <= (layer1_outputs(11802)) and not (layer1_outputs(7649));
    layer2_outputs(7328) <= not(layer1_outputs(2285));
    layer2_outputs(7329) <= not(layer1_outputs(2741));
    layer2_outputs(7330) <= layer1_outputs(8972);
    layer2_outputs(7331) <= not(layer1_outputs(797));
    layer2_outputs(7332) <= '0';
    layer2_outputs(7333) <= not(layer1_outputs(10725));
    layer2_outputs(7334) <= not(layer1_outputs(9172));
    layer2_outputs(7335) <= not(layer1_outputs(10719));
    layer2_outputs(7336) <= (layer1_outputs(5593)) and not (layer1_outputs(11221));
    layer2_outputs(7337) <= not((layer1_outputs(4042)) xor (layer1_outputs(10282)));
    layer2_outputs(7338) <= not(layer1_outputs(11441));
    layer2_outputs(7339) <= not(layer1_outputs(11473));
    layer2_outputs(7340) <= (layer1_outputs(7956)) xor (layer1_outputs(7195));
    layer2_outputs(7341) <= not(layer1_outputs(1329));
    layer2_outputs(7342) <= '1';
    layer2_outputs(7343) <= not((layer1_outputs(8059)) xor (layer1_outputs(12457)));
    layer2_outputs(7344) <= not(layer1_outputs(11360));
    layer2_outputs(7345) <= not(layer1_outputs(6877));
    layer2_outputs(7346) <= not(layer1_outputs(11773));
    layer2_outputs(7347) <= not(layer1_outputs(12772));
    layer2_outputs(7348) <= (layer1_outputs(1522)) xor (layer1_outputs(6623));
    layer2_outputs(7349) <= layer1_outputs(5220);
    layer2_outputs(7350) <= not(layer1_outputs(6044));
    layer2_outputs(7351) <= (layer1_outputs(8161)) xor (layer1_outputs(8660));
    layer2_outputs(7352) <= not((layer1_outputs(976)) and (layer1_outputs(2436)));
    layer2_outputs(7353) <= not(layer1_outputs(3492));
    layer2_outputs(7354) <= not(layer1_outputs(760)) or (layer1_outputs(1957));
    layer2_outputs(7355) <= (layer1_outputs(10425)) and not (layer1_outputs(2228));
    layer2_outputs(7356) <= not(layer1_outputs(7534));
    layer2_outputs(7357) <= layer1_outputs(954);
    layer2_outputs(7358) <= layer1_outputs(2771);
    layer2_outputs(7359) <= not(layer1_outputs(4649));
    layer2_outputs(7360) <= layer1_outputs(9094);
    layer2_outputs(7361) <= (layer1_outputs(6628)) xor (layer1_outputs(12089));
    layer2_outputs(7362) <= (layer1_outputs(4765)) xor (layer1_outputs(11904));
    layer2_outputs(7363) <= layer1_outputs(9455);
    layer2_outputs(7364) <= not(layer1_outputs(1810)) or (layer1_outputs(5080));
    layer2_outputs(7365) <= not(layer1_outputs(1134));
    layer2_outputs(7366) <= (layer1_outputs(11697)) or (layer1_outputs(9047));
    layer2_outputs(7367) <= not(layer1_outputs(8888));
    layer2_outputs(7368) <= layer1_outputs(7811);
    layer2_outputs(7369) <= not(layer1_outputs(8625));
    layer2_outputs(7370) <= layer1_outputs(618);
    layer2_outputs(7371) <= not(layer1_outputs(8254)) or (layer1_outputs(7263));
    layer2_outputs(7372) <= not(layer1_outputs(2926));
    layer2_outputs(7373) <= (layer1_outputs(2075)) xor (layer1_outputs(5741));
    layer2_outputs(7374) <= not(layer1_outputs(6419));
    layer2_outputs(7375) <= not(layer1_outputs(8821)) or (layer1_outputs(2115));
    layer2_outputs(7376) <= layer1_outputs(4908);
    layer2_outputs(7377) <= layer1_outputs(4553);
    layer2_outputs(7378) <= (layer1_outputs(1368)) xor (layer1_outputs(8715));
    layer2_outputs(7379) <= not(layer1_outputs(2920)) or (layer1_outputs(6462));
    layer2_outputs(7380) <= layer1_outputs(7941);
    layer2_outputs(7381) <= layer1_outputs(1888);
    layer2_outputs(7382) <= layer1_outputs(7961);
    layer2_outputs(7383) <= not(layer1_outputs(5559)) or (layer1_outputs(6127));
    layer2_outputs(7384) <= (layer1_outputs(2870)) and (layer1_outputs(10784));
    layer2_outputs(7385) <= not((layer1_outputs(9746)) or (layer1_outputs(12550)));
    layer2_outputs(7386) <= not((layer1_outputs(4358)) xor (layer1_outputs(1885)));
    layer2_outputs(7387) <= (layer1_outputs(1504)) and not (layer1_outputs(5349));
    layer2_outputs(7388) <= not((layer1_outputs(6694)) xor (layer1_outputs(7898)));
    layer2_outputs(7389) <= not((layer1_outputs(5836)) or (layer1_outputs(1432)));
    layer2_outputs(7390) <= not(layer1_outputs(438));
    layer2_outputs(7391) <= (layer1_outputs(501)) and not (layer1_outputs(1458));
    layer2_outputs(7392) <= not((layer1_outputs(5876)) xor (layer1_outputs(9103)));
    layer2_outputs(7393) <= not(layer1_outputs(8458)) or (layer1_outputs(739));
    layer2_outputs(7394) <= (layer1_outputs(3407)) or (layer1_outputs(2286));
    layer2_outputs(7395) <= (layer1_outputs(3563)) and not (layer1_outputs(4641));
    layer2_outputs(7396) <= layer1_outputs(7860);
    layer2_outputs(7397) <= not((layer1_outputs(2807)) or (layer1_outputs(12457)));
    layer2_outputs(7398) <= not(layer1_outputs(6703));
    layer2_outputs(7399) <= not((layer1_outputs(12563)) or (layer1_outputs(5945)));
    layer2_outputs(7400) <= not(layer1_outputs(12255));
    layer2_outputs(7401) <= not((layer1_outputs(6642)) and (layer1_outputs(3529)));
    layer2_outputs(7402) <= (layer1_outputs(10061)) xor (layer1_outputs(2902));
    layer2_outputs(7403) <= (layer1_outputs(3081)) and not (layer1_outputs(11328));
    layer2_outputs(7404) <= not(layer1_outputs(6179)) or (layer1_outputs(10553));
    layer2_outputs(7405) <= layer1_outputs(9506);
    layer2_outputs(7406) <= (layer1_outputs(4268)) xor (layer1_outputs(150));
    layer2_outputs(7407) <= layer1_outputs(11043);
    layer2_outputs(7408) <= layer1_outputs(12229);
    layer2_outputs(7409) <= layer1_outputs(3646);
    layer2_outputs(7410) <= not(layer1_outputs(8492));
    layer2_outputs(7411) <= (layer1_outputs(11536)) xor (layer1_outputs(7984));
    layer2_outputs(7412) <= not((layer1_outputs(8272)) xor (layer1_outputs(3301)));
    layer2_outputs(7413) <= layer1_outputs(1649);
    layer2_outputs(7414) <= not(layer1_outputs(9745));
    layer2_outputs(7415) <= not(layer1_outputs(9888));
    layer2_outputs(7416) <= not(layer1_outputs(5528));
    layer2_outputs(7417) <= layer1_outputs(6771);
    layer2_outputs(7418) <= not((layer1_outputs(1447)) or (layer1_outputs(7424)));
    layer2_outputs(7419) <= not(layer1_outputs(5767));
    layer2_outputs(7420) <= not(layer1_outputs(11722)) or (layer1_outputs(12162));
    layer2_outputs(7421) <= not(layer1_outputs(4912));
    layer2_outputs(7422) <= layer1_outputs(2810);
    layer2_outputs(7423) <= (layer1_outputs(2218)) and (layer1_outputs(6950));
    layer2_outputs(7424) <= not((layer1_outputs(12426)) and (layer1_outputs(9617)));
    layer2_outputs(7425) <= (layer1_outputs(10317)) and not (layer1_outputs(2535));
    layer2_outputs(7426) <= layer1_outputs(11733);
    layer2_outputs(7427) <= layer1_outputs(79);
    layer2_outputs(7428) <= '0';
    layer2_outputs(7429) <= (layer1_outputs(5426)) or (layer1_outputs(10203));
    layer2_outputs(7430) <= not(layer1_outputs(381)) or (layer1_outputs(8781));
    layer2_outputs(7431) <= not(layer1_outputs(7776));
    layer2_outputs(7432) <= not((layer1_outputs(10430)) xor (layer1_outputs(9518)));
    layer2_outputs(7433) <= not((layer1_outputs(5700)) and (layer1_outputs(3559)));
    layer2_outputs(7434) <= (layer1_outputs(5853)) and not (layer1_outputs(8746));
    layer2_outputs(7435) <= layer1_outputs(421);
    layer2_outputs(7436) <= not((layer1_outputs(3768)) xor (layer1_outputs(7262)));
    layer2_outputs(7437) <= not((layer1_outputs(7476)) xor (layer1_outputs(3467)));
    layer2_outputs(7438) <= not(layer1_outputs(10372));
    layer2_outputs(7439) <= not(layer1_outputs(10305));
    layer2_outputs(7440) <= layer1_outputs(12170);
    layer2_outputs(7441) <= not((layer1_outputs(3396)) xor (layer1_outputs(2172)));
    layer2_outputs(7442) <= not(layer1_outputs(8623));
    layer2_outputs(7443) <= not(layer1_outputs(12193));
    layer2_outputs(7444) <= (layer1_outputs(11838)) xor (layer1_outputs(11039));
    layer2_outputs(7445) <= layer1_outputs(240);
    layer2_outputs(7446) <= (layer1_outputs(7785)) xor (layer1_outputs(5825));
    layer2_outputs(7447) <= (layer1_outputs(10216)) xor (layer1_outputs(5175));
    layer2_outputs(7448) <= not((layer1_outputs(7692)) xor (layer1_outputs(7794)));
    layer2_outputs(7449) <= not(layer1_outputs(11230)) or (layer1_outputs(4237));
    layer2_outputs(7450) <= not((layer1_outputs(9806)) xor (layer1_outputs(7068)));
    layer2_outputs(7451) <= not(layer1_outputs(3793));
    layer2_outputs(7452) <= not(layer1_outputs(8000)) or (layer1_outputs(1901));
    layer2_outputs(7453) <= layer1_outputs(7781);
    layer2_outputs(7454) <= not(layer1_outputs(9248));
    layer2_outputs(7455) <= not(layer1_outputs(3429));
    layer2_outputs(7456) <= not((layer1_outputs(8345)) and (layer1_outputs(4574)));
    layer2_outputs(7457) <= (layer1_outputs(2071)) xor (layer1_outputs(11727));
    layer2_outputs(7458) <= layer1_outputs(9136);
    layer2_outputs(7459) <= not(layer1_outputs(4657));
    layer2_outputs(7460) <= (layer1_outputs(4679)) or (layer1_outputs(6843));
    layer2_outputs(7461) <= not((layer1_outputs(3618)) and (layer1_outputs(7016)));
    layer2_outputs(7462) <= not(layer1_outputs(5937)) or (layer1_outputs(5352));
    layer2_outputs(7463) <= not(layer1_outputs(5362)) or (layer1_outputs(11976));
    layer2_outputs(7464) <= layer1_outputs(12164);
    layer2_outputs(7465) <= (layer1_outputs(2023)) xor (layer1_outputs(9167));
    layer2_outputs(7466) <= not(layer1_outputs(2521));
    layer2_outputs(7467) <= layer1_outputs(572);
    layer2_outputs(7468) <= (layer1_outputs(1612)) xor (layer1_outputs(838));
    layer2_outputs(7469) <= not(layer1_outputs(7489)) or (layer1_outputs(8812));
    layer2_outputs(7470) <= layer1_outputs(6452);
    layer2_outputs(7471) <= (layer1_outputs(7719)) xor (layer1_outputs(8199));
    layer2_outputs(7472) <= (layer1_outputs(12483)) xor (layer1_outputs(8114));
    layer2_outputs(7473) <= layer1_outputs(5291);
    layer2_outputs(7474) <= layer1_outputs(1428);
    layer2_outputs(7475) <= not(layer1_outputs(10318));
    layer2_outputs(7476) <= not(layer1_outputs(2617));
    layer2_outputs(7477) <= '0';
    layer2_outputs(7478) <= not(layer1_outputs(6908));
    layer2_outputs(7479) <= not((layer1_outputs(4738)) xor (layer1_outputs(8360)));
    layer2_outputs(7480) <= layer1_outputs(3347);
    layer2_outputs(7481) <= not(layer1_outputs(8690));
    layer2_outputs(7482) <= (layer1_outputs(7276)) xor (layer1_outputs(5883));
    layer2_outputs(7483) <= layer1_outputs(8393);
    layer2_outputs(7484) <= (layer1_outputs(7042)) xor (layer1_outputs(7028));
    layer2_outputs(7485) <= (layer1_outputs(7564)) and not (layer1_outputs(4902));
    layer2_outputs(7486) <= not(layer1_outputs(1124));
    layer2_outputs(7487) <= not(layer1_outputs(2957)) or (layer1_outputs(11897));
    layer2_outputs(7488) <= '0';
    layer2_outputs(7489) <= (layer1_outputs(8633)) and (layer1_outputs(12039));
    layer2_outputs(7490) <= not(layer1_outputs(3786)) or (layer1_outputs(7748));
    layer2_outputs(7491) <= not(layer1_outputs(6643));
    layer2_outputs(7492) <= (layer1_outputs(7188)) and not (layer1_outputs(4436));
    layer2_outputs(7493) <= not((layer1_outputs(5334)) xor (layer1_outputs(9221)));
    layer2_outputs(7494) <= not(layer1_outputs(9194)) or (layer1_outputs(11683));
    layer2_outputs(7495) <= (layer1_outputs(11070)) and not (layer1_outputs(9432));
    layer2_outputs(7496) <= layer1_outputs(2732);
    layer2_outputs(7497) <= not(layer1_outputs(6025));
    layer2_outputs(7498) <= layer1_outputs(5187);
    layer2_outputs(7499) <= layer1_outputs(4977);
    layer2_outputs(7500) <= not(layer1_outputs(160));
    layer2_outputs(7501) <= (layer1_outputs(12005)) and not (layer1_outputs(3759));
    layer2_outputs(7502) <= layer1_outputs(434);
    layer2_outputs(7503) <= not(layer1_outputs(7254));
    layer2_outputs(7504) <= layer1_outputs(624);
    layer2_outputs(7505) <= layer1_outputs(4341);
    layer2_outputs(7506) <= not(layer1_outputs(2263)) or (layer1_outputs(8124));
    layer2_outputs(7507) <= layer1_outputs(3240);
    layer2_outputs(7508) <= not(layer1_outputs(3426));
    layer2_outputs(7509) <= (layer1_outputs(5837)) xor (layer1_outputs(1925));
    layer2_outputs(7510) <= not((layer1_outputs(4952)) xor (layer1_outputs(11817)));
    layer2_outputs(7511) <= not((layer1_outputs(10390)) xor (layer1_outputs(6324)));
    layer2_outputs(7512) <= (layer1_outputs(980)) xor (layer1_outputs(5746));
    layer2_outputs(7513) <= not(layer1_outputs(8496)) or (layer1_outputs(7954));
    layer2_outputs(7514) <= (layer1_outputs(9353)) and (layer1_outputs(10643));
    layer2_outputs(7515) <= not(layer1_outputs(8773));
    layer2_outputs(7516) <= not(layer1_outputs(7731));
    layer2_outputs(7517) <= (layer1_outputs(2284)) and (layer1_outputs(10370));
    layer2_outputs(7518) <= (layer1_outputs(7593)) and not (layer1_outputs(2269));
    layer2_outputs(7519) <= not(layer1_outputs(2558));
    layer2_outputs(7520) <= layer1_outputs(2301);
    layer2_outputs(7521) <= (layer1_outputs(6707)) and (layer1_outputs(12671));
    layer2_outputs(7522) <= not(layer1_outputs(868));
    layer2_outputs(7523) <= (layer1_outputs(5041)) and not (layer1_outputs(2834));
    layer2_outputs(7524) <= not(layer1_outputs(843));
    layer2_outputs(7525) <= layer1_outputs(6497);
    layer2_outputs(7526) <= (layer1_outputs(492)) xor (layer1_outputs(11196));
    layer2_outputs(7527) <= not(layer1_outputs(1227));
    layer2_outputs(7528) <= (layer1_outputs(664)) and (layer1_outputs(755));
    layer2_outputs(7529) <= not(layer1_outputs(6644));
    layer2_outputs(7530) <= layer1_outputs(12134);
    layer2_outputs(7531) <= not(layer1_outputs(9999)) or (layer1_outputs(9639));
    layer2_outputs(7532) <= (layer1_outputs(5057)) xor (layer1_outputs(8362));
    layer2_outputs(7533) <= not(layer1_outputs(12766));
    layer2_outputs(7534) <= layer1_outputs(12127);
    layer2_outputs(7535) <= not(layer1_outputs(7821)) or (layer1_outputs(11082));
    layer2_outputs(7536) <= (layer1_outputs(8200)) or (layer1_outputs(3317));
    layer2_outputs(7537) <= not(layer1_outputs(1218));
    layer2_outputs(7538) <= layer1_outputs(1167);
    layer2_outputs(7539) <= (layer1_outputs(3901)) and not (layer1_outputs(10182));
    layer2_outputs(7540) <= (layer1_outputs(5771)) and (layer1_outputs(6183));
    layer2_outputs(7541) <= (layer1_outputs(404)) and not (layer1_outputs(7520));
    layer2_outputs(7542) <= (layer1_outputs(9782)) or (layer1_outputs(10617));
    layer2_outputs(7543) <= not(layer1_outputs(12485));
    layer2_outputs(7544) <= not((layer1_outputs(1086)) xor (layer1_outputs(8002)));
    layer2_outputs(7545) <= (layer1_outputs(2751)) xor (layer1_outputs(12006));
    layer2_outputs(7546) <= layer1_outputs(9437);
    layer2_outputs(7547) <= layer1_outputs(2095);
    layer2_outputs(7548) <= not(layer1_outputs(12777));
    layer2_outputs(7549) <= layer1_outputs(2656);
    layer2_outputs(7550) <= (layer1_outputs(3679)) and not (layer1_outputs(6288));
    layer2_outputs(7551) <= not(layer1_outputs(11630));
    layer2_outputs(7552) <= not(layer1_outputs(1052));
    layer2_outputs(7553) <= not(layer1_outputs(12451));
    layer2_outputs(7554) <= not(layer1_outputs(11945));
    layer2_outputs(7555) <= (layer1_outputs(4423)) and not (layer1_outputs(4907));
    layer2_outputs(7556) <= not(layer1_outputs(7705)) or (layer1_outputs(12196));
    layer2_outputs(7557) <= layer1_outputs(7510);
    layer2_outputs(7558) <= not((layer1_outputs(6670)) or (layer1_outputs(5325)));
    layer2_outputs(7559) <= not((layer1_outputs(11411)) or (layer1_outputs(8403)));
    layer2_outputs(7560) <= layer1_outputs(11013);
    layer2_outputs(7561) <= layer1_outputs(10373);
    layer2_outputs(7562) <= (layer1_outputs(8172)) and (layer1_outputs(5491));
    layer2_outputs(7563) <= layer1_outputs(4304);
    layer2_outputs(7564) <= (layer1_outputs(1895)) and not (layer1_outputs(8882));
    layer2_outputs(7565) <= not(layer1_outputs(6009));
    layer2_outputs(7566) <= not(layer1_outputs(10611)) or (layer1_outputs(3269));
    layer2_outputs(7567) <= (layer1_outputs(2213)) and not (layer1_outputs(9490));
    layer2_outputs(7568) <= layer1_outputs(5745);
    layer2_outputs(7569) <= not(layer1_outputs(4522)) or (layer1_outputs(4110));
    layer2_outputs(7570) <= not(layer1_outputs(8079)) or (layer1_outputs(850));
    layer2_outputs(7571) <= not(layer1_outputs(5975));
    layer2_outputs(7572) <= not(layer1_outputs(3749)) or (layer1_outputs(576));
    layer2_outputs(7573) <= not((layer1_outputs(11818)) and (layer1_outputs(2941)));
    layer2_outputs(7574) <= layer1_outputs(4709);
    layer2_outputs(7575) <= layer1_outputs(2975);
    layer2_outputs(7576) <= (layer1_outputs(5675)) or (layer1_outputs(7082));
    layer2_outputs(7577) <= (layer1_outputs(999)) and (layer1_outputs(8988));
    layer2_outputs(7578) <= (layer1_outputs(4487)) or (layer1_outputs(9865));
    layer2_outputs(7579) <= (layer1_outputs(1126)) or (layer1_outputs(2420));
    layer2_outputs(7580) <= layer1_outputs(12724);
    layer2_outputs(7581) <= not(layer1_outputs(11664)) or (layer1_outputs(4559));
    layer2_outputs(7582) <= layer1_outputs(10235);
    layer2_outputs(7583) <= not(layer1_outputs(3682));
    layer2_outputs(7584) <= not(layer1_outputs(2777));
    layer2_outputs(7585) <= layer1_outputs(3852);
    layer2_outputs(7586) <= not((layer1_outputs(2524)) xor (layer1_outputs(5641)));
    layer2_outputs(7587) <= (layer1_outputs(7026)) and (layer1_outputs(6996));
    layer2_outputs(7588) <= (layer1_outputs(629)) and (layer1_outputs(2890));
    layer2_outputs(7589) <= not(layer1_outputs(12776)) or (layer1_outputs(8633));
    layer2_outputs(7590) <= layer1_outputs(2852);
    layer2_outputs(7591) <= '0';
    layer2_outputs(7592) <= not(layer1_outputs(5536)) or (layer1_outputs(10980));
    layer2_outputs(7593) <= not(layer1_outputs(3611));
    layer2_outputs(7594) <= not((layer1_outputs(12050)) xor (layer1_outputs(11527)));
    layer2_outputs(7595) <= not(layer1_outputs(4213));
    layer2_outputs(7596) <= not((layer1_outputs(2019)) xor (layer1_outputs(3430)));
    layer2_outputs(7597) <= not(layer1_outputs(2850)) or (layer1_outputs(4784));
    layer2_outputs(7598) <= layer1_outputs(7349);
    layer2_outputs(7599) <= not((layer1_outputs(7670)) xor (layer1_outputs(5053)));
    layer2_outputs(7600) <= layer1_outputs(6695);
    layer2_outputs(7601) <= (layer1_outputs(3094)) and (layer1_outputs(4116));
    layer2_outputs(7602) <= not(layer1_outputs(11668));
    layer2_outputs(7603) <= not((layer1_outputs(12236)) or (layer1_outputs(11798)));
    layer2_outputs(7604) <= layer1_outputs(9165);
    layer2_outputs(7605) <= not(layer1_outputs(10180));
    layer2_outputs(7606) <= layer1_outputs(698);
    layer2_outputs(7607) <= not(layer1_outputs(7730)) or (layer1_outputs(8348));
    layer2_outputs(7608) <= (layer1_outputs(8979)) and (layer1_outputs(4790));
    layer2_outputs(7609) <= not((layer1_outputs(2140)) and (layer1_outputs(1371)));
    layer2_outputs(7610) <= (layer1_outputs(2472)) or (layer1_outputs(99));
    layer2_outputs(7611) <= layer1_outputs(7812);
    layer2_outputs(7612) <= (layer1_outputs(5950)) and not (layer1_outputs(1620));
    layer2_outputs(7613) <= not(layer1_outputs(5661));
    layer2_outputs(7614) <= not(layer1_outputs(2965));
    layer2_outputs(7615) <= not(layer1_outputs(5921));
    layer2_outputs(7616) <= not((layer1_outputs(7002)) and (layer1_outputs(7613)));
    layer2_outputs(7617) <= layer1_outputs(2676);
    layer2_outputs(7618) <= not((layer1_outputs(1696)) and (layer1_outputs(4309)));
    layer2_outputs(7619) <= layer1_outputs(257);
    layer2_outputs(7620) <= not((layer1_outputs(12676)) xor (layer1_outputs(491)));
    layer2_outputs(7621) <= not((layer1_outputs(11458)) or (layer1_outputs(7094)));
    layer2_outputs(7622) <= not((layer1_outputs(9388)) and (layer1_outputs(5956)));
    layer2_outputs(7623) <= not(layer1_outputs(3578));
    layer2_outputs(7624) <= not(layer1_outputs(11127));
    layer2_outputs(7625) <= not((layer1_outputs(7898)) or (layer1_outputs(6170)));
    layer2_outputs(7626) <= not((layer1_outputs(4617)) xor (layer1_outputs(2318)));
    layer2_outputs(7627) <= layer1_outputs(2897);
    layer2_outputs(7628) <= layer1_outputs(9264);
    layer2_outputs(7629) <= not((layer1_outputs(6012)) and (layer1_outputs(7638)));
    layer2_outputs(7630) <= not((layer1_outputs(6585)) xor (layer1_outputs(3587)));
    layer2_outputs(7631) <= (layer1_outputs(9242)) xor (layer1_outputs(7924));
    layer2_outputs(7632) <= (layer1_outputs(4262)) and not (layer1_outputs(123));
    layer2_outputs(7633) <= not(layer1_outputs(4283)) or (layer1_outputs(6821));
    layer2_outputs(7634) <= not(layer1_outputs(3866));
    layer2_outputs(7635) <= not(layer1_outputs(9685));
    layer2_outputs(7636) <= not(layer1_outputs(9256));
    layer2_outputs(7637) <= not(layer1_outputs(2690)) or (layer1_outputs(5573));
    layer2_outputs(7638) <= (layer1_outputs(3212)) xor (layer1_outputs(2512));
    layer2_outputs(7639) <= not(layer1_outputs(8723));
    layer2_outputs(7640) <= not((layer1_outputs(2847)) and (layer1_outputs(7478)));
    layer2_outputs(7641) <= layer1_outputs(5130);
    layer2_outputs(7642) <= not(layer1_outputs(922));
    layer2_outputs(7643) <= layer1_outputs(12424);
    layer2_outputs(7644) <= not((layer1_outputs(11860)) xor (layer1_outputs(1910)));
    layer2_outputs(7645) <= (layer1_outputs(10897)) and not (layer1_outputs(8031));
    layer2_outputs(7646) <= not(layer1_outputs(242));
    layer2_outputs(7647) <= (layer1_outputs(9941)) and (layer1_outputs(9518));
    layer2_outputs(7648) <= layer1_outputs(4751);
    layer2_outputs(7649) <= not((layer1_outputs(1191)) and (layer1_outputs(1704)));
    layer2_outputs(7650) <= layer1_outputs(6613);
    layer2_outputs(7651) <= not((layer1_outputs(5706)) xor (layer1_outputs(3128)));
    layer2_outputs(7652) <= layer1_outputs(8422);
    layer2_outputs(7653) <= (layer1_outputs(2204)) and not (layer1_outputs(6628));
    layer2_outputs(7654) <= not((layer1_outputs(5271)) xor (layer1_outputs(2887)));
    layer2_outputs(7655) <= not((layer1_outputs(7925)) xor (layer1_outputs(5628)));
    layer2_outputs(7656) <= layer1_outputs(6415);
    layer2_outputs(7657) <= not((layer1_outputs(6681)) xor (layer1_outputs(1869)));
    layer2_outputs(7658) <= not(layer1_outputs(7527));
    layer2_outputs(7659) <= not(layer1_outputs(8415));
    layer2_outputs(7660) <= not((layer1_outputs(7646)) or (layer1_outputs(6120)));
    layer2_outputs(7661) <= layer1_outputs(2439);
    layer2_outputs(7662) <= layer1_outputs(11070);
    layer2_outputs(7663) <= not(layer1_outputs(6370));
    layer2_outputs(7664) <= not(layer1_outputs(6673));
    layer2_outputs(7665) <= (layer1_outputs(424)) xor (layer1_outputs(3636));
    layer2_outputs(7666) <= (layer1_outputs(10400)) and not (layer1_outputs(8766));
    layer2_outputs(7667) <= layer1_outputs(4909);
    layer2_outputs(7668) <= not(layer1_outputs(4168));
    layer2_outputs(7669) <= layer1_outputs(787);
    layer2_outputs(7670) <= not(layer1_outputs(1077));
    layer2_outputs(7671) <= (layer1_outputs(4662)) and not (layer1_outputs(3948));
    layer2_outputs(7672) <= layer1_outputs(6137);
    layer2_outputs(7673) <= not((layer1_outputs(2953)) xor (layer1_outputs(12584)));
    layer2_outputs(7674) <= layer1_outputs(1700);
    layer2_outputs(7675) <= not(layer1_outputs(4641));
    layer2_outputs(7676) <= (layer1_outputs(3538)) and (layer1_outputs(6886));
    layer2_outputs(7677) <= layer1_outputs(2108);
    layer2_outputs(7678) <= not(layer1_outputs(3835));
    layer2_outputs(7679) <= '1';
    layer2_outputs(7680) <= not((layer1_outputs(12175)) and (layer1_outputs(180)));
    layer2_outputs(7681) <= layer1_outputs(9545);
    layer2_outputs(7682) <= not(layer1_outputs(11479)) or (layer1_outputs(8846));
    layer2_outputs(7683) <= not(layer1_outputs(9805));
    layer2_outputs(7684) <= layer1_outputs(10717);
    layer2_outputs(7685) <= (layer1_outputs(11622)) and (layer1_outputs(7797));
    layer2_outputs(7686) <= layer1_outputs(137);
    layer2_outputs(7687) <= not((layer1_outputs(6726)) xor (layer1_outputs(2934)));
    layer2_outputs(7688) <= (layer1_outputs(455)) and not (layer1_outputs(7868));
    layer2_outputs(7689) <= not((layer1_outputs(6053)) xor (layer1_outputs(4869)));
    layer2_outputs(7690) <= (layer1_outputs(7113)) or (layer1_outputs(5693));
    layer2_outputs(7691) <= not((layer1_outputs(12552)) xor (layer1_outputs(5118)));
    layer2_outputs(7692) <= (layer1_outputs(2698)) xor (layer1_outputs(11823));
    layer2_outputs(7693) <= not(layer1_outputs(2384));
    layer2_outputs(7694) <= not(layer1_outputs(4504));
    layer2_outputs(7695) <= layer1_outputs(9034);
    layer2_outputs(7696) <= not(layer1_outputs(3087)) or (layer1_outputs(4067));
    layer2_outputs(7697) <= (layer1_outputs(32)) or (layer1_outputs(196));
    layer2_outputs(7698) <= layer1_outputs(5897);
    layer2_outputs(7699) <= (layer1_outputs(6738)) xor (layer1_outputs(11103));
    layer2_outputs(7700) <= (layer1_outputs(4336)) and (layer1_outputs(10422));
    layer2_outputs(7701) <= not(layer1_outputs(7975)) or (layer1_outputs(7441));
    layer2_outputs(7702) <= not(layer1_outputs(5410)) or (layer1_outputs(10701));
    layer2_outputs(7703) <= (layer1_outputs(7496)) and not (layer1_outputs(10451));
    layer2_outputs(7704) <= layer1_outputs(12798);
    layer2_outputs(7705) <= not((layer1_outputs(9636)) and (layer1_outputs(3234)));
    layer2_outputs(7706) <= not(layer1_outputs(787));
    layer2_outputs(7707) <= not(layer1_outputs(7609)) or (layer1_outputs(2905));
    layer2_outputs(7708) <= (layer1_outputs(8775)) or (layer1_outputs(12348));
    layer2_outputs(7709) <= (layer1_outputs(8141)) and not (layer1_outputs(5735));
    layer2_outputs(7710) <= (layer1_outputs(9890)) and not (layer1_outputs(7584));
    layer2_outputs(7711) <= not(layer1_outputs(10296)) or (layer1_outputs(1854));
    layer2_outputs(7712) <= (layer1_outputs(7869)) xor (layer1_outputs(1133));
    layer2_outputs(7713) <= not((layer1_outputs(3724)) xor (layer1_outputs(4924)));
    layer2_outputs(7714) <= not(layer1_outputs(5506)) or (layer1_outputs(7495));
    layer2_outputs(7715) <= layer1_outputs(413);
    layer2_outputs(7716) <= layer1_outputs(9279);
    layer2_outputs(7717) <= not(layer1_outputs(11767));
    layer2_outputs(7718) <= (layer1_outputs(6600)) and (layer1_outputs(1658));
    layer2_outputs(7719) <= layer1_outputs(2129);
    layer2_outputs(7720) <= not((layer1_outputs(10965)) or (layer1_outputs(5597)));
    layer2_outputs(7721) <= not((layer1_outputs(1476)) and (layer1_outputs(11470)));
    layer2_outputs(7722) <= (layer1_outputs(256)) or (layer1_outputs(8368));
    layer2_outputs(7723) <= layer1_outputs(10391);
    layer2_outputs(7724) <= layer1_outputs(6814);
    layer2_outputs(7725) <= not((layer1_outputs(10065)) or (layer1_outputs(829)));
    layer2_outputs(7726) <= not(layer1_outputs(4917));
    layer2_outputs(7727) <= layer1_outputs(12605);
    layer2_outputs(7728) <= not(layer1_outputs(5980));
    layer2_outputs(7729) <= not(layer1_outputs(9243)) or (layer1_outputs(5855));
    layer2_outputs(7730) <= not((layer1_outputs(10318)) and (layer1_outputs(12654)));
    layer2_outputs(7731) <= not((layer1_outputs(5067)) or (layer1_outputs(8815)));
    layer2_outputs(7732) <= layer1_outputs(4903);
    layer2_outputs(7733) <= not(layer1_outputs(12609));
    layer2_outputs(7734) <= not((layer1_outputs(7038)) xor (layer1_outputs(4371)));
    layer2_outputs(7735) <= (layer1_outputs(4996)) or (layer1_outputs(7810));
    layer2_outputs(7736) <= not(layer1_outputs(11004));
    layer2_outputs(7737) <= (layer1_outputs(11724)) and not (layer1_outputs(3696));
    layer2_outputs(7738) <= not(layer1_outputs(2685)) or (layer1_outputs(1002));
    layer2_outputs(7739) <= layer1_outputs(5853);
    layer2_outputs(7740) <= not(layer1_outputs(801));
    layer2_outputs(7741) <= not(layer1_outputs(1365));
    layer2_outputs(7742) <= not(layer1_outputs(856));
    layer2_outputs(7743) <= not(layer1_outputs(855));
    layer2_outputs(7744) <= not(layer1_outputs(4877));
    layer2_outputs(7745) <= layer1_outputs(3062);
    layer2_outputs(7746) <= (layer1_outputs(2054)) and (layer1_outputs(7129));
    layer2_outputs(7747) <= not(layer1_outputs(9329));
    layer2_outputs(7748) <= (layer1_outputs(11443)) and not (layer1_outputs(10825));
    layer2_outputs(7749) <= not(layer1_outputs(6046));
    layer2_outputs(7750) <= not(layer1_outputs(10720)) or (layer1_outputs(11564));
    layer2_outputs(7751) <= not(layer1_outputs(7092));
    layer2_outputs(7752) <= (layer1_outputs(1336)) and not (layer1_outputs(6916));
    layer2_outputs(7753) <= layer1_outputs(1773);
    layer2_outputs(7754) <= layer1_outputs(1309);
    layer2_outputs(7755) <= (layer1_outputs(6842)) and (layer1_outputs(9892));
    layer2_outputs(7756) <= layer1_outputs(5307);
    layer2_outputs(7757) <= not(layer1_outputs(9355));
    layer2_outputs(7758) <= not((layer1_outputs(9592)) xor (layer1_outputs(7062)));
    layer2_outputs(7759) <= layer1_outputs(9930);
    layer2_outputs(7760) <= not(layer1_outputs(5150));
    layer2_outputs(7761) <= (layer1_outputs(6778)) and not (layer1_outputs(807));
    layer2_outputs(7762) <= not((layer1_outputs(4491)) or (layer1_outputs(12522)));
    layer2_outputs(7763) <= not((layer1_outputs(3236)) and (layer1_outputs(7191)));
    layer2_outputs(7764) <= layer1_outputs(7444);
    layer2_outputs(7765) <= (layer1_outputs(1021)) and not (layer1_outputs(4677));
    layer2_outputs(7766) <= layer1_outputs(9009);
    layer2_outputs(7767) <= not((layer1_outputs(5116)) or (layer1_outputs(4661)));
    layer2_outputs(7768) <= layer1_outputs(8357);
    layer2_outputs(7769) <= layer1_outputs(4610);
    layer2_outputs(7770) <= (layer1_outputs(7405)) and not (layer1_outputs(5069));
    layer2_outputs(7771) <= not(layer1_outputs(9077));
    layer2_outputs(7772) <= (layer1_outputs(3475)) and not (layer1_outputs(10867));
    layer2_outputs(7773) <= (layer1_outputs(10206)) and (layer1_outputs(9601));
    layer2_outputs(7774) <= not(layer1_outputs(6966));
    layer2_outputs(7775) <= (layer1_outputs(4774)) and (layer1_outputs(7396));
    layer2_outputs(7776) <= not((layer1_outputs(8155)) xor (layer1_outputs(8503)));
    layer2_outputs(7777) <= (layer1_outputs(7836)) and not (layer1_outputs(2015));
    layer2_outputs(7778) <= not(layer1_outputs(7586)) or (layer1_outputs(6986));
    layer2_outputs(7779) <= (layer1_outputs(295)) or (layer1_outputs(9350));
    layer2_outputs(7780) <= not(layer1_outputs(7799)) or (layer1_outputs(2633));
    layer2_outputs(7781) <= not(layer1_outputs(4384)) or (layer1_outputs(894));
    layer2_outputs(7782) <= (layer1_outputs(8422)) and (layer1_outputs(346));
    layer2_outputs(7783) <= layer1_outputs(12370);
    layer2_outputs(7784) <= not((layer1_outputs(1558)) or (layer1_outputs(9236)));
    layer2_outputs(7785) <= layer1_outputs(3693);
    layer2_outputs(7786) <= (layer1_outputs(3086)) and not (layer1_outputs(5887));
    layer2_outputs(7787) <= (layer1_outputs(3744)) or (layer1_outputs(10002));
    layer2_outputs(7788) <= not(layer1_outputs(7554)) or (layer1_outputs(7432));
    layer2_outputs(7789) <= layer1_outputs(8037);
    layer2_outputs(7790) <= not(layer1_outputs(6915));
    layer2_outputs(7791) <= not((layer1_outputs(4426)) or (layer1_outputs(3188)));
    layer2_outputs(7792) <= not(layer1_outputs(8167));
    layer2_outputs(7793) <= not(layer1_outputs(10432));
    layer2_outputs(7794) <= not((layer1_outputs(11566)) or (layer1_outputs(1176)));
    layer2_outputs(7795) <= layer1_outputs(3440);
    layer2_outputs(7796) <= not((layer1_outputs(10263)) or (layer1_outputs(8609)));
    layer2_outputs(7797) <= (layer1_outputs(8253)) and not (layer1_outputs(1087));
    layer2_outputs(7798) <= (layer1_outputs(486)) and not (layer1_outputs(2617));
    layer2_outputs(7799) <= not((layer1_outputs(2053)) or (layer1_outputs(12169)));
    layer2_outputs(7800) <= layer1_outputs(3635);
    layer2_outputs(7801) <= not(layer1_outputs(5568)) or (layer1_outputs(1178));
    layer2_outputs(7802) <= not(layer1_outputs(10592));
    layer2_outputs(7803) <= layer1_outputs(7049);
    layer2_outputs(7804) <= not(layer1_outputs(626));
    layer2_outputs(7805) <= not(layer1_outputs(4263));
    layer2_outputs(7806) <= not(layer1_outputs(10020));
    layer2_outputs(7807) <= not(layer1_outputs(7710)) or (layer1_outputs(8365));
    layer2_outputs(7808) <= not((layer1_outputs(5508)) xor (layer1_outputs(4235)));
    layer2_outputs(7809) <= layer1_outputs(277);
    layer2_outputs(7810) <= not(layer1_outputs(1876));
    layer2_outputs(7811) <= (layer1_outputs(10731)) xor (layer1_outputs(6373));
    layer2_outputs(7812) <= layer1_outputs(11390);
    layer2_outputs(7813) <= not(layer1_outputs(1205));
    layer2_outputs(7814) <= not((layer1_outputs(5098)) xor (layer1_outputs(841)));
    layer2_outputs(7815) <= not((layer1_outputs(1362)) or (layer1_outputs(8905)));
    layer2_outputs(7816) <= (layer1_outputs(5760)) xor (layer1_outputs(7625));
    layer2_outputs(7817) <= layer1_outputs(519);
    layer2_outputs(7818) <= not(layer1_outputs(1285)) or (layer1_outputs(7890));
    layer2_outputs(7819) <= not((layer1_outputs(1447)) xor (layer1_outputs(3976)));
    layer2_outputs(7820) <= layer1_outputs(6809);
    layer2_outputs(7821) <= (layer1_outputs(4534)) or (layer1_outputs(4934));
    layer2_outputs(7822) <= (layer1_outputs(3435)) or (layer1_outputs(8809));
    layer2_outputs(7823) <= layer1_outputs(3340);
    layer2_outputs(7824) <= layer1_outputs(7803);
    layer2_outputs(7825) <= not(layer1_outputs(6267));
    layer2_outputs(7826) <= layer1_outputs(2306);
    layer2_outputs(7827) <= layer1_outputs(8455);
    layer2_outputs(7828) <= not(layer1_outputs(7764));
    layer2_outputs(7829) <= (layer1_outputs(11391)) xor (layer1_outputs(7020));
    layer2_outputs(7830) <= not(layer1_outputs(1006));
    layer2_outputs(7831) <= (layer1_outputs(934)) and not (layer1_outputs(3419));
    layer2_outputs(7832) <= (layer1_outputs(1708)) and not (layer1_outputs(9014));
    layer2_outputs(7833) <= not(layer1_outputs(874));
    layer2_outputs(7834) <= not(layer1_outputs(4201));
    layer2_outputs(7835) <= not((layer1_outputs(2339)) and (layer1_outputs(3719)));
    layer2_outputs(7836) <= (layer1_outputs(12497)) or (layer1_outputs(5497));
    layer2_outputs(7837) <= (layer1_outputs(12512)) xor (layer1_outputs(672));
    layer2_outputs(7838) <= not(layer1_outputs(8708));
    layer2_outputs(7839) <= layer1_outputs(6358);
    layer2_outputs(7840) <= not((layer1_outputs(9792)) xor (layer1_outputs(6578)));
    layer2_outputs(7841) <= not((layer1_outputs(8402)) and (layer1_outputs(5215)));
    layer2_outputs(7842) <= (layer1_outputs(10122)) and not (layer1_outputs(12385));
    layer2_outputs(7843) <= (layer1_outputs(10574)) xor (layer1_outputs(8771));
    layer2_outputs(7844) <= not((layer1_outputs(5591)) or (layer1_outputs(7689)));
    layer2_outputs(7845) <= not((layer1_outputs(1660)) and (layer1_outputs(8357)));
    layer2_outputs(7846) <= (layer1_outputs(1370)) and not (layer1_outputs(10936));
    layer2_outputs(7847) <= not((layer1_outputs(7133)) xor (layer1_outputs(411)));
    layer2_outputs(7848) <= (layer1_outputs(37)) xor (layer1_outputs(8653));
    layer2_outputs(7849) <= (layer1_outputs(4381)) and not (layer1_outputs(12448));
    layer2_outputs(7850) <= not(layer1_outputs(2373));
    layer2_outputs(7851) <= not(layer1_outputs(11343));
    layer2_outputs(7852) <= layer1_outputs(3048);
    layer2_outputs(7853) <= (layer1_outputs(2989)) and not (layer1_outputs(10966));
    layer2_outputs(7854) <= layer1_outputs(7660);
    layer2_outputs(7855) <= not(layer1_outputs(6383));
    layer2_outputs(7856) <= layer1_outputs(4788);
    layer2_outputs(7857) <= (layer1_outputs(7981)) or (layer1_outputs(9861));
    layer2_outputs(7858) <= not((layer1_outputs(12244)) and (layer1_outputs(2508)));
    layer2_outputs(7859) <= layer1_outputs(5080);
    layer2_outputs(7860) <= not(layer1_outputs(3612));
    layer2_outputs(7861) <= layer1_outputs(6384);
    layer2_outputs(7862) <= not(layer1_outputs(11944));
    layer2_outputs(7863) <= (layer1_outputs(7851)) and not (layer1_outputs(1952));
    layer2_outputs(7864) <= not((layer1_outputs(2377)) and (layer1_outputs(9111)));
    layer2_outputs(7865) <= not((layer1_outputs(5934)) or (layer1_outputs(10820)));
    layer2_outputs(7866) <= layer1_outputs(533);
    layer2_outputs(7867) <= (layer1_outputs(5461)) xor (layer1_outputs(110));
    layer2_outputs(7868) <= not(layer1_outputs(8619));
    layer2_outputs(7869) <= not((layer1_outputs(8282)) and (layer1_outputs(8578)));
    layer2_outputs(7870) <= (layer1_outputs(11544)) xor (layer1_outputs(5961));
    layer2_outputs(7871) <= not(layer1_outputs(12258));
    layer2_outputs(7872) <= not(layer1_outputs(1059));
    layer2_outputs(7873) <= layer1_outputs(9409);
    layer2_outputs(7874) <= layer1_outputs(11362);
    layer2_outputs(7875) <= not((layer1_outputs(10792)) or (layer1_outputs(6180)));
    layer2_outputs(7876) <= not(layer1_outputs(7021));
    layer2_outputs(7877) <= (layer1_outputs(315)) and (layer1_outputs(4343));
    layer2_outputs(7878) <= layer1_outputs(9195);
    layer2_outputs(7879) <= (layer1_outputs(8844)) xor (layer1_outputs(6789));
    layer2_outputs(7880) <= (layer1_outputs(6270)) and (layer1_outputs(12154));
    layer2_outputs(7881) <= layer1_outputs(3957);
    layer2_outputs(7882) <= (layer1_outputs(10925)) and not (layer1_outputs(11382));
    layer2_outputs(7883) <= layer1_outputs(2869);
    layer2_outputs(7884) <= layer1_outputs(12473);
    layer2_outputs(7885) <= not((layer1_outputs(12139)) or (layer1_outputs(8204)));
    layer2_outputs(7886) <= (layer1_outputs(777)) xor (layer1_outputs(5775));
    layer2_outputs(7887) <= not(layer1_outputs(1130));
    layer2_outputs(7888) <= not(layer1_outputs(12031)) or (layer1_outputs(3267));
    layer2_outputs(7889) <= not(layer1_outputs(7620));
    layer2_outputs(7890) <= not(layer1_outputs(4925));
    layer2_outputs(7891) <= (layer1_outputs(4321)) or (layer1_outputs(3689));
    layer2_outputs(7892) <= (layer1_outputs(11154)) and not (layer1_outputs(1188));
    layer2_outputs(7893) <= (layer1_outputs(3078)) and not (layer1_outputs(10413));
    layer2_outputs(7894) <= layer1_outputs(12131);
    layer2_outputs(7895) <= not(layer1_outputs(3055)) or (layer1_outputs(5347));
    layer2_outputs(7896) <= not(layer1_outputs(12233));
    layer2_outputs(7897) <= not(layer1_outputs(4470)) or (layer1_outputs(3986));
    layer2_outputs(7898) <= (layer1_outputs(3778)) and not (layer1_outputs(5337));
    layer2_outputs(7899) <= not(layer1_outputs(3944));
    layer2_outputs(7900) <= layer1_outputs(3953);
    layer2_outputs(7901) <= not((layer1_outputs(8308)) or (layer1_outputs(2898)));
    layer2_outputs(7902) <= layer1_outputs(7476);
    layer2_outputs(7903) <= not(layer1_outputs(1157)) or (layer1_outputs(10628));
    layer2_outputs(7904) <= not(layer1_outputs(3330));
    layer2_outputs(7905) <= not((layer1_outputs(11863)) or (layer1_outputs(5629)));
    layer2_outputs(7906) <= layer1_outputs(10423);
    layer2_outputs(7907) <= (layer1_outputs(6972)) xor (layer1_outputs(3695));
    layer2_outputs(7908) <= not((layer1_outputs(1348)) and (layer1_outputs(10018)));
    layer2_outputs(7909) <= layer1_outputs(9648);
    layer2_outputs(7910) <= layer1_outputs(1549);
    layer2_outputs(7911) <= (layer1_outputs(8158)) or (layer1_outputs(2265));
    layer2_outputs(7912) <= not((layer1_outputs(9837)) xor (layer1_outputs(463)));
    layer2_outputs(7913) <= layer1_outputs(10834);
    layer2_outputs(7914) <= (layer1_outputs(1452)) and (layer1_outputs(9049));
    layer2_outputs(7915) <= not(layer1_outputs(428));
    layer2_outputs(7916) <= not(layer1_outputs(1827));
    layer2_outputs(7917) <= not(layer1_outputs(3934)) or (layer1_outputs(12110));
    layer2_outputs(7918) <= not((layer1_outputs(2103)) xor (layer1_outputs(5246)));
    layer2_outputs(7919) <= (layer1_outputs(5985)) and not (layer1_outputs(10304));
    layer2_outputs(7920) <= not(layer1_outputs(8937));
    layer2_outputs(7921) <= not(layer1_outputs(8057));
    layer2_outputs(7922) <= (layer1_outputs(7360)) or (layer1_outputs(10266));
    layer2_outputs(7923) <= not((layer1_outputs(5030)) and (layer1_outputs(8285)));
    layer2_outputs(7924) <= (layer1_outputs(10298)) and not (layer1_outputs(12636));
    layer2_outputs(7925) <= not(layer1_outputs(3768));
    layer2_outputs(7926) <= (layer1_outputs(284)) or (layer1_outputs(5951));
    layer2_outputs(7927) <= not((layer1_outputs(12394)) and (layer1_outputs(5666)));
    layer2_outputs(7928) <= layer1_outputs(3906);
    layer2_outputs(7929) <= layer1_outputs(1508);
    layer2_outputs(7930) <= not((layer1_outputs(2132)) xor (layer1_outputs(2773)));
    layer2_outputs(7931) <= layer1_outputs(6548);
    layer2_outputs(7932) <= (layer1_outputs(10362)) and not (layer1_outputs(1285));
    layer2_outputs(7933) <= layer1_outputs(12306);
    layer2_outputs(7934) <= '1';
    layer2_outputs(7935) <= (layer1_outputs(5596)) and not (layer1_outputs(5206));
    layer2_outputs(7936) <= (layer1_outputs(2609)) or (layer1_outputs(11922));
    layer2_outputs(7937) <= not(layer1_outputs(2723));
    layer2_outputs(7938) <= (layer1_outputs(5121)) xor (layer1_outputs(11474));
    layer2_outputs(7939) <= layer1_outputs(3612);
    layer2_outputs(7940) <= layer1_outputs(5594);
    layer2_outputs(7941) <= layer1_outputs(3199);
    layer2_outputs(7942) <= not(layer1_outputs(2872));
    layer2_outputs(7943) <= not((layer1_outputs(830)) or (layer1_outputs(1456)));
    layer2_outputs(7944) <= not(layer1_outputs(8532));
    layer2_outputs(7945) <= layer1_outputs(11557);
    layer2_outputs(7946) <= not(layer1_outputs(6699)) or (layer1_outputs(10249));
    layer2_outputs(7947) <= layer1_outputs(7951);
    layer2_outputs(7948) <= layer1_outputs(5002);
    layer2_outputs(7949) <= not(layer1_outputs(10729));
    layer2_outputs(7950) <= not(layer1_outputs(815));
    layer2_outputs(7951) <= layer1_outputs(208);
    layer2_outputs(7952) <= layer1_outputs(8457);
    layer2_outputs(7953) <= not((layer1_outputs(314)) or (layer1_outputs(689)));
    layer2_outputs(7954) <= layer1_outputs(1473);
    layer2_outputs(7955) <= (layer1_outputs(12219)) and (layer1_outputs(5404));
    layer2_outputs(7956) <= not(layer1_outputs(554));
    layer2_outputs(7957) <= not((layer1_outputs(12413)) xor (layer1_outputs(2290)));
    layer2_outputs(7958) <= not((layer1_outputs(65)) xor (layer1_outputs(11180)));
    layer2_outputs(7959) <= not(layer1_outputs(11602));
    layer2_outputs(7960) <= not(layer1_outputs(6297));
    layer2_outputs(7961) <= not(layer1_outputs(8088)) or (layer1_outputs(2915));
    layer2_outputs(7962) <= not(layer1_outputs(11375));
    layer2_outputs(7963) <= not(layer1_outputs(7368));
    layer2_outputs(7964) <= not(layer1_outputs(10647));
    layer2_outputs(7965) <= not(layer1_outputs(11658));
    layer2_outputs(7966) <= not(layer1_outputs(9963));
    layer2_outputs(7967) <= not((layer1_outputs(221)) or (layer1_outputs(1654)));
    layer2_outputs(7968) <= (layer1_outputs(1480)) xor (layer1_outputs(209));
    layer2_outputs(7969) <= layer1_outputs(8302);
    layer2_outputs(7970) <= (layer1_outputs(11361)) and not (layer1_outputs(1032));
    layer2_outputs(7971) <= not(layer1_outputs(1774));
    layer2_outputs(7972) <= not(layer1_outputs(12750));
    layer2_outputs(7973) <= '0';
    layer2_outputs(7974) <= (layer1_outputs(450)) and not (layer1_outputs(7966));
    layer2_outputs(7975) <= not(layer1_outputs(9758));
    layer2_outputs(7976) <= (layer1_outputs(1204)) xor (layer1_outputs(6677));
    layer2_outputs(7977) <= not((layer1_outputs(3055)) or (layer1_outputs(4545)));
    layer2_outputs(7978) <= not(layer1_outputs(9681));
    layer2_outputs(7979) <= (layer1_outputs(1500)) and not (layer1_outputs(2652));
    layer2_outputs(7980) <= not(layer1_outputs(5632)) or (layer1_outputs(6479));
    layer2_outputs(7981) <= layer1_outputs(11537);
    layer2_outputs(7982) <= not((layer1_outputs(9037)) xor (layer1_outputs(6808)));
    layer2_outputs(7983) <= not(layer1_outputs(10690)) or (layer1_outputs(599));
    layer2_outputs(7984) <= not((layer1_outputs(7263)) and (layer1_outputs(4604)));
    layer2_outputs(7985) <= (layer1_outputs(12511)) or (layer1_outputs(3371));
    layer2_outputs(7986) <= layer1_outputs(3067);
    layer2_outputs(7987) <= (layer1_outputs(689)) xor (layer1_outputs(10155));
    layer2_outputs(7988) <= not(layer1_outputs(1682));
    layer2_outputs(7989) <= not((layer1_outputs(2854)) or (layer1_outputs(9933)));
    layer2_outputs(7990) <= layer1_outputs(12165);
    layer2_outputs(7991) <= layer1_outputs(750);
    layer2_outputs(7992) <= not((layer1_outputs(1580)) xor (layer1_outputs(5341)));
    layer2_outputs(7993) <= not((layer1_outputs(5023)) xor (layer1_outputs(6841)));
    layer2_outputs(7994) <= not(layer1_outputs(6838));
    layer2_outputs(7995) <= (layer1_outputs(11873)) and (layer1_outputs(1312));
    layer2_outputs(7996) <= layer1_outputs(7093);
    layer2_outputs(7997) <= not(layer1_outputs(183));
    layer2_outputs(7998) <= not(layer1_outputs(3386)) or (layer1_outputs(856));
    layer2_outputs(7999) <= not(layer1_outputs(11933));
    layer2_outputs(8000) <= layer1_outputs(7259);
    layer2_outputs(8001) <= (layer1_outputs(1175)) and not (layer1_outputs(2999));
    layer2_outputs(8002) <= not(layer1_outputs(9204));
    layer2_outputs(8003) <= not(layer1_outputs(10447));
    layer2_outputs(8004) <= not(layer1_outputs(6735));
    layer2_outputs(8005) <= not(layer1_outputs(9169));
    layer2_outputs(8006) <= not(layer1_outputs(8639)) or (layer1_outputs(2761));
    layer2_outputs(8007) <= layer1_outputs(881);
    layer2_outputs(8008) <= (layer1_outputs(11242)) and not (layer1_outputs(12636));
    layer2_outputs(8009) <= not(layer1_outputs(10258)) or (layer1_outputs(12187));
    layer2_outputs(8010) <= not(layer1_outputs(8041));
    layer2_outputs(8011) <= not(layer1_outputs(10207));
    layer2_outputs(8012) <= layer1_outputs(2311);
    layer2_outputs(8013) <= not((layer1_outputs(5804)) xor (layer1_outputs(12787)));
    layer2_outputs(8014) <= not(layer1_outputs(10803));
    layer2_outputs(8015) <= (layer1_outputs(4697)) xor (layer1_outputs(3134));
    layer2_outputs(8016) <= (layer1_outputs(7388)) and not (layer1_outputs(4053));
    layer2_outputs(8017) <= not(layer1_outputs(4667));
    layer2_outputs(8018) <= (layer1_outputs(1883)) and not (layer1_outputs(1871));
    layer2_outputs(8019) <= '0';
    layer2_outputs(8020) <= layer1_outputs(9145);
    layer2_outputs(8021) <= not(layer1_outputs(11765));
    layer2_outputs(8022) <= not(layer1_outputs(1915));
    layer2_outputs(8023) <= not((layer1_outputs(12481)) xor (layer1_outputs(5803)));
    layer2_outputs(8024) <= layer1_outputs(1592);
    layer2_outputs(8025) <= layer1_outputs(12393);
    layer2_outputs(8026) <= not(layer1_outputs(9061)) or (layer1_outputs(4637));
    layer2_outputs(8027) <= layer1_outputs(7075);
    layer2_outputs(8028) <= not(layer1_outputs(1817));
    layer2_outputs(8029) <= (layer1_outputs(6002)) or (layer1_outputs(6513));
    layer2_outputs(8030) <= not(layer1_outputs(6692));
    layer2_outputs(8031) <= not((layer1_outputs(4371)) xor (layer1_outputs(1079)));
    layer2_outputs(8032) <= layer1_outputs(8694);
    layer2_outputs(8033) <= not(layer1_outputs(7060));
    layer2_outputs(8034) <= layer1_outputs(7565);
    layer2_outputs(8035) <= not((layer1_outputs(7497)) xor (layer1_outputs(1830)));
    layer2_outputs(8036) <= (layer1_outputs(7292)) or (layer1_outputs(11113));
    layer2_outputs(8037) <= (layer1_outputs(12369)) xor (layer1_outputs(11649));
    layer2_outputs(8038) <= layer1_outputs(7930);
    layer2_outputs(8039) <= not(layer1_outputs(6240));
    layer2_outputs(8040) <= (layer1_outputs(6928)) and not (layer1_outputs(9966));
    layer2_outputs(8041) <= layer1_outputs(11462);
    layer2_outputs(8042) <= not(layer1_outputs(2359)) or (layer1_outputs(6523));
    layer2_outputs(8043) <= not(layer1_outputs(3790));
    layer2_outputs(8044) <= not((layer1_outputs(3016)) xor (layer1_outputs(11323)));
    layer2_outputs(8045) <= layer1_outputs(8064);
    layer2_outputs(8046) <= (layer1_outputs(2538)) xor (layer1_outputs(9900));
    layer2_outputs(8047) <= layer1_outputs(7633);
    layer2_outputs(8048) <= not(layer1_outputs(218));
    layer2_outputs(8049) <= (layer1_outputs(4887)) xor (layer1_outputs(6947));
    layer2_outputs(8050) <= not(layer1_outputs(4185));
    layer2_outputs(8051) <= layer1_outputs(2559);
    layer2_outputs(8052) <= (layer1_outputs(1821)) and (layer1_outputs(11108));
    layer2_outputs(8053) <= (layer1_outputs(1278)) xor (layer1_outputs(549));
    layer2_outputs(8054) <= not(layer1_outputs(3747));
    layer2_outputs(8055) <= not(layer1_outputs(1741));
    layer2_outputs(8056) <= not(layer1_outputs(7150));
    layer2_outputs(8057) <= layer1_outputs(9185);
    layer2_outputs(8058) <= not(layer1_outputs(2962)) or (layer1_outputs(6535));
    layer2_outputs(8059) <= (layer1_outputs(9386)) or (layer1_outputs(11188));
    layer2_outputs(8060) <= (layer1_outputs(11063)) and not (layer1_outputs(4833));
    layer2_outputs(8061) <= not(layer1_outputs(12616)) or (layer1_outputs(5241));
    layer2_outputs(8062) <= not(layer1_outputs(12095)) or (layer1_outputs(803));
    layer2_outputs(8063) <= layer1_outputs(9540);
    layer2_outputs(8064) <= layer1_outputs(6814);
    layer2_outputs(8065) <= not(layer1_outputs(5797)) or (layer1_outputs(514));
    layer2_outputs(8066) <= (layer1_outputs(11120)) and (layer1_outputs(5733));
    layer2_outputs(8067) <= not(layer1_outputs(6238)) or (layer1_outputs(5658));
    layer2_outputs(8068) <= layer1_outputs(6486);
    layer2_outputs(8069) <= layer1_outputs(4687);
    layer2_outputs(8070) <= (layer1_outputs(3025)) or (layer1_outputs(12100));
    layer2_outputs(8071) <= layer1_outputs(8528);
    layer2_outputs(8072) <= not((layer1_outputs(1265)) and (layer1_outputs(9700)));
    layer2_outputs(8073) <= (layer1_outputs(3515)) or (layer1_outputs(11560));
    layer2_outputs(8074) <= not((layer1_outputs(1301)) or (layer1_outputs(7691)));
    layer2_outputs(8075) <= (layer1_outputs(10168)) and (layer1_outputs(8965));
    layer2_outputs(8076) <= '0';
    layer2_outputs(8077) <= (layer1_outputs(4333)) or (layer1_outputs(28));
    layer2_outputs(8078) <= not(layer1_outputs(906)) or (layer1_outputs(6100));
    layer2_outputs(8079) <= layer1_outputs(6392);
    layer2_outputs(8080) <= not(layer1_outputs(5196)) or (layer1_outputs(5972));
    layer2_outputs(8081) <= not((layer1_outputs(12697)) or (layer1_outputs(6519)));
    layer2_outputs(8082) <= layer1_outputs(4573);
    layer2_outputs(8083) <= not(layer1_outputs(4214));
    layer2_outputs(8084) <= layer1_outputs(1870);
    layer2_outputs(8085) <= not(layer1_outputs(1095)) or (layer1_outputs(6076));
    layer2_outputs(8086) <= not(layer1_outputs(7096));
    layer2_outputs(8087) <= layer1_outputs(8696);
    layer2_outputs(8088) <= (layer1_outputs(7967)) xor (layer1_outputs(10577));
    layer2_outputs(8089) <= not(layer1_outputs(9385));
    layer2_outputs(8090) <= not(layer1_outputs(10117)) or (layer1_outputs(8381));
    layer2_outputs(8091) <= not(layer1_outputs(2246));
    layer2_outputs(8092) <= (layer1_outputs(1978)) and not (layer1_outputs(5594));
    layer2_outputs(8093) <= layer1_outputs(2995);
    layer2_outputs(8094) <= not((layer1_outputs(2428)) xor (layer1_outputs(6967)));
    layer2_outputs(8095) <= layer1_outputs(1443);
    layer2_outputs(8096) <= not((layer1_outputs(11988)) xor (layer1_outputs(7382)));
    layer2_outputs(8097) <= not((layer1_outputs(11431)) xor (layer1_outputs(2877)));
    layer2_outputs(8098) <= (layer1_outputs(5200)) and not (layer1_outputs(7362));
    layer2_outputs(8099) <= not(layer1_outputs(3313));
    layer2_outputs(8100) <= not(layer1_outputs(6092));
    layer2_outputs(8101) <= not((layer1_outputs(11485)) and (layer1_outputs(6793)));
    layer2_outputs(8102) <= not(layer1_outputs(4308)) or (layer1_outputs(12439));
    layer2_outputs(8103) <= (layer1_outputs(11016)) or (layer1_outputs(245));
    layer2_outputs(8104) <= layer1_outputs(8753);
    layer2_outputs(8105) <= (layer1_outputs(11203)) xor (layer1_outputs(7559));
    layer2_outputs(8106) <= (layer1_outputs(704)) xor (layer1_outputs(1516));
    layer2_outputs(8107) <= (layer1_outputs(3404)) and not (layer1_outputs(6590));
    layer2_outputs(8108) <= (layer1_outputs(260)) or (layer1_outputs(10137));
    layer2_outputs(8109) <= not(layer1_outputs(10015)) or (layer1_outputs(3375));
    layer2_outputs(8110) <= not(layer1_outputs(4087)) or (layer1_outputs(5566));
    layer2_outputs(8111) <= layer1_outputs(6278);
    layer2_outputs(8112) <= not(layer1_outputs(3279));
    layer2_outputs(8113) <= not(layer1_outputs(1305)) or (layer1_outputs(11526));
    layer2_outputs(8114) <= not(layer1_outputs(12118));
    layer2_outputs(8115) <= layer1_outputs(819);
    layer2_outputs(8116) <= not(layer1_outputs(673));
    layer2_outputs(8117) <= layer1_outputs(5245);
    layer2_outputs(8118) <= not(layer1_outputs(6874));
    layer2_outputs(8119) <= layer1_outputs(1406);
    layer2_outputs(8120) <= layer1_outputs(7661);
    layer2_outputs(8121) <= not(layer1_outputs(9744));
    layer2_outputs(8122) <= not((layer1_outputs(7158)) or (layer1_outputs(7261)));
    layer2_outputs(8123) <= not(layer1_outputs(10111));
    layer2_outputs(8124) <= (layer1_outputs(1985)) xor (layer1_outputs(587));
    layer2_outputs(8125) <= layer1_outputs(1131);
    layer2_outputs(8126) <= not(layer1_outputs(4286)) or (layer1_outputs(641));
    layer2_outputs(8127) <= (layer1_outputs(10964)) and (layer1_outputs(5895));
    layer2_outputs(8128) <= layer1_outputs(3653);
    layer2_outputs(8129) <= (layer1_outputs(10716)) or (layer1_outputs(4022));
    layer2_outputs(8130) <= not(layer1_outputs(6509));
    layer2_outputs(8131) <= layer1_outputs(1268);
    layer2_outputs(8132) <= not((layer1_outputs(8978)) xor (layer1_outputs(7147)));
    layer2_outputs(8133) <= layer1_outputs(5679);
    layer2_outputs(8134) <= not((layer1_outputs(1761)) xor (layer1_outputs(2002)));
    layer2_outputs(8135) <= (layer1_outputs(9541)) xor (layer1_outputs(1574));
    layer2_outputs(8136) <= layer1_outputs(4200);
    layer2_outputs(8137) <= layer1_outputs(1579);
    layer2_outputs(8138) <= not((layer1_outputs(11291)) or (layer1_outputs(11507)));
    layer2_outputs(8139) <= not(layer1_outputs(942)) or (layer1_outputs(12594));
    layer2_outputs(8140) <= not((layer1_outputs(11094)) and (layer1_outputs(366)));
    layer2_outputs(8141) <= not(layer1_outputs(634));
    layer2_outputs(8142) <= not((layer1_outputs(3112)) or (layer1_outputs(4376)));
    layer2_outputs(8143) <= not((layer1_outputs(7714)) and (layer1_outputs(12230)));
    layer2_outputs(8144) <= (layer1_outputs(2130)) and not (layer1_outputs(7865));
    layer2_outputs(8145) <= layer1_outputs(9355);
    layer2_outputs(8146) <= layer1_outputs(12582);
    layer2_outputs(8147) <= layer1_outputs(3229);
    layer2_outputs(8148) <= layer1_outputs(11707);
    layer2_outputs(8149) <= not(layer1_outputs(1335));
    layer2_outputs(8150) <= layer1_outputs(6805);
    layer2_outputs(8151) <= not(layer1_outputs(10636));
    layer2_outputs(8152) <= not(layer1_outputs(11001)) or (layer1_outputs(2256));
    layer2_outputs(8153) <= layer1_outputs(1370);
    layer2_outputs(8154) <= not(layer1_outputs(6093)) or (layer1_outputs(5860));
    layer2_outputs(8155) <= (layer1_outputs(9041)) or (layer1_outputs(6945));
    layer2_outputs(8156) <= not(layer1_outputs(12663)) or (layer1_outputs(8168));
    layer2_outputs(8157) <= not(layer1_outputs(199));
    layer2_outputs(8158) <= (layer1_outputs(5858)) xor (layer1_outputs(12425));
    layer2_outputs(8159) <= (layer1_outputs(3710)) or (layer1_outputs(8117));
    layer2_outputs(8160) <= layer1_outputs(4769);
    layer2_outputs(8161) <= not((layer1_outputs(952)) xor (layer1_outputs(978)));
    layer2_outputs(8162) <= not((layer1_outputs(6327)) xor (layer1_outputs(9940)));
    layer2_outputs(8163) <= layer1_outputs(4524);
    layer2_outputs(8164) <= not((layer1_outputs(7862)) and (layer1_outputs(10379)));
    layer2_outputs(8165) <= not((layer1_outputs(2322)) and (layer1_outputs(3091)));
    layer2_outputs(8166) <= not(layer1_outputs(2348)) or (layer1_outputs(3755));
    layer2_outputs(8167) <= not(layer1_outputs(1590));
    layer2_outputs(8168) <= (layer1_outputs(11912)) or (layer1_outputs(1785));
    layer2_outputs(8169) <= not(layer1_outputs(12633));
    layer2_outputs(8170) <= not(layer1_outputs(2396));
    layer2_outputs(8171) <= (layer1_outputs(3202)) or (layer1_outputs(11173));
    layer2_outputs(8172) <= not(layer1_outputs(5927));
    layer2_outputs(8173) <= not(layer1_outputs(9561)) or (layer1_outputs(30));
    layer2_outputs(8174) <= not((layer1_outputs(9657)) and (layer1_outputs(4916)));
    layer2_outputs(8175) <= layer1_outputs(12108);
    layer2_outputs(8176) <= not((layer1_outputs(10132)) and (layer1_outputs(3192)));
    layer2_outputs(8177) <= layer1_outputs(11631);
    layer2_outputs(8178) <= not(layer1_outputs(4408));
    layer2_outputs(8179) <= not(layer1_outputs(12741)) or (layer1_outputs(8050));
    layer2_outputs(8180) <= layer1_outputs(895);
    layer2_outputs(8181) <= layer1_outputs(11953);
    layer2_outputs(8182) <= not(layer1_outputs(2528)) or (layer1_outputs(12649));
    layer2_outputs(8183) <= (layer1_outputs(7486)) or (layer1_outputs(11815));
    layer2_outputs(8184) <= not(layer1_outputs(7725));
    layer2_outputs(8185) <= not(layer1_outputs(12169));
    layer2_outputs(8186) <= (layer1_outputs(11251)) and not (layer1_outputs(1442));
    layer2_outputs(8187) <= not((layer1_outputs(2430)) or (layer1_outputs(2489)));
    layer2_outputs(8188) <= not(layer1_outputs(1196)) or (layer1_outputs(6120));
    layer2_outputs(8189) <= layer1_outputs(949);
    layer2_outputs(8190) <= layer1_outputs(6675);
    layer2_outputs(8191) <= not((layer1_outputs(4093)) and (layer1_outputs(975)));
    layer2_outputs(8192) <= not(layer1_outputs(2197));
    layer2_outputs(8193) <= not((layer1_outputs(6503)) xor (layer1_outputs(949)));
    layer2_outputs(8194) <= not(layer1_outputs(5725));
    layer2_outputs(8195) <= not((layer1_outputs(11644)) xor (layer1_outputs(1316)));
    layer2_outputs(8196) <= layer1_outputs(11539);
    layer2_outputs(8197) <= not(layer1_outputs(44));
    layer2_outputs(8198) <= layer1_outputs(8631);
    layer2_outputs(8199) <= layer1_outputs(12069);
    layer2_outputs(8200) <= not(layer1_outputs(7239));
    layer2_outputs(8201) <= not((layer1_outputs(10028)) xor (layer1_outputs(4406)));
    layer2_outputs(8202) <= (layer1_outputs(6424)) xor (layer1_outputs(12400));
    layer2_outputs(8203) <= (layer1_outputs(12061)) or (layer1_outputs(2066));
    layer2_outputs(8204) <= not(layer1_outputs(2505)) or (layer1_outputs(10340));
    layer2_outputs(8205) <= (layer1_outputs(2143)) xor (layer1_outputs(1989));
    layer2_outputs(8206) <= not((layer1_outputs(11573)) xor (layer1_outputs(6525)));
    layer2_outputs(8207) <= not(layer1_outputs(9254));
    layer2_outputs(8208) <= not(layer1_outputs(8060)) or (layer1_outputs(709));
    layer2_outputs(8209) <= (layer1_outputs(7732)) and not (layer1_outputs(4250));
    layer2_outputs(8210) <= layer1_outputs(4205);
    layer2_outputs(8211) <= not(layer1_outputs(11606)) or (layer1_outputs(10968));
    layer2_outputs(8212) <= (layer1_outputs(10157)) or (layer1_outputs(6573));
    layer2_outputs(8213) <= (layer1_outputs(7482)) or (layer1_outputs(8676));
    layer2_outputs(8214) <= (layer1_outputs(11445)) and not (layer1_outputs(4242));
    layer2_outputs(8215) <= not(layer1_outputs(2505)) or (layer1_outputs(2782));
    layer2_outputs(8216) <= (layer1_outputs(7908)) xor (layer1_outputs(9318));
    layer2_outputs(8217) <= not(layer1_outputs(6114)) or (layer1_outputs(8083));
    layer2_outputs(8218) <= (layer1_outputs(711)) or (layer1_outputs(10066));
    layer2_outputs(8219) <= layer1_outputs(11387);
    layer2_outputs(8220) <= (layer1_outputs(9292)) or (layer1_outputs(2055));
    layer2_outputs(8221) <= not((layer1_outputs(3722)) xor (layer1_outputs(6601)));
    layer2_outputs(8222) <= not(layer1_outputs(7067)) or (layer1_outputs(11336));
    layer2_outputs(8223) <= layer1_outputs(2260);
    layer2_outputs(8224) <= layer1_outputs(7783);
    layer2_outputs(8225) <= not((layer1_outputs(11738)) xor (layer1_outputs(11750)));
    layer2_outputs(8226) <= not(layer1_outputs(12351));
    layer2_outputs(8227) <= not(layer1_outputs(8042));
    layer2_outputs(8228) <= not(layer1_outputs(2423));
    layer2_outputs(8229) <= (layer1_outputs(4474)) and not (layer1_outputs(7587));
    layer2_outputs(8230) <= not((layer1_outputs(10303)) xor (layer1_outputs(5894)));
    layer2_outputs(8231) <= layer1_outputs(11367);
    layer2_outputs(8232) <= layer1_outputs(4290);
    layer2_outputs(8233) <= layer1_outputs(12451);
    layer2_outputs(8234) <= not(layer1_outputs(4845));
    layer2_outputs(8235) <= layer1_outputs(474);
    layer2_outputs(8236) <= not(layer1_outputs(423));
    layer2_outputs(8237) <= layer1_outputs(421);
    layer2_outputs(8238) <= not(layer1_outputs(5191)) or (layer1_outputs(3162));
    layer2_outputs(8239) <= not((layer1_outputs(8203)) and (layer1_outputs(5086)));
    layer2_outputs(8240) <= layer1_outputs(2724);
    layer2_outputs(8241) <= not(layer1_outputs(3593));
    layer2_outputs(8242) <= (layer1_outputs(3085)) and not (layer1_outputs(11283));
    layer2_outputs(8243) <= not(layer1_outputs(10683));
    layer2_outputs(8244) <= not((layer1_outputs(4945)) or (layer1_outputs(11151)));
    layer2_outputs(8245) <= not((layer1_outputs(12407)) and (layer1_outputs(3971)));
    layer2_outputs(8246) <= layer1_outputs(8593);
    layer2_outputs(8247) <= not((layer1_outputs(507)) and (layer1_outputs(11567)));
    layer2_outputs(8248) <= layer1_outputs(805);
    layer2_outputs(8249) <= layer1_outputs(481);
    layer2_outputs(8250) <= not(layer1_outputs(9762));
    layer2_outputs(8251) <= (layer1_outputs(6033)) and not (layer1_outputs(6816));
    layer2_outputs(8252) <= (layer1_outputs(5567)) xor (layer1_outputs(3687));
    layer2_outputs(8253) <= not(layer1_outputs(126));
    layer2_outputs(8254) <= '1';
    layer2_outputs(8255) <= layer1_outputs(5882);
    layer2_outputs(8256) <= not(layer1_outputs(12373)) or (layer1_outputs(9931));
    layer2_outputs(8257) <= (layer1_outputs(334)) and not (layer1_outputs(12768));
    layer2_outputs(8258) <= not(layer1_outputs(9833));
    layer2_outputs(8259) <= not(layer1_outputs(12580)) or (layer1_outputs(4839));
    layer2_outputs(8260) <= not((layer1_outputs(10752)) or (layer1_outputs(8882)));
    layer2_outputs(8261) <= not(layer1_outputs(661));
    layer2_outputs(8262) <= not(layer1_outputs(12138));
    layer2_outputs(8263) <= not((layer1_outputs(8155)) or (layer1_outputs(12670)));
    layer2_outputs(8264) <= layer1_outputs(1486);
    layer2_outputs(8265) <= (layer1_outputs(5738)) and (layer1_outputs(8574));
    layer2_outputs(8266) <= not(layer1_outputs(5642));
    layer2_outputs(8267) <= not(layer1_outputs(6458)) or (layer1_outputs(313));
    layer2_outputs(8268) <= not(layer1_outputs(2252));
    layer2_outputs(8269) <= (layer1_outputs(3932)) and (layer1_outputs(12201));
    layer2_outputs(8270) <= layer1_outputs(5838);
    layer2_outputs(8271) <= layer1_outputs(5104);
    layer2_outputs(8272) <= layer1_outputs(7408);
    layer2_outputs(8273) <= not((layer1_outputs(135)) and (layer1_outputs(8477)));
    layer2_outputs(8274) <= not(layer1_outputs(9778));
    layer2_outputs(8275) <= (layer1_outputs(1623)) or (layer1_outputs(4534));
    layer2_outputs(8276) <= layer1_outputs(7521);
    layer2_outputs(8277) <= (layer1_outputs(10578)) or (layer1_outputs(5063));
    layer2_outputs(8278) <= layer1_outputs(11593);
    layer2_outputs(8279) <= not(layer1_outputs(12667)) or (layer1_outputs(11389));
    layer2_outputs(8280) <= not((layer1_outputs(4991)) xor (layer1_outputs(10086)));
    layer2_outputs(8281) <= layer1_outputs(7009);
    layer2_outputs(8282) <= (layer1_outputs(7024)) and not (layer1_outputs(8216));
    layer2_outputs(8283) <= not(layer1_outputs(6230));
    layer2_outputs(8284) <= (layer1_outputs(12231)) or (layer1_outputs(9231));
    layer2_outputs(8285) <= not(layer1_outputs(8457));
    layer2_outputs(8286) <= (layer1_outputs(4670)) xor (layer1_outputs(6021));
    layer2_outputs(8287) <= layer1_outputs(7839);
    layer2_outputs(8288) <= not((layer1_outputs(8788)) and (layer1_outputs(4953)));
    layer2_outputs(8289) <= not((layer1_outputs(4166)) and (layer1_outputs(770)));
    layer2_outputs(8290) <= not(layer1_outputs(7620));
    layer2_outputs(8291) <= not(layer1_outputs(8748)) or (layer1_outputs(9714));
    layer2_outputs(8292) <= layer1_outputs(5921);
    layer2_outputs(8293) <= not(layer1_outputs(2508));
    layer2_outputs(8294) <= layer1_outputs(7977);
    layer2_outputs(8295) <= (layer1_outputs(12030)) xor (layer1_outputs(2429));
    layer2_outputs(8296) <= not(layer1_outputs(7127)) or (layer1_outputs(12350));
    layer2_outputs(8297) <= not(layer1_outputs(11639)) or (layer1_outputs(67));
    layer2_outputs(8298) <= layer1_outputs(7239);
    layer2_outputs(8299) <= layer1_outputs(12310);
    layer2_outputs(8300) <= (layer1_outputs(7298)) and not (layer1_outputs(1148));
    layer2_outputs(8301) <= (layer1_outputs(9458)) and (layer1_outputs(3961));
    layer2_outputs(8302) <= layer1_outputs(5640);
    layer2_outputs(8303) <= not(layer1_outputs(786));
    layer2_outputs(8304) <= layer1_outputs(5348);
    layer2_outputs(8305) <= layer1_outputs(12052);
    layer2_outputs(8306) <= layer1_outputs(3452);
    layer2_outputs(8307) <= not(layer1_outputs(2646)) or (layer1_outputs(9040));
    layer2_outputs(8308) <= not(layer1_outputs(8525));
    layer2_outputs(8309) <= (layer1_outputs(3852)) and (layer1_outputs(10660));
    layer2_outputs(8310) <= not(layer1_outputs(4554));
    layer2_outputs(8311) <= layer1_outputs(1902);
    layer2_outputs(8312) <= (layer1_outputs(11881)) and not (layer1_outputs(9064));
    layer2_outputs(8313) <= not(layer1_outputs(11026));
    layer2_outputs(8314) <= layer1_outputs(471);
    layer2_outputs(8315) <= layer1_outputs(6047);
    layer2_outputs(8316) <= not((layer1_outputs(10922)) or (layer1_outputs(1368)));
    layer2_outputs(8317) <= (layer1_outputs(9998)) and not (layer1_outputs(1980));
    layer2_outputs(8318) <= (layer1_outputs(9740)) and (layer1_outputs(12394));
    layer2_outputs(8319) <= layer1_outputs(11240);
    layer2_outputs(8320) <= not((layer1_outputs(4989)) and (layer1_outputs(1288)));
    layer2_outputs(8321) <= not(layer1_outputs(7278));
    layer2_outputs(8322) <= layer1_outputs(12682);
    layer2_outputs(8323) <= not(layer1_outputs(6538)) or (layer1_outputs(5674));
    layer2_outputs(8324) <= (layer1_outputs(8742)) and (layer1_outputs(6712));
    layer2_outputs(8325) <= not((layer1_outputs(9179)) xor (layer1_outputs(8076)));
    layer2_outputs(8326) <= layer1_outputs(248);
    layer2_outputs(8327) <= layer1_outputs(11136);
    layer2_outputs(8328) <= not(layer1_outputs(10596));
    layer2_outputs(8329) <= not(layer1_outputs(7179));
    layer2_outputs(8330) <= (layer1_outputs(10565)) and (layer1_outputs(4785));
    layer2_outputs(8331) <= layer1_outputs(462);
    layer2_outputs(8332) <= not(layer1_outputs(5015));
    layer2_outputs(8333) <= not(layer1_outputs(12437)) or (layer1_outputs(7383));
    layer2_outputs(8334) <= layer1_outputs(11355);
    layer2_outputs(8335) <= not(layer1_outputs(3952));
    layer2_outputs(8336) <= layer1_outputs(9085);
    layer2_outputs(8337) <= layer1_outputs(8524);
    layer2_outputs(8338) <= not(layer1_outputs(8778));
    layer2_outputs(8339) <= (layer1_outputs(1117)) and (layer1_outputs(865));
    layer2_outputs(8340) <= (layer1_outputs(8501)) or (layer1_outputs(8665));
    layer2_outputs(8341) <= layer1_outputs(418);
    layer2_outputs(8342) <= layer1_outputs(887);
    layer2_outputs(8343) <= not((layer1_outputs(7010)) or (layer1_outputs(9333)));
    layer2_outputs(8344) <= layer1_outputs(12660);
    layer2_outputs(8345) <= not(layer1_outputs(8521));
    layer2_outputs(8346) <= not(layer1_outputs(4502)) or (layer1_outputs(8231));
    layer2_outputs(8347) <= layer1_outputs(2672);
    layer2_outputs(8348) <= not(layer1_outputs(3214));
    layer2_outputs(8349) <= not((layer1_outputs(1562)) and (layer1_outputs(1605)));
    layer2_outputs(8350) <= not(layer1_outputs(1122));
    layer2_outputs(8351) <= not(layer1_outputs(11492));
    layer2_outputs(8352) <= (layer1_outputs(4036)) and not (layer1_outputs(1842));
    layer2_outputs(8353) <= not(layer1_outputs(11281)) or (layer1_outputs(12117));
    layer2_outputs(8354) <= not(layer1_outputs(3862));
    layer2_outputs(8355) <= (layer1_outputs(10037)) and (layer1_outputs(3944));
    layer2_outputs(8356) <= not((layer1_outputs(9933)) and (layer1_outputs(5470)));
    layer2_outputs(8357) <= not((layer1_outputs(4059)) and (layer1_outputs(10359)));
    layer2_outputs(8358) <= layer1_outputs(9265);
    layer2_outputs(8359) <= not(layer1_outputs(12642));
    layer2_outputs(8360) <= not(layer1_outputs(3096)) or (layer1_outputs(745));
    layer2_outputs(8361) <= not((layer1_outputs(9926)) or (layer1_outputs(3581)));
    layer2_outputs(8362) <= '0';
    layer2_outputs(8363) <= (layer1_outputs(12737)) and not (layer1_outputs(10988));
    layer2_outputs(8364) <= layer1_outputs(10045);
    layer2_outputs(8365) <= layer1_outputs(11410);
    layer2_outputs(8366) <= not(layer1_outputs(11404));
    layer2_outputs(8367) <= not(layer1_outputs(4672));
    layer2_outputs(8368) <= not((layer1_outputs(10352)) or (layer1_outputs(10100)));
    layer2_outputs(8369) <= not(layer1_outputs(3300));
    layer2_outputs(8370) <= not(layer1_outputs(4598));
    layer2_outputs(8371) <= not((layer1_outputs(4692)) or (layer1_outputs(4980)));
    layer2_outputs(8372) <= not((layer1_outputs(4045)) or (layer1_outputs(2153)));
    layer2_outputs(8373) <= not((layer1_outputs(9504)) xor (layer1_outputs(11747)));
    layer2_outputs(8374) <= layer1_outputs(855);
    layer2_outputs(8375) <= (layer1_outputs(651)) or (layer1_outputs(9016));
    layer2_outputs(8376) <= not((layer1_outputs(9843)) xor (layer1_outputs(10208)));
    layer2_outputs(8377) <= not((layer1_outputs(652)) xor (layer1_outputs(5328)));
    layer2_outputs(8378) <= not((layer1_outputs(299)) and (layer1_outputs(6936)));
    layer2_outputs(8379) <= (layer1_outputs(6226)) and not (layer1_outputs(5805));
    layer2_outputs(8380) <= not(layer1_outputs(3928));
    layer2_outputs(8381) <= layer1_outputs(1055);
    layer2_outputs(8382) <= not(layer1_outputs(1897));
    layer2_outputs(8383) <= layer1_outputs(7715);
    layer2_outputs(8384) <= layer1_outputs(7267);
    layer2_outputs(8385) <= layer1_outputs(1955);
    layer2_outputs(8386) <= (layer1_outputs(11104)) or (layer1_outputs(5500));
    layer2_outputs(8387) <= not(layer1_outputs(10050)) or (layer1_outputs(11077));
    layer2_outputs(8388) <= layer1_outputs(12090);
    layer2_outputs(8389) <= (layer1_outputs(2352)) xor (layer1_outputs(702));
    layer2_outputs(8390) <= not(layer1_outputs(10953));
    layer2_outputs(8391) <= not(layer1_outputs(10930)) or (layer1_outputs(9741));
    layer2_outputs(8392) <= not(layer1_outputs(996));
    layer2_outputs(8393) <= not((layer1_outputs(3466)) or (layer1_outputs(9765)));
    layer2_outputs(8394) <= (layer1_outputs(2329)) and not (layer1_outputs(11447));
    layer2_outputs(8395) <= not(layer1_outputs(6200));
    layer2_outputs(8396) <= not(layer1_outputs(1325)) or (layer1_outputs(6750));
    layer2_outputs(8397) <= not(layer1_outputs(10192)) or (layer1_outputs(4093));
    layer2_outputs(8398) <= (layer1_outputs(4467)) xor (layer1_outputs(5174));
    layer2_outputs(8399) <= not(layer1_outputs(3314));
    layer2_outputs(8400) <= (layer1_outputs(4829)) xor (layer1_outputs(11995));
    layer2_outputs(8401) <= not(layer1_outputs(2562));
    layer2_outputs(8402) <= not(layer1_outputs(7344));
    layer2_outputs(8403) <= (layer1_outputs(133)) xor (layer1_outputs(4249));
    layer2_outputs(8404) <= not(layer1_outputs(8401));
    layer2_outputs(8405) <= layer1_outputs(628);
    layer2_outputs(8406) <= not(layer1_outputs(2315)) or (layer1_outputs(6224));
    layer2_outputs(8407) <= layer1_outputs(2345);
    layer2_outputs(8408) <= not((layer1_outputs(2605)) or (layer1_outputs(12166)));
    layer2_outputs(8409) <= layer1_outputs(11056);
    layer2_outputs(8410) <= (layer1_outputs(3249)) or (layer1_outputs(5612));
    layer2_outputs(8411) <= layer1_outputs(7903);
    layer2_outputs(8412) <= (layer1_outputs(12290)) xor (layer1_outputs(11779));
    layer2_outputs(8413) <= not(layer1_outputs(11901));
    layer2_outputs(8414) <= layer1_outputs(1555);
    layer2_outputs(8415) <= (layer1_outputs(4288)) and not (layer1_outputs(9683));
    layer2_outputs(8416) <= layer1_outputs(10346);
    layer2_outputs(8417) <= not((layer1_outputs(5138)) or (layer1_outputs(4507)));
    layer2_outputs(8418) <= not((layer1_outputs(5566)) or (layer1_outputs(8939)));
    layer2_outputs(8419) <= not((layer1_outputs(8363)) and (layer1_outputs(6836)));
    layer2_outputs(8420) <= (layer1_outputs(11252)) xor (layer1_outputs(1942));
    layer2_outputs(8421) <= layer1_outputs(699);
    layer2_outputs(8422) <= (layer1_outputs(11010)) xor (layer1_outputs(11834));
    layer2_outputs(8423) <= not(layer1_outputs(7416)) or (layer1_outputs(9557));
    layer2_outputs(8424) <= not(layer1_outputs(6072)) or (layer1_outputs(130));
    layer2_outputs(8425) <= not(layer1_outputs(3641));
    layer2_outputs(8426) <= layer1_outputs(10575);
    layer2_outputs(8427) <= (layer1_outputs(4265)) and not (layer1_outputs(5588));
    layer2_outputs(8428) <= not((layer1_outputs(8329)) and (layer1_outputs(6976)));
    layer2_outputs(8429) <= (layer1_outputs(6994)) and not (layer1_outputs(7242));
    layer2_outputs(8430) <= (layer1_outputs(5673)) and not (layer1_outputs(1052));
    layer2_outputs(8431) <= not(layer1_outputs(4126));
    layer2_outputs(8432) <= not((layer1_outputs(11491)) or (layer1_outputs(11787)));
    layer2_outputs(8433) <= not(layer1_outputs(5551)) or (layer1_outputs(6202));
    layer2_outputs(8434) <= layer1_outputs(5101);
    layer2_outputs(8435) <= layer1_outputs(1009);
    layer2_outputs(8436) <= '0';
    layer2_outputs(8437) <= layer1_outputs(4090);
    layer2_outputs(8438) <= not(layer1_outputs(1300));
    layer2_outputs(8439) <= not(layer1_outputs(11043));
    layer2_outputs(8440) <= not((layer1_outputs(6801)) or (layer1_outputs(8175)));
    layer2_outputs(8441) <= layer1_outputs(10215);
    layer2_outputs(8442) <= layer1_outputs(12057);
    layer2_outputs(8443) <= not(layer1_outputs(9131));
    layer2_outputs(8444) <= not(layer1_outputs(1470)) or (layer1_outputs(3246));
    layer2_outputs(8445) <= not(layer1_outputs(10321));
    layer2_outputs(8446) <= layer1_outputs(1000);
    layer2_outputs(8447) <= not(layer1_outputs(9154)) or (layer1_outputs(5301));
    layer2_outputs(8448) <= not(layer1_outputs(2829));
    layer2_outputs(8449) <= layer1_outputs(4326);
    layer2_outputs(8450) <= not(layer1_outputs(10938)) or (layer1_outputs(7759));
    layer2_outputs(8451) <= layer1_outputs(11316);
    layer2_outputs(8452) <= (layer1_outputs(12602)) and not (layer1_outputs(6088));
    layer2_outputs(8453) <= not((layer1_outputs(11195)) or (layer1_outputs(10673)));
    layer2_outputs(8454) <= (layer1_outputs(2715)) xor (layer1_outputs(4361));
    layer2_outputs(8455) <= '0';
    layer2_outputs(8456) <= layer1_outputs(2223);
    layer2_outputs(8457) <= (layer1_outputs(1616)) or (layer1_outputs(9971));
    layer2_outputs(8458) <= (layer1_outputs(1937)) and not (layer1_outputs(4716));
    layer2_outputs(8459) <= (layer1_outputs(1610)) xor (layer1_outputs(12542));
    layer2_outputs(8460) <= not(layer1_outputs(4783));
    layer2_outputs(8461) <= not(layer1_outputs(6075));
    layer2_outputs(8462) <= not(layer1_outputs(2370));
    layer2_outputs(8463) <= layer1_outputs(156);
    layer2_outputs(8464) <= layer1_outputs(2795);
    layer2_outputs(8465) <= layer1_outputs(523);
    layer2_outputs(8466) <= layer1_outputs(11321);
    layer2_outputs(8467) <= not(layer1_outputs(1560)) or (layer1_outputs(6430));
    layer2_outputs(8468) <= (layer1_outputs(7636)) and (layer1_outputs(7933));
    layer2_outputs(8469) <= not(layer1_outputs(12476));
    layer2_outputs(8470) <= layer1_outputs(6686);
    layer2_outputs(8471) <= (layer1_outputs(7041)) and (layer1_outputs(3120));
    layer2_outputs(8472) <= not((layer1_outputs(3497)) xor (layer1_outputs(8548)));
    layer2_outputs(8473) <= layer1_outputs(3449);
    layer2_outputs(8474) <= not(layer1_outputs(7730)) or (layer1_outputs(2520));
    layer2_outputs(8475) <= (layer1_outputs(10392)) or (layer1_outputs(3153));
    layer2_outputs(8476) <= layer1_outputs(530);
    layer2_outputs(8477) <= not(layer1_outputs(5190)) or (layer1_outputs(12225));
    layer2_outputs(8478) <= (layer1_outputs(6937)) and not (layer1_outputs(11208));
    layer2_outputs(8479) <= not((layer1_outputs(6199)) xor (layer1_outputs(11709)));
    layer2_outputs(8480) <= (layer1_outputs(512)) and not (layer1_outputs(2893));
    layer2_outputs(8481) <= not(layer1_outputs(2070));
    layer2_outputs(8482) <= (layer1_outputs(5759)) and (layer1_outputs(3897));
    layer2_outputs(8483) <= (layer1_outputs(1732)) and (layer1_outputs(149));
    layer2_outputs(8484) <= not((layer1_outputs(6442)) xor (layer1_outputs(7823)));
    layer2_outputs(8485) <= (layer1_outputs(7795)) xor (layer1_outputs(3995));
    layer2_outputs(8486) <= (layer1_outputs(6621)) and not (layer1_outputs(5269));
    layer2_outputs(8487) <= not((layer1_outputs(9525)) or (layer1_outputs(35)));
    layer2_outputs(8488) <= layer1_outputs(9295);
    layer2_outputs(8489) <= not((layer1_outputs(11413)) or (layer1_outputs(7206)));
    layer2_outputs(8490) <= (layer1_outputs(3319)) and not (layer1_outputs(10148));
    layer2_outputs(8491) <= not(layer1_outputs(2042));
    layer2_outputs(8492) <= not(layer1_outputs(4903));
    layer2_outputs(8493) <= layer1_outputs(8467);
    layer2_outputs(8494) <= (layer1_outputs(9096)) and not (layer1_outputs(9985));
    layer2_outputs(8495) <= layer1_outputs(10354);
    layer2_outputs(8496) <= not(layer1_outputs(7085));
    layer2_outputs(8497) <= not(layer1_outputs(762));
    layer2_outputs(8498) <= not(layer1_outputs(5740)) or (layer1_outputs(1336));
    layer2_outputs(8499) <= (layer1_outputs(7611)) and (layer1_outputs(1158));
    layer2_outputs(8500) <= (layer1_outputs(1265)) or (layer1_outputs(5672));
    layer2_outputs(8501) <= layer1_outputs(8707);
    layer2_outputs(8502) <= layer1_outputs(9445);
    layer2_outputs(8503) <= not((layer1_outputs(588)) xor (layer1_outputs(3090)));
    layer2_outputs(8504) <= (layer1_outputs(12621)) or (layer1_outputs(12396));
    layer2_outputs(8505) <= (layer1_outputs(10414)) xor (layer1_outputs(2817));
    layer2_outputs(8506) <= (layer1_outputs(3845)) xor (layer1_outputs(11111));
    layer2_outputs(8507) <= not(layer1_outputs(9830)) or (layer1_outputs(3158));
    layer2_outputs(8508) <= layer1_outputs(11804);
    layer2_outputs(8509) <= (layer1_outputs(4558)) xor (layer1_outputs(11920));
    layer2_outputs(8510) <= not(layer1_outputs(4963));
    layer2_outputs(8511) <= not(layer1_outputs(2049)) or (layer1_outputs(9122));
    layer2_outputs(8512) <= (layer1_outputs(2790)) and not (layer1_outputs(4455));
    layer2_outputs(8513) <= (layer1_outputs(1185)) and (layer1_outputs(6797));
    layer2_outputs(8514) <= (layer1_outputs(863)) xor (layer1_outputs(7689));
    layer2_outputs(8515) <= layer1_outputs(10903);
    layer2_outputs(8516) <= not(layer1_outputs(6112));
    layer2_outputs(8517) <= not(layer1_outputs(4927)) or (layer1_outputs(11811));
    layer2_outputs(8518) <= not(layer1_outputs(12618));
    layer2_outputs(8519) <= not(layer1_outputs(9497));
    layer2_outputs(8520) <= not((layer1_outputs(6758)) and (layer1_outputs(6919)));
    layer2_outputs(8521) <= layer1_outputs(6091);
    layer2_outputs(8522) <= layer1_outputs(1444);
    layer2_outputs(8523) <= (layer1_outputs(8203)) and (layer1_outputs(415));
    layer2_outputs(8524) <= '0';
    layer2_outputs(8525) <= not(layer1_outputs(6587)) or (layer1_outputs(4325));
    layer2_outputs(8526) <= (layer1_outputs(389)) or (layer1_outputs(5060));
    layer2_outputs(8527) <= (layer1_outputs(4932)) and not (layer1_outputs(3615));
    layer2_outputs(8528) <= layer1_outputs(10526);
    layer2_outputs(8529) <= (layer1_outputs(1928)) and not (layer1_outputs(57));
    layer2_outputs(8530) <= not((layer1_outputs(8975)) xor (layer1_outputs(3966)));
    layer2_outputs(8531) <= (layer1_outputs(6836)) and not (layer1_outputs(1822));
    layer2_outputs(8532) <= not(layer1_outputs(10932));
    layer2_outputs(8533) <= not(layer1_outputs(2912)) or (layer1_outputs(2075));
    layer2_outputs(8534) <= layer1_outputs(8868);
    layer2_outputs(8535) <= not(layer1_outputs(4669));
    layer2_outputs(8536) <= not(layer1_outputs(4424));
    layer2_outputs(8537) <= layer1_outputs(5664);
    layer2_outputs(8538) <= (layer1_outputs(635)) or (layer1_outputs(12440));
    layer2_outputs(8539) <= layer1_outputs(12347);
    layer2_outputs(8540) <= layer1_outputs(7905);
    layer2_outputs(8541) <= not(layer1_outputs(1915));
    layer2_outputs(8542) <= layer1_outputs(1737);
    layer2_outputs(8543) <= not(layer1_outputs(710));
    layer2_outputs(8544) <= (layer1_outputs(5580)) or (layer1_outputs(7232));
    layer2_outputs(8545) <= not((layer1_outputs(5686)) or (layer1_outputs(4255)));
    layer2_outputs(8546) <= layer1_outputs(6335);
    layer2_outputs(8547) <= (layer1_outputs(7514)) xor (layer1_outputs(6652));
    layer2_outputs(8548) <= not(layer1_outputs(3278)) or (layer1_outputs(9162));
    layer2_outputs(8549) <= not(layer1_outputs(1635));
    layer2_outputs(8550) <= layer1_outputs(663);
    layer2_outputs(8551) <= (layer1_outputs(12547)) and not (layer1_outputs(3750));
    layer2_outputs(8552) <= not(layer1_outputs(726));
    layer2_outputs(8553) <= (layer1_outputs(782)) xor (layer1_outputs(5494));
    layer2_outputs(8554) <= not(layer1_outputs(8313));
    layer2_outputs(8555) <= (layer1_outputs(9322)) and not (layer1_outputs(7941));
    layer2_outputs(8556) <= not(layer1_outputs(1496));
    layer2_outputs(8557) <= layer1_outputs(4415);
    layer2_outputs(8558) <= layer1_outputs(8114);
    layer2_outputs(8559) <= (layer1_outputs(7183)) and not (layer1_outputs(3568));
    layer2_outputs(8560) <= (layer1_outputs(5118)) or (layer1_outputs(9549));
    layer2_outputs(8561) <= not(layer1_outputs(9290));
    layer2_outputs(8562) <= not(layer1_outputs(11437));
    layer2_outputs(8563) <= not(layer1_outputs(5768));
    layer2_outputs(8564) <= (layer1_outputs(3573)) and not (layer1_outputs(7533));
    layer2_outputs(8565) <= not((layer1_outputs(1715)) and (layer1_outputs(6484)));
    layer2_outputs(8566) <= layer1_outputs(2699);
    layer2_outputs(8567) <= (layer1_outputs(8712)) xor (layer1_outputs(621));
    layer2_outputs(8568) <= (layer1_outputs(113)) and (layer1_outputs(5763));
    layer2_outputs(8569) <= not(layer1_outputs(4719)) or (layer1_outputs(9783));
    layer2_outputs(8570) <= not((layer1_outputs(8517)) xor (layer1_outputs(9675)));
    layer2_outputs(8571) <= (layer1_outputs(654)) xor (layer1_outputs(5794));
    layer2_outputs(8572) <= (layer1_outputs(4510)) xor (layer1_outputs(4350));
    layer2_outputs(8573) <= not(layer1_outputs(4245));
    layer2_outputs(8574) <= not((layer1_outputs(1399)) xor (layer1_outputs(9902)));
    layer2_outputs(8575) <= not(layer1_outputs(11760));
    layer2_outputs(8576) <= (layer1_outputs(7658)) and (layer1_outputs(749));
    layer2_outputs(8577) <= not((layer1_outputs(1141)) and (layer1_outputs(9890)));
    layer2_outputs(8578) <= layer1_outputs(4043);
    layer2_outputs(8579) <= (layer1_outputs(5510)) and not (layer1_outputs(6139));
    layer2_outputs(8580) <= layer1_outputs(7734);
    layer2_outputs(8581) <= not(layer1_outputs(11219));
    layer2_outputs(8582) <= layer1_outputs(10772);
    layer2_outputs(8583) <= (layer1_outputs(11384)) or (layer1_outputs(8073));
    layer2_outputs(8584) <= not((layer1_outputs(683)) xor (layer1_outputs(7835)));
    layer2_outputs(8585) <= not(layer1_outputs(6303));
    layer2_outputs(8586) <= layer1_outputs(756);
    layer2_outputs(8587) <= (layer1_outputs(10129)) and (layer1_outputs(1748));
    layer2_outputs(8588) <= (layer1_outputs(12197)) and not (layer1_outputs(6843));
    layer2_outputs(8589) <= (layer1_outputs(2697)) and not (layer1_outputs(7244));
    layer2_outputs(8590) <= not(layer1_outputs(2808));
    layer2_outputs(8591) <= not(layer1_outputs(1001));
    layer2_outputs(8592) <= (layer1_outputs(1643)) and not (layer1_outputs(9608));
    layer2_outputs(8593) <= (layer1_outputs(6982)) and not (layer1_outputs(6803));
    layer2_outputs(8594) <= layer1_outputs(6069);
    layer2_outputs(8595) <= layer1_outputs(6017);
    layer2_outputs(8596) <= not(layer1_outputs(1921));
    layer2_outputs(8597) <= (layer1_outputs(12202)) xor (layer1_outputs(2342));
    layer2_outputs(8598) <= not((layer1_outputs(11432)) and (layer1_outputs(9584)));
    layer2_outputs(8599) <= not(layer1_outputs(11140)) or (layer1_outputs(3674));
    layer2_outputs(8600) <= (layer1_outputs(2931)) and (layer1_outputs(7351));
    layer2_outputs(8601) <= layer1_outputs(4466);
    layer2_outputs(8602) <= not((layer1_outputs(5718)) or (layer1_outputs(5284)));
    layer2_outputs(8603) <= not(layer1_outputs(6554)) or (layer1_outputs(212));
    layer2_outputs(8604) <= not(layer1_outputs(4345));
    layer2_outputs(8605) <= not(layer1_outputs(10039));
    layer2_outputs(8606) <= not((layer1_outputs(10844)) or (layer1_outputs(1111)));
    layer2_outputs(8607) <= not(layer1_outputs(11680));
    layer2_outputs(8608) <= (layer1_outputs(11142)) and not (layer1_outputs(5460));
    layer2_outputs(8609) <= layer1_outputs(373);
    layer2_outputs(8610) <= not((layer1_outputs(3976)) or (layer1_outputs(6639)));
    layer2_outputs(8611) <= not(layer1_outputs(314));
    layer2_outputs(8612) <= not(layer1_outputs(4000));
    layer2_outputs(8613) <= not(layer1_outputs(1171));
    layer2_outputs(8614) <= (layer1_outputs(7614)) or (layer1_outputs(11341));
    layer2_outputs(8615) <= layer1_outputs(8082);
    layer2_outputs(8616) <= layer1_outputs(10822);
    layer2_outputs(8617) <= (layer1_outputs(11912)) or (layer1_outputs(9763));
    layer2_outputs(8618) <= (layer1_outputs(11720)) and (layer1_outputs(3564));
    layer2_outputs(8619) <= not((layer1_outputs(10214)) and (layer1_outputs(4914)));
    layer2_outputs(8620) <= not(layer1_outputs(1816));
    layer2_outputs(8621) <= (layer1_outputs(4252)) and (layer1_outputs(11894));
    layer2_outputs(8622) <= not(layer1_outputs(4962));
    layer2_outputs(8623) <= (layer1_outputs(4865)) and (layer1_outputs(6401));
    layer2_outputs(8624) <= not(layer1_outputs(9138)) or (layer1_outputs(3814));
    layer2_outputs(8625) <= not((layer1_outputs(7366)) xor (layer1_outputs(4587)));
    layer2_outputs(8626) <= layer1_outputs(2450);
    layer2_outputs(8627) <= not(layer1_outputs(1229));
    layer2_outputs(8628) <= (layer1_outputs(4929)) and not (layer1_outputs(3888));
    layer2_outputs(8629) <= '0';
    layer2_outputs(8630) <= layer1_outputs(3108);
    layer2_outputs(8631) <= (layer1_outputs(984)) or (layer1_outputs(3547));
    layer2_outputs(8632) <= not(layer1_outputs(591));
    layer2_outputs(8633) <= layer1_outputs(8067);
    layer2_outputs(8634) <= not(layer1_outputs(9665));
    layer2_outputs(8635) <= (layer1_outputs(1851)) and (layer1_outputs(3713));
    layer2_outputs(8636) <= layer1_outputs(7501);
    layer2_outputs(8637) <= layer1_outputs(10931);
    layer2_outputs(8638) <= (layer1_outputs(4721)) or (layer1_outputs(1983));
    layer2_outputs(8639) <= layer1_outputs(7949);
    layer2_outputs(8640) <= not(layer1_outputs(913)) or (layer1_outputs(8132));
    layer2_outputs(8641) <= (layer1_outputs(1960)) or (layer1_outputs(2667));
    layer2_outputs(8642) <= layer1_outputs(6394);
    layer2_outputs(8643) <= (layer1_outputs(12318)) and not (layer1_outputs(7459));
    layer2_outputs(8644) <= (layer1_outputs(1398)) and not (layer1_outputs(3894));
    layer2_outputs(8645) <= layer1_outputs(5969);
    layer2_outputs(8646) <= layer1_outputs(2946);
    layer2_outputs(8647) <= (layer1_outputs(5772)) xor (layer1_outputs(7014));
    layer2_outputs(8648) <= (layer1_outputs(448)) and not (layer1_outputs(178));
    layer2_outputs(8649) <= layer1_outputs(2638);
    layer2_outputs(8650) <= not(layer1_outputs(4928));
    layer2_outputs(8651) <= not((layer1_outputs(2210)) and (layer1_outputs(6943)));
    layer2_outputs(8652) <= not((layer1_outputs(3636)) and (layer1_outputs(5692)));
    layer2_outputs(8653) <= (layer1_outputs(3306)) and (layer1_outputs(7250));
    layer2_outputs(8654) <= layer1_outputs(6108);
    layer2_outputs(8655) <= not((layer1_outputs(5954)) xor (layer1_outputs(8389)));
    layer2_outputs(8656) <= (layer1_outputs(12040)) and not (layer1_outputs(9697));
    layer2_outputs(8657) <= not((layer1_outputs(8835)) xor (layer1_outputs(3271)));
    layer2_outputs(8658) <= layer1_outputs(10581);
    layer2_outputs(8659) <= '1';
    layer2_outputs(8660) <= not((layer1_outputs(5335)) and (layer1_outputs(6141)));
    layer2_outputs(8661) <= not(layer1_outputs(11662));
    layer2_outputs(8662) <= (layer1_outputs(4412)) and not (layer1_outputs(4771));
    layer2_outputs(8663) <= '0';
    layer2_outputs(8664) <= not(layer1_outputs(3719));
    layer2_outputs(8665) <= layer1_outputs(12619);
    layer2_outputs(8666) <= not(layer1_outputs(8381)) or (layer1_outputs(7271));
    layer2_outputs(8667) <= layer1_outputs(5237);
    layer2_outputs(8668) <= not(layer1_outputs(11372)) or (layer1_outputs(9801));
    layer2_outputs(8669) <= not((layer1_outputs(6443)) xor (layer1_outputs(10818)));
    layer2_outputs(8670) <= not((layer1_outputs(8195)) xor (layer1_outputs(577)));
    layer2_outputs(8671) <= not(layer1_outputs(9108)) or (layer1_outputs(3648));
    layer2_outputs(8672) <= layer1_outputs(12370);
    layer2_outputs(8673) <= (layer1_outputs(12726)) and not (layer1_outputs(2840));
    layer2_outputs(8674) <= not((layer1_outputs(677)) or (layer1_outputs(6365)));
    layer2_outputs(8675) <= not(layer1_outputs(4749)) or (layer1_outputs(2567));
    layer2_outputs(8676) <= (layer1_outputs(10264)) xor (layer1_outputs(8100));
    layer2_outputs(8677) <= not((layer1_outputs(9171)) or (layer1_outputs(3769)));
    layer2_outputs(8678) <= not((layer1_outputs(3642)) xor (layer1_outputs(879)));
    layer2_outputs(8679) <= not(layer1_outputs(12386));
    layer2_outputs(8680) <= layer1_outputs(7419);
    layer2_outputs(8681) <= not(layer1_outputs(11929));
    layer2_outputs(8682) <= (layer1_outputs(4261)) and not (layer1_outputs(2952));
    layer2_outputs(8683) <= (layer1_outputs(3802)) xor (layer1_outputs(1468));
    layer2_outputs(8684) <= layer1_outputs(5292);
    layer2_outputs(8685) <= layer1_outputs(12412);
    layer2_outputs(8686) <= layer1_outputs(1342);
    layer2_outputs(8687) <= (layer1_outputs(11986)) or (layer1_outputs(11429));
    layer2_outputs(8688) <= not(layer1_outputs(5189));
    layer2_outputs(8689) <= not((layer1_outputs(10876)) or (layer1_outputs(65)));
    layer2_outputs(8690) <= not(layer1_outputs(2099));
    layer2_outputs(8691) <= not(layer1_outputs(8336)) or (layer1_outputs(9470));
    layer2_outputs(8692) <= layer1_outputs(7789);
    layer2_outputs(8693) <= not(layer1_outputs(6948));
    layer2_outputs(8694) <= not(layer1_outputs(1240));
    layer2_outputs(8695) <= (layer1_outputs(1179)) xor (layer1_outputs(4418));
    layer2_outputs(8696) <= (layer1_outputs(2290)) and (layer1_outputs(7152));
    layer2_outputs(8697) <= layer1_outputs(6291);
    layer2_outputs(8698) <= not((layer1_outputs(9481)) and (layer1_outputs(11375)));
    layer2_outputs(8699) <= (layer1_outputs(9400)) and not (layer1_outputs(8990));
    layer2_outputs(8700) <= (layer1_outputs(9564)) xor (layer1_outputs(3072));
    layer2_outputs(8701) <= (layer1_outputs(272)) xor (layer1_outputs(9473));
    layer2_outputs(8702) <= '1';
    layer2_outputs(8703) <= (layer1_outputs(5970)) or (layer1_outputs(10516));
    layer2_outputs(8704) <= not(layer1_outputs(10195)) or (layer1_outputs(8522));
    layer2_outputs(8705) <= not(layer1_outputs(6329)) or (layer1_outputs(9226));
    layer2_outputs(8706) <= not((layer1_outputs(10606)) xor (layer1_outputs(4605)));
    layer2_outputs(8707) <= (layer1_outputs(4895)) and (layer1_outputs(9113));
    layer2_outputs(8708) <= layer1_outputs(6910);
    layer2_outputs(8709) <= (layer1_outputs(5161)) or (layer1_outputs(2025));
    layer2_outputs(8710) <= not(layer1_outputs(6788));
    layer2_outputs(8711) <= layer1_outputs(864);
    layer2_outputs(8712) <= (layer1_outputs(3295)) or (layer1_outputs(11068));
    layer2_outputs(8713) <= (layer1_outputs(2940)) and not (layer1_outputs(568));
    layer2_outputs(8714) <= layer1_outputs(2781);
    layer2_outputs(8715) <= '1';
    layer2_outputs(8716) <= (layer1_outputs(6037)) or (layer1_outputs(4905));
    layer2_outputs(8717) <= not(layer1_outputs(4015));
    layer2_outputs(8718) <= not(layer1_outputs(17));
    layer2_outputs(8719) <= (layer1_outputs(9690)) and not (layer1_outputs(10279));
    layer2_outputs(8720) <= layer1_outputs(1685);
    layer2_outputs(8721) <= not((layer1_outputs(8421)) and (layer1_outputs(8123)));
    layer2_outputs(8722) <= not(layer1_outputs(559)) or (layer1_outputs(10294));
    layer2_outputs(8723) <= not(layer1_outputs(7872));
    layer2_outputs(8724) <= layer1_outputs(6128);
    layer2_outputs(8725) <= not((layer1_outputs(9561)) or (layer1_outputs(509)));
    layer2_outputs(8726) <= not(layer1_outputs(5345)) or (layer1_outputs(9083));
    layer2_outputs(8727) <= not(layer1_outputs(5217));
    layer2_outputs(8728) <= not((layer1_outputs(3614)) or (layer1_outputs(10268)));
    layer2_outputs(8729) <= (layer1_outputs(1714)) xor (layer1_outputs(4061));
    layer2_outputs(8730) <= not(layer1_outputs(3859)) or (layer1_outputs(5962));
    layer2_outputs(8731) <= layer1_outputs(1255);
    layer2_outputs(8732) <= not((layer1_outputs(11445)) xor (layer1_outputs(12614)));
    layer2_outputs(8733) <= layer1_outputs(4992);
    layer2_outputs(8734) <= not(layer1_outputs(2702));
    layer2_outputs(8735) <= (layer1_outputs(4591)) and not (layer1_outputs(5320));
    layer2_outputs(8736) <= not((layer1_outputs(5571)) or (layer1_outputs(11970)));
    layer2_outputs(8737) <= (layer1_outputs(5775)) and not (layer1_outputs(3505));
    layer2_outputs(8738) <= (layer1_outputs(436)) xor (layer1_outputs(10891));
    layer2_outputs(8739) <= not(layer1_outputs(4413));
    layer2_outputs(8740) <= (layer1_outputs(3907)) and not (layer1_outputs(8424));
    layer2_outputs(8741) <= not((layer1_outputs(1840)) xor (layer1_outputs(10924)));
    layer2_outputs(8742) <= not(layer1_outputs(6334));
    layer2_outputs(8743) <= (layer1_outputs(8962)) and (layer1_outputs(8845));
    layer2_outputs(8744) <= not((layer1_outputs(6098)) and (layer1_outputs(3481)));
    layer2_outputs(8745) <= layer1_outputs(4017);
    layer2_outputs(8746) <= layer1_outputs(3069);
    layer2_outputs(8747) <= layer1_outputs(3708);
    layer2_outputs(8748) <= not(layer1_outputs(7759));
    layer2_outputs(8749) <= (layer1_outputs(584)) and not (layer1_outputs(9924));
    layer2_outputs(8750) <= (layer1_outputs(4975)) or (layer1_outputs(5182));
    layer2_outputs(8751) <= (layer1_outputs(1744)) and not (layer1_outputs(1995));
    layer2_outputs(8752) <= not(layer1_outputs(2421));
    layer2_outputs(8753) <= not(layer1_outputs(6360)) or (layer1_outputs(6754));
    layer2_outputs(8754) <= (layer1_outputs(4725)) and (layer1_outputs(1987));
    layer2_outputs(8755) <= not(layer1_outputs(7027)) or (layer1_outputs(1244));
    layer2_outputs(8756) <= not(layer1_outputs(781));
    layer2_outputs(8757) <= not((layer1_outputs(5428)) or (layer1_outputs(2806)));
    layer2_outputs(8758) <= layer1_outputs(936);
    layer2_outputs(8759) <= not(layer1_outputs(1637));
    layer2_outputs(8760) <= (layer1_outputs(11971)) and not (layer1_outputs(3448));
    layer2_outputs(8761) <= '1';
    layer2_outputs(8762) <= (layer1_outputs(5681)) xor (layer1_outputs(1361));
    layer2_outputs(8763) <= (layer1_outputs(10016)) and (layer1_outputs(10200));
    layer2_outputs(8764) <= layer1_outputs(12107);
    layer2_outputs(8765) <= (layer1_outputs(7347)) and not (layer1_outputs(10149));
    layer2_outputs(8766) <= layer1_outputs(5336);
    layer2_outputs(8767) <= layer1_outputs(10833);
    layer2_outputs(8768) <= not(layer1_outputs(1269)) or (layer1_outputs(9599));
    layer2_outputs(8769) <= not((layer1_outputs(7243)) and (layer1_outputs(5524)));
    layer2_outputs(8770) <= layer1_outputs(7582);
    layer2_outputs(8771) <= (layer1_outputs(2846)) and (layer1_outputs(4867));
    layer2_outputs(8772) <= not((layer1_outputs(6765)) xor (layer1_outputs(11741)));
    layer2_outputs(8773) <= layer1_outputs(11077);
    layer2_outputs(8774) <= not(layer1_outputs(2296));
    layer2_outputs(8775) <= (layer1_outputs(7029)) and not (layer1_outputs(5931));
    layer2_outputs(8776) <= (layer1_outputs(4178)) and (layer1_outputs(735));
    layer2_outputs(8777) <= not(layer1_outputs(12773)) or (layer1_outputs(779));
    layer2_outputs(8778) <= (layer1_outputs(6536)) or (layer1_outputs(7237));
    layer2_outputs(8779) <= not(layer1_outputs(12400)) or (layer1_outputs(4147));
    layer2_outputs(8780) <= (layer1_outputs(7929)) or (layer1_outputs(4967));
    layer2_outputs(8781) <= (layer1_outputs(2496)) and not (layer1_outputs(6956));
    layer2_outputs(8782) <= not((layer1_outputs(2947)) or (layer1_outputs(10026)));
    layer2_outputs(8783) <= (layer1_outputs(8287)) and not (layer1_outputs(6818));
    layer2_outputs(8784) <= (layer1_outputs(6526)) and (layer1_outputs(4327));
    layer2_outputs(8785) <= layer1_outputs(3652);
    layer2_outputs(8786) <= layer1_outputs(12099);
    layer2_outputs(8787) <= not(layer1_outputs(1202));
    layer2_outputs(8788) <= layer1_outputs(9303);
    layer2_outputs(8789) <= not(layer1_outputs(5597));
    layer2_outputs(8790) <= not(layer1_outputs(8228)) or (layer1_outputs(9770));
    layer2_outputs(8791) <= not(layer1_outputs(2407));
    layer2_outputs(8792) <= not(layer1_outputs(9));
    layer2_outputs(8793) <= not((layer1_outputs(2503)) and (layer1_outputs(2122)));
    layer2_outputs(8794) <= layer1_outputs(1779);
    layer2_outputs(8795) <= (layer1_outputs(1394)) or (layer1_outputs(3675));
    layer2_outputs(8796) <= layer1_outputs(1819);
    layer2_outputs(8797) <= not(layer1_outputs(5488));
    layer2_outputs(8798) <= not((layer1_outputs(11579)) and (layer1_outputs(3197)));
    layer2_outputs(8799) <= not(layer1_outputs(10112)) or (layer1_outputs(4266));
    layer2_outputs(8800) <= (layer1_outputs(7160)) xor (layer1_outputs(4882));
    layer2_outputs(8801) <= not(layer1_outputs(460));
    layer2_outputs(8802) <= (layer1_outputs(8870)) xor (layer1_outputs(6658));
    layer2_outputs(8803) <= (layer1_outputs(5421)) and not (layer1_outputs(2264));
    layer2_outputs(8804) <= layer1_outputs(2128);
    layer2_outputs(8805) <= (layer1_outputs(10960)) xor (layer1_outputs(11582));
    layer2_outputs(8806) <= layer1_outputs(7726);
    layer2_outputs(8807) <= layer1_outputs(12248);
    layer2_outputs(8808) <= not(layer1_outputs(3514));
    layer2_outputs(8809) <= (layer1_outputs(11055)) xor (layer1_outputs(9979));
    layer2_outputs(8810) <= (layer1_outputs(7959)) xor (layer1_outputs(9736));
    layer2_outputs(8811) <= (layer1_outputs(5758)) or (layer1_outputs(12116));
    layer2_outputs(8812) <= not((layer1_outputs(10512)) xor (layer1_outputs(10637)));
    layer2_outputs(8813) <= not((layer1_outputs(737)) xor (layer1_outputs(10662)));
    layer2_outputs(8814) <= (layer1_outputs(7048)) or (layer1_outputs(1890));
    layer2_outputs(8815) <= not((layer1_outputs(6720)) xor (layer1_outputs(12271)));
    layer2_outputs(8816) <= not(layer1_outputs(10093)) or (layer1_outputs(6472));
    layer2_outputs(8817) <= layer1_outputs(5603);
    layer2_outputs(8818) <= not((layer1_outputs(10395)) xor (layer1_outputs(3873)));
    layer2_outputs(8819) <= not(layer1_outputs(3241));
    layer2_outputs(8820) <= layer1_outputs(11655);
    layer2_outputs(8821) <= not(layer1_outputs(739)) or (layer1_outputs(9180));
    layer2_outputs(8822) <= layer1_outputs(8504);
    layer2_outputs(8823) <= not(layer1_outputs(163));
    layer2_outputs(8824) <= not((layer1_outputs(12353)) or (layer1_outputs(11041)));
    layer2_outputs(8825) <= (layer1_outputs(4232)) and (layer1_outputs(2940));
    layer2_outputs(8826) <= not((layer1_outputs(6087)) xor (layer1_outputs(2921)));
    layer2_outputs(8827) <= not(layer1_outputs(1144));
    layer2_outputs(8828) <= not((layer1_outputs(8547)) xor (layer1_outputs(9652)));
    layer2_outputs(8829) <= (layer1_outputs(11511)) and (layer1_outputs(859));
    layer2_outputs(8830) <= not((layer1_outputs(8230)) and (layer1_outputs(4379)));
    layer2_outputs(8831) <= not(layer1_outputs(5333));
    layer2_outputs(8832) <= layer1_outputs(11705);
    layer2_outputs(8833) <= layer1_outputs(3142);
    layer2_outputs(8834) <= layer1_outputs(9365);
    layer2_outputs(8835) <= not(layer1_outputs(6068));
    layer2_outputs(8836) <= not((layer1_outputs(4785)) and (layer1_outputs(9745)));
    layer2_outputs(8837) <= not(layer1_outputs(660));
    layer2_outputs(8838) <= layer1_outputs(112);
    layer2_outputs(8839) <= not(layer1_outputs(11005));
    layer2_outputs(8840) <= not(layer1_outputs(2645)) or (layer1_outputs(3574));
    layer2_outputs(8841) <= not(layer1_outputs(11459));
    layer2_outputs(8842) <= (layer1_outputs(2186)) and not (layer1_outputs(897));
    layer2_outputs(8843) <= layer1_outputs(325);
    layer2_outputs(8844) <= (layer1_outputs(9258)) and (layer1_outputs(7439));
    layer2_outputs(8845) <= not(layer1_outputs(6039));
    layer2_outputs(8846) <= (layer1_outputs(9670)) and (layer1_outputs(7409));
    layer2_outputs(8847) <= not(layer1_outputs(6042)) or (layer1_outputs(1321));
    layer2_outputs(8848) <= not(layer1_outputs(7217));
    layer2_outputs(8849) <= not(layer1_outputs(6904));
    layer2_outputs(8850) <= not(layer1_outputs(1546));
    layer2_outputs(8851) <= (layer1_outputs(6603)) xor (layer1_outputs(4973));
    layer2_outputs(8852) <= layer1_outputs(3118);
    layer2_outputs(8853) <= layer1_outputs(2492);
    layer2_outputs(8854) <= (layer1_outputs(7748)) or (layer1_outputs(562));
    layer2_outputs(8855) <= not((layer1_outputs(12358)) xor (layer1_outputs(1274)));
    layer2_outputs(8856) <= not(layer1_outputs(5193)) or (layer1_outputs(6676));
    layer2_outputs(8857) <= layer1_outputs(1847);
    layer2_outputs(8858) <= not(layer1_outputs(5370));
    layer2_outputs(8859) <= layer1_outputs(6465);
    layer2_outputs(8860) <= not((layer1_outputs(3179)) xor (layer1_outputs(12630)));
    layer2_outputs(8861) <= '1';
    layer2_outputs(8862) <= not((layer1_outputs(11431)) and (layer1_outputs(11201)));
    layer2_outputs(8863) <= layer1_outputs(8244);
    layer2_outputs(8864) <= not(layer1_outputs(3375));
    layer2_outputs(8865) <= layer1_outputs(4990);
    layer2_outputs(8866) <= not((layer1_outputs(2908)) or (layer1_outputs(10290)));
    layer2_outputs(8867) <= not((layer1_outputs(10301)) and (layer1_outputs(4642)));
    layer2_outputs(8868) <= (layer1_outputs(2747)) xor (layer1_outputs(11560));
    layer2_outputs(8869) <= (layer1_outputs(12415)) xor (layer1_outputs(8734));
    layer2_outputs(8870) <= not(layer1_outputs(6626)) or (layer1_outputs(1406));
    layer2_outputs(8871) <= layer1_outputs(8709);
    layer2_outputs(8872) <= (layer1_outputs(5499)) and (layer1_outputs(12446));
    layer2_outputs(8873) <= not((layer1_outputs(12392)) xor (layer1_outputs(1397)));
    layer2_outputs(8874) <= (layer1_outputs(193)) xor (layer1_outputs(5208));
    layer2_outputs(8875) <= layer1_outputs(503);
    layer2_outputs(8876) <= (layer1_outputs(2682)) or (layer1_outputs(8382));
    layer2_outputs(8877) <= (layer1_outputs(4543)) and not (layer1_outputs(11435));
    layer2_outputs(8878) <= not(layer1_outputs(7955));
    layer2_outputs(8879) <= (layer1_outputs(9389)) and (layer1_outputs(229));
    layer2_outputs(8880) <= layer1_outputs(2291);
    layer2_outputs(8881) <= not(layer1_outputs(11520));
    layer2_outputs(8882) <= layer1_outputs(6208);
    layer2_outputs(8883) <= not(layer1_outputs(5561));
    layer2_outputs(8884) <= layer1_outputs(9842);
    layer2_outputs(8885) <= not(layer1_outputs(11635));
    layer2_outputs(8886) <= not(layer1_outputs(1988));
    layer2_outputs(8887) <= (layer1_outputs(1166)) and (layer1_outputs(9393));
    layer2_outputs(8888) <= (layer1_outputs(1675)) and not (layer1_outputs(2767));
    layer2_outputs(8889) <= not(layer1_outputs(246));
    layer2_outputs(8890) <= '1';
    layer2_outputs(8891) <= '1';
    layer2_outputs(8892) <= not((layer1_outputs(8031)) and (layer1_outputs(9181)));
    layer2_outputs(8893) <= not(layer1_outputs(4259));
    layer2_outputs(8894) <= (layer1_outputs(9779)) or (layer1_outputs(7091));
    layer2_outputs(8895) <= (layer1_outputs(973)) xor (layer1_outputs(727));
    layer2_outputs(8896) <= (layer1_outputs(688)) or (layer1_outputs(8151));
    layer2_outputs(8897) <= not(layer1_outputs(2751));
    layer2_outputs(8898) <= not(layer1_outputs(648)) or (layer1_outputs(11642));
    layer2_outputs(8899) <= (layer1_outputs(9290)) and not (layer1_outputs(8680));
    layer2_outputs(8900) <= not((layer1_outputs(2826)) xor (layer1_outputs(9586)));
    layer2_outputs(8901) <= (layer1_outputs(5858)) xor (layer1_outputs(3624));
    layer2_outputs(8902) <= (layer1_outputs(5235)) xor (layer1_outputs(6722));
    layer2_outputs(8903) <= not(layer1_outputs(7415));
    layer2_outputs(8904) <= not((layer1_outputs(4939)) xor (layer1_outputs(12585)));
    layer2_outputs(8905) <= not(layer1_outputs(4461));
    layer2_outputs(8906) <= (layer1_outputs(4864)) or (layer1_outputs(4194));
    layer2_outputs(8907) <= layer1_outputs(9771);
    layer2_outputs(8908) <= layer1_outputs(3129);
    layer2_outputs(8909) <= layer1_outputs(4282);
    layer2_outputs(8910) <= not(layer1_outputs(3247)) or (layer1_outputs(5360));
    layer2_outputs(8911) <= layer1_outputs(1281);
    layer2_outputs(8912) <= not((layer1_outputs(12352)) xor (layer1_outputs(3594)));
    layer2_outputs(8913) <= layer1_outputs(11370);
    layer2_outputs(8914) <= (layer1_outputs(73)) and (layer1_outputs(3165));
    layer2_outputs(8915) <= layer1_outputs(6034);
    layer2_outputs(8916) <= (layer1_outputs(3990)) and not (layer1_outputs(10849));
    layer2_outputs(8917) <= not(layer1_outputs(6835));
    layer2_outputs(8918) <= not((layer1_outputs(11053)) and (layer1_outputs(30)));
    layer2_outputs(8919) <= not((layer1_outputs(9440)) and (layer1_outputs(9017)));
    layer2_outputs(8920) <= (layer1_outputs(8573)) xor (layer1_outputs(8720));
    layer2_outputs(8921) <= (layer1_outputs(5204)) xor (layer1_outputs(5236));
    layer2_outputs(8922) <= not(layer1_outputs(8244));
    layer2_outputs(8923) <= not((layer1_outputs(5646)) xor (layer1_outputs(834)));
    layer2_outputs(8924) <= layer1_outputs(6259);
    layer2_outputs(8925) <= layer1_outputs(2684);
    layer2_outputs(8926) <= not((layer1_outputs(3706)) or (layer1_outputs(10918)));
    layer2_outputs(8927) <= not(layer1_outputs(8818));
    layer2_outputs(8928) <= (layer1_outputs(7202)) and not (layer1_outputs(1478));
    layer2_outputs(8929) <= not(layer1_outputs(1668));
    layer2_outputs(8930) <= (layer1_outputs(12104)) and (layer1_outputs(7178));
    layer2_outputs(8931) <= not((layer1_outputs(12123)) xor (layer1_outputs(509)));
    layer2_outputs(8932) <= (layer1_outputs(3738)) xor (layer1_outputs(840));
    layer2_outputs(8933) <= not(layer1_outputs(6011)) or (layer1_outputs(2563));
    layer2_outputs(8934) <= not(layer1_outputs(135)) or (layer1_outputs(2653));
    layer2_outputs(8935) <= not(layer1_outputs(1424));
    layer2_outputs(8936) <= not(layer1_outputs(12540));
    layer2_outputs(8937) <= layer1_outputs(12528);
    layer2_outputs(8938) <= layer1_outputs(11872);
    layer2_outputs(8939) <= not(layer1_outputs(10617));
    layer2_outputs(8940) <= not(layer1_outputs(10853));
    layer2_outputs(8941) <= (layer1_outputs(1374)) xor (layer1_outputs(6204));
    layer2_outputs(8942) <= not(layer1_outputs(6823));
    layer2_outputs(8943) <= layer1_outputs(3074);
    layer2_outputs(8944) <= not(layer1_outputs(2816));
    layer2_outputs(8945) <= (layer1_outputs(7087)) or (layer1_outputs(10764));
    layer2_outputs(8946) <= layer1_outputs(4960);
    layer2_outputs(8947) <= (layer1_outputs(7870)) or (layer1_outputs(10806));
    layer2_outputs(8948) <= not(layer1_outputs(2545)) or (layer1_outputs(1309));
    layer2_outputs(8949) <= not(layer1_outputs(7942));
    layer2_outputs(8950) <= not(layer1_outputs(9742));
    layer2_outputs(8951) <= layer1_outputs(3294);
    layer2_outputs(8952) <= '1';
    layer2_outputs(8953) <= not(layer1_outputs(11548));
    layer2_outputs(8954) <= (layer1_outputs(4529)) and not (layer1_outputs(4525));
    layer2_outputs(8955) <= (layer1_outputs(4529)) xor (layer1_outputs(8554));
    layer2_outputs(8956) <= not(layer1_outputs(6355));
    layer2_outputs(8957) <= not(layer1_outputs(7216)) or (layer1_outputs(6887));
    layer2_outputs(8958) <= not((layer1_outputs(5442)) or (layer1_outputs(5501)));
    layer2_outputs(8959) <= not((layer1_outputs(9691)) or (layer1_outputs(6111)));
    layer2_outputs(8960) <= not(layer1_outputs(4060));
    layer2_outputs(8961) <= not(layer1_outputs(4624));
    layer2_outputs(8962) <= not((layer1_outputs(1122)) or (layer1_outputs(6117)));
    layer2_outputs(8963) <= layer1_outputs(1272);
    layer2_outputs(8964) <= not(layer1_outputs(2558));
    layer2_outputs(8965) <= not(layer1_outputs(5332)) or (layer1_outputs(12790));
    layer2_outputs(8966) <= not((layer1_outputs(11940)) or (layer1_outputs(8514)));
    layer2_outputs(8967) <= not((layer1_outputs(2636)) xor (layer1_outputs(1179)));
    layer2_outputs(8968) <= '1';
    layer2_outputs(8969) <= not(layer1_outputs(11995));
    layer2_outputs(8970) <= (layer1_outputs(12786)) and (layer1_outputs(2709));
    layer2_outputs(8971) <= not(layer1_outputs(9667));
    layer2_outputs(8972) <= not(layer1_outputs(6580));
    layer2_outputs(8973) <= layer1_outputs(4088);
    layer2_outputs(8974) <= (layer1_outputs(7058)) xor (layer1_outputs(9186));
    layer2_outputs(8975) <= layer1_outputs(7924);
    layer2_outputs(8976) <= layer1_outputs(7323);
    layer2_outputs(8977) <= not(layer1_outputs(3779)) or (layer1_outputs(4270));
    layer2_outputs(8978) <= (layer1_outputs(11116)) xor (layer1_outputs(12580));
    layer2_outputs(8979) <= (layer1_outputs(8856)) and not (layer1_outputs(911));
    layer2_outputs(8980) <= not((layer1_outputs(9805)) or (layer1_outputs(2668)));
    layer2_outputs(8981) <= not(layer1_outputs(2983));
    layer2_outputs(8982) <= (layer1_outputs(3856)) and (layer1_outputs(5997));
    layer2_outputs(8983) <= not((layer1_outputs(10620)) or (layer1_outputs(3454)));
    layer2_outputs(8984) <= not(layer1_outputs(3499));
    layer2_outputs(8985) <= not((layer1_outputs(7549)) xor (layer1_outputs(213)));
    layer2_outputs(8986) <= (layer1_outputs(10852)) xor (layer1_outputs(2973));
    layer2_outputs(8987) <= not(layer1_outputs(8192));
    layer2_outputs(8988) <= not(layer1_outputs(3476));
    layer2_outputs(8989) <= not(layer1_outputs(10210)) or (layer1_outputs(4253));
    layer2_outputs(8990) <= not(layer1_outputs(7969));
    layer2_outputs(8991) <= layer1_outputs(972);
    layer2_outputs(8992) <= not((layer1_outputs(7702)) xor (layer1_outputs(7640)));
    layer2_outputs(8993) <= (layer1_outputs(4400)) and (layer1_outputs(4468));
    layer2_outputs(8994) <= layer1_outputs(6397);
    layer2_outputs(8995) <= (layer1_outputs(5670)) xor (layer1_outputs(9728));
    layer2_outputs(8996) <= not(layer1_outputs(4245));
    layer2_outputs(8997) <= (layer1_outputs(9239)) or (layer1_outputs(2459));
    layer2_outputs(8998) <= layer1_outputs(6388);
    layer2_outputs(8999) <= not(layer1_outputs(2877));
    layer2_outputs(9000) <= not(layer1_outputs(4447)) or (layer1_outputs(2816));
    layer2_outputs(9001) <= (layer1_outputs(3982)) and not (layer1_outputs(8927));
    layer2_outputs(9002) <= not(layer1_outputs(11351)) or (layer1_outputs(6235));
    layer2_outputs(9003) <= layer1_outputs(9912);
    layer2_outputs(9004) <= not((layer1_outputs(11592)) xor (layer1_outputs(10909)));
    layer2_outputs(9005) <= layer1_outputs(10169);
    layer2_outputs(9006) <= not(layer1_outputs(6674)) or (layer1_outputs(7003));
    layer2_outputs(9007) <= not((layer1_outputs(4309)) xor (layer1_outputs(9894)));
    layer2_outputs(9008) <= layer1_outputs(7148);
    layer2_outputs(9009) <= (layer1_outputs(10705)) and not (layer1_outputs(5692));
    layer2_outputs(9010) <= not(layer1_outputs(1626));
    layer2_outputs(9011) <= not(layer1_outputs(2763));
    layer2_outputs(9012) <= not((layer1_outputs(5337)) xor (layer1_outputs(10552)));
    layer2_outputs(9013) <= layer1_outputs(10022);
    layer2_outputs(9014) <= (layer1_outputs(11117)) and (layer1_outputs(859));
    layer2_outputs(9015) <= not((layer1_outputs(12000)) or (layer1_outputs(5934)));
    layer2_outputs(9016) <= not(layer1_outputs(5226));
    layer2_outputs(9017) <= (layer1_outputs(6017)) and (layer1_outputs(24));
    layer2_outputs(9018) <= (layer1_outputs(6796)) or (layer1_outputs(1112));
    layer2_outputs(9019) <= (layer1_outputs(5881)) and (layer1_outputs(9174));
    layer2_outputs(9020) <= not((layer1_outputs(9771)) and (layer1_outputs(10816)));
    layer2_outputs(9021) <= layer1_outputs(10544);
    layer2_outputs(9022) <= not(layer1_outputs(1815)) or (layer1_outputs(6336));
    layer2_outputs(9023) <= (layer1_outputs(4181)) and not (layer1_outputs(6711));
    layer2_outputs(9024) <= layer1_outputs(4590);
    layer2_outputs(9025) <= layer1_outputs(11692);
    layer2_outputs(9026) <= (layer1_outputs(9796)) or (layer1_outputs(4612));
    layer2_outputs(9027) <= not(layer1_outputs(7339));
    layer2_outputs(9028) <= not(layer1_outputs(8991));
    layer2_outputs(9029) <= (layer1_outputs(1041)) or (layer1_outputs(8270));
    layer2_outputs(9030) <= not((layer1_outputs(6961)) and (layer1_outputs(12567)));
    layer2_outputs(9031) <= layer1_outputs(9374);
    layer2_outputs(9032) <= layer1_outputs(12071);
    layer2_outputs(9033) <= layer1_outputs(9618);
    layer2_outputs(9034) <= not(layer1_outputs(1768));
    layer2_outputs(9035) <= not(layer1_outputs(5274));
    layer2_outputs(9036) <= not((layer1_outputs(4787)) and (layer1_outputs(3267)));
    layer2_outputs(9037) <= layer1_outputs(2700);
    layer2_outputs(9038) <= not((layer1_outputs(1249)) xor (layer1_outputs(3109)));
    layer2_outputs(9039) <= not((layer1_outputs(3565)) xor (layer1_outputs(10475)));
    layer2_outputs(9040) <= not(layer1_outputs(1178));
    layer2_outputs(9041) <= (layer1_outputs(6411)) xor (layer1_outputs(9671));
    layer2_outputs(9042) <= (layer1_outputs(4555)) and not (layer1_outputs(3881));
    layer2_outputs(9043) <= layer1_outputs(10224);
    layer2_outputs(9044) <= (layer1_outputs(4679)) and not (layer1_outputs(12637));
    layer2_outputs(9045) <= layer1_outputs(935);
    layer2_outputs(9046) <= not(layer1_outputs(4816));
    layer2_outputs(9047) <= (layer1_outputs(3881)) or (layer1_outputs(11081));
    layer2_outputs(9048) <= (layer1_outputs(4092)) or (layer1_outputs(4403));
    layer2_outputs(9049) <= layer1_outputs(7596);
    layer2_outputs(9050) <= not(layer1_outputs(3083));
    layer2_outputs(9051) <= (layer1_outputs(5400)) and (layer1_outputs(9876));
    layer2_outputs(9052) <= layer1_outputs(12489);
    layer2_outputs(9053) <= not(layer1_outputs(10737));
    layer2_outputs(9054) <= not(layer1_outputs(904));
    layer2_outputs(9055) <= not(layer1_outputs(12626));
    layer2_outputs(9056) <= not((layer1_outputs(3258)) or (layer1_outputs(6817)));
    layer2_outputs(9057) <= not(layer1_outputs(2813));
    layer2_outputs(9058) <= layer1_outputs(1945);
    layer2_outputs(9059) <= layer1_outputs(6765);
    layer2_outputs(9060) <= not(layer1_outputs(4837));
    layer2_outputs(9061) <= (layer1_outputs(10711)) and not (layer1_outputs(9708));
    layer2_outputs(9062) <= not((layer1_outputs(4123)) and (layer1_outputs(6898)));
    layer2_outputs(9063) <= not(layer1_outputs(7042));
    layer2_outputs(9064) <= not(layer1_outputs(1587));
    layer2_outputs(9065) <= (layer1_outputs(3539)) and (layer1_outputs(10051));
    layer2_outputs(9066) <= not(layer1_outputs(5222));
    layer2_outputs(9067) <= (layer1_outputs(11778)) xor (layer1_outputs(2105));
    layer2_outputs(9068) <= not((layer1_outputs(2107)) and (layer1_outputs(2103)));
    layer2_outputs(9069) <= not(layer1_outputs(8475)) or (layer1_outputs(3059));
    layer2_outputs(9070) <= not((layer1_outputs(1250)) and (layer1_outputs(6745)));
    layer2_outputs(9071) <= not(layer1_outputs(10874)) or (layer1_outputs(9002));
    layer2_outputs(9072) <= (layer1_outputs(9546)) and not (layer1_outputs(1956));
    layer2_outputs(9073) <= layer1_outputs(11209);
    layer2_outputs(9074) <= (layer1_outputs(3389)) xor (layer1_outputs(8670));
    layer2_outputs(9075) <= not(layer1_outputs(8922));
    layer2_outputs(9076) <= (layer1_outputs(7139)) xor (layer1_outputs(2043));
    layer2_outputs(9077) <= (layer1_outputs(8599)) xor (layer1_outputs(6408));
    layer2_outputs(9078) <= (layer1_outputs(12642)) and not (layer1_outputs(5269));
    layer2_outputs(9079) <= not(layer1_outputs(3403));
    layer2_outputs(9080) <= layer1_outputs(51);
    layer2_outputs(9081) <= (layer1_outputs(5224)) and not (layer1_outputs(6136));
    layer2_outputs(9082) <= not(layer1_outputs(6988));
    layer2_outputs(9083) <= not(layer1_outputs(6188));
    layer2_outputs(9084) <= not((layer1_outputs(1088)) or (layer1_outputs(4370)));
    layer2_outputs(9085) <= not((layer1_outputs(9133)) and (layer1_outputs(1350)));
    layer2_outputs(9086) <= (layer1_outputs(2026)) or (layer1_outputs(7268));
    layer2_outputs(9087) <= not(layer1_outputs(3378)) or (layer1_outputs(4805));
    layer2_outputs(9088) <= not((layer1_outputs(8342)) xor (layer1_outputs(8077)));
    layer2_outputs(9089) <= (layer1_outputs(1267)) and (layer1_outputs(5781));
    layer2_outputs(9090) <= (layer1_outputs(3912)) and (layer1_outputs(12502));
    layer2_outputs(9091) <= layer1_outputs(10026);
    layer2_outputs(9092) <= layer1_outputs(4284);
    layer2_outputs(9093) <= layer1_outputs(7806);
    layer2_outputs(9094) <= (layer1_outputs(5014)) and not (layer1_outputs(5238));
    layer2_outputs(9095) <= (layer1_outputs(10183)) xor (layer1_outputs(5716));
    layer2_outputs(9096) <= not(layer1_outputs(11178));
    layer2_outputs(9097) <= layer1_outputs(2200);
    layer2_outputs(9098) <= (layer1_outputs(623)) and not (layer1_outputs(7997));
    layer2_outputs(9099) <= (layer1_outputs(1110)) and not (layer1_outputs(6054));
    layer2_outputs(9100) <= (layer1_outputs(7252)) or (layer1_outputs(12429));
    layer2_outputs(9101) <= not(layer1_outputs(445));
    layer2_outputs(9102) <= layer1_outputs(10007);
    layer2_outputs(9103) <= layer1_outputs(11005);
    layer2_outputs(9104) <= not(layer1_outputs(1997));
    layer2_outputs(9105) <= layer1_outputs(1235);
    layer2_outputs(9106) <= not(layer1_outputs(12551));
    layer2_outputs(9107) <= (layer1_outputs(2160)) and not (layer1_outputs(8664));
    layer2_outputs(9108) <= not(layer1_outputs(8341));
    layer2_outputs(9109) <= (layer1_outputs(7283)) and not (layer1_outputs(9702));
    layer2_outputs(9110) <= layer1_outputs(6299);
    layer2_outputs(9111) <= layer1_outputs(1005);
    layer2_outputs(9112) <= layer1_outputs(6927);
    layer2_outputs(9113) <= (layer1_outputs(8570)) and not (layer1_outputs(11004));
    layer2_outputs(9114) <= not(layer1_outputs(3268));
    layer2_outputs(9115) <= not((layer1_outputs(11125)) and (layer1_outputs(4205)));
    layer2_outputs(9116) <= (layer1_outputs(845)) and not (layer1_outputs(12629));
    layer2_outputs(9117) <= layer1_outputs(7087);
    layer2_outputs(9118) <= not((layer1_outputs(12331)) or (layer1_outputs(6755)));
    layer2_outputs(9119) <= not(layer1_outputs(2713));
    layer2_outputs(9120) <= not(layer1_outputs(5262)) or (layer1_outputs(4892));
    layer2_outputs(9121) <= not(layer1_outputs(4258)) or (layer1_outputs(4808));
    layer2_outputs(9122) <= layer1_outputs(3941);
    layer2_outputs(9123) <= layer1_outputs(6052);
    layer2_outputs(9124) <= not(layer1_outputs(8138));
    layer2_outputs(9125) <= not(layer1_outputs(4890));
    layer2_outputs(9126) <= not((layer1_outputs(6928)) and (layer1_outputs(10027)));
    layer2_outputs(9127) <= (layer1_outputs(9521)) xor (layer1_outputs(7264));
    layer2_outputs(9128) <= not((layer1_outputs(7511)) xor (layer1_outputs(2119)));
    layer2_outputs(9129) <= layer1_outputs(4324);
    layer2_outputs(9130) <= not(layer1_outputs(6078));
    layer2_outputs(9131) <= layer1_outputs(9167);
    layer2_outputs(9132) <= not(layer1_outputs(326));
    layer2_outputs(9133) <= layer1_outputs(11947);
    layer2_outputs(9134) <= (layer1_outputs(8530)) xor (layer1_outputs(9396));
    layer2_outputs(9135) <= (layer1_outputs(4616)) and (layer1_outputs(3265));
    layer2_outputs(9136) <= (layer1_outputs(10651)) or (layer1_outputs(11612));
    layer2_outputs(9137) <= not(layer1_outputs(11286)) or (layer1_outputs(10025));
    layer2_outputs(9138) <= not(layer1_outputs(12011)) or (layer1_outputs(2720));
    layer2_outputs(9139) <= not(layer1_outputs(4027));
    layer2_outputs(9140) <= (layer1_outputs(2860)) xor (layer1_outputs(9811));
    layer2_outputs(9141) <= not((layer1_outputs(2326)) and (layer1_outputs(8802)));
    layer2_outputs(9142) <= (layer1_outputs(11463)) and not (layer1_outputs(6052));
    layer2_outputs(9143) <= (layer1_outputs(12331)) and not (layer1_outputs(6275));
    layer2_outputs(9144) <= not(layer1_outputs(11038));
    layer2_outputs(9145) <= layer1_outputs(5403);
    layer2_outputs(9146) <= not(layer1_outputs(10174));
    layer2_outputs(9147) <= (layer1_outputs(12689)) and (layer1_outputs(749));
    layer2_outputs(9148) <= not((layer1_outputs(3691)) xor (layer1_outputs(3014)));
    layer2_outputs(9149) <= layer1_outputs(1435);
    layer2_outputs(9150) <= layer1_outputs(6432);
    layer2_outputs(9151) <= layer1_outputs(1253);
    layer2_outputs(9152) <= not((layer1_outputs(1624)) xor (layer1_outputs(9269)));
    layer2_outputs(9153) <= layer1_outputs(6103);
    layer2_outputs(9154) <= not((layer1_outputs(1354)) xor (layer1_outputs(714)));
    layer2_outputs(9155) <= not(layer1_outputs(4287)) or (layer1_outputs(9701));
    layer2_outputs(9156) <= not((layer1_outputs(2597)) xor (layer1_outputs(1968)));
    layer2_outputs(9157) <= layer1_outputs(1004);
    layer2_outputs(9158) <= (layer1_outputs(2110)) and not (layer1_outputs(3046));
    layer2_outputs(9159) <= (layer1_outputs(8695)) and not (layer1_outputs(12365));
    layer2_outputs(9160) <= layer1_outputs(10119);
    layer2_outputs(9161) <= (layer1_outputs(11048)) and (layer1_outputs(9824));
    layer2_outputs(9162) <= (layer1_outputs(3161)) and not (layer1_outputs(109));
    layer2_outputs(9163) <= layer1_outputs(3741);
    layer2_outputs(9164) <= not(layer1_outputs(1145));
    layer2_outputs(9165) <= not(layer1_outputs(6347));
    layer2_outputs(9166) <= not(layer1_outputs(9257));
    layer2_outputs(9167) <= layer1_outputs(544);
    layer2_outputs(9168) <= (layer1_outputs(9981)) xor (layer1_outputs(7774));
    layer2_outputs(9169) <= (layer1_outputs(597)) and not (layer1_outputs(2370));
    layer2_outputs(9170) <= not(layer1_outputs(8760));
    layer2_outputs(9171) <= layer1_outputs(1327);
    layer2_outputs(9172) <= not((layer1_outputs(7028)) xor (layer1_outputs(9660)));
    layer2_outputs(9173) <= (layer1_outputs(80)) and not (layer1_outputs(5034));
    layer2_outputs(9174) <= layer1_outputs(9077);
    layer2_outputs(9175) <= not(layer1_outputs(2975));
    layer2_outputs(9176) <= layer1_outputs(6083);
    layer2_outputs(9177) <= layer1_outputs(8467);
    layer2_outputs(9178) <= (layer1_outputs(5718)) xor (layer1_outputs(10171));
    layer2_outputs(9179) <= not(layer1_outputs(1363));
    layer2_outputs(9180) <= not(layer1_outputs(7706));
    layer2_outputs(9181) <= (layer1_outputs(2081)) and (layer1_outputs(5097));
    layer2_outputs(9182) <= not((layer1_outputs(9178)) xor (layer1_outputs(7973)));
    layer2_outputs(9183) <= (layer1_outputs(9880)) or (layer1_outputs(4466));
    layer2_outputs(9184) <= not(layer1_outputs(7335));
    layer2_outputs(9185) <= not(layer1_outputs(6768));
    layer2_outputs(9186) <= layer1_outputs(4673);
    layer2_outputs(9187) <= not((layer1_outputs(7197)) and (layer1_outputs(3846)));
    layer2_outputs(9188) <= (layer1_outputs(10695)) and not (layer1_outputs(3351));
    layer2_outputs(9189) <= layer1_outputs(9069);
    layer2_outputs(9190) <= not(layer1_outputs(7055));
    layer2_outputs(9191) <= layer1_outputs(3472);
    layer2_outputs(9192) <= not((layer1_outputs(2097)) xor (layer1_outputs(3357)));
    layer2_outputs(9193) <= layer1_outputs(12701);
    layer2_outputs(9194) <= (layer1_outputs(3730)) and (layer1_outputs(3415));
    layer2_outputs(9195) <= not((layer1_outputs(11530)) xor (layer1_outputs(12534)));
    layer2_outputs(9196) <= '1';
    layer2_outputs(9197) <= layer1_outputs(5705);
    layer2_outputs(9198) <= not(layer1_outputs(3309));
    layer2_outputs(9199) <= (layer1_outputs(12747)) or (layer1_outputs(9944));
    layer2_outputs(9200) <= not(layer1_outputs(6194));
    layer2_outputs(9201) <= layer1_outputs(4807);
    layer2_outputs(9202) <= not(layer1_outputs(1824));
    layer2_outputs(9203) <= not(layer1_outputs(2312));
    layer2_outputs(9204) <= not(layer1_outputs(10295));
    layer2_outputs(9205) <= not(layer1_outputs(1378));
    layer2_outputs(9206) <= not(layer1_outputs(6521));
    layer2_outputs(9207) <= not((layer1_outputs(12048)) and (layer1_outputs(11583)));
    layer2_outputs(9208) <= not(layer1_outputs(9503)) or (layer1_outputs(6827));
    layer2_outputs(9209) <= (layer1_outputs(4969)) and (layer1_outputs(3151));
    layer2_outputs(9210) <= not(layer1_outputs(12209));
    layer2_outputs(9211) <= not((layer1_outputs(4034)) and (layer1_outputs(2730)));
    layer2_outputs(9212) <= layer1_outputs(543);
    layer2_outputs(9213) <= not((layer1_outputs(4109)) or (layer1_outputs(538)));
    layer2_outputs(9214) <= layer1_outputs(11676);
    layer2_outputs(9215) <= not(layer1_outputs(3511)) or (layer1_outputs(8004));
    layer2_outputs(9216) <= not(layer1_outputs(5676)) or (layer1_outputs(2838));
    layer2_outputs(9217) <= not(layer1_outputs(2688));
    layer2_outputs(9218) <= not(layer1_outputs(7049)) or (layer1_outputs(3908));
    layer2_outputs(9219) <= layer1_outputs(5248);
    layer2_outputs(9220) <= not((layer1_outputs(10572)) or (layer1_outputs(6223)));
    layer2_outputs(9221) <= (layer1_outputs(12087)) and (layer1_outputs(10109));
    layer2_outputs(9222) <= layer1_outputs(6917);
    layer2_outputs(9223) <= not(layer1_outputs(8804)) or (layer1_outputs(9438));
    layer2_outputs(9224) <= not(layer1_outputs(9866)) or (layer1_outputs(8174));
    layer2_outputs(9225) <= not((layer1_outputs(8793)) xor (layer1_outputs(1976)));
    layer2_outputs(9226) <= (layer1_outputs(7245)) xor (layer1_outputs(5014));
    layer2_outputs(9227) <= (layer1_outputs(4811)) and (layer1_outputs(66));
    layer2_outputs(9228) <= not(layer1_outputs(12240));
    layer2_outputs(9229) <= (layer1_outputs(9957)) and not (layer1_outputs(2734));
    layer2_outputs(9230) <= layer1_outputs(12030);
    layer2_outputs(9231) <= not((layer1_outputs(3315)) and (layer1_outputs(2275)));
    layer2_outputs(9232) <= layer1_outputs(11095);
    layer2_outputs(9233) <= not(layer1_outputs(4700));
    layer2_outputs(9234) <= not((layer1_outputs(10644)) or (layer1_outputs(2623)));
    layer2_outputs(9235) <= not((layer1_outputs(12412)) or (layer1_outputs(2969)));
    layer2_outputs(9236) <= '0';
    layer2_outputs(9237) <= not((layer1_outputs(6614)) xor (layer1_outputs(4923)));
    layer2_outputs(9238) <= (layer1_outputs(660)) and not (layer1_outputs(6870));
    layer2_outputs(9239) <= (layer1_outputs(12638)) or (layer1_outputs(5620));
    layer2_outputs(9240) <= (layer1_outputs(554)) and (layer1_outputs(2647));
    layer2_outputs(9241) <= layer1_outputs(2518);
    layer2_outputs(9242) <= not((layer1_outputs(8715)) xor (layer1_outputs(915)));
    layer2_outputs(9243) <= not(layer1_outputs(4523));
    layer2_outputs(9244) <= not((layer1_outputs(3242)) xor (layer1_outputs(7450)));
    layer2_outputs(9245) <= (layer1_outputs(9183)) xor (layer1_outputs(7151));
    layer2_outputs(9246) <= not(layer1_outputs(5028));
    layer2_outputs(9247) <= not(layer1_outputs(2620));
    layer2_outputs(9248) <= layer1_outputs(4736);
    layer2_outputs(9249) <= layer1_outputs(4252);
    layer2_outputs(9250) <= not(layer1_outputs(11428)) or (layer1_outputs(9563));
    layer2_outputs(9251) <= not((layer1_outputs(4821)) or (layer1_outputs(6028)));
    layer2_outputs(9252) <= (layer1_outputs(7808)) or (layer1_outputs(9485));
    layer2_outputs(9253) <= not(layer1_outputs(3002));
    layer2_outputs(9254) <= not(layer1_outputs(9335));
    layer2_outputs(9255) <= not(layer1_outputs(543));
    layer2_outputs(9256) <= layer1_outputs(8993);
    layer2_outputs(9257) <= (layer1_outputs(4496)) and not (layer1_outputs(5134));
    layer2_outputs(9258) <= layer1_outputs(210);
    layer2_outputs(9259) <= not(layer1_outputs(12167));
    layer2_outputs(9260) <= not(layer1_outputs(10778));
    layer2_outputs(9261) <= layer1_outputs(7582);
    layer2_outputs(9262) <= not((layer1_outputs(8984)) and (layer1_outputs(11712)));
    layer2_outputs(9263) <= (layer1_outputs(11607)) and (layer1_outputs(12368));
    layer2_outputs(9264) <= (layer1_outputs(7555)) or (layer1_outputs(4067));
    layer2_outputs(9265) <= not(layer1_outputs(4166));
    layer2_outputs(9266) <= layer1_outputs(3451);
    layer2_outputs(9267) <= not((layer1_outputs(12001)) or (layer1_outputs(12384)));
    layer2_outputs(9268) <= not(layer1_outputs(9445));
    layer2_outputs(9269) <= not(layer1_outputs(10055));
    layer2_outputs(9270) <= not((layer1_outputs(12261)) and (layer1_outputs(5328)));
    layer2_outputs(9271) <= (layer1_outputs(11415)) xor (layer1_outputs(7691));
    layer2_outputs(9272) <= not(layer1_outputs(12769));
    layer2_outputs(9273) <= (layer1_outputs(12056)) and not (layer1_outputs(11073));
    layer2_outputs(9274) <= not((layer1_outputs(1553)) xor (layer1_outputs(6966)));
    layer2_outputs(9275) <= (layer1_outputs(7422)) and not (layer1_outputs(1941));
    layer2_outputs(9276) <= layer1_outputs(3400);
    layer2_outputs(9277) <= (layer1_outputs(7927)) and not (layer1_outputs(8518));
    layer2_outputs(9278) <= layer1_outputs(12500);
    layer2_outputs(9279) <= (layer1_outputs(9804)) and not (layer1_outputs(4736));
    layer2_outputs(9280) <= not((layer1_outputs(3914)) and (layer1_outputs(2850)));
    layer2_outputs(9281) <= (layer1_outputs(12489)) and (layer1_outputs(7529));
    layer2_outputs(9282) <= layer1_outputs(8802);
    layer2_outputs(9283) <= not((layer1_outputs(442)) and (layer1_outputs(11047)));
    layer2_outputs(9284) <= (layer1_outputs(9924)) xor (layer1_outputs(2263));
    layer2_outputs(9285) <= (layer1_outputs(7884)) or (layer1_outputs(5486));
    layer2_outputs(9286) <= layer1_outputs(6829);
    layer2_outputs(9287) <= layer1_outputs(4297);
    layer2_outputs(9288) <= not(layer1_outputs(8253)) or (layer1_outputs(370));
    layer2_outputs(9289) <= not(layer1_outputs(610));
    layer2_outputs(9290) <= not((layer1_outputs(3917)) or (layer1_outputs(12494)));
    layer2_outputs(9291) <= layer1_outputs(8609);
    layer2_outputs(9292) <= layer1_outputs(5931);
    layer2_outputs(9293) <= not(layer1_outputs(10586));
    layer2_outputs(9294) <= not(layer1_outputs(10394)) or (layer1_outputs(7508));
    layer2_outputs(9295) <= (layer1_outputs(7701)) xor (layer1_outputs(1680));
    layer2_outputs(9296) <= (layer1_outputs(5416)) and not (layer1_outputs(9728));
    layer2_outputs(9297) <= (layer1_outputs(8231)) or (layer1_outputs(1586));
    layer2_outputs(9298) <= not(layer1_outputs(2432)) or (layer1_outputs(5407));
    layer2_outputs(9299) <= layer1_outputs(1874);
    layer2_outputs(9300) <= layer1_outputs(9358);
    layer2_outputs(9301) <= not((layer1_outputs(6927)) xor (layer1_outputs(11121)));
    layer2_outputs(9302) <= (layer1_outputs(3134)) or (layer1_outputs(1090));
    layer2_outputs(9303) <= layer1_outputs(10488);
    layer2_outputs(9304) <= layer1_outputs(4439);
    layer2_outputs(9305) <= not(layer1_outputs(9688));
    layer2_outputs(9306) <= layer1_outputs(277);
    layer2_outputs(9307) <= (layer1_outputs(7325)) and not (layer1_outputs(5666));
    layer2_outputs(9308) <= '1';
    layer2_outputs(9309) <= layer1_outputs(7131);
    layer2_outputs(9310) <= not(layer1_outputs(7220));
    layer2_outputs(9311) <= not(layer1_outputs(5220));
    layer2_outputs(9312) <= (layer1_outputs(615)) xor (layer1_outputs(11119));
    layer2_outputs(9313) <= not((layer1_outputs(2334)) xor (layer1_outputs(11284)));
    layer2_outputs(9314) <= (layer1_outputs(3607)) or (layer1_outputs(1290));
    layer2_outputs(9315) <= layer1_outputs(10948);
    layer2_outputs(9316) <= (layer1_outputs(9928)) xor (layer1_outputs(3308));
    layer2_outputs(9317) <= layer1_outputs(12677);
    layer2_outputs(9318) <= not(layer1_outputs(8234)) or (layer1_outputs(2254));
    layer2_outputs(9319) <= layer1_outputs(6359);
    layer2_outputs(9320) <= not(layer1_outputs(4314));
    layer2_outputs(9321) <= not((layer1_outputs(10362)) xor (layer1_outputs(9927)));
    layer2_outputs(9322) <= layer1_outputs(3960);
    layer2_outputs(9323) <= layer1_outputs(11865);
    layer2_outputs(9324) <= (layer1_outputs(2638)) or (layer1_outputs(2138));
    layer2_outputs(9325) <= not((layer1_outputs(11903)) xor (layer1_outputs(8356)));
    layer2_outputs(9326) <= (layer1_outputs(430)) and not (layer1_outputs(2016));
    layer2_outputs(9327) <= (layer1_outputs(3889)) and not (layer1_outputs(3405));
    layer2_outputs(9328) <= layer1_outputs(2621);
    layer2_outputs(9329) <= not(layer1_outputs(12748));
    layer2_outputs(9330) <= (layer1_outputs(6265)) and not (layer1_outputs(8433));
    layer2_outputs(9331) <= not((layer1_outputs(10517)) or (layer1_outputs(3567)));
    layer2_outputs(9332) <= not(layer1_outputs(459));
    layer2_outputs(9333) <= not(layer1_outputs(12452));
    layer2_outputs(9334) <= not((layer1_outputs(10922)) and (layer1_outputs(11732)));
    layer2_outputs(9335) <= layer1_outputs(2513);
    layer2_outputs(9336) <= not(layer1_outputs(10507));
    layer2_outputs(9337) <= (layer1_outputs(2798)) and (layer1_outputs(12342));
    layer2_outputs(9338) <= not((layer1_outputs(7438)) xor (layer1_outputs(9128)));
    layer2_outputs(9339) <= not(layer1_outputs(1194));
    layer2_outputs(9340) <= not(layer1_outputs(2859));
    layer2_outputs(9341) <= layer1_outputs(10454);
    layer2_outputs(9342) <= layer1_outputs(1968);
    layer2_outputs(9343) <= (layer1_outputs(3235)) and not (layer1_outputs(9120));
    layer2_outputs(9344) <= (layer1_outputs(4645)) and (layer1_outputs(4595));
    layer2_outputs(9345) <= not(layer1_outputs(8468)) or (layer1_outputs(4280));
    layer2_outputs(9346) <= not((layer1_outputs(6364)) and (layer1_outputs(8055)));
    layer2_outputs(9347) <= layer1_outputs(9960);
    layer2_outputs(9348) <= not(layer1_outputs(3936));
    layer2_outputs(9349) <= not(layer1_outputs(10747));
    layer2_outputs(9350) <= not(layer1_outputs(1625));
    layer2_outputs(9351) <= layer1_outputs(6544);
    layer2_outputs(9352) <= layer1_outputs(3883);
    layer2_outputs(9353) <= (layer1_outputs(789)) and (layer1_outputs(4231));
    layer2_outputs(9354) <= not((layer1_outputs(5459)) and (layer1_outputs(1245)));
    layer2_outputs(9355) <= not(layer1_outputs(2609));
    layer2_outputs(9356) <= (layer1_outputs(7069)) and not (layer1_outputs(3217));
    layer2_outputs(9357) <= not((layer1_outputs(10557)) xor (layer1_outputs(3933)));
    layer2_outputs(9358) <= layer1_outputs(5993);
    layer2_outputs(9359) <= not(layer1_outputs(10958));
    layer2_outputs(9360) <= layer1_outputs(7451);
    layer2_outputs(9361) <= not(layer1_outputs(11821));
    layer2_outputs(9362) <= (layer1_outputs(10353)) and not (layer1_outputs(6813));
    layer2_outputs(9363) <= not(layer1_outputs(7775));
    layer2_outputs(9364) <= '1';
    layer2_outputs(9365) <= not((layer1_outputs(12593)) and (layer1_outputs(6968)));
    layer2_outputs(9366) <= layer1_outputs(10626);
    layer2_outputs(9367) <= not(layer1_outputs(1212));
    layer2_outputs(9368) <= not((layer1_outputs(1508)) xor (layer1_outputs(2029)));
    layer2_outputs(9369) <= layer1_outputs(11528);
    layer2_outputs(9370) <= (layer1_outputs(8363)) or (layer1_outputs(7676));
    layer2_outputs(9371) <= not(layer1_outputs(2418)) or (layer1_outputs(2127));
    layer2_outputs(9372) <= layer1_outputs(225);
    layer2_outputs(9373) <= not(layer1_outputs(10037));
    layer2_outputs(9374) <= not((layer1_outputs(359)) xor (layer1_outputs(5235)));
    layer2_outputs(9375) <= (layer1_outputs(279)) xor (layer1_outputs(11035));
    layer2_outputs(9376) <= (layer1_outputs(8588)) or (layer1_outputs(19));
    layer2_outputs(9377) <= not(layer1_outputs(11572));
    layer2_outputs(9378) <= not(layer1_outputs(8650));
    layer2_outputs(9379) <= layer1_outputs(6045);
    layer2_outputs(9380) <= not((layer1_outputs(1087)) xor (layer1_outputs(3933)));
    layer2_outputs(9381) <= (layer1_outputs(12657)) and (layer1_outputs(9447));
    layer2_outputs(9382) <= not((layer1_outputs(4422)) xor (layer1_outputs(11418)));
    layer2_outputs(9383) <= layer1_outputs(4780);
    layer2_outputs(9384) <= '1';
    layer2_outputs(9385) <= not(layer1_outputs(12653));
    layer2_outputs(9386) <= not((layer1_outputs(6104)) and (layer1_outputs(3326)));
    layer2_outputs(9387) <= not((layer1_outputs(11216)) xor (layer1_outputs(12315)));
    layer2_outputs(9388) <= '0';
    layer2_outputs(9389) <= (layer1_outputs(7741)) and not (layer1_outputs(8963));
    layer2_outputs(9390) <= layer1_outputs(9863);
    layer2_outputs(9391) <= layer1_outputs(8209);
    layer2_outputs(9392) <= layer1_outputs(12517);
    layer2_outputs(9393) <= not(layer1_outputs(1785));
    layer2_outputs(9394) <= layer1_outputs(5482);
    layer2_outputs(9395) <= layer1_outputs(9535);
    layer2_outputs(9396) <= layer1_outputs(9742);
    layer2_outputs(9397) <= not(layer1_outputs(3469));
    layer2_outputs(9398) <= (layer1_outputs(5876)) xor (layer1_outputs(7140));
    layer2_outputs(9399) <= (layer1_outputs(11029)) and not (layer1_outputs(12711));
    layer2_outputs(9400) <= layer1_outputs(4782);
    layer2_outputs(9401) <= (layer1_outputs(10895)) xor (layer1_outputs(4667));
    layer2_outputs(9402) <= not((layer1_outputs(4952)) xor (layer1_outputs(3864)));
    layer2_outputs(9403) <= (layer1_outputs(6804)) and not (layer1_outputs(3720));
    layer2_outputs(9404) <= (layer1_outputs(220)) xor (layer1_outputs(2778));
    layer2_outputs(9405) <= not(layer1_outputs(778));
    layer2_outputs(9406) <= layer1_outputs(12792);
    layer2_outputs(9407) <= not((layer1_outputs(9115)) or (layer1_outputs(11239)));
    layer2_outputs(9408) <= (layer1_outputs(516)) or (layer1_outputs(12020));
    layer2_outputs(9409) <= not((layer1_outputs(12447)) xor (layer1_outputs(5663)));
    layer2_outputs(9410) <= not(layer1_outputs(4857));
    layer2_outputs(9411) <= (layer1_outputs(10659)) and not (layer1_outputs(5873));
    layer2_outputs(9412) <= (layer1_outputs(6086)) and not (layer1_outputs(669));
    layer2_outputs(9413) <= layer1_outputs(7718);
    layer2_outputs(9414) <= (layer1_outputs(11302)) and not (layer1_outputs(5832));
    layer2_outputs(9415) <= layer1_outputs(2199);
    layer2_outputs(9416) <= not((layer1_outputs(5038)) xor (layer1_outputs(2618)));
    layer2_outputs(9417) <= layer1_outputs(3464);
    layer2_outputs(9418) <= not(layer1_outputs(10371));
    layer2_outputs(9419) <= (layer1_outputs(8814)) and not (layer1_outputs(4651));
    layer2_outputs(9420) <= (layer1_outputs(11146)) and not (layer1_outputs(461));
    layer2_outputs(9421) <= not((layer1_outputs(2151)) xor (layer1_outputs(8909)));
    layer2_outputs(9422) <= (layer1_outputs(17)) and not (layer1_outputs(11150));
    layer2_outputs(9423) <= (layer1_outputs(12791)) xor (layer1_outputs(2961));
    layer2_outputs(9424) <= not((layer1_outputs(1618)) and (layer1_outputs(7149)));
    layer2_outputs(9425) <= (layer1_outputs(10075)) xor (layer1_outputs(3087));
    layer2_outputs(9426) <= not(layer1_outputs(6170)) or (layer1_outputs(10429));
    layer2_outputs(9427) <= not(layer1_outputs(11742));
    layer2_outputs(9428) <= not((layer1_outputs(5377)) and (layer1_outputs(8702)));
    layer2_outputs(9429) <= (layer1_outputs(2297)) and not (layer1_outputs(8727));
    layer2_outputs(9430) <= (layer1_outputs(1556)) and not (layer1_outputs(770));
    layer2_outputs(9431) <= not((layer1_outputs(7484)) xor (layer1_outputs(8583)));
    layer2_outputs(9432) <= layer1_outputs(6262);
    layer2_outputs(9433) <= (layer1_outputs(8278)) xor (layer1_outputs(1417));
    layer2_outputs(9434) <= not(layer1_outputs(10559));
    layer2_outputs(9435) <= not(layer1_outputs(11610));
    layer2_outputs(9436) <= (layer1_outputs(5754)) and (layer1_outputs(11621));
    layer2_outputs(9437) <= '0';
    layer2_outputs(9438) <= (layer1_outputs(11218)) and not (layer1_outputs(1323));
    layer2_outputs(9439) <= not(layer1_outputs(12613));
    layer2_outputs(9440) <= '1';
    layer2_outputs(9441) <= not(layer1_outputs(9542));
    layer2_outputs(9442) <= (layer1_outputs(6210)) and (layer1_outputs(2442));
    layer2_outputs(9443) <= layer1_outputs(7992);
    layer2_outputs(9444) <= (layer1_outputs(10969)) xor (layer1_outputs(3484));
    layer2_outputs(9445) <= layer1_outputs(5375);
    layer2_outputs(9446) <= (layer1_outputs(6466)) and (layer1_outputs(7838));
    layer2_outputs(9447) <= (layer1_outputs(1121)) xor (layer1_outputs(11096));
    layer2_outputs(9448) <= not(layer1_outputs(10039));
    layer2_outputs(9449) <= (layer1_outputs(1057)) or (layer1_outputs(9992));
    layer2_outputs(9450) <= layer1_outputs(8059);
    layer2_outputs(9451) <= not(layer1_outputs(12546));
    layer2_outputs(9452) <= layer1_outputs(3819);
    layer2_outputs(9453) <= not((layer1_outputs(9810)) or (layer1_outputs(9835)));
    layer2_outputs(9454) <= not(layer1_outputs(11789));
    layer2_outputs(9455) <= (layer1_outputs(10798)) xor (layer1_outputs(10068));
    layer2_outputs(9456) <= not(layer1_outputs(4756));
    layer2_outputs(9457) <= not((layer1_outputs(11318)) and (layer1_outputs(7943)));
    layer2_outputs(9458) <= not(layer1_outputs(10956)) or (layer1_outputs(4940));
    layer2_outputs(9459) <= layer1_outputs(10415);
    layer2_outputs(9460) <= layer1_outputs(7137);
    layer2_outputs(9461) <= not((layer1_outputs(2635)) and (layer1_outputs(11787)));
    layer2_outputs(9462) <= not((layer1_outputs(335)) xor (layer1_outputs(11076)));
    layer2_outputs(9463) <= (layer1_outputs(6648)) and not (layer1_outputs(6083));
    layer2_outputs(9464) <= (layer1_outputs(1751)) and (layer1_outputs(2643));
    layer2_outputs(9465) <= (layer1_outputs(10863)) xor (layer1_outputs(8175));
    layer2_outputs(9466) <= not(layer1_outputs(3471));
    layer2_outputs(9467) <= (layer1_outputs(236)) xor (layer1_outputs(4630));
    layer2_outputs(9468) <= (layer1_outputs(617)) xor (layer1_outputs(7423));
    layer2_outputs(9469) <= layer1_outputs(5157);
    layer2_outputs(9470) <= not((layer1_outputs(7593)) and (layer1_outputs(6477)));
    layer2_outputs(9471) <= layer1_outputs(6251);
    layer2_outputs(9472) <= layer1_outputs(3296);
    layer2_outputs(9473) <= not(layer1_outputs(7006));
    layer2_outputs(9474) <= (layer1_outputs(737)) xor (layer1_outputs(6026));
    layer2_outputs(9475) <= not(layer1_outputs(10104));
    layer2_outputs(9476) <= not(layer1_outputs(2187));
    layer2_outputs(9477) <= (layer1_outputs(9367)) and (layer1_outputs(11871));
    layer2_outputs(9478) <= (layer1_outputs(8679)) or (layer1_outputs(6436));
    layer2_outputs(9479) <= not((layer1_outputs(4489)) and (layer1_outputs(9256)));
    layer2_outputs(9480) <= (layer1_outputs(6991)) xor (layer1_outputs(924));
    layer2_outputs(9481) <= not(layer1_outputs(1573));
    layer2_outputs(9482) <= layer1_outputs(4);
    layer2_outputs(9483) <= not(layer1_outputs(10072));
    layer2_outputs(9484) <= not(layer1_outputs(2277));
    layer2_outputs(9485) <= not(layer1_outputs(2105)) or (layer1_outputs(9803));
    layer2_outputs(9486) <= layer1_outputs(6165);
    layer2_outputs(9487) <= not(layer1_outputs(2052));
    layer2_outputs(9488) <= layer1_outputs(2444);
    layer2_outputs(9489) <= not(layer1_outputs(6894));
    layer2_outputs(9490) <= not(layer1_outputs(11124)) or (layer1_outputs(2643));
    layer2_outputs(9491) <= (layer1_outputs(6245)) xor (layer1_outputs(2752));
    layer2_outputs(9492) <= layer1_outputs(5693);
    layer2_outputs(9493) <= (layer1_outputs(2207)) or (layer1_outputs(2529));
    layer2_outputs(9494) <= not((layer1_outputs(6641)) and (layer1_outputs(10377)));
    layer2_outputs(9495) <= (layer1_outputs(8197)) xor (layer1_outputs(892));
    layer2_outputs(9496) <= layer1_outputs(6282);
    layer2_outputs(9497) <= (layer1_outputs(9671)) and not (layer1_outputs(9287));
    layer2_outputs(9498) <= not(layer1_outputs(885)) or (layer1_outputs(3310));
    layer2_outputs(9499) <= layer1_outputs(7299);
    layer2_outputs(9500) <= (layer1_outputs(5089)) and (layer1_outputs(9881));
    layer2_outputs(9501) <= (layer1_outputs(8966)) and (layer1_outputs(3776));
    layer2_outputs(9502) <= layer1_outputs(2804);
    layer2_outputs(9503) <= not(layer1_outputs(4771));
    layer2_outputs(9504) <= not((layer1_outputs(8655)) or (layer1_outputs(5162)));
    layer2_outputs(9505) <= not(layer1_outputs(1140)) or (layer1_outputs(7030));
    layer2_outputs(9506) <= layer1_outputs(7834);
    layer2_outputs(9507) <= (layer1_outputs(11845)) and not (layer1_outputs(11339));
    layer2_outputs(9508) <= not((layer1_outputs(8812)) and (layer1_outputs(1272)));
    layer2_outputs(9509) <= not((layer1_outputs(9761)) or (layer1_outputs(1624)));
    layer2_outputs(9510) <= layer1_outputs(10411);
    layer2_outputs(9511) <= layer1_outputs(1945);
    layer2_outputs(9512) <= not((layer1_outputs(3890)) and (layer1_outputs(12752)));
    layer2_outputs(9513) <= layer1_outputs(5445);
    layer2_outputs(9514) <= not(layer1_outputs(11637));
    layer2_outputs(9515) <= (layer1_outputs(8916)) and (layer1_outputs(6453));
    layer2_outputs(9516) <= (layer1_outputs(10352)) xor (layer1_outputs(7679));
    layer2_outputs(9517) <= not(layer1_outputs(9649)) or (layer1_outputs(9215));
    layer2_outputs(9518) <= layer1_outputs(4453);
    layer2_outputs(9519) <= not(layer1_outputs(10237));
    layer2_outputs(9520) <= layer1_outputs(1010);
    layer2_outputs(9521) <= layer1_outputs(11956);
    layer2_outputs(9522) <= layer1_outputs(5492);
    layer2_outputs(9523) <= (layer1_outputs(3817)) and (layer1_outputs(5864));
    layer2_outputs(9524) <= not((layer1_outputs(8534)) and (layer1_outputs(2979)));
    layer2_outputs(9525) <= not(layer1_outputs(9178));
    layer2_outputs(9526) <= not(layer1_outputs(3657));
    layer2_outputs(9527) <= layer1_outputs(6497);
    layer2_outputs(9528) <= not(layer1_outputs(6963)) or (layer1_outputs(3148));
    layer2_outputs(9529) <= not(layer1_outputs(1914));
    layer2_outputs(9530) <= (layer1_outputs(2211)) xor (layer1_outputs(12793));
    layer2_outputs(9531) <= not(layer1_outputs(11877));
    layer2_outputs(9532) <= not(layer1_outputs(5167)) or (layer1_outputs(4768));
    layer2_outputs(9533) <= (layer1_outputs(12388)) and not (layer1_outputs(8249));
    layer2_outputs(9534) <= not(layer1_outputs(5824));
    layer2_outputs(9535) <= not(layer1_outputs(8184));
    layer2_outputs(9536) <= layer1_outputs(12720);
    layer2_outputs(9537) <= not(layer1_outputs(4822));
    layer2_outputs(9538) <= (layer1_outputs(2176)) xor (layer1_outputs(5025));
    layer2_outputs(9539) <= layer1_outputs(12664);
    layer2_outputs(9540) <= not(layer1_outputs(5948));
    layer2_outputs(9541) <= not(layer1_outputs(8911)) or (layer1_outputs(4441));
    layer2_outputs(9542) <= not((layer1_outputs(7341)) or (layer1_outputs(9190)));
    layer2_outputs(9543) <= layer1_outputs(12087);
    layer2_outputs(9544) <= (layer1_outputs(11981)) or (layer1_outputs(12348));
    layer2_outputs(9545) <= not((layer1_outputs(5103)) or (layer1_outputs(10843)));
    layer2_outputs(9546) <= (layer1_outputs(7211)) xor (layer1_outputs(12366));
    layer2_outputs(9547) <= layer1_outputs(2413);
    layer2_outputs(9548) <= (layer1_outputs(2226)) xor (layer1_outputs(4592));
    layer2_outputs(9549) <= not(layer1_outputs(3777));
    layer2_outputs(9550) <= (layer1_outputs(10067)) and not (layer1_outputs(10005));
    layer2_outputs(9551) <= (layer1_outputs(7486)) xor (layer1_outputs(2964));
    layer2_outputs(9552) <= layer1_outputs(7982);
    layer2_outputs(9553) <= layer1_outputs(9243);
    layer2_outputs(9554) <= not(layer1_outputs(9991));
    layer2_outputs(9555) <= layer1_outputs(3761);
    layer2_outputs(9556) <= (layer1_outputs(6237)) and not (layer1_outputs(11872));
    layer2_outputs(9557) <= (layer1_outputs(11476)) xor (layer1_outputs(8449));
    layer2_outputs(9558) <= not(layer1_outputs(2785));
    layer2_outputs(9559) <= layer1_outputs(3033);
    layer2_outputs(9560) <= not(layer1_outputs(5147));
    layer2_outputs(9561) <= layer1_outputs(11218);
    layer2_outputs(9562) <= not((layer1_outputs(6219)) and (layer1_outputs(12648)));
    layer2_outputs(9563) <= (layer1_outputs(11523)) xor (layer1_outputs(12623));
    layer2_outputs(9564) <= not(layer1_outputs(12279));
    layer2_outputs(9565) <= not(layer1_outputs(2475));
    layer2_outputs(9566) <= (layer1_outputs(12213)) and not (layer1_outputs(8983));
    layer2_outputs(9567) <= not((layer1_outputs(11718)) or (layer1_outputs(6513)));
    layer2_outputs(9568) <= layer1_outputs(4506);
    layer2_outputs(9569) <= layer1_outputs(3695);
    layer2_outputs(9570) <= not(layer1_outputs(2610)) or (layer1_outputs(5188));
    layer2_outputs(9571) <= not(layer1_outputs(7604)) or (layer1_outputs(2773));
    layer2_outputs(9572) <= not(layer1_outputs(10219));
    layer2_outputs(9573) <= not(layer1_outputs(1938)) or (layer1_outputs(4127));
    layer2_outputs(9574) <= not(layer1_outputs(6620));
    layer2_outputs(9575) <= not(layer1_outputs(3653));
    layer2_outputs(9576) <= not(layer1_outputs(457));
    layer2_outputs(9577) <= layer1_outputs(11282);
    layer2_outputs(9578) <= (layer1_outputs(12780)) and not (layer1_outputs(4333));
    layer2_outputs(9579) <= not(layer1_outputs(9013));
    layer2_outputs(9580) <= not((layer1_outputs(3823)) and (layer1_outputs(629)));
    layer2_outputs(9581) <= (layer1_outputs(11939)) xor (layer1_outputs(8508));
    layer2_outputs(9582) <= (layer1_outputs(10945)) and not (layer1_outputs(10201));
    layer2_outputs(9583) <= not((layer1_outputs(10779)) and (layer1_outputs(8291)));
    layer2_outputs(9584) <= (layer1_outputs(330)) and not (layer1_outputs(11347));
    layer2_outputs(9585) <= '1';
    layer2_outputs(9586) <= layer1_outputs(2428);
    layer2_outputs(9587) <= not(layer1_outputs(4462));
    layer2_outputs(9588) <= layer1_outputs(9705);
    layer2_outputs(9589) <= not(layer1_outputs(4114));
    layer2_outputs(9590) <= not(layer1_outputs(11708));
    layer2_outputs(9591) <= not(layer1_outputs(6914));
    layer2_outputs(9592) <= (layer1_outputs(1020)) and not (layer1_outputs(4611));
    layer2_outputs(9593) <= layer1_outputs(2796);
    layer2_outputs(9594) <= not(layer1_outputs(5338)) or (layer1_outputs(6787));
    layer2_outputs(9595) <= (layer1_outputs(7664)) and (layer1_outputs(10162));
    layer2_outputs(9596) <= layer1_outputs(7895);
    layer2_outputs(9597) <= layer1_outputs(7887);
    layer2_outputs(9598) <= not(layer1_outputs(2424));
    layer2_outputs(9599) <= '1';
    layer2_outputs(9600) <= not((layer1_outputs(6613)) xor (layer1_outputs(9642)));
    layer2_outputs(9601) <= not(layer1_outputs(3632));
    layer2_outputs(9602) <= not(layer1_outputs(4711));
    layer2_outputs(9603) <= (layer1_outputs(3872)) or (layer1_outputs(5660));
    layer2_outputs(9604) <= not(layer1_outputs(11439));
    layer2_outputs(9605) <= not(layer1_outputs(10708));
    layer2_outputs(9606) <= (layer1_outputs(1791)) xor (layer1_outputs(10941));
    layer2_outputs(9607) <= (layer1_outputs(4338)) xor (layer1_outputs(7450));
    layer2_outputs(9608) <= not((layer1_outputs(6592)) xor (layer1_outputs(7849)));
    layer2_outputs(9609) <= not(layer1_outputs(5144)) or (layer1_outputs(12422));
    layer2_outputs(9610) <= layer1_outputs(6141);
    layer2_outputs(9611) <= not(layer1_outputs(125)) or (layer1_outputs(2358));
    layer2_outputs(9612) <= not((layer1_outputs(5462)) xor (layer1_outputs(11793)));
    layer2_outputs(9613) <= not((layer1_outputs(526)) xor (layer1_outputs(11506)));
    layer2_outputs(9614) <= not((layer1_outputs(9467)) and (layer1_outputs(9747)));
    layer2_outputs(9615) <= layer1_outputs(2415);
    layer2_outputs(9616) <= not(layer1_outputs(703));
    layer2_outputs(9617) <= layer1_outputs(7311);
    layer2_outputs(9618) <= layer1_outputs(10049);
    layer2_outputs(9619) <= not((layer1_outputs(11127)) or (layer1_outputs(620)));
    layer2_outputs(9620) <= layer1_outputs(9537);
    layer2_outputs(9621) <= (layer1_outputs(170)) and not (layer1_outputs(6581));
    layer2_outputs(9622) <= not(layer1_outputs(7001));
    layer2_outputs(9623) <= (layer1_outputs(10447)) and not (layer1_outputs(3163));
    layer2_outputs(9624) <= (layer1_outputs(3551)) and (layer1_outputs(6233));
    layer2_outputs(9625) <= (layer1_outputs(11171)) xor (layer1_outputs(11164));
    layer2_outputs(9626) <= layer1_outputs(10116);
    layer2_outputs(9627) <= not((layer1_outputs(3641)) xor (layer1_outputs(10989)));
    layer2_outputs(9628) <= (layer1_outputs(7618)) xor (layer1_outputs(2524));
    layer2_outputs(9629) <= (layer1_outputs(10335)) and not (layer1_outputs(12654));
    layer2_outputs(9630) <= (layer1_outputs(9244)) or (layer1_outputs(11602));
    layer2_outputs(9631) <= layer1_outputs(10591);
    layer2_outputs(9632) <= (layer1_outputs(3084)) or (layer1_outputs(4581));
    layer2_outputs(9633) <= not((layer1_outputs(5253)) xor (layer1_outputs(79)));
    layer2_outputs(9634) <= not(layer1_outputs(6420));
    layer2_outputs(9635) <= (layer1_outputs(11503)) and not (layer1_outputs(5834));
    layer2_outputs(9636) <= not(layer1_outputs(12228));
    layer2_outputs(9637) <= (layer1_outputs(95)) xor (layer1_outputs(758));
    layer2_outputs(9638) <= layer1_outputs(3272);
    layer2_outputs(9639) <= not((layer1_outputs(6377)) or (layer1_outputs(10508)));
    layer2_outputs(9640) <= not(layer1_outputs(10175));
    layer2_outputs(9641) <= (layer1_outputs(5557)) and not (layer1_outputs(12378));
    layer2_outputs(9642) <= (layer1_outputs(6456)) and not (layer1_outputs(9323));
    layer2_outputs(9643) <= (layer1_outputs(9662)) and not (layer1_outputs(472));
    layer2_outputs(9644) <= (layer1_outputs(7763)) xor (layer1_outputs(6199));
    layer2_outputs(9645) <= not((layer1_outputs(7698)) xor (layer1_outputs(391)));
    layer2_outputs(9646) <= not(layer1_outputs(2443));
    layer2_outputs(9647) <= (layer1_outputs(3250)) xor (layer1_outputs(7634));
    layer2_outputs(9648) <= layer1_outputs(4118);
    layer2_outputs(9649) <= not(layer1_outputs(6344));
    layer2_outputs(9650) <= not((layer1_outputs(1013)) and (layer1_outputs(5532)));
    layer2_outputs(9651) <= not(layer1_outputs(5912));
    layer2_outputs(9652) <= not(layer1_outputs(4435));
    layer2_outputs(9653) <= not((layer1_outputs(5755)) xor (layer1_outputs(3861)));
    layer2_outputs(9654) <= not(layer1_outputs(12067)) or (layer1_outputs(4170));
    layer2_outputs(9655) <= not((layer1_outputs(11310)) xor (layer1_outputs(11504)));
    layer2_outputs(9656) <= not((layer1_outputs(872)) xor (layer1_outputs(11166)));
    layer2_outputs(9657) <= not(layer1_outputs(2955));
    layer2_outputs(9658) <= not(layer1_outputs(407)) or (layer1_outputs(4028));
    layer2_outputs(9659) <= layer1_outputs(9421);
    layer2_outputs(9660) <= not((layer1_outputs(9923)) xor (layer1_outputs(8223)));
    layer2_outputs(9661) <= not(layer1_outputs(6174));
    layer2_outputs(9662) <= layer1_outputs(11770);
    layer2_outputs(9663) <= not(layer1_outputs(6805)) or (layer1_outputs(7506));
    layer2_outputs(9664) <= not(layer1_outputs(2871)) or (layer1_outputs(4708));
    layer2_outputs(9665) <= not(layer1_outputs(10031)) or (layer1_outputs(3413));
    layer2_outputs(9666) <= (layer1_outputs(11485)) or (layer1_outputs(9552));
    layer2_outputs(9667) <= layer1_outputs(7645);
    layer2_outputs(9668) <= layer1_outputs(1677);
    layer2_outputs(9669) <= not((layer1_outputs(12298)) or (layer1_outputs(11148)));
    layer2_outputs(9670) <= layer1_outputs(5990);
    layer2_outputs(9671) <= (layer1_outputs(460)) and not (layer1_outputs(12527));
    layer2_outputs(9672) <= '0';
    layer2_outputs(9673) <= not(layer1_outputs(7367));
    layer2_outputs(9674) <= not(layer1_outputs(5343));
    layer2_outputs(9675) <= layer1_outputs(12607);
    layer2_outputs(9676) <= layer1_outputs(7218);
    layer2_outputs(9677) <= layer1_outputs(6800);
    layer2_outputs(9678) <= layer1_outputs(11729);
    layer2_outputs(9679) <= not(layer1_outputs(7865));
    layer2_outputs(9680) <= (layer1_outputs(4226)) and (layer1_outputs(5628));
    layer2_outputs(9681) <= layer1_outputs(8173);
    layer2_outputs(9682) <= not(layer1_outputs(6042)) or (layer1_outputs(7321));
    layer2_outputs(9683) <= layer1_outputs(11803);
    layer2_outputs(9684) <= layer1_outputs(4049);
    layer2_outputs(9685) <= (layer1_outputs(4190)) or (layer1_outputs(1518));
    layer2_outputs(9686) <= not(layer1_outputs(2214)) or (layer1_outputs(251));
    layer2_outputs(9687) <= (layer1_outputs(2291)) or (layer1_outputs(9506));
    layer2_outputs(9688) <= not(layer1_outputs(4179)) or (layer1_outputs(8493));
    layer2_outputs(9689) <= layer1_outputs(8617);
    layer2_outputs(9690) <= not(layer1_outputs(5454)) or (layer1_outputs(12674));
    layer2_outputs(9691) <= (layer1_outputs(1600)) and (layer1_outputs(5139));
    layer2_outputs(9692) <= not(layer1_outputs(3662));
    layer2_outputs(9693) <= layer1_outputs(40);
    layer2_outputs(9694) <= layer1_outputs(6410);
    layer2_outputs(9695) <= not((layer1_outputs(12150)) or (layer1_outputs(8240)));
    layer2_outputs(9696) <= layer1_outputs(9061);
    layer2_outputs(9697) <= not(layer1_outputs(11113));
    layer2_outputs(9698) <= not((layer1_outputs(7600)) and (layer1_outputs(2268)));
    layer2_outputs(9699) <= layer1_outputs(8631);
    layer2_outputs(9700) <= not(layer1_outputs(7552)) or (layer1_outputs(11307));
    layer2_outputs(9701) <= not(layer1_outputs(10172));
    layer2_outputs(9702) <= layer1_outputs(5653);
    layer2_outputs(9703) <= not(layer1_outputs(4872)) or (layer1_outputs(11554));
    layer2_outputs(9704) <= not(layer1_outputs(8739));
    layer2_outputs(9705) <= not(layer1_outputs(11282)) or (layer1_outputs(4559));
    layer2_outputs(9706) <= (layer1_outputs(7378)) and (layer1_outputs(9291));
    layer2_outputs(9707) <= not(layer1_outputs(10232));
    layer2_outputs(9708) <= (layer1_outputs(9846)) and not (layer1_outputs(1629));
    layer2_outputs(9709) <= (layer1_outputs(2727)) and not (layer1_outputs(5722));
    layer2_outputs(9710) <= not(layer1_outputs(977));
    layer2_outputs(9711) <= layer1_outputs(8119);
    layer2_outputs(9712) <= not(layer1_outputs(5910));
    layer2_outputs(9713) <= (layer1_outputs(4050)) and (layer1_outputs(5766));
    layer2_outputs(9714) <= not((layer1_outputs(1936)) or (layer1_outputs(3991)));
    layer2_outputs(9715) <= not(layer1_outputs(11252));
    layer2_outputs(9716) <= layer1_outputs(738);
    layer2_outputs(9717) <= (layer1_outputs(713)) or (layer1_outputs(9453));
    layer2_outputs(9718) <= not(layer1_outputs(4492)) or (layer1_outputs(6074));
    layer2_outputs(9719) <= layer1_outputs(1848);
    layer2_outputs(9720) <= (layer1_outputs(9989)) and not (layer1_outputs(8024));
    layer2_outputs(9721) <= not((layer1_outputs(11274)) xor (layer1_outputs(5928)));
    layer2_outputs(9722) <= not((layer1_outputs(3220)) xor (layer1_outputs(8459)));
    layer2_outputs(9723) <= not(layer1_outputs(5650));
    layer2_outputs(9724) <= (layer1_outputs(8486)) xor (layer1_outputs(12176));
    layer2_outputs(9725) <= not(layer1_outputs(4571));
    layer2_outputs(9726) <= (layer1_outputs(7190)) or (layer1_outputs(1537));
    layer2_outputs(9727) <= not((layer1_outputs(12581)) xor (layer1_outputs(9555)));
    layer2_outputs(9728) <= layer1_outputs(6399);
    layer2_outputs(9729) <= (layer1_outputs(1542)) and not (layer1_outputs(7667));
    layer2_outputs(9730) <= '0';
    layer2_outputs(9731) <= (layer1_outputs(3916)) xor (layer1_outputs(1411));
    layer2_outputs(9732) <= layer1_outputs(8708);
    layer2_outputs(9733) <= not(layer1_outputs(8048));
    layer2_outputs(9734) <= not(layer1_outputs(2146));
    layer2_outputs(9735) <= not(layer1_outputs(8372));
    layer2_outputs(9736) <= not(layer1_outputs(1413));
    layer2_outputs(9737) <= layer1_outputs(2260);
    layer2_outputs(9738) <= not(layer1_outputs(8738));
    layer2_outputs(9739) <= not(layer1_outputs(514));
    layer2_outputs(9740) <= not(layer1_outputs(5940));
    layer2_outputs(9741) <= not(layer1_outputs(11857));
    layer2_outputs(9742) <= not((layer1_outputs(1544)) and (layer1_outputs(5709)));
    layer2_outputs(9743) <= not((layer1_outputs(12747)) or (layer1_outputs(4142)));
    layer2_outputs(9744) <= not(layer1_outputs(7827));
    layer2_outputs(9745) <= not((layer1_outputs(3857)) xor (layer1_outputs(3490)));
    layer2_outputs(9746) <= not((layer1_outputs(3175)) xor (layer1_outputs(10478)));
    layer2_outputs(9747) <= not(layer1_outputs(12142));
    layer2_outputs(9748) <= not((layer1_outputs(625)) xor (layer1_outputs(2818)));
    layer2_outputs(9749) <= not(layer1_outputs(3286));
    layer2_outputs(9750) <= not(layer1_outputs(3621));
    layer2_outputs(9751) <= layer1_outputs(6923);
    layer2_outputs(9752) <= layer1_outputs(8063);
    layer2_outputs(9753) <= not(layer1_outputs(8339));
    layer2_outputs(9754) <= not((layer1_outputs(11224)) or (layer1_outputs(3550)));
    layer2_outputs(9755) <= (layer1_outputs(1479)) xor (layer1_outputs(1664));
    layer2_outputs(9756) <= not(layer1_outputs(12242));
    layer2_outputs(9757) <= not(layer1_outputs(4288));
    layer2_outputs(9758) <= not(layer1_outputs(3185)) or (layer1_outputs(2702));
    layer2_outputs(9759) <= layer1_outputs(6036);
    layer2_outputs(9760) <= not(layer1_outputs(7365));
    layer2_outputs(9761) <= layer1_outputs(10809);
    layer2_outputs(9762) <= layer1_outputs(212);
    layer2_outputs(9763) <= (layer1_outputs(12188)) and (layer1_outputs(6361));
    layer2_outputs(9764) <= layer1_outputs(761);
    layer2_outputs(9765) <= not(layer1_outputs(3790));
    layer2_outputs(9766) <= layer1_outputs(1994);
    layer2_outputs(9767) <= layer1_outputs(4195);
    layer2_outputs(9768) <= (layer1_outputs(12546)) xor (layer1_outputs(2655));
    layer2_outputs(9769) <= not(layer1_outputs(10229));
    layer2_outputs(9770) <= layer1_outputs(4599);
    layer2_outputs(9771) <= (layer1_outputs(5633)) and (layer1_outputs(631));
    layer2_outputs(9772) <= not(layer1_outputs(6532));
    layer2_outputs(9773) <= not(layer1_outputs(10553));
    layer2_outputs(9774) <= layer1_outputs(8526);
    layer2_outputs(9775) <= not(layer1_outputs(5737));
    layer2_outputs(9776) <= not((layer1_outputs(3376)) or (layer1_outputs(9207)));
    layer2_outputs(9777) <= not((layer1_outputs(4452)) xor (layer1_outputs(12726)));
    layer2_outputs(9778) <= layer1_outputs(8674);
    layer2_outputs(9779) <= layer1_outputs(3800);
    layer2_outputs(9780) <= not(layer1_outputs(6636)) or (layer1_outputs(362));
    layer2_outputs(9781) <= not((layer1_outputs(8762)) xor (layer1_outputs(520)));
    layer2_outputs(9782) <= layer1_outputs(1416);
    layer2_outputs(9783) <= (layer1_outputs(8586)) xor (layer1_outputs(10739));
    layer2_outputs(9784) <= (layer1_outputs(4286)) and not (layer1_outputs(11089));
    layer2_outputs(9785) <= (layer1_outputs(9309)) and not (layer1_outputs(11937));
    layer2_outputs(9786) <= not(layer1_outputs(4668));
    layer2_outputs(9787) <= layer1_outputs(9308);
    layer2_outputs(9788) <= (layer1_outputs(1804)) and not (layer1_outputs(6089));
    layer2_outputs(9789) <= (layer1_outputs(2118)) and not (layer1_outputs(11045));
    layer2_outputs(9790) <= (layer1_outputs(3909)) and (layer1_outputs(5401));
    layer2_outputs(9791) <= (layer1_outputs(9031)) and not (layer1_outputs(8025));
    layer2_outputs(9792) <= (layer1_outputs(4038)) xor (layer1_outputs(6223));
    layer2_outputs(9793) <= (layer1_outputs(4341)) and (layer1_outputs(10595));
    layer2_outputs(9794) <= (layer1_outputs(8214)) and not (layer1_outputs(9264));
    layer2_outputs(9795) <= not((layer1_outputs(733)) or (layer1_outputs(12484)));
    layer2_outputs(9796) <= not(layer1_outputs(3464)) or (layer1_outputs(6883));
    layer2_outputs(9797) <= (layer1_outputs(7630)) and not (layer1_outputs(10537));
    layer2_outputs(9798) <= not(layer1_outputs(3690));
    layer2_outputs(9799) <= (layer1_outputs(8404)) and not (layer1_outputs(1123));
    layer2_outputs(9800) <= (layer1_outputs(8831)) and (layer1_outputs(5935));
    layer2_outputs(9801) <= not((layer1_outputs(5529)) xor (layer1_outputs(2674)));
    layer2_outputs(9802) <= not(layer1_outputs(11197));
    layer2_outputs(9803) <= not(layer1_outputs(7436));
    layer2_outputs(9804) <= not(layer1_outputs(2362)) or (layer1_outputs(569));
    layer2_outputs(9805) <= not(layer1_outputs(11901)) or (layer1_outputs(12446));
    layer2_outputs(9806) <= layer1_outputs(2009);
    layer2_outputs(9807) <= not(layer1_outputs(11715));
    layer2_outputs(9808) <= not(layer1_outputs(6187)) or (layer1_outputs(3980));
    layer2_outputs(9809) <= (layer1_outputs(5149)) xor (layer1_outputs(4752));
    layer2_outputs(9810) <= not((layer1_outputs(2071)) or (layer1_outputs(10890)));
    layer2_outputs(9811) <= (layer1_outputs(2053)) and not (layer1_outputs(4437));
    layer2_outputs(9812) <= not(layer1_outputs(640));
    layer2_outputs(9813) <= not((layer1_outputs(7580)) or (layer1_outputs(5631)));
    layer2_outputs(9814) <= layer1_outputs(8284);
    layer2_outputs(9815) <= not(layer1_outputs(12008));
    layer2_outputs(9816) <= (layer1_outputs(8406)) and not (layer1_outputs(8512));
    layer2_outputs(9817) <= (layer1_outputs(2804)) and not (layer1_outputs(8199));
    layer2_outputs(9818) <= (layer1_outputs(8698)) and (layer1_outputs(7006));
    layer2_outputs(9819) <= layer1_outputs(4460);
    layer2_outputs(9820) <= not(layer1_outputs(5217));
    layer2_outputs(9821) <= not((layer1_outputs(11130)) xor (layer1_outputs(5977)));
    layer2_outputs(9822) <= not((layer1_outputs(6008)) or (layer1_outputs(7465)));
    layer2_outputs(9823) <= (layer1_outputs(558)) or (layer1_outputs(1146));
    layer2_outputs(9824) <= not(layer1_outputs(1828)) or (layer1_outputs(5671));
    layer2_outputs(9825) <= (layer1_outputs(11244)) and not (layer1_outputs(5448));
    layer2_outputs(9826) <= not(layer1_outputs(11386));
    layer2_outputs(9827) <= not((layer1_outputs(7336)) xor (layer1_outputs(6466)));
    layer2_outputs(9828) <= not(layer1_outputs(8169)) or (layer1_outputs(5736));
    layer2_outputs(9829) <= layer1_outputs(6186);
    layer2_outputs(9830) <= layer1_outputs(6426);
    layer2_outputs(9831) <= not(layer1_outputs(4239)) or (layer1_outputs(11621));
    layer2_outputs(9832) <= layer1_outputs(12397);
    layer2_outputs(9833) <= (layer1_outputs(10642)) and not (layer1_outputs(3739));
    layer2_outputs(9834) <= not((layer1_outputs(8176)) or (layer1_outputs(5619)));
    layer2_outputs(9835) <= (layer1_outputs(9032)) and (layer1_outputs(12745));
    layer2_outputs(9836) <= '0';
    layer2_outputs(9837) <= not(layer1_outputs(12199));
    layer2_outputs(9838) <= not(layer1_outputs(2100));
    layer2_outputs(9839) <= layer1_outputs(7120);
    layer2_outputs(9840) <= not(layer1_outputs(8672)) or (layer1_outputs(670));
    layer2_outputs(9841) <= not(layer1_outputs(1957));
    layer2_outputs(9842) <= (layer1_outputs(1384)) and (layer1_outputs(6362));
    layer2_outputs(9843) <= (layer1_outputs(9124)) xor (layer1_outputs(3169));
    layer2_outputs(9844) <= (layer1_outputs(10835)) xor (layer1_outputs(2366));
    layer2_outputs(9845) <= layer1_outputs(565);
    layer2_outputs(9846) <= not(layer1_outputs(10106));
    layer2_outputs(9847) <= (layer1_outputs(10677)) xor (layer1_outputs(5389));
    layer2_outputs(9848) <= '1';
    layer2_outputs(9849) <= not(layer1_outputs(7204)) or (layer1_outputs(5387));
    layer2_outputs(9850) <= layer1_outputs(6157);
    layer2_outputs(9851) <= (layer1_outputs(10272)) and (layer1_outputs(3771));
    layer2_outputs(9852) <= not(layer1_outputs(3822));
    layer2_outputs(9853) <= (layer1_outputs(10698)) xor (layer1_outputs(87));
    layer2_outputs(9854) <= not(layer1_outputs(1866)) or (layer1_outputs(3977));
    layer2_outputs(9855) <= (layer1_outputs(3545)) and not (layer1_outputs(5939));
    layer2_outputs(9856) <= not((layer1_outputs(6663)) xor (layer1_outputs(2299)));
    layer2_outputs(9857) <= (layer1_outputs(8168)) xor (layer1_outputs(12186));
    layer2_outputs(9858) <= not(layer1_outputs(7300));
    layer2_outputs(9859) <= (layer1_outputs(11175)) xor (layer1_outputs(10488));
    layer2_outputs(9860) <= (layer1_outputs(5920)) and not (layer1_outputs(5800));
    layer2_outputs(9861) <= (layer1_outputs(5607)) xor (layer1_outputs(4568));
    layer2_outputs(9862) <= not((layer1_outputs(89)) xor (layer1_outputs(3590)));
    layer2_outputs(9863) <= layer1_outputs(11870);
    layer2_outputs(9864) <= not(layer1_outputs(11570)) or (layer1_outputs(5401));
    layer2_outputs(9865) <= not(layer1_outputs(12712));
    layer2_outputs(9866) <= not((layer1_outputs(5281)) xor (layer1_outputs(11247)));
    layer2_outputs(9867) <= not(layer1_outputs(575));
    layer2_outputs(9868) <= layer1_outputs(3175);
    layer2_outputs(9869) <= layer1_outputs(8077);
    layer2_outputs(9870) <= (layer1_outputs(9197)) and (layer1_outputs(12597));
    layer2_outputs(9871) <= (layer1_outputs(10699)) and not (layer1_outputs(5323));
    layer2_outputs(9872) <= (layer1_outputs(12185)) or (layer1_outputs(143));
    layer2_outputs(9873) <= not(layer1_outputs(6709));
    layer2_outputs(9874) <= not(layer1_outputs(793));
    layer2_outputs(9875) <= not((layer1_outputs(9475)) or (layer1_outputs(5996)));
    layer2_outputs(9876) <= not(layer1_outputs(8841)) or (layer1_outputs(58));
    layer2_outputs(9877) <= not(layer1_outputs(132));
    layer2_outputs(9878) <= not((layer1_outputs(10945)) and (layer1_outputs(1980)));
    layer2_outputs(9879) <= not((layer1_outputs(7612)) xor (layer1_outputs(1474)));
    layer2_outputs(9880) <= (layer1_outputs(4530)) and (layer1_outputs(9632));
    layer2_outputs(9881) <= (layer1_outputs(42)) and not (layer1_outputs(7012));
    layer2_outputs(9882) <= not(layer1_outputs(5423));
    layer2_outputs(9883) <= not((layer1_outputs(7009)) xor (layer1_outputs(10722)));
    layer2_outputs(9884) <= not(layer1_outputs(3089));
    layer2_outputs(9885) <= not((layer1_outputs(8924)) and (layer1_outputs(78)));
    layer2_outputs(9886) <= (layer1_outputs(1402)) or (layer1_outputs(4578));
    layer2_outputs(9887) <= not(layer1_outputs(3546));
    layer2_outputs(9888) <= not(layer1_outputs(6616));
    layer2_outputs(9889) <= (layer1_outputs(1337)) and not (layer1_outputs(7413));
    layer2_outputs(9890) <= not(layer1_outputs(3913)) or (layer1_outputs(11339));
    layer2_outputs(9891) <= not(layer1_outputs(5600));
    layer2_outputs(9892) <= not(layer1_outputs(12383));
    layer2_outputs(9893) <= layer1_outputs(8328);
    layer2_outputs(9894) <= not((layer1_outputs(88)) or (layer1_outputs(252)));
    layer2_outputs(9895) <= not(layer1_outputs(5434));
    layer2_outputs(9896) <= (layer1_outputs(9266)) or (layer1_outputs(11030));
    layer2_outputs(9897) <= not(layer1_outputs(3874));
    layer2_outputs(9898) <= (layer1_outputs(10354)) xor (layer1_outputs(2666));
    layer2_outputs(9899) <= not((layer1_outputs(10919)) xor (layer1_outputs(8418)));
    layer2_outputs(9900) <= not(layer1_outputs(8066));
    layer2_outputs(9901) <= not(layer1_outputs(2598));
    layer2_outputs(9902) <= not(layer1_outputs(4356));
    layer2_outputs(9903) <= not(layer1_outputs(446));
    layer2_outputs(9904) <= layer1_outputs(8138);
    layer2_outputs(9905) <= not(layer1_outputs(5924));
    layer2_outputs(9906) <= (layer1_outputs(7833)) and not (layer1_outputs(1612));
    layer2_outputs(9907) <= (layer1_outputs(3949)) and (layer1_outputs(7837));
    layer2_outputs(9908) <= (layer1_outputs(12587)) and not (layer1_outputs(8761));
    layer2_outputs(9909) <= layer1_outputs(4201);
    layer2_outputs(9910) <= layer1_outputs(1579);
    layer2_outputs(9911) <= layer1_outputs(11857);
    layer2_outputs(9912) <= not(layer1_outputs(10332));
    layer2_outputs(9913) <= layer1_outputs(5896);
    layer2_outputs(9914) <= not(layer1_outputs(10482));
    layer2_outputs(9915) <= (layer1_outputs(6737)) and not (layer1_outputs(7351));
    layer2_outputs(9916) <= (layer1_outputs(5783)) or (layer1_outputs(7337));
    layer2_outputs(9917) <= not(layer1_outputs(1003));
    layer2_outputs(9918) <= not(layer1_outputs(12055)) or (layer1_outputs(6351));
    layer2_outputs(9919) <= (layer1_outputs(1234)) or (layer1_outputs(6208));
    layer2_outputs(9920) <= not(layer1_outputs(3415));
    layer2_outputs(9921) <= '1';
    layer2_outputs(9922) <= not(layer1_outputs(3805)) or (layer1_outputs(295));
    layer2_outputs(9923) <= not((layer1_outputs(11962)) and (layer1_outputs(2980)));
    layer2_outputs(9924) <= not(layer1_outputs(8129)) or (layer1_outputs(6987));
    layer2_outputs(9925) <= not((layer1_outputs(12167)) or (layer1_outputs(11279)));
    layer2_outputs(9926) <= (layer1_outputs(9214)) and (layer1_outputs(12323));
    layer2_outputs(9927) <= not(layer1_outputs(5465)) or (layer1_outputs(10813));
    layer2_outputs(9928) <= layer1_outputs(5667);
    layer2_outputs(9929) <= (layer1_outputs(9570)) xor (layer1_outputs(9023));
    layer2_outputs(9930) <= layer1_outputs(11259);
    layer2_outputs(9931) <= not(layer1_outputs(8816));
    layer2_outputs(9932) <= not(layer1_outputs(2830));
    layer2_outputs(9933) <= (layer1_outputs(12624)) and not (layer1_outputs(7666));
    layer2_outputs(9934) <= not(layer1_outputs(2948));
    layer2_outputs(9935) <= (layer1_outputs(4351)) xor (layer1_outputs(1478));
    layer2_outputs(9936) <= (layer1_outputs(5397)) and not (layer1_outputs(10496));
    layer2_outputs(9937) <= not(layer1_outputs(6892));
    layer2_outputs(9938) <= layer1_outputs(10014);
    layer2_outputs(9939) <= (layer1_outputs(3152)) xor (layer1_outputs(12509));
    layer2_outputs(9940) <= (layer1_outputs(3189)) and not (layer1_outputs(7635));
    layer2_outputs(9941) <= layer1_outputs(8929);
    layer2_outputs(9942) <= not(layer1_outputs(4801));
    layer2_outputs(9943) <= (layer1_outputs(1787)) or (layer1_outputs(10465));
    layer2_outputs(9944) <= not(layer1_outputs(10879));
    layer2_outputs(9945) <= (layer1_outputs(5668)) and (layer1_outputs(6722));
    layer2_outputs(9946) <= (layer1_outputs(10099)) xor (layer1_outputs(12550));
    layer2_outputs(9947) <= layer1_outputs(4503);
    layer2_outputs(9948) <= (layer1_outputs(278)) and (layer1_outputs(3358));
    layer2_outputs(9949) <= not(layer1_outputs(3817));
    layer2_outputs(9950) <= (layer1_outputs(12233)) and (layer1_outputs(11488));
    layer2_outputs(9951) <= layer1_outputs(1039);
    layer2_outputs(9952) <= (layer1_outputs(12286)) and (layer1_outputs(2982));
    layer2_outputs(9953) <= not(layer1_outputs(7817)) or (layer1_outputs(7385));
    layer2_outputs(9954) <= not((layer1_outputs(2464)) xor (layer1_outputs(3486)));
    layer2_outputs(9955) <= not((layer1_outputs(6566)) and (layer1_outputs(140)));
    layer2_outputs(9956) <= not(layer1_outputs(5538));
    layer2_outputs(9957) <= not(layer1_outputs(9041));
    layer2_outputs(9958) <= (layer1_outputs(896)) xor (layer1_outputs(860));
    layer2_outputs(9959) <= not((layer1_outputs(5752)) xor (layer1_outputs(1742)));
    layer2_outputs(9960) <= layer1_outputs(9986);
    layer2_outputs(9961) <= not(layer1_outputs(2376));
    layer2_outputs(9962) <= (layer1_outputs(6584)) and not (layer1_outputs(3164));
    layer2_outputs(9963) <= not(layer1_outputs(7923));
    layer2_outputs(9964) <= (layer1_outputs(4106)) and not (layer1_outputs(2837));
    layer2_outputs(9965) <= (layer1_outputs(9086)) xor (layer1_outputs(7739));
    layer2_outputs(9966) <= layer1_outputs(5437);
    layer2_outputs(9967) <= not(layer1_outputs(1219)) or (layer1_outputs(4464));
    layer2_outputs(9968) <= layer1_outputs(2125);
    layer2_outputs(9969) <= layer1_outputs(10861);
    layer2_outputs(9970) <= layer1_outputs(234);
    layer2_outputs(9971) <= (layer1_outputs(3640)) and not (layer1_outputs(11068));
    layer2_outputs(9972) <= not((layer1_outputs(3039)) xor (layer1_outputs(1186)));
    layer2_outputs(9973) <= layer1_outputs(8782);
    layer2_outputs(9974) <= layer1_outputs(3270);
    layer2_outputs(9975) <= layer1_outputs(206);
    layer2_outputs(9976) <= not((layer1_outputs(7697)) or (layer1_outputs(11963)));
    layer2_outputs(9977) <= not(layer1_outputs(5578)) or (layer1_outputs(6353));
    layer2_outputs(9978) <= layer1_outputs(3703);
    layer2_outputs(9979) <= not((layer1_outputs(11973)) xor (layer1_outputs(4497)));
    layer2_outputs(9980) <= not(layer1_outputs(10860));
    layer2_outputs(9981) <= (layer1_outputs(12115)) or (layer1_outputs(5037));
    layer2_outputs(9982) <= (layer1_outputs(2666)) xor (layer1_outputs(7871));
    layer2_outputs(9983) <= not(layer1_outputs(432)) or (layer1_outputs(2163));
    layer2_outputs(9984) <= not((layer1_outputs(11285)) and (layer1_outputs(888)));
    layer2_outputs(9985) <= (layer1_outputs(8954)) and (layer1_outputs(6885));
    layer2_outputs(9986) <= layer1_outputs(11481);
    layer2_outputs(9987) <= layer1_outputs(340);
    layer2_outputs(9988) <= layer1_outputs(10755);
    layer2_outputs(9989) <= not((layer1_outputs(2453)) xor (layer1_outputs(6402)));
    layer2_outputs(9990) <= not(layer1_outputs(7184));
    layer2_outputs(9991) <= (layer1_outputs(3035)) and not (layer1_outputs(1355));
    layer2_outputs(9992) <= layer1_outputs(6934);
    layer2_outputs(9993) <= not(layer1_outputs(676)) or (layer1_outputs(11253));
    layer2_outputs(9994) <= not(layer1_outputs(6931));
    layer2_outputs(9995) <= layer1_outputs(1539);
    layer2_outputs(9996) <= layer1_outputs(4192);
    layer2_outputs(9997) <= not((layer1_outputs(5410)) xor (layer1_outputs(7804)));
    layer2_outputs(9998) <= not((layer1_outputs(468)) and (layer1_outputs(1423)));
    layer2_outputs(9999) <= (layer1_outputs(8261)) and not (layer1_outputs(7402));
    layer2_outputs(10000) <= not(layer1_outputs(8959));
    layer2_outputs(10001) <= (layer1_outputs(7506)) and (layer1_outputs(1397));
    layer2_outputs(10002) <= not(layer1_outputs(9786));
    layer2_outputs(10003) <= (layer1_outputs(1005)) and not (layer1_outputs(11130));
    layer2_outputs(10004) <= layer1_outputs(9969);
    layer2_outputs(10005) <= layer1_outputs(3721);
    layer2_outputs(10006) <= not(layer1_outputs(2215)) or (layer1_outputs(7199));
    layer2_outputs(10007) <= not(layer1_outputs(10387)) or (layer1_outputs(6293));
    layer2_outputs(10008) <= (layer1_outputs(9075)) or (layer1_outputs(173));
    layer2_outputs(10009) <= (layer1_outputs(341)) and (layer1_outputs(2404));
    layer2_outputs(10010) <= not(layer1_outputs(12679));
    layer2_outputs(10011) <= layer1_outputs(7828);
    layer2_outputs(10012) <= (layer1_outputs(1053)) and (layer1_outputs(1852));
    layer2_outputs(10013) <= (layer1_outputs(3147)) and not (layer1_outputs(4850));
    layer2_outputs(10014) <= not(layer1_outputs(1093));
    layer2_outputs(10015) <= layer1_outputs(10573);
    layer2_outputs(10016) <= layer1_outputs(3418);
    layer2_outputs(10017) <= (layer1_outputs(9220)) and not (layer1_outputs(5216));
    layer2_outputs(10018) <= not(layer1_outputs(6917));
    layer2_outputs(10019) <= (layer1_outputs(5986)) and not (layer1_outputs(4701));
    layer2_outputs(10020) <= (layer1_outputs(4366)) and not (layer1_outputs(4018));
    layer2_outputs(10021) <= (layer1_outputs(7320)) and not (layer1_outputs(1863));
    layer2_outputs(10022) <= layer1_outputs(1476);
    layer2_outputs(10023) <= not((layer1_outputs(3354)) xor (layer1_outputs(2366)));
    layer2_outputs(10024) <= layer1_outputs(5616);
    layer2_outputs(10025) <= not(layer1_outputs(8768));
    layer2_outputs(10026) <= (layer1_outputs(1892)) or (layer1_outputs(198));
    layer2_outputs(10027) <= not((layer1_outputs(4383)) or (layer1_outputs(10875)));
    layer2_outputs(10028) <= layer1_outputs(6627);
    layer2_outputs(10029) <= not(layer1_outputs(1975)) or (layer1_outputs(9333));
    layer2_outputs(10030) <= not((layer1_outputs(7144)) xor (layer1_outputs(1635)));
    layer2_outputs(10031) <= (layer1_outputs(513)) xor (layer1_outputs(6142));
    layer2_outputs(10032) <= (layer1_outputs(9241)) or (layer1_outputs(3417));
    layer2_outputs(10033) <= layer1_outputs(3787);
    layer2_outputs(10034) <= not((layer1_outputs(5270)) xor (layer1_outputs(2375)));
    layer2_outputs(10035) <= not(layer1_outputs(4966));
    layer2_outputs(10036) <= not((layer1_outputs(1420)) and (layer1_outputs(8355)));
    layer2_outputs(10037) <= not(layer1_outputs(449)) or (layer1_outputs(3126));
    layer2_outputs(10038) <= layer1_outputs(6934);
    layer2_outputs(10039) <= not(layer1_outputs(6677)) or (layer1_outputs(5526));
    layer2_outputs(10040) <= (layer1_outputs(2421)) and not (layer1_outputs(10943));
    layer2_outputs(10041) <= (layer1_outputs(8557)) or (layer1_outputs(12123));
    layer2_outputs(10042) <= layer1_outputs(10603);
    layer2_outputs(10043) <= not(layer1_outputs(8318));
    layer2_outputs(10044) <= not(layer1_outputs(1260));
    layer2_outputs(10045) <= not(layer1_outputs(3650)) or (layer1_outputs(11929));
    layer2_outputs(10046) <= (layer1_outputs(6343)) or (layer1_outputs(4027));
    layer2_outputs(10047) <= not((layer1_outputs(1718)) or (layer1_outputs(2215)));
    layer2_outputs(10048) <= not((layer1_outputs(4965)) and (layer1_outputs(2392)));
    layer2_outputs(10049) <= not(layer1_outputs(2970));
    layer2_outputs(10050) <= layer1_outputs(1694);
    layer2_outputs(10051) <= not(layer1_outputs(12535));
    layer2_outputs(10052) <= not(layer1_outputs(1692));
    layer2_outputs(10053) <= not(layer1_outputs(3794));
    layer2_outputs(10054) <= layer1_outputs(9994);
    layer2_outputs(10055) <= (layer1_outputs(12212)) and not (layer1_outputs(8677));
    layer2_outputs(10056) <= not(layer1_outputs(2769));
    layer2_outputs(10057) <= layer1_outputs(5481);
    layer2_outputs(10058) <= (layer1_outputs(7010)) and (layer1_outputs(3333));
    layer2_outputs(10059) <= (layer1_outputs(11054)) xor (layer1_outputs(4577));
    layer2_outputs(10060) <= layer1_outputs(8264);
    layer2_outputs(10061) <= not(layer1_outputs(12178));
    layer2_outputs(10062) <= not(layer1_outputs(7225));
    layer2_outputs(10063) <= layer1_outputs(10133);
    layer2_outputs(10064) <= (layer1_outputs(5455)) xor (layer1_outputs(10615));
    layer2_outputs(10065) <= layer1_outputs(11555);
    layer2_outputs(10066) <= not(layer1_outputs(152));
    layer2_outputs(10067) <= (layer1_outputs(2239)) xor (layer1_outputs(2232));
    layer2_outputs(10068) <= (layer1_outputs(7876)) and not (layer1_outputs(90));
    layer2_outputs(10069) <= (layer1_outputs(6671)) and not (layer1_outputs(339));
    layer2_outputs(10070) <= not(layer1_outputs(10458));
    layer2_outputs(10071) <= layer1_outputs(5609);
    layer2_outputs(10072) <= (layer1_outputs(6242)) and not (layer1_outputs(3576));
    layer2_outputs(10073) <= not((layer1_outputs(3902)) or (layer1_outputs(1460)));
    layer2_outputs(10074) <= layer1_outputs(7631);
    layer2_outputs(10075) <= not(layer1_outputs(6463));
    layer2_outputs(10076) <= (layer1_outputs(9731)) or (layer1_outputs(11471));
    layer2_outputs(10077) <= (layer1_outputs(3124)) and not (layer1_outputs(12141));
    layer2_outputs(10078) <= not((layer1_outputs(367)) or (layer1_outputs(5439)));
    layer2_outputs(10079) <= not(layer1_outputs(9348));
    layer2_outputs(10080) <= layer1_outputs(8777);
    layer2_outputs(10081) <= layer1_outputs(12146);
    layer2_outputs(10082) <= (layer1_outputs(592)) and not (layer1_outputs(3125));
    layer2_outputs(10083) <= (layer1_outputs(790)) xor (layer1_outputs(4065));
    layer2_outputs(10084) <= (layer1_outputs(1084)) and not (layer1_outputs(4509));
    layer2_outputs(10085) <= (layer1_outputs(5485)) and not (layer1_outputs(8042));
    layer2_outputs(10086) <= not(layer1_outputs(4300));
    layer2_outputs(10087) <= not((layer1_outputs(101)) xor (layer1_outputs(8584)));
    layer2_outputs(10088) <= (layer1_outputs(4444)) or (layer1_outputs(9694));
    layer2_outputs(10089) <= not((layer1_outputs(3920)) xor (layer1_outputs(9529)));
    layer2_outputs(10090) <= (layer1_outputs(4099)) xor (layer1_outputs(10347));
    layer2_outputs(10091) <= not((layer1_outputs(11891)) and (layer1_outputs(5755)));
    layer2_outputs(10092) <= not(layer1_outputs(2750));
    layer2_outputs(10093) <= not(layer1_outputs(1597));
    layer2_outputs(10094) <= not(layer1_outputs(1895)) or (layer1_outputs(10775));
    layer2_outputs(10095) <= not(layer1_outputs(235));
    layer2_outputs(10096) <= not((layer1_outputs(5729)) and (layer1_outputs(3690)));
    layer2_outputs(10097) <= (layer1_outputs(8506)) xor (layer1_outputs(11986));
    layer2_outputs(10098) <= layer1_outputs(9404);
    layer2_outputs(10099) <= not(layer1_outputs(1997)) or (layer1_outputs(11202));
    layer2_outputs(10100) <= not(layer1_outputs(8855)) or (layer1_outputs(10160));
    layer2_outputs(10101) <= layer1_outputs(2757);
    layer2_outputs(10102) <= layer1_outputs(10668);
    layer2_outputs(10103) <= layer1_outputs(11998);
    layer2_outputs(10104) <= (layer1_outputs(7363)) and (layer1_outputs(4988));
    layer2_outputs(10105) <= '1';
    layer2_outputs(10106) <= layer1_outputs(12159);
    layer2_outputs(10107) <= (layer1_outputs(9340)) or (layer1_outputs(782));
    layer2_outputs(10108) <= layer1_outputs(1509);
    layer2_outputs(10109) <= layer1_outputs(1641);
    layer2_outputs(10110) <= not(layer1_outputs(2030));
    layer2_outputs(10111) <= (layer1_outputs(2815)) or (layer1_outputs(10252));
    layer2_outputs(10112) <= (layer1_outputs(7830)) and (layer1_outputs(9832));
    layer2_outputs(10113) <= not((layer1_outputs(1768)) and (layer1_outputs(3598)));
    layer2_outputs(10114) <= not(layer1_outputs(156));
    layer2_outputs(10115) <= not(layer1_outputs(1949)) or (layer1_outputs(11633));
    layer2_outputs(10116) <= not(layer1_outputs(6909)) or (layer1_outputs(7019));
    layer2_outputs(10117) <= (layer1_outputs(6144)) and (layer1_outputs(5346));
    layer2_outputs(10118) <= layer1_outputs(3378);
    layer2_outputs(10119) <= layer1_outputs(1825);
    layer2_outputs(10120) <= not((layer1_outputs(7733)) xor (layer1_outputs(8649)));
    layer2_outputs(10121) <= (layer1_outputs(5898)) xor (layer1_outputs(5588));
    layer2_outputs(10122) <= (layer1_outputs(8475)) xor (layer1_outputs(11585));
    layer2_outputs(10123) <= not((layer1_outputs(4794)) xor (layer1_outputs(11295)));
    layer2_outputs(10124) <= (layer1_outputs(1745)) and (layer1_outputs(8143));
    layer2_outputs(10125) <= layer1_outputs(11666);
    layer2_outputs(10126) <= (layer1_outputs(3989)) xor (layer1_outputs(8065));
    layer2_outputs(10127) <= '0';
    layer2_outputs(10128) <= layer1_outputs(12407);
    layer2_outputs(10129) <= (layer1_outputs(5976)) xor (layer1_outputs(6852));
    layer2_outputs(10130) <= not(layer1_outputs(4627));
    layer2_outputs(10131) <= not(layer1_outputs(4084));
    layer2_outputs(10132) <= not(layer1_outputs(3038));
    layer2_outputs(10133) <= layer1_outputs(10418);
    layer2_outputs(10134) <= layer1_outputs(11325);
    layer2_outputs(10135) <= layer1_outputs(3499);
    layer2_outputs(10136) <= not(layer1_outputs(12734));
    layer2_outputs(10137) <= (layer1_outputs(7915)) and not (layer1_outputs(12264));
    layer2_outputs(10138) <= '0';
    layer2_outputs(10139) <= (layer1_outputs(5452)) and not (layer1_outputs(1260));
    layer2_outputs(10140) <= (layer1_outputs(7431)) xor (layer1_outputs(9140));
    layer2_outputs(10141) <= not((layer1_outputs(12110)) xor (layer1_outputs(11417)));
    layer2_outputs(10142) <= layer1_outputs(940);
    layer2_outputs(10143) <= (layer1_outputs(11515)) xor (layer1_outputs(8523));
    layer2_outputs(10144) <= not(layer1_outputs(5517));
    layer2_outputs(10145) <= not((layer1_outputs(5135)) xor (layer1_outputs(1197)));
    layer2_outputs(10146) <= layer1_outputs(7541);
    layer2_outputs(10147) <= layer1_outputs(9839);
    layer2_outputs(10148) <= not(layer1_outputs(3905)) or (layer1_outputs(9623));
    layer2_outputs(10149) <= not(layer1_outputs(6346)) or (layer1_outputs(11304));
    layer2_outputs(10150) <= not(layer1_outputs(3784));
    layer2_outputs(10151) <= layer1_outputs(10503);
    layer2_outputs(10152) <= not(layer1_outputs(4203));
    layer2_outputs(10153) <= layer1_outputs(1465);
    layer2_outputs(10154) <= not(layer1_outputs(910));
    layer2_outputs(10155) <= layer1_outputs(372);
    layer2_outputs(10156) <= not((layer1_outputs(9172)) and (layer1_outputs(4662)));
    layer2_outputs(10157) <= not(layer1_outputs(8229));
    layer2_outputs(10158) <= not(layer1_outputs(62)) or (layer1_outputs(4955));
    layer2_outputs(10159) <= not(layer1_outputs(162));
    layer2_outputs(10160) <= (layer1_outputs(2458)) xor (layer1_outputs(1714));
    layer2_outputs(10161) <= (layer1_outputs(9528)) or (layer1_outputs(9831));
    layer2_outputs(10162) <= not(layer1_outputs(10652));
    layer2_outputs(10163) <= not(layer1_outputs(9026));
    layer2_outputs(10164) <= not((layer1_outputs(5643)) and (layer1_outputs(3560)));
    layer2_outputs(10165) <= not(layer1_outputs(6879));
    layer2_outputs(10166) <= layer1_outputs(10837);
    layer2_outputs(10167) <= layer1_outputs(11287);
    layer2_outputs(10168) <= layer1_outputs(12652);
    layer2_outputs(10169) <= (layer1_outputs(8341)) and not (layer1_outputs(11392));
    layer2_outputs(10170) <= not((layer1_outputs(3553)) or (layer1_outputs(6678)));
    layer2_outputs(10171) <= not(layer1_outputs(12205));
    layer2_outputs(10172) <= layer1_outputs(7985);
    layer2_outputs(10173) <= (layer1_outputs(8320)) xor (layer1_outputs(2168));
    layer2_outputs(10174) <= (layer1_outputs(897)) and not (layer1_outputs(4348));
    layer2_outputs(10175) <= not(layer1_outputs(5742)) or (layer1_outputs(6101));
    layer2_outputs(10176) <= not(layer1_outputs(7141));
    layer2_outputs(10177) <= layer1_outputs(1843);
    layer2_outputs(10178) <= not(layer1_outputs(6494));
    layer2_outputs(10179) <= (layer1_outputs(10052)) or (layer1_outputs(10353));
    layer2_outputs(10180) <= not(layer1_outputs(6970)) or (layer1_outputs(8333));
    layer2_outputs(10181) <= (layer1_outputs(1256)) and not (layer1_outputs(7286));
    layer2_outputs(10182) <= not(layer1_outputs(12316)) or (layer1_outputs(8297));
    layer2_outputs(10183) <= (layer1_outputs(5186)) and (layer1_outputs(3344));
    layer2_outputs(10184) <= layer1_outputs(465);
    layer2_outputs(10185) <= (layer1_outputs(7211)) xor (layer1_outputs(3327));
    layer2_outputs(10186) <= not(layer1_outputs(9454));
    layer2_outputs(10187) <= layer1_outputs(6480);
    layer2_outputs(10188) <= not(layer1_outputs(11395));
    layer2_outputs(10189) <= (layer1_outputs(7495)) and not (layer1_outputs(4867));
    layer2_outputs(10190) <= layer1_outputs(636);
    layer2_outputs(10191) <= (layer1_outputs(9480)) and not (layer1_outputs(10292));
    layer2_outputs(10192) <= not(layer1_outputs(2728));
    layer2_outputs(10193) <= (layer1_outputs(12610)) or (layer1_outputs(12748));
    layer2_outputs(10194) <= not(layer1_outputs(5425));
    layer2_outputs(10195) <= layer1_outputs(1096);
    layer2_outputs(10196) <= (layer1_outputs(8324)) xor (layer1_outputs(4452));
    layer2_outputs(10197) <= layer1_outputs(9570);
    layer2_outputs(10198) <= (layer1_outputs(1517)) or (layer1_outputs(200));
    layer2_outputs(10199) <= layer1_outputs(10311);
    layer2_outputs(10200) <= not((layer1_outputs(7384)) xor (layer1_outputs(10307)));
    layer2_outputs(10201) <= not(layer1_outputs(4085));
    layer2_outputs(10202) <= layer1_outputs(5509);
    layer2_outputs(10203) <= layer1_outputs(8714);
    layer2_outputs(10204) <= (layer1_outputs(12163)) and not (layer1_outputs(5771));
    layer2_outputs(10205) <= not((layer1_outputs(10084)) or (layer1_outputs(11746)));
    layer2_outputs(10206) <= not(layer1_outputs(7000));
    layer2_outputs(10207) <= (layer1_outputs(5966)) xor (layer1_outputs(12151));
    layer2_outputs(10208) <= not(layer1_outputs(1707)) or (layer1_outputs(5513));
    layer2_outputs(10209) <= not(layer1_outputs(7578)) or (layer1_outputs(10501));
    layer2_outputs(10210) <= not(layer1_outputs(5252));
    layer2_outputs(10211) <= not((layer1_outputs(8758)) xor (layer1_outputs(9526)));
    layer2_outputs(10212) <= layer1_outputs(10923);
    layer2_outputs(10213) <= not(layer1_outputs(121));
    layer2_outputs(10214) <= layer1_outputs(4467);
    layer2_outputs(10215) <= not(layer1_outputs(8898)) or (layer1_outputs(4892));
    layer2_outputs(10216) <= not(layer1_outputs(3155));
    layer2_outputs(10217) <= (layer1_outputs(8151)) or (layer1_outputs(3190));
    layer2_outputs(10218) <= not(layer1_outputs(10208)) or (layer1_outputs(9087));
    layer2_outputs(10219) <= not(layer1_outputs(2937));
    layer2_outputs(10220) <= not(layer1_outputs(7989));
    layer2_outputs(10221) <= (layer1_outputs(10232)) xor (layer1_outputs(1395));
    layer2_outputs(10222) <= layer1_outputs(8269);
    layer2_outputs(10223) <= (layer1_outputs(7259)) and (layer1_outputs(2494));
    layer2_outputs(10224) <= not(layer1_outputs(9335));
    layer2_outputs(10225) <= (layer1_outputs(2441)) and not (layer1_outputs(2161));
    layer2_outputs(10226) <= not((layer1_outputs(567)) and (layer1_outputs(6474)));
    layer2_outputs(10227) <= not(layer1_outputs(1899));
    layer2_outputs(10228) <= layer1_outputs(7529);
    layer2_outputs(10229) <= not(layer1_outputs(2391));
    layer2_outputs(10230) <= not((layer1_outputs(6837)) and (layer1_outputs(411)));
    layer2_outputs(10231) <= layer1_outputs(9114);
    layer2_outputs(10232) <= not(layer1_outputs(10150)) or (layer1_outputs(7335));
    layer2_outputs(10233) <= not(layer1_outputs(12597));
    layer2_outputs(10234) <= layer1_outputs(8626);
    layer2_outputs(10235) <= layer1_outputs(4124);
    layer2_outputs(10236) <= not((layer1_outputs(6873)) xor (layer1_outputs(2173)));
    layer2_outputs(10237) <= not(layer1_outputs(4875)) or (layer1_outputs(8719));
    layer2_outputs(10238) <= (layer1_outputs(12268)) and (layer1_outputs(510));
    layer2_outputs(10239) <= (layer1_outputs(9450)) and not (layer1_outputs(7498));
    layer2_outputs(10240) <= not((layer1_outputs(5857)) and (layer1_outputs(6140)));
    layer2_outputs(10241) <= not(layer1_outputs(10203));
    layer2_outputs(10242) <= layer1_outputs(12449);
    layer2_outputs(10243) <= layer1_outputs(6328);
    layer2_outputs(10244) <= (layer1_outputs(12149)) xor (layer1_outputs(7013));
    layer2_outputs(10245) <= not(layer1_outputs(6656)) or (layer1_outputs(8836));
    layer2_outputs(10246) <= not((layer1_outputs(12380)) xor (layer1_outputs(7074)));
    layer2_outputs(10247) <= not(layer1_outputs(3261));
    layer2_outputs(10248) <= (layer1_outputs(12309)) and not (layer1_outputs(10873));
    layer2_outputs(10249) <= (layer1_outputs(3167)) and (layer1_outputs(2477));
    layer2_outputs(10250) <= not(layer1_outputs(2028)) or (layer1_outputs(12109));
    layer2_outputs(10251) <= layer1_outputs(11439);
    layer2_outputs(10252) <= (layer1_outputs(9388)) and not (layer1_outputs(11977));
    layer2_outputs(10253) <= not((layer1_outputs(1213)) and (layer1_outputs(9171)));
    layer2_outputs(10254) <= not((layer1_outputs(12337)) or (layer1_outputs(10800)));
    layer2_outputs(10255) <= layer1_outputs(9269);
    layer2_outputs(10256) <= not(layer1_outputs(2644));
    layer2_outputs(10257) <= layer1_outputs(9030);
    layer2_outputs(10258) <= layer1_outputs(4995);
    layer2_outputs(10259) <= (layer1_outputs(9410)) and not (layer1_outputs(4869));
    layer2_outputs(10260) <= not((layer1_outputs(2090)) and (layer1_outputs(7636)));
    layer2_outputs(10261) <= not((layer1_outputs(8636)) xor (layer1_outputs(7380)));
    layer2_outputs(10262) <= not((layer1_outputs(7840)) or (layer1_outputs(5493)));
    layer2_outputs(10263) <= not((layer1_outputs(12408)) or (layer1_outputs(227)));
    layer2_outputs(10264) <= (layer1_outputs(10452)) xor (layer1_outputs(6227));
    layer2_outputs(10265) <= not(layer1_outputs(3097)) or (layer1_outputs(3797));
    layer2_outputs(10266) <= not(layer1_outputs(8692)) or (layer1_outputs(10259));
    layer2_outputs(10267) <= not((layer1_outputs(10501)) or (layer1_outputs(5368)));
    layer2_outputs(10268) <= not((layer1_outputs(10125)) and (layer1_outputs(9399)));
    layer2_outputs(10269) <= (layer1_outputs(7662)) or (layer1_outputs(7316));
    layer2_outputs(10270) <= layer1_outputs(10226);
    layer2_outputs(10271) <= layer1_outputs(6567);
    layer2_outputs(10272) <= layer1_outputs(10470);
    layer2_outputs(10273) <= (layer1_outputs(8961)) or (layer1_outputs(7879));
    layer2_outputs(10274) <= (layer1_outputs(3829)) and (layer1_outputs(3839));
    layer2_outputs(10275) <= layer1_outputs(11931);
    layer2_outputs(10276) <= (layer1_outputs(3482)) or (layer1_outputs(9137));
    layer2_outputs(10277) <= not(layer1_outputs(3939));
    layer2_outputs(10278) <= not(layer1_outputs(3596)) or (layer1_outputs(11654));
    layer2_outputs(10279) <= (layer1_outputs(3133)) and (layer1_outputs(10206));
    layer2_outputs(10280) <= layer1_outputs(2591);
    layer2_outputs(10281) <= not(layer1_outputs(1416));
    layer2_outputs(10282) <= layer1_outputs(7548);
    layer2_outputs(10283) <= layer1_outputs(2412);
    layer2_outputs(10284) <= not((layer1_outputs(268)) xor (layer1_outputs(6800)));
    layer2_outputs(10285) <= not((layer1_outputs(7519)) or (layer1_outputs(1450)));
    layer2_outputs(10286) <= layer1_outputs(11125);
    layer2_outputs(10287) <= (layer1_outputs(11571)) and (layer1_outputs(8020));
    layer2_outputs(10288) <= not((layer1_outputs(8897)) xor (layer1_outputs(2693)));
    layer2_outputs(10289) <= not(layer1_outputs(5811));
    layer2_outputs(10290) <= not(layer1_outputs(8965));
    layer2_outputs(10291) <= not(layer1_outputs(11476));
    layer2_outputs(10292) <= layer1_outputs(4285);
    layer2_outputs(10293) <= not(layer1_outputs(2904));
    layer2_outputs(10294) <= not(layer1_outputs(9712));
    layer2_outputs(10295) <= (layer1_outputs(1347)) and (layer1_outputs(12));
    layer2_outputs(10296) <= (layer1_outputs(256)) or (layer1_outputs(6338));
    layer2_outputs(10297) <= (layer1_outputs(5584)) or (layer1_outputs(3974));
    layer2_outputs(10298) <= not(layer1_outputs(2595));
    layer2_outputs(10299) <= (layer1_outputs(2151)) xor (layer1_outputs(6350));
    layer2_outputs(10300) <= not((layer1_outputs(9619)) xor (layer1_outputs(8466)));
    layer2_outputs(10301) <= layer1_outputs(11556);
    layer2_outputs(10302) <= not(layer1_outputs(579));
    layer2_outputs(10303) <= layer1_outputs(6429);
    layer2_outputs(10304) <= (layer1_outputs(8750)) and (layer1_outputs(2588));
    layer2_outputs(10305) <= not(layer1_outputs(499)) or (layer1_outputs(3156));
    layer2_outputs(10306) <= layer1_outputs(6280);
    layer2_outputs(10307) <= (layer1_outputs(6680)) and (layer1_outputs(6011));
    layer2_outputs(10308) <= (layer1_outputs(9676)) xor (layer1_outputs(5394));
    layer2_outputs(10309) <= (layer1_outputs(5502)) or (layer1_outputs(262));
    layer2_outputs(10310) <= (layer1_outputs(11034)) and (layer1_outputs(3362));
    layer2_outputs(10311) <= not(layer1_outputs(6155)) or (layer1_outputs(5821));
    layer2_outputs(10312) <= not(layer1_outputs(11049));
    layer2_outputs(10313) <= (layer1_outputs(7129)) and not (layer1_outputs(3651));
    layer2_outputs(10314) <= not(layer1_outputs(2104));
    layer2_outputs(10315) <= not(layer1_outputs(5386)) or (layer1_outputs(4523));
    layer2_outputs(10316) <= (layer1_outputs(11334)) and not (layer1_outputs(4967));
    layer2_outputs(10317) <= layer1_outputs(511);
    layer2_outputs(10318) <= not((layer1_outputs(11131)) or (layer1_outputs(8835)));
    layer2_outputs(10319) <= layer1_outputs(2109);
    layer2_outputs(10320) <= layer1_outputs(6578);
    layer2_outputs(10321) <= not(layer1_outputs(11563));
    layer2_outputs(10322) <= layer1_outputs(4741);
    layer2_outputs(10323) <= layer1_outputs(9634);
    layer2_outputs(10324) <= not(layer1_outputs(1156));
    layer2_outputs(10325) <= (layer1_outputs(8414)) and (layer1_outputs(7713));
    layer2_outputs(10326) <= layer1_outputs(2085);
    layer2_outputs(10327) <= layer1_outputs(10583);
    layer2_outputs(10328) <= not((layer1_outputs(6292)) and (layer1_outputs(11871)));
    layer2_outputs(10329) <= not(layer1_outputs(1827)) or (layer1_outputs(1808));
    layer2_outputs(10330) <= layer1_outputs(10977);
    layer2_outputs(10331) <= not(layer1_outputs(6960));
    layer2_outputs(10332) <= layer1_outputs(5004);
    layer2_outputs(10333) <= not(layer1_outputs(5125));
    layer2_outputs(10334) <= not((layer1_outputs(6982)) and (layer1_outputs(3259)));
    layer2_outputs(10335) <= not(layer1_outputs(7391));
    layer2_outputs(10336) <= not(layer1_outputs(9571));
    layer2_outputs(10337) <= (layer1_outputs(10720)) and (layer1_outputs(8513));
    layer2_outputs(10338) <= not(layer1_outputs(9740));
    layer2_outputs(10339) <= (layer1_outputs(5938)) and not (layer1_outputs(1407));
    layer2_outputs(10340) <= not(layer1_outputs(10862));
    layer2_outputs(10341) <= layer1_outputs(10054);
    layer2_outputs(10342) <= not(layer1_outputs(6304)) or (layer1_outputs(12091));
    layer2_outputs(10343) <= not(layer1_outputs(1083)) or (layer1_outputs(9461));
    layer2_outputs(10344) <= not((layer1_outputs(3411)) or (layer1_outputs(6163)));
    layer2_outputs(10345) <= layer1_outputs(3526);
    layer2_outputs(10346) <= not(layer1_outputs(6787));
    layer2_outputs(10347) <= not((layer1_outputs(3426)) or (layer1_outputs(540)));
    layer2_outputs(10348) <= not((layer1_outputs(11678)) and (layer1_outputs(8797)));
    layer2_outputs(10349) <= not(layer1_outputs(4607)) or (layer1_outputs(8951));
    layer2_outputs(10350) <= (layer1_outputs(2897)) and not (layer1_outputs(5138));
    layer2_outputs(10351) <= (layer1_outputs(2278)) xor (layer1_outputs(5613));
    layer2_outputs(10352) <= not(layer1_outputs(6005));
    layer2_outputs(10353) <= layer1_outputs(10599);
    layer2_outputs(10354) <= not(layer1_outputs(11685)) or (layer1_outputs(1240));
    layer2_outputs(10355) <= layer1_outputs(10056);
    layer2_outputs(10356) <= layer1_outputs(11845);
    layer2_outputs(10357) <= not(layer1_outputs(7370));
    layer2_outputs(10358) <= layer1_outputs(9046);
    layer2_outputs(10359) <= not(layer1_outputs(9307));
    layer2_outputs(10360) <= not(layer1_outputs(8545));
    layer2_outputs(10361) <= layer1_outputs(8563);
    layer2_outputs(10362) <= not((layer1_outputs(3108)) xor (layer1_outputs(12780)));
    layer2_outputs(10363) <= not(layer1_outputs(3516)) or (layer1_outputs(7292));
    layer2_outputs(10364) <= not(layer1_outputs(2224));
    layer2_outputs(10365) <= not(layer1_outputs(10966));
    layer2_outputs(10366) <= layer1_outputs(11242);
    layer2_outputs(10367) <= layer1_outputs(3424);
    layer2_outputs(10368) <= not(layer1_outputs(11166));
    layer2_outputs(10369) <= not((layer1_outputs(1556)) xor (layer1_outputs(10888)));
    layer2_outputs(10370) <= (layer1_outputs(9473)) xor (layer1_outputs(10972));
    layer2_outputs(10371) <= (layer1_outputs(11502)) and not (layer1_outputs(5079));
    layer2_outputs(10372) <= layer1_outputs(10417);
    layer2_outputs(10373) <= not(layer1_outputs(8953));
    layer2_outputs(10374) <= (layer1_outputs(4546)) and not (layer1_outputs(1775));
    layer2_outputs(10375) <= not((layer1_outputs(11183)) and (layer1_outputs(1779)));
    layer2_outputs(10376) <= (layer1_outputs(11211)) and not (layer1_outputs(9313));
    layer2_outputs(10377) <= (layer1_outputs(6598)) and not (layer1_outputs(5571));
    layer2_outputs(10378) <= (layer1_outputs(1504)) and not (layer1_outputs(12332));
    layer2_outputs(10379) <= layer1_outputs(3244);
    layer2_outputs(10380) <= layer1_outputs(9275);
    layer2_outputs(10381) <= (layer1_outputs(3328)) xor (layer1_outputs(2475));
    layer2_outputs(10382) <= layer1_outputs(1547);
    layer2_outputs(10383) <= not(layer1_outputs(7571));
    layer2_outputs(10384) <= not(layer1_outputs(12701));
    layer2_outputs(10385) <= '0';
    layer2_outputs(10386) <= not((layer1_outputs(4200)) xor (layer1_outputs(6090)));
    layer2_outputs(10387) <= not((layer1_outputs(3116)) and (layer1_outputs(3424)));
    layer2_outputs(10388) <= layer1_outputs(9816);
    layer2_outputs(10389) <= (layer1_outputs(4350)) and not (layer1_outputs(5120));
    layer2_outputs(10390) <= not(layer1_outputs(9616));
    layer2_outputs(10391) <= not((layer1_outputs(1132)) or (layer1_outputs(1047)));
    layer2_outputs(10392) <= not(layer1_outputs(2032));
    layer2_outputs(10393) <= not(layer1_outputs(443));
    layer2_outputs(10394) <= not((layer1_outputs(5020)) and (layer1_outputs(11671)));
    layer2_outputs(10395) <= layer1_outputs(10226);
    layer2_outputs(10396) <= (layer1_outputs(6565)) or (layer1_outputs(1711));
    layer2_outputs(10397) <= not(layer1_outputs(5815));
    layer2_outputs(10398) <= layer1_outputs(12402);
    layer2_outputs(10399) <= not(layer1_outputs(1278));
    layer2_outputs(10400) <= not(layer1_outputs(2539));
    layer2_outputs(10401) <= not(layer1_outputs(6993));
    layer2_outputs(10402) <= not(layer1_outputs(2896));
    layer2_outputs(10403) <= (layer1_outputs(8879)) and not (layer1_outputs(6146));
    layer2_outputs(10404) <= (layer1_outputs(6779)) and not (layer1_outputs(11401));
    layer2_outputs(10405) <= not(layer1_outputs(1046));
    layer2_outputs(10406) <= not(layer1_outputs(1887));
    layer2_outputs(10407) <= not(layer1_outputs(6822)) or (layer1_outputs(11734));
    layer2_outputs(10408) <= not(layer1_outputs(12223));
    layer2_outputs(10409) <= not(layer1_outputs(5508));
    layer2_outputs(10410) <= not((layer1_outputs(254)) and (layer1_outputs(1099)));
    layer2_outputs(10411) <= (layer1_outputs(12545)) and (layer1_outputs(4729));
    layer2_outputs(10412) <= not((layer1_outputs(521)) and (layer1_outputs(6318)));
    layer2_outputs(10413) <= not(layer1_outputs(5955));
    layer2_outputs(10414) <= layer1_outputs(4168);
    layer2_outputs(10415) <= not((layer1_outputs(7574)) xor (layer1_outputs(1129)));
    layer2_outputs(10416) <= not(layer1_outputs(9812));
    layer2_outputs(10417) <= not((layer1_outputs(10585)) xor (layer1_outputs(5550)));
    layer2_outputs(10418) <= not(layer1_outputs(446));
    layer2_outputs(10419) <= (layer1_outputs(2942)) xor (layer1_outputs(11450));
    layer2_outputs(10420) <= layer1_outputs(5734);
    layer2_outputs(10421) <= layer1_outputs(2325);
    layer2_outputs(10422) <= (layer1_outputs(10355)) and not (layer1_outputs(12234));
    layer2_outputs(10423) <= not(layer1_outputs(2431)) or (layer1_outputs(3677));
    layer2_outputs(10424) <= not(layer1_outputs(2895));
    layer2_outputs(10425) <= layer1_outputs(4849);
    layer2_outputs(10426) <= (layer1_outputs(1861)) and not (layer1_outputs(4656));
    layer2_outputs(10427) <= (layer1_outputs(11310)) xor (layer1_outputs(9850));
    layer2_outputs(10428) <= not(layer1_outputs(12362));
    layer2_outputs(10429) <= layer1_outputs(10485);
    layer2_outputs(10430) <= layer1_outputs(8811);
    layer2_outputs(10431) <= (layer1_outputs(11898)) or (layer1_outputs(5195));
    layer2_outputs(10432) <= not((layer1_outputs(9903)) and (layer1_outputs(430)));
    layer2_outputs(10433) <= not((layer1_outputs(6328)) or (layer1_outputs(6844)));
    layer2_outputs(10434) <= (layer1_outputs(7408)) and (layer1_outputs(7920));
    layer2_outputs(10435) <= layer1_outputs(3149);
    layer2_outputs(10436) <= (layer1_outputs(5922)) or (layer1_outputs(10752));
    layer2_outputs(10437) <= (layer1_outputs(12605)) or (layer1_outputs(11381));
    layer2_outputs(10438) <= (layer1_outputs(5928)) and not (layer1_outputs(8529));
    layer2_outputs(10439) <= (layer1_outputs(7720)) and (layer1_outputs(4921));
    layer2_outputs(10440) <= (layer1_outputs(7626)) and not (layer1_outputs(12189));
    layer2_outputs(10441) <= layer1_outputs(1102);
    layer2_outputs(10442) <= layer1_outputs(11644);
    layer2_outputs(10443) <= (layer1_outputs(1844)) xor (layer1_outputs(9653));
    layer2_outputs(10444) <= layer1_outputs(8719);
    layer2_outputs(10445) <= layer1_outputs(6572);
    layer2_outputs(10446) <= not((layer1_outputs(10737)) or (layer1_outputs(1763)));
    layer2_outputs(10447) <= layer1_outputs(857);
    layer2_outputs(10448) <= layer1_outputs(12554);
    layer2_outputs(10449) <= not((layer1_outputs(4594)) or (layer1_outputs(8392)));
    layer2_outputs(10450) <= not((layer1_outputs(2360)) or (layer1_outputs(10681)));
    layer2_outputs(10451) <= not(layer1_outputs(11689)) or (layer1_outputs(11899));
    layer2_outputs(10452) <= layer1_outputs(9074);
    layer2_outputs(10453) <= not(layer1_outputs(3401));
    layer2_outputs(10454) <= layer1_outputs(12404);
    layer2_outputs(10455) <= (layer1_outputs(12183)) or (layer1_outputs(10625));
    layer2_outputs(10456) <= not(layer1_outputs(2864));
    layer2_outputs(10457) <= not(layer1_outputs(2120));
    layer2_outputs(10458) <= not(layer1_outputs(3572));
    layer2_outputs(10459) <= not(layer1_outputs(1719));
    layer2_outputs(10460) <= not((layer1_outputs(9923)) or (layer1_outputs(5243)));
    layer2_outputs(10461) <= not((layer1_outputs(1222)) or (layer1_outputs(6073)));
    layer2_outputs(10462) <= layer1_outputs(7443);
    layer2_outputs(10463) <= not((layer1_outputs(4111)) or (layer1_outputs(1906)));
    layer2_outputs(10464) <= layer1_outputs(10690);
    layer2_outputs(10465) <= layer1_outputs(1068);
    layer2_outputs(10466) <= not(layer1_outputs(3421));
    layer2_outputs(10467) <= layer1_outputs(3616);
    layer2_outputs(10468) <= not(layer1_outputs(9766));
    layer2_outputs(10469) <= not(layer1_outputs(5547));
    layer2_outputs(10470) <= '0';
    layer2_outputs(10471) <= (layer1_outputs(10420)) and not (layer1_outputs(7762));
    layer2_outputs(10472) <= not((layer1_outputs(9235)) or (layer1_outputs(811)));
    layer2_outputs(10473) <= not((layer1_outputs(9589)) or (layer1_outputs(4138)));
    layer2_outputs(10474) <= (layer1_outputs(7452)) or (layer1_outputs(664));
    layer2_outputs(10475) <= not((layer1_outputs(11858)) or (layer1_outputs(9602)));
    layer2_outputs(10476) <= not(layer1_outputs(233));
    layer2_outputs(10477) <= layer1_outputs(4956);
    layer2_outputs(10478) <= not((layer1_outputs(1877)) xor (layer1_outputs(3753)));
    layer2_outputs(10479) <= layer1_outputs(4044);
    layer2_outputs(10480) <= not(layer1_outputs(12659)) or (layer1_outputs(6762));
    layer2_outputs(10481) <= not(layer1_outputs(1877));
    layer2_outputs(10482) <= (layer1_outputs(10011)) and not (layer1_outputs(5081));
    layer2_outputs(10483) <= layer1_outputs(1434);
    layer2_outputs(10484) <= not((layer1_outputs(5778)) and (layer1_outputs(10983)));
    layer2_outputs(10485) <= not(layer1_outputs(741));
    layer2_outputs(10486) <= not(layer1_outputs(9710)) or (layer1_outputs(928));
    layer2_outputs(10487) <= layer1_outputs(7914);
    layer2_outputs(10488) <= layer1_outputs(11191);
    layer2_outputs(10489) <= layer1_outputs(8937);
    layer2_outputs(10490) <= not((layer1_outputs(4029)) or (layer1_outputs(6718)));
    layer2_outputs(10491) <= (layer1_outputs(1926)) and not (layer1_outputs(6590));
    layer2_outputs(10492) <= not(layer1_outputs(1666));
    layer2_outputs(10493) <= layer1_outputs(12608);
    layer2_outputs(10494) <= not(layer1_outputs(1615));
    layer2_outputs(10495) <= (layer1_outputs(9325)) xor (layer1_outputs(8010));
    layer2_outputs(10496) <= layer1_outputs(4092);
    layer2_outputs(10497) <= (layer1_outputs(12360)) xor (layer1_outputs(2392));
    layer2_outputs(10498) <= layer1_outputs(4210);
    layer2_outputs(10499) <= layer1_outputs(769);
    layer2_outputs(10500) <= not((layer1_outputs(1100)) xor (layer1_outputs(3964)));
    layer2_outputs(10501) <= layer1_outputs(4761);
    layer2_outputs(10502) <= '1';
    layer2_outputs(10503) <= not(layer1_outputs(11023)) or (layer1_outputs(10135));
    layer2_outputs(10504) <= not((layer1_outputs(677)) and (layer1_outputs(7996)));
    layer2_outputs(10505) <= layer1_outputs(12308);
    layer2_outputs(10506) <= layer1_outputs(11695);
    layer2_outputs(10507) <= (layer1_outputs(3383)) xor (layer1_outputs(10485));
    layer2_outputs(10508) <= (layer1_outputs(6280)) or (layer1_outputs(5507));
    layer2_outputs(10509) <= layer1_outputs(10046);
    layer2_outputs(10510) <= (layer1_outputs(3940)) and not (layer1_outputs(11378));
    layer2_outputs(10511) <= not(layer1_outputs(8958));
    layer2_outputs(10512) <= (layer1_outputs(71)) or (layer1_outputs(7920));
    layer2_outputs(10513) <= layer1_outputs(9249);
    layer2_outputs(10514) <= not(layer1_outputs(948));
    layer2_outputs(10515) <= layer1_outputs(11183);
    layer2_outputs(10516) <= (layer1_outputs(9097)) xor (layer1_outputs(3474));
    layer2_outputs(10517) <= layer1_outputs(4946);
    layer2_outputs(10518) <= not(layer1_outputs(63));
    layer2_outputs(10519) <= (layer1_outputs(11910)) and not (layer1_outputs(10913));
    layer2_outputs(10520) <= not((layer1_outputs(12798)) and (layer1_outputs(1850)));
    layer2_outputs(10521) <= not(layer1_outputs(203));
    layer2_outputs(10522) <= not(layer1_outputs(11952));
    layer2_outputs(10523) <= layer1_outputs(7374);
    layer2_outputs(10524) <= layer1_outputs(8900);
    layer2_outputs(10525) <= not((layer1_outputs(2145)) xor (layer1_outputs(9304)));
    layer2_outputs(10526) <= layer1_outputs(5537);
    layer2_outputs(10527) <= not((layer1_outputs(1171)) or (layer1_outputs(8370)));
    layer2_outputs(10528) <= not((layer1_outputs(8294)) xor (layer1_outputs(974)));
    layer2_outputs(10529) <= not(layer1_outputs(7672));
    layer2_outputs(10530) <= not(layer1_outputs(6649));
    layer2_outputs(10531) <= layer1_outputs(9500);
    layer2_outputs(10532) <= not((layer1_outputs(4625)) and (layer1_outputs(7911)));
    layer2_outputs(10533) <= (layer1_outputs(5065)) or (layer1_outputs(4587));
    layer2_outputs(10534) <= not(layer1_outputs(5848));
    layer2_outputs(10535) <= not(layer1_outputs(8638)) or (layer1_outputs(12195));
    layer2_outputs(10536) <= layer1_outputs(5817);
    layer2_outputs(10537) <= not(layer1_outputs(7283)) or (layer1_outputs(2622));
    layer2_outputs(10538) <= (layer1_outputs(9120)) and not (layer1_outputs(3714));
    layer2_outputs(10539) <= (layer1_outputs(5114)) and not (layer1_outputs(5521));
    layer2_outputs(10540) <= layer1_outputs(11801);
    layer2_outputs(10541) <= not(layer1_outputs(7881));
    layer2_outputs(10542) <= (layer1_outputs(6434)) or (layer1_outputs(10409));
    layer2_outputs(10543) <= (layer1_outputs(10115)) and (layer1_outputs(3507));
    layer2_outputs(10544) <= not(layer1_outputs(11171));
    layer2_outputs(10545) <= layer1_outputs(11292);
    layer2_outputs(10546) <= (layer1_outputs(4263)) and not (layer1_outputs(5308));
    layer2_outputs(10547) <= (layer1_outputs(10013)) and (layer1_outputs(4046));
    layer2_outputs(10548) <= not((layer1_outputs(1550)) xor (layer1_outputs(11255)));
    layer2_outputs(10549) <= not((layer1_outputs(4119)) xor (layer1_outputs(7394)));
    layer2_outputs(10550) <= (layer1_outputs(11899)) xor (layer1_outputs(406));
    layer2_outputs(10551) <= layer1_outputs(1237);
    layer2_outputs(10552) <= not(layer1_outputs(3128));
    layer2_outputs(10553) <= not(layer1_outputs(10778));
    layer2_outputs(10554) <= layer1_outputs(560);
    layer2_outputs(10555) <= not((layer1_outputs(7963)) xor (layer1_outputs(6030)));
    layer2_outputs(10556) <= layer1_outputs(12353);
    layer2_outputs(10557) <= layer1_outputs(5207);
    layer2_outputs(10558) <= not((layer1_outputs(4732)) or (layer1_outputs(12059)));
    layer2_outputs(10559) <= not(layer1_outputs(3663));
    layer2_outputs(10560) <= not(layer1_outputs(10120));
    layer2_outputs(10561) <= not(layer1_outputs(7778));
    layer2_outputs(10562) <= (layer1_outputs(2121)) and not (layer1_outputs(10183));
    layer2_outputs(10563) <= (layer1_outputs(5767)) and not (layer1_outputs(238));
    layer2_outputs(10564) <= layer1_outputs(2288);
    layer2_outputs(10565) <= not(layer1_outputs(2906));
    layer2_outputs(10566) <= not(layer1_outputs(1328));
    layer2_outputs(10567) <= layer1_outputs(2022);
    layer2_outputs(10568) <= not(layer1_outputs(590));
    layer2_outputs(10569) <= layer1_outputs(563);
    layer2_outputs(10570) <= not((layer1_outputs(10421)) or (layer1_outputs(9874)));
    layer2_outputs(10571) <= not((layer1_outputs(6050)) and (layer1_outputs(2243)));
    layer2_outputs(10572) <= not((layer1_outputs(6540)) xor (layer1_outputs(12453)));
    layer2_outputs(10573) <= not((layer1_outputs(3346)) or (layer1_outputs(4463)));
    layer2_outputs(10574) <= not(layer1_outputs(1917));
    layer2_outputs(10575) <= (layer1_outputs(5100)) or (layer1_outputs(6700));
    layer2_outputs(10576) <= layer1_outputs(1896);
    layer2_outputs(10577) <= (layer1_outputs(3373)) and not (layer1_outputs(5185));
    layer2_outputs(10578) <= (layer1_outputs(8854)) and not (layer1_outputs(7341));
    layer2_outputs(10579) <= not(layer1_outputs(9180));
    layer2_outputs(10580) <= (layer1_outputs(3035)) or (layer1_outputs(1414));
    layer2_outputs(10581) <= not(layer1_outputs(5483));
    layer2_outputs(10582) <= (layer1_outputs(4876)) or (layer1_outputs(3660));
    layer2_outputs(10583) <= '0';
    layer2_outputs(10584) <= (layer1_outputs(2339)) and (layer1_outputs(11279));
    layer2_outputs(10585) <= not((layer1_outputs(6080)) or (layer1_outputs(9224)));
    layer2_outputs(10586) <= not((layer1_outputs(4722)) and (layer1_outputs(7275)));
    layer2_outputs(10587) <= (layer1_outputs(5330)) and (layer1_outputs(1726));
    layer2_outputs(10588) <= (layer1_outputs(1008)) xor (layer1_outputs(2727));
    layer2_outputs(10589) <= layer1_outputs(12499);
    layer2_outputs(10590) <= layer1_outputs(1614);
    layer2_outputs(10591) <= not(layer1_outputs(12694)) or (layer1_outputs(5946));
    layer2_outputs(10592) <= layer1_outputs(2517);
    layer2_outputs(10593) <= layer1_outputs(7709);
    layer2_outputs(10594) <= layer1_outputs(10967);
    layer2_outputs(10595) <= not((layer1_outputs(7962)) xor (layer1_outputs(12756)));
    layer2_outputs(10596) <= not(layer1_outputs(12606));
    layer2_outputs(10597) <= (layer1_outputs(6492)) and (layer1_outputs(475));
    layer2_outputs(10598) <= not(layer1_outputs(7516));
    layer2_outputs(10599) <= layer1_outputs(6575);
    layer2_outputs(10600) <= layer1_outputs(8309);
    layer2_outputs(10601) <= layer1_outputs(6364);
    layer2_outputs(10602) <= (layer1_outputs(3312)) and not (layer1_outputs(4779));
    layer2_outputs(10603) <= not(layer1_outputs(2364));
    layer2_outputs(10604) <= (layer1_outputs(808)) and not (layer1_outputs(2639));
    layer2_outputs(10605) <= (layer1_outputs(10249)) or (layer1_outputs(5505));
    layer2_outputs(10606) <= layer1_outputs(1820);
    layer2_outputs(10607) <= not(layer1_outputs(8644));
    layer2_outputs(10608) <= (layer1_outputs(1891)) and not (layer1_outputs(12577));
    layer2_outputs(10609) <= not(layer1_outputs(746));
    layer2_outputs(10610) <= (layer1_outputs(12769)) and not (layer1_outputs(6266));
    layer2_outputs(10611) <= layer1_outputs(2965);
    layer2_outputs(10612) <= layer1_outputs(9644);
    layer2_outputs(10613) <= not((layer1_outputs(7662)) and (layer1_outputs(6334)));
    layer2_outputs(10614) <= layer1_outputs(5239);
    layer2_outputs(10615) <= (layer1_outputs(7666)) xor (layer1_outputs(12751));
    layer2_outputs(10616) <= not(layer1_outputs(10847)) or (layer1_outputs(5016));
    layer2_outputs(10617) <= not(layer1_outputs(2760));
    layer2_outputs(10618) <= not((layer1_outputs(3150)) xor (layer1_outputs(302)));
    layer2_outputs(10619) <= (layer1_outputs(4274)) and not (layer1_outputs(3927));
    layer2_outputs(10620) <= not(layer1_outputs(12283));
    layer2_outputs(10621) <= not(layer1_outputs(11660));
    layer2_outputs(10622) <= (layer1_outputs(5437)) and not (layer1_outputs(11624));
    layer2_outputs(10623) <= layer1_outputs(1702);
    layer2_outputs(10624) <= not(layer1_outputs(11425));
    layer2_outputs(10625) <= layer1_outputs(4454);
    layer2_outputs(10626) <= not(layer1_outputs(676));
    layer2_outputs(10627) <= not(layer1_outputs(600));
    layer2_outputs(10628) <= layer1_outputs(4797);
    layer2_outputs(10629) <= not(layer1_outputs(1115));
    layer2_outputs(10630) <= layer1_outputs(415);
    layer2_outputs(10631) <= (layer1_outputs(8404)) and not (layer1_outputs(9380));
    layer2_outputs(10632) <= (layer1_outputs(3693)) and (layer1_outputs(2721));
    layer2_outputs(10633) <= (layer1_outputs(8595)) xor (layer1_outputs(3436));
    layer2_outputs(10634) <= (layer1_outputs(7394)) xor (layer1_outputs(7683));
    layer2_outputs(10635) <= not(layer1_outputs(10080));
    layer2_outputs(10636) <= (layer1_outputs(7725)) xor (layer1_outputs(454));
    layer2_outputs(10637) <= not((layer1_outputs(11152)) or (layer1_outputs(11065)));
    layer2_outputs(10638) <= (layer1_outputs(9683)) or (layer1_outputs(1811));
    layer2_outputs(10639) <= layer1_outputs(12584);
    layer2_outputs(10640) <= (layer1_outputs(9087)) and (layer1_outputs(6091));
    layer2_outputs(10641) <= (layer1_outputs(8637)) xor (layer1_outputs(3969));
    layer2_outputs(10642) <= not((layer1_outputs(6063)) xor (layer1_outputs(8700)));
    layer2_outputs(10643) <= not(layer1_outputs(6731));
    layer2_outputs(10644) <= (layer1_outputs(6822)) xor (layer1_outputs(3892));
    layer2_outputs(10645) <= (layer1_outputs(7063)) xor (layer1_outputs(6897));
    layer2_outputs(10646) <= not(layer1_outputs(4041));
    layer2_outputs(10647) <= layer1_outputs(12737);
    layer2_outputs(10648) <= not(layer1_outputs(3402));
    layer2_outputs(10649) <= not(layer1_outputs(2728));
    layer2_outputs(10650) <= not(layer1_outputs(8183)) or (layer1_outputs(138));
    layer2_outputs(10651) <= not(layer1_outputs(6557));
    layer2_outputs(10652) <= (layer1_outputs(10149)) xor (layer1_outputs(2859));
    layer2_outputs(10653) <= (layer1_outputs(5557)) xor (layer1_outputs(8951));
    layer2_outputs(10654) <= (layer1_outputs(5798)) xor (layer1_outputs(8612));
    layer2_outputs(10655) <= (layer1_outputs(12358)) xor (layer1_outputs(1080));
    layer2_outputs(10656) <= not(layer1_outputs(6342)) or (layer1_outputs(944));
    layer2_outputs(10657) <= layer1_outputs(12316);
    layer2_outputs(10658) <= not((layer1_outputs(574)) xor (layer1_outputs(9568)));
    layer2_outputs(10659) <= not((layer1_outputs(6361)) and (layer1_outputs(5893)));
    layer2_outputs(10660) <= layer1_outputs(10368);
    layer2_outputs(10661) <= not(layer1_outputs(4164));
    layer2_outputs(10662) <= (layer1_outputs(4513)) and not (layer1_outputs(8541));
    layer2_outputs(10663) <= (layer1_outputs(2014)) and (layer1_outputs(4047));
    layer2_outputs(10664) <= (layer1_outputs(2225)) or (layer1_outputs(9646));
    layer2_outputs(10665) <= (layer1_outputs(11603)) xor (layer1_outputs(12608));
    layer2_outputs(10666) <= (layer1_outputs(11653)) xor (layer1_outputs(8170));
    layer2_outputs(10667) <= layer1_outputs(2608);
    layer2_outputs(10668) <= (layer1_outputs(10583)) xor (layer1_outputs(8102));
    layer2_outputs(10669) <= (layer1_outputs(10898)) and not (layer1_outputs(3592));
    layer2_outputs(10670) <= not(layer1_outputs(6454));
    layer2_outputs(10671) <= (layer1_outputs(10977)) and not (layer1_outputs(4524));
    layer2_outputs(10672) <= (layer1_outputs(10999)) and not (layer1_outputs(9140));
    layer2_outputs(10673) <= not(layer1_outputs(986));
    layer2_outputs(10674) <= layer1_outputs(3591);
    layer2_outputs(10675) <= not(layer1_outputs(1288));
    layer2_outputs(10676) <= not(layer1_outputs(7780));
    layer2_outputs(10677) <= not((layer1_outputs(11636)) and (layer1_outputs(3970)));
    layer2_outputs(10678) <= (layer1_outputs(5315)) or (layer1_outputs(4863));
    layer2_outputs(10679) <= (layer1_outputs(4737)) and (layer1_outputs(11607));
    layer2_outputs(10680) <= not((layer1_outputs(4540)) xor (layer1_outputs(7052)));
    layer2_outputs(10681) <= not((layer1_outputs(11961)) xor (layer1_outputs(11236)));
    layer2_outputs(10682) <= not((layer1_outputs(1034)) or (layer1_outputs(4856)));
    layer2_outputs(10683) <= not(layer1_outputs(3600));
    layer2_outputs(10684) <= not(layer1_outputs(1064));
    layer2_outputs(10685) <= not(layer1_outputs(6495));
    layer2_outputs(10686) <= not((layer1_outputs(9707)) and (layer1_outputs(10751)));
    layer2_outputs(10687) <= not((layer1_outputs(6499)) or (layer1_outputs(10139)));
    layer2_outputs(10688) <= not(layer1_outputs(6337));
    layer2_outputs(10689) <= layer1_outputs(9716);
    layer2_outputs(10690) <= not(layer1_outputs(9863));
    layer2_outputs(10691) <= (layer1_outputs(99)) and not (layer1_outputs(7400));
    layer2_outputs(10692) <= not((layer1_outputs(5276)) xor (layer1_outputs(11123)));
    layer2_outputs(10693) <= not(layer1_outputs(6953)) or (layer1_outputs(2735));
    layer2_outputs(10694) <= layer1_outputs(5691);
    layer2_outputs(10695) <= not(layer1_outputs(4725));
    layer2_outputs(10696) <= not(layer1_outputs(5687)) or (layer1_outputs(2507));
    layer2_outputs(10697) <= not((layer1_outputs(11866)) and (layer1_outputs(2284)));
    layer2_outputs(10698) <= not(layer1_outputs(9276)) or (layer1_outputs(10098));
    layer2_outputs(10699) <= not(layer1_outputs(2839));
    layer2_outputs(10700) <= not((layer1_outputs(5729)) xor (layer1_outputs(6225)));
    layer2_outputs(10701) <= not(layer1_outputs(12416));
    layer2_outputs(10702) <= layer1_outputs(8538);
    layer2_outputs(10703) <= layer1_outputs(6381);
    layer2_outputs(10704) <= not((layer1_outputs(4789)) or (layer1_outputs(8277)));
    layer2_outputs(10705) <= layer1_outputs(306);
    layer2_outputs(10706) <= not(layer1_outputs(10815));
    layer2_outputs(10707) <= (layer1_outputs(8618)) or (layer1_outputs(6213));
    layer2_outputs(10708) <= not((layer1_outputs(1574)) and (layer1_outputs(4777)));
    layer2_outputs(10709) <= not(layer1_outputs(5302));
    layer2_outputs(10710) <= not((layer1_outputs(1217)) and (layer1_outputs(2237)));
    layer2_outputs(10711) <= layer1_outputs(6856);
    layer2_outputs(10712) <= not((layer1_outputs(5845)) and (layer1_outputs(10676)));
    layer2_outputs(10713) <= layer1_outputs(12025);
    layer2_outputs(10714) <= (layer1_outputs(9337)) xor (layer1_outputs(9218));
    layer2_outputs(10715) <= not(layer1_outputs(705));
    layer2_outputs(10716) <= (layer1_outputs(7563)) or (layer1_outputs(5151));
    layer2_outputs(10717) <= layer1_outputs(8439);
    layer2_outputs(10718) <= not((layer1_outputs(7742)) xor (layer1_outputs(5555)));
    layer2_outputs(10719) <= '0';
    layer2_outputs(10720) <= not(layer1_outputs(5657));
    layer2_outputs(10721) <= layer1_outputs(6368);
    layer2_outputs(10722) <= not((layer1_outputs(3408)) xor (layer1_outputs(2189)));
    layer2_outputs(10723) <= not((layer1_outputs(11945)) or (layer1_outputs(401)));
    layer2_outputs(10724) <= not((layer1_outputs(500)) and (layer1_outputs(2562)));
    layer2_outputs(10725) <= not((layer1_outputs(3221)) xor (layer1_outputs(1711)));
    layer2_outputs(10726) <= (layer1_outputs(688)) and not (layer1_outputs(12710));
    layer2_outputs(10727) <= (layer1_outputs(4975)) and (layer1_outputs(5809));
    layer2_outputs(10728) <= layer1_outputs(2640);
    layer2_outputs(10729) <= not(layer1_outputs(10629));
    layer2_outputs(10730) <= not(layer1_outputs(4136)) or (layer1_outputs(12665));
    layer2_outputs(10731) <= not(layer1_outputs(286));
    layer2_outputs(10732) <= not(layer1_outputs(2509)) or (layer1_outputs(11359));
    layer2_outputs(10733) <= layer1_outputs(6606);
    layer2_outputs(10734) <= (layer1_outputs(5670)) xor (layer1_outputs(11863));
    layer2_outputs(10735) <= not(layer1_outputs(10071));
    layer2_outputs(10736) <= not((layer1_outputs(6102)) xor (layer1_outputs(9268)));
    layer2_outputs(10737) <= not(layer1_outputs(9057));
    layer2_outputs(10738) <= (layer1_outputs(1073)) and not (layer1_outputs(5395));
    layer2_outputs(10739) <= not((layer1_outputs(11224)) xor (layer1_outputs(4108)));
    layer2_outputs(10740) <= layer1_outputs(8646);
    layer2_outputs(10741) <= layer1_outputs(1568);
    layer2_outputs(10742) <= (layer1_outputs(5703)) xor (layer1_outputs(3416));
    layer2_outputs(10743) <= (layer1_outputs(1602)) and not (layer1_outputs(2973));
    layer2_outputs(10744) <= not((layer1_outputs(4375)) and (layer1_outputs(780)));
    layer2_outputs(10745) <= (layer1_outputs(9605)) xor (layer1_outputs(3962));
    layer2_outputs(10746) <= layer1_outputs(4048);
    layer2_outputs(10747) <= (layer1_outputs(8908)) and (layer1_outputs(1441));
    layer2_outputs(10748) <= layer1_outputs(12555);
    layer2_outputs(10749) <= layer1_outputs(6764);
    layer2_outputs(10750) <= not(layer1_outputs(12439));
    layer2_outputs(10751) <= not(layer1_outputs(8101));
    layer2_outputs(10752) <= layer1_outputs(5857);
    layer2_outputs(10753) <= not((layer1_outputs(9031)) and (layer1_outputs(7786)));
    layer2_outputs(10754) <= layer1_outputs(6851);
    layer2_outputs(10755) <= not(layer1_outputs(2630)) or (layer1_outputs(3379));
    layer2_outputs(10756) <= not(layer1_outputs(4418));
    layer2_outputs(10757) <= layer1_outputs(6496);
    layer2_outputs(10758) <= (layer1_outputs(1051)) and (layer1_outputs(8072));
    layer2_outputs(10759) <= layer1_outputs(4276);
    layer2_outputs(10760) <= not(layer1_outputs(8055));
    layer2_outputs(10761) <= not((layer1_outputs(11426)) and (layer1_outputs(9606)));
    layer2_outputs(10762) <= not(layer1_outputs(9299)) or (layer1_outputs(3631));
    layer2_outputs(10763) <= layer1_outputs(2894);
    layer2_outputs(10764) <= not(layer1_outputs(6003));
    layer2_outputs(10765) <= not(layer1_outputs(3849));
    layer2_outputs(10766) <= not(layer1_outputs(1789));
    layer2_outputs(10767) <= (layer1_outputs(1096)) and not (layer1_outputs(4031));
    layer2_outputs(10768) <= layer1_outputs(3931);
    layer2_outputs(10769) <= not(layer1_outputs(7078));
    layer2_outputs(10770) <= not(layer1_outputs(9592));
    layer2_outputs(10771) <= (layer1_outputs(9919)) and not (layer1_outputs(8185));
    layer2_outputs(10772) <= (layer1_outputs(6354)) or (layer1_outputs(9665));
    layer2_outputs(10773) <= not((layer1_outputs(7568)) xor (layer1_outputs(2114)));
    layer2_outputs(10774) <= not(layer1_outputs(5168));
    layer2_outputs(10775) <= (layer1_outputs(6030)) and (layer1_outputs(150));
    layer2_outputs(10776) <= layer1_outputs(1776);
    layer2_outputs(10777) <= layer1_outputs(5710);
    layer2_outputs(10778) <= layer1_outputs(9286);
    layer2_outputs(10779) <= layer1_outputs(2394);
    layer2_outputs(10780) <= not((layer1_outputs(7836)) and (layer1_outputs(9858)));
    layer2_outputs(10781) <= not(layer1_outputs(9687));
    layer2_outputs(10782) <= (layer1_outputs(10365)) or (layer1_outputs(1164));
    layer2_outputs(10783) <= not((layer1_outputs(924)) or (layer1_outputs(10272)));
    layer2_outputs(10784) <= layer1_outputs(3527);
    layer2_outputs(10785) <= not(layer1_outputs(506)) or (layer1_outputs(10534));
    layer2_outputs(10786) <= (layer1_outputs(9377)) and (layer1_outputs(9059));
    layer2_outputs(10787) <= (layer1_outputs(11510)) and not (layer1_outputs(8683));
    layer2_outputs(10788) <= not((layer1_outputs(12344)) xor (layer1_outputs(6685)));
    layer2_outputs(10789) <= layer1_outputs(1452);
    layer2_outputs(10790) <= layer1_outputs(8847);
    layer2_outputs(10791) <= not(layer1_outputs(7707)) or (layer1_outputs(5072));
    layer2_outputs(10792) <= layer1_outputs(785);
    layer2_outputs(10793) <= (layer1_outputs(9079)) and (layer1_outputs(9869));
    layer2_outputs(10794) <= (layer1_outputs(122)) or (layer1_outputs(12787));
    layer2_outputs(10795) <= not(layer1_outputs(4270)) or (layer1_outputs(5285));
    layer2_outputs(10796) <= not(layer1_outputs(1200));
    layer2_outputs(10797) <= not(layer1_outputs(12736)) or (layer1_outputs(12723));
    layer2_outputs(10798) <= not(layer1_outputs(3456));
    layer2_outputs(10799) <= not(layer1_outputs(3225));
    layer2_outputs(10800) <= not((layer1_outputs(10656)) xor (layer1_outputs(8729)));
    layer2_outputs(10801) <= not((layer1_outputs(3479)) or (layer1_outputs(2454)));
    layer2_outputs(10802) <= not((layer1_outputs(8672)) xor (layer1_outputs(966)));
    layer2_outputs(10803) <= (layer1_outputs(8678)) xor (layer1_outputs(7316));
    layer2_outputs(10804) <= not((layer1_outputs(2186)) and (layer1_outputs(4106)));
    layer2_outputs(10805) <= (layer1_outputs(3370)) xor (layer1_outputs(3251));
    layer2_outputs(10806) <= not(layer1_outputs(3253));
    layer2_outputs(10807) <= (layer1_outputs(7277)) xor (layer1_outputs(6451));
    layer2_outputs(10808) <= not(layer1_outputs(10003));
    layer2_outputs(10809) <= not(layer1_outputs(5031));
    layer2_outputs(10810) <= not((layer1_outputs(10194)) xor (layer1_outputs(12624)));
    layer2_outputs(10811) <= not(layer1_outputs(4638));
    layer2_outputs(10812) <= not((layer1_outputs(2887)) xor (layer1_outputs(3090)));
    layer2_outputs(10813) <= (layer1_outputs(3765)) and (layer1_outputs(7511));
    layer2_outputs(10814) <= layer1_outputs(5077);
    layer2_outputs(10815) <= not(layer1_outputs(3393));
    layer2_outputs(10816) <= not(layer1_outputs(5116)) or (layer1_outputs(1936));
    layer2_outputs(10817) <= not(layer1_outputs(2664));
    layer2_outputs(10818) <= not(layer1_outputs(11759));
    layer2_outputs(10819) <= not(layer1_outputs(8753));
    layer2_outputs(10820) <= not((layer1_outputs(1669)) and (layer1_outputs(11856)));
    layer2_outputs(10821) <= not(layer1_outputs(6932));
    layer2_outputs(10822) <= (layer1_outputs(4712)) and not (layer1_outputs(7669));
    layer2_outputs(10823) <= not(layer1_outputs(900));
    layer2_outputs(10824) <= not(layer1_outputs(11247)) or (layer1_outputs(5822));
    layer2_outputs(10825) <= not(layer1_outputs(9808));
    layer2_outputs(10826) <= '0';
    layer2_outputs(10827) <= layer1_outputs(980);
    layer2_outputs(10828) <= not(layer1_outputs(4712));
    layer2_outputs(10829) <= not(layer1_outputs(7877)) or (layer1_outputs(249));
    layer2_outputs(10830) <= not(layer1_outputs(9963)) or (layer1_outputs(5607));
    layer2_outputs(10831) <= (layer1_outputs(11852)) and (layer1_outputs(9829));
    layer2_outputs(10832) <= not((layer1_outputs(10023)) or (layer1_outputs(128)));
    layer2_outputs(10833) <= not((layer1_outputs(9417)) or (layer1_outputs(2264)));
    layer2_outputs(10834) <= layer1_outputs(3819);
    layer2_outputs(10835) <= (layer1_outputs(9556)) xor (layer1_outputs(8701));
    layer2_outputs(10836) <= layer1_outputs(74);
    layer2_outputs(10837) <= not(layer1_outputs(4674));
    layer2_outputs(10838) <= layer1_outputs(278);
    layer2_outputs(10839) <= not(layer1_outputs(12463));
    layer2_outputs(10840) <= layer1_outputs(879);
    layer2_outputs(10841) <= not(layer1_outputs(2914)) or (layer1_outputs(379));
    layer2_outputs(10842) <= not(layer1_outputs(12052));
    layer2_outputs(10843) <= not(layer1_outputs(9459));
    layer2_outputs(10844) <= not((layer1_outputs(2526)) xor (layer1_outputs(1961)));
    layer2_outputs(10845) <= not(layer1_outputs(4535));
    layer2_outputs(10846) <= layer1_outputs(2578);
    layer2_outputs(10847) <= not(layer1_outputs(10611));
    layer2_outputs(10848) <= not(layer1_outputs(4802));
    layer2_outputs(10849) <= not((layer1_outputs(6178)) xor (layer1_outputs(1879)));
    layer2_outputs(10850) <= not(layer1_outputs(11768));
    layer2_outputs(10851) <= not(layer1_outputs(3757));
    layer2_outputs(10852) <= layer1_outputs(2112);
    layer2_outputs(10853) <= (layer1_outputs(2920)) xor (layer1_outputs(11150));
    layer2_outputs(10854) <= (layer1_outputs(11996)) or (layer1_outputs(9948));
    layer2_outputs(10855) <= layer1_outputs(6295);
    layer2_outputs(10856) <= not((layer1_outputs(8432)) or (layer1_outputs(9802)));
    layer2_outputs(10857) <= layer1_outputs(4178);
    layer2_outputs(10858) <= not((layer1_outputs(12763)) or (layer1_outputs(237)));
    layer2_outputs(10859) <= not((layer1_outputs(4181)) xor (layer1_outputs(11419)));
    layer2_outputs(10860) <= layer1_outputs(2181);
    layer2_outputs(10861) <= (layer1_outputs(9559)) xor (layer1_outputs(4544));
    layer2_outputs(10862) <= not((layer1_outputs(8845)) xor (layer1_outputs(1671)));
    layer2_outputs(10863) <= layer1_outputs(2472);
    layer2_outputs(10864) <= not((layer1_outputs(7099)) and (layer1_outputs(1725)));
    layer2_outputs(10865) <= not(layer1_outputs(2882));
    layer2_outputs(10866) <= not(layer1_outputs(976));
    layer2_outputs(10867) <= not((layer1_outputs(12438)) or (layer1_outputs(2469)));
    layer2_outputs(10868) <= not(layer1_outputs(1420)) or (layer1_outputs(11509));
    layer2_outputs(10869) <= not((layer1_outputs(8179)) xor (layer1_outputs(8039)));
    layer2_outputs(10870) <= layer1_outputs(4707);
    layer2_outputs(10871) <= (layer1_outputs(621)) and (layer1_outputs(2441));
    layer2_outputs(10872) <= not(layer1_outputs(6354));
    layer2_outputs(10873) <= not((layer1_outputs(2696)) xor (layer1_outputs(3517)));
    layer2_outputs(10874) <= not(layer1_outputs(124));
    layer2_outputs(10875) <= layer1_outputs(3845);
    layer2_outputs(10876) <= not(layer1_outputs(8105));
    layer2_outputs(10877) <= layer1_outputs(11698);
    layer2_outputs(10878) <= not((layer1_outputs(11234)) and (layer1_outputs(98)));
    layer2_outputs(10879) <= (layer1_outputs(2718)) or (layer1_outputs(108));
    layer2_outputs(10880) <= not((layer1_outputs(11629)) and (layer1_outputs(6295)));
    layer2_outputs(10881) <= not(layer1_outputs(4498));
    layer2_outputs(10882) <= (layer1_outputs(10748)) and not (layer1_outputs(7715));
    layer2_outputs(10883) <= (layer1_outputs(2051)) xor (layer1_outputs(7358));
    layer2_outputs(10884) <= not(layer1_outputs(6213));
    layer2_outputs(10885) <= (layer1_outputs(2347)) and (layer1_outputs(1492));
    layer2_outputs(10886) <= (layer1_outputs(4640)) and (layer1_outputs(4084));
    layer2_outputs(10887) <= not((layer1_outputs(12387)) xor (layer1_outputs(10138)));
    layer2_outputs(10888) <= (layer1_outputs(5202)) and not (layer1_outputs(2896));
    layer2_outputs(10889) <= layer1_outputs(2079);
    layer2_outputs(10890) <= layer1_outputs(9343);
    layer2_outputs(10891) <= layer1_outputs(11229);
    layer2_outputs(10892) <= not(layer1_outputs(11752));
    layer2_outputs(10893) <= layer1_outputs(4061);
    layer2_outputs(10894) <= not(layer1_outputs(3747));
    layer2_outputs(10895) <= not(layer1_outputs(2012)) or (layer1_outputs(3264));
    layer2_outputs(10896) <= not((layer1_outputs(5466)) xor (layer1_outputs(929)));
    layer2_outputs(10897) <= (layer1_outputs(9407)) xor (layer1_outputs(11964));
    layer2_outputs(10898) <= (layer1_outputs(7877)) xor (layer1_outputs(5639));
    layer2_outputs(10899) <= layer1_outputs(6658);
    layer2_outputs(10900) <= not(layer1_outputs(3550));
    layer2_outputs(10901) <= layer1_outputs(10545);
    layer2_outputs(10902) <= not((layer1_outputs(4749)) or (layer1_outputs(10645)));
    layer2_outputs(10903) <= not(layer1_outputs(5960));
    layer2_outputs(10904) <= not(layer1_outputs(10712));
    layer2_outputs(10905) <= not(layer1_outputs(12427));
    layer2_outputs(10906) <= not(layer1_outputs(11189));
    layer2_outputs(10907) <= not(layer1_outputs(1079));
    layer2_outputs(10908) <= not(layer1_outputs(7798));
    layer2_outputs(10909) <= (layer1_outputs(11915)) and not (layer1_outputs(4912));
    layer2_outputs(10910) <= not(layer1_outputs(7103));
    layer2_outputs(10911) <= not((layer1_outputs(5066)) and (layer1_outputs(2983)));
    layer2_outputs(10912) <= not(layer1_outputs(2093));
    layer2_outputs(10913) <= layer1_outputs(10718);
    layer2_outputs(10914) <= (layer1_outputs(10057)) and not (layer1_outputs(9627));
    layer2_outputs(10915) <= not(layer1_outputs(5349));
    layer2_outputs(10916) <= not(layer1_outputs(10689));
    layer2_outputs(10917) <= not(layer1_outputs(9868)) or (layer1_outputs(8989));
    layer2_outputs(10918) <= not(layer1_outputs(10765)) or (layer1_outputs(10154));
    layer2_outputs(10919) <= layer1_outputs(5155);
    layer2_outputs(10920) <= layer1_outputs(8085);
    layer2_outputs(10921) <= not(layer1_outputs(7758));
    layer2_outputs(10922) <= not(layer1_outputs(4439));
    layer2_outputs(10923) <= not((layer1_outputs(6879)) or (layer1_outputs(7289)));
    layer2_outputs(10924) <= layer1_outputs(6853);
    layer2_outputs(10925) <= not((layer1_outputs(286)) xor (layer1_outputs(1287)));
    layer2_outputs(10926) <= (layer1_outputs(450)) xor (layer1_outputs(4450));
    layer2_outputs(10927) <= (layer1_outputs(3639)) and (layer1_outputs(6994));
    layer2_outputs(10928) <= not((layer1_outputs(6535)) or (layer1_outputs(6409)));
    layer2_outputs(10929) <= (layer1_outputs(1904)) xor (layer1_outputs(7906));
    layer2_outputs(10930) <= not(layer1_outputs(8512));
    layer2_outputs(10931) <= layer1_outputs(12367);
    layer2_outputs(10932) <= not(layer1_outputs(4836)) or (layer1_outputs(4189));
    layer2_outputs(10933) <= layer1_outputs(10659);
    layer2_outputs(10934) <= layer1_outputs(5918);
    layer2_outputs(10935) <= not((layer1_outputs(6713)) xor (layer1_outputs(11923)));
    layer2_outputs(10936) <= not((layer1_outputs(3352)) or (layer1_outputs(4769)));
    layer2_outputs(10937) <= layer1_outputs(2204);
    layer2_outputs(10938) <= not(layer1_outputs(5223));
    layer2_outputs(10939) <= (layer1_outputs(5334)) and (layer1_outputs(6858));
    layer2_outputs(10940) <= not((layer1_outputs(7592)) xor (layer1_outputs(8252)));
    layer2_outputs(10941) <= not(layer1_outputs(685));
    layer2_outputs(10942) <= layer1_outputs(9597);
    layer2_outputs(10943) <= layer1_outputs(955);
    layer2_outputs(10944) <= not(layer1_outputs(8782)) or (layer1_outputs(307));
    layer2_outputs(10945) <= layer1_outputs(6750);
    layer2_outputs(10946) <= layer1_outputs(4003);
    layer2_outputs(10947) <= not((layer1_outputs(2016)) xor (layer1_outputs(8447)));
    layer2_outputs(10948) <= not(layer1_outputs(5075));
    layer2_outputs(10949) <= not(layer1_outputs(1870));
    layer2_outputs(10950) <= not(layer1_outputs(10185)) or (layer1_outputs(10620));
    layer2_outputs(10951) <= not(layer1_outputs(8220));
    layer2_outputs(10952) <= not(layer1_outputs(2531));
    layer2_outputs(10953) <= layer1_outputs(8641);
    layer2_outputs(10954) <= not(layer1_outputs(12220));
    layer2_outputs(10955) <= layer1_outputs(10813);
    layer2_outputs(10956) <= not((layer1_outputs(6520)) xor (layer1_outputs(12100)));
    layer2_outputs(10957) <= (layer1_outputs(2248)) and not (layer1_outputs(11979));
    layer2_outputs(10958) <= layer1_outputs(6064);
    layer2_outputs(10959) <= not(layer1_outputs(11619));
    layer2_outputs(10960) <= (layer1_outputs(11896)) xor (layer1_outputs(11854));
    layer2_outputs(10961) <= not(layer1_outputs(4883));
    layer2_outputs(10962) <= (layer1_outputs(4413)) xor (layer1_outputs(5836));
    layer2_outputs(10963) <= not((layer1_outputs(4829)) xor (layer1_outputs(6939)));
    layer2_outputs(10964) <= not(layer1_outputs(2572));
    layer2_outputs(10965) <= (layer1_outputs(12441)) and not (layer1_outputs(11448));
    layer2_outputs(10966) <= not(layer1_outputs(4582)) or (layer1_outputs(1932));
    layer2_outputs(10967) <= (layer1_outputs(9433)) or (layer1_outputs(2415));
    layer2_outputs(10968) <= not((layer1_outputs(6680)) xor (layer1_outputs(959)));
    layer2_outputs(10969) <= not((layer1_outputs(1757)) xor (layer1_outputs(4074)));
    layer2_outputs(10970) <= (layer1_outputs(4561)) and not (layer1_outputs(6238));
    layer2_outputs(10971) <= layer1_outputs(9723);
    layer2_outputs(10972) <= layer1_outputs(8811);
    layer2_outputs(10973) <= (layer1_outputs(9705)) or (layer1_outputs(12450));
    layer2_outputs(10974) <= (layer1_outputs(7756)) and not (layer1_outputs(3700));
    layer2_outputs(10975) <= layer1_outputs(6367);
    layer2_outputs(10976) <= layer1_outputs(10022);
    layer2_outputs(10977) <= layer1_outputs(4577);
    layer2_outputs(10978) <= (layer1_outputs(1954)) xor (layer1_outputs(9828));
    layer2_outputs(10979) <= layer1_outputs(2087);
    layer2_outputs(10980) <= not(layer1_outputs(12764));
    layer2_outputs(10981) <= (layer1_outputs(1710)) and not (layer1_outputs(979));
    layer2_outputs(10982) <= layer1_outputs(1532);
    layer2_outputs(10983) <= layer1_outputs(7330);
    layer2_outputs(10984) <= not(layer1_outputs(2911)) or (layer1_outputs(12650));
    layer2_outputs(10985) <= layer1_outputs(10907);
    layer2_outputs(10986) <= not(layer1_outputs(4985));
    layer2_outputs(10987) <= layer1_outputs(718);
    layer2_outputs(10988) <= layer1_outputs(7041);
    layer2_outputs(10989) <= not(layer1_outputs(10665));
    layer2_outputs(10990) <= layer1_outputs(12699);
    layer2_outputs(10991) <= not((layer1_outputs(7240)) xor (layer1_outputs(3178)));
    layer2_outputs(10992) <= layer1_outputs(6723);
    layer2_outputs(10993) <= layer1_outputs(6018);
    layer2_outputs(10994) <= (layer1_outputs(6168)) and not (layer1_outputs(167));
    layer2_outputs(10995) <= not(layer1_outputs(8033));
    layer2_outputs(10996) <= (layer1_outputs(11861)) and (layer1_outputs(5792));
    layer2_outputs(10997) <= (layer1_outputs(4693)) or (layer1_outputs(3924));
    layer2_outputs(10998) <= not((layer1_outputs(2010)) xor (layer1_outputs(7995)));
    layer2_outputs(10999) <= not((layer1_outputs(9236)) xor (layer1_outputs(6552)));
    layer2_outputs(11000) <= layer1_outputs(10725);
    layer2_outputs(11001) <= not(layer1_outputs(12417));
    layer2_outputs(11002) <= (layer1_outputs(2078)) and not (layer1_outputs(7787));
    layer2_outputs(11003) <= not(layer1_outputs(4631));
    layer2_outputs(11004) <= (layer1_outputs(1098)) or (layer1_outputs(4830));
    layer2_outputs(11005) <= layer1_outputs(4752);
    layer2_outputs(11006) <= not(layer1_outputs(8567));
    layer2_outputs(11007) <= layer1_outputs(11373);
    layer2_outputs(11008) <= not((layer1_outputs(8942)) and (layer1_outputs(10379)));
    layer2_outputs(11009) <= not(layer1_outputs(11198)) or (layer1_outputs(2177));
    layer2_outputs(11010) <= not(layer1_outputs(1017));
    layer2_outputs(11011) <= not(layer1_outputs(4654)) or (layer1_outputs(11935));
    layer2_outputs(11012) <= (layer1_outputs(2924)) and (layer1_outputs(9427));
    layer2_outputs(11013) <= (layer1_outputs(216)) and not (layer1_outputs(5407));
    layer2_outputs(11014) <= not((layer1_outputs(2073)) and (layer1_outputs(591)));
    layer2_outputs(11015) <= (layer1_outputs(2141)) and (layer1_outputs(4722));
    layer2_outputs(11016) <= (layer1_outputs(3730)) and not (layer1_outputs(2209));
    layer2_outputs(11017) <= not((layer1_outputs(3720)) and (layer1_outputs(4069)));
    layer2_outputs(11018) <= not((layer1_outputs(11277)) and (layer1_outputs(7950)));
    layer2_outputs(11019) <= (layer1_outputs(3288)) or (layer1_outputs(12153));
    layer2_outputs(11020) <= (layer1_outputs(10827)) and not (layer1_outputs(1037));
    layer2_outputs(11021) <= not(layer1_outputs(11732));
    layer2_outputs(11022) <= layer1_outputs(2550);
    layer2_outputs(11023) <= not(layer1_outputs(11353));
    layer2_outputs(11024) <= (layer1_outputs(4272)) and not (layer1_outputs(7054));
    layer2_outputs(11025) <= not((layer1_outputs(465)) xor (layer1_outputs(2938)));
    layer2_outputs(11026) <= not(layer1_outputs(5933)) or (layer1_outputs(696));
    layer2_outputs(11027) <= not((layer1_outputs(12218)) and (layer1_outputs(7823)));
    layer2_outputs(11028) <= layer1_outputs(8661);
    layer2_outputs(11029) <= layer1_outputs(3394);
    layer2_outputs(11030) <= (layer1_outputs(6390)) xor (layer1_outputs(8005));
    layer2_outputs(11031) <= '0';
    layer2_outputs(11032) <= not(layer1_outputs(5457));
    layer2_outputs(11033) <= (layer1_outputs(1655)) xor (layer1_outputs(3076));
    layer2_outputs(11034) <= not((layer1_outputs(5867)) or (layer1_outputs(1507)));
    layer2_outputs(11035) <= not((layer1_outputs(5884)) or (layer1_outputs(12582)));
    layer2_outputs(11036) <= not(layer1_outputs(7735));
    layer2_outputs(11037) <= not((layer1_outputs(3380)) xor (layer1_outputs(11676)));
    layer2_outputs(11038) <= not(layer1_outputs(11177));
    layer2_outputs(11039) <= not(layer1_outputs(12078));
    layer2_outputs(11040) <= (layer1_outputs(1069)) xor (layer1_outputs(498));
    layer2_outputs(11041) <= not(layer1_outputs(8287));
    layer2_outputs(11042) <= not(layer1_outputs(6585));
    layer2_outputs(11043) <= '1';
    layer2_outputs(11044) <= not(layer1_outputs(4088));
    layer2_outputs(11045) <= (layer1_outputs(12288)) and not (layer1_outputs(10560));
    layer2_outputs(11046) <= not(layer1_outputs(8017));
    layer2_outputs(11047) <= (layer1_outputs(259)) and not (layer1_outputs(70));
    layer2_outputs(11048) <= not(layer1_outputs(9155));
    layer2_outputs(11049) <= layer1_outputs(11144);
    layer2_outputs(11050) <= layer1_outputs(10912);
    layer2_outputs(11051) <= layer1_outputs(6965);
    layer2_outputs(11052) <= not((layer1_outputs(6324)) and (layer1_outputs(9159)));
    layer2_outputs(11053) <= not(layer1_outputs(525));
    layer2_outputs(11054) <= not((layer1_outputs(3955)) xor (layer1_outputs(7329)));
    layer2_outputs(11055) <= layer1_outputs(6760);
    layer2_outputs(11056) <= not(layer1_outputs(4792)) or (layer1_outputs(1885));
    layer2_outputs(11057) <= not(layer1_outputs(10051));
    layer2_outputs(11058) <= layer1_outputs(977);
    layer2_outputs(11059) <= layer1_outputs(5598);
    layer2_outputs(11060) <= not(layer1_outputs(2753));
    layer2_outputs(11061) <= (layer1_outputs(2797)) and not (layer1_outputs(1594));
    layer2_outputs(11062) <= (layer1_outputs(5665)) xor (layer1_outputs(8343));
    layer2_outputs(11063) <= (layer1_outputs(9389)) and (layer1_outputs(8013));
    layer2_outputs(11064) <= (layer1_outputs(10978)) and not (layer1_outputs(9158));
    layer2_outputs(11065) <= (layer1_outputs(5298)) and not (layer1_outputs(2062));
    layer2_outputs(11066) <= layer1_outputs(10077);
    layer2_outputs(11067) <= not(layer1_outputs(2117));
    layer2_outputs(11068) <= not(layer1_outputs(1307));
    layer2_outputs(11069) <= layer1_outputs(3363);
    layer2_outputs(11070) <= not((layer1_outputs(97)) and (layer1_outputs(4134)));
    layer2_outputs(11071) <= (layer1_outputs(11155)) xor (layer1_outputs(6160));
    layer2_outputs(11072) <= not(layer1_outputs(4680));
    layer2_outputs(11073) <= not(layer1_outputs(9233)) or (layer1_outputs(2665));
    layer2_outputs(11074) <= (layer1_outputs(7788)) xor (layer1_outputs(7095));
    layer2_outputs(11075) <= layer1_outputs(663);
    layer2_outputs(11076) <= (layer1_outputs(9000)) or (layer1_outputs(1578));
    layer2_outputs(11077) <= not((layer1_outputs(8759)) and (layer1_outputs(7824)));
    layer2_outputs(11078) <= not(layer1_outputs(2201));
    layer2_outputs(11079) <= not(layer1_outputs(9432));
    layer2_outputs(11080) <= (layer1_outputs(7607)) and not (layer1_outputs(2494));
    layer2_outputs(11081) <= not(layer1_outputs(918));
    layer2_outputs(11082) <= layer1_outputs(6206);
    layer2_outputs(11083) <= not((layer1_outputs(5490)) xor (layer1_outputs(3844)));
    layer2_outputs(11084) <= layer1_outputs(10649);
    layer2_outputs(11085) <= (layer1_outputs(4909)) or (layer1_outputs(6923));
    layer2_outputs(11086) <= not(layer1_outputs(8717)) or (layer1_outputs(11165));
    layer2_outputs(11087) <= not((layer1_outputs(3520)) or (layer1_outputs(9042)));
    layer2_outputs(11088) <= not(layer1_outputs(11374)) or (layer1_outputs(3299));
    layer2_outputs(11089) <= layer1_outputs(1335);
    layer2_outputs(11090) <= not(layer1_outputs(10805));
    layer2_outputs(11091) <= not((layer1_outputs(21)) and (layer1_outputs(7106)));
    layer2_outputs(11092) <= not(layer1_outputs(4532));
    layer2_outputs(11093) <= layer1_outputs(4530);
    layer2_outputs(11094) <= (layer1_outputs(10798)) and not (layer1_outputs(7965));
    layer2_outputs(11095) <= not(layer1_outputs(5915)) or (layer1_outputs(10233));
    layer2_outputs(11096) <= (layer1_outputs(1729)) or (layer1_outputs(12738));
    layer2_outputs(11097) <= (layer1_outputs(9419)) and not (layer1_outputs(7602));
    layer2_outputs(11098) <= layer1_outputs(6487);
    layer2_outputs(11099) <= not((layer1_outputs(1037)) xor (layer1_outputs(2672)));
    layer2_outputs(11100) <= not(layer1_outputs(9763));
    layer2_outputs(11101) <= not((layer1_outputs(7342)) or (layer1_outputs(11316)));
    layer2_outputs(11102) <= layer1_outputs(1281);
    layer2_outputs(11103) <= not(layer1_outputs(4596));
    layer2_outputs(11104) <= not(layer1_outputs(5357));
    layer2_outputs(11105) <= (layer1_outputs(10)) xor (layer1_outputs(6557));
    layer2_outputs(11106) <= layer1_outputs(12444);
    layer2_outputs(11107) <= not(layer1_outputs(4987));
    layer2_outputs(11108) <= '1';
    layer2_outputs(11109) <= not((layer1_outputs(11582)) or (layer1_outputs(3986)));
    layer2_outputs(11110) <= layer1_outputs(6618);
    layer2_outputs(11111) <= (layer1_outputs(1506)) xor (layer1_outputs(11565));
    layer2_outputs(11112) <= (layer1_outputs(332)) and (layer1_outputs(6159));
    layer2_outputs(11113) <= not(layer1_outputs(172));
    layer2_outputs(11114) <= (layer1_outputs(3236)) and not (layer1_outputs(1911));
    layer2_outputs(11115) <= not((layer1_outputs(8999)) and (layer1_outputs(8711)));
    layer2_outputs(11116) <= (layer1_outputs(2802)) xor (layer1_outputs(7319));
    layer2_outputs(11117) <= (layer1_outputs(2081)) and not (layer1_outputs(9313));
    layer2_outputs(11118) <= not((layer1_outputs(2232)) xor (layer1_outputs(6073)));
    layer2_outputs(11119) <= layer1_outputs(12596);
    layer2_outputs(11120) <= not((layer1_outputs(847)) xor (layer1_outputs(1814)));
    layer2_outputs(11121) <= layer1_outputs(9738);
    layer2_outputs(11122) <= not((layer1_outputs(6023)) xor (layer1_outputs(2432)));
    layer2_outputs(11123) <= not(layer1_outputs(7480)) or (layer1_outputs(8757));
    layer2_outputs(11124) <= (layer1_outputs(11479)) xor (layer1_outputs(10196));
    layer2_outputs(11125) <= (layer1_outputs(3922)) xor (layer1_outputs(4423));
    layer2_outputs(11126) <= (layer1_outputs(11957)) and (layer1_outputs(1867));
    layer2_outputs(11127) <= not((layer1_outputs(9434)) xor (layer1_outputs(8247)));
    layer2_outputs(11128) <= not(layer1_outputs(2674));
    layer2_outputs(11129) <= layer1_outputs(6322);
    layer2_outputs(11130) <= layer1_outputs(10019);
    layer2_outputs(11131) <= (layer1_outputs(6935)) and not (layer1_outputs(8997));
    layer2_outputs(11132) <= not((layer1_outputs(11078)) xor (layer1_outputs(5686)));
    layer2_outputs(11133) <= layer1_outputs(6958);
    layer2_outputs(11134) <= not(layer1_outputs(12054));
    layer2_outputs(11135) <= layer1_outputs(5256);
    layer2_outputs(11136) <= (layer1_outputs(10987)) xor (layer1_outputs(9424));
    layer2_outputs(11137) <= not(layer1_outputs(4012));
    layer2_outputs(11138) <= not(layer1_outputs(9902));
    layer2_outputs(11139) <= layer1_outputs(1535);
    layer2_outputs(11140) <= not((layer1_outputs(6369)) or (layer1_outputs(3523)));
    layer2_outputs(11141) <= not(layer1_outputs(614)) or (layer1_outputs(1393));
    layer2_outputs(11142) <= layer1_outputs(1740);
    layer2_outputs(11143) <= layer1_outputs(11094);
    layer2_outputs(11144) <= (layer1_outputs(1289)) xor (layer1_outputs(9945));
    layer2_outputs(11145) <= (layer1_outputs(9722)) and (layer1_outputs(3323));
    layer2_outputs(11146) <= not(layer1_outputs(6059)) or (layer1_outputs(10958));
    layer2_outputs(11147) <= not(layer1_outputs(10166));
    layer2_outputs(11148) <= not((layer1_outputs(11605)) or (layer1_outputs(8499)));
    layer2_outputs(11149) <= layer1_outputs(6273);
    layer2_outputs(11150) <= layer1_outputs(1251);
    layer2_outputs(11151) <= not(layer1_outputs(377));
    layer2_outputs(11152) <= not(layer1_outputs(7271));
    layer2_outputs(11153) <= layer1_outputs(12230);
    layer2_outputs(11154) <= layer1_outputs(439);
    layer2_outputs(11155) <= not(layer1_outputs(5429));
    layer2_outputs(11156) <= not(layer1_outputs(1241));
    layer2_outputs(11157) <= layer1_outputs(11919);
    layer2_outputs(11158) <= (layer1_outputs(5608)) or (layer1_outputs(1445));
    layer2_outputs(11159) <= layer1_outputs(5433);
    layer2_outputs(11160) <= not(layer1_outputs(5871)) or (layer1_outputs(6088));
    layer2_outputs(11161) <= layer1_outputs(981);
    layer2_outputs(11162) <= layer1_outputs(6040);
    layer2_outputs(11163) <= (layer1_outputs(10610)) or (layer1_outputs(8678));
    layer2_outputs(11164) <= (layer1_outputs(7637)) xor (layer1_outputs(7381));
    layer2_outputs(11165) <= layer1_outputs(4244);
    layer2_outputs(11166) <= layer1_outputs(7601);
    layer2_outputs(11167) <= layer1_outputs(9285);
    layer2_outputs(11168) <= not(layer1_outputs(31));
    layer2_outputs(11169) <= layer1_outputs(5131);
    layer2_outputs(11170) <= layer1_outputs(12033);
    layer2_outputs(11171) <= not(layer1_outputs(12692));
    layer2_outputs(11172) <= (layer1_outputs(9858)) and not (layer1_outputs(4605));
    layer2_outputs(11173) <= (layer1_outputs(5309)) xor (layer1_outputs(84));
    layer2_outputs(11174) <= layer1_outputs(4689);
    layer2_outputs(11175) <= (layer1_outputs(7257)) xor (layer1_outputs(587));
    layer2_outputs(11176) <= layer1_outputs(9267);
    layer2_outputs(11177) <= (layer1_outputs(6188)) or (layer1_outputs(6569));
    layer2_outputs(11178) <= layer1_outputs(6632);
    layer2_outputs(11179) <= (layer1_outputs(5031)) and not (layer1_outputs(4984));
    layer2_outputs(11180) <= not((layer1_outputs(2094)) and (layer1_outputs(12691)));
    layer2_outputs(11181) <= not((layer1_outputs(9304)) xor (layer1_outputs(7656)));
    layer2_outputs(11182) <= not(layer1_outputs(1981));
    layer2_outputs(11183) <= layer1_outputs(11832);
    layer2_outputs(11184) <= not(layer1_outputs(385));
    layer2_outputs(11185) <= not((layer1_outputs(10445)) xor (layer1_outputs(10631)));
    layer2_outputs(11186) <= (layer1_outputs(5139)) and not (layer1_outputs(11862));
    layer2_outputs(11187) <= not(layer1_outputs(11521)) or (layer1_outputs(10520));
    layer2_outputs(11188) <= (layer1_outputs(10900)) and (layer1_outputs(3751));
    layer2_outputs(11189) <= layer1_outputs(4776);
    layer2_outputs(11190) <= (layer1_outputs(7305)) and not (layer1_outputs(920));
    layer2_outputs(11191) <= layer1_outputs(6231);
    layer2_outputs(11192) <= (layer1_outputs(7831)) or (layer1_outputs(4241));
    layer2_outputs(11193) <= (layer1_outputs(767)) and not (layer1_outputs(9397));
    layer2_outputs(11194) <= layer1_outputs(9663);
    layer2_outputs(11195) <= '1';
    layer2_outputs(11196) <= (layer1_outputs(10521)) xor (layer1_outputs(11955));
    layer2_outputs(11197) <= not((layer1_outputs(11251)) xor (layer1_outputs(8746)));
    layer2_outputs(11198) <= (layer1_outputs(145)) xor (layer1_outputs(3496));
    layer2_outputs(11199) <= (layer1_outputs(6711)) and (layer1_outputs(11492));
    layer2_outputs(11200) <= layer1_outputs(1499);
    layer2_outputs(11201) <= not((layer1_outputs(12536)) and (layer1_outputs(7866)));
    layer2_outputs(11202) <= (layer1_outputs(11244)) and (layer1_outputs(8316));
    layer2_outputs(11203) <= (layer1_outputs(11822)) and not (layer1_outputs(6849));
    layer2_outputs(11204) <= not(layer1_outputs(5899)) or (layer1_outputs(2913));
    layer2_outputs(11205) <= not((layer1_outputs(2144)) xor (layer1_outputs(1905)));
    layer2_outputs(11206) <= not(layer1_outputs(47));
    layer2_outputs(11207) <= not(layer1_outputs(6363));
    layer2_outputs(11208) <= not(layer1_outputs(11909));
    layer2_outputs(11209) <= layer1_outputs(3256);
    layer2_outputs(11210) <= not(layer1_outputs(380));
    layer2_outputs(11211) <= layer1_outputs(8127);
    layer2_outputs(11212) <= not((layer1_outputs(9785)) or (layer1_outputs(12414)));
    layer2_outputs(11213) <= not((layer1_outputs(12133)) xor (layer1_outputs(8659)));
    layer2_outputs(11214) <= not(layer1_outputs(9582));
    layer2_outputs(11215) <= not(layer1_outputs(5096)) or (layer1_outputs(12289));
    layer2_outputs(11216) <= (layer1_outputs(2927)) and not (layer1_outputs(2984));
    layer2_outputs(11217) <= not((layer1_outputs(10669)) or (layer1_outputs(7183)));
    layer2_outputs(11218) <= layer1_outputs(3037);
    layer2_outputs(11219) <= (layer1_outputs(871)) and not (layer1_outputs(4911));
    layer2_outputs(11220) <= (layer1_outputs(1706)) xor (layer1_outputs(6012));
    layer2_outputs(11221) <= layer1_outputs(3704);
    layer2_outputs(11222) <= not(layer1_outputs(3901));
    layer2_outputs(11223) <= not(layer1_outputs(10607));
    layer2_outputs(11224) <= (layer1_outputs(5035)) xor (layer1_outputs(5044));
    layer2_outputs(11225) <= not((layer1_outputs(1611)) or (layer1_outputs(12349)));
    layer2_outputs(11226) <= layer1_outputs(560);
    layer2_outputs(11227) <= not((layer1_outputs(6482)) and (layer1_outputs(11059)));
    layer2_outputs(11228) <= layer1_outputs(5887);
    layer2_outputs(11229) <= layer1_outputs(5286);
    layer2_outputs(11230) <= not((layer1_outputs(177)) xor (layer1_outputs(5058)));
    layer2_outputs(11231) <= (layer1_outputs(11701)) and (layer1_outputs(12361));
    layer2_outputs(11232) <= not((layer1_outputs(2328)) or (layer1_outputs(9912)));
    layer2_outputs(11233) <= not(layer1_outputs(4056));
    layer2_outputs(11234) <= not(layer1_outputs(1068));
    layer2_outputs(11235) <= not(layer1_outputs(4726)) or (layer1_outputs(10406));
    layer2_outputs(11236) <= (layer1_outputs(9658)) xor (layer1_outputs(2160));
    layer2_outputs(11237) <= not(layer1_outputs(11079));
    layer2_outputs(11238) <= layer1_outputs(12736);
    layer2_outputs(11239) <= not((layer1_outputs(10818)) and (layer1_outputs(3350)));
    layer2_outputs(11240) <= layer1_outputs(11227);
    layer2_outputs(11241) <= not(layer1_outputs(7739));
    layer2_outputs(11242) <= (layer1_outputs(8087)) xor (layer1_outputs(10673));
    layer2_outputs(11243) <= (layer1_outputs(3235)) and not (layer1_outputs(106));
    layer2_outputs(11244) <= (layer1_outputs(1226)) and not (layer1_outputs(3737));
    layer2_outputs(11245) <= (layer1_outputs(7193)) and not (layer1_outputs(7625));
    layer2_outputs(11246) <= not(layer1_outputs(7978)) or (layer1_outputs(988));
    layer2_outputs(11247) <= not(layer1_outputs(613)) or (layer1_outputs(8567));
    layer2_outputs(11248) <= not((layer1_outputs(5405)) xor (layer1_outputs(9156)));
    layer2_outputs(11249) <= layer1_outputs(11792);
    layer2_outputs(11250) <= (layer1_outputs(3367)) or (layer1_outputs(7274));
    layer2_outputs(11251) <= layer1_outputs(2766);
    layer2_outputs(11252) <= not(layer1_outputs(8276));
    layer2_outputs(11253) <= not(layer1_outputs(4580));
    layer2_outputs(11254) <= not(layer1_outputs(2731));
    layer2_outputs(11255) <= (layer1_outputs(1626)) and (layer1_outputs(2692));
    layer2_outputs(11256) <= layer1_outputs(9339);
    layer2_outputs(11257) <= layer1_outputs(3004);
    layer2_outputs(11258) <= not(layer1_outputs(8293)) or (layer1_outputs(6345));
    layer2_outputs(11259) <= (layer1_outputs(7301)) or (layer1_outputs(11364));
    layer2_outputs(11260) <= (layer1_outputs(9182)) or (layer1_outputs(11744));
    layer2_outputs(11261) <= (layer1_outputs(11535)) and (layer1_outputs(10455));
    layer2_outputs(11262) <= not(layer1_outputs(1733));
    layer2_outputs(11263) <= not((layer1_outputs(1034)) or (layer1_outputs(4016)));
    layer2_outputs(11264) <= layer1_outputs(11522);
    layer2_outputs(11265) <= layer1_outputs(3311);
    layer2_outputs(11266) <= layer1_outputs(2402);
    layer2_outputs(11267) <= not(layer1_outputs(5132));
    layer2_outputs(11268) <= not((layer1_outputs(8838)) or (layer1_outputs(1975)));
    layer2_outputs(11269) <= not(layer1_outputs(11990)) or (layer1_outputs(11301));
    layer2_outputs(11270) <= (layer1_outputs(9046)) and (layer1_outputs(12010));
    layer2_outputs(11271) <= layer1_outputs(8540);
    layer2_outputs(11272) <= layer1_outputs(9878);
    layer2_outputs(11273) <= '0';
    layer2_outputs(11274) <= layer1_outputs(12718);
    layer2_outputs(11275) <= (layer1_outputs(2993)) or (layer1_outputs(9834));
    layer2_outputs(11276) <= not((layer1_outputs(11272)) xor (layer1_outputs(754)));
    layer2_outputs(11277) <= not((layer1_outputs(12254)) xor (layer1_outputs(6921)));
    layer2_outputs(11278) <= (layer1_outputs(9616)) and (layer1_outputs(6517));
    layer2_outputs(11279) <= layer1_outputs(6212);
    layer2_outputs(11280) <= not(layer1_outputs(9282));
    layer2_outputs(11281) <= layer1_outputs(5951);
    layer2_outputs(11282) <= not((layer1_outputs(10908)) xor (layer1_outputs(3089)));
    layer2_outputs(11283) <= (layer1_outputs(346)) and not (layer1_outputs(9266));
    layer2_outputs(11284) <= not((layer1_outputs(7848)) xor (layer1_outputs(1317)));
    layer2_outputs(11285) <= not(layer1_outputs(5527));
    layer2_outputs(11286) <= not((layer1_outputs(12354)) xor (layer1_outputs(11008)));
    layer2_outputs(11287) <= (layer1_outputs(9569)) or (layer1_outputs(10774));
    layer2_outputs(11288) <= not((layer1_outputs(5111)) xor (layer1_outputs(2111)));
    layer2_outputs(11289) <= not(layer1_outputs(2998));
    layer2_outputs(11290) <= not(layer1_outputs(11349));
    layer2_outputs(11291) <= layer1_outputs(2007);
    layer2_outputs(11292) <= (layer1_outputs(2072)) and not (layer1_outputs(10329));
    layer2_outputs(11293) <= not(layer1_outputs(7522));
    layer2_outputs(11294) <= not(layer1_outputs(5943));
    layer2_outputs(11295) <= not(layer1_outputs(6309));
    layer2_outputs(11296) <= (layer1_outputs(7946)) xor (layer1_outputs(4156));
    layer2_outputs(11297) <= (layer1_outputs(12735)) and (layer1_outputs(11654));
    layer2_outputs(11298) <= not(layer1_outputs(6551));
    layer2_outputs(11299) <= not(layer1_outputs(12249));
    layer2_outputs(11300) <= layer1_outputs(3238);
    layer2_outputs(11301) <= not(layer1_outputs(6864));
    layer2_outputs(11302) <= not(layer1_outputs(12479));
    layer2_outputs(11303) <= not(layer1_outputs(6826)) or (layer1_outputs(10667));
    layer2_outputs(11304) <= not((layer1_outputs(8433)) or (layer1_outputs(1672)));
    layer2_outputs(11305) <= not((layer1_outputs(8330)) or (layer1_outputs(12032)));
    layer2_outputs(11306) <= (layer1_outputs(12454)) and (layer1_outputs(6337));
    layer2_outputs(11307) <= layer1_outputs(3879);
    layer2_outputs(11308) <= not((layer1_outputs(1361)) and (layer1_outputs(9543)));
    layer2_outputs(11309) <= not(layer1_outputs(11657));
    layer2_outputs(11310) <= layer1_outputs(6247);
    layer2_outputs(11311) <= not((layer1_outputs(5458)) xor (layer1_outputs(11448)));
    layer2_outputs(11312) <= not(layer1_outputs(7044));
    layer2_outputs(11313) <= layer1_outputs(6743);
    layer2_outputs(11314) <= (layer1_outputs(5531)) and not (layer1_outputs(2294));
    layer2_outputs(11315) <= (layer1_outputs(7747)) xor (layer1_outputs(12379));
    layer2_outputs(11316) <= (layer1_outputs(2310)) xor (layer1_outputs(8580));
    layer2_outputs(11317) <= not(layer1_outputs(11684)) or (layer1_outputs(4621));
    layer2_outputs(11318) <= (layer1_outputs(1897)) xor (layer1_outputs(9793));
    layer2_outputs(11319) <= layer1_outputs(6049);
    layer2_outputs(11320) <= '1';
    layer2_outputs(11321) <= layer1_outputs(5491);
    layer2_outputs(11322) <= not(layer1_outputs(5469));
    layer2_outputs(11323) <= (layer1_outputs(9768)) or (layer1_outputs(1));
    layer2_outputs(11324) <= not(layer1_outputs(5992));
    layer2_outputs(11325) <= layer1_outputs(8509);
    layer2_outputs(11326) <= (layer1_outputs(6619)) and not (layer1_outputs(4367));
    layer2_outputs(11327) <= layer1_outputs(5310);
    layer2_outputs(11328) <= not(layer1_outputs(9429));
    layer2_outputs(11329) <= not(layer1_outputs(4915));
    layer2_outputs(11330) <= (layer1_outputs(7749)) or (layer1_outputs(5000));
    layer2_outputs(11331) <= not(layer1_outputs(6197));
    layer2_outputs(11332) <= not(layer1_outputs(11724));
    layer2_outputs(11333) <= not(layer1_outputs(6655));
    layer2_outputs(11334) <= layer1_outputs(3878);
    layer2_outputs(11335) <= not(layer1_outputs(12632));
    layer2_outputs(11336) <= (layer1_outputs(9555)) or (layer1_outputs(6903));
    layer2_outputs(11337) <= not(layer1_outputs(147));
    layer2_outputs(11338) <= not((layer1_outputs(1757)) xor (layer1_outputs(6316)));
    layer2_outputs(11339) <= layer1_outputs(12259);
    layer2_outputs(11340) <= not((layer1_outputs(5719)) xor (layer1_outputs(6065)));
    layer2_outputs(11341) <= not(layer1_outputs(12129));
    layer2_outputs(11342) <= (layer1_outputs(3519)) xor (layer1_outputs(5810));
    layer2_outputs(11343) <= layer1_outputs(12157);
    layer2_outputs(11344) <= not(layer1_outputs(4208));
    layer2_outputs(11345) <= not(layer1_outputs(3960)) or (layer1_outputs(11906));
    layer2_outputs(11346) <= not((layer1_outputs(4905)) xor (layer1_outputs(3584)));
    layer2_outputs(11347) <= not(layer1_outputs(8179));
    layer2_outputs(11348) <= layer1_outputs(2882);
    layer2_outputs(11349) <= not(layer1_outputs(3496));
    layer2_outputs(11350) <= layer1_outputs(3679);
    layer2_outputs(11351) <= not((layer1_outputs(1378)) or (layer1_outputs(4223)));
    layer2_outputs(11352) <= layer1_outputs(5451);
    layer2_outputs(11353) <= not((layer1_outputs(10814)) and (layer1_outputs(531)));
    layer2_outputs(11354) <= layer1_outputs(10024);
    layer2_outputs(11355) <= not(layer1_outputs(4175));
    layer2_outputs(11356) <= (layer1_outputs(3199)) or (layer1_outputs(10557));
    layer2_outputs(11357) <= (layer1_outputs(1695)) and not (layer1_outputs(9935));
    layer2_outputs(11358) <= not(layer1_outputs(2546));
    layer2_outputs(11359) <= (layer1_outputs(1293)) or (layer1_outputs(2282));
    layer2_outputs(11360) <= layer1_outputs(12103);
    layer2_outputs(11361) <= not((layer1_outputs(11796)) or (layer1_outputs(2820)));
    layer2_outputs(11362) <= not(layer1_outputs(12355)) or (layer1_outputs(1851));
    layer2_outputs(11363) <= not((layer1_outputs(2323)) xor (layer1_outputs(11761)));
    layer2_outputs(11364) <= not(layer1_outputs(2017));
    layer2_outputs(11365) <= not((layer1_outputs(4187)) or (layer1_outputs(5662)));
    layer2_outputs(11366) <= layer1_outputs(8062);
    layer2_outputs(11367) <= not(layer1_outputs(1275)) or (layer1_outputs(11313));
    layer2_outputs(11368) <= layer1_outputs(9098);
    layer2_outputs(11369) <= (layer1_outputs(12465)) and (layer1_outputs(9177));
    layer2_outputs(11370) <= not(layer1_outputs(1598));
    layer2_outputs(11371) <= not((layer1_outputs(2357)) and (layer1_outputs(6315)));
    layer2_outputs(11372) <= (layer1_outputs(10472)) and not (layer1_outputs(6531));
    layer2_outputs(11373) <= layer1_outputs(8917);
    layer2_outputs(11374) <= not(layer1_outputs(9230));
    layer2_outputs(11375) <= not(layer1_outputs(3562));
    layer2_outputs(11376) <= not(layer1_outputs(3201));
    layer2_outputs(11377) <= (layer1_outputs(10121)) and (layer1_outputs(10231));
    layer2_outputs(11378) <= not(layer1_outputs(10536));
    layer2_outputs(11379) <= layer1_outputs(8076);
    layer2_outputs(11380) <= (layer1_outputs(2543)) and not (layer1_outputs(11349));
    layer2_outputs(11381) <= not(layer1_outputs(5714)) or (layer1_outputs(4134));
    layer2_outputs(11382) <= (layer1_outputs(7131)) and (layer1_outputs(8669));
    layer2_outputs(11383) <= layer1_outputs(11019);
    layer2_outputs(11384) <= (layer1_outputs(3029)) xor (layer1_outputs(11438));
    layer2_outputs(11385) <= not(layer1_outputs(1790));
    layer2_outputs(11386) <= not(layer1_outputs(611));
    layer2_outputs(11387) <= layer1_outputs(3680);
    layer2_outputs(11388) <= not(layer1_outputs(11645)) or (layer1_outputs(9607));
    layer2_outputs(11389) <= layer1_outputs(6545);
    layer2_outputs(11390) <= (layer1_outputs(7822)) and (layer1_outputs(3285));
    layer2_outputs(11391) <= (layer1_outputs(2809)) and not (layer1_outputs(4553));
    layer2_outputs(11392) <= not(layer1_outputs(6290));
    layer2_outputs(11393) <= (layer1_outputs(11467)) and not (layer1_outputs(11714));
    layer2_outputs(11394) <= (layer1_outputs(2010)) and not (layer1_outputs(5833));
    layer2_outputs(11395) <= (layer1_outputs(12768)) xor (layer1_outputs(5094));
    layer2_outputs(11396) <= layer1_outputs(324);
    layer2_outputs(11397) <= not((layer1_outputs(10654)) and (layer1_outputs(12121)));
    layer2_outputs(11398) <= layer1_outputs(9376);
    layer2_outputs(11399) <= (layer1_outputs(8652)) xor (layer1_outputs(11012));
    layer2_outputs(11400) <= not((layer1_outputs(10952)) or (layer1_outputs(11090)));
    layer2_outputs(11401) <= not(layer1_outputs(8399));
    layer2_outputs(11402) <= layer1_outputs(6709);
    layer2_outputs(11403) <= layer1_outputs(9723);
    layer2_outputs(11404) <= not(layer1_outputs(9704));
    layer2_outputs(11405) <= not((layer1_outputs(12482)) or (layer1_outputs(8166)));
    layer2_outputs(11406) <= not(layer1_outputs(2729));
    layer2_outputs(11407) <= layer1_outputs(3102);
    layer2_outputs(11408) <= not((layer1_outputs(10121)) xor (layer1_outputs(10346)));
    layer2_outputs(11409) <= (layer1_outputs(10365)) or (layer1_outputs(11982));
    layer2_outputs(11410) <= not(layer1_outputs(1321));
    layer2_outputs(11411) <= not((layer1_outputs(990)) or (layer1_outputs(1109)));
    layer2_outputs(11412) <= (layer1_outputs(1103)) and not (layer1_outputs(375));
    layer2_outputs(11413) <= (layer1_outputs(12351)) and not (layer1_outputs(12464));
    layer2_outputs(11414) <= (layer1_outputs(1104)) xor (layer1_outputs(556));
    layer2_outputs(11415) <= not((layer1_outputs(2501)) or (layer1_outputs(10590)));
    layer2_outputs(11416) <= not((layer1_outputs(8297)) or (layer1_outputs(7340)));
    layer2_outputs(11417) <= not(layer1_outputs(10351));
    layer2_outputs(11418) <= (layer1_outputs(3796)) xor (layer1_outputs(2627));
    layer2_outputs(11419) <= '1';
    layer2_outputs(11420) <= (layer1_outputs(5342)) and (layer1_outputs(12117));
    layer2_outputs(11421) <= not(layer1_outputs(9901)) or (layer1_outputs(2314));
    layer2_outputs(11422) <= not(layer1_outputs(10429));
    layer2_outputs(11423) <= not(layer1_outputs(678));
    layer2_outputs(11424) <= not(layer1_outputs(7577));
    layer2_outputs(11425) <= not(layer1_outputs(1522)) or (layer1_outputs(6774));
    layer2_outputs(11426) <= layer1_outputs(4481);
    layer2_outputs(11427) <= (layer1_outputs(3406)) and not (layer1_outputs(6774));
    layer2_outputs(11428) <= not(layer1_outputs(12503));
    layer2_outputs(11429) <= not((layer1_outputs(906)) or (layer1_outputs(360)));
    layer2_outputs(11430) <= (layer1_outputs(8873)) and not (layer1_outputs(6844));
    layer2_outputs(11431) <= (layer1_outputs(12765)) xor (layer1_outputs(3076));
    layer2_outputs(11432) <= not(layer1_outputs(10047)) or (layer1_outputs(8021));
    layer2_outputs(11433) <= not(layer1_outputs(11134));
    layer2_outputs(11434) <= layer1_outputs(5344);
    layer2_outputs(11435) <= not(layer1_outputs(1593));
    layer2_outputs(11436) <= (layer1_outputs(10376)) and (layer1_outputs(11797));
    layer2_outputs(11437) <= (layer1_outputs(4484)) and not (layer1_outputs(8310));
    layer2_outputs(11438) <= (layer1_outputs(5263)) xor (layer1_outputs(7785));
    layer2_outputs(11439) <= '0';
    layer2_outputs(11440) <= (layer1_outputs(10295)) xor (layer1_outputs(8926));
    layer2_outputs(11441) <= (layer1_outputs(12774)) or (layer1_outputs(10676));
    layer2_outputs(11442) <= not(layer1_outputs(2568));
    layer2_outputs(11443) <= not(layer1_outputs(1857));
    layer2_outputs(11444) <= not(layer1_outputs(11289));
    layer2_outputs(11445) <= not(layer1_outputs(6132));
    layer2_outputs(11446) <= not((layer1_outputs(2320)) xor (layer1_outputs(6312)));
    layer2_outputs(11447) <= layer1_outputs(4537);
    layer2_outputs(11448) <= layer1_outputs(5968);
    layer2_outputs(11449) <= layer1_outputs(5249);
    layer2_outputs(11450) <= not((layer1_outputs(8147)) or (layer1_outputs(9519)));
    layer2_outputs(11451) <= layer1_outputs(11176);
    layer2_outputs(11452) <= layer1_outputs(3811);
    layer2_outputs(11453) <= (layer1_outputs(310)) or (layer1_outputs(7712));
    layer2_outputs(11454) <= layer1_outputs(9995);
    layer2_outputs(11455) <= not((layer1_outputs(3776)) or (layer1_outputs(1284)));
    layer2_outputs(11456) <= not(layer1_outputs(7116));
    layer2_outputs(11457) <= layer1_outputs(832);
    layer2_outputs(11458) <= not(layer1_outputs(298));
    layer2_outputs(11459) <= not(layer1_outputs(3732));
    layer2_outputs(11460) <= not(layer1_outputs(12274));
    layer2_outputs(11461) <= not(layer1_outputs(5577));
    layer2_outputs(11462) <= layer1_outputs(6575);
    layer2_outputs(11463) <= layer1_outputs(8021);
    layer2_outputs(11464) <= not((layer1_outputs(128)) and (layer1_outputs(12632)));
    layer2_outputs(11465) <= (layer1_outputs(848)) xor (layer1_outputs(54));
    layer2_outputs(11466) <= not(layer1_outputs(8279));
    layer2_outputs(11467) <= not(layer1_outputs(518)) or (layer1_outputs(10533));
    layer2_outputs(11468) <= layer1_outputs(1305);
    layer2_outputs(11469) <= not(layer1_outputs(16));
    layer2_outputs(11470) <= (layer1_outputs(4493)) and not (layer1_outputs(2361));
    layer2_outputs(11471) <= not(layer1_outputs(3349));
    layer2_outputs(11472) <= not((layer1_outputs(7523)) or (layer1_outputs(4311)));
    layer2_outputs(11473) <= layer1_outputs(4627);
    layer2_outputs(11474) <= not(layer1_outputs(2041));
    layer2_outputs(11475) <= not((layer1_outputs(10106)) or (layer1_outputs(3823)));
    layer2_outputs(11476) <= not(layer1_outputs(1992));
    layer2_outputs(11477) <= not((layer1_outputs(6719)) or (layer1_outputs(5958)));
    layer2_outputs(11478) <= not(layer1_outputs(5074));
    layer2_outputs(11479) <= not(layer1_outputs(6935));
    layer2_outputs(11480) <= not(layer1_outputs(12255));
    layer2_outputs(11481) <= layer1_outputs(10614);
    layer2_outputs(11482) <= not(layer1_outputs(4891));
    layer2_outputs(11483) <= not((layer1_outputs(6598)) or (layer1_outputs(5141)));
    layer2_outputs(11484) <= layer1_outputs(10594);
    layer2_outputs(11485) <= not((layer1_outputs(5768)) and (layer1_outputs(8726)));
    layer2_outputs(11486) <= layer1_outputs(7179);
    layer2_outputs(11487) <= not(layer1_outputs(5197)) or (layer1_outputs(11574));
    layer2_outputs(11488) <= not(layer1_outputs(9251));
    layer2_outputs(11489) <= not(layer1_outputs(12715));
    layer2_outputs(11490) <= not(layer1_outputs(264));
    layer2_outputs(11491) <= (layer1_outputs(6483)) and not (layer1_outputs(4007));
    layer2_outputs(11492) <= layer1_outputs(7864);
    layer2_outputs(11493) <= (layer1_outputs(1107)) and not (layer1_outputs(8947));
    layer2_outputs(11494) <= layer1_outputs(12278);
    layer2_outputs(11495) <= (layer1_outputs(8303)) and not (layer1_outputs(363));
    layer2_outputs(11496) <= not(layer1_outputs(8647));
    layer2_outputs(11497) <= layer1_outputs(3057);
    layer2_outputs(11498) <= not(layer1_outputs(4363));
    layer2_outputs(11499) <= layer1_outputs(7461);
    layer2_outputs(11500) <= layer1_outputs(858);
    layer2_outputs(11501) <= not(layer1_outputs(2544));
    layer2_outputs(11502) <= layer1_outputs(2363);
    layer2_outputs(11503) <= not((layer1_outputs(3281)) or (layer1_outputs(11354)));
    layer2_outputs(11504) <= layer1_outputs(8144);
    layer2_outputs(11505) <= layer1_outputs(11058);
    layer2_outputs(11506) <= (layer1_outputs(10820)) or (layer1_outputs(7767));
    layer2_outputs(11507) <= (layer1_outputs(10243)) xor (layer1_outputs(4630));
    layer2_outputs(11508) <= not(layer1_outputs(7414));
    layer2_outputs(11509) <= not((layer1_outputs(7377)) and (layer1_outputs(9686)));
    layer2_outputs(11510) <= not(layer1_outputs(6234));
    layer2_outputs(11511) <= layer1_outputs(2251);
    layer2_outputs(11512) <= not((layer1_outputs(7937)) and (layer1_outputs(7462)));
    layer2_outputs(11513) <= (layer1_outputs(1033)) or (layer1_outputs(1408));
    layer2_outputs(11514) <= (layer1_outputs(700)) xor (layer1_outputs(9193));
    layer2_outputs(11515) <= layer1_outputs(3446);
    layer2_outputs(11516) <= (layer1_outputs(8014)) xor (layer1_outputs(2242));
    layer2_outputs(11517) <= layer1_outputs(11114);
    layer2_outputs(11518) <= (layer1_outputs(5173)) xor (layer1_outputs(6385));
    layer2_outputs(11519) <= layer1_outputs(2909);
    layer2_outputs(11520) <= not(layer1_outputs(6403));
    layer2_outputs(11521) <= (layer1_outputs(7170)) and (layer1_outputs(7298));
    layer2_outputs(11522) <= not((layer1_outputs(2242)) xor (layer1_outputs(302)));
    layer2_outputs(11523) <= layer1_outputs(5861);
    layer2_outputs(11524) <= not((layer1_outputs(8614)) and (layer1_outputs(8196)));
    layer2_outputs(11525) <= not((layer1_outputs(4443)) or (layer1_outputs(6037)));
    layer2_outputs(11526) <= not((layer1_outputs(9341)) xor (layer1_outputs(12343)));
    layer2_outputs(11527) <= layer1_outputs(4957);
    layer2_outputs(11528) <= layer1_outputs(11859);
    layer2_outputs(11529) <= layer1_outputs(1340);
    layer2_outputs(11530) <= layer1_outputs(1389);
    layer2_outputs(11531) <= not(layer1_outputs(7050)) or (layer1_outputs(4893));
    layer2_outputs(11532) <= not(layer1_outputs(6349));
    layer2_outputs(11533) <= not(layer1_outputs(4223));
    layer2_outputs(11534) <= layer1_outputs(328);
    layer2_outputs(11535) <= layer1_outputs(7876);
    layer2_outputs(11536) <= (layer1_outputs(5242)) xor (layer1_outputs(8535));
    layer2_outputs(11537) <= not((layer1_outputs(1380)) and (layer1_outputs(7643)));
    layer2_outputs(11538) <= (layer1_outputs(4976)) and not (layer1_outputs(2425));
    layer2_outputs(11539) <= not(layer1_outputs(269)) or (layer1_outputs(7155));
    layer2_outputs(11540) <= (layer1_outputs(10091)) or (layer1_outputs(11135));
    layer2_outputs(11541) <= not(layer1_outputs(5066));
    layer2_outputs(11542) <= (layer1_outputs(7421)) xor (layer1_outputs(2463));
    layer2_outputs(11543) <= not(layer1_outputs(11080));
    layer2_outputs(11544) <= layer1_outputs(4233);
    layer2_outputs(11545) <= not((layer1_outputs(1572)) or (layer1_outputs(1023)));
    layer2_outputs(11546) <= not(layer1_outputs(12268));
    layer2_outputs(11547) <= layer1_outputs(3821);
    layer2_outputs(11548) <= layer1_outputs(7363);
    layer2_outputs(11549) <= (layer1_outputs(6779)) and not (layer1_outputs(1174));
    layer2_outputs(11550) <= (layer1_outputs(8340)) xor (layer1_outputs(5082));
    layer2_outputs(11551) <= layer1_outputs(2517);
    layer2_outputs(11552) <= not((layer1_outputs(4675)) xor (layer1_outputs(11753)));
    layer2_outputs(11553) <= (layer1_outputs(743)) and (layer1_outputs(1857));
    layer2_outputs(11554) <= (layer1_outputs(6374)) and not (layer1_outputs(1161));
    layer2_outputs(11555) <= not((layer1_outputs(10916)) and (layer1_outputs(3598)));
    layer2_outputs(11556) <= not(layer1_outputs(9959));
    layer2_outputs(11557) <= layer1_outputs(727);
    layer2_outputs(11558) <= not(layer1_outputs(4569)) or (layer1_outputs(285));
    layer2_outputs(11559) <= not(layer1_outputs(528)) or (layer1_outputs(4961));
    layer2_outputs(11560) <= not((layer1_outputs(6290)) or (layer1_outputs(10486)));
    layer2_outputs(11561) <= (layer1_outputs(12302)) and (layer1_outputs(11059));
    layer2_outputs(11562) <= layer1_outputs(8081);
    layer2_outputs(11563) <= not((layer1_outputs(324)) and (layer1_outputs(9983)));
    layer2_outputs(11564) <= not((layer1_outputs(9533)) xor (layer1_outputs(5477)));
    layer2_outputs(11565) <= layer1_outputs(11088);
    layer2_outputs(11566) <= not(layer1_outputs(964)) or (layer1_outputs(10032));
    layer2_outputs(11567) <= (layer1_outputs(9349)) and not (layer1_outputs(451));
    layer2_outputs(11568) <= not((layer1_outputs(1063)) xor (layer1_outputs(477)));
    layer2_outputs(11569) <= not(layer1_outputs(2878));
    layer2_outputs(11570) <= (layer1_outputs(3030)) and not (layer1_outputs(7190));
    layer2_outputs(11571) <= (layer1_outputs(9330)) and not (layer1_outputs(12566));
    layer2_outputs(11572) <= not(layer1_outputs(8701));
    layer2_outputs(11573) <= (layer1_outputs(5975)) and (layer1_outputs(6962));
    layer2_outputs(11574) <= not(layer1_outputs(10545)) or (layer1_outputs(5841));
    layer2_outputs(11575) <= not(layer1_outputs(10749));
    layer2_outputs(11576) <= layer1_outputs(3396);
    layer2_outputs(11577) <= (layer1_outputs(5323)) and (layer1_outputs(1577));
    layer2_outputs(11578) <= not(layer1_outputs(1571));
    layer2_outputs(11579) <= (layer1_outputs(12347)) xor (layer1_outputs(4344));
    layer2_outputs(11580) <= not(layer1_outputs(8156)) or (layer1_outputs(7427));
    layer2_outputs(11581) <= (layer1_outputs(4538)) xor (layer1_outputs(9707));
    layer2_outputs(11582) <= not(layer1_outputs(1969));
    layer2_outputs(11583) <= not(layer1_outputs(10090));
    layer2_outputs(11584) <= not((layer1_outputs(10363)) or (layer1_outputs(1540)));
    layer2_outputs(11585) <= layer1_outputs(5464);
    layer2_outputs(11586) <= layer1_outputs(10902);
    layer2_outputs(11587) <= not(layer1_outputs(9601));
    layer2_outputs(11588) <= layer1_outputs(7251);
    layer2_outputs(11589) <= not(layer1_outputs(1412));
    layer2_outputs(11590) <= layer1_outputs(1078);
    layer2_outputs(11591) <= (layer1_outputs(9943)) and not (layer1_outputs(11270));
    layer2_outputs(11592) <= layer1_outputs(6488);
    layer2_outputs(11593) <= (layer1_outputs(12059)) xor (layer1_outputs(4389));
    layer2_outputs(11594) <= not(layer1_outputs(2710)) or (layer1_outputs(747));
    layer2_outputs(11595) <= layer1_outputs(1576);
    layer2_outputs(11596) <= layer1_outputs(9146);
    layer2_outputs(11597) <= not(layer1_outputs(10771));
    layer2_outputs(11598) <= layer1_outputs(1310);
    layer2_outputs(11599) <= not(layer1_outputs(3530));
    layer2_outputs(11600) <= (layer1_outputs(7607)) xor (layer1_outputs(10036));
    layer2_outputs(11601) <= layer1_outputs(12500);
    layer2_outputs(11602) <= not(layer1_outputs(5944));
    layer2_outputs(11603) <= not(layer1_outputs(3548));
    layer2_outputs(11604) <= layer1_outputs(9149);
    layer2_outputs(11605) <= layer1_outputs(12511);
    layer2_outputs(11606) <= not(layer1_outputs(11979));
    layer2_outputs(11607) <= (layer1_outputs(6255)) and not (layer1_outputs(8400));
    layer2_outputs(11608) <= layer1_outputs(10098);
    layer2_outputs(11609) <= layer1_outputs(11482);
    layer2_outputs(11610) <= layer1_outputs(6102);
    layer2_outputs(11611) <= not(layer1_outputs(9806));
    layer2_outputs(11612) <= not(layer1_outputs(2943)) or (layer1_outputs(5829));
    layer2_outputs(11613) <= layer1_outputs(1937);
    layer2_outputs(11614) <= not(layer1_outputs(3231));
    layer2_outputs(11615) <= (layer1_outputs(11685)) and not (layer1_outputs(4763));
    layer2_outputs(11616) <= layer1_outputs(11885);
    layer2_outputs(11617) <= not(layer1_outputs(10906)) or (layer1_outputs(7926));
    layer2_outputs(11618) <= (layer1_outputs(2607)) and not (layer1_outputs(4852));
    layer2_outputs(11619) <= not(layer1_outputs(3461));
    layer2_outputs(11620) <= (layer1_outputs(10174)) xor (layer1_outputs(10283));
    layer2_outputs(11621) <= layer1_outputs(11932);
    layer2_outputs(11622) <= not((layer1_outputs(943)) xor (layer1_outputs(3609)));
    layer2_outputs(11623) <= layer1_outputs(3900);
    layer2_outputs(11624) <= layer1_outputs(11280);
    layer2_outputs(11625) <= (layer1_outputs(1017)) and (layer1_outputs(11725));
    layer2_outputs(11626) <= not(layer1_outputs(2515));
    layer2_outputs(11627) <= (layer1_outputs(9568)) and (layer1_outputs(1563));
    layer2_outputs(11628) <= (layer1_outputs(3057)) xor (layer1_outputs(2056));
    layer2_outputs(11629) <= not((layer1_outputs(10883)) xor (layer1_outputs(9370)));
    layer2_outputs(11630) <= layer1_outputs(1211);
    layer2_outputs(11631) <= layer1_outputs(9139);
    layer2_outputs(11632) <= layer1_outputs(7611);
    layer2_outputs(11633) <= not(layer1_outputs(1772));
    layer2_outputs(11634) <= layer1_outputs(12594);
    layer2_outputs(11635) <= (layer1_outputs(4281)) or (layer1_outputs(10887));
    layer2_outputs(11636) <= layer1_outputs(597);
    layer2_outputs(11637) <= not(layer1_outputs(11613));
    layer2_outputs(11638) <= (layer1_outputs(5488)) xor (layer1_outputs(8181));
    layer2_outputs(11639) <= layer1_outputs(10384);
    layer2_outputs(11640) <= (layer1_outputs(4485)) and not (layer1_outputs(4499));
    layer2_outputs(11641) <= (layer1_outputs(344)) xor (layer1_outputs(715));
    layer2_outputs(11642) <= layer1_outputs(12253);
    layer2_outputs(11643) <= layer1_outputs(6973);
    layer2_outputs(11644) <= layer1_outputs(5145);
    layer2_outputs(11645) <= not(layer1_outputs(7806));
    layer2_outputs(11646) <= layer1_outputs(1189);
    layer2_outputs(11647) <= layer1_outputs(9070);
    layer2_outputs(11648) <= not(layer1_outputs(8626));
    layer2_outputs(11649) <= not((layer1_outputs(3664)) xor (layer1_outputs(1813)));
    layer2_outputs(11650) <= not(layer1_outputs(3646));
    layer2_outputs(11651) <= not(layer1_outputs(8150));
    layer2_outputs(11652) <= layer1_outputs(6003);
    layer2_outputs(11653) <= layer1_outputs(10302);
    layer2_outputs(11654) <= not((layer1_outputs(12286)) and (layer1_outputs(4954)));
    layer2_outputs(11655) <= not(layer1_outputs(11641));
    layer2_outputs(11656) <= not((layer1_outputs(698)) and (layer1_outputs(10637)));
    layer2_outputs(11657) <= not(layer1_outputs(1512));
    layer2_outputs(11658) <= (layer1_outputs(7810)) and not (layer1_outputs(6278));
    layer2_outputs(11659) <= not(layer1_outputs(3746));
    layer2_outputs(11660) <= not((layer1_outputs(11996)) xor (layer1_outputs(10759)));
    layer2_outputs(11661) <= not(layer1_outputs(12473));
    layer2_outputs(11662) <= (layer1_outputs(12699)) and not (layer1_outputs(12287));
    layer2_outputs(11663) <= not((layer1_outputs(2560)) xor (layer1_outputs(7812)));
    layer2_outputs(11664) <= (layer1_outputs(1213)) and not (layer1_outputs(1527));
    layer2_outputs(11665) <= layer1_outputs(4303);
    layer2_outputs(11666) <= layer1_outputs(12144);
    layer2_outputs(11667) <= layer1_outputs(4799);
    layer2_outputs(11668) <= not(layer1_outputs(10435));
    layer2_outputs(11669) <= not(layer1_outputs(6014));
    layer2_outputs(11670) <= not(layer1_outputs(12250));
    layer2_outputs(11671) <= (layer1_outputs(2414)) or (layer1_outputs(5949));
    layer2_outputs(11672) <= (layer1_outputs(8559)) and (layer1_outputs(2446));
    layer2_outputs(11673) <= not(layer1_outputs(10310));
    layer2_outputs(11674) <= (layer1_outputs(5765)) xor (layer1_outputs(9429));
    layer2_outputs(11675) <= not((layer1_outputs(12499)) xor (layer1_outputs(4487)));
    layer2_outputs(11676) <= layer1_outputs(1237);
    layer2_outputs(11677) <= not(layer1_outputs(5869));
    layer2_outputs(11678) <= not(layer1_outputs(1048)) or (layer1_outputs(11122));
    layer2_outputs(11679) <= (layer1_outputs(1510)) or (layer1_outputs(10522));
    layer2_outputs(11680) <= layer1_outputs(1914);
    layer2_outputs(11681) <= not((layer1_outputs(2766)) xor (layer1_outputs(7059)));
    layer2_outputs(11682) <= not(layer1_outputs(5525));
    layer2_outputs(11683) <= layer1_outputs(6820);
    layer2_outputs(11684) <= not(layer1_outputs(867));
    layer2_outputs(11685) <= not(layer1_outputs(10838)) or (layer1_outputs(9635));
    layer2_outputs(11686) <= (layer1_outputs(6875)) and not (layer1_outputs(2373));
    layer2_outputs(11687) <= not((layer1_outputs(5808)) and (layer1_outputs(9936)));
    layer2_outputs(11688) <= (layer1_outputs(1498)) and not (layer1_outputs(4330));
    layer2_outputs(11689) <= not((layer1_outputs(2050)) or (layer1_outputs(8485)));
    layer2_outputs(11690) <= not(layer1_outputs(8953));
    layer2_outputs(11691) <= layer1_outputs(8144);
    layer2_outputs(11692) <= (layer1_outputs(5908)) and not (layer1_outputs(236));
    layer2_outputs(11693) <= not((layer1_outputs(6869)) xor (layer1_outputs(7824)));
    layer2_outputs(11694) <= not((layer1_outputs(7628)) or (layer1_outputs(7562)));
    layer2_outputs(11695) <= layer1_outputs(1598);
    layer2_outputs(11696) <= layer1_outputs(11547);
    layer2_outputs(11697) <= not((layer1_outputs(3593)) xor (layer1_outputs(5806)));
    layer2_outputs(11698) <= not(layer1_outputs(11646));
    layer2_outputs(11699) <= layer1_outputs(11020);
    layer2_outputs(11700) <= not(layer1_outputs(8027));
    layer2_outputs(11701) <= not((layer1_outputs(12270)) and (layer1_outputs(10663)));
    layer2_outputs(11702) <= (layer1_outputs(479)) and not (layer1_outputs(1459));
    layer2_outputs(11703) <= layer1_outputs(5008);
    layer2_outputs(11704) <= (layer1_outputs(10508)) xor (layer1_outputs(1199));
    layer2_outputs(11705) <= not(layer1_outputs(5494));
    layer2_outputs(11706) <= not(layer1_outputs(4411));
    layer2_outputs(11707) <= layer1_outputs(287);
    layer2_outputs(11708) <= (layer1_outputs(423)) and (layer1_outputs(3194));
    layer2_outputs(11709) <= layer1_outputs(4978);
    layer2_outputs(11710) <= not(layer1_outputs(8327));
    layer2_outputs(11711) <= layer1_outputs(792);
    layer2_outputs(11712) <= not(layer1_outputs(3676));
    layer2_outputs(11713) <= not(layer1_outputs(9143));
    layer2_outputs(11714) <= layer1_outputs(7256);
    layer2_outputs(11715) <= not(layer1_outputs(10151));
    layer2_outputs(11716) <= layer1_outputs(6710);
    layer2_outputs(11717) <= layer1_outputs(10452);
    layer2_outputs(11718) <= not((layer1_outputs(1961)) xor (layer1_outputs(3321)));
    layer2_outputs(11719) <= layer1_outputs(5721);
    layer2_outputs(11720) <= not(layer1_outputs(8494)) or (layer1_outputs(6672));
    layer2_outputs(11721) <= not(layer1_outputs(5440));
    layer2_outputs(11722) <= layer1_outputs(5635);
    layer2_outputs(11723) <= not(layer1_outputs(10444));
    layer2_outputs(11724) <= layer1_outputs(4009);
    layer2_outputs(11725) <= not((layer1_outputs(8295)) or (layer1_outputs(3855)));
    layer2_outputs(11726) <= not(layer1_outputs(11342));
    layer2_outputs(11727) <= layer1_outputs(545);
    layer2_outputs(11728) <= (layer1_outputs(2059)) and (layer1_outputs(3973));
    layer2_outputs(11729) <= not(layer1_outputs(12700)) or (layer1_outputs(231));
    layer2_outputs(11730) <= layer1_outputs(8270);
    layer2_outputs(11731) <= layer1_outputs(11507);
    layer2_outputs(11732) <= (layer1_outputs(4611)) and not (layer1_outputs(8703));
    layer2_outputs(11733) <= not((layer1_outputs(7776)) and (layer1_outputs(5694)));
    layer2_outputs(11734) <= (layer1_outputs(4859)) xor (layer1_outputs(3335));
    layer2_outputs(11735) <= not(layer1_outputs(7777));
    layer2_outputs(11736) <= layer1_outputs(9659);
    layer2_outputs(11737) <= layer1_outputs(5509);
    layer2_outputs(11738) <= layer1_outputs(4974);
    layer2_outputs(11739) <= not(layer1_outputs(4563)) or (layer1_outputs(10797));
    layer2_outputs(11740) <= not((layer1_outputs(10891)) or (layer1_outputs(8048)));
    layer2_outputs(11741) <= not(layer1_outputs(827));
    layer2_outputs(11742) <= not(layer1_outputs(4986));
    layer2_outputs(11743) <= (layer1_outputs(6714)) xor (layer1_outputs(11418));
    layer2_outputs(11744) <= not(layer1_outputs(6913));
    layer2_outputs(11745) <= layer1_outputs(5630);
    layer2_outputs(11746) <= not((layer1_outputs(10556)) xor (layer1_outputs(8658)));
    layer2_outputs(11747) <= (layer1_outputs(203)) and not (layer1_outputs(6004));
    layer2_outputs(11748) <= layer1_outputs(9274);
    layer2_outputs(11749) <= layer1_outputs(7107);
    layer2_outputs(11750) <= not(layer1_outputs(10714)) or (layer1_outputs(4570));
    layer2_outputs(11751) <= not(layer1_outputs(3772));
    layer2_outputs(11752) <= '0';
    layer2_outputs(11753) <= not(layer1_outputs(10355));
    layer2_outputs(11754) <= layer1_outputs(6230);
    layer2_outputs(11755) <= not((layer1_outputs(765)) or (layer1_outputs(1538)));
    layer2_outputs(11756) <= not((layer1_outputs(10728)) xor (layer1_outputs(9123)));
    layer2_outputs(11757) <= not(layer1_outputs(5268));
    layer2_outputs(11758) <= not((layer1_outputs(8776)) and (layer1_outputs(10609)));
    layer2_outputs(11759) <= not(layer1_outputs(9915)) or (layer1_outputs(8450));
    layer2_outputs(11760) <= (layer1_outputs(1376)) and not (layer1_outputs(834));
    layer2_outputs(11761) <= not(layer1_outputs(908));
    layer2_outputs(11762) <= layer1_outputs(1491);
    layer2_outputs(11763) <= layer1_outputs(3370);
    layer2_outputs(11764) <= layer1_outputs(11377);
    layer2_outputs(11765) <= not(layer1_outputs(11165)) or (layer1_outputs(3587));
    layer2_outputs(11766) <= not((layer1_outputs(1713)) xor (layer1_outputs(185)));
    layer2_outputs(11767) <= layer1_outputs(7629);
    layer2_outputs(11768) <= layer1_outputs(1318);
    layer2_outputs(11769) <= layer1_outputs(6020);
    layer2_outputs(11770) <= not((layer1_outputs(11731)) xor (layer1_outputs(4997)));
    layer2_outputs(11771) <= (layer1_outputs(9065)) xor (layer1_outputs(10076));
    layer2_outputs(11772) <= not(layer1_outputs(5749));
    layer2_outputs(11773) <= not((layer1_outputs(3428)) xor (layer1_outputs(7863)));
    layer2_outputs(11774) <= not(layer1_outputs(6639));
    layer2_outputs(11775) <= not(layer1_outputs(1491));
    layer2_outputs(11776) <= layer1_outputs(8751);
    layer2_outputs(11777) <= (layer1_outputs(6759)) and not (layer1_outputs(4968));
    layer2_outputs(11778) <= layer1_outputs(8162);
    layer2_outputs(11779) <= (layer1_outputs(8743)) and not (layer1_outputs(2557));
    layer2_outputs(11780) <= not(layer1_outputs(2398));
    layer2_outputs(11781) <= (layer1_outputs(2308)) xor (layer1_outputs(12433));
    layer2_outputs(11782) <= (layer1_outputs(8890)) and not (layer1_outputs(12513));
    layer2_outputs(11783) <= not((layer1_outputs(4590)) and (layer1_outputs(11223)));
    layer2_outputs(11784) <= not((layer1_outputs(12231)) or (layer1_outputs(3086)));
    layer2_outputs(11785) <= layer1_outputs(9866);
    layer2_outputs(11786) <= not((layer1_outputs(11332)) xor (layer1_outputs(12356)));
    layer2_outputs(11787) <= not(layer1_outputs(11066));
    layer2_outputs(11788) <= not(layer1_outputs(7599));
    layer2_outputs(11789) <= not(layer1_outputs(12402)) or (layer1_outputs(11449));
    layer2_outputs(11790) <= (layer1_outputs(2014)) and not (layer1_outputs(2916));
    layer2_outputs(11791) <= layer1_outputs(9471);
    layer2_outputs(11792) <= layer1_outputs(8649);
    layer2_outputs(11793) <= layer1_outputs(10198);
    layer2_outputs(11794) <= not(layer1_outputs(1998));
    layer2_outputs(11795) <= layer1_outputs(2026);
    layer2_outputs(11796) <= not(layer1_outputs(11496));
    layer2_outputs(11797) <= not(layer1_outputs(5637));
    layer2_outputs(11798) <= (layer1_outputs(12024)) xor (layer1_outputs(12427));
    layer2_outputs(11799) <= not(layer1_outputs(3625));
    layer2_outputs(11800) <= not(layer1_outputs(10689));
    layer2_outputs(11801) <= not((layer1_outputs(4760)) and (layer1_outputs(10539)));
    layer2_outputs(11802) <= (layer1_outputs(41)) and not (layer1_outputs(5408));
    layer2_outputs(11803) <= not((layer1_outputs(8704)) xor (layer1_outputs(4827)));
    layer2_outputs(11804) <= layer1_outputs(14);
    layer2_outputs(11805) <= not(layer1_outputs(8705));
    layer2_outputs(11806) <= not(layer1_outputs(6776));
    layer2_outputs(11807) <= not((layer1_outputs(11751)) and (layer1_outputs(3617)));
    layer2_outputs(11808) <= (layer1_outputs(2086)) xor (layer1_outputs(7410));
    layer2_outputs(11809) <= not(layer1_outputs(11616));
    layer2_outputs(11810) <= (layer1_outputs(1028)) and not (layer1_outputs(6661));
    layer2_outputs(11811) <= not((layer1_outputs(11515)) or (layer1_outputs(11006)));
    layer2_outputs(11812) <= layer1_outputs(9436);
    layer2_outputs(11813) <= not((layer1_outputs(2193)) xor (layer1_outputs(10471)));
    layer2_outputs(11814) <= layer1_outputs(12543);
    layer2_outputs(11815) <= (layer1_outputs(3592)) and (layer1_outputs(1766));
    layer2_outputs(11816) <= not(layer1_outputs(5354)) or (layer1_outputs(9235));
    layer2_outputs(11817) <= not(layer1_outputs(12789)) or (layer1_outputs(4267));
    layer2_outputs(11818) <= not(layer1_outputs(7987));
    layer2_outputs(11819) <= not(layer1_outputs(12468));
    layer2_outputs(11820) <= not(layer1_outputs(6690)) or (layer1_outputs(5304));
    layer2_outputs(11821) <= (layer1_outputs(2462)) and (layer1_outputs(1674));
    layer2_outputs(11822) <= (layer1_outputs(7309)) and (layer1_outputs(5651));
    layer2_outputs(11823) <= (layer1_outputs(814)) xor (layer1_outputs(3917));
    layer2_outputs(11824) <= layer1_outputs(3210);
    layer2_outputs(11825) <= not(layer1_outputs(7686));
    layer2_outputs(11826) <= (layer1_outputs(7994)) or (layer1_outputs(8336));
    layer2_outputs(11827) <= not(layer1_outputs(9067));
    layer2_outputs(11828) <= not(layer1_outputs(11993));
    layer2_outputs(11829) <= not(layer1_outputs(12650));
    layer2_outputs(11830) <= '0';
    layer2_outputs(11831) <= (layer1_outputs(1796)) xor (layer1_outputs(8408));
    layer2_outputs(11832) <= (layer1_outputs(12673)) and (layer1_outputs(204));
    layer2_outputs(11833) <= (layer1_outputs(1838)) and not (layer1_outputs(1990));
    layer2_outputs(11834) <= not(layer1_outputs(4065));
    layer2_outputs(11835) <= layer1_outputs(9914);
    layer2_outputs(11836) <= (layer1_outputs(4960)) or (layer1_outputs(12431));
    layer2_outputs(11837) <= not(layer1_outputs(5321));
    layer2_outputs(11838) <= layer1_outputs(5723);
    layer2_outputs(11839) <= not(layer1_outputs(8261));
    layer2_outputs(11840) <= layer1_outputs(4236);
    layer2_outputs(11841) <= layer1_outputs(8830);
    layer2_outputs(11842) <= layer1_outputs(4874);
    layer2_outputs(11843) <= not(layer1_outputs(2111));
    layer2_outputs(11844) <= (layer1_outputs(5667)) and (layer1_outputs(3529));
    layer2_outputs(11845) <= not(layer1_outputs(7112)) or (layer1_outputs(12788));
    layer2_outputs(11846) <= (layer1_outputs(2654)) xor (layer1_outputs(2997));
    layer2_outputs(11847) <= (layer1_outputs(5897)) and (layer1_outputs(2029));
    layer2_outputs(11848) <= not((layer1_outputs(443)) or (layer1_outputs(3053)));
    layer2_outputs(11849) <= layer1_outputs(907);
    layer2_outputs(11850) <= not(layer1_outputs(5364));
    layer2_outputs(11851) <= not(layer1_outputs(11968));
    layer2_outputs(11852) <= (layer1_outputs(2065)) and (layer1_outputs(171));
    layer2_outputs(11853) <= not(layer1_outputs(9778));
    layer2_outputs(11854) <= (layer1_outputs(10470)) and not (layer1_outputs(9379));
    layer2_outputs(11855) <= not((layer1_outputs(7080)) xor (layer1_outputs(10151)));
    layer2_outputs(11856) <= layer1_outputs(4949);
    layer2_outputs(11857) <= not(layer1_outputs(4420));
    layer2_outputs(11858) <= layer1_outputs(9028);
    layer2_outputs(11859) <= not((layer1_outputs(4373)) xor (layer1_outputs(6184)));
    layer2_outputs(11860) <= layer1_outputs(5831);
    layer2_outputs(11861) <= (layer1_outputs(12639)) or (layer1_outputs(12165));
    layer2_outputs(11862) <= layer1_outputs(5989);
    layer2_outputs(11863) <= not(layer1_outputs(757));
    layer2_outputs(11864) <= not(layer1_outputs(8061)) or (layer1_outputs(7116));
    layer2_outputs(11865) <= (layer1_outputs(5819)) or (layer1_outputs(5902));
    layer2_outputs(11866) <= layer1_outputs(8288);
    layer2_outputs(11867) <= not(layer1_outputs(8364));
    layer2_outputs(11868) <= not((layer1_outputs(1843)) or (layer1_outputs(606)));
    layer2_outputs(11869) <= (layer1_outputs(3799)) or (layer1_outputs(2552));
    layer2_outputs(11870) <= not((layer1_outputs(8495)) xor (layer1_outputs(3391)));
    layer2_outputs(11871) <= not((layer1_outputs(708)) and (layer1_outputs(6698)));
    layer2_outputs(11872) <= not(layer1_outputs(12531));
    layer2_outputs(11873) <= not(layer1_outputs(8760));
    layer2_outputs(11874) <= (layer1_outputs(1953)) and (layer1_outputs(11055));
    layer2_outputs(11875) <= not(layer1_outputs(1421));
    layer2_outputs(11876) <= (layer1_outputs(9228)) and not (layer1_outputs(8482));
    layer2_outputs(11877) <= not(layer1_outputs(7796));
    layer2_outputs(11878) <= layer1_outputs(3065);
    layer2_outputs(11879) <= not(layer1_outputs(1875)) or (layer1_outputs(7282));
    layer2_outputs(11880) <= (layer1_outputs(12355)) and (layer1_outputs(8756));
    layer2_outputs(11881) <= (layer1_outputs(11917)) xor (layer1_outputs(5516));
    layer2_outputs(11882) <= not(layer1_outputs(10001)) or (layer1_outputs(4383));
    layer2_outputs(11883) <= not(layer1_outputs(2047)) or (layer1_outputs(8438));
    layer2_outputs(11884) <= (layer1_outputs(5909)) or (layer1_outputs(9310));
    layer2_outputs(11885) <= layer1_outputs(365);
    layer2_outputs(11886) <= (layer1_outputs(5372)) and not (layer1_outputs(3833));
    layer2_outputs(11887) <= not(layer1_outputs(5796));
    layer2_outputs(11888) <= not((layer1_outputs(11914)) or (layer1_outputs(9813)));
    layer2_outputs(11889) <= layer1_outputs(6957);
    layer2_outputs(11890) <= not((layer1_outputs(200)) or (layer1_outputs(9440)));
    layer2_outputs(11891) <= not(layer1_outputs(4241));
    layer2_outputs(11892) <= not(layer1_outputs(11875));
    layer2_outputs(11893) <= not((layer1_outputs(10056)) xor (layer1_outputs(7257)));
    layer2_outputs(11894) <= not(layer1_outputs(11513));
    layer2_outputs(11895) <= (layer1_outputs(8793)) and not (layer1_outputs(5431));
    layer2_outputs(11896) <= (layer1_outputs(9675)) or (layer1_outputs(5799));
    layer2_outputs(11897) <= not(layer1_outputs(12011));
    layer2_outputs(11898) <= not(layer1_outputs(1832));
    layer2_outputs(11899) <= (layer1_outputs(10854)) xor (layer1_outputs(4212));
    layer2_outputs(11900) <= (layer1_outputs(11057)) and not (layer1_outputs(3374));
    layer2_outputs(11901) <= not(layer1_outputs(8684)) or (layer1_outputs(10840));
    layer2_outputs(11902) <= not((layer1_outputs(7650)) and (layer1_outputs(817)));
    layer2_outputs(11903) <= not(layer1_outputs(9667));
    layer2_outputs(11904) <= (layer1_outputs(4376)) and not (layer1_outputs(4386));
    layer2_outputs(11905) <= layer1_outputs(6204);
    layer2_outputs(11906) <= layer1_outputs(10814);
    layer2_outputs(11907) <= layer1_outputs(138);
    layer2_outputs(11908) <= (layer1_outputs(8771)) xor (layer1_outputs(5965));
    layer2_outputs(11909) <= not(layer1_outputs(4410)) or (layer1_outputs(3921));
    layer2_outputs(11910) <= not(layer1_outputs(8304));
    layer2_outputs(11911) <= layer1_outputs(11143);
    layer2_outputs(11912) <= layer1_outputs(4584);
    layer2_outputs(11913) <= (layer1_outputs(10140)) or (layer1_outputs(1901));
    layer2_outputs(11914) <= not((layer1_outputs(4545)) or (layer1_outputs(5540)));
    layer2_outputs(11915) <= not(layer1_outputs(7236));
    layer2_outputs(11916) <= not((layer1_outputs(12343)) xor (layer1_outputs(2800)));
    layer2_outputs(11917) <= not(layer1_outputs(6666)) or (layer1_outputs(1358));
    layer2_outputs(11918) <= not((layer1_outputs(11684)) or (layer1_outputs(6151)));
    layer2_outputs(11919) <= (layer1_outputs(10161)) and (layer1_outputs(3479));
    layer2_outputs(11920) <= not(layer1_outputs(11098));
    layer2_outputs(11921) <= layer1_outputs(5048);
    layer2_outputs(11922) <= (layer1_outputs(3314)) or (layer1_outputs(8125));
    layer2_outputs(11923) <= layer1_outputs(11036);
    layer2_outputs(11924) <= not(layer1_outputs(8153));
    layer2_outputs(11925) <= not(layer1_outputs(12529));
    layer2_outputs(11926) <= not((layer1_outputs(3699)) or (layer1_outputs(5425)));
    layer2_outputs(11927) <= not((layer1_outputs(6032)) and (layer1_outputs(12092)));
    layer2_outputs(11928) <= (layer1_outputs(5345)) xor (layer1_outputs(9593));
    layer2_outputs(11929) <= layer1_outputs(4025);
    layer2_outputs(11930) <= layer1_outputs(4622);
    layer2_outputs(11931) <= layer1_outputs(5645);
    layer2_outputs(11932) <= not(layer1_outputs(10220));
    layer2_outputs(11933) <= not(layer1_outputs(8516)) or (layer1_outputs(272));
    layer2_outputs(11934) <= not(layer1_outputs(11672)) or (layer1_outputs(5629));
    layer2_outputs(11935) <= not((layer1_outputs(12009)) xor (layer1_outputs(6096)));
    layer2_outputs(11936) <= not((layer1_outputs(2061)) xor (layer1_outputs(6395)));
    layer2_outputs(11937) <= (layer1_outputs(4505)) or (layer1_outputs(4191));
    layer2_outputs(11938) <= not(layer1_outputs(12277));
    layer2_outputs(11939) <= not(layer1_outputs(590));
    layer2_outputs(11940) <= not(layer1_outputs(2133));
    layer2_outputs(11941) <= not((layer1_outputs(10804)) or (layer1_outputs(5310)));
    layer2_outputs(11942) <= layer1_outputs(8437);
    layer2_outputs(11943) <= (layer1_outputs(8029)) and (layer1_outputs(2553));
    layer2_outputs(11944) <= layer1_outputs(4868);
    layer2_outputs(11945) <= (layer1_outputs(9005)) and not (layer1_outputs(1910));
    layer2_outputs(11946) <= not(layer1_outputs(8446)) or (layer1_outputs(10474));
    layer2_outputs(11947) <= not((layer1_outputs(11342)) xor (layer1_outputs(10768)));
    layer2_outputs(11948) <= layer1_outputs(2221);
    layer2_outputs(11949) <= not(layer1_outputs(1364));
    layer2_outputs(11950) <= not(layer1_outputs(6015));
    layer2_outputs(11951) <= not((layer1_outputs(7535)) and (layer1_outputs(2181)));
    layer2_outputs(11952) <= (layer1_outputs(6662)) xor (layer1_outputs(9280));
    layer2_outputs(11953) <= layer1_outputs(7126);
    layer2_outputs(11954) <= layer1_outputs(3910);
    layer2_outputs(11955) <= layer1_outputs(11954);
    layer2_outputs(11956) <= not(layer1_outputs(1765));
    layer2_outputs(11957) <= not(layer1_outputs(1520)) or (layer1_outputs(10146));
    layer2_outputs(11958) <= layer1_outputs(8442);
    layer2_outputs(11959) <= not(layer1_outputs(552));
    layer2_outputs(11960) <= (layer1_outputs(8053)) xor (layer1_outputs(8883));
    layer2_outputs(11961) <= (layer1_outputs(6678)) and not (layer1_outputs(12461));
    layer2_outputs(11962) <= not(layer1_outputs(404));
    layer2_outputs(11963) <= (layer1_outputs(9425)) and (layer1_outputs(5576));
    layer2_outputs(11964) <= (layer1_outputs(12396)) and not (layer1_outputs(1930));
    layer2_outputs(11965) <= not(layer1_outputs(8800));
    layer2_outputs(11966) <= (layer1_outputs(1807)) xor (layer1_outputs(12301));
    layer2_outputs(11967) <= not(layer1_outputs(8300));
    layer2_outputs(11968) <= layer1_outputs(11652);
    layer2_outputs(11969) <= not(layer1_outputs(12161));
    layer2_outputs(11970) <= layer1_outputs(2745);
    layer2_outputs(11971) <= not((layer1_outputs(8180)) or (layer1_outputs(369)));
    layer2_outputs(11972) <= (layer1_outputs(6485)) and not (layer1_outputs(6257));
    layer2_outputs(11973) <= not(layer1_outputs(7050)) or (layer1_outputs(1209));
    layer2_outputs(11974) <= not(layer1_outputs(5779)) or (layer1_outputs(9309));
    layer2_outputs(11975) <= not(layer1_outputs(8152)) or (layer1_outputs(1514));
    layer2_outputs(11976) <= not(layer1_outputs(7461)) or (layer1_outputs(8408));
    layer2_outputs(11977) <= layer1_outputs(1297);
    layer2_outputs(11978) <= layer1_outputs(4234);
    layer2_outputs(11979) <= layer1_outputs(9604);
    layer2_outputs(11980) <= layer1_outputs(1283);
    layer2_outputs(11981) <= not((layer1_outputs(3395)) xor (layer1_outputs(9481)));
    layer2_outputs(11982) <= layer1_outputs(11398);
    layer2_outputs(11983) <= layer1_outputs(7609);
    layer2_outputs(11984) <= layer1_outputs(833);
    layer2_outputs(11985) <= (layer1_outputs(933)) and not (layer1_outputs(5373));
    layer2_outputs(11986) <= not(layer1_outputs(1984));
    layer2_outputs(11987) <= not(layer1_outputs(6493)) or (layer1_outputs(4442));
    layer2_outputs(11988) <= layer1_outputs(12782);
    layer2_outputs(11989) <= (layer1_outputs(1029)) and not (layer1_outputs(9974));
    layer2_outputs(11990) <= (layer1_outputs(720)) and (layer1_outputs(5127));
    layer2_outputs(11991) <= not(layer1_outputs(2554));
    layer2_outputs(11992) <= not((layer1_outputs(2230)) or (layer1_outputs(4746)));
    layer2_outputs(11993) <= layer1_outputs(8099);
    layer2_outputs(11994) <= '0';
    layer2_outputs(11995) <= not(layer1_outputs(2145));
    layer2_outputs(11996) <= not(layer1_outputs(8766));
    layer2_outputs(11997) <= not(layer1_outputs(2218));
    layer2_outputs(11998) <= not(layer1_outputs(11754));
    layer2_outputs(11999) <= layer1_outputs(2767);
    layer2_outputs(12000) <= not((layer1_outputs(7475)) and (layer1_outputs(5679)));
    layer2_outputs(12001) <= not((layer1_outputs(3946)) or (layer1_outputs(935)));
    layer2_outputs(12002) <= layer1_outputs(9229);
    layer2_outputs(12003) <= layer1_outputs(6715);
    layer2_outputs(12004) <= (layer1_outputs(4832)) xor (layer1_outputs(7483));
    layer2_outputs(12005) <= not(layer1_outputs(9133));
    layer2_outputs(12006) <= (layer1_outputs(12578)) xor (layer1_outputs(9337));
    layer2_outputs(12007) <= not(layer1_outputs(2239)) or (layer1_outputs(1027));
    layer2_outputs(12008) <= (layer1_outputs(12214)) xor (layer1_outputs(10621));
    layer2_outputs(12009) <= (layer1_outputs(4805)) and not (layer1_outputs(11152));
    layer2_outputs(12010) <= not(layer1_outputs(6878));
    layer2_outputs(12011) <= not(layer1_outputs(5503));
    layer2_outputs(12012) <= not(layer1_outputs(6150));
    layer2_outputs(12013) <= not(layer1_outputs(3868));
    layer2_outputs(12014) <= (layer1_outputs(5183)) and not (layer1_outputs(7795));
    layer2_outputs(12015) <= layer1_outputs(11423);
    layer2_outputs(12016) <= (layer1_outputs(8008)) or (layer1_outputs(6125));
    layer2_outputs(12017) <= layer1_outputs(5082);
    layer2_outputs(12018) <= '0';
    layer2_outputs(12019) <= (layer1_outputs(11565)) and not (layer1_outputs(763));
    layer2_outputs(12020) <= (layer1_outputs(7234)) xor (layer1_outputs(8443));
    layer2_outputs(12021) <= not(layer1_outputs(957));
    layer2_outputs(12022) <= '1';
    layer2_outputs(12023) <= layer1_outputs(5015);
    layer2_outputs(12024) <= layer1_outputs(11762);
    layer2_outputs(12025) <= not(layer1_outputs(7526));
    layer2_outputs(12026) <= (layer1_outputs(7275)) or (layer1_outputs(8234));
    layer2_outputs(12027) <= (layer1_outputs(2039)) xor (layer1_outputs(6186));
    layer2_outputs(12028) <= (layer1_outputs(11543)) and not (layer1_outputs(11452));
    layer2_outputs(12029) <= not(layer1_outputs(3645));
    layer2_outputs(12030) <= (layer1_outputs(4265)) or (layer1_outputs(10073));
    layer2_outputs(12031) <= layer1_outputs(12206);
    layer2_outputs(12032) <= not(layer1_outputs(2525));
    layer2_outputs(12033) <= not(layer1_outputs(9111));
    layer2_outputs(12034) <= not((layer1_outputs(4229)) or (layer1_outputs(10601)));
    layer2_outputs(12035) <= (layer1_outputs(4157)) xor (layer1_outputs(3213));
    layer2_outputs(12036) <= not((layer1_outputs(1480)) xor (layer1_outputs(3833)));
    layer2_outputs(12037) <= not((layer1_outputs(10946)) xor (layer1_outputs(9947)));
    layer2_outputs(12038) <= not(layer1_outputs(6284)) or (layer1_outputs(11776));
    layer2_outputs(12039) <= layer1_outputs(10535);
    layer2_outputs(12040) <= not((layer1_outputs(849)) xor (layer1_outputs(9772)));
    layer2_outputs(12041) <= layer1_outputs(9774);
    layer2_outputs(12042) <= not(layer1_outputs(1428)) or (layer1_outputs(11854));
    layer2_outputs(12043) <= not(layer1_outputs(8375));
    layer2_outputs(12044) <= layer1_outputs(10010);
    layer2_outputs(12045) <= not(layer1_outputs(3310));
    layer2_outputs(12046) <= layer1_outputs(5487);
    layer2_outputs(12047) <= not(layer1_outputs(5481)) or (layer1_outputs(4540));
    layer2_outputs(12048) <= not(layer1_outputs(5991));
    layer2_outputs(12049) <= not((layer1_outputs(10923)) or (layer1_outputs(8415)));
    layer2_outputs(12050) <= layer1_outputs(7433);
    layer2_outputs(12051) <= not((layer1_outputs(3985)) or (layer1_outputs(9670)));
    layer2_outputs(12052) <= not(layer1_outputs(5471));
    layer2_outputs(12053) <= (layer1_outputs(7853)) or (layer1_outputs(12078));
    layer2_outputs(12054) <= not(layer1_outputs(1330)) or (layer1_outputs(8078));
    layer2_outputs(12055) <= layer1_outputs(3082);
    layer2_outputs(12056) <= layer1_outputs(10350);
    layer2_outputs(12057) <= not((layer1_outputs(7329)) and (layer1_outputs(12131)));
    layer2_outputs(12058) <= layer1_outputs(11771);
    layer2_outputs(12059) <= (layer1_outputs(8398)) and not (layer1_outputs(4486));
    layer2_outputs(12060) <= not(layer1_outputs(5515)) or (layer1_outputs(8255));
    layer2_outputs(12061) <= not(layer1_outputs(9586));
    layer2_outputs(12062) <= not(layer1_outputs(12401));
    layer2_outputs(12063) <= not(layer1_outputs(7947)) or (layer1_outputs(4784));
    layer2_outputs(12064) <= layer1_outputs(9556);
    layer2_outputs(12065) <= layer1_outputs(6381);
    layer2_outputs(12066) <= not(layer1_outputs(729)) or (layer1_outputs(4747));
    layer2_outputs(12067) <= not(layer1_outputs(10341)) or (layer1_outputs(7983));
    layer2_outputs(12068) <= not((layer1_outputs(8443)) and (layer1_outputs(2241)));
    layer2_outputs(12069) <= not((layer1_outputs(8247)) xor (layer1_outputs(504)));
    layer2_outputs(12070) <= not((layer1_outputs(6272)) and (layer1_outputs(7958)));
    layer2_outputs(12071) <= not(layer1_outputs(6243));
    layer2_outputs(12072) <= not((layer1_outputs(637)) xor (layer1_outputs(8941)));
    layer2_outputs(12073) <= not(layer1_outputs(11011));
    layer2_outputs(12074) <= (layer1_outputs(4256)) or (layer1_outputs(10981));
    layer2_outputs(12075) <= (layer1_outputs(5756)) and not (layer1_outputs(8207));
    layer2_outputs(12076) <= layer1_outputs(3884);
    layer2_outputs(12077) <= layer1_outputs(10641);
    layer2_outputs(12078) <= (layer1_outputs(25)) xor (layer1_outputs(6326));
    layer2_outputs(12079) <= layer1_outputs(10895);
    layer2_outputs(12080) <= layer1_outputs(1343);
    layer2_outputs(12081) <= (layer1_outputs(1662)) xor (layer1_outputs(9168));
    layer2_outputs(12082) <= not(layer1_outputs(7746));
    layer2_outputs(12083) <= (layer1_outputs(6423)) xor (layer1_outputs(4388));
    layer2_outputs(12084) <= layer1_outputs(253);
    layer2_outputs(12085) <= (layer1_outputs(2604)) and not (layer1_outputs(3422));
    layer2_outputs(12086) <= (layer1_outputs(10715)) and not (layer1_outputs(2174));
    layer2_outputs(12087) <= not(layer1_outputs(12340));
    layer2_outputs(12088) <= not(layer1_outputs(3158));
    layer2_outputs(12089) <= not((layer1_outputs(2776)) xor (layer1_outputs(3526)));
    layer2_outputs(12090) <= not(layer1_outputs(12058));
    layer2_outputs(12091) <= (layer1_outputs(10382)) or (layer1_outputs(1225));
    layer2_outputs(12092) <= layer1_outputs(8556);
    layer2_outputs(12093) <= layer1_outputs(681);
    layer2_outputs(12094) <= not((layer1_outputs(9035)) xor (layer1_outputs(5109)));
    layer2_outputs(12095) <= not(layer1_outputs(12477));
    layer2_outputs(12096) <= not(layer1_outputs(5341)) or (layer1_outputs(10341));
    layer2_outputs(12097) <= (layer1_outputs(86)) and not (layer1_outputs(10163));
    layer2_outputs(12098) <= layer1_outputs(9614);
    layer2_outputs(12099) <= layer1_outputs(2783);
    layer2_outputs(12100) <= (layer1_outputs(9321)) or (layer1_outputs(10082));
    layer2_outputs(12101) <= layer1_outputs(2021);
    layer2_outputs(12102) <= not((layer1_outputs(847)) and (layer1_outputs(11790)));
    layer2_outputs(12103) <= (layer1_outputs(3977)) xor (layer1_outputs(796));
    layer2_outputs(12104) <= (layer1_outputs(2135)) and not (layer1_outputs(2261));
    layer2_outputs(12105) <= (layer1_outputs(3443)) and (layer1_outputs(8908));
    layer2_outputs(12106) <= not(layer1_outputs(5647)) or (layer1_outputs(2481));
    layer2_outputs(12107) <= layer1_outputs(7693);
    layer2_outputs(12108) <= not(layer1_outputs(3248)) or (layer1_outputs(7479));
    layer2_outputs(12109) <= not((layer1_outputs(4713)) xor (layer1_outputs(11380)));
    layer2_outputs(12110) <= layer1_outputs(1927);
    layer2_outputs(12111) <= (layer1_outputs(12145)) xor (layer1_outputs(1164));
    layer2_outputs(12112) <= not(layer1_outputs(122)) or (layer1_outputs(6746));
    layer2_outputs(12113) <= layer1_outputs(10468);
    layer2_outputs(12114) <= layer1_outputs(740);
    layer2_outputs(12115) <= not((layer1_outputs(2388)) and (layer1_outputs(11544)));
    layer2_outputs(12116) <= not(layer1_outputs(2815));
    layer2_outputs(12117) <= layer1_outputs(10210);
    layer2_outputs(12118) <= layer1_outputs(3349);
    layer2_outputs(12119) <= not(layer1_outputs(2064));
    layer2_outputs(12120) <= layer1_outputs(2866);
    layer2_outputs(12121) <= not(layer1_outputs(3474)) or (layer1_outputs(10242));
    layer2_outputs(12122) <= not(layer1_outputs(9627)) or (layer1_outputs(3886));
    layer2_outputs(12123) <= (layer1_outputs(2551)) and not (layer1_outputs(12164));
    layer2_outputs(12124) <= (layer1_outputs(8600)) xor (layer1_outputs(11618));
    layer2_outputs(12125) <= layer1_outputs(9479);
    layer2_outputs(12126) <= (layer1_outputs(3631)) and (layer1_outputs(6495));
    layer2_outputs(12127) <= not((layer1_outputs(6870)) xor (layer1_outputs(3733)));
    layer2_outputs(12128) <= layer1_outputs(8137);
    layer2_outputs(12129) <= not((layer1_outputs(10746)) and (layer1_outputs(5203)));
    layer2_outputs(12130) <= not((layer1_outputs(4920)) xor (layer1_outputs(7813)));
    layer2_outputs(12131) <= not((layer1_outputs(4801)) xor (layer1_outputs(5732)));
    layer2_outputs(12132) <= not((layer1_outputs(1438)) or (layer1_outputs(578)));
    layer2_outputs(12133) <= not((layer1_outputs(9209)) and (layer1_outputs(8682)));
    layer2_outputs(12134) <= not(layer1_outputs(8335));
    layer2_outputs(12135) <= layer1_outputs(11815);
    layer2_outputs(12136) <= layer1_outputs(9656);
    layer2_outputs(12137) <= not(layer1_outputs(9093)) or (layer1_outputs(1919));
    layer2_outputs(12138) <= layer1_outputs(2683);
    layer2_outputs(12139) <= not((layer1_outputs(3353)) or (layer1_outputs(7209)));
    layer2_outputs(12140) <= (layer1_outputs(6458)) and not (layer1_outputs(0));
    layer2_outputs(12141) <= not(layer1_outputs(1697)) or (layer1_outputs(147));
    layer2_outputs(12142) <= layer1_outputs(3077);
    layer2_outputs(12143) <= not(layer1_outputs(1803));
    layer2_outputs(12144) <= layer1_outputs(2787);
    layer2_outputs(12145) <= not(layer1_outputs(4609));
    layer2_outputs(12146) <= not(layer1_outputs(6562));
    layer2_outputs(12147) <= not(layer1_outputs(6248)) or (layer1_outputs(1607));
    layer2_outputs(12148) <= not((layer1_outputs(6862)) and (layer1_outputs(7401)));
    layer2_outputs(12149) <= layer1_outputs(2144);
    layer2_outputs(12150) <= layer1_outputs(6867);
    layer2_outputs(12151) <= layer1_outputs(2742);
    layer2_outputs(12152) <= not(layer1_outputs(10639));
    layer2_outputs(12153) <= not(layer1_outputs(11719)) or (layer1_outputs(4268));
    layer2_outputs(12154) <= layer1_outputs(11391);
    layer2_outputs(12155) <= layer1_outputs(3638);
    layer2_outputs(12156) <= (layer1_outputs(9731)) and (layer1_outputs(8905));
    layer2_outputs(12157) <= layer1_outputs(7034);
    layer2_outputs(12158) <= not((layer1_outputs(4105)) xor (layer1_outputs(12581)));
    layer2_outputs(12159) <= (layer1_outputs(5190)) and (layer1_outputs(8303));
    layer2_outputs(12160) <= not((layer1_outputs(5598)) or (layer1_outputs(7756)));
    layer2_outputs(12161) <= not(layer1_outputs(211)) or (layer1_outputs(5312));
    layer2_outputs(12162) <= (layer1_outputs(6734)) xor (layer1_outputs(10516));
    layer2_outputs(12163) <= (layer1_outputs(4483)) and (layer1_outputs(4931));
    layer2_outputs(12164) <= (layer1_outputs(358)) and not (layer1_outputs(8424));
    layer2_outputs(12165) <= layer1_outputs(9794);
    layer2_outputs(12166) <= (layer1_outputs(12062)) and not (layer1_outputs(2868));
    layer2_outputs(12167) <= not(layer1_outputs(5507));
    layer2_outputs(12168) <= not(layer1_outputs(2236)) or (layer1_outputs(474));
    layer2_outputs(12169) <= (layer1_outputs(1631)) and not (layer1_outputs(5165));
    layer2_outputs(12170) <= not((layer1_outputs(2889)) xor (layer1_outputs(6410)));
    layer2_outputs(12171) <= not(layer1_outputs(11191));
    layer2_outputs(12172) <= not(layer1_outputs(11182)) or (layer1_outputs(7364));
    layer2_outputs(12173) <= layer1_outputs(851);
    layer2_outputs(12174) <= layer1_outputs(2484);
    layer2_outputs(12175) <= not(layer1_outputs(5264));
    layer2_outputs(12176) <= not(layer1_outputs(6319));
    layer2_outputs(12177) <= not(layer1_outputs(1162));
    layer2_outputs(12178) <= not(layer1_outputs(8370));
    layer2_outputs(12179) <= not(layer1_outputs(9324));
    layer2_outputs(12180) <= not((layer1_outputs(7246)) or (layer1_outputs(12601)));
    layer2_outputs(12181) <= not((layer1_outputs(7960)) or (layer1_outputs(9245)));
    layer2_outputs(12182) <= (layer1_outputs(1616)) and (layer1_outputs(11542));
    layer2_outputs(12183) <= not(layer1_outputs(9123));
    layer2_outputs(12184) <= (layer1_outputs(10942)) xor (layer1_outputs(10883));
    layer2_outputs(12185) <= not(layer1_outputs(4386));
    layer2_outputs(12186) <= layer1_outputs(7542);
    layer2_outputs(12187) <= layer1_outputs(9369);
    layer2_outputs(12188) <= not(layer1_outputs(2278));
    layer2_outputs(12189) <= layer1_outputs(9468);
    layer2_outputs(12190) <= layer1_outputs(694);
    layer2_outputs(12191) <= layer1_outputs(8561);
    layer2_outputs(12192) <= not(layer1_outputs(6386));
    layer2_outputs(12193) <= not(layer1_outputs(3428)) or (layer1_outputs(12161));
    layer2_outputs(12194) <= not(layer1_outputs(247));
    layer2_outputs(12195) <= (layer1_outputs(8724)) xor (layer1_outputs(7076));
    layer2_outputs(12196) <= layer1_outputs(8843);
    layer2_outputs(12197) <= not(layer1_outputs(8012));
    layer2_outputs(12198) <= layer1_outputs(10247);
    layer2_outputs(12199) <= not(layer1_outputs(10571));
    layer2_outputs(12200) <= (layer1_outputs(7187)) xor (layer1_outputs(5572));
    layer2_outputs(12201) <= not((layer1_outputs(4091)) and (layer1_outputs(10910)));
    layer2_outputs(12202) <= not((layer1_outputs(1137)) xor (layer1_outputs(1562)));
    layer2_outputs(12203) <= (layer1_outputs(7445)) xor (layer1_outputs(6439));
    layer2_outputs(12204) <= not((layer1_outputs(7948)) and (layer1_outputs(611)));
    layer2_outputs(12205) <= not((layer1_outputs(3899)) and (layer1_outputs(2929)));
    layer2_outputs(12206) <= not((layer1_outputs(2492)) or (layer1_outputs(9034)));
    layer2_outputs(12207) <= (layer1_outputs(5205)) and not (layer1_outputs(6171));
    layer2_outputs(12208) <= not(layer1_outputs(5530));
    layer2_outputs(12209) <= not(layer1_outputs(7862));
    layer2_outputs(12210) <= not((layer1_outputs(8886)) xor (layer1_outputs(11461)));
    layer2_outputs(12211) <= layer1_outputs(2743);
    layer2_outputs(12212) <= not(layer1_outputs(7097)) or (layer1_outputs(1912));
    layer2_outputs(12213) <= not(layer1_outputs(2330)) or (layer1_outputs(5448));
    layer2_outputs(12214) <= not(layer1_outputs(11525));
    layer2_outputs(12215) <= layer1_outputs(3427);
    layer2_outputs(12216) <= (layer1_outputs(11465)) xor (layer1_outputs(6297));
    layer2_outputs(12217) <= layer1_outputs(2565);
    layer2_outputs(12218) <= layer1_outputs(3893);
    layer2_outputs(12219) <= layer1_outputs(10254);
    layer2_outputs(12220) <= not((layer1_outputs(12595)) and (layer1_outputs(12063)));
    layer2_outputs(12221) <= not((layer1_outputs(1661)) xor (layer1_outputs(12693)));
    layer2_outputs(12222) <= not(layer1_outputs(11913));
    layer2_outputs(12223) <= not(layer1_outputs(8402));
    layer2_outputs(12224) <= not((layer1_outputs(6861)) and (layer1_outputs(11935)));
    layer2_outputs(12225) <= (layer1_outputs(2544)) and (layer1_outputs(1575));
    layer2_outputs(12226) <= not((layer1_outputs(10763)) or (layer1_outputs(6345)));
    layer2_outputs(12227) <= (layer1_outputs(6409)) xor (layer1_outputs(1833));
    layer2_outputs(12228) <= not(layer1_outputs(10523)) or (layer1_outputs(6846));
    layer2_outputs(12229) <= not(layer1_outputs(835));
    layer2_outputs(12230) <= not(layer1_outputs(5273));
    layer2_outputs(12231) <= (layer1_outputs(12057)) and not (layer1_outputs(3524));
    layer2_outputs(12232) <= not(layer1_outputs(12694)) or (layer1_outputs(6202));
    layer2_outputs(12233) <= not(layer1_outputs(12643)) or (layer1_outputs(6629));
    layer2_outputs(12234) <= not(layer1_outputs(8116));
    layer2_outputs(12235) <= not(layer1_outputs(3522));
    layer2_outputs(12236) <= not((layer1_outputs(4854)) or (layer1_outputs(175)));
    layer2_outputs(12237) <= layer1_outputs(6821);
    layer2_outputs(12238) <= not(layer1_outputs(96));
    layer2_outputs(12239) <= layer1_outputs(5713);
    layer2_outputs(12240) <= layer1_outputs(11691);
    layer2_outputs(12241) <= not(layer1_outputs(271));
    layer2_outputs(12242) <= layer1_outputs(2203);
    layer2_outputs(12243) <= not((layer1_outputs(1043)) xor (layer1_outputs(1435)));
    layer2_outputs(12244) <= (layer1_outputs(7135)) and (layer1_outputs(3571));
    layer2_outputs(12245) <= not((layer1_outputs(585)) and (layer1_outputs(6296)));
    layer2_outputs(12246) <= (layer1_outputs(7125)) xor (layer1_outputs(11844));
    layer2_outputs(12247) <= not(layer1_outputs(2689));
    layer2_outputs(12248) <= not(layer1_outputs(7146)) or (layer1_outputs(8436));
    layer2_outputs(12249) <= not(layer1_outputs(11905));
    layer2_outputs(12250) <= not(layer1_outputs(62));
    layer2_outputs(12251) <= (layer1_outputs(9607)) xor (layer1_outputs(8668));
    layer2_outputs(12252) <= not((layer1_outputs(10124)) xor (layer1_outputs(8191)));
    layer2_outputs(12253) <= not((layer1_outputs(1749)) and (layer1_outputs(171)));
    layer2_outputs(12254) <= (layer1_outputs(10439)) xor (layer1_outputs(4225));
    layer2_outputs(12255) <= layer1_outputs(11099);
    layer2_outputs(12256) <= not((layer1_outputs(3897)) xor (layer1_outputs(12557)));
    layer2_outputs(12257) <= (layer1_outputs(639)) and (layer1_outputs(9899));
    layer2_outputs(12258) <= layer1_outputs(7974);
    layer2_outputs(12259) <= not((layer1_outputs(8699)) or (layer1_outputs(5420)));
    layer2_outputs(12260) <= not((layer1_outputs(1613)) or (layer1_outputs(6498)));
    layer2_outputs(12261) <= (layer1_outputs(813)) and not (layer1_outputs(12340));
    layer2_outputs(12262) <= (layer1_outputs(3497)) or (layer1_outputs(1198));
    layer2_outputs(12263) <= layer1_outputs(6165);
    layer2_outputs(12264) <= not(layer1_outputs(5279));
    layer2_outputs(12265) <= not(layer1_outputs(2275));
    layer2_outputs(12266) <= not(layer1_outputs(5995));
    layer2_outputs(12267) <= layer1_outputs(11190);
    layer2_outputs(12268) <= not(layer1_outputs(4295));
    layer2_outputs(12269) <= (layer1_outputs(1532)) xor (layer1_outputs(7543));
    layer2_outputs(12270) <= not(layer1_outputs(5495));
    layer2_outputs(12271) <= not((layer1_outputs(11136)) and (layer1_outputs(3715)));
    layer2_outputs(12272) <= (layer1_outputs(5489)) and (layer1_outputs(5583));
    layer2_outputs(12273) <= not((layer1_outputs(11749)) or (layer1_outputs(5791)));
    layer2_outputs(12274) <= (layer1_outputs(2976)) or (layer1_outputs(2981));
    layer2_outputs(12275) <= layer1_outputs(9038);
    layer2_outputs(12276) <= not(layer1_outputs(5911));
    layer2_outputs(12277) <= not(layer1_outputs(5382)) or (layer1_outputs(9602));
    layer2_outputs(12278) <= not(layer1_outputs(5441)) or (layer1_outputs(7846));
    layer2_outputs(12279) <= layer1_outputs(1080);
    layer2_outputs(12280) <= not((layer1_outputs(8661)) xor (layer1_outputs(4790)));
    layer2_outputs(12281) <= layer1_outputs(809);
    layer2_outputs(12282) <= (layer1_outputs(11311)) xor (layer1_outputs(8491));
    layer2_outputs(12283) <= not(layer1_outputs(7477)) or (layer1_outputs(3297));
    layer2_outputs(12284) <= not(layer1_outputs(8121));
    layer2_outputs(12285) <= not((layer1_outputs(340)) xor (layer1_outputs(3548)));
    layer2_outputs(12286) <= (layer1_outputs(12035)) xor (layer1_outputs(9861));
    layer2_outputs(12287) <= not(layer1_outputs(5603));
    layer2_outputs(12288) <= layer1_outputs(9674);
    layer2_outputs(12289) <= (layer1_outputs(6469)) and not (layer1_outputs(5761));
    layer2_outputs(12290) <= layer1_outputs(11811);
    layer2_outputs(12291) <= not(layer1_outputs(3208));
    layer2_outputs(12292) <= not(layer1_outputs(7671));
    layer2_outputs(12293) <= not(layer1_outputs(93));
    layer2_outputs(12294) <= (layer1_outputs(2618)) xor (layer1_outputs(4830));
    layer2_outputs(12295) <= layer1_outputs(9231);
    layer2_outputs(12296) <= not(layer1_outputs(12683)) or (layer1_outputs(3093));
    layer2_outputs(12297) <= not((layer1_outputs(8643)) and (layer1_outputs(2170)));
    layer2_outputs(12298) <= not(layer1_outputs(8930));
    layer2_outputs(12299) <= (layer1_outputs(5453)) xor (layer1_outputs(10388));
    layer2_outputs(12300) <= not((layer1_outputs(9619)) xor (layer1_outputs(5918)));
    layer2_outputs(12301) <= not(layer1_outputs(9531));
    layer2_outputs(12302) <= (layer1_outputs(9836)) or (layer1_outputs(4325));
    layer2_outputs(12303) <= not(layer1_outputs(11268));
    layer2_outputs(12304) <= layer1_outputs(11430);
    layer2_outputs(12305) <= (layer1_outputs(9110)) xor (layer1_outputs(5277));
    layer2_outputs(12306) <= layer1_outputs(2785);
    layer2_outputs(12307) <= layer1_outputs(3280);
    layer2_outputs(12308) <= not((layer1_outputs(4767)) xor (layer1_outputs(2189)));
    layer2_outputs(12309) <= layer1_outputs(3532);
    layer2_outputs(12310) <= (layer1_outputs(4177)) xor (layer1_outputs(11663));
    layer2_outputs(12311) <= not(layer1_outputs(5952)) or (layer1_outputs(2851));
    layer2_outputs(12312) <= not(layer1_outputs(6520));
    layer2_outputs(12313) <= layer1_outputs(1837);
    layer2_outputs(12314) <= not((layer1_outputs(4428)) xor (layer1_outputs(2216)));
    layer2_outputs(12315) <= layer1_outputs(11843);
    layer2_outputs(12316) <= not(layer1_outputs(7579));
    layer2_outputs(12317) <= not(layer1_outputs(2378));
    layer2_outputs(12318) <= '1';
    layer2_outputs(12319) <= not(layer1_outputs(10029)) or (layer1_outputs(1437));
    layer2_outputs(12320) <= not((layer1_outputs(3902)) xor (layer1_outputs(1629)));
    layer2_outputs(12321) <= (layer1_outputs(11376)) xor (layer1_outputs(5783));
    layer2_outputs(12322) <= layer1_outputs(3337);
    layer2_outputs(12323) <= not(layer1_outputs(12475)) or (layer1_outputs(206));
    layer2_outputs(12324) <= not((layer1_outputs(6544)) or (layer1_outputs(5498)));
    layer2_outputs(12325) <= (layer1_outputs(11193)) and (layer1_outputs(2293));
    layer2_outputs(12326) <= '1';
    layer2_outputs(12327) <= layer1_outputs(7936);
    layer2_outputs(12328) <= not((layer1_outputs(12492)) or (layer1_outputs(2463)));
    layer2_outputs(12329) <= not(layer1_outputs(9729));
    layer2_outputs(12330) <= not(layer1_outputs(3812));
    layer2_outputs(12331) <= (layer1_outputs(1341)) xor (layer1_outputs(12527));
    layer2_outputs(12332) <= layer1_outputs(10195);
    layer2_outputs(12333) <= layer1_outputs(11694);
    layer2_outputs(12334) <= (layer1_outputs(9225)) and not (layer1_outputs(10479));
    layer2_outputs(12335) <= not(layer1_outputs(8662));
    layer2_outputs(12336) <= layer1_outputs(5953);
    layer2_outputs(12337) <= layer1_outputs(15);
    layer2_outputs(12338) <= layer1_outputs(1795);
    layer2_outputs(12339) <= (layer1_outputs(8019)) or (layer1_outputs(3868));
    layer2_outputs(12340) <= (layer1_outputs(300)) and (layer1_outputs(8235));
    layer2_outputs(12341) <= layer1_outputs(12523);
    layer2_outputs(12342) <= not((layer1_outputs(8689)) xor (layer1_outputs(8202)));
    layer2_outputs(12343) <= not(layer1_outputs(6683)) or (layer1_outputs(3009));
    layer2_outputs(12344) <= layer1_outputs(1404);
    layer2_outputs(12345) <= layer1_outputs(8);
    layer2_outputs(12346) <= not(layer1_outputs(12313)) or (layer1_outputs(2937));
    layer2_outputs(12347) <= not(layer1_outputs(2837));
    layer2_outputs(12348) <= (layer1_outputs(11174)) xor (layer1_outputs(4589));
    layer2_outputs(12349) <= layer1_outputs(1541);
    layer2_outputs(12350) <= not((layer1_outputs(6736)) or (layer1_outputs(1411)));
    layer2_outputs(12351) <= layer1_outputs(6450);
    layer2_outputs(12352) <= '1';
    layer2_outputs(12353) <= layer1_outputs(11384);
    layer2_outputs(12354) <= layer1_outputs(4706);
    layer2_outputs(12355) <= (layer1_outputs(7229)) xor (layer1_outputs(11949));
    layer2_outputs(12356) <= (layer1_outputs(12645)) xor (layer1_outputs(8624));
    layer2_outputs(12357) <= layer1_outputs(4696);
    layer2_outputs(12358) <= (layer1_outputs(9484)) and not (layer1_outputs(7218));
    layer2_outputs(12359) <= (layer1_outputs(1455)) and not (layer1_outputs(279));
    layer2_outputs(12360) <= not(layer1_outputs(6313)) or (layer1_outputs(3036));
    layer2_outputs(12361) <= not(layer1_outputs(4970)) or (layer1_outputs(4984));
    layer2_outputs(12362) <= (layer1_outputs(9222)) and (layer1_outputs(11799));
    layer2_outputs(12363) <= not(layer1_outputs(9247)) or (layer1_outputs(11340));
    layer2_outputs(12364) <= not(layer1_outputs(2018));
    layer2_outputs(12365) <= layer1_outputs(11284);
    layer2_outputs(12366) <= (layer1_outputs(3001)) xor (layer1_outputs(10101));
    layer2_outputs(12367) <= layer1_outputs(11323);
    layer2_outputs(12368) <= not(layer1_outputs(5699));
    layer2_outputs(12369) <= not((layer1_outputs(6001)) or (layer1_outputs(488)));
    layer2_outputs(12370) <= not(layer1_outputs(7207)) or (layer1_outputs(3672));
    layer2_outputs(12371) <= (layer1_outputs(752)) xor (layer1_outputs(12181));
    layer2_outputs(12372) <= layer1_outputs(10200);
    layer2_outputs(12373) <= not(layer1_outputs(10281));
    layer2_outputs(12374) <= not(layer1_outputs(12084)) or (layer1_outputs(7917));
    layer2_outputs(12375) <= not((layer1_outputs(7078)) or (layer1_outputs(6331)));
    layer2_outputs(12376) <= not(layer1_outputs(3033));
    layer2_outputs(12377) <= not(layer1_outputs(3282));
    layer2_outputs(12378) <= '1';
    layer2_outputs(12379) <= layer1_outputs(2898);
    layer2_outputs(12380) <= not((layer1_outputs(3116)) xor (layer1_outputs(1495)));
    layer2_outputs(12381) <= layer1_outputs(5648);
    layer2_outputs(12382) <= not(layer1_outputs(1282));
    layer2_outputs(12383) <= not(layer1_outputs(11658)) or (layer1_outputs(7458));
    layer2_outputs(12384) <= (layer1_outputs(1273)) and not (layer1_outputs(92));
    layer2_outputs(12385) <= (layer1_outputs(3109)) xor (layer1_outputs(6785));
    layer2_outputs(12386) <= layer1_outputs(2486);
    layer2_outputs(12387) <= (layer1_outputs(3261)) and not (layer1_outputs(8227));
    layer2_outputs(12388) <= not(layer1_outputs(2357));
    layer2_outputs(12389) <= not(layer1_outputs(3979)) or (layer1_outputs(10238));
    layer2_outputs(12390) <= (layer1_outputs(5061)) and not (layer1_outputs(2295));
    layer2_outputs(12391) <= layer1_outputs(3556);
    layer2_outputs(12392) <= not(layer1_outputs(10579)) or (layer1_outputs(4412));
    layer2_outputs(12393) <= (layer1_outputs(10523)) and not (layer1_outputs(12545));
    layer2_outputs(12394) <= not(layer1_outputs(4233));
    layer2_outputs(12395) <= not(layer1_outputs(1893));
    layer2_outputs(12396) <= (layer1_outputs(8493)) xor (layer1_outputs(816));
    layer2_outputs(12397) <= not(layer1_outputs(1790));
    layer2_outputs(12398) <= (layer1_outputs(6118)) xor (layer1_outputs(5124));
    layer2_outputs(12399) <= not(layer1_outputs(8916));
    layer2_outputs(12400) <= not(layer1_outputs(2992));
    layer2_outputs(12401) <= not(layer1_outputs(3816));
    layer2_outputs(12402) <= not(layer1_outputs(9365));
    layer2_outputs(12403) <= (layer1_outputs(4822)) and not (layer1_outputs(4646));
    layer2_outputs(12404) <= not((layer1_outputs(12764)) or (layer1_outputs(686)));
    layer2_outputs(12405) <= not((layer1_outputs(7999)) xor (layer1_outputs(8832)));
    layer2_outputs(12406) <= (layer1_outputs(7909)) or (layer1_outputs(8880));
    layer2_outputs(12407) <= not(layer1_outputs(2886));
    layer2_outputs(12408) <= layer1_outputs(4135);
    layer2_outputs(12409) <= (layer1_outputs(547)) or (layer1_outputs(8667));
    layer2_outputs(12410) <= not(layer1_outputs(4819)) or (layer1_outputs(3381));
    layer2_outputs(12411) <= not((layer1_outputs(7338)) or (layer1_outputs(11392)));
    layer2_outputs(12412) <= (layer1_outputs(632)) and (layer1_outputs(7561));
    layer2_outputs(12413) <= layer1_outputs(10426);
    layer2_outputs(12414) <= layer1_outputs(6606);
    layer2_outputs(12415) <= layer1_outputs(908);
    layer2_outputs(12416) <= not(layer1_outputs(9021)) or (layer1_outputs(7765));
    layer2_outputs(12417) <= not((layer1_outputs(3872)) xor (layer1_outputs(2487)));
    layer2_outputs(12418) <= (layer1_outputs(11862)) and not (layer1_outputs(6393));
    layer2_outputs(12419) <= not(layer1_outputs(7182));
    layer2_outputs(12420) <= not((layer1_outputs(6263)) or (layer1_outputs(10732)));
    layer2_outputs(12421) <= layer1_outputs(7740);
    layer2_outputs(12422) <= layer1_outputs(11775);
    layer2_outputs(12423) <= '1';
    layer2_outputs(12424) <= not(layer1_outputs(1958));
    layer2_outputs(12425) <= layer1_outputs(7567);
    layer2_outputs(12426) <= not(layer1_outputs(12479)) or (layer1_outputs(1035));
    layer2_outputs(12427) <= (layer1_outputs(5096)) and not (layer1_outputs(1363));
    layer2_outputs(12428) <= not(layer1_outputs(6479));
    layer2_outputs(12429) <= not(layer1_outputs(9693)) or (layer1_outputs(5904));
    layer2_outputs(12430) <= not(layer1_outputs(3249)) or (layer1_outputs(7716));
    layer2_outputs(12431) <= not((layer1_outputs(3535)) xor (layer1_outputs(12666)));
    layer2_outputs(12432) <= not(layer1_outputs(139)) or (layer1_outputs(3998));
    layer2_outputs(12433) <= not((layer1_outputs(8733)) xor (layer1_outputs(10984)));
    layer2_outputs(12434) <= layer1_outputs(1765);
    layer2_outputs(12435) <= not(layer1_outputs(2295));
    layer2_outputs(12436) <= not((layer1_outputs(1066)) xor (layer1_outputs(4745)));
    layer2_outputs(12437) <= layer1_outputs(10642);
    layer2_outputs(12438) <= not(layer1_outputs(53));
    layer2_outputs(12439) <= not((layer1_outputs(8545)) xor (layer1_outputs(2202)));
    layer2_outputs(12440) <= not(layer1_outputs(880)) or (layer1_outputs(5558));
    layer2_outputs(12441) <= not((layer1_outputs(2371)) or (layer1_outputs(2001)));
    layer2_outputs(12442) <= (layer1_outputs(4023)) and not (layer1_outputs(4594));
    layer2_outputs(12443) <= (layer1_outputs(6026)) and (layer1_outputs(8221));
    layer2_outputs(12444) <= layer1_outputs(7853);
    layer2_outputs(12445) <= not(layer1_outputs(11742)) or (layer1_outputs(8426));
    layer2_outputs(12446) <= layer1_outputs(1462);
    layer2_outputs(12447) <= layer1_outputs(3079);
    layer2_outputs(12448) <= (layer1_outputs(12267)) xor (layer1_outputs(2600));
    layer2_outputs(12449) <= not((layer1_outputs(7376)) and (layer1_outputs(4894)));
    layer2_outputs(12450) <= (layer1_outputs(1648)) and not (layer1_outputs(7556));
    layer2_outputs(12451) <= not(layer1_outputs(7717));
    layer2_outputs(12452) <= (layer1_outputs(7575)) and (layer1_outputs(5249));
    layer2_outputs(12453) <= layer1_outputs(7431);
    layer2_outputs(12454) <= not((layer1_outputs(8981)) xor (layer1_outputs(7569)));
    layer2_outputs(12455) <= not(layer1_outputs(12643));
    layer2_outputs(12456) <= not(layer1_outputs(3493)) or (layer1_outputs(831));
    layer2_outputs(12457) <= (layer1_outputs(6798)) xor (layer1_outputs(2803));
    layer2_outputs(12458) <= not((layer1_outputs(5560)) xor (layer1_outputs(11812)));
    layer2_outputs(12459) <= layer1_outputs(10497);
    layer2_outputs(12460) <= layer1_outputs(10324);
    layer2_outputs(12461) <= (layer1_outputs(4139)) and not (layer1_outputs(3895));
    layer2_outputs(12462) <= layer1_outputs(9777);
    layer2_outputs(12463) <= (layer1_outputs(5114)) xor (layer1_outputs(7181));
    layer2_outputs(12464) <= not((layer1_outputs(3321)) xor (layer1_outputs(3480)));
    layer2_outputs(12465) <= '0';
    layer2_outputs(12466) <= not(layer1_outputs(4481));
    layer2_outputs(12467) <= (layer1_outputs(7260)) and (layer1_outputs(7696));
    layer2_outputs(12468) <= (layer1_outputs(9415)) or (layer1_outputs(1928));
    layer2_outputs(12469) <= not(layer1_outputs(1638));
    layer2_outputs(12470) <= not((layer1_outputs(6256)) and (layer1_outputs(9760)));
    layer2_outputs(12471) <= not(layer1_outputs(2367));
    layer2_outputs(12472) <= layer1_outputs(7644);
    layer2_outputs(12473) <= not(layer1_outputs(2271)) or (layer1_outputs(10360));
    layer2_outputs(12474) <= layer1_outputs(10654);
    layer2_outputs(12475) <= layer1_outputs(4882);
    layer2_outputs(12476) <= not(layer1_outputs(1138));
    layer2_outputs(12477) <= layer1_outputs(6768);
    layer2_outputs(12478) <= not(layer1_outputs(10461)) or (layer1_outputs(12101));
    layer2_outputs(12479) <= (layer1_outputs(6241)) and not (layer1_outputs(7589));
    layer2_outputs(12480) <= not(layer1_outputs(2642)) or (layer1_outputs(6181));
    layer2_outputs(12481) <= not((layer1_outputs(5933)) xor (layer1_outputs(11220)));
    layer2_outputs(12482) <= (layer1_outputs(7326)) and not (layer1_outputs(7916));
    layer2_outputs(12483) <= layer1_outputs(3136);
    layer2_outputs(12484) <= not(layer1_outputs(11910));
    layer2_outputs(12485) <= layer1_outputs(3431);
    layer2_outputs(12486) <= layer1_outputs(5541);
    layer2_outputs(12487) <= (layer1_outputs(3332)) and (layer1_outputs(3100));
    layer2_outputs(12488) <= not(layer1_outputs(8054)) or (layer1_outputs(459));
    layer2_outputs(12489) <= not((layer1_outputs(2306)) or (layer1_outputs(679)));
    layer2_outputs(12490) <= layer1_outputs(7672);
    layer2_outputs(12491) <= (layer1_outputs(5344)) and not (layer1_outputs(8219));
    layer2_outputs(12492) <= (layer1_outputs(540)) and not (layer1_outputs(5626));
    layer2_outputs(12493) <= layer1_outputs(1133);
    layer2_outputs(12494) <= layer1_outputs(12746);
    layer2_outputs(12495) <= not(layer1_outputs(4982));
    layer2_outputs(12496) <= (layer1_outputs(384)) and not (layer1_outputs(1868));
    layer2_outputs(12497) <= not(layer1_outputs(11120));
    layer2_outputs(12498) <= (layer1_outputs(844)) or (layer1_outputs(9769));
    layer2_outputs(12499) <= not((layer1_outputs(2333)) and (layer1_outputs(10357)));
    layer2_outputs(12500) <= not(layer1_outputs(1112)) or (layer1_outputs(11409));
    layer2_outputs(12501) <= (layer1_outputs(2977)) xor (layer1_outputs(4062));
    layer2_outputs(12502) <= (layer1_outputs(11394)) and (layer1_outputs(10860));
    layer2_outputs(12503) <= (layer1_outputs(2369)) and not (layer1_outputs(3323));
    layer2_outputs(12504) <= not(layer1_outputs(10564));
    layer2_outputs(12505) <= layer1_outputs(1847);
    layer2_outputs(12506) <= not((layer1_outputs(2599)) and (layer1_outputs(1898)));
    layer2_outputs(12507) <= not(layer1_outputs(4391));
    layer2_outputs(12508) <= not(layer1_outputs(7499)) or (layer1_outputs(2860));
    layer2_outputs(12509) <= layer1_outputs(8046);
    layer2_outputs(12510) <= not((layer1_outputs(7557)) and (layer1_outputs(4863)));
    layer2_outputs(12511) <= not((layer1_outputs(1028)) xor (layer1_outputs(9444)));
    layer2_outputs(12512) <= (layer1_outputs(1849)) and not (layer1_outputs(11090));
    layer2_outputs(12513) <= not(layer1_outputs(6933)) or (layer1_outputs(4344));
    layer2_outputs(12514) <= (layer1_outputs(12013)) xor (layer1_outputs(11172));
    layer2_outputs(12515) <= layer1_outputs(1739);
    layer2_outputs(12516) <= not(layer1_outputs(3006));
    layer2_outputs(12517) <= not((layer1_outputs(12094)) and (layer1_outputs(7615)));
    layer2_outputs(12518) <= layer1_outputs(5108);
    layer2_outputs(12519) <= layer1_outputs(11330);
    layer2_outputs(12520) <= not((layer1_outputs(3032)) and (layer1_outputs(4613)));
    layer2_outputs(12521) <= (layer1_outputs(3821)) and not (layer1_outputs(3836));
    layer2_outputs(12522) <= not(layer1_outputs(7953)) or (layer1_outputs(5856));
    layer2_outputs(12523) <= not(layer1_outputs(5812));
    layer2_outputs(12524) <= layer1_outputs(11189);
    layer2_outputs(12525) <= layer1_outputs(2953);
    layer2_outputs(12526) <= not(layer1_outputs(9054)) or (layer1_outputs(396));
    layer2_outputs(12527) <= not(layer1_outputs(8437));
    layer2_outputs(12528) <= not(layer1_outputs(5586)) or (layer1_outputs(2387));
    layer2_outputs(12529) <= layer1_outputs(989);
    layer2_outputs(12530) <= not(layer1_outputs(8957));
    layer2_outputs(12531) <= (layer1_outputs(10799)) or (layer1_outputs(9126));
    layer2_outputs(12532) <= not((layer1_outputs(6761)) or (layer1_outputs(8588)));
    layer2_outputs(12533) <= (layer1_outputs(11669)) and (layer1_outputs(6485));
    layer2_outputs(12534) <= not((layer1_outputs(2984)) and (layer1_outputs(9532)));
    layer2_outputs(12535) <= (layer1_outputs(108)) xor (layer1_outputs(8124));
    layer2_outputs(12536) <= (layer1_outputs(11951)) or (layer1_outputs(12179));
    layer2_outputs(12537) <= not((layer1_outputs(2918)) or (layer1_outputs(6461)));
    layer2_outputs(12538) <= layer1_outputs(12004);
    layer2_outputs(12539) <= not(layer1_outputs(10873)) or (layer1_outputs(5036));
    layer2_outputs(12540) <= (layer1_outputs(11876)) xor (layer1_outputs(9253));
    layer2_outputs(12541) <= (layer1_outputs(11663)) or (layer1_outputs(3659));
    layer2_outputs(12542) <= not(layer1_outputs(8268));
    layer2_outputs(12543) <= not(layer1_outputs(5210));
    layer2_outputs(12544) <= not(layer1_outputs(3943));
    layer2_outputs(12545) <= not((layer1_outputs(12575)) or (layer1_outputs(3172)));
    layer2_outputs(12546) <= (layer1_outputs(3148)) xor (layer1_outputs(3856));
    layer2_outputs(12547) <= not(layer1_outputs(6289));
    layer2_outputs(12548) <= (layer1_outputs(10973)) and not (layer1_outputs(7968));
    layer2_outputs(12549) <= layer1_outputs(2495);
    layer2_outputs(12550) <= not(layer1_outputs(1981)) or (layer1_outputs(1426));
    layer2_outputs(12551) <= layer1_outputs(12390);
    layer2_outputs(12552) <= not(layer1_outputs(12005));
    layer2_outputs(12553) <= not(layer1_outputs(12312));
    layer2_outputs(12554) <= not(layer1_outputs(10758)) or (layer1_outputs(7829));
    layer2_outputs(12555) <= layer1_outputs(8478);
    layer2_outputs(12556) <= not(layer1_outputs(10228));
    layer2_outputs(12557) <= not(layer1_outputs(8860));
    layer2_outputs(12558) <= (layer1_outputs(3959)) and not (layer1_outputs(951));
    layer2_outputs(12559) <= not((layer1_outputs(7303)) xor (layer1_outputs(6908)));
    layer2_outputs(12560) <= not((layer1_outputs(3251)) and (layer1_outputs(878)));
    layer2_outputs(12561) <= (layer1_outputs(11133)) and (layer1_outputs(12220));
    layer2_outputs(12562) <= (layer1_outputs(288)) or (layer1_outputs(9934));
    layer2_outputs(12563) <= layer1_outputs(10185);
    layer2_outputs(12564) <= (layer1_outputs(6543)) xor (layer1_outputs(232));
    layer2_outputs(12565) <= layer1_outputs(9604);
    layer2_outputs(12566) <= not(layer1_outputs(12634));
    layer2_outputs(12567) <= (layer1_outputs(10537)) and not (layer1_outputs(11327));
    layer2_outputs(12568) <= layer1_outputs(469);
    layer2_outputs(12569) <= (layer1_outputs(1062)) or (layer1_outputs(5406));
    layer2_outputs(12570) <= not((layer1_outputs(2385)) xor (layer1_outputs(9246)));
    layer2_outputs(12571) <= layer1_outputs(735);
    layer2_outputs(12572) <= not(layer1_outputs(11917));
    layer2_outputs(12573) <= (layer1_outputs(872)) and not (layer1_outputs(6977));
    layer2_outputs(12574) <= not(layer1_outputs(11368));
    layer2_outputs(12575) <= not(layer1_outputs(1085));
    layer2_outputs(12576) <= not((layer1_outputs(383)) and (layer1_outputs(4436)));
    layer2_outputs(12577) <= (layer1_outputs(3120)) and not (layer1_outputs(1986));
    layer2_outputs(12578) <= layer1_outputs(3926);
    layer2_outputs(12579) <= not((layer1_outputs(9085)) and (layer1_outputs(12265)));
    layer2_outputs(12580) <= not((layer1_outputs(7942)) and (layer1_outputs(10188)));
    layer2_outputs(12581) <= (layer1_outputs(11237)) xor (layer1_outputs(1960));
    layer2_outputs(12582) <= not(layer1_outputs(7652));
    layer2_outputs(12583) <= (layer1_outputs(10851)) xor (layer1_outputs(2005));
    layer2_outputs(12584) <= layer1_outputs(10087);
    layer2_outputs(12585) <= not(layer1_outputs(6284));
    layer2_outputs(12586) <= not((layer1_outputs(9457)) and (layer1_outputs(6250)));
    layer2_outputs(12587) <= not(layer1_outputs(9331));
    layer2_outputs(12588) <= not(layer1_outputs(9737));
    layer2_outputs(12589) <= layer1_outputs(3542);
    layer2_outputs(12590) <= (layer1_outputs(1086)) and not (layer1_outputs(10995));
    layer2_outputs(12591) <= not((layer1_outputs(4972)) xor (layer1_outputs(9554)));
    layer2_outputs(12592) <= not(layer1_outputs(7890));
    layer2_outputs(12593) <= not(layer1_outputs(8799));
    layer2_outputs(12594) <= not(layer1_outputs(7814));
    layer2_outputs(12595) <= (layer1_outputs(463)) xor (layer1_outputs(11715));
    layer2_outputs(12596) <= (layer1_outputs(11601)) and not (layer1_outputs(9342));
    layer2_outputs(12597) <= not(layer1_outputs(9764));
    layer2_outputs(12598) <= layer1_outputs(5586);
    layer2_outputs(12599) <= not((layer1_outputs(7982)) xor (layer1_outputs(1106)));
    layer2_outputs(12600) <= not((layer1_outputs(3630)) and (layer1_outputs(8505)));
    layer2_outputs(12601) <= (layer1_outputs(569)) and (layer1_outputs(2169));
    layer2_outputs(12602) <= (layer1_outputs(2532)) xor (layer1_outputs(12113));
    layer2_outputs(12603) <= (layer1_outputs(647)) and not (layer1_outputs(7788));
    layer2_outputs(12604) <= not(layer1_outputs(11622));
    layer2_outputs(12605) <= layer1_outputs(4781);
    layer2_outputs(12606) <= (layer1_outputs(6412)) xor (layer1_outputs(2234));
    layer2_outputs(12607) <= (layer1_outputs(5170)) xor (layer1_outputs(12247));
    layer2_outputs(12608) <= layer1_outputs(2184);
    layer2_outputs(12609) <= not((layer1_outputs(9993)) xor (layer1_outputs(816)));
    layer2_outputs(12610) <= not(layer1_outputs(8594));
    layer2_outputs(12611) <= layer1_outputs(1082);
    layer2_outputs(12612) <= layer1_outputs(1239);
    layer2_outputs(12613) <= layer1_outputs(12727);
    layer2_outputs(12614) <= layer1_outputs(5948);
    layer2_outputs(12615) <= layer1_outputs(804);
    layer2_outputs(12616) <= not(layer1_outputs(4874));
    layer2_outputs(12617) <= not(layer1_outputs(9183));
    layer2_outputs(12618) <= layer1_outputs(5379);
    layer2_outputs(12619) <= not(layer1_outputs(9942)) or (layer1_outputs(2679));
    layer2_outputs(12620) <= (layer1_outputs(2606)) and not (layer1_outputs(48));
    layer2_outputs(12621) <= not(layer1_outputs(10349));
    layer2_outputs(12622) <= layer1_outputs(11123);
    layer2_outputs(12623) <= (layer1_outputs(4842)) xor (layer1_outputs(11772));
    layer2_outputs(12624) <= layer1_outputs(1402);
    layer2_outputs(12625) <= (layer1_outputs(1888)) xor (layer1_outputs(12598));
    layer2_outputs(12626) <= (layer1_outputs(230)) and not (layer1_outputs(3702));
    layer2_outputs(12627) <= not((layer1_outputs(9160)) xor (layer1_outputs(9751)));
    layer2_outputs(12628) <= layer1_outputs(4335);
    layer2_outputs(12629) <= layer1_outputs(11739);
    layer2_outputs(12630) <= not((layer1_outputs(10994)) xor (layer1_outputs(12063)));
    layer2_outputs(12631) <= not(layer1_outputs(6674)) or (layer1_outputs(2571));
    layer2_outputs(12632) <= not(layer1_outputs(5788));
    layer2_outputs(12633) <= not((layer1_outputs(348)) xor (layer1_outputs(4778)));
    layer2_outputs(12634) <= layer1_outputs(9471);
    layer2_outputs(12635) <= '0';
    layer2_outputs(12636) <= (layer1_outputs(4171)) and not (layer1_outputs(2763));
    layer2_outputs(12637) <= not(layer1_outputs(3044));
    layer2_outputs(12638) <= (layer1_outputs(9144)) and (layer1_outputs(4716));
    layer2_outputs(12639) <= not(layer1_outputs(230));
    layer2_outputs(12640) <= not(layer1_outputs(5049)) or (layer1_outputs(11959));
    layer2_outputs(12641) <= layer1_outputs(5739);
    layer2_outputs(12642) <= '1';
    layer2_outputs(12643) <= not(layer1_outputs(1455)) or (layer1_outputs(3789));
    layer2_outputs(12644) <= not(layer1_outputs(11812));
    layer2_outputs(12645) <= not((layer1_outputs(6094)) and (layer1_outputs(4678)));
    layer2_outputs(12646) <= not((layer1_outputs(11355)) and (layer1_outputs(6502)));
    layer2_outputs(12647) <= (layer1_outputs(6139)) and (layer1_outputs(11528));
    layer2_outputs(12648) <= layer1_outputs(6503);
    layer2_outputs(12649) <= not(layer1_outputs(6154));
    layer2_outputs(12650) <= (layer1_outputs(12567)) and not (layer1_outputs(475));
    layer2_outputs(12651) <= (layer1_outputs(10839)) xor (layer1_outputs(4087));
    layer2_outputs(12652) <= (layer1_outputs(5303)) xor (layer1_outputs(7207));
    layer2_outputs(12653) <= not(layer1_outputs(2966)) or (layer1_outputs(10526));
    layer2_outputs(12654) <= (layer1_outputs(5851)) or (layer1_outputs(5231));
    layer2_outputs(12655) <= not(layer1_outputs(478)) or (layer1_outputs(10107));
    layer2_outputs(12656) <= not((layer1_outputs(1521)) xor (layer1_outputs(10809)));
    layer2_outputs(12657) <= (layer1_outputs(8376)) or (layer1_outputs(673));
    layer2_outputs(12658) <= layer1_outputs(6263);
    layer2_outputs(12659) <= (layer1_outputs(9018)) and not (layer1_outputs(9574));
    layer2_outputs(12660) <= not(layer1_outputs(3911)) or (layer1_outputs(7368));
    layer2_outputs(12661) <= not((layer1_outputs(1431)) or (layer1_outputs(5613)));
    layer2_outputs(12662) <= not(layer1_outputs(2240));
    layer2_outputs(12663) <= not((layer1_outputs(5154)) or (layer1_outputs(11147)));
    layer2_outputs(12664) <= (layer1_outputs(3571)) xor (layer1_outputs(2208));
    layer2_outputs(12665) <= not(layer1_outputs(8249)) or (layer1_outputs(8403));
    layer2_outputs(12666) <= not((layer1_outputs(2891)) or (layer1_outputs(6602)));
    layer2_outputs(12667) <= layer1_outputs(9312);
    layer2_outputs(12668) <= layer1_outputs(4202);
    layer2_outputs(12669) <= (layer1_outputs(2466)) and (layer1_outputs(2991));
    layer2_outputs(12670) <= not(layer1_outputs(5035));
    layer2_outputs(12671) <= (layer1_outputs(9493)) xor (layer1_outputs(10164));
    layer2_outputs(12672) <= (layer1_outputs(1654)) and not (layer1_outputs(8575));
    layer2_outputs(12673) <= layer1_outputs(4670);
    layer2_outputs(12674) <= layer1_outputs(685);
    layer2_outputs(12675) <= (layer1_outputs(7186)) xor (layer1_outputs(5576));
    layer2_outputs(12676) <= not((layer1_outputs(3573)) or (layer1_outputs(2680)));
    layer2_outputs(12677) <= layer1_outputs(433);
    layer2_outputs(12678) <= layer1_outputs(12497);
    layer2_outputs(12679) <= not(layer1_outputs(2797)) or (layer1_outputs(11636));
    layer2_outputs(12680) <= (layer1_outputs(1823)) or (layer1_outputs(7343));
    layer2_outputs(12681) <= (layer1_outputs(10257)) and not (layer1_outputs(11486));
    layer2_outputs(12682) <= (layer1_outputs(9079)) and (layer1_outputs(5099));
    layer2_outputs(12683) <= (layer1_outputs(3691)) or (layer1_outputs(10584));
    layer2_outputs(12684) <= (layer1_outputs(1875)) and not (layer1_outputs(3580));
    layer2_outputs(12685) <= not(layer1_outputs(12393));
    layer2_outputs(12686) <= not(layer1_outputs(3591)) or (layer1_outputs(9560));
    layer2_outputs(12687) <= not(layer1_outputs(10458));
    layer2_outputs(12688) <= (layer1_outputs(8240)) xor (layer1_outputs(92));
    layer2_outputs(12689) <= not(layer1_outputs(853));
    layer2_outputs(12690) <= layer1_outputs(10969);
    layer2_outputs(12691) <= not(layer1_outputs(7074));
    layer2_outputs(12692) <= not(layer1_outputs(10340));
    layer2_outputs(12693) <= (layer1_outputs(6912)) or (layer1_outputs(8696));
    layer2_outputs(12694) <= layer1_outputs(12612);
    layer2_outputs(12695) <= layer1_outputs(3334);
    layer2_outputs(12696) <= not((layer1_outputs(6464)) xor (layer1_outputs(3453)));
    layer2_outputs(12697) <= layer1_outputs(10000);
    layer2_outputs(12698) <= layer1_outputs(7479);
    layer2_outputs(12699) <= (layer1_outputs(759)) and (layer1_outputs(3017));
    layer2_outputs(12700) <= '0';
    layer2_outputs(12701) <= (layer1_outputs(11160)) and not (layer1_outputs(6527));
    layer2_outputs(12702) <= not(layer1_outputs(89));
    layer2_outputs(12703) <= (layer1_outputs(11126)) and not (layer1_outputs(4755));
    layer2_outputs(12704) <= '0';
    layer2_outputs(12705) <= layer1_outputs(9867);
    layer2_outputs(12706) <= (layer1_outputs(736)) and (layer1_outputs(4544));
    layer2_outputs(12707) <= (layer1_outputs(11888)) and not (layer1_outputs(3036));
    layer2_outputs(12708) <= layer1_outputs(4776);
    layer2_outputs(12709) <= layer1_outputs(905);
    layer2_outputs(12710) <= layer1_outputs(11671);
    layer2_outputs(12711) <= not(layer1_outputs(11264));
    layer2_outputs(12712) <= (layer1_outputs(8239)) xor (layer1_outputs(4596));
    layer2_outputs(12713) <= layer1_outputs(9889);
    layer2_outputs(12714) <= layer1_outputs(10111);
    layer2_outputs(12715) <= not(layer1_outputs(2008));
    layer2_outputs(12716) <= not(layer1_outputs(7596)) or (layer1_outputs(2981));
    layer2_outputs(12717) <= not((layer1_outputs(227)) and (layer1_outputs(11457)));
    layer2_outputs(12718) <= not(layer1_outputs(7633)) or (layer1_outputs(7247));
    layer2_outputs(12719) <= not((layer1_outputs(11679)) and (layer1_outputs(8599)));
    layer2_outputs(12720) <= not(layer1_outputs(11914));
    layer2_outputs(12721) <= not(layer1_outputs(11073));
    layer2_outputs(12722) <= layer1_outputs(6916);
    layer2_outputs(12723) <= not(layer1_outputs(9142));
    layer2_outputs(12724) <= (layer1_outputs(8544)) and not (layer1_outputs(9025));
    layer2_outputs(12725) <= layer1_outputs(11604);
    layer2_outputs(12726) <= (layer1_outputs(7457)) xor (layer1_outputs(12501));
    layer2_outputs(12727) <= layer1_outputs(6893);
    layer2_outputs(12728) <= layer1_outputs(7150);
    layer2_outputs(12729) <= not(layer1_outputs(6529));
    layer2_outputs(12730) <= layer1_outputs(2206);
    layer2_outputs(12731) <= (layer1_outputs(12192)) xor (layer1_outputs(10633));
    layer2_outputs(12732) <= layer1_outputs(6607);
    layer2_outputs(12733) <= not((layer1_outputs(4108)) or (layer1_outputs(1879)));
    layer2_outputs(12734) <= layer1_outputs(9092);
    layer2_outputs(12735) <= not(layer1_outputs(9496));
    layer2_outputs(12736) <= not(layer1_outputs(1810)) or (layer1_outputs(2985));
    layer2_outputs(12737) <= (layer1_outputs(3008)) xor (layer1_outputs(11465));
    layer2_outputs(12738) <= layer1_outputs(9720);
    layer2_outputs(12739) <= not(layer1_outputs(7956)) or (layer1_outputs(368));
    layer2_outputs(12740) <= (layer1_outputs(10708)) and not (layer1_outputs(8583));
    layer2_outputs(12741) <= (layer1_outputs(1058)) xor (layer1_outputs(5058));
    layer2_outputs(12742) <= (layer1_outputs(4117)) xor (layer1_outputs(4302));
    layer2_outputs(12743) <= not(layer1_outputs(11789));
    layer2_outputs(12744) <= layer1_outputs(9937);
    layer2_outputs(12745) <= layer1_outputs(10247);
    layer2_outputs(12746) <= (layer1_outputs(1540)) and (layer1_outputs(10491));
    layer2_outputs(12747) <= not((layer1_outputs(7085)) xor (layer1_outputs(4323)));
    layer2_outputs(12748) <= not(layer1_outputs(10463)) or (layer1_outputs(9799));
    layer2_outputs(12749) <= not(layer1_outputs(7328));
    layer2_outputs(12750) <= layer1_outputs(1523);
    layer2_outputs(12751) <= '1';
    layer2_outputs(12752) <= layer1_outputs(1473);
    layer2_outputs(12753) <= (layer1_outputs(2046)) and not (layer1_outputs(9091));
    layer2_outputs(12754) <= (layer1_outputs(5976)) xor (layer1_outputs(1921));
    layer2_outputs(12755) <= (layer1_outputs(5662)) and not (layer1_outputs(1304));
    layer2_outputs(12756) <= layer1_outputs(8418);
    layer2_outputs(12757) <= '1';
    layer2_outputs(12758) <= not(layer1_outputs(3105)) or (layer1_outputs(10657));
    layer2_outputs(12759) <= (layer1_outputs(3940)) and not (layer1_outputs(10128));
    layer2_outputs(12760) <= (layer1_outputs(10154)) or (layer1_outputs(4800));
    layer2_outputs(12761) <= (layer1_outputs(9281)) xor (layer1_outputs(903));
    layer2_outputs(12762) <= not(layer1_outputs(1923)) or (layer1_outputs(6944));
    layer2_outputs(12763) <= layer1_outputs(10803);
    layer2_outputs(12764) <= not(layer1_outputs(992));
    layer2_outputs(12765) <= not((layer1_outputs(12543)) or (layer1_outputs(5013)));
    layer2_outputs(12766) <= not(layer1_outputs(1326));
    layer2_outputs(12767) <= layer1_outputs(9060);
    layer2_outputs(12768) <= not((layer1_outputs(10973)) or (layer1_outputs(10812)));
    layer2_outputs(12769) <= layer1_outputs(178);
    layer2_outputs(12770) <= not(layer1_outputs(5458)) or (layer1_outputs(1566));
    layer2_outputs(12771) <= not((layer1_outputs(3628)) or (layer1_outputs(4639)));
    layer2_outputs(12772) <= (layer1_outputs(11229)) xor (layer1_outputs(9773));
    layer2_outputs(12773) <= (layer1_outputs(6620)) or (layer1_outputs(11919));
    layer2_outputs(12774) <= not((layer1_outputs(674)) and (layer1_outputs(1318)));
    layer2_outputs(12775) <= not(layer1_outputs(7578));
    layer2_outputs(12776) <= layer1_outputs(11824);
    layer2_outputs(12777) <= not(layer1_outputs(8987));
    layer2_outputs(12778) <= (layer1_outputs(3043)) and not (layer1_outputs(1036));
    layer2_outputs(12779) <= not((layer1_outputs(12150)) xor (layer1_outputs(3405)));
    layer2_outputs(12780) <= (layer1_outputs(8045)) xor (layer1_outputs(4422));
    layer2_outputs(12781) <= (layer1_outputs(7449)) xor (layer1_outputs(6419));
    layer2_outputs(12782) <= (layer1_outputs(9594)) and (layer1_outputs(11141));
    layer2_outputs(12783) <= not((layer1_outputs(11157)) or (layer1_outputs(1701)));
    layer2_outputs(12784) <= layer1_outputs(11455);
    layer2_outputs(12785) <= layer1_outputs(479);
    layer2_outputs(12786) <= not(layer1_outputs(5311)) or (layer1_outputs(11902));
    layer2_outputs(12787) <= (layer1_outputs(8628)) xor (layer1_outputs(12245));
    layer2_outputs(12788) <= not((layer1_outputs(4161)) xor (layer1_outputs(5694)));
    layer2_outputs(12789) <= not(layer1_outputs(3244));
    layer2_outputs(12790) <= not((layer1_outputs(7249)) and (layer1_outputs(9985)));
    layer2_outputs(12791) <= not(layer1_outputs(9527));
    layer2_outputs(12792) <= (layer1_outputs(8998)) and (layer1_outputs(11298));
    layer2_outputs(12793) <= not(layer1_outputs(11509));
    layer2_outputs(12794) <= not(layer1_outputs(5500));
    layer2_outputs(12795) <= layer1_outputs(2129);
    layer2_outputs(12796) <= layer1_outputs(10281);
    layer2_outputs(12797) <= not((layer1_outputs(10693)) and (layer1_outputs(5774)));
    layer2_outputs(12798) <= not((layer1_outputs(8605)) xor (layer1_outputs(10213)));
    layer2_outputs(12799) <= (layer1_outputs(4616)) or (layer1_outputs(7352));
    outputs(0) <= (layer2_outputs(3241)) and not (layer2_outputs(40));
    outputs(1) <= not((layer2_outputs(11896)) xor (layer2_outputs(5388)));
    outputs(2) <= (layer2_outputs(12741)) xor (layer2_outputs(4720));
    outputs(3) <= not(layer2_outputs(9654)) or (layer2_outputs(787));
    outputs(4) <= (layer2_outputs(7134)) xor (layer2_outputs(4556));
    outputs(5) <= layer2_outputs(1508);
    outputs(6) <= not(layer2_outputs(5909));
    outputs(7) <= layer2_outputs(12707);
    outputs(8) <= layer2_outputs(192);
    outputs(9) <= layer2_outputs(4244);
    outputs(10) <= not(layer2_outputs(8345));
    outputs(11) <= not(layer2_outputs(12373));
    outputs(12) <= not(layer2_outputs(5295)) or (layer2_outputs(3894));
    outputs(13) <= (layer2_outputs(11018)) xor (layer2_outputs(3391));
    outputs(14) <= layer2_outputs(921);
    outputs(15) <= (layer2_outputs(12528)) xor (layer2_outputs(2984));
    outputs(16) <= not(layer2_outputs(10802));
    outputs(17) <= layer2_outputs(7337);
    outputs(18) <= layer2_outputs(8746);
    outputs(19) <= not((layer2_outputs(7257)) or (layer2_outputs(12123)));
    outputs(20) <= not(layer2_outputs(2053));
    outputs(21) <= (layer2_outputs(12135)) and not (layer2_outputs(10556));
    outputs(22) <= (layer2_outputs(6674)) xor (layer2_outputs(1633));
    outputs(23) <= (layer2_outputs(3684)) and (layer2_outputs(10142));
    outputs(24) <= (layer2_outputs(671)) or (layer2_outputs(3030));
    outputs(25) <= not(layer2_outputs(11018));
    outputs(26) <= layer2_outputs(1171);
    outputs(27) <= (layer2_outputs(12384)) xor (layer2_outputs(6870));
    outputs(28) <= not(layer2_outputs(11074));
    outputs(29) <= not(layer2_outputs(4273));
    outputs(30) <= not((layer2_outputs(7397)) xor (layer2_outputs(10243)));
    outputs(31) <= (layer2_outputs(6742)) and not (layer2_outputs(10906));
    outputs(32) <= not(layer2_outputs(11964));
    outputs(33) <= not(layer2_outputs(10954));
    outputs(34) <= not(layer2_outputs(12150));
    outputs(35) <= (layer2_outputs(9233)) and not (layer2_outputs(9256));
    outputs(36) <= not((layer2_outputs(6547)) xor (layer2_outputs(3808)));
    outputs(37) <= layer2_outputs(11473);
    outputs(38) <= not(layer2_outputs(9081));
    outputs(39) <= (layer2_outputs(7205)) and (layer2_outputs(8433));
    outputs(40) <= layer2_outputs(5770);
    outputs(41) <= not(layer2_outputs(7859));
    outputs(42) <= (layer2_outputs(2806)) or (layer2_outputs(7050));
    outputs(43) <= layer2_outputs(3237);
    outputs(44) <= not(layer2_outputs(12017));
    outputs(45) <= not(layer2_outputs(10537)) or (layer2_outputs(10977));
    outputs(46) <= layer2_outputs(8009);
    outputs(47) <= not(layer2_outputs(3456));
    outputs(48) <= layer2_outputs(8932);
    outputs(49) <= layer2_outputs(4272);
    outputs(50) <= layer2_outputs(5572);
    outputs(51) <= (layer2_outputs(1675)) and (layer2_outputs(9045));
    outputs(52) <= not(layer2_outputs(116));
    outputs(53) <= not(layer2_outputs(10048));
    outputs(54) <= (layer2_outputs(3937)) xor (layer2_outputs(2994));
    outputs(55) <= not((layer2_outputs(10065)) xor (layer2_outputs(5155)));
    outputs(56) <= layer2_outputs(6539);
    outputs(57) <= not(layer2_outputs(6900));
    outputs(58) <= layer2_outputs(2874);
    outputs(59) <= (layer2_outputs(2786)) xor (layer2_outputs(540));
    outputs(60) <= not(layer2_outputs(9297));
    outputs(61) <= layer2_outputs(7414);
    outputs(62) <= (layer2_outputs(8491)) and not (layer2_outputs(7037));
    outputs(63) <= not((layer2_outputs(507)) xor (layer2_outputs(6996)));
    outputs(64) <= not((layer2_outputs(477)) or (layer2_outputs(11495)));
    outputs(65) <= (layer2_outputs(4224)) and not (layer2_outputs(4887));
    outputs(66) <= layer2_outputs(6769);
    outputs(67) <= layer2_outputs(961);
    outputs(68) <= not((layer2_outputs(1616)) xor (layer2_outputs(3505)));
    outputs(69) <= not(layer2_outputs(4935));
    outputs(70) <= not(layer2_outputs(9874));
    outputs(71) <= (layer2_outputs(3463)) or (layer2_outputs(7498));
    outputs(72) <= not((layer2_outputs(3770)) xor (layer2_outputs(207)));
    outputs(73) <= not(layer2_outputs(2040));
    outputs(74) <= not((layer2_outputs(10065)) xor (layer2_outputs(2134)));
    outputs(75) <= not((layer2_outputs(3235)) and (layer2_outputs(11906)));
    outputs(76) <= (layer2_outputs(6215)) and not (layer2_outputs(11074));
    outputs(77) <= (layer2_outputs(10163)) and not (layer2_outputs(1720));
    outputs(78) <= layer2_outputs(9944);
    outputs(79) <= (layer2_outputs(8760)) xor (layer2_outputs(6173));
    outputs(80) <= not(layer2_outputs(30));
    outputs(81) <= not((layer2_outputs(5958)) or (layer2_outputs(12347)));
    outputs(82) <= layer2_outputs(8443);
    outputs(83) <= not((layer2_outputs(1785)) xor (layer2_outputs(9919)));
    outputs(84) <= layer2_outputs(10781);
    outputs(85) <= not(layer2_outputs(7501));
    outputs(86) <= layer2_outputs(708);
    outputs(87) <= not((layer2_outputs(5205)) and (layer2_outputs(7545)));
    outputs(88) <= layer2_outputs(11570);
    outputs(89) <= not(layer2_outputs(9842));
    outputs(90) <= not((layer2_outputs(4510)) xor (layer2_outputs(5340)));
    outputs(91) <= not(layer2_outputs(5288));
    outputs(92) <= not(layer2_outputs(9684));
    outputs(93) <= not((layer2_outputs(7306)) xor (layer2_outputs(9397)));
    outputs(94) <= not(layer2_outputs(5773));
    outputs(95) <= not(layer2_outputs(4957));
    outputs(96) <= (layer2_outputs(5497)) xor (layer2_outputs(3393));
    outputs(97) <= not((layer2_outputs(9573)) xor (layer2_outputs(10858)));
    outputs(98) <= not(layer2_outputs(11831));
    outputs(99) <= layer2_outputs(2088);
    outputs(100) <= not(layer2_outputs(11799));
    outputs(101) <= (layer2_outputs(2310)) and not (layer2_outputs(11090));
    outputs(102) <= not(layer2_outputs(2450));
    outputs(103) <= (layer2_outputs(12430)) xor (layer2_outputs(6329));
    outputs(104) <= not((layer2_outputs(5506)) xor (layer2_outputs(7677)));
    outputs(105) <= not(layer2_outputs(5108));
    outputs(106) <= (layer2_outputs(11783)) xor (layer2_outputs(5017));
    outputs(107) <= not(layer2_outputs(11834));
    outputs(108) <= layer2_outputs(5756);
    outputs(109) <= layer2_outputs(7062);
    outputs(110) <= layer2_outputs(159);
    outputs(111) <= not(layer2_outputs(11712)) or (layer2_outputs(7851));
    outputs(112) <= (layer2_outputs(6409)) and not (layer2_outputs(2006));
    outputs(113) <= layer2_outputs(7326);
    outputs(114) <= (layer2_outputs(1131)) xor (layer2_outputs(6265));
    outputs(115) <= not(layer2_outputs(8369));
    outputs(116) <= not(layer2_outputs(4957));
    outputs(117) <= not(layer2_outputs(6237));
    outputs(118) <= not(layer2_outputs(12303));
    outputs(119) <= layer2_outputs(3697);
    outputs(120) <= not((layer2_outputs(9319)) xor (layer2_outputs(11654)));
    outputs(121) <= layer2_outputs(11418);
    outputs(122) <= not(layer2_outputs(11179)) or (layer2_outputs(6907));
    outputs(123) <= layer2_outputs(7482);
    outputs(124) <= not((layer2_outputs(7736)) xor (layer2_outputs(3181)));
    outputs(125) <= layer2_outputs(9609);
    outputs(126) <= not((layer2_outputs(2313)) and (layer2_outputs(3056)));
    outputs(127) <= not(layer2_outputs(2081));
    outputs(128) <= layer2_outputs(11197);
    outputs(129) <= not(layer2_outputs(11391));
    outputs(130) <= layer2_outputs(1800);
    outputs(131) <= not(layer2_outputs(593));
    outputs(132) <= not(layer2_outputs(2147));
    outputs(133) <= layer2_outputs(11214);
    outputs(134) <= layer2_outputs(1913);
    outputs(135) <= not((layer2_outputs(6581)) and (layer2_outputs(11961)));
    outputs(136) <= not(layer2_outputs(9130)) or (layer2_outputs(327));
    outputs(137) <= not(layer2_outputs(7935));
    outputs(138) <= layer2_outputs(6208);
    outputs(139) <= not((layer2_outputs(7488)) xor (layer2_outputs(7116)));
    outputs(140) <= (layer2_outputs(8941)) and not (layer2_outputs(86));
    outputs(141) <= layer2_outputs(9858);
    outputs(142) <= layer2_outputs(11197);
    outputs(143) <= layer2_outputs(7839);
    outputs(144) <= not(layer2_outputs(4637));
    outputs(145) <= not((layer2_outputs(11475)) xor (layer2_outputs(7229)));
    outputs(146) <= not(layer2_outputs(5767));
    outputs(147) <= layer2_outputs(8801);
    outputs(148) <= not((layer2_outputs(11630)) xor (layer2_outputs(6371)));
    outputs(149) <= not(layer2_outputs(6179));
    outputs(150) <= layer2_outputs(126);
    outputs(151) <= layer2_outputs(3609);
    outputs(152) <= not((layer2_outputs(10254)) xor (layer2_outputs(7070)));
    outputs(153) <= not(layer2_outputs(11190));
    outputs(154) <= (layer2_outputs(9111)) and not (layer2_outputs(10023));
    outputs(155) <= not(layer2_outputs(1720)) or (layer2_outputs(6313));
    outputs(156) <= not(layer2_outputs(10229));
    outputs(157) <= not(layer2_outputs(7076));
    outputs(158) <= layer2_outputs(3102);
    outputs(159) <= not(layer2_outputs(6760));
    outputs(160) <= not(layer2_outputs(10307));
    outputs(161) <= layer2_outputs(3731);
    outputs(162) <= layer2_outputs(3616);
    outputs(163) <= layer2_outputs(6723);
    outputs(164) <= layer2_outputs(7118);
    outputs(165) <= not(layer2_outputs(12480));
    outputs(166) <= layer2_outputs(10703);
    outputs(167) <= (layer2_outputs(1040)) and not (layer2_outputs(8059));
    outputs(168) <= not(layer2_outputs(3849));
    outputs(169) <= layer2_outputs(11490);
    outputs(170) <= (layer2_outputs(3552)) xor (layer2_outputs(9264));
    outputs(171) <= layer2_outputs(6231);
    outputs(172) <= not(layer2_outputs(8822));
    outputs(173) <= not((layer2_outputs(3492)) xor (layer2_outputs(7744)));
    outputs(174) <= (layer2_outputs(3423)) and (layer2_outputs(10267));
    outputs(175) <= (layer2_outputs(12422)) and (layer2_outputs(5648));
    outputs(176) <= (layer2_outputs(2922)) xor (layer2_outputs(10695));
    outputs(177) <= layer2_outputs(4462);
    outputs(178) <= not(layer2_outputs(9727));
    outputs(179) <= layer2_outputs(11451);
    outputs(180) <= layer2_outputs(10133);
    outputs(181) <= not((layer2_outputs(3244)) or (layer2_outputs(8678)));
    outputs(182) <= layer2_outputs(12403);
    outputs(183) <= (layer2_outputs(5870)) xor (layer2_outputs(11549));
    outputs(184) <= not(layer2_outputs(6125));
    outputs(185) <= layer2_outputs(4234);
    outputs(186) <= not(layer2_outputs(2640));
    outputs(187) <= not(layer2_outputs(11276));
    outputs(188) <= not((layer2_outputs(12766)) xor (layer2_outputs(6022)));
    outputs(189) <= not(layer2_outputs(11947));
    outputs(190) <= not(layer2_outputs(7666));
    outputs(191) <= not(layer2_outputs(7173));
    outputs(192) <= not((layer2_outputs(11345)) xor (layer2_outputs(8537)));
    outputs(193) <= not(layer2_outputs(7167)) or (layer2_outputs(3540));
    outputs(194) <= layer2_outputs(12184);
    outputs(195) <= (layer2_outputs(9942)) xor (layer2_outputs(11176));
    outputs(196) <= not((layer2_outputs(12153)) xor (layer2_outputs(6354)));
    outputs(197) <= layer2_outputs(122);
    outputs(198) <= not(layer2_outputs(10683));
    outputs(199) <= not((layer2_outputs(5603)) xor (layer2_outputs(4161)));
    outputs(200) <= layer2_outputs(1550);
    outputs(201) <= (layer2_outputs(11988)) or (layer2_outputs(11876));
    outputs(202) <= not(layer2_outputs(4324));
    outputs(203) <= not(layer2_outputs(3597));
    outputs(204) <= not(layer2_outputs(1615));
    outputs(205) <= layer2_outputs(12161);
    outputs(206) <= not(layer2_outputs(5260));
    outputs(207) <= layer2_outputs(715);
    outputs(208) <= not(layer2_outputs(10810));
    outputs(209) <= not(layer2_outputs(4993));
    outputs(210) <= (layer2_outputs(9688)) and (layer2_outputs(4373));
    outputs(211) <= (layer2_outputs(3214)) and not (layer2_outputs(2739));
    outputs(212) <= (layer2_outputs(10916)) and not (layer2_outputs(6137));
    outputs(213) <= (layer2_outputs(2296)) xor (layer2_outputs(1932));
    outputs(214) <= not(layer2_outputs(3156));
    outputs(215) <= not((layer2_outputs(6922)) xor (layer2_outputs(2729)));
    outputs(216) <= not((layer2_outputs(3862)) xor (layer2_outputs(9933)));
    outputs(217) <= (layer2_outputs(8733)) xor (layer2_outputs(10465));
    outputs(218) <= layer2_outputs(10413);
    outputs(219) <= not((layer2_outputs(10589)) xor (layer2_outputs(6698)));
    outputs(220) <= (layer2_outputs(1746)) and not (layer2_outputs(186));
    outputs(221) <= not(layer2_outputs(12150));
    outputs(222) <= (layer2_outputs(6509)) and not (layer2_outputs(4882));
    outputs(223) <= layer2_outputs(7816);
    outputs(224) <= (layer2_outputs(8385)) and not (layer2_outputs(9665));
    outputs(225) <= not(layer2_outputs(11319));
    outputs(226) <= not(layer2_outputs(9268));
    outputs(227) <= not((layer2_outputs(12390)) xor (layer2_outputs(6636)));
    outputs(228) <= (layer2_outputs(3598)) xor (layer2_outputs(8165));
    outputs(229) <= layer2_outputs(822);
    outputs(230) <= not((layer2_outputs(843)) and (layer2_outputs(1688)));
    outputs(231) <= not(layer2_outputs(9137));
    outputs(232) <= not(layer2_outputs(5773));
    outputs(233) <= not(layer2_outputs(2607));
    outputs(234) <= (layer2_outputs(8307)) and (layer2_outputs(5517));
    outputs(235) <= layer2_outputs(1620);
    outputs(236) <= (layer2_outputs(7376)) and (layer2_outputs(8711));
    outputs(237) <= layer2_outputs(244);
    outputs(238) <= not(layer2_outputs(7813));
    outputs(239) <= (layer2_outputs(9439)) and (layer2_outputs(10345));
    outputs(240) <= layer2_outputs(6877);
    outputs(241) <= not(layer2_outputs(8376));
    outputs(242) <= (layer2_outputs(11807)) and (layer2_outputs(9488));
    outputs(243) <= (layer2_outputs(8067)) and not (layer2_outputs(7020));
    outputs(244) <= layer2_outputs(8611);
    outputs(245) <= layer2_outputs(10981);
    outputs(246) <= layer2_outputs(3105);
    outputs(247) <= layer2_outputs(10439);
    outputs(248) <= layer2_outputs(11769);
    outputs(249) <= not(layer2_outputs(586));
    outputs(250) <= layer2_outputs(9922);
    outputs(251) <= not(layer2_outputs(2410));
    outputs(252) <= not(layer2_outputs(9459));
    outputs(253) <= (layer2_outputs(7681)) xor (layer2_outputs(6327));
    outputs(254) <= (layer2_outputs(2462)) and (layer2_outputs(10890));
    outputs(255) <= not((layer2_outputs(10499)) and (layer2_outputs(3788)));
    outputs(256) <= (layer2_outputs(5772)) and (layer2_outputs(131));
    outputs(257) <= layer2_outputs(5941);
    outputs(258) <= not((layer2_outputs(2500)) xor (layer2_outputs(456)));
    outputs(259) <= layer2_outputs(4475);
    outputs(260) <= not((layer2_outputs(8603)) xor (layer2_outputs(10805)));
    outputs(261) <= layer2_outputs(11285);
    outputs(262) <= (layer2_outputs(9152)) and not (layer2_outputs(1680));
    outputs(263) <= layer2_outputs(638);
    outputs(264) <= not((layer2_outputs(5709)) xor (layer2_outputs(10341)));
    outputs(265) <= layer2_outputs(10204);
    outputs(266) <= layer2_outputs(3900);
    outputs(267) <= not(layer2_outputs(2747));
    outputs(268) <= layer2_outputs(10752);
    outputs(269) <= not((layer2_outputs(6672)) or (layer2_outputs(519)));
    outputs(270) <= not(layer2_outputs(19));
    outputs(271) <= layer2_outputs(10959);
    outputs(272) <= layer2_outputs(8511);
    outputs(273) <= layer2_outputs(4155);
    outputs(274) <= not((layer2_outputs(3807)) xor (layer2_outputs(6775)));
    outputs(275) <= not(layer2_outputs(7462));
    outputs(276) <= (layer2_outputs(6700)) and (layer2_outputs(8360));
    outputs(277) <= not((layer2_outputs(7374)) xor (layer2_outputs(6459)));
    outputs(278) <= not(layer2_outputs(7855)) or (layer2_outputs(3441));
    outputs(279) <= not((layer2_outputs(825)) xor (layer2_outputs(829)));
    outputs(280) <= not(layer2_outputs(1150));
    outputs(281) <= not(layer2_outputs(7565));
    outputs(282) <= not(layer2_outputs(1283));
    outputs(283) <= not(layer2_outputs(10946));
    outputs(284) <= not(layer2_outputs(2634));
    outputs(285) <= layer2_outputs(2834);
    outputs(286) <= not(layer2_outputs(5672));
    outputs(287) <= not(layer2_outputs(9950));
    outputs(288) <= layer2_outputs(10227);
    outputs(289) <= not(layer2_outputs(10430));
    outputs(290) <= (layer2_outputs(5964)) and (layer2_outputs(3025));
    outputs(291) <= layer2_outputs(4227);
    outputs(292) <= layer2_outputs(3034);
    outputs(293) <= layer2_outputs(907);
    outputs(294) <= layer2_outputs(591);
    outputs(295) <= not(layer2_outputs(1373));
    outputs(296) <= (layer2_outputs(1454)) xor (layer2_outputs(10551));
    outputs(297) <= not((layer2_outputs(5297)) xor (layer2_outputs(1019)));
    outputs(298) <= not((layer2_outputs(3381)) or (layer2_outputs(5807)));
    outputs(299) <= not((layer2_outputs(10383)) xor (layer2_outputs(9540)));
    outputs(300) <= layer2_outputs(439);
    outputs(301) <= not((layer2_outputs(3374)) xor (layer2_outputs(8626)));
    outputs(302) <= layer2_outputs(12259);
    outputs(303) <= (layer2_outputs(7226)) and (layer2_outputs(8752));
    outputs(304) <= layer2_outputs(5196);
    outputs(305) <= not(layer2_outputs(6852));
    outputs(306) <= not((layer2_outputs(7575)) xor (layer2_outputs(12060)));
    outputs(307) <= not((layer2_outputs(11599)) xor (layer2_outputs(10301)));
    outputs(308) <= not((layer2_outputs(5881)) and (layer2_outputs(3387)));
    outputs(309) <= layer2_outputs(2048);
    outputs(310) <= not(layer2_outputs(12139));
    outputs(311) <= not(layer2_outputs(5339));
    outputs(312) <= (layer2_outputs(10265)) and not (layer2_outputs(2128));
    outputs(313) <= (layer2_outputs(9979)) and (layer2_outputs(2305));
    outputs(314) <= layer2_outputs(8502);
    outputs(315) <= not(layer2_outputs(7874));
    outputs(316) <= layer2_outputs(4082);
    outputs(317) <= layer2_outputs(4960);
    outputs(318) <= layer2_outputs(8731);
    outputs(319) <= not((layer2_outputs(269)) xor (layer2_outputs(6218)));
    outputs(320) <= not(layer2_outputs(3582));
    outputs(321) <= layer2_outputs(7617);
    outputs(322) <= not((layer2_outputs(6832)) or (layer2_outputs(3531)));
    outputs(323) <= layer2_outputs(910);
    outputs(324) <= not(layer2_outputs(5172));
    outputs(325) <= (layer2_outputs(5057)) xor (layer2_outputs(9674));
    outputs(326) <= (layer2_outputs(3212)) and not (layer2_outputs(1869));
    outputs(327) <= not(layer2_outputs(8345));
    outputs(328) <= not(layer2_outputs(3141));
    outputs(329) <= layer2_outputs(1915);
    outputs(330) <= not((layer2_outputs(12740)) xor (layer2_outputs(9435)));
    outputs(331) <= layer2_outputs(2188);
    outputs(332) <= layer2_outputs(2026);
    outputs(333) <= (layer2_outputs(4672)) xor (layer2_outputs(6094));
    outputs(334) <= layer2_outputs(10481);
    outputs(335) <= not((layer2_outputs(2944)) xor (layer2_outputs(11247)));
    outputs(336) <= layer2_outputs(9240);
    outputs(337) <= layer2_outputs(6174);
    outputs(338) <= (layer2_outputs(4966)) xor (layer2_outputs(10464));
    outputs(339) <= layer2_outputs(3559);
    outputs(340) <= not(layer2_outputs(1862));
    outputs(341) <= not(layer2_outputs(11516)) or (layer2_outputs(784));
    outputs(342) <= not((layer2_outputs(3148)) xor (layer2_outputs(1425)));
    outputs(343) <= not(layer2_outputs(3930));
    outputs(344) <= (layer2_outputs(10733)) xor (layer2_outputs(9918));
    outputs(345) <= not(layer2_outputs(2921)) or (layer2_outputs(8806));
    outputs(346) <= layer2_outputs(467);
    outputs(347) <= layer2_outputs(7287);
    outputs(348) <= not(layer2_outputs(1383));
    outputs(349) <= not(layer2_outputs(725));
    outputs(350) <= not((layer2_outputs(6807)) xor (layer2_outputs(11702)));
    outputs(351) <= not((layer2_outputs(3837)) and (layer2_outputs(9741)));
    outputs(352) <= not((layer2_outputs(1979)) xor (layer2_outputs(11129)));
    outputs(353) <= not(layer2_outputs(7291));
    outputs(354) <= not(layer2_outputs(9906));
    outputs(355) <= not(layer2_outputs(9245));
    outputs(356) <= not((layer2_outputs(12090)) xor (layer2_outputs(10768)));
    outputs(357) <= not(layer2_outputs(2677));
    outputs(358) <= layer2_outputs(652);
    outputs(359) <= not((layer2_outputs(12091)) xor (layer2_outputs(11405)));
    outputs(360) <= not(layer2_outputs(5915));
    outputs(361) <= not((layer2_outputs(3969)) xor (layer2_outputs(5284)));
    outputs(362) <= not(layer2_outputs(1187)) or (layer2_outputs(6064));
    outputs(363) <= (layer2_outputs(7152)) and not (layer2_outputs(8220));
    outputs(364) <= not((layer2_outputs(10195)) xor (layer2_outputs(5548)));
    outputs(365) <= layer2_outputs(10866);
    outputs(366) <= not(layer2_outputs(6315));
    outputs(367) <= (layer2_outputs(183)) and not (layer2_outputs(6371));
    outputs(368) <= not((layer2_outputs(10587)) xor (layer2_outputs(5989)));
    outputs(369) <= not(layer2_outputs(1346));
    outputs(370) <= layer2_outputs(4029);
    outputs(371) <= layer2_outputs(9703);
    outputs(372) <= not((layer2_outputs(9080)) xor (layer2_outputs(9777)));
    outputs(373) <= not(layer2_outputs(11647));
    outputs(374) <= not(layer2_outputs(7636));
    outputs(375) <= not(layer2_outputs(11598));
    outputs(376) <= not(layer2_outputs(10363));
    outputs(377) <= layer2_outputs(5042);
    outputs(378) <= '0';
    outputs(379) <= (layer2_outputs(10743)) and (layer2_outputs(4376));
    outputs(380) <= not((layer2_outputs(5355)) or (layer2_outputs(8342)));
    outputs(381) <= not((layer2_outputs(8644)) or (layer2_outputs(8285)));
    outputs(382) <= not(layer2_outputs(8377));
    outputs(383) <= layer2_outputs(7212);
    outputs(384) <= not(layer2_outputs(5062));
    outputs(385) <= not((layer2_outputs(1870)) or (layer2_outputs(9594)));
    outputs(386) <= (layer2_outputs(6121)) and (layer2_outputs(11628));
    outputs(387) <= (layer2_outputs(7179)) xor (layer2_outputs(12035));
    outputs(388) <= not((layer2_outputs(4847)) xor (layer2_outputs(4073)));
    outputs(389) <= (layer2_outputs(6443)) and not (layer2_outputs(10789));
    outputs(390) <= layer2_outputs(11196);
    outputs(391) <= (layer2_outputs(21)) xor (layer2_outputs(9482));
    outputs(392) <= not(layer2_outputs(5146));
    outputs(393) <= (layer2_outputs(12543)) and (layer2_outputs(12579));
    outputs(394) <= (layer2_outputs(4843)) xor (layer2_outputs(1051));
    outputs(395) <= layer2_outputs(6443);
    outputs(396) <= not((layer2_outputs(11514)) and (layer2_outputs(7838)));
    outputs(397) <= layer2_outputs(2158);
    outputs(398) <= layer2_outputs(1891);
    outputs(399) <= layer2_outputs(9135);
    outputs(400) <= not(layer2_outputs(3344));
    outputs(401) <= not((layer2_outputs(4720)) and (layer2_outputs(11345)));
    outputs(402) <= not(layer2_outputs(11610));
    outputs(403) <= not(layer2_outputs(12787));
    outputs(404) <= not((layer2_outputs(12162)) xor (layer2_outputs(9708)));
    outputs(405) <= (layer2_outputs(79)) xor (layer2_outputs(10436));
    outputs(406) <= not((layer2_outputs(12386)) xor (layer2_outputs(5952)));
    outputs(407) <= not(layer2_outputs(1473)) or (layer2_outputs(8842));
    outputs(408) <= layer2_outputs(8698);
    outputs(409) <= not(layer2_outputs(2492)) or (layer2_outputs(10882));
    outputs(410) <= not(layer2_outputs(1678));
    outputs(411) <= layer2_outputs(2539);
    outputs(412) <= layer2_outputs(8947);
    outputs(413) <= layer2_outputs(1368);
    outputs(414) <= (layer2_outputs(9345)) and (layer2_outputs(6778));
    outputs(415) <= not((layer2_outputs(12179)) xor (layer2_outputs(4133)));
    outputs(416) <= not(layer2_outputs(8147));
    outputs(417) <= not(layer2_outputs(5541));
    outputs(418) <= not(layer2_outputs(3962)) or (layer2_outputs(701));
    outputs(419) <= not(layer2_outputs(1553));
    outputs(420) <= layer2_outputs(5843);
    outputs(421) <= layer2_outputs(9215);
    outputs(422) <= not((layer2_outputs(2334)) xor (layer2_outputs(63)));
    outputs(423) <= not(layer2_outputs(10437));
    outputs(424) <= (layer2_outputs(1868)) and not (layer2_outputs(6402));
    outputs(425) <= layer2_outputs(3904);
    outputs(426) <= not(layer2_outputs(10239));
    outputs(427) <= layer2_outputs(1506);
    outputs(428) <= layer2_outputs(3102);
    outputs(429) <= not(layer2_outputs(212));
    outputs(430) <= (layer2_outputs(1317)) xor (layer2_outputs(10102));
    outputs(431) <= not(layer2_outputs(3155));
    outputs(432) <= not(layer2_outputs(1192));
    outputs(433) <= layer2_outputs(2412);
    outputs(434) <= layer2_outputs(8418);
    outputs(435) <= not(layer2_outputs(12251));
    outputs(436) <= not((layer2_outputs(1086)) xor (layer2_outputs(11918)));
    outputs(437) <= not((layer2_outputs(7829)) or (layer2_outputs(12066)));
    outputs(438) <= not(layer2_outputs(8262));
    outputs(439) <= (layer2_outputs(10403)) and not (layer2_outputs(6117));
    outputs(440) <= (layer2_outputs(9334)) and (layer2_outputs(5018));
    outputs(441) <= layer2_outputs(5028);
    outputs(442) <= layer2_outputs(726);
    outputs(443) <= not(layer2_outputs(554));
    outputs(444) <= (layer2_outputs(9614)) xor (layer2_outputs(12063));
    outputs(445) <= not(layer2_outputs(10295));
    outputs(446) <= not((layer2_outputs(10992)) or (layer2_outputs(12357)));
    outputs(447) <= not((layer2_outputs(2963)) xor (layer2_outputs(8038)));
    outputs(448) <= layer2_outputs(8916);
    outputs(449) <= not(layer2_outputs(2156));
    outputs(450) <= layer2_outputs(5553);
    outputs(451) <= layer2_outputs(3649);
    outputs(452) <= not((layer2_outputs(103)) xor (layer2_outputs(9742)));
    outputs(453) <= not(layer2_outputs(12556)) or (layer2_outputs(1168));
    outputs(454) <= layer2_outputs(7626);
    outputs(455) <= not((layer2_outputs(270)) xor (layer2_outputs(11581)));
    outputs(456) <= (layer2_outputs(9905)) xor (layer2_outputs(4732));
    outputs(457) <= not(layer2_outputs(8757));
    outputs(458) <= not((layer2_outputs(1409)) and (layer2_outputs(2303)));
    outputs(459) <= not(layer2_outputs(2049));
    outputs(460) <= not((layer2_outputs(443)) xor (layer2_outputs(4164)));
    outputs(461) <= layer2_outputs(9413);
    outputs(462) <= layer2_outputs(5140);
    outputs(463) <= not((layer2_outputs(622)) xor (layer2_outputs(7720)));
    outputs(464) <= not(layer2_outputs(8215));
    outputs(465) <= layer2_outputs(6431);
    outputs(466) <= (layer2_outputs(4931)) and not (layer2_outputs(826));
    outputs(467) <= not((layer2_outputs(8850)) xor (layer2_outputs(9289)));
    outputs(468) <= not(layer2_outputs(9034));
    outputs(469) <= layer2_outputs(2705);
    outputs(470) <= (layer2_outputs(1248)) or (layer2_outputs(74));
    outputs(471) <= (layer2_outputs(9438)) and not (layer2_outputs(10284));
    outputs(472) <= not(layer2_outputs(4039));
    outputs(473) <= layer2_outputs(4399);
    outputs(474) <= layer2_outputs(1391);
    outputs(475) <= not(layer2_outputs(2888));
    outputs(476) <= layer2_outputs(7920);
    outputs(477) <= not((layer2_outputs(10186)) xor (layer2_outputs(5739)));
    outputs(478) <= not(layer2_outputs(5060));
    outputs(479) <= layer2_outputs(10244);
    outputs(480) <= (layer2_outputs(12694)) or (layer2_outputs(6407));
    outputs(481) <= (layer2_outputs(2882)) xor (layer2_outputs(5659));
    outputs(482) <= layer2_outputs(1699);
    outputs(483) <= layer2_outputs(806);
    outputs(484) <= not(layer2_outputs(12263));
    outputs(485) <= not((layer2_outputs(12497)) xor (layer2_outputs(10687)));
    outputs(486) <= layer2_outputs(9872);
    outputs(487) <= (layer2_outputs(5845)) xor (layer2_outputs(11013));
    outputs(488) <= not(layer2_outputs(9678));
    outputs(489) <= layer2_outputs(12223);
    outputs(490) <= not(layer2_outputs(9280));
    outputs(491) <= not(layer2_outputs(9365)) or (layer2_outputs(9868));
    outputs(492) <= not(layer2_outputs(12589));
    outputs(493) <= (layer2_outputs(3025)) and not (layer2_outputs(1213));
    outputs(494) <= not(layer2_outputs(6894));
    outputs(495) <= not(layer2_outputs(11072));
    outputs(496) <= (layer2_outputs(9929)) xor (layer2_outputs(2334));
    outputs(497) <= layer2_outputs(2406);
    outputs(498) <= not((layer2_outputs(73)) xor (layer2_outputs(10345)));
    outputs(499) <= layer2_outputs(3626);
    outputs(500) <= (layer2_outputs(11530)) xor (layer2_outputs(5925));
    outputs(501) <= layer2_outputs(4288);
    outputs(502) <= not(layer2_outputs(11686));
    outputs(503) <= (layer2_outputs(223)) or (layer2_outputs(9051));
    outputs(504) <= not(layer2_outputs(12407));
    outputs(505) <= layer2_outputs(8726);
    outputs(506) <= not((layer2_outputs(3474)) xor (layer2_outputs(8042)));
    outputs(507) <= not((layer2_outputs(8275)) xor (layer2_outputs(1896)));
    outputs(508) <= not(layer2_outputs(4492));
    outputs(509) <= (layer2_outputs(3649)) and not (layer2_outputs(5413));
    outputs(510) <= (layer2_outputs(12133)) xor (layer2_outputs(9231));
    outputs(511) <= (layer2_outputs(5467)) and (layer2_outputs(163));
    outputs(512) <= not(layer2_outputs(3631));
    outputs(513) <= (layer2_outputs(11889)) xor (layer2_outputs(3355));
    outputs(514) <= not((layer2_outputs(1977)) xor (layer2_outputs(11760)));
    outputs(515) <= not(layer2_outputs(7310));
    outputs(516) <= (layer2_outputs(7877)) xor (layer2_outputs(12448));
    outputs(517) <= layer2_outputs(8365);
    outputs(518) <= layer2_outputs(11228);
    outputs(519) <= not((layer2_outputs(12064)) xor (layer2_outputs(10396)));
    outputs(520) <= layer2_outputs(4060);
    outputs(521) <= not(layer2_outputs(2747));
    outputs(522) <= not(layer2_outputs(3349));
    outputs(523) <= (layer2_outputs(6272)) and (layer2_outputs(10273));
    outputs(524) <= not(layer2_outputs(496));
    outputs(525) <= not(layer2_outputs(10492));
    outputs(526) <= not(layer2_outputs(7254)) or (layer2_outputs(4894));
    outputs(527) <= (layer2_outputs(5653)) and not (layer2_outputs(9593));
    outputs(528) <= layer2_outputs(10961);
    outputs(529) <= layer2_outputs(616);
    outputs(530) <= layer2_outputs(10627);
    outputs(531) <= not((layer2_outputs(11249)) or (layer2_outputs(9943)));
    outputs(532) <= (layer2_outputs(2257)) and not (layer2_outputs(10233));
    outputs(533) <= (layer2_outputs(6166)) or (layer2_outputs(395));
    outputs(534) <= not(layer2_outputs(3768));
    outputs(535) <= layer2_outputs(1388);
    outputs(536) <= (layer2_outputs(12590)) xor (layer2_outputs(11468));
    outputs(537) <= not(layer2_outputs(8738));
    outputs(538) <= (layer2_outputs(125)) xor (layer2_outputs(7734));
    outputs(539) <= layer2_outputs(7861);
    outputs(540) <= (layer2_outputs(6966)) and (layer2_outputs(9909));
    outputs(541) <= not((layer2_outputs(12011)) and (layer2_outputs(4760)));
    outputs(542) <= not(layer2_outputs(6455));
    outputs(543) <= not(layer2_outputs(8086));
    outputs(544) <= not(layer2_outputs(1396)) or (layer2_outputs(6436));
    outputs(545) <= not(layer2_outputs(5835)) or (layer2_outputs(11379));
    outputs(546) <= not(layer2_outputs(353));
    outputs(547) <= not(layer2_outputs(3185));
    outputs(548) <= (layer2_outputs(31)) xor (layer2_outputs(9336));
    outputs(549) <= layer2_outputs(1507);
    outputs(550) <= layer2_outputs(258);
    outputs(551) <= not(layer2_outputs(4001)) or (layer2_outputs(2388));
    outputs(552) <= not(layer2_outputs(10460));
    outputs(553) <= not(layer2_outputs(5012));
    outputs(554) <= layer2_outputs(9765);
    outputs(555) <= (layer2_outputs(10782)) or (layer2_outputs(5643));
    outputs(556) <= not(layer2_outputs(3163)) or (layer2_outputs(4572));
    outputs(557) <= not(layer2_outputs(837));
    outputs(558) <= not(layer2_outputs(1613));
    outputs(559) <= layer2_outputs(6183);
    outputs(560) <= not(layer2_outputs(10620));
    outputs(561) <= not(layer2_outputs(1534));
    outputs(562) <= layer2_outputs(465);
    outputs(563) <= (layer2_outputs(6480)) and not (layer2_outputs(562));
    outputs(564) <= layer2_outputs(4127);
    outputs(565) <= (layer2_outputs(1599)) and not (layer2_outputs(9864));
    outputs(566) <= not(layer2_outputs(5742)) or (layer2_outputs(12316));
    outputs(567) <= not((layer2_outputs(426)) xor (layer2_outputs(11826)));
    outputs(568) <= layer2_outputs(3010);
    outputs(569) <= not(layer2_outputs(1754));
    outputs(570) <= (layer2_outputs(4180)) xor (layer2_outputs(2096));
    outputs(571) <= not(layer2_outputs(1797));
    outputs(572) <= not(layer2_outputs(8287));
    outputs(573) <= (layer2_outputs(10493)) and not (layer2_outputs(4156));
    outputs(574) <= not(layer2_outputs(3916)) or (layer2_outputs(9129));
    outputs(575) <= (layer2_outputs(5052)) xor (layer2_outputs(2776));
    outputs(576) <= not(layer2_outputs(6173)) or (layer2_outputs(8022));
    outputs(577) <= layer2_outputs(11196);
    outputs(578) <= layer2_outputs(9832);
    outputs(579) <= (layer2_outputs(10378)) xor (layer2_outputs(10570));
    outputs(580) <= not(layer2_outputs(10027));
    outputs(581) <= not(layer2_outputs(6611));
    outputs(582) <= not(layer2_outputs(11226));
    outputs(583) <= (layer2_outputs(3751)) xor (layer2_outputs(4793));
    outputs(584) <= not(layer2_outputs(10636));
    outputs(585) <= not(layer2_outputs(6422));
    outputs(586) <= (layer2_outputs(7645)) or (layer2_outputs(10385));
    outputs(587) <= layer2_outputs(6282);
    outputs(588) <= layer2_outputs(4833);
    outputs(589) <= not(layer2_outputs(4905));
    outputs(590) <= not(layer2_outputs(11865));
    outputs(591) <= not(layer2_outputs(3748));
    outputs(592) <= not((layer2_outputs(7199)) and (layer2_outputs(10321)));
    outputs(593) <= not((layer2_outputs(2778)) xor (layer2_outputs(8193)));
    outputs(594) <= not(layer2_outputs(3204)) or (layer2_outputs(6073));
    outputs(595) <= layer2_outputs(10273);
    outputs(596) <= (layer2_outputs(3079)) or (layer2_outputs(5439));
    outputs(597) <= (layer2_outputs(11480)) and not (layer2_outputs(3018));
    outputs(598) <= not(layer2_outputs(5814)) or (layer2_outputs(3101));
    outputs(599) <= not(layer2_outputs(5846));
    outputs(600) <= not(layer2_outputs(7027));
    outputs(601) <= not(layer2_outputs(1627)) or (layer2_outputs(5196));
    outputs(602) <= layer2_outputs(7683);
    outputs(603) <= (layer2_outputs(6926)) xor (layer2_outputs(3270));
    outputs(604) <= not((layer2_outputs(7316)) xor (layer2_outputs(3150)));
    outputs(605) <= (layer2_outputs(9849)) and not (layer2_outputs(6209));
    outputs(606) <= layer2_outputs(2478);
    outputs(607) <= (layer2_outputs(667)) xor (layer2_outputs(7629));
    outputs(608) <= not(layer2_outputs(8970));
    outputs(609) <= layer2_outputs(11128);
    outputs(610) <= layer2_outputs(12023);
    outputs(611) <= layer2_outputs(8403);
    outputs(612) <= (layer2_outputs(21)) and not (layer2_outputs(1143));
    outputs(613) <= not(layer2_outputs(1264));
    outputs(614) <= not(layer2_outputs(11237));
    outputs(615) <= layer2_outputs(9170);
    outputs(616) <= (layer2_outputs(6925)) and not (layer2_outputs(9562));
    outputs(617) <= not(layer2_outputs(5504));
    outputs(618) <= layer2_outputs(6415);
    outputs(619) <= layer2_outputs(10488);
    outputs(620) <= not((layer2_outputs(4896)) xor (layer2_outputs(5916)));
    outputs(621) <= not((layer2_outputs(2397)) xor (layer2_outputs(2716)));
    outputs(622) <= not((layer2_outputs(5417)) xor (layer2_outputs(9582)));
    outputs(623) <= (layer2_outputs(6669)) xor (layer2_outputs(5826));
    outputs(624) <= not((layer2_outputs(4055)) xor (layer2_outputs(4968)));
    outputs(625) <= not((layer2_outputs(5375)) xor (layer2_outputs(11650)));
    outputs(626) <= layer2_outputs(5988);
    outputs(627) <= not(layer2_outputs(12035));
    outputs(628) <= (layer2_outputs(10953)) xor (layer2_outputs(495));
    outputs(629) <= not(layer2_outputs(7502));
    outputs(630) <= layer2_outputs(10515);
    outputs(631) <= not(layer2_outputs(9706));
    outputs(632) <= layer2_outputs(8375);
    outputs(633) <= not(layer2_outputs(10389));
    outputs(634) <= not((layer2_outputs(6400)) and (layer2_outputs(12125)));
    outputs(635) <= not(layer2_outputs(132));
    outputs(636) <= not(layer2_outputs(1180)) or (layer2_outputs(93));
    outputs(637) <= layer2_outputs(1935);
    outputs(638) <= layer2_outputs(3910);
    outputs(639) <= not(layer2_outputs(2948));
    outputs(640) <= (layer2_outputs(10525)) and not (layer2_outputs(6146));
    outputs(641) <= not((layer2_outputs(3785)) and (layer2_outputs(4573)));
    outputs(642) <= not(layer2_outputs(2246));
    outputs(643) <= layer2_outputs(9318);
    outputs(644) <= not(layer2_outputs(6011));
    outputs(645) <= layer2_outputs(11988);
    outputs(646) <= layer2_outputs(2749);
    outputs(647) <= layer2_outputs(3441);
    outputs(648) <= not(layer2_outputs(12738)) or (layer2_outputs(6466));
    outputs(649) <= not(layer2_outputs(6558));
    outputs(650) <= not(layer2_outputs(3062));
    outputs(651) <= layer2_outputs(7285);
    outputs(652) <= layer2_outputs(10005);
    outputs(653) <= not(layer2_outputs(1680));
    outputs(654) <= (layer2_outputs(99)) and not (layer2_outputs(12496));
    outputs(655) <= layer2_outputs(2874);
    outputs(656) <= (layer2_outputs(9673)) or (layer2_outputs(5675));
    outputs(657) <= not((layer2_outputs(10030)) xor (layer2_outputs(3912)));
    outputs(658) <= (layer2_outputs(2266)) and not (layer2_outputs(5617));
    outputs(659) <= not(layer2_outputs(6849));
    outputs(660) <= not((layer2_outputs(6765)) xor (layer2_outputs(10803)));
    outputs(661) <= not(layer2_outputs(6575));
    outputs(662) <= not(layer2_outputs(5991));
    outputs(663) <= layer2_outputs(8316);
    outputs(664) <= not((layer2_outputs(8782)) or (layer2_outputs(935)));
    outputs(665) <= not(layer2_outputs(7828));
    outputs(666) <= layer2_outputs(3528);
    outputs(667) <= not((layer2_outputs(5286)) or (layer2_outputs(1095)));
    outputs(668) <= not(layer2_outputs(12763));
    outputs(669) <= not(layer2_outputs(2292));
    outputs(670) <= not((layer2_outputs(11437)) or (layer2_outputs(8018)));
    outputs(671) <= not((layer2_outputs(3882)) xor (layer2_outputs(4667)));
    outputs(672) <= layer2_outputs(3604);
    outputs(673) <= (layer2_outputs(10520)) xor (layer2_outputs(11259));
    outputs(674) <= not(layer2_outputs(6612));
    outputs(675) <= layer2_outputs(5799);
    outputs(676) <= layer2_outputs(8641);
    outputs(677) <= not(layer2_outputs(1956));
    outputs(678) <= layer2_outputs(3729);
    outputs(679) <= (layer2_outputs(5660)) and not (layer2_outputs(1053));
    outputs(680) <= not((layer2_outputs(3211)) xor (layer2_outputs(6985)));
    outputs(681) <= layer2_outputs(6283);
    outputs(682) <= not((layer2_outputs(7786)) and (layer2_outputs(10387)));
    outputs(683) <= not(layer2_outputs(5963));
    outputs(684) <= (layer2_outputs(9497)) and not (layer2_outputs(9741));
    outputs(685) <= (layer2_outputs(3674)) and not (layer2_outputs(12696));
    outputs(686) <= (layer2_outputs(7771)) or (layer2_outputs(1558));
    outputs(687) <= (layer2_outputs(11729)) and (layer2_outputs(7247));
    outputs(688) <= not(layer2_outputs(2147));
    outputs(689) <= layer2_outputs(2036);
    outputs(690) <= layer2_outputs(8006);
    outputs(691) <= layer2_outputs(12204);
    outputs(692) <= not((layer2_outputs(10553)) xor (layer2_outputs(3308)));
    outputs(693) <= not(layer2_outputs(5406));
    outputs(694) <= not(layer2_outputs(11552));
    outputs(695) <= not(layer2_outputs(379)) or (layer2_outputs(3536));
    outputs(696) <= not((layer2_outputs(3478)) or (layer2_outputs(8531)));
    outputs(697) <= not(layer2_outputs(927));
    outputs(698) <= not(layer2_outputs(8911));
    outputs(699) <= not(layer2_outputs(458));
    outputs(700) <= layer2_outputs(27);
    outputs(701) <= not((layer2_outputs(10209)) xor (layer2_outputs(3005)));
    outputs(702) <= layer2_outputs(4215);
    outputs(703) <= layer2_outputs(8029);
    outputs(704) <= not(layer2_outputs(3314));
    outputs(705) <= not(layer2_outputs(5188));
    outputs(706) <= not((layer2_outputs(9265)) xor (layer2_outputs(6379)));
    outputs(707) <= not(layer2_outputs(9231));
    outputs(708) <= not(layer2_outputs(12605));
    outputs(709) <= (layer2_outputs(4824)) xor (layer2_outputs(11559));
    outputs(710) <= not(layer2_outputs(3732));
    outputs(711) <= not((layer2_outputs(1581)) or (layer2_outputs(355)));
    outputs(712) <= (layer2_outputs(2062)) xor (layer2_outputs(4379));
    outputs(713) <= layer2_outputs(961);
    outputs(714) <= layer2_outputs(656);
    outputs(715) <= not(layer2_outputs(1966));
    outputs(716) <= not(layer2_outputs(12069));
    outputs(717) <= not((layer2_outputs(8462)) xor (layer2_outputs(6791)));
    outputs(718) <= not(layer2_outputs(7061));
    outputs(719) <= layer2_outputs(520);
    outputs(720) <= not((layer2_outputs(11218)) xor (layer2_outputs(153)));
    outputs(721) <= not((layer2_outputs(2853)) xor (layer2_outputs(3702)));
    outputs(722) <= layer2_outputs(8706);
    outputs(723) <= layer2_outputs(12213);
    outputs(724) <= (layer2_outputs(5974)) xor (layer2_outputs(4424));
    outputs(725) <= (layer2_outputs(10121)) and not (layer2_outputs(9816));
    outputs(726) <= (layer2_outputs(10746)) xor (layer2_outputs(4816));
    outputs(727) <= (layer2_outputs(5247)) xor (layer2_outputs(710));
    outputs(728) <= layer2_outputs(7234);
    outputs(729) <= layer2_outputs(11008);
    outputs(730) <= not(layer2_outputs(1277));
    outputs(731) <= not(layer2_outputs(12268));
    outputs(732) <= (layer2_outputs(10783)) or (layer2_outputs(364));
    outputs(733) <= not(layer2_outputs(3732));
    outputs(734) <= not(layer2_outputs(12106)) or (layer2_outputs(7294));
    outputs(735) <= not(layer2_outputs(3307));
    outputs(736) <= layer2_outputs(4695);
    outputs(737) <= not(layer2_outputs(2932));
    outputs(738) <= (layer2_outputs(6003)) or (layer2_outputs(7144));
    outputs(739) <= not((layer2_outputs(5574)) xor (layer2_outputs(3971)));
    outputs(740) <= layer2_outputs(5137);
    outputs(741) <= layer2_outputs(8929);
    outputs(742) <= layer2_outputs(5920);
    outputs(743) <= layer2_outputs(5704);
    outputs(744) <= layer2_outputs(10651);
    outputs(745) <= not(layer2_outputs(1682));
    outputs(746) <= not((layer2_outputs(8889)) xor (layer2_outputs(9100)));
    outputs(747) <= not(layer2_outputs(3564));
    outputs(748) <= not(layer2_outputs(2508));
    outputs(749) <= not(layer2_outputs(10970));
    outputs(750) <= not((layer2_outputs(8066)) and (layer2_outputs(4548)));
    outputs(751) <= layer2_outputs(2585);
    outputs(752) <= layer2_outputs(11465);
    outputs(753) <= (layer2_outputs(5621)) or (layer2_outputs(570));
    outputs(754) <= not((layer2_outputs(3255)) and (layer2_outputs(11993)));
    outputs(755) <= (layer2_outputs(10814)) and (layer2_outputs(9374));
    outputs(756) <= layer2_outputs(5149);
    outputs(757) <= layer2_outputs(9519);
    outputs(758) <= layer2_outputs(2860);
    outputs(759) <= (layer2_outputs(3709)) and not (layer2_outputs(1166));
    outputs(760) <= not(layer2_outputs(7850));
    outputs(761) <= layer2_outputs(4804);
    outputs(762) <= layer2_outputs(2998);
    outputs(763) <= (layer2_outputs(5477)) xor (layer2_outputs(1893));
    outputs(764) <= not((layer2_outputs(2010)) xor (layer2_outputs(3341)));
    outputs(765) <= (layer2_outputs(2460)) xor (layer2_outputs(6224));
    outputs(766) <= not(layer2_outputs(9201));
    outputs(767) <= layer2_outputs(8080);
    outputs(768) <= not(layer2_outputs(12607));
    outputs(769) <= (layer2_outputs(4026)) xor (layer2_outputs(8020));
    outputs(770) <= not((layer2_outputs(8735)) xor (layer2_outputs(7335)));
    outputs(771) <= (layer2_outputs(1850)) and not (layer2_outputs(6686));
    outputs(772) <= not((layer2_outputs(7180)) xor (layer2_outputs(7710)));
    outputs(773) <= layer2_outputs(9916);
    outputs(774) <= not(layer2_outputs(10976));
    outputs(775) <= (layer2_outputs(5682)) and not (layer2_outputs(1425));
    outputs(776) <= layer2_outputs(11629);
    outputs(777) <= layer2_outputs(9894);
    outputs(778) <= not(layer2_outputs(9355));
    outputs(779) <= not((layer2_outputs(10039)) xor (layer2_outputs(8888)));
    outputs(780) <= (layer2_outputs(12330)) and not (layer2_outputs(2943));
    outputs(781) <= (layer2_outputs(11867)) and (layer2_outputs(9863));
    outputs(782) <= not((layer2_outputs(8107)) xor (layer2_outputs(2047)));
    outputs(783) <= not((layer2_outputs(3952)) xor (layer2_outputs(4215)));
    outputs(784) <= not((layer2_outputs(7789)) xor (layer2_outputs(50)));
    outputs(785) <= not(layer2_outputs(205));
    outputs(786) <= not(layer2_outputs(11009)) or (layer2_outputs(9908));
    outputs(787) <= layer2_outputs(9046);
    outputs(788) <= not((layer2_outputs(8628)) xor (layer2_outputs(5002)));
    outputs(789) <= not(layer2_outputs(9587));
    outputs(790) <= not(layer2_outputs(11069)) or (layer2_outputs(10084));
    outputs(791) <= not(layer2_outputs(11189)) or (layer2_outputs(3638));
    outputs(792) <= (layer2_outputs(12307)) xor (layer2_outputs(2303));
    outputs(793) <= layer2_outputs(2998);
    outputs(794) <= (layer2_outputs(9272)) or (layer2_outputs(4860));
    outputs(795) <= (layer2_outputs(10703)) or (layer2_outputs(2243));
    outputs(796) <= not((layer2_outputs(2383)) or (layer2_outputs(7016)));
    outputs(797) <= not((layer2_outputs(3428)) xor (layer2_outputs(11846)));
    outputs(798) <= not(layer2_outputs(2503)) or (layer2_outputs(7528));
    outputs(799) <= (layer2_outputs(2624)) or (layer2_outputs(1285));
    outputs(800) <= layer2_outputs(1604);
    outputs(801) <= (layer2_outputs(2437)) or (layer2_outputs(12329));
    outputs(802) <= (layer2_outputs(4240)) or (layer2_outputs(1610));
    outputs(803) <= not(layer2_outputs(9992));
    outputs(804) <= layer2_outputs(11958);
    outputs(805) <= layer2_outputs(198);
    outputs(806) <= (layer2_outputs(6659)) xor (layer2_outputs(10010));
    outputs(807) <= not(layer2_outputs(12159));
    outputs(808) <= (layer2_outputs(6941)) xor (layer2_outputs(5366));
    outputs(809) <= (layer2_outputs(4120)) and (layer2_outputs(924));
    outputs(810) <= (layer2_outputs(8300)) and not (layer2_outputs(11254));
    outputs(811) <= not((layer2_outputs(11375)) xor (layer2_outputs(9569)));
    outputs(812) <= not(layer2_outputs(3711));
    outputs(813) <= (layer2_outputs(3285)) and not (layer2_outputs(6750));
    outputs(814) <= not((layer2_outputs(5364)) xor (layer2_outputs(12369)));
    outputs(815) <= (layer2_outputs(11777)) xor (layer2_outputs(11691));
    outputs(816) <= not((layer2_outputs(9131)) xor (layer2_outputs(10322)));
    outputs(817) <= layer2_outputs(8457);
    outputs(818) <= not(layer2_outputs(10373));
    outputs(819) <= (layer2_outputs(1559)) and not (layer2_outputs(3677));
    outputs(820) <= not(layer2_outputs(960));
    outputs(821) <= not(layer2_outputs(12178));
    outputs(822) <= not((layer2_outputs(2357)) xor (layer2_outputs(6666)));
    outputs(823) <= (layer2_outputs(9299)) xor (layer2_outputs(10033));
    outputs(824) <= layer2_outputs(1221);
    outputs(825) <= (layer2_outputs(3764)) xor (layer2_outputs(9247));
    outputs(826) <= (layer2_outputs(7745)) xor (layer2_outputs(3001));
    outputs(827) <= not((layer2_outputs(5635)) or (layer2_outputs(276)));
    outputs(828) <= (layer2_outputs(5402)) xor (layer2_outputs(8304));
    outputs(829) <= not(layer2_outputs(8207));
    outputs(830) <= not(layer2_outputs(2089));
    outputs(831) <= not(layer2_outputs(796));
    outputs(832) <= (layer2_outputs(8055)) xor (layer2_outputs(637));
    outputs(833) <= (layer2_outputs(6883)) and not (layer2_outputs(10565));
    outputs(834) <= (layer2_outputs(2449)) and not (layer2_outputs(1050));
    outputs(835) <= layer2_outputs(9290);
    outputs(836) <= not((layer2_outputs(3051)) xor (layer2_outputs(7481)));
    outputs(837) <= layer2_outputs(5213);
    outputs(838) <= not(layer2_outputs(12367));
    outputs(839) <= layer2_outputs(12223);
    outputs(840) <= layer2_outputs(12172);
    outputs(841) <= (layer2_outputs(2435)) xor (layer2_outputs(2058));
    outputs(842) <= layer2_outputs(7484);
    outputs(843) <= layer2_outputs(11942);
    outputs(844) <= not((layer2_outputs(5879)) or (layer2_outputs(11650)));
    outputs(845) <= layer2_outputs(1809);
    outputs(846) <= not(layer2_outputs(5688));
    outputs(847) <= (layer2_outputs(7645)) and not (layer2_outputs(6658));
    outputs(848) <= not(layer2_outputs(382));
    outputs(849) <= not((layer2_outputs(1930)) and (layer2_outputs(3575)));
    outputs(850) <= not(layer2_outputs(11448));
    outputs(851) <= not((layer2_outputs(2508)) xor (layer2_outputs(11104)));
    outputs(852) <= not(layer2_outputs(2094));
    outputs(853) <= not((layer2_outputs(2802)) xor (layer2_outputs(8225)));
    outputs(854) <= not(layer2_outputs(9864));
    outputs(855) <= layer2_outputs(2827);
    outputs(856) <= (layer2_outputs(9676)) and (layer2_outputs(8179));
    outputs(857) <= layer2_outputs(11388);
    outputs(858) <= not((layer2_outputs(10172)) xor (layer2_outputs(10151)));
    outputs(859) <= layer2_outputs(12204);
    outputs(860) <= layer2_outputs(3644);
    outputs(861) <= not(layer2_outputs(2946));
    outputs(862) <= not(layer2_outputs(3014));
    outputs(863) <= not(layer2_outputs(67));
    outputs(864) <= not(layer2_outputs(3228));
    outputs(865) <= not(layer2_outputs(5358));
    outputs(866) <= layer2_outputs(3489);
    outputs(867) <= not(layer2_outputs(1141));
    outputs(868) <= layer2_outputs(9190);
    outputs(869) <= (layer2_outputs(4519)) xor (layer2_outputs(11534));
    outputs(870) <= (layer2_outputs(10639)) xor (layer2_outputs(7247));
    outputs(871) <= not(layer2_outputs(896));
    outputs(872) <= layer2_outputs(9127);
    outputs(873) <= (layer2_outputs(4077)) xor (layer2_outputs(8781));
    outputs(874) <= not((layer2_outputs(1012)) xor (layer2_outputs(6481)));
    outputs(875) <= not((layer2_outputs(11342)) xor (layer2_outputs(2326)));
    outputs(876) <= layer2_outputs(1599);
    outputs(877) <= (layer2_outputs(234)) or (layer2_outputs(2767));
    outputs(878) <= layer2_outputs(3558);
    outputs(879) <= layer2_outputs(2562);
    outputs(880) <= not((layer2_outputs(7004)) xor (layer2_outputs(3685)));
    outputs(881) <= layer2_outputs(5953);
    outputs(882) <= not(layer2_outputs(809));
    outputs(883) <= layer2_outputs(11990);
    outputs(884) <= not(layer2_outputs(8136));
    outputs(885) <= not(layer2_outputs(11312));
    outputs(886) <= not(layer2_outputs(11122));
    outputs(887) <= layer2_outputs(8448);
    outputs(888) <= not((layer2_outputs(5201)) or (layer2_outputs(11377)));
    outputs(889) <= not((layer2_outputs(7345)) xor (layer2_outputs(1858)));
    outputs(890) <= not(layer2_outputs(3026));
    outputs(891) <= layer2_outputs(4294);
    outputs(892) <= not(layer2_outputs(8965));
    outputs(893) <= not((layer2_outputs(2500)) xor (layer2_outputs(8521)));
    outputs(894) <= not((layer2_outputs(12592)) xor (layer2_outputs(1376)));
    outputs(895) <= layer2_outputs(8241);
    outputs(896) <= (layer2_outputs(7430)) and not (layer2_outputs(4370));
    outputs(897) <= not((layer2_outputs(7183)) xor (layer2_outputs(9897)));
    outputs(898) <= layer2_outputs(7790);
    outputs(899) <= (layer2_outputs(6029)) xor (layer2_outputs(4930));
    outputs(900) <= (layer2_outputs(4822)) xor (layer2_outputs(1553));
    outputs(901) <= not((layer2_outputs(10347)) or (layer2_outputs(10846)));
    outputs(902) <= not(layer2_outputs(1134));
    outputs(903) <= (layer2_outputs(976)) xor (layer2_outputs(10098));
    outputs(904) <= layer2_outputs(6525);
    outputs(905) <= (layer2_outputs(11171)) xor (layer2_outputs(12123));
    outputs(906) <= layer2_outputs(137);
    outputs(907) <= not(layer2_outputs(291)) or (layer2_outputs(12274));
    outputs(908) <= not(layer2_outputs(11213));
    outputs(909) <= layer2_outputs(1926);
    outputs(910) <= layer2_outputs(3709);
    outputs(911) <= (layer2_outputs(550)) and (layer2_outputs(8515));
    outputs(912) <= not(layer2_outputs(7713));
    outputs(913) <= layer2_outputs(5140);
    outputs(914) <= (layer2_outputs(6085)) and (layer2_outputs(12489));
    outputs(915) <= not(layer2_outputs(5688));
    outputs(916) <= not((layer2_outputs(8497)) xor (layer2_outputs(7702)));
    outputs(917) <= (layer2_outputs(945)) xor (layer2_outputs(3579));
    outputs(918) <= layer2_outputs(8043);
    outputs(919) <= (layer2_outputs(12408)) and not (layer2_outputs(7914));
    outputs(920) <= not((layer2_outputs(10289)) and (layer2_outputs(1047)));
    outputs(921) <= not((layer2_outputs(7935)) xor (layer2_outputs(326)));
    outputs(922) <= not(layer2_outputs(8074)) or (layer2_outputs(10061));
    outputs(923) <= layer2_outputs(6710);
    outputs(924) <= not(layer2_outputs(9779));
    outputs(925) <= (layer2_outputs(3179)) and (layer2_outputs(9266));
    outputs(926) <= (layer2_outputs(8357)) and not (layer2_outputs(186));
    outputs(927) <= not(layer2_outputs(2049));
    outputs(928) <= (layer2_outputs(6139)) xor (layer2_outputs(8526));
    outputs(929) <= not(layer2_outputs(5647));
    outputs(930) <= layer2_outputs(4438);
    outputs(931) <= not(layer2_outputs(5539));
    outputs(932) <= not(layer2_outputs(7451)) or (layer2_outputs(890));
    outputs(933) <= layer2_outputs(8347);
    outputs(934) <= not(layer2_outputs(2297));
    outputs(935) <= (layer2_outputs(2221)) and not (layer2_outputs(3421));
    outputs(936) <= not((layer2_outputs(3987)) xor (layer2_outputs(9564)));
    outputs(937) <= (layer2_outputs(4823)) xor (layer2_outputs(5164));
    outputs(938) <= (layer2_outputs(1574)) xor (layer2_outputs(5420));
    outputs(939) <= (layer2_outputs(7046)) and not (layer2_outputs(10885));
    outputs(940) <= layer2_outputs(7217);
    outputs(941) <= layer2_outputs(12600);
    outputs(942) <= layer2_outputs(10670);
    outputs(943) <= (layer2_outputs(7303)) and (layer2_outputs(5480));
    outputs(944) <= not(layer2_outputs(1798));
    outputs(945) <= not((layer2_outputs(12494)) xor (layer2_outputs(11974)));
    outputs(946) <= layer2_outputs(10739);
    outputs(947) <= layer2_outputs(11637);
    outputs(948) <= layer2_outputs(11892);
    outputs(949) <= not((layer2_outputs(5759)) xor (layer2_outputs(11620)));
    outputs(950) <= layer2_outputs(4682);
    outputs(951) <= layer2_outputs(12056);
    outputs(952) <= not(layer2_outputs(3243)) or (layer2_outputs(1086));
    outputs(953) <= not(layer2_outputs(1918));
    outputs(954) <= (layer2_outputs(2870)) or (layer2_outputs(683));
    outputs(955) <= layer2_outputs(8295);
    outputs(956) <= (layer2_outputs(1584)) xor (layer2_outputs(3287));
    outputs(957) <= not(layer2_outputs(11102));
    outputs(958) <= not((layer2_outputs(8191)) and (layer2_outputs(5191)));
    outputs(959) <= not(layer2_outputs(35));
    outputs(960) <= not(layer2_outputs(7157)) or (layer2_outputs(7989));
    outputs(961) <= not(layer2_outputs(11079));
    outputs(962) <= layer2_outputs(1486);
    outputs(963) <= not((layer2_outputs(3603)) and (layer2_outputs(7836)));
    outputs(964) <= not(layer2_outputs(11617)) or (layer2_outputs(6466));
    outputs(965) <= not(layer2_outputs(1962));
    outputs(966) <= not(layer2_outputs(6060));
    outputs(967) <= not(layer2_outputs(11003));
    outputs(968) <= not((layer2_outputs(11160)) and (layer2_outputs(11677)));
    outputs(969) <= layer2_outputs(1637);
    outputs(970) <= not(layer2_outputs(8741));
    outputs(971) <= not(layer2_outputs(11102));
    outputs(972) <= layer2_outputs(9260);
    outputs(973) <= not(layer2_outputs(6484)) or (layer2_outputs(5231));
    outputs(974) <= layer2_outputs(3843);
    outputs(975) <= (layer2_outputs(7432)) xor (layer2_outputs(1251));
    outputs(976) <= not((layer2_outputs(5368)) xor (layer2_outputs(6841)));
    outputs(977) <= layer2_outputs(4209);
    outputs(978) <= (layer2_outputs(9197)) or (layer2_outputs(1344));
    outputs(979) <= layer2_outputs(7038);
    outputs(980) <= layer2_outputs(6380);
    outputs(981) <= not(layer2_outputs(7823));
    outputs(982) <= not(layer2_outputs(3958));
    outputs(983) <= layer2_outputs(4595);
    outputs(984) <= not(layer2_outputs(6754));
    outputs(985) <= not(layer2_outputs(6580));
    outputs(986) <= not(layer2_outputs(12565));
    outputs(987) <= (layer2_outputs(9698)) and (layer2_outputs(6364));
    outputs(988) <= not(layer2_outputs(1264));
    outputs(989) <= not(layer2_outputs(7112)) or (layer2_outputs(2894));
    outputs(990) <= layer2_outputs(11870);
    outputs(991) <= not(layer2_outputs(7092)) or (layer2_outputs(530));
    outputs(992) <= layer2_outputs(3984);
    outputs(993) <= (layer2_outputs(12021)) xor (layer2_outputs(8388));
    outputs(994) <= layer2_outputs(9785);
    outputs(995) <= layer2_outputs(9397);
    outputs(996) <= not((layer2_outputs(3555)) or (layer2_outputs(8045)));
    outputs(997) <= (layer2_outputs(2337)) xor (layer2_outputs(3968));
    outputs(998) <= (layer2_outputs(2010)) and (layer2_outputs(7122));
    outputs(999) <= layer2_outputs(11569);
    outputs(1000) <= (layer2_outputs(3666)) and not (layer2_outputs(3398));
    outputs(1001) <= layer2_outputs(4543);
    outputs(1002) <= not(layer2_outputs(352));
    outputs(1003) <= not(layer2_outputs(7840));
    outputs(1004) <= not(layer2_outputs(2350));
    outputs(1005) <= layer2_outputs(11154);
    outputs(1006) <= not(layer2_outputs(7562));
    outputs(1007) <= layer2_outputs(3569);
    outputs(1008) <= not(layer2_outputs(9876));
    outputs(1009) <= not(layer2_outputs(10975));
    outputs(1010) <= not((layer2_outputs(3370)) xor (layer2_outputs(12248)));
    outputs(1011) <= not(layer2_outputs(10745));
    outputs(1012) <= (layer2_outputs(11219)) or (layer2_outputs(11843));
    outputs(1013) <= layer2_outputs(4067);
    outputs(1014) <= layer2_outputs(1447);
    outputs(1015) <= layer2_outputs(213);
    outputs(1016) <= (layer2_outputs(7899)) and (layer2_outputs(10331));
    outputs(1017) <= not(layer2_outputs(8901));
    outputs(1018) <= not(layer2_outputs(5504));
    outputs(1019) <= not(layer2_outputs(416));
    outputs(1020) <= not(layer2_outputs(7740));
    outputs(1021) <= not(layer2_outputs(3627));
    outputs(1022) <= (layer2_outputs(7670)) xor (layer2_outputs(5090));
    outputs(1023) <= (layer2_outputs(3451)) or (layer2_outputs(9230));
    outputs(1024) <= not(layer2_outputs(11158));
    outputs(1025) <= layer2_outputs(6898);
    outputs(1026) <= not(layer2_outputs(12678));
    outputs(1027) <= layer2_outputs(7373);
    outputs(1028) <= not(layer2_outputs(11094));
    outputs(1029) <= layer2_outputs(12127);
    outputs(1030) <= (layer2_outputs(1333)) xor (layer2_outputs(1858));
    outputs(1031) <= (layer2_outputs(9410)) and not (layer2_outputs(7520));
    outputs(1032) <= not((layer2_outputs(7400)) xor (layer2_outputs(8245)));
    outputs(1033) <= layer2_outputs(12624);
    outputs(1034) <= not(layer2_outputs(4620));
    outputs(1035) <= layer2_outputs(1250);
    outputs(1036) <= layer2_outputs(1275);
    outputs(1037) <= not(layer2_outputs(12254));
    outputs(1038) <= not((layer2_outputs(316)) or (layer2_outputs(7820)));
    outputs(1039) <= (layer2_outputs(8972)) xor (layer2_outputs(11951));
    outputs(1040) <= not((layer2_outputs(5170)) or (layer2_outputs(3238)));
    outputs(1041) <= (layer2_outputs(5721)) or (layer2_outputs(7644));
    outputs(1042) <= layer2_outputs(9532);
    outputs(1043) <= (layer2_outputs(7291)) xor (layer2_outputs(11518));
    outputs(1044) <= not(layer2_outputs(11029)) or (layer2_outputs(10720));
    outputs(1045) <= not(layer2_outputs(9960));
    outputs(1046) <= not((layer2_outputs(4927)) xor (layer2_outputs(7282)));
    outputs(1047) <= not((layer2_outputs(2320)) xor (layer2_outputs(1975)));
    outputs(1048) <= not((layer2_outputs(3881)) xor (layer2_outputs(8380)));
    outputs(1049) <= layer2_outputs(8472);
    outputs(1050) <= not(layer2_outputs(124));
    outputs(1051) <= not(layer2_outputs(4369));
    outputs(1052) <= not(layer2_outputs(3121));
    outputs(1053) <= not(layer2_outputs(5245));
    outputs(1054) <= (layer2_outputs(769)) and not (layer2_outputs(12555));
    outputs(1055) <= not(layer2_outputs(6624));
    outputs(1056) <= not(layer2_outputs(9466));
    outputs(1057) <= (layer2_outputs(11882)) and not (layer2_outputs(5674));
    outputs(1058) <= not(layer2_outputs(7536));
    outputs(1059) <= not(layer2_outputs(7165));
    outputs(1060) <= not(layer2_outputs(10193));
    outputs(1061) <= not(layer2_outputs(3267));
    outputs(1062) <= layer2_outputs(10662);
    outputs(1063) <= (layer2_outputs(9136)) and not (layer2_outputs(777));
    outputs(1064) <= not(layer2_outputs(12719));
    outputs(1065) <= layer2_outputs(7527);
    outputs(1066) <= layer2_outputs(5763);
    outputs(1067) <= not((layer2_outputs(3873)) xor (layer2_outputs(12495)));
    outputs(1068) <= not((layer2_outputs(1524)) xor (layer2_outputs(6491)));
    outputs(1069) <= (layer2_outputs(9885)) xor (layer2_outputs(9846));
    outputs(1070) <= not(layer2_outputs(11403));
    outputs(1071) <= layer2_outputs(10336);
    outputs(1072) <= (layer2_outputs(9901)) and (layer2_outputs(5725));
    outputs(1073) <= layer2_outputs(6185);
    outputs(1074) <= not(layer2_outputs(12671));
    outputs(1075) <= not((layer2_outputs(11830)) xor (layer2_outputs(6735)));
    outputs(1076) <= not(layer2_outputs(2493));
    outputs(1077) <= (layer2_outputs(8572)) and (layer2_outputs(7236));
    outputs(1078) <= not((layer2_outputs(4415)) xor (layer2_outputs(7898)));
    outputs(1079) <= layer2_outputs(9762);
    outputs(1080) <= not((layer2_outputs(2762)) and (layer2_outputs(1304)));
    outputs(1081) <= not(layer2_outputs(7269)) or (layer2_outputs(11886));
    outputs(1082) <= layer2_outputs(12472);
    outputs(1083) <= layer2_outputs(3790);
    outputs(1084) <= layer2_outputs(5379);
    outputs(1085) <= not(layer2_outputs(1955));
    outputs(1086) <= not(layer2_outputs(8324)) or (layer2_outputs(1030));
    outputs(1087) <= (layer2_outputs(7073)) and (layer2_outputs(9824));
    outputs(1088) <= layer2_outputs(2201);
    outputs(1089) <= not((layer2_outputs(4132)) or (layer2_outputs(3425)));
    outputs(1090) <= layer2_outputs(12585);
    outputs(1091) <= layer2_outputs(5333);
    outputs(1092) <= (layer2_outputs(8922)) and not (layer2_outputs(7588));
    outputs(1093) <= (layer2_outputs(1593)) and (layer2_outputs(8477));
    outputs(1094) <= layer2_outputs(9862);
    outputs(1095) <= layer2_outputs(12301);
    outputs(1096) <= layer2_outputs(10002);
    outputs(1097) <= (layer2_outputs(5067)) and not (layer2_outputs(2715));
    outputs(1098) <= (layer2_outputs(2800)) xor (layer2_outputs(8391));
    outputs(1099) <= layer2_outputs(11829);
    outputs(1100) <= layer2_outputs(11880);
    outputs(1101) <= not((layer2_outputs(269)) or (layer2_outputs(4103)));
    outputs(1102) <= layer2_outputs(5251);
    outputs(1103) <= (layer2_outputs(5389)) xor (layer2_outputs(12052));
    outputs(1104) <= not(layer2_outputs(10748));
    outputs(1105) <= (layer2_outputs(3943)) and not (layer2_outputs(3089));
    outputs(1106) <= layer2_outputs(4251);
    outputs(1107) <= not(layer2_outputs(1857)) or (layer2_outputs(11411));
    outputs(1108) <= (layer2_outputs(6483)) and not (layer2_outputs(9143));
    outputs(1109) <= layer2_outputs(1025);
    outputs(1110) <= not((layer2_outputs(3753)) and (layer2_outputs(6455)));
    outputs(1111) <= (layer2_outputs(8185)) and not (layer2_outputs(3591));
    outputs(1112) <= (layer2_outputs(10872)) or (layer2_outputs(5744));
    outputs(1113) <= layer2_outputs(2420);
    outputs(1114) <= not((layer2_outputs(7951)) or (layer2_outputs(5208)));
    outputs(1115) <= layer2_outputs(4006);
    outputs(1116) <= layer2_outputs(828);
    outputs(1117) <= (layer2_outputs(5455)) and not (layer2_outputs(10457));
    outputs(1118) <= layer2_outputs(10134);
    outputs(1119) <= not(layer2_outputs(1270));
    outputs(1120) <= not((layer2_outputs(10904)) xor (layer2_outputs(10521)));
    outputs(1121) <= (layer2_outputs(2990)) xor (layer2_outputs(12399));
    outputs(1122) <= not((layer2_outputs(326)) xor (layer2_outputs(7123)));
    outputs(1123) <= not(layer2_outputs(4700));
    outputs(1124) <= not(layer2_outputs(10971));
    outputs(1125) <= not((layer2_outputs(2891)) xor (layer2_outputs(2687)));
    outputs(1126) <= not(layer2_outputs(12264));
    outputs(1127) <= not(layer2_outputs(5984));
    outputs(1128) <= layer2_outputs(225);
    outputs(1129) <= (layer2_outputs(4767)) and not (layer2_outputs(12548));
    outputs(1130) <= layer2_outputs(3146);
    outputs(1131) <= (layer2_outputs(3568)) and not (layer2_outputs(1882));
    outputs(1132) <= not(layer2_outputs(10924)) or (layer2_outputs(11228));
    outputs(1133) <= not(layer2_outputs(5159));
    outputs(1134) <= layer2_outputs(9385);
    outputs(1135) <= (layer2_outputs(6162)) and (layer2_outputs(5666));
    outputs(1136) <= layer2_outputs(12405);
    outputs(1137) <= layer2_outputs(5869);
    outputs(1138) <= layer2_outputs(8013);
    outputs(1139) <= (layer2_outputs(87)) and (layer2_outputs(7466));
    outputs(1140) <= not(layer2_outputs(4013));
    outputs(1141) <= (layer2_outputs(4120)) and not (layer2_outputs(10865));
    outputs(1142) <= not(layer2_outputs(1307));
    outputs(1143) <= not((layer2_outputs(10895)) xor (layer2_outputs(7949)));
    outputs(1144) <= layer2_outputs(10503);
    outputs(1145) <= not(layer2_outputs(4678)) or (layer2_outputs(5599));
    outputs(1146) <= (layer2_outputs(12317)) and not (layer2_outputs(951));
    outputs(1147) <= not(layer2_outputs(3842));
    outputs(1148) <= not((layer2_outputs(9738)) xor (layer2_outputs(6748)));
    outputs(1149) <= not(layer2_outputs(10441));
    outputs(1150) <= not(layer2_outputs(8182));
    outputs(1151) <= layer2_outputs(10278);
    outputs(1152) <= not(layer2_outputs(8423));
    outputs(1153) <= (layer2_outputs(5929)) and (layer2_outputs(11502));
    outputs(1154) <= layer2_outputs(9064);
    outputs(1155) <= layer2_outputs(9127);
    outputs(1156) <= not((layer2_outputs(6310)) xor (layer2_outputs(892)));
    outputs(1157) <= layer2_outputs(2427);
    outputs(1158) <= not(layer2_outputs(3712));
    outputs(1159) <= not(layer2_outputs(5182));
    outputs(1160) <= not((layer2_outputs(4347)) xor (layer2_outputs(11635)));
    outputs(1161) <= layer2_outputs(7503);
    outputs(1162) <= not((layer2_outputs(11121)) xor (layer2_outputs(915)));
    outputs(1163) <= (layer2_outputs(8991)) and not (layer2_outputs(10461));
    outputs(1164) <= not(layer2_outputs(5531)) or (layer2_outputs(9570));
    outputs(1165) <= not((layer2_outputs(11505)) xor (layer2_outputs(4653)));
    outputs(1166) <= layer2_outputs(4912);
    outputs(1167) <= not((layer2_outputs(6161)) xor (layer2_outputs(4245)));
    outputs(1168) <= layer2_outputs(9012);
    outputs(1169) <= not(layer2_outputs(4692));
    outputs(1170) <= not((layer2_outputs(2236)) and (layer2_outputs(7325)));
    outputs(1171) <= not((layer2_outputs(5621)) xor (layer2_outputs(9963)));
    outputs(1172) <= layer2_outputs(10217);
    outputs(1173) <= not(layer2_outputs(4546));
    outputs(1174) <= not((layer2_outputs(2567)) and (layer2_outputs(11944)));
    outputs(1175) <= not((layer2_outputs(5934)) xor (layer2_outputs(6328)));
    outputs(1176) <= not(layer2_outputs(7682)) or (layer2_outputs(1098));
    outputs(1177) <= (layer2_outputs(6314)) xor (layer2_outputs(374));
    outputs(1178) <= not(layer2_outputs(11321));
    outputs(1179) <= layer2_outputs(4107);
    outputs(1180) <= layer2_outputs(10102);
    outputs(1181) <= layer2_outputs(1903);
    outputs(1182) <= layer2_outputs(4138);
    outputs(1183) <= not(layer2_outputs(5580));
    outputs(1184) <= not(layer2_outputs(3654));
    outputs(1185) <= (layer2_outputs(289)) or (layer2_outputs(12015));
    outputs(1186) <= not(layer2_outputs(9210));
    outputs(1187) <= layer2_outputs(8687);
    outputs(1188) <= not(layer2_outputs(8412)) or (layer2_outputs(11876));
    outputs(1189) <= (layer2_outputs(611)) xor (layer2_outputs(1722));
    outputs(1190) <= (layer2_outputs(6845)) xor (layer2_outputs(3496));
    outputs(1191) <= not(layer2_outputs(5876));
    outputs(1192) <= (layer2_outputs(1314)) xor (layer2_outputs(3832));
    outputs(1193) <= layer2_outputs(8401);
    outputs(1194) <= not(layer2_outputs(6697));
    outputs(1195) <= layer2_outputs(9287);
    outputs(1196) <= layer2_outputs(4756);
    outputs(1197) <= not(layer2_outputs(8878));
    outputs(1198) <= not(layer2_outputs(7755));
    outputs(1199) <= (layer2_outputs(4329)) xor (layer2_outputs(11438));
    outputs(1200) <= not(layer2_outputs(12564));
    outputs(1201) <= not((layer2_outputs(7496)) xor (layer2_outputs(3848)));
    outputs(1202) <= not(layer2_outputs(7991));
    outputs(1203) <= not((layer2_outputs(9757)) xor (layer2_outputs(9829)));
    outputs(1204) <= not((layer2_outputs(1987)) and (layer2_outputs(8367)));
    outputs(1205) <= (layer2_outputs(9097)) xor (layer2_outputs(10202));
    outputs(1206) <= not(layer2_outputs(10984));
    outputs(1207) <= (layer2_outputs(5787)) and not (layer2_outputs(1696));
    outputs(1208) <= not(layer2_outputs(731));
    outputs(1209) <= not((layer2_outputs(8578)) xor (layer2_outputs(8864)));
    outputs(1210) <= layer2_outputs(12535);
    outputs(1211) <= layer2_outputs(6262);
    outputs(1212) <= layer2_outputs(4100);
    outputs(1213) <= not((layer2_outputs(2995)) xor (layer2_outputs(7931)));
    outputs(1214) <= not(layer2_outputs(4635));
    outputs(1215) <= not((layer2_outputs(7672)) or (layer2_outputs(1567)));
    outputs(1216) <= (layer2_outputs(4753)) and (layer2_outputs(3099));
    outputs(1217) <= layer2_outputs(2482);
    outputs(1218) <= layer2_outputs(1644);
    outputs(1219) <= not((layer2_outputs(3676)) xor (layer2_outputs(3503)));
    outputs(1220) <= (layer2_outputs(1839)) and (layer2_outputs(5475));
    outputs(1221) <= layer2_outputs(581);
    outputs(1222) <= (layer2_outputs(6277)) xor (layer2_outputs(9696));
    outputs(1223) <= layer2_outputs(6158);
    outputs(1224) <= not((layer2_outputs(2661)) xor (layer2_outputs(5334)));
    outputs(1225) <= not(layer2_outputs(2782));
    outputs(1226) <= not(layer2_outputs(5747)) or (layer2_outputs(4643));
    outputs(1227) <= layer2_outputs(3870);
    outputs(1228) <= layer2_outputs(11088);
    outputs(1229) <= not((layer2_outputs(1930)) and (layer2_outputs(3444)));
    outputs(1230) <= not((layer2_outputs(10363)) and (layer2_outputs(1924)));
    outputs(1231) <= not(layer2_outputs(3176)) or (layer2_outputs(9778));
    outputs(1232) <= layer2_outputs(2363);
    outputs(1233) <= not(layer2_outputs(8389)) or (layer2_outputs(11148));
    outputs(1234) <= not(layer2_outputs(6984));
    outputs(1235) <= not(layer2_outputs(3390));
    outputs(1236) <= not(layer2_outputs(8095)) or (layer2_outputs(3058));
    outputs(1237) <= (layer2_outputs(2839)) and not (layer2_outputs(6982));
    outputs(1238) <= (layer2_outputs(28)) xor (layer2_outputs(7689));
    outputs(1239) <= (layer2_outputs(8004)) xor (layer2_outputs(7559));
    outputs(1240) <= not(layer2_outputs(9619));
    outputs(1241) <= (layer2_outputs(2787)) and (layer2_outputs(7721));
    outputs(1242) <= not(layer2_outputs(3196));
    outputs(1243) <= not(layer2_outputs(3301));
    outputs(1244) <= (layer2_outputs(11596)) xor (layer2_outputs(4757));
    outputs(1245) <= not(layer2_outputs(12155));
    outputs(1246) <= not((layer2_outputs(9921)) xor (layer2_outputs(84)));
    outputs(1247) <= (layer2_outputs(11531)) and (layer2_outputs(10452));
    outputs(1248) <= layer2_outputs(2742);
    outputs(1249) <= not(layer2_outputs(4388)) or (layer2_outputs(6798));
    outputs(1250) <= not(layer2_outputs(10342)) or (layer2_outputs(2090));
    outputs(1251) <= not((layer2_outputs(6630)) xor (layer2_outputs(11429)));
    outputs(1252) <= not(layer2_outputs(8282));
    outputs(1253) <= (layer2_outputs(10900)) xor (layer2_outputs(3353));
    outputs(1254) <= not(layer2_outputs(8234));
    outputs(1255) <= not(layer2_outputs(3822)) or (layer2_outputs(3384));
    outputs(1256) <= not((layer2_outputs(9503)) or (layer2_outputs(5944)));
    outputs(1257) <= not(layer2_outputs(1786));
    outputs(1258) <= (layer2_outputs(7831)) or (layer2_outputs(696));
    outputs(1259) <= layer2_outputs(7735);
    outputs(1260) <= not(layer2_outputs(9406));
    outputs(1261) <= (layer2_outputs(5853)) xor (layer2_outputs(8442));
    outputs(1262) <= (layer2_outputs(11067)) or (layer2_outputs(8498));
    outputs(1263) <= not(layer2_outputs(1255));
    outputs(1264) <= not((layer2_outputs(8817)) xor (layer2_outputs(357)));
    outputs(1265) <= not(layer2_outputs(1883));
    outputs(1266) <= not((layer2_outputs(10728)) xor (layer2_outputs(11787)));
    outputs(1267) <= (layer2_outputs(3566)) or (layer2_outputs(2074));
    outputs(1268) <= not(layer2_outputs(10514));
    outputs(1269) <= not(layer2_outputs(4088));
    outputs(1270) <= (layer2_outputs(4501)) and not (layer2_outputs(12729));
    outputs(1271) <= (layer2_outputs(11957)) and not (layer2_outputs(11216));
    outputs(1272) <= not(layer2_outputs(9481)) or (layer2_outputs(8164));
    outputs(1273) <= not((layer2_outputs(2829)) xor (layer2_outputs(3634)));
    outputs(1274) <= not(layer2_outputs(5423));
    outputs(1275) <= (layer2_outputs(9823)) and (layer2_outputs(1709));
    outputs(1276) <= not(layer2_outputs(1986));
    outputs(1277) <= not(layer2_outputs(2903));
    outputs(1278) <= layer2_outputs(10630);
    outputs(1279) <= (layer2_outputs(7641)) xor (layer2_outputs(701));
    outputs(1280) <= (layer2_outputs(1851)) xor (layer2_outputs(4266));
    outputs(1281) <= not((layer2_outputs(7225)) or (layer2_outputs(8351)));
    outputs(1282) <= (layer2_outputs(11478)) and not (layer2_outputs(10389));
    outputs(1283) <= not(layer2_outputs(178));
    outputs(1284) <= (layer2_outputs(3265)) and not (layer2_outputs(2368));
    outputs(1285) <= not((layer2_outputs(2323)) xor (layer2_outputs(10024)));
    outputs(1286) <= layer2_outputs(147);
    outputs(1287) <= layer2_outputs(11618);
    outputs(1288) <= (layer2_outputs(5616)) and (layer2_outputs(11786));
    outputs(1289) <= layer2_outputs(7609);
    outputs(1290) <= (layer2_outputs(5733)) and not (layer2_outputs(9521));
    outputs(1291) <= not(layer2_outputs(10707));
    outputs(1292) <= not(layer2_outputs(6407));
    outputs(1293) <= not((layer2_outputs(2784)) xor (layer2_outputs(7913)));
    outputs(1294) <= (layer2_outputs(7777)) xor (layer2_outputs(8181));
    outputs(1295) <= layer2_outputs(2953);
    outputs(1296) <= layer2_outputs(10489);
    outputs(1297) <= not((layer2_outputs(7930)) xor (layer2_outputs(541)));
    outputs(1298) <= (layer2_outputs(4372)) and (layer2_outputs(11422));
    outputs(1299) <= (layer2_outputs(12659)) and not (layer2_outputs(234));
    outputs(1300) <= (layer2_outputs(1478)) xor (layer2_outputs(107));
    outputs(1301) <= not((layer2_outputs(5447)) xor (layer2_outputs(4778)));
    outputs(1302) <= not((layer2_outputs(11396)) xor (layer2_outputs(7950)));
    outputs(1303) <= not((layer2_outputs(7126)) xor (layer2_outputs(12217)));
    outputs(1304) <= not((layer2_outputs(8065)) or (layer2_outputs(5805)));
    outputs(1305) <= not((layer2_outputs(3053)) or (layer2_outputs(2720)));
    outputs(1306) <= not((layer2_outputs(8671)) xor (layer2_outputs(10251)));
    outputs(1307) <= not((layer2_outputs(8123)) or (layer2_outputs(5312)));
    outputs(1308) <= not(layer2_outputs(9965));
    outputs(1309) <= layer2_outputs(1810);
    outputs(1310) <= layer2_outputs(12781);
    outputs(1311) <= (layer2_outputs(8192)) and not (layer2_outputs(8048));
    outputs(1312) <= not(layer2_outputs(910));
    outputs(1313) <= (layer2_outputs(6842)) xor (layer2_outputs(5629));
    outputs(1314) <= not((layer2_outputs(11238)) xor (layer2_outputs(12138)));
    outputs(1315) <= not((layer2_outputs(5677)) xor (layer2_outputs(6067)));
    outputs(1316) <= not((layer2_outputs(417)) xor (layer2_outputs(11866)));
    outputs(1317) <= (layer2_outputs(9008)) xor (layer2_outputs(7458));
    outputs(1318) <= layer2_outputs(5862);
    outputs(1319) <= not((layer2_outputs(12642)) and (layer2_outputs(3503)));
    outputs(1320) <= not(layer2_outputs(1462)) or (layer2_outputs(5632));
    outputs(1321) <= (layer2_outputs(10450)) and (layer2_outputs(6445));
    outputs(1322) <= layer2_outputs(9362);
    outputs(1323) <= not((layer2_outputs(2236)) xor (layer2_outputs(4295)));
    outputs(1324) <= (layer2_outputs(7539)) and (layer2_outputs(7610));
    outputs(1325) <= (layer2_outputs(686)) xor (layer2_outputs(12701));
    outputs(1326) <= not((layer2_outputs(4566)) and (layer2_outputs(969)));
    outputs(1327) <= (layer2_outputs(5175)) and not (layer2_outputs(10750));
    outputs(1328) <= not(layer2_outputs(8990));
    outputs(1329) <= layer2_outputs(12505);
    outputs(1330) <= (layer2_outputs(9212)) xor (layer2_outputs(12497));
    outputs(1331) <= not((layer2_outputs(5109)) and (layer2_outputs(9371)));
    outputs(1332) <= not(layer2_outputs(8870));
    outputs(1333) <= not((layer2_outputs(7606)) xor (layer2_outputs(10649)));
    outputs(1334) <= not(layer2_outputs(3275));
    outputs(1335) <= (layer2_outputs(1232)) and not (layer2_outputs(2434));
    outputs(1336) <= not(layer2_outputs(2735));
    outputs(1337) <= not(layer2_outputs(734));
    outputs(1338) <= not(layer2_outputs(9622));
    outputs(1339) <= not((layer2_outputs(10624)) xor (layer2_outputs(12711)));
    outputs(1340) <= not(layer2_outputs(6347));
    outputs(1341) <= (layer2_outputs(8242)) and not (layer2_outputs(3593));
    outputs(1342) <= not((layer2_outputs(9024)) or (layer2_outputs(1183)));
    outputs(1343) <= not((layer2_outputs(7431)) xor (layer2_outputs(4913)));
    outputs(1344) <= not(layer2_outputs(7044));
    outputs(1345) <= not((layer2_outputs(3633)) xor (layer2_outputs(9460)));
    outputs(1346) <= layer2_outputs(5421);
    outputs(1347) <= layer2_outputs(5365);
    outputs(1348) <= layer2_outputs(2627);
    outputs(1349) <= layer2_outputs(12734);
    outputs(1350) <= layer2_outputs(10862);
    outputs(1351) <= (layer2_outputs(12188)) xor (layer2_outputs(12582));
    outputs(1352) <= layer2_outputs(6773);
    outputs(1353) <= (layer2_outputs(3517)) xor (layer2_outputs(2501));
    outputs(1354) <= not(layer2_outputs(3181));
    outputs(1355) <= (layer2_outputs(11476)) xor (layer2_outputs(4779));
    outputs(1356) <= layer2_outputs(4180);
    outputs(1357) <= not((layer2_outputs(5933)) or (layer2_outputs(8603)));
    outputs(1358) <= not(layer2_outputs(7290)) or (layer2_outputs(8774));
    outputs(1359) <= not(layer2_outputs(10750));
    outputs(1360) <= (layer2_outputs(6774)) and (layer2_outputs(1814));
    outputs(1361) <= (layer2_outputs(1758)) xor (layer2_outputs(4856));
    outputs(1362) <= not(layer2_outputs(8563)) or (layer2_outputs(1030));
    outputs(1363) <= not((layer2_outputs(451)) or (layer2_outputs(8054)));
    outputs(1364) <= not(layer2_outputs(2451));
    outputs(1365) <= not((layer2_outputs(5411)) or (layer2_outputs(5755)));
    outputs(1366) <= (layer2_outputs(9361)) and not (layer2_outputs(5681));
    outputs(1367) <= layer2_outputs(4013);
    outputs(1368) <= not((layer2_outputs(6389)) or (layer2_outputs(4532)));
    outputs(1369) <= (layer2_outputs(7147)) and not (layer2_outputs(11569));
    outputs(1370) <= (layer2_outputs(6411)) and not (layer2_outputs(5503));
    outputs(1371) <= layer2_outputs(11113);
    outputs(1372) <= not((layer2_outputs(10839)) xor (layer2_outputs(6088)));
    outputs(1373) <= layer2_outputs(3078);
    outputs(1374) <= not((layer2_outputs(7615)) xor (layer2_outputs(5082)));
    outputs(1375) <= (layer2_outputs(5695)) and not (layer2_outputs(7557));
    outputs(1376) <= not((layer2_outputs(9446)) xor (layer2_outputs(6544)));
    outputs(1377) <= (layer2_outputs(8736)) or (layer2_outputs(2208));
    outputs(1378) <= not((layer2_outputs(4312)) xor (layer2_outputs(1444)));
    outputs(1379) <= not((layer2_outputs(3523)) or (layer2_outputs(5103)));
    outputs(1380) <= (layer2_outputs(6671)) and not (layer2_outputs(1507));
    outputs(1381) <= layer2_outputs(159);
    outputs(1382) <= (layer2_outputs(5601)) xor (layer2_outputs(1361));
    outputs(1383) <= not(layer2_outputs(11973));
    outputs(1384) <= (layer2_outputs(11295)) xor (layer2_outputs(9103));
    outputs(1385) <= (layer2_outputs(137)) xor (layer2_outputs(10185));
    outputs(1386) <= not((layer2_outputs(7350)) xor (layer2_outputs(10104)));
    outputs(1387) <= not(layer2_outputs(4424));
    outputs(1388) <= not((layer2_outputs(1015)) xor (layer2_outputs(9009)));
    outputs(1389) <= not(layer2_outputs(6649));
    outputs(1390) <= not((layer2_outputs(1833)) and (layer2_outputs(6345)));
    outputs(1391) <= not((layer2_outputs(7103)) or (layer2_outputs(1261)));
    outputs(1392) <= not(layer2_outputs(5174));
    outputs(1393) <= (layer2_outputs(10874)) and (layer2_outputs(5985));
    outputs(1394) <= (layer2_outputs(7619)) xor (layer2_outputs(5363));
    outputs(1395) <= not((layer2_outputs(11589)) xor (layer2_outputs(6663)));
    outputs(1396) <= not(layer2_outputs(11698));
    outputs(1397) <= (layer2_outputs(4904)) and not (layer2_outputs(2420));
    outputs(1398) <= layer2_outputs(11179);
    outputs(1399) <= not((layer2_outputs(9834)) xor (layer2_outputs(569)));
    outputs(1400) <= (layer2_outputs(9651)) and (layer2_outputs(56));
    outputs(1401) <= layer2_outputs(5302);
    outputs(1402) <= not(layer2_outputs(10549)) or (layer2_outputs(10833));
    outputs(1403) <= not(layer2_outputs(12542));
    outputs(1404) <= not(layer2_outputs(6910));
    outputs(1405) <= (layer2_outputs(5911)) and not (layer2_outputs(7086));
    outputs(1406) <= not((layer2_outputs(10315)) xor (layer2_outputs(10816)));
    outputs(1407) <= layer2_outputs(2224);
    outputs(1408) <= not((layer2_outputs(10180)) xor (layer2_outputs(2660)));
    outputs(1409) <= (layer2_outputs(8695)) and not (layer2_outputs(9348));
    outputs(1410) <= not(layer2_outputs(8011));
    outputs(1411) <= layer2_outputs(6534);
    outputs(1412) <= not((layer2_outputs(1306)) xor (layer2_outputs(5986)));
    outputs(1413) <= not(layer2_outputs(2059));
    outputs(1414) <= not(layer2_outputs(8624)) or (layer2_outputs(2286));
    outputs(1415) <= not(layer2_outputs(11198));
    outputs(1416) <= (layer2_outputs(7076)) and (layer2_outputs(11217));
    outputs(1417) <= not((layer2_outputs(3158)) and (layer2_outputs(914)));
    outputs(1418) <= layer2_outputs(11052);
    outputs(1419) <= (layer2_outputs(5634)) and not (layer2_outputs(748));
    outputs(1420) <= not((layer2_outputs(7874)) and (layer2_outputs(10951)));
    outputs(1421) <= not((layer2_outputs(2840)) xor (layer2_outputs(1790)));
    outputs(1422) <= not(layer2_outputs(2025));
    outputs(1423) <= (layer2_outputs(1273)) and not (layer2_outputs(334));
    outputs(1424) <= (layer2_outputs(2184)) xor (layer2_outputs(2231));
    outputs(1425) <= not(layer2_outputs(4852));
    outputs(1426) <= (layer2_outputs(11879)) and not (layer2_outputs(4014));
    outputs(1427) <= not((layer2_outputs(11735)) or (layer2_outputs(8770)));
    outputs(1428) <= not((layer2_outputs(6059)) or (layer2_outputs(10419)));
    outputs(1429) <= (layer2_outputs(7105)) xor (layer2_outputs(4585));
    outputs(1430) <= not(layer2_outputs(11160));
    outputs(1431) <= layer2_outputs(3667);
    outputs(1432) <= not((layer2_outputs(20)) xor (layer2_outputs(1331)));
    outputs(1433) <= not(layer2_outputs(4042)) or (layer2_outputs(9842));
    outputs(1434) <= (layer2_outputs(10319)) xor (layer2_outputs(5335));
    outputs(1435) <= layer2_outputs(4077);
    outputs(1436) <= (layer2_outputs(12001)) and (layer2_outputs(3280));
    outputs(1437) <= layer2_outputs(6693);
    outputs(1438) <= (layer2_outputs(10045)) and not (layer2_outputs(3999));
    outputs(1439) <= (layer2_outputs(10966)) xor (layer2_outputs(8748));
    outputs(1440) <= not((layer2_outputs(9420)) or (layer2_outputs(3033)));
    outputs(1441) <= (layer2_outputs(5119)) and not (layer2_outputs(1564));
    outputs(1442) <= layer2_outputs(2876);
    outputs(1443) <= layer2_outputs(3977);
    outputs(1444) <= layer2_outputs(9656);
    outputs(1445) <= layer2_outputs(5823);
    outputs(1446) <= (layer2_outputs(10960)) and not (layer2_outputs(11313));
    outputs(1447) <= (layer2_outputs(9558)) and not (layer2_outputs(58));
    outputs(1448) <= layer2_outputs(5541);
    outputs(1449) <= (layer2_outputs(8217)) xor (layer2_outputs(11168));
    outputs(1450) <= (layer2_outputs(11922)) xor (layer2_outputs(8885));
    outputs(1451) <= (layer2_outputs(12085)) and not (layer2_outputs(4322));
    outputs(1452) <= not(layer2_outputs(4886));
    outputs(1453) <= not((layer2_outputs(5006)) xor (layer2_outputs(12009)));
    outputs(1454) <= (layer2_outputs(4071)) xor (layer2_outputs(5265));
    outputs(1455) <= not(layer2_outputs(1691));
    outputs(1456) <= (layer2_outputs(11733)) or (layer2_outputs(3263));
    outputs(1457) <= layer2_outputs(1560);
    outputs(1458) <= (layer2_outputs(5372)) xor (layer2_outputs(5740));
    outputs(1459) <= (layer2_outputs(3343)) xor (layer2_outputs(9128));
    outputs(1460) <= (layer2_outputs(10147)) xor (layer2_outputs(12067));
    outputs(1461) <= (layer2_outputs(2614)) and not (layer2_outputs(3599));
    outputs(1462) <= (layer2_outputs(9681)) and (layer2_outputs(8608));
    outputs(1463) <= (layer2_outputs(8671)) and (layer2_outputs(5428));
    outputs(1464) <= not((layer2_outputs(6421)) xor (layer2_outputs(9947)));
    outputs(1465) <= not((layer2_outputs(7860)) xor (layer2_outputs(1936)));
    outputs(1466) <= not(layer2_outputs(12528));
    outputs(1467) <= not((layer2_outputs(11280)) or (layer2_outputs(10778)));
    outputs(1468) <= (layer2_outputs(2960)) xor (layer2_outputs(12082));
    outputs(1469) <= (layer2_outputs(10152)) xor (layer2_outputs(9195));
    outputs(1470) <= not(layer2_outputs(3170));
    outputs(1471) <= not((layer2_outputs(7877)) xor (layer2_outputs(2752)));
    outputs(1472) <= not(layer2_outputs(2506));
    outputs(1473) <= not(layer2_outputs(1103));
    outputs(1474) <= not((layer2_outputs(8989)) or (layer2_outputs(4291)));
    outputs(1475) <= (layer2_outputs(958)) and not (layer2_outputs(801));
    outputs(1476) <= not((layer2_outputs(10713)) xor (layer2_outputs(288)));
    outputs(1477) <= not((layer2_outputs(3227)) xor (layer2_outputs(255)));
    outputs(1478) <= (layer2_outputs(9758)) and (layer2_outputs(12087));
    outputs(1479) <= (layer2_outputs(3754)) and (layer2_outputs(9858));
    outputs(1480) <= not((layer2_outputs(12207)) xor (layer2_outputs(8074)));
    outputs(1481) <= not((layer2_outputs(459)) xor (layer2_outputs(6955)));
    outputs(1482) <= (layer2_outputs(7155)) xor (layer2_outputs(7818));
    outputs(1483) <= not((layer2_outputs(8571)) xor (layer2_outputs(9926)));
    outputs(1484) <= not((layer2_outputs(3129)) xor (layer2_outputs(9228)));
    outputs(1485) <= not(layer2_outputs(11905));
    outputs(1486) <= layer2_outputs(9845);
    outputs(1487) <= '0';
    outputs(1488) <= (layer2_outputs(8354)) xor (layer2_outputs(5639));
    outputs(1489) <= layer2_outputs(12461);
    outputs(1490) <= (layer2_outputs(3805)) and not (layer2_outputs(8469));
    outputs(1491) <= (layer2_outputs(2572)) and not (layer2_outputs(11485));
    outputs(1492) <= layer2_outputs(3019);
    outputs(1493) <= (layer2_outputs(8211)) and not (layer2_outputs(10258));
    outputs(1494) <= layer2_outputs(6145);
    outputs(1495) <= (layer2_outputs(5309)) and not (layer2_outputs(149));
    outputs(1496) <= not(layer2_outputs(3382));
    outputs(1497) <= (layer2_outputs(2654)) xor (layer2_outputs(689));
    outputs(1498) <= not(layer2_outputs(8768));
    outputs(1499) <= not(layer2_outputs(9368));
    outputs(1500) <= layer2_outputs(8929);
    outputs(1501) <= not((layer2_outputs(323)) and (layer2_outputs(2159)));
    outputs(1502) <= (layer2_outputs(11361)) and not (layer2_outputs(5815));
    outputs(1503) <= (layer2_outputs(9016)) or (layer2_outputs(4896));
    outputs(1504) <= not(layer2_outputs(3322));
    outputs(1505) <= not((layer2_outputs(11591)) or (layer2_outputs(5638)));
    outputs(1506) <= layer2_outputs(221);
    outputs(1507) <= (layer2_outputs(7343)) and not (layer2_outputs(290));
    outputs(1508) <= not((layer2_outputs(1230)) xor (layer2_outputs(10425)));
    outputs(1509) <= (layer2_outputs(8987)) xor (layer2_outputs(2459));
    outputs(1510) <= not(layer2_outputs(698));
    outputs(1511) <= (layer2_outputs(6963)) xor (layer2_outputs(12778));
    outputs(1512) <= not(layer2_outputs(11174));
    outputs(1513) <= not(layer2_outputs(3717));
    outputs(1514) <= layer2_outputs(4665);
    outputs(1515) <= layer2_outputs(8503);
    outputs(1516) <= not((layer2_outputs(6611)) or (layer2_outputs(8117)));
    outputs(1517) <= layer2_outputs(874);
    outputs(1518) <= layer2_outputs(4942);
    outputs(1519) <= not((layer2_outputs(5731)) or (layer2_outputs(3875)));
    outputs(1520) <= (layer2_outputs(6096)) and not (layer2_outputs(11815));
    outputs(1521) <= not((layer2_outputs(4409)) xor (layer2_outputs(6541)));
    outputs(1522) <= not(layer2_outputs(3715));
    outputs(1523) <= not(layer2_outputs(5831));
    outputs(1524) <= layer2_outputs(4471);
    outputs(1525) <= (layer2_outputs(1358)) or (layer2_outputs(10933));
    outputs(1526) <= (layer2_outputs(1971)) and (layer2_outputs(10740));
    outputs(1527) <= (layer2_outputs(12745)) xor (layer2_outputs(7561));
    outputs(1528) <= not(layer2_outputs(5703));
    outputs(1529) <= not((layer2_outputs(5429)) xor (layer2_outputs(7653)));
    outputs(1530) <= not((layer2_outputs(1611)) xor (layer2_outputs(8937)));
    outputs(1531) <= not(layer2_outputs(8205));
    outputs(1532) <= not((layer2_outputs(8405)) xor (layer2_outputs(962)));
    outputs(1533) <= layer2_outputs(7601);
    outputs(1534) <= not((layer2_outputs(5893)) xor (layer2_outputs(4681)));
    outputs(1535) <= (layer2_outputs(7202)) xor (layer2_outputs(2015));
    outputs(1536) <= (layer2_outputs(2024)) and not (layer2_outputs(2343));
    outputs(1537) <= layer2_outputs(12662);
    outputs(1538) <= not((layer2_outputs(653)) xor (layer2_outputs(6650)));
    outputs(1539) <= (layer2_outputs(7057)) and not (layer2_outputs(5010));
    outputs(1540) <= layer2_outputs(9866);
    outputs(1541) <= not((layer2_outputs(6384)) xor (layer2_outputs(8138)));
    outputs(1542) <= layer2_outputs(3043);
    outputs(1543) <= not((layer2_outputs(2524)) or (layer2_outputs(9542)));
    outputs(1544) <= not(layer2_outputs(11290));
    outputs(1545) <= not((layer2_outputs(9606)) xor (layer2_outputs(1514)));
    outputs(1546) <= not((layer2_outputs(4257)) xor (layer2_outputs(10936)));
    outputs(1547) <= layer2_outputs(6780);
    outputs(1548) <= (layer2_outputs(7317)) and not (layer2_outputs(12129));
    outputs(1549) <= not((layer2_outputs(4404)) xor (layer2_outputs(11117)));
    outputs(1550) <= (layer2_outputs(2871)) and not (layer2_outputs(523));
    outputs(1551) <= layer2_outputs(312);
    outputs(1552) <= (layer2_outputs(12297)) xor (layer2_outputs(2768));
    outputs(1553) <= (layer2_outputs(3692)) or (layer2_outputs(2520));
    outputs(1554) <= layer2_outputs(10054);
    outputs(1555) <= (layer2_outputs(7720)) xor (layer2_outputs(11798));
    outputs(1556) <= (layer2_outputs(9259)) and not (layer2_outputs(7809));
    outputs(1557) <= (layer2_outputs(11121)) and not (layer2_outputs(1541));
    outputs(1558) <= not(layer2_outputs(10327));
    outputs(1559) <= layer2_outputs(11636);
    outputs(1560) <= not(layer2_outputs(4676));
    outputs(1561) <= (layer2_outputs(1023)) and not (layer2_outputs(9806));
    outputs(1562) <= not((layer2_outputs(901)) xor (layer2_outputs(1803)));
    outputs(1563) <= not(layer2_outputs(1754));
    outputs(1564) <= (layer2_outputs(3859)) and not (layer2_outputs(821));
    outputs(1565) <= layer2_outputs(2503);
    outputs(1566) <= not(layer2_outputs(5025));
    outputs(1567) <= not(layer2_outputs(1926));
    outputs(1568) <= (layer2_outputs(12212)) xor (layer2_outputs(8704));
    outputs(1569) <= (layer2_outputs(5084)) and not (layer2_outputs(11751));
    outputs(1570) <= not(layer2_outputs(4945)) or (layer2_outputs(12325));
    outputs(1571) <= (layer2_outputs(3870)) and not (layer2_outputs(2197));
    outputs(1572) <= (layer2_outputs(1683)) and (layer2_outputs(3809));
    outputs(1573) <= layer2_outputs(4302);
    outputs(1574) <= layer2_outputs(44);
    outputs(1575) <= (layer2_outputs(4213)) and (layer2_outputs(9718));
    outputs(1576) <= (layer2_outputs(3947)) or (layer2_outputs(6266));
    outputs(1577) <= not(layer2_outputs(1944));
    outputs(1578) <= (layer2_outputs(6486)) and (layer2_outputs(1706));
    outputs(1579) <= not((layer2_outputs(9938)) or (layer2_outputs(161)));
    outputs(1580) <= not(layer2_outputs(4878));
    outputs(1581) <= not((layer2_outputs(9791)) xor (layer2_outputs(12272)));
    outputs(1582) <= (layer2_outputs(8546)) xor (layer2_outputs(5055));
    outputs(1583) <= not(layer2_outputs(1906));
    outputs(1584) <= not(layer2_outputs(945));
    outputs(1585) <= not(layer2_outputs(1895));
    outputs(1586) <= (layer2_outputs(11112)) or (layer2_outputs(5818));
    outputs(1587) <= not((layer2_outputs(8089)) xor (layer2_outputs(67)));
    outputs(1588) <= not(layer2_outputs(4566));
    outputs(1589) <= not(layer2_outputs(4722));
    outputs(1590) <= not((layer2_outputs(4176)) xor (layer2_outputs(1783)));
    outputs(1591) <= (layer2_outputs(7616)) and not (layer2_outputs(9827));
    outputs(1592) <= layer2_outputs(4796);
    outputs(1593) <= not(layer2_outputs(8821));
    outputs(1594) <= layer2_outputs(12002);
    outputs(1595) <= layer2_outputs(7209);
    outputs(1596) <= not((layer2_outputs(10138)) xor (layer2_outputs(3112)));
    outputs(1597) <= not(layer2_outputs(2578));
    outputs(1598) <= not((layer2_outputs(109)) xor (layer2_outputs(10320)));
    outputs(1599) <= layer2_outputs(10453);
    outputs(1600) <= not((layer2_outputs(5413)) or (layer2_outputs(8536)));
    outputs(1601) <= layer2_outputs(9501);
    outputs(1602) <= (layer2_outputs(3068)) or (layer2_outputs(4718));
    outputs(1603) <= layer2_outputs(3782);
    outputs(1604) <= not(layer2_outputs(2342));
    outputs(1605) <= not(layer2_outputs(2403));
    outputs(1606) <= (layer2_outputs(9528)) and (layer2_outputs(53));
    outputs(1607) <= layer2_outputs(12324);
    outputs(1608) <= not(layer2_outputs(6356));
    outputs(1609) <= not((layer2_outputs(9393)) or (layer2_outputs(3832)));
    outputs(1610) <= not(layer2_outputs(11769));
    outputs(1611) <= not(layer2_outputs(8152));
    outputs(1612) <= not((layer2_outputs(7334)) or (layer2_outputs(2741)));
    outputs(1613) <= not(layer2_outputs(12449)) or (layer2_outputs(442));
    outputs(1614) <= (layer2_outputs(1665)) and not (layer2_outputs(7590));
    outputs(1615) <= not((layer2_outputs(596)) xor (layer2_outputs(7777)));
    outputs(1616) <= layer2_outputs(3548);
    outputs(1617) <= layer2_outputs(8303);
    outputs(1618) <= (layer2_outputs(8568)) and (layer2_outputs(6839));
    outputs(1619) <= not((layer2_outputs(11358)) xor (layer2_outputs(10324)));
    outputs(1620) <= not(layer2_outputs(2373)) or (layer2_outputs(832));
    outputs(1621) <= (layer2_outputs(6621)) and not (layer2_outputs(10773));
    outputs(1622) <= not(layer2_outputs(3071));
    outputs(1623) <= not((layer2_outputs(11556)) xor (layer2_outputs(9810)));
    outputs(1624) <= not(layer2_outputs(12775));
    outputs(1625) <= (layer2_outputs(5616)) xor (layer2_outputs(5941));
    outputs(1626) <= (layer2_outputs(4323)) or (layer2_outputs(6473));
    outputs(1627) <= layer2_outputs(3606);
    outputs(1628) <= (layer2_outputs(5073)) and (layer2_outputs(9932));
    outputs(1629) <= layer2_outputs(8454);
    outputs(1630) <= (layer2_outputs(9165)) and not (layer2_outputs(2000));
    outputs(1631) <= (layer2_outputs(12007)) xor (layer2_outputs(6774));
    outputs(1632) <= layer2_outputs(8100);
    outputs(1633) <= not(layer2_outputs(7569));
    outputs(1634) <= (layer2_outputs(9609)) and not (layer2_outputs(2325));
    outputs(1635) <= (layer2_outputs(5482)) xor (layer2_outputs(11336));
    outputs(1636) <= not(layer2_outputs(6408)) or (layer2_outputs(2416));
    outputs(1637) <= layer2_outputs(10047);
    outputs(1638) <= not((layer2_outputs(12140)) xor (layer2_outputs(12520)));
    outputs(1639) <= (layer2_outputs(970)) and (layer2_outputs(7209));
    outputs(1640) <= not((layer2_outputs(10974)) xor (layer2_outputs(8504)));
    outputs(1641) <= (layer2_outputs(6580)) xor (layer2_outputs(1376));
    outputs(1642) <= (layer2_outputs(8848)) xor (layer2_outputs(2466));
    outputs(1643) <= not(layer2_outputs(10759));
    outputs(1644) <= layer2_outputs(10506);
    outputs(1645) <= not((layer2_outputs(8925)) and (layer2_outputs(10166)));
    outputs(1646) <= not((layer2_outputs(358)) xor (layer2_outputs(11269)));
    outputs(1647) <= (layer2_outputs(578)) and (layer2_outputs(7520));
    outputs(1648) <= layer2_outputs(8336);
    outputs(1649) <= not(layer2_outputs(4579));
    outputs(1650) <= (layer2_outputs(9658)) xor (layer2_outputs(9705));
    outputs(1651) <= layer2_outputs(7834);
    outputs(1652) <= not(layer2_outputs(1160));
    outputs(1653) <= not((layer2_outputs(6759)) xor (layer2_outputs(5774)));
    outputs(1654) <= not((layer2_outputs(8407)) xor (layer2_outputs(11865)));
    outputs(1655) <= not((layer2_outputs(12079)) xor (layer2_outputs(11360)));
    outputs(1656) <= not(layer2_outputs(12158));
    outputs(1657) <= not((layer2_outputs(2470)) or (layer2_outputs(1500)));
    outputs(1658) <= not(layer2_outputs(4759));
    outputs(1659) <= not(layer2_outputs(6890));
    outputs(1660) <= not(layer2_outputs(10829));
    outputs(1661) <= (layer2_outputs(9237)) and not (layer2_outputs(12006));
    outputs(1662) <= not((layer2_outputs(2004)) xor (layer2_outputs(2127)));
    outputs(1663) <= (layer2_outputs(3289)) and (layer2_outputs(12366));
    outputs(1664) <= not((layer2_outputs(7563)) or (layer2_outputs(6190)));
    outputs(1665) <= (layer2_outputs(2002)) or (layer2_outputs(4378));
    outputs(1666) <= not(layer2_outputs(7340));
    outputs(1667) <= not(layer2_outputs(1299));
    outputs(1668) <= not(layer2_outputs(3676));
    outputs(1669) <= not(layer2_outputs(12012));
    outputs(1670) <= (layer2_outputs(2541)) and (layer2_outputs(10112));
    outputs(1671) <= (layer2_outputs(10320)) xor (layer2_outputs(6103));
    outputs(1672) <= (layer2_outputs(11026)) and not (layer2_outputs(4265));
    outputs(1673) <= not(layer2_outputs(6648));
    outputs(1674) <= not((layer2_outputs(9164)) xor (layer2_outputs(1881)));
    outputs(1675) <= (layer2_outputs(12521)) and not (layer2_outputs(6739));
    outputs(1676) <= not(layer2_outputs(6480));
    outputs(1677) <= not(layer2_outputs(12572));
    outputs(1678) <= layer2_outputs(1883);
    outputs(1679) <= (layer2_outputs(9732)) xor (layer2_outputs(7640));
    outputs(1680) <= layer2_outputs(6086);
    outputs(1681) <= (layer2_outputs(2034)) and (layer2_outputs(7878));
    outputs(1682) <= not((layer2_outputs(10648)) xor (layer2_outputs(2877)));
    outputs(1683) <= (layer2_outputs(941)) and not (layer2_outputs(1538));
    outputs(1684) <= (layer2_outputs(3816)) or (layer2_outputs(11629));
    outputs(1685) <= not((layer2_outputs(8359)) and (layer2_outputs(8714)));
    outputs(1686) <= (layer2_outputs(5159)) and (layer2_outputs(8387));
    outputs(1687) <= not(layer2_outputs(8119));
    outputs(1688) <= not(layer2_outputs(1299));
    outputs(1689) <= (layer2_outputs(1998)) and not (layer2_outputs(9517));
    outputs(1690) <= layer2_outputs(9099);
    outputs(1691) <= not(layer2_outputs(3719));
    outputs(1692) <= not(layer2_outputs(470));
    outputs(1693) <= not(layer2_outputs(1461));
    outputs(1694) <= layer2_outputs(8600);
    outputs(1695) <= not((layer2_outputs(4017)) xor (layer2_outputs(2403)));
    outputs(1696) <= (layer2_outputs(11354)) xor (layer2_outputs(12550));
    outputs(1697) <= not((layer2_outputs(4051)) or (layer2_outputs(8945)));
    outputs(1698) <= not(layer2_outputs(7352));
    outputs(1699) <= not((layer2_outputs(5891)) or (layer2_outputs(4970)));
    outputs(1700) <= not(layer2_outputs(3668));
    outputs(1701) <= not((layer2_outputs(5087)) or (layer2_outputs(702)));
    outputs(1702) <= not(layer2_outputs(3834));
    outputs(1703) <= not((layer2_outputs(2712)) or (layer2_outputs(11331)));
    outputs(1704) <= not((layer2_outputs(9837)) xor (layer2_outputs(922)));
    outputs(1705) <= (layer2_outputs(10252)) and not (layer2_outputs(11856));
    outputs(1706) <= not((layer2_outputs(1447)) xor (layer2_outputs(4980)));
    outputs(1707) <= layer2_outputs(124);
    outputs(1708) <= layer2_outputs(11152);
    outputs(1709) <= (layer2_outputs(8327)) and not (layer2_outputs(1563));
    outputs(1710) <= (layer2_outputs(9714)) or (layer2_outputs(2696));
    outputs(1711) <= (layer2_outputs(3366)) and not (layer2_outputs(2409));
    outputs(1712) <= not(layer2_outputs(4885));
    outputs(1713) <= (layer2_outputs(1252)) and not (layer2_outputs(9180));
    outputs(1714) <= layer2_outputs(7388);
    outputs(1715) <= not(layer2_outputs(11914));
    outputs(1716) <= layer2_outputs(12351);
    outputs(1717) <= not(layer2_outputs(12453));
    outputs(1718) <= layer2_outputs(12668);
    outputs(1719) <= (layer2_outputs(11399)) and (layer2_outputs(7491));
    outputs(1720) <= not((layer2_outputs(507)) xor (layer2_outputs(6961)));
    outputs(1721) <= not((layer2_outputs(3333)) or (layer2_outputs(11033)));
    outputs(1722) <= (layer2_outputs(6978)) and (layer2_outputs(3942));
    outputs(1723) <= (layer2_outputs(8220)) xor (layer2_outputs(11205));
    outputs(1724) <= (layer2_outputs(10871)) xor (layer2_outputs(11757));
    outputs(1725) <= not(layer2_outputs(1943));
    outputs(1726) <= not(layer2_outputs(1512));
    outputs(1727) <= (layer2_outputs(1611)) and not (layer2_outputs(1274));
    outputs(1728) <= layer2_outputs(9046);
    outputs(1729) <= not(layer2_outputs(3438));
    outputs(1730) <= (layer2_outputs(2603)) xor (layer2_outputs(12177));
    outputs(1731) <= layer2_outputs(10008);
    outputs(1732) <= (layer2_outputs(8664)) and (layer2_outputs(4826));
    outputs(1733) <= layer2_outputs(4113);
    outputs(1734) <= not(layer2_outputs(8997));
    outputs(1735) <= (layer2_outputs(3016)) xor (layer2_outputs(868));
    outputs(1736) <= (layer2_outputs(5010)) xor (layer2_outputs(447));
    outputs(1737) <= layer2_outputs(3576);
    outputs(1738) <= not(layer2_outputs(8036));
    outputs(1739) <= not(layer2_outputs(12050));
    outputs(1740) <= layer2_outputs(2619);
    outputs(1741) <= layer2_outputs(10377);
    outputs(1742) <= not((layer2_outputs(1780)) and (layer2_outputs(8983)));
    outputs(1743) <= (layer2_outputs(11832)) and (layer2_outputs(2371));
    outputs(1744) <= not((layer2_outputs(7621)) xor (layer2_outputs(7369)));
    outputs(1745) <= (layer2_outputs(7691)) xor (layer2_outputs(10968));
    outputs(1746) <= not((layer2_outputs(1537)) xor (layer2_outputs(11083)));
    outputs(1747) <= not((layer2_outputs(7177)) or (layer2_outputs(9074)));
    outputs(1748) <= layer2_outputs(11472);
    outputs(1749) <= not((layer2_outputs(11873)) xor (layer2_outputs(497)));
    outputs(1750) <= (layer2_outputs(4597)) xor (layer2_outputs(8474));
    outputs(1751) <= '1';
    outputs(1752) <= not((layer2_outputs(1788)) xor (layer2_outputs(5990)));
    outputs(1753) <= not(layer2_outputs(5065));
    outputs(1754) <= layer2_outputs(4072);
    outputs(1755) <= not(layer2_outputs(11253));
    outputs(1756) <= not((layer2_outputs(3108)) or (layer2_outputs(5689)));
    outputs(1757) <= (layer2_outputs(9222)) and (layer2_outputs(6082));
    outputs(1758) <= not((layer2_outputs(8899)) xor (layer2_outputs(1828)));
    outputs(1759) <= not(layer2_outputs(7818));
    outputs(1760) <= layer2_outputs(5242);
    outputs(1761) <= not((layer2_outputs(1058)) xor (layer2_outputs(2548)));
    outputs(1762) <= not(layer2_outputs(6141));
    outputs(1763) <= layer2_outputs(7161);
    outputs(1764) <= not((layer2_outputs(4740)) or (layer2_outputs(6654)));
    outputs(1765) <= not(layer2_outputs(352));
    outputs(1766) <= (layer2_outputs(10149)) and (layer2_outputs(8303));
    outputs(1767) <= not(layer2_outputs(10088));
    outputs(1768) <= (layer2_outputs(6011)) and (layer2_outputs(9556));
    outputs(1769) <= not(layer2_outputs(10901));
    outputs(1770) <= (layer2_outputs(10101)) xor (layer2_outputs(5094));
    outputs(1771) <= not((layer2_outputs(7066)) xor (layer2_outputs(5193)));
    outputs(1772) <= (layer2_outputs(4975)) and (layer2_outputs(6206));
    outputs(1773) <= (layer2_outputs(4403)) and (layer2_outputs(7219));
    outputs(1774) <= not((layer2_outputs(8782)) xor (layer2_outputs(6628)));
    outputs(1775) <= not((layer2_outputs(7465)) xor (layer2_outputs(9485)));
    outputs(1776) <= not(layer2_outputs(11930));
    outputs(1777) <= layer2_outputs(9239);
    outputs(1778) <= layer2_outputs(3327);
    outputs(1779) <= not((layer2_outputs(10398)) xor (layer2_outputs(6310)));
    outputs(1780) <= (layer2_outputs(4700)) xor (layer2_outputs(9455));
    outputs(1781) <= (layer2_outputs(1762)) xor (layer2_outputs(1794));
    outputs(1782) <= (layer2_outputs(2353)) and not (layer2_outputs(11563));
    outputs(1783) <= (layer2_outputs(6446)) xor (layer2_outputs(2407));
    outputs(1784) <= not(layer2_outputs(11928));
    outputs(1785) <= not((layer2_outputs(157)) xor (layer2_outputs(11887)));
    outputs(1786) <= not((layer2_outputs(6259)) or (layer2_outputs(9058)));
    outputs(1787) <= not(layer2_outputs(12162));
    outputs(1788) <= not((layer2_outputs(3356)) or (layer2_outputs(5830)));
    outputs(1789) <= not(layer2_outputs(5717));
    outputs(1790) <= (layer2_outputs(2613)) xor (layer2_outputs(1433));
    outputs(1791) <= (layer2_outputs(3771)) and not (layer2_outputs(1697));
    outputs(1792) <= not((layer2_outputs(11099)) or (layer2_outputs(4911)));
    outputs(1793) <= layer2_outputs(2284);
    outputs(1794) <= not((layer2_outputs(272)) or (layer2_outputs(11093)));
    outputs(1795) <= (layer2_outputs(3825)) and not (layer2_outputs(12397));
    outputs(1796) <= (layer2_outputs(7485)) and (layer2_outputs(12741));
    outputs(1797) <= layer2_outputs(3177);
    outputs(1798) <= (layer2_outputs(4774)) xor (layer2_outputs(885));
    outputs(1799) <= (layer2_outputs(8095)) xor (layer2_outputs(6642));
    outputs(1800) <= (layer2_outputs(1094)) xor (layer2_outputs(6108));
    outputs(1801) <= not((layer2_outputs(5155)) or (layer2_outputs(105)));
    outputs(1802) <= (layer2_outputs(11938)) xor (layer2_outputs(7225));
    outputs(1803) <= not(layer2_outputs(5209));
    outputs(1804) <= not(layer2_outputs(2172));
    outputs(1805) <= layer2_outputs(6421);
    outputs(1806) <= not((layer2_outputs(12315)) xor (layer2_outputs(9187)));
    outputs(1807) <= not((layer2_outputs(10942)) or (layer2_outputs(8140)));
    outputs(1808) <= layer2_outputs(12147);
    outputs(1809) <= (layer2_outputs(742)) and not (layer2_outputs(1866));
    outputs(1810) <= not(layer2_outputs(1472));
    outputs(1811) <= not(layer2_outputs(8252));
    outputs(1812) <= not(layer2_outputs(6150));
    outputs(1813) <= (layer2_outputs(5981)) xor (layer2_outputs(7421));
    outputs(1814) <= layer2_outputs(6621);
    outputs(1815) <= not(layer2_outputs(6656));
    outputs(1816) <= (layer2_outputs(1123)) xor (layer2_outputs(9512));
    outputs(1817) <= (layer2_outputs(9389)) and not (layer2_outputs(11689));
    outputs(1818) <= not(layer2_outputs(1046));
    outputs(1819) <= (layer2_outputs(875)) xor (layer2_outputs(12621));
    outputs(1820) <= not(layer2_outputs(7017)) or (layer2_outputs(3366));
    outputs(1821) <= (layer2_outputs(5048)) xor (layer2_outputs(11932));
    outputs(1822) <= not((layer2_outputs(9188)) xor (layer2_outputs(11420)));
    outputs(1823) <= not((layer2_outputs(7781)) or (layer2_outputs(3547)));
    outputs(1824) <= (layer2_outputs(653)) and not (layer2_outputs(1919));
    outputs(1825) <= not((layer2_outputs(2443)) or (layer2_outputs(162)));
    outputs(1826) <= not((layer2_outputs(8417)) or (layer2_outputs(2054)));
    outputs(1827) <= not((layer2_outputs(10704)) or (layer2_outputs(9140)));
    outputs(1828) <= not(layer2_outputs(2692));
    outputs(1829) <= (layer2_outputs(10744)) xor (layer2_outputs(5797));
    outputs(1830) <= not((layer2_outputs(1400)) xor (layer2_outputs(6691)));
    outputs(1831) <= not((layer2_outputs(8550)) xor (layer2_outputs(7957)));
    outputs(1832) <= layer2_outputs(5957);
    outputs(1833) <= not((layer2_outputs(1347)) or (layer2_outputs(11060)));
    outputs(1834) <= layer2_outputs(3539);
    outputs(1835) <= not(layer2_outputs(3589));
    outputs(1836) <= not(layer2_outputs(5369));
    outputs(1837) <= not((layer2_outputs(7403)) xor (layer2_outputs(4214)));
    outputs(1838) <= layer2_outputs(8092);
    outputs(1839) <= not(layer2_outputs(1948));
    outputs(1840) <= not((layer2_outputs(1401)) or (layer2_outputs(11886)));
    outputs(1841) <= layer2_outputs(974);
    outputs(1842) <= layer2_outputs(2693);
    outputs(1843) <= not(layer2_outputs(3574));
    outputs(1844) <= layer2_outputs(12573);
    outputs(1845) <= layer2_outputs(7149);
    outputs(1846) <= not(layer2_outputs(516));
    outputs(1847) <= not((layer2_outputs(1894)) xor (layer2_outputs(758)));
    outputs(1848) <= not((layer2_outputs(3231)) xor (layer2_outputs(5980)));
    outputs(1849) <= not(layer2_outputs(10476));
    outputs(1850) <= layer2_outputs(5564);
    outputs(1851) <= (layer2_outputs(7804)) and (layer2_outputs(11187));
    outputs(1852) <= layer2_outputs(9646);
    outputs(1853) <= layer2_outputs(7614);
    outputs(1854) <= not(layer2_outputs(1552));
    outputs(1855) <= (layer2_outputs(8052)) and (layer2_outputs(8588));
    outputs(1856) <= layer2_outputs(9014);
    outputs(1857) <= layer2_outputs(10791);
    outputs(1858) <= (layer2_outputs(9926)) xor (layer2_outputs(6428));
    outputs(1859) <= not((layer2_outputs(5261)) xor (layer2_outputs(10762)));
    outputs(1860) <= layer2_outputs(12502);
    outputs(1861) <= (layer2_outputs(11131)) and (layer2_outputs(10681));
    outputs(1862) <= not((layer2_outputs(4450)) xor (layer2_outputs(4346)));
    outputs(1863) <= (layer2_outputs(10187)) and (layer2_outputs(1266));
    outputs(1864) <= (layer2_outputs(9161)) and not (layer2_outputs(11822));
    outputs(1865) <= layer2_outputs(9398);
    outputs(1866) <= (layer2_outputs(3481)) xor (layer2_outputs(7774));
    outputs(1867) <= not((layer2_outputs(1590)) or (layer2_outputs(10014)));
    outputs(1868) <= not(layer2_outputs(420));
    outputs(1869) <= not((layer2_outputs(1121)) or (layer2_outputs(1848)));
    outputs(1870) <= layer2_outputs(6125);
    outputs(1871) <= not((layer2_outputs(1919)) xor (layer2_outputs(10749)));
    outputs(1872) <= not(layer2_outputs(1010));
    outputs(1873) <= (layer2_outputs(6679)) xor (layer2_outputs(325));
    outputs(1874) <= (layer2_outputs(7573)) xor (layer2_outputs(5782));
    outputs(1875) <= not((layer2_outputs(4246)) xor (layer2_outputs(12072)));
    outputs(1876) <= (layer2_outputs(7125)) and not (layer2_outputs(9083));
    outputs(1877) <= not((layer2_outputs(11507)) xor (layer2_outputs(3065)));
    outputs(1878) <= not(layer2_outputs(691));
    outputs(1879) <= layer2_outputs(2828);
    outputs(1880) <= not(layer2_outputs(1310));
    outputs(1881) <= (layer2_outputs(1487)) and not (layer2_outputs(7454));
    outputs(1882) <= not(layer2_outputs(7337));
    outputs(1883) <= (layer2_outputs(7262)) and (layer2_outputs(12201));
    outputs(1884) <= (layer2_outputs(2663)) xor (layer2_outputs(766));
    outputs(1885) <= not((layer2_outputs(11695)) xor (layer2_outputs(8524)));
    outputs(1886) <= not(layer2_outputs(7440)) or (layer2_outputs(1850));
    outputs(1887) <= not(layer2_outputs(3890));
    outputs(1888) <= not((layer2_outputs(9686)) xor (layer2_outputs(6495)));
    outputs(1889) <= (layer2_outputs(12084)) xor (layer2_outputs(11335));
    outputs(1890) <= not((layer2_outputs(3705)) xor (layer2_outputs(4537)));
    outputs(1891) <= (layer2_outputs(5221)) and not (layer2_outputs(3189));
    outputs(1892) <= layer2_outputs(12587);
    outputs(1893) <= not(layer2_outputs(10763));
    outputs(1894) <= (layer2_outputs(431)) and (layer2_outputs(5748));
    outputs(1895) <= (layer2_outputs(1952)) and not (layer2_outputs(10084));
    outputs(1896) <= (layer2_outputs(9643)) or (layer2_outputs(4211));
    outputs(1897) <= not(layer2_outputs(6827)) or (layer2_outputs(6493));
    outputs(1898) <= not((layer2_outputs(7182)) xor (layer2_outputs(562)));
    outputs(1899) <= not(layer2_outputs(266));
    outputs(1900) <= (layer2_outputs(12666)) xor (layer2_outputs(6037));
    outputs(1901) <= not((layer2_outputs(10490)) or (layer2_outputs(7657)));
    outputs(1902) <= (layer2_outputs(4379)) and not (layer2_outputs(8751));
    outputs(1903) <= (layer2_outputs(2072)) xor (layer2_outputs(1255));
    outputs(1904) <= not(layer2_outputs(9485));
    outputs(1905) <= (layer2_outputs(10936)) xor (layer2_outputs(2522));
    outputs(1906) <= not(layer2_outputs(4006));
    outputs(1907) <= not((layer2_outputs(2760)) or (layer2_outputs(4643)));
    outputs(1908) <= not((layer2_outputs(11561)) xor (layer2_outputs(2322)));
    outputs(1909) <= not((layer2_outputs(6001)) or (layer2_outputs(684)));
    outputs(1910) <= not((layer2_outputs(11625)) or (layer2_outputs(2834)));
    outputs(1911) <= (layer2_outputs(11982)) and not (layer2_outputs(10080));
    outputs(1912) <= layer2_outputs(12567);
    outputs(1913) <= not((layer2_outputs(1834)) xor (layer2_outputs(3524)));
    outputs(1914) <= (layer2_outputs(10731)) xor (layer2_outputs(5700));
    outputs(1915) <= (layer2_outputs(2710)) and not (layer2_outputs(4673));
    outputs(1916) <= not(layer2_outputs(4880));
    outputs(1917) <= not(layer2_outputs(10737));
    outputs(1918) <= not(layer2_outputs(983));
    outputs(1919) <= not(layer2_outputs(12122));
    outputs(1920) <= layer2_outputs(7827);
    outputs(1921) <= not(layer2_outputs(10663));
    outputs(1922) <= layer2_outputs(7574);
    outputs(1923) <= (layer2_outputs(9865)) xor (layer2_outputs(10446));
    outputs(1924) <= not((layer2_outputs(4172)) or (layer2_outputs(9859)));
    outputs(1925) <= not((layer2_outputs(10441)) xor (layer2_outputs(8594)));
    outputs(1926) <= layer2_outputs(5256);
    outputs(1927) <= not((layer2_outputs(11477)) xor (layer2_outputs(12224)));
    outputs(1928) <= not(layer2_outputs(2961));
    outputs(1929) <= not(layer2_outputs(2087));
    outputs(1930) <= (layer2_outputs(12764)) and not (layer2_outputs(7099));
    outputs(1931) <= (layer2_outputs(4341)) and not (layer2_outputs(9208));
    outputs(1932) <= not((layer2_outputs(2685)) or (layer2_outputs(10087)));
    outputs(1933) <= (layer2_outputs(12750)) and not (layer2_outputs(9837));
    outputs(1934) <= not((layer2_outputs(8850)) xor (layer2_outputs(11938)));
    outputs(1935) <= (layer2_outputs(7919)) xor (layer2_outputs(2840));
    outputs(1936) <= layer2_outputs(4816);
    outputs(1937) <= not((layer2_outputs(9292)) xor (layer2_outputs(7178)));
    outputs(1938) <= not((layer2_outputs(1108)) xor (layer2_outputs(8159)));
    outputs(1939) <= layer2_outputs(10651);
    outputs(1940) <= layer2_outputs(12238);
    outputs(1941) <= not(layer2_outputs(9476));
    outputs(1942) <= (layer2_outputs(2596)) xor (layer2_outputs(242));
    outputs(1943) <= not((layer2_outputs(10231)) xor (layer2_outputs(8946)));
    outputs(1944) <= (layer2_outputs(8609)) xor (layer2_outputs(9152));
    outputs(1945) <= (layer2_outputs(11803)) and (layer2_outputs(8855));
    outputs(1946) <= layer2_outputs(3367);
    outputs(1947) <= (layer2_outputs(3702)) xor (layer2_outputs(3063));
    outputs(1948) <= not((layer2_outputs(3368)) xor (layer2_outputs(12434)));
    outputs(1949) <= layer2_outputs(995);
    outputs(1950) <= not(layer2_outputs(7693));
    outputs(1951) <= not((layer2_outputs(12009)) xor (layer2_outputs(7103)));
    outputs(1952) <= (layer2_outputs(6355)) xor (layer2_outputs(11061));
    outputs(1953) <= layer2_outputs(1526);
    outputs(1954) <= not((layer2_outputs(5974)) or (layer2_outputs(4759)));
    outputs(1955) <= (layer2_outputs(7432)) and not (layer2_outputs(1833));
    outputs(1956) <= not(layer2_outputs(7890));
    outputs(1957) <= (layer2_outputs(7441)) and not (layer2_outputs(2461));
    outputs(1958) <= not((layer2_outputs(1999)) xor (layer2_outputs(8310)));
    outputs(1959) <= layer2_outputs(6970);
    outputs(1960) <= not((layer2_outputs(6191)) or (layer2_outputs(7942)));
    outputs(1961) <= not(layer2_outputs(3236));
    outputs(1962) <= not(layer2_outputs(297));
    outputs(1963) <= layer2_outputs(7525);
    outputs(1964) <= not(layer2_outputs(7708));
    outputs(1965) <= not((layer2_outputs(11801)) and (layer2_outputs(5390)));
    outputs(1966) <= not((layer2_outputs(77)) xor (layer2_outputs(6836)));
    outputs(1967) <= not(layer2_outputs(8821));
    outputs(1968) <= not((layer2_outputs(8597)) xor (layer2_outputs(5291)));
    outputs(1969) <= layer2_outputs(9588);
    outputs(1970) <= (layer2_outputs(9866)) xor (layer2_outputs(754));
    outputs(1971) <= not(layer2_outputs(9796));
    outputs(1972) <= not((layer2_outputs(1349)) xor (layer2_outputs(3713)));
    outputs(1973) <= not(layer2_outputs(4252));
    outputs(1974) <= not((layer2_outputs(8356)) or (layer2_outputs(714)));
    outputs(1975) <= not((layer2_outputs(5456)) and (layer2_outputs(5099)));
    outputs(1976) <= not((layer2_outputs(10368)) xor (layer2_outputs(6748)));
    outputs(1977) <= not(layer2_outputs(9935));
    outputs(1978) <= layer2_outputs(4782);
    outputs(1979) <= (layer2_outputs(2438)) and (layer2_outputs(9890));
    outputs(1980) <= layer2_outputs(8804);
    outputs(1981) <= (layer2_outputs(4982)) and not (layer2_outputs(2581));
    outputs(1982) <= not((layer2_outputs(5515)) xor (layer2_outputs(1525)));
    outputs(1983) <= not((layer2_outputs(436)) xor (layer2_outputs(4708)));
    outputs(1984) <= not(layer2_outputs(4526));
    outputs(1985) <= (layer2_outputs(4770)) and (layer2_outputs(4230));
    outputs(1986) <= not((layer2_outputs(4825)) or (layer2_outputs(2130)));
    outputs(1987) <= (layer2_outputs(3403)) xor (layer2_outputs(4939));
    outputs(1988) <= not(layer2_outputs(1448));
    outputs(1989) <= not(layer2_outputs(3384)) or (layer2_outputs(7775));
    outputs(1990) <= not((layer2_outputs(9405)) xor (layer2_outputs(5669)));
    outputs(1991) <= (layer2_outputs(10865)) xor (layer2_outputs(9474));
    outputs(1992) <= not(layer2_outputs(8213));
    outputs(1993) <= not((layer2_outputs(12207)) xor (layer2_outputs(4987)));
    outputs(1994) <= not((layer2_outputs(2754)) xor (layer2_outputs(121)));
    outputs(1995) <= layer2_outputs(8388);
    outputs(1996) <= (layer2_outputs(10049)) and not (layer2_outputs(861));
    outputs(1997) <= (layer2_outputs(11797)) xor (layer2_outputs(2041));
    outputs(1998) <= not(layer2_outputs(11048));
    outputs(1999) <= layer2_outputs(8921);
    outputs(2000) <= not(layer2_outputs(7735));
    outputs(2001) <= not((layer2_outputs(5676)) or (layer2_outputs(10428)));
    outputs(2002) <= not((layer2_outputs(1697)) or (layer2_outputs(7001)));
    outputs(2003) <= layer2_outputs(4951);
    outputs(2004) <= not(layer2_outputs(8195));
    outputs(2005) <= not(layer2_outputs(2157));
    outputs(2006) <= layer2_outputs(1092);
    outputs(2007) <= (layer2_outputs(8355)) and not (layer2_outputs(3257));
    outputs(2008) <= not((layer2_outputs(9107)) or (layer2_outputs(6724)));
    outputs(2009) <= not(layer2_outputs(1063));
    outputs(2010) <= (layer2_outputs(5326)) and not (layer2_outputs(4407));
    outputs(2011) <= not(layer2_outputs(1604));
    outputs(2012) <= not((layer2_outputs(8145)) or (layer2_outputs(7992)));
    outputs(2013) <= not(layer2_outputs(4886));
    outputs(2014) <= layer2_outputs(6068);
    outputs(2015) <= not(layer2_outputs(3150));
    outputs(2016) <= (layer2_outputs(5608)) and not (layer2_outputs(1464));
    outputs(2017) <= (layer2_outputs(6861)) and not (layer2_outputs(4831));
    outputs(2018) <= not((layer2_outputs(83)) or (layer2_outputs(11465)));
    outputs(2019) <= not(layer2_outputs(11456));
    outputs(2020) <= layer2_outputs(9870);
    outputs(2021) <= not(layer2_outputs(11885)) or (layer2_outputs(9953));
    outputs(2022) <= layer2_outputs(1435);
    outputs(2023) <= not((layer2_outputs(1276)) or (layer2_outputs(528)));
    outputs(2024) <= (layer2_outputs(6271)) xor (layer2_outputs(12231));
    outputs(2025) <= not(layer2_outputs(5076));
    outputs(2026) <= not((layer2_outputs(10206)) or (layer2_outputs(7439)));
    outputs(2027) <= layer2_outputs(4060);
    outputs(2028) <= (layer2_outputs(7982)) xor (layer2_outputs(7521));
    outputs(2029) <= layer2_outputs(4242);
    outputs(2030) <= not((layer2_outputs(1394)) xor (layer2_outputs(7602)));
    outputs(2031) <= (layer2_outputs(7112)) and not (layer2_outputs(4468));
    outputs(2032) <= not(layer2_outputs(12570));
    outputs(2033) <= (layer2_outputs(8149)) xor (layer2_outputs(664));
    outputs(2034) <= layer2_outputs(4950);
    outputs(2035) <= layer2_outputs(3554);
    outputs(2036) <= layer2_outputs(5440);
    outputs(2037) <= not((layer2_outputs(3915)) or (layer2_outputs(6654)));
    outputs(2038) <= not((layer2_outputs(11659)) xor (layer2_outputs(6768)));
    outputs(2039) <= not((layer2_outputs(284)) or (layer2_outputs(12625)));
    outputs(2040) <= layer2_outputs(9785);
    outputs(2041) <= not(layer2_outputs(6448));
    outputs(2042) <= not(layer2_outputs(10156));
    outputs(2043) <= not((layer2_outputs(5144)) or (layer2_outputs(2942)));
    outputs(2044) <= (layer2_outputs(4704)) and not (layer2_outputs(10050));
    outputs(2045) <= (layer2_outputs(10585)) xor (layer2_outputs(59));
    outputs(2046) <= not((layer2_outputs(215)) xor (layer2_outputs(9840)));
    outputs(2047) <= not(layer2_outputs(4866));
    outputs(2048) <= (layer2_outputs(9204)) and not (layer2_outputs(11958));
    outputs(2049) <= layer2_outputs(6852);
    outputs(2050) <= (layer2_outputs(5952)) xor (layer2_outputs(12733));
    outputs(2051) <= (layer2_outputs(9853)) xor (layer2_outputs(11357));
    outputs(2052) <= layer2_outputs(1673);
    outputs(2053) <= not((layer2_outputs(5026)) or (layer2_outputs(7655)));
    outputs(2054) <= layer2_outputs(11788);
    outputs(2055) <= not(layer2_outputs(8275));
    outputs(2056) <= not(layer2_outputs(11366));
    outputs(2057) <= (layer2_outputs(3632)) and not (layer2_outputs(4220));
    outputs(2058) <= not(layer2_outputs(6554));
    outputs(2059) <= layer2_outputs(749);
    outputs(2060) <= not((layer2_outputs(1176)) xor (layer2_outputs(10976)));
    outputs(2061) <= not(layer2_outputs(3741));
    outputs(2062) <= (layer2_outputs(5409)) and (layer2_outputs(3985));
    outputs(2063) <= (layer2_outputs(3545)) and not (layer2_outputs(11291));
    outputs(2064) <= (layer2_outputs(2446)) and (layer2_outputs(751));
    outputs(2065) <= layer2_outputs(5605);
    outputs(2066) <= not(layer2_outputs(5274));
    outputs(2067) <= (layer2_outputs(11835)) xor (layer2_outputs(2481));
    outputs(2068) <= not((layer2_outputs(799)) and (layer2_outputs(3729)));
    outputs(2069) <= not((layer2_outputs(12121)) or (layer2_outputs(6522)));
    outputs(2070) <= not((layer2_outputs(2326)) or (layer2_outputs(6609)));
    outputs(2071) <= not((layer2_outputs(10546)) xor (layer2_outputs(6995)));
    outputs(2072) <= not((layer2_outputs(5910)) xor (layer2_outputs(5863)));
    outputs(2073) <= layer2_outputs(9615);
    outputs(2074) <= layer2_outputs(10440);
    outputs(2075) <= (layer2_outputs(4609)) and (layer2_outputs(4469));
    outputs(2076) <= (layer2_outputs(6099)) and not (layer2_outputs(385));
    outputs(2077) <= (layer2_outputs(965)) xor (layer2_outputs(9399));
    outputs(2078) <= layer2_outputs(8270);
    outputs(2079) <= (layer2_outputs(6413)) and (layer2_outputs(11728));
    outputs(2080) <= not(layer2_outputs(8413));
    outputs(2081) <= not((layer2_outputs(6562)) or (layer2_outputs(11775)));
    outputs(2082) <= layer2_outputs(6129);
    outputs(2083) <= layer2_outputs(1815);
    outputs(2084) <= (layer2_outputs(4560)) xor (layer2_outputs(8507));
    outputs(2085) <= layer2_outputs(12065);
    outputs(2086) <= (layer2_outputs(4084)) and not (layer2_outputs(580));
    outputs(2087) <= not(layer2_outputs(5015));
    outputs(2088) <= (layer2_outputs(4318)) and not (layer2_outputs(8569));
    outputs(2089) <= layer2_outputs(6091);
    outputs(2090) <= not(layer2_outputs(6212));
    outputs(2091) <= (layer2_outputs(7428)) xor (layer2_outputs(2893));
    outputs(2092) <= (layer2_outputs(4961)) and (layer2_outputs(8786));
    outputs(2093) <= (layer2_outputs(8400)) and not (layer2_outputs(12163));
    outputs(2094) <= not((layer2_outputs(6767)) xor (layer2_outputs(11651)));
    outputs(2095) <= not(layer2_outputs(6316));
    outputs(2096) <= layer2_outputs(180);
    outputs(2097) <= not((layer2_outputs(4486)) xor (layer2_outputs(4442)));
    outputs(2098) <= not((layer2_outputs(10123)) xor (layer2_outputs(1718)));
    outputs(2099) <= not((layer2_outputs(4191)) xor (layer2_outputs(8527)));
    outputs(2100) <= (layer2_outputs(4045)) xor (layer2_outputs(10694));
    outputs(2101) <= layer2_outputs(4384);
    outputs(2102) <= layer2_outputs(9772);
    outputs(2103) <= not((layer2_outputs(11973)) or (layer2_outputs(5785)));
    outputs(2104) <= not(layer2_outputs(11134));
    outputs(2105) <= not(layer2_outputs(7582));
    outputs(2106) <= not((layer2_outputs(2043)) xor (layer2_outputs(3592)));
    outputs(2107) <= not((layer2_outputs(11909)) xor (layer2_outputs(1643)));
    outputs(2108) <= not((layer2_outputs(11751)) xor (layer2_outputs(7656)));
    outputs(2109) <= (layer2_outputs(4960)) and (layer2_outputs(8627));
    outputs(2110) <= (layer2_outputs(4097)) and not (layer2_outputs(6529));
    outputs(2111) <= (layer2_outputs(4721)) or (layer2_outputs(5618));
    outputs(2112) <= layer2_outputs(3259);
    outputs(2113) <= (layer2_outputs(8249)) and not (layer2_outputs(1001));
    outputs(2114) <= (layer2_outputs(6675)) and not (layer2_outputs(5982));
    outputs(2115) <= (layer2_outputs(12427)) or (layer2_outputs(9249));
    outputs(2116) <= not(layer2_outputs(6714));
    outputs(2117) <= not(layer2_outputs(1664));
    outputs(2118) <= layer2_outputs(9362);
    outputs(2119) <= not((layer2_outputs(10806)) xor (layer2_outputs(9083)));
    outputs(2120) <= (layer2_outputs(3208)) and (layer2_outputs(9398));
    outputs(2121) <= not((layer2_outputs(4937)) or (layer2_outputs(11791)));
    outputs(2122) <= layer2_outputs(8844);
    outputs(2123) <= layer2_outputs(1153);
    outputs(2124) <= (layer2_outputs(8625)) and not (layer2_outputs(4236));
    outputs(2125) <= layer2_outputs(11561);
    outputs(2126) <= not(layer2_outputs(4339));
    outputs(2127) <= not(layer2_outputs(7897));
    outputs(2128) <= not((layer2_outputs(12769)) xor (layer2_outputs(2275)));
    outputs(2129) <= not((layer2_outputs(8143)) xor (layer2_outputs(423)));
    outputs(2130) <= (layer2_outputs(2366)) xor (layer2_outputs(820));
    outputs(2131) <= not((layer2_outputs(5854)) xor (layer2_outputs(11034)));
    outputs(2132) <= not((layer2_outputs(5148)) or (layer2_outputs(5812)));
    outputs(2133) <= not((layer2_outputs(8621)) xor (layer2_outputs(5393)));
    outputs(2134) <= (layer2_outputs(9052)) xor (layer2_outputs(6322));
    outputs(2135) <= not(layer2_outputs(9936));
    outputs(2136) <= (layer2_outputs(9148)) and not (layer2_outputs(11066));
    outputs(2137) <= (layer2_outputs(7139)) and not (layer2_outputs(1415));
    outputs(2138) <= not((layer2_outputs(6356)) xor (layer2_outputs(10482)));
    outputs(2139) <= not(layer2_outputs(10704));
    outputs(2140) <= not(layer2_outputs(4301));
    outputs(2141) <= not((layer2_outputs(1287)) xor (layer2_outputs(5619)));
    outputs(2142) <= (layer2_outputs(4844)) and not (layer2_outputs(747));
    outputs(2143) <= (layer2_outputs(8783)) and (layer2_outputs(4427));
    outputs(2144) <= not((layer2_outputs(4048)) xor (layer2_outputs(4600)));
    outputs(2145) <= not(layer2_outputs(10226));
    outputs(2146) <= not((layer2_outputs(6197)) xor (layer2_outputs(583)));
    outputs(2147) <= (layer2_outputs(9464)) xor (layer2_outputs(4092));
    outputs(2148) <= (layer2_outputs(10365)) or (layer2_outputs(8189));
    outputs(2149) <= layer2_outputs(3816);
    outputs(2150) <= (layer2_outputs(5998)) and (layer2_outputs(6289));
    outputs(2151) <= (layer2_outputs(9809)) and not (layer2_outputs(4518));
    outputs(2152) <= layer2_outputs(6559);
    outputs(2153) <= not(layer2_outputs(8956)) or (layer2_outputs(3383));
    outputs(2154) <= not(layer2_outputs(3578));
    outputs(2155) <= not(layer2_outputs(536));
    outputs(2156) <= not((layer2_outputs(7156)) or (layer2_outputs(5167)));
    outputs(2157) <= not((layer2_outputs(898)) or (layer2_outputs(3605)));
    outputs(2158) <= (layer2_outputs(1728)) xor (layer2_outputs(10003));
    outputs(2159) <= not(layer2_outputs(6844));
    outputs(2160) <= not((layer2_outputs(5842)) xor (layer2_outputs(12026)));
    outputs(2161) <= not((layer2_outputs(2848)) xor (layer2_outputs(2187)));
    outputs(2162) <= layer2_outputs(4984);
    outputs(2163) <= (layer2_outputs(1781)) and not (layer2_outputs(10298));
    outputs(2164) <= (layer2_outputs(7500)) xor (layer2_outputs(12374));
    outputs(2165) <= (layer2_outputs(4773)) and not (layer2_outputs(2622));
    outputs(2166) <= not(layer2_outputs(11676));
    outputs(2167) <= not((layer2_outputs(1842)) xor (layer2_outputs(1441)));
    outputs(2168) <= (layer2_outputs(11193)) or (layer2_outputs(5468));
    outputs(2169) <= (layer2_outputs(5521)) and not (layer2_outputs(11764));
    outputs(2170) <= not(layer2_outputs(9630));
    outputs(2171) <= (layer2_outputs(10958)) xor (layer2_outputs(6986));
    outputs(2172) <= not((layer2_outputs(5165)) xor (layer2_outputs(7758)));
    outputs(2173) <= layer2_outputs(2586);
    outputs(2174) <= not(layer2_outputs(8212));
    outputs(2175) <= (layer2_outputs(5993)) xor (layer2_outputs(3020));
    outputs(2176) <= not((layer2_outputs(10719)) or (layer2_outputs(12153)));
    outputs(2177) <= (layer2_outputs(2021)) and not (layer2_outputs(8329));
    outputs(2178) <= (layer2_outputs(3632)) and (layer2_outputs(177));
    outputs(2179) <= (layer2_outputs(12661)) and not (layer2_outputs(12676));
    outputs(2180) <= layer2_outputs(1772);
    outputs(2181) <= layer2_outputs(4792);
    outputs(2182) <= (layer2_outputs(305)) and not (layer2_outputs(6043));
    outputs(2183) <= (layer2_outputs(1826)) and not (layer2_outputs(6355));
    outputs(2184) <= not(layer2_outputs(2319));
    outputs(2185) <= not((layer2_outputs(10475)) xor (layer2_outputs(5986)));
    outputs(2186) <= (layer2_outputs(2162)) xor (layer2_outputs(9242));
    outputs(2187) <= layer2_outputs(3514);
    outputs(2188) <= not(layer2_outputs(1702));
    outputs(2189) <= not(layer2_outputs(9104));
    outputs(2190) <= (layer2_outputs(8670)) xor (layer2_outputs(12689));
    outputs(2191) <= (layer2_outputs(5425)) xor (layer2_outputs(921));
    outputs(2192) <= not(layer2_outputs(2391));
    outputs(2193) <= layer2_outputs(3067);
    outputs(2194) <= layer2_outputs(6556);
    outputs(2195) <= not((layer2_outputs(4601)) xor (layer2_outputs(5097)));
    outputs(2196) <= not(layer2_outputs(1872));
    outputs(2197) <= (layer2_outputs(3029)) xor (layer2_outputs(3443));
    outputs(2198) <= (layer2_outputs(10369)) xor (layer2_outputs(3701));
    outputs(2199) <= (layer2_outputs(8294)) and (layer2_outputs(2555));
    outputs(2200) <= (layer2_outputs(10279)) and not (layer2_outputs(3135));
    outputs(2201) <= not(layer2_outputs(6546));
    outputs(2202) <= not(layer2_outputs(12754));
    outputs(2203) <= not(layer2_outputs(4578));
    outputs(2204) <= (layer2_outputs(5852)) and not (layer2_outputs(1865));
    outputs(2205) <= layer2_outputs(2318);
    outputs(2206) <= not(layer2_outputs(2189));
    outputs(2207) <= (layer2_outputs(12790)) and not (layer2_outputs(3560));
    outputs(2208) <= not((layer2_outputs(10034)) xor (layer2_outputs(9996)));
    outputs(2209) <= (layer2_outputs(10621)) xor (layer2_outputs(5775));
    outputs(2210) <= layer2_outputs(11736);
    outputs(2211) <= not(layer2_outputs(1990)) or (layer2_outputs(10019));
    outputs(2212) <= layer2_outputs(8539);
    outputs(2213) <= not(layer2_outputs(398));
    outputs(2214) <= (layer2_outputs(10049)) and not (layer2_outputs(12137));
    outputs(2215) <= not((layer2_outputs(7018)) xor (layer2_outputs(5122)));
    outputs(2216) <= (layer2_outputs(4041)) and (layer2_outputs(6560));
    outputs(2217) <= (layer2_outputs(11574)) and not (layer2_outputs(96));
    outputs(2218) <= (layer2_outputs(233)) xor (layer2_outputs(11077));
    outputs(2219) <= not(layer2_outputs(8665));
    outputs(2220) <= not(layer2_outputs(12175));
    outputs(2221) <= layer2_outputs(12471);
    outputs(2222) <= (layer2_outputs(12498)) and (layer2_outputs(10918));
    outputs(2223) <= (layer2_outputs(2599)) and not (layer2_outputs(2575));
    outputs(2224) <= (layer2_outputs(11098)) xor (layer2_outputs(11668));
    outputs(2225) <= (layer2_outputs(4317)) xor (layer2_outputs(11203));
    outputs(2226) <= layer2_outputs(2119);
    outputs(2227) <= not(layer2_outputs(3900));
    outputs(2228) <= not(layer2_outputs(10919));
    outputs(2229) <= not((layer2_outputs(2504)) or (layer2_outputs(8762)));
    outputs(2230) <= (layer2_outputs(3199)) xor (layer2_outputs(8691));
    outputs(2231) <= not(layer2_outputs(8666));
    outputs(2232) <= not(layer2_outputs(12559));
    outputs(2233) <= (layer2_outputs(1722)) and not (layer2_outputs(10602));
    outputs(2234) <= (layer2_outputs(8779)) and not (layer2_outputs(4662));
    outputs(2235) <= (layer2_outputs(6391)) and not (layer2_outputs(7201));
    outputs(2236) <= (layer2_outputs(5427)) and (layer2_outputs(10058));
    outputs(2237) <= (layer2_outputs(2222)) and (layer2_outputs(8532));
    outputs(2238) <= not(layer2_outputs(12215));
    outputs(2239) <= (layer2_outputs(5354)) xor (layer2_outputs(8020));
    outputs(2240) <= not(layer2_outputs(8517));
    outputs(2241) <= (layer2_outputs(8364)) and not (layer2_outputs(4352));
    outputs(2242) <= (layer2_outputs(1172)) xor (layer2_outputs(12024));
    outputs(2243) <= not(layer2_outputs(3708));
    outputs(2244) <= (layer2_outputs(3120)) and not (layer2_outputs(6921));
    outputs(2245) <= not(layer2_outputs(12389));
    outputs(2246) <= (layer2_outputs(401)) and not (layer2_outputs(4671));
    outputs(2247) <= (layer2_outputs(10264)) xor (layer2_outputs(239));
    outputs(2248) <= (layer2_outputs(271)) and not (layer2_outputs(11533));
    outputs(2249) <= layer2_outputs(5599);
    outputs(2250) <= not((layer2_outputs(10112)) xor (layer2_outputs(11344)));
    outputs(2251) <= layer2_outputs(5049);
    outputs(2252) <= not(layer2_outputs(4441));
    outputs(2253) <= not(layer2_outputs(11040));
    outputs(2254) <= layer2_outputs(3838);
    outputs(2255) <= not(layer2_outputs(9614));
    outputs(2256) <= (layer2_outputs(7824)) and not (layer2_outputs(7864));
    outputs(2257) <= not(layer2_outputs(3407));
    outputs(2258) <= not(layer2_outputs(7706));
    outputs(2259) <= not(layer2_outputs(8676));
    outputs(2260) <= not(layer2_outputs(1381));
    outputs(2261) <= layer2_outputs(5597);
    outputs(2262) <= (layer2_outputs(7107)) and not (layer2_outputs(8759));
    outputs(2263) <= layer2_outputs(7403);
    outputs(2264) <= not((layer2_outputs(1608)) xor (layer2_outputs(2886)));
    outputs(2265) <= (layer2_outputs(2117)) xor (layer2_outputs(1906));
    outputs(2266) <= (layer2_outputs(5210)) xor (layer2_outputs(7000));
    outputs(2267) <= (layer2_outputs(1032)) xor (layer2_outputs(6302));
    outputs(2268) <= not((layer2_outputs(6387)) xor (layer2_outputs(4289)));
    outputs(2269) <= (layer2_outputs(5561)) and (layer2_outputs(10386));
    outputs(2270) <= layer2_outputs(1576);
    outputs(2271) <= not((layer2_outputs(10561)) xor (layer2_outputs(8913)));
    outputs(2272) <= not(layer2_outputs(12145));
    outputs(2273) <= not((layer2_outputs(5435)) xor (layer2_outputs(1247)));
    outputs(2274) <= (layer2_outputs(2447)) xor (layer2_outputs(5294));
    outputs(2275) <= layer2_outputs(12201);
    outputs(2276) <= (layer2_outputs(10184)) xor (layer2_outputs(2405));
    outputs(2277) <= not((layer2_outputs(2093)) xor (layer2_outputs(1004)));
    outputs(2278) <= not((layer2_outputs(4522)) xor (layer2_outputs(5945)));
    outputs(2279) <= not(layer2_outputs(11795));
    outputs(2280) <= (layer2_outputs(8749)) xor (layer2_outputs(2005));
    outputs(2281) <= (layer2_outputs(12495)) or (layer2_outputs(8427));
    outputs(2282) <= (layer2_outputs(11270)) xor (layer2_outputs(4576));
    outputs(2283) <= layer2_outputs(1031);
    outputs(2284) <= (layer2_outputs(1847)) or (layer2_outputs(2576));
    outputs(2285) <= not(layer2_outputs(7297)) or (layer2_outputs(8251));
    outputs(2286) <= (layer2_outputs(1847)) or (layer2_outputs(4044));
    outputs(2287) <= not((layer2_outputs(5392)) or (layer2_outputs(5312)));
    outputs(2288) <= layer2_outputs(11276);
    outputs(2289) <= not(layer2_outputs(5194));
    outputs(2290) <= layer2_outputs(6863);
    outputs(2291) <= layer2_outputs(10434);
    outputs(2292) <= (layer2_outputs(12731)) and (layer2_outputs(6669));
    outputs(2293) <= (layer2_outputs(12454)) xor (layer2_outputs(7391));
    outputs(2294) <= (layer2_outputs(1594)) and (layer2_outputs(8269));
    outputs(2295) <= (layer2_outputs(5323)) xor (layer2_outputs(12576));
    outputs(2296) <= layer2_outputs(6326);
    outputs(2297) <= not((layer2_outputs(5646)) and (layer2_outputs(11149)));
    outputs(2298) <= (layer2_outputs(5178)) xor (layer2_outputs(126));
    outputs(2299) <= (layer2_outputs(7908)) xor (layer2_outputs(5082));
    outputs(2300) <= (layer2_outputs(737)) and (layer2_outputs(3902));
    outputs(2301) <= layer2_outputs(658);
    outputs(2302) <= layer2_outputs(9656);
    outputs(2303) <= layer2_outputs(826);
    outputs(2304) <= (layer2_outputs(3749)) xor (layer2_outputs(82));
    outputs(2305) <= not(layer2_outputs(11056));
    outputs(2306) <= not(layer2_outputs(11960));
    outputs(2307) <= (layer2_outputs(2154)) xor (layer2_outputs(10568));
    outputs(2308) <= (layer2_outputs(2616)) xor (layer2_outputs(11823));
    outputs(2309) <= not(layer2_outputs(1161));
    outputs(2310) <= not(layer2_outputs(8477));
    outputs(2311) <= (layer2_outputs(3203)) xor (layer2_outputs(9407));
    outputs(2312) <= not((layer2_outputs(859)) xor (layer2_outputs(8514)));
    outputs(2313) <= (layer2_outputs(1293)) and (layer2_outputs(1886));
    outputs(2314) <= not((layer2_outputs(5426)) xor (layer2_outputs(11192)));
    outputs(2315) <= layer2_outputs(8567);
    outputs(2316) <= not((layer2_outputs(3341)) and (layer2_outputs(1270)));
    outputs(2317) <= (layer2_outputs(3807)) and (layer2_outputs(7149));
    outputs(2318) <= layer2_outputs(10926);
    outputs(2319) <= not(layer2_outputs(3380));
    outputs(2320) <= (layer2_outputs(4034)) xor (layer2_outputs(2013));
    outputs(2321) <= (layer2_outputs(11639)) xor (layer2_outputs(1603));
    outputs(2322) <= layer2_outputs(1470);
    outputs(2323) <= not((layer2_outputs(9373)) xor (layer2_outputs(9098)));
    outputs(2324) <= not(layer2_outputs(5297));
    outputs(2325) <= (layer2_outputs(7675)) xor (layer2_outputs(4211));
    outputs(2326) <= layer2_outputs(8361);
    outputs(2327) <= not(layer2_outputs(3376));
    outputs(2328) <= layer2_outputs(5715);
    outputs(2329) <= not(layer2_outputs(1373));
    outputs(2330) <= (layer2_outputs(5522)) and not (layer2_outputs(169));
    outputs(2331) <= (layer2_outputs(6753)) and not (layer2_outputs(8730));
    outputs(2332) <= (layer2_outputs(576)) xor (layer2_outputs(2045));
    outputs(2333) <= layer2_outputs(9105);
    outputs(2334) <= layer2_outputs(8740);
    outputs(2335) <= not((layer2_outputs(6279)) or (layer2_outputs(7195)));
    outputs(2336) <= (layer2_outputs(3688)) and not (layer2_outputs(2341));
    outputs(2337) <= (layer2_outputs(9339)) and (layer2_outputs(3436));
    outputs(2338) <= not((layer2_outputs(42)) xor (layer2_outputs(6188)));
    outputs(2339) <= not(layer2_outputs(3099));
    outputs(2340) <= (layer2_outputs(12029)) xor (layer2_outputs(9363));
    outputs(2341) <= not(layer2_outputs(9367));
    outputs(2342) <= (layer2_outputs(8629)) and (layer2_outputs(9311));
    outputs(2343) <= layer2_outputs(8341);
    outputs(2344) <= not(layer2_outputs(11298));
    outputs(2345) <= (layer2_outputs(4029)) xor (layer2_outputs(8460));
    outputs(2346) <= layer2_outputs(9946);
    outputs(2347) <= (layer2_outputs(6093)) and (layer2_outputs(1456));
    outputs(2348) <= not(layer2_outputs(11037));
    outputs(2349) <= not(layer2_outputs(11526));
    outputs(2350) <= layer2_outputs(10566);
    outputs(2351) <= layer2_outputs(6232);
    outputs(2352) <= not(layer2_outputs(12241));
    outputs(2353) <= (layer2_outputs(11903)) xor (layer2_outputs(11819));
    outputs(2354) <= not(layer2_outputs(12485));
    outputs(2355) <= not((layer2_outputs(8945)) or (layer2_outputs(11606)));
    outputs(2356) <= layer2_outputs(12502);
    outputs(2357) <= layer2_outputs(12048);
    outputs(2358) <= not(layer2_outputs(4645));
    outputs(2359) <= (layer2_outputs(12782)) xor (layer2_outputs(4872));
    outputs(2360) <= not((layer2_outputs(8134)) or (layer2_outputs(4593)));
    outputs(2361) <= (layer2_outputs(5486)) and not (layer2_outputs(6730));
    outputs(2362) <= (layer2_outputs(8907)) xor (layer2_outputs(11311));
    outputs(2363) <= not(layer2_outputs(9020));
    outputs(2364) <= layer2_outputs(257);
    outputs(2365) <= not(layer2_outputs(1457));
    outputs(2366) <= (layer2_outputs(1393)) and not (layer2_outputs(733));
    outputs(2367) <= (layer2_outputs(11437)) and not (layer2_outputs(8046));
    outputs(2368) <= layer2_outputs(7060);
    outputs(2369) <= not((layer2_outputs(6819)) xor (layer2_outputs(7453)));
    outputs(2370) <= not(layer2_outputs(8072));
    outputs(2371) <= (layer2_outputs(9119)) and not (layer2_outputs(1992));
    outputs(2372) <= (layer2_outputs(11601)) and not (layer2_outputs(10860));
    outputs(2373) <= (layer2_outputs(2527)) xor (layer2_outputs(1707));
    outputs(2374) <= layer2_outputs(4264);
    outputs(2375) <= (layer2_outputs(3479)) and not (layer2_outputs(4955));
    outputs(2376) <= not((layer2_outputs(7475)) xor (layer2_outputs(1915)));
    outputs(2377) <= not((layer2_outputs(3851)) or (layer2_outputs(10602)));
    outputs(2378) <= (layer2_outputs(8286)) and not (layer2_outputs(647));
    outputs(2379) <= (layer2_outputs(3554)) and not (layer2_outputs(57));
    outputs(2380) <= (layer2_outputs(11605)) and (layer2_outputs(1814));
    outputs(2381) <= not((layer2_outputs(9382)) xor (layer2_outputs(5030)));
    outputs(2382) <= not(layer2_outputs(8853));
    outputs(2383) <= (layer2_outputs(4076)) xor (layer2_outputs(5598));
    outputs(2384) <= not((layer2_outputs(8155)) or (layer2_outputs(6317)));
    outputs(2385) <= (layer2_outputs(3980)) and not (layer2_outputs(12050));
    outputs(2386) <= (layer2_outputs(9835)) and not (layer2_outputs(11002));
    outputs(2387) <= (layer2_outputs(4359)) xor (layer2_outputs(12163));
    outputs(2388) <= not(layer2_outputs(1492));
    outputs(2389) <= layer2_outputs(11713);
    outputs(2390) <= (layer2_outputs(9244)) and not (layer2_outputs(4336));
    outputs(2391) <= (layer2_outputs(4267)) xor (layer2_outputs(10624));
    outputs(2392) <= not((layer2_outputs(5399)) and (layer2_outputs(10606)));
    outputs(2393) <= (layer2_outputs(5)) and (layer2_outputs(9941));
    outputs(2394) <= not((layer2_outputs(11186)) or (layer2_outputs(4286)));
    outputs(2395) <= (layer2_outputs(5014)) and not (layer2_outputs(10866));
    outputs(2396) <= layer2_outputs(9566);
    outputs(2397) <= not(layer2_outputs(2276));
    outputs(2398) <= not(layer2_outputs(7730));
    outputs(2399) <= not((layer2_outputs(7361)) or (layer2_outputs(1000)));
    outputs(2400) <= layer2_outputs(3565);
    outputs(2401) <= not((layer2_outputs(12114)) xor (layer2_outputs(12421)));
    outputs(2402) <= layer2_outputs(10078);
    outputs(2403) <= (layer2_outputs(7691)) and not (layer2_outputs(733));
    outputs(2404) <= not(layer2_outputs(10214));
    outputs(2405) <= not(layer2_outputs(9041));
    outputs(2406) <= (layer2_outputs(9281)) or (layer2_outputs(11715));
    outputs(2407) <= (layer2_outputs(5991)) and not (layer2_outputs(9725));
    outputs(2408) <= not(layer2_outputs(10635));
    outputs(2409) <= (layer2_outputs(4028)) or (layer2_outputs(11220));
    outputs(2410) <= not(layer2_outputs(11660));
    outputs(2411) <= not(layer2_outputs(928));
    outputs(2412) <= layer2_outputs(10228);
    outputs(2413) <= not((layer2_outputs(2227)) or (layer2_outputs(11464)));
    outputs(2414) <= not(layer2_outputs(11927));
    outputs(2415) <= (layer2_outputs(5168)) xor (layer2_outputs(10917));
    outputs(2416) <= (layer2_outputs(7424)) and not (layer2_outputs(1317));
    outputs(2417) <= not(layer2_outputs(9213));
    outputs(2418) <= not(layer2_outputs(5125));
    outputs(2419) <= (layer2_outputs(5664)) and not (layer2_outputs(10701));
    outputs(2420) <= not(layer2_outputs(10160));
    outputs(2421) <= layer2_outputs(10044);
    outputs(2422) <= not(layer2_outputs(5303)) or (layer2_outputs(10261));
    outputs(2423) <= not(layer2_outputs(10428));
    outputs(2424) <= layer2_outputs(6660);
    outputs(2425) <= not(layer2_outputs(6856));
    outputs(2426) <= (layer2_outputs(8636)) xor (layer2_outputs(2584));
    outputs(2427) <= (layer2_outputs(574)) xor (layer2_outputs(5827));
    outputs(2428) <= not(layer2_outputs(2791));
    outputs(2429) <= (layer2_outputs(11740)) and not (layer2_outputs(6085));
    outputs(2430) <= (layer2_outputs(11401)) and not (layer2_outputs(9729));
    outputs(2431) <= not((layer2_outputs(8910)) or (layer2_outputs(9554)));
    outputs(2432) <= not(layer2_outputs(5090));
    outputs(2433) <= not(layer2_outputs(10989));
    outputs(2434) <= layer2_outputs(2924);
    outputs(2435) <= layer2_outputs(10758);
    outputs(2436) <= (layer2_outputs(2673)) xor (layer2_outputs(9287));
    outputs(2437) <= not((layer2_outputs(9520)) or (layer2_outputs(5884)));
    outputs(2438) <= (layer2_outputs(8825)) and not (layer2_outputs(10523));
    outputs(2439) <= layer2_outputs(3486);
    outputs(2440) <= (layer2_outputs(6946)) and not (layer2_outputs(5609));
    outputs(2441) <= (layer2_outputs(639)) and not (layer2_outputs(1257));
    outputs(2442) <= not(layer2_outputs(9900));
    outputs(2443) <= (layer2_outputs(6637)) xor (layer2_outputs(8699));
    outputs(2444) <= not(layer2_outputs(5956));
    outputs(2445) <= '0';
    outputs(2446) <= layer2_outputs(5551);
    outputs(2447) <= (layer2_outputs(8310)) xor (layer2_outputs(11557));
    outputs(2448) <= not(layer2_outputs(11767)) or (layer2_outputs(9752));
    outputs(2449) <= not((layer2_outputs(3267)) xor (layer2_outputs(6542)));
    outputs(2450) <= not((layer2_outputs(11070)) xor (layer2_outputs(4771)));
    outputs(2451) <= (layer2_outputs(5905)) and not (layer2_outputs(691));
    outputs(2452) <= not((layer2_outputs(10738)) or (layer2_outputs(3693)));
    outputs(2453) <= (layer2_outputs(7371)) xor (layer2_outputs(6515));
    outputs(2454) <= (layer2_outputs(1917)) and (layer2_outputs(3597));
    outputs(2455) <= not(layer2_outputs(12033));
    outputs(2456) <= not((layer2_outputs(12023)) xor (layer2_outputs(619)));
    outputs(2457) <= (layer2_outputs(9634)) and (layer2_outputs(852));
    outputs(2458) <= not((layer2_outputs(12005)) xor (layer2_outputs(1410)));
    outputs(2459) <= (layer2_outputs(7752)) and (layer2_outputs(5995));
    outputs(2460) <= layer2_outputs(9655);
    outputs(2461) <= (layer2_outputs(9788)) or (layer2_outputs(1679));
    outputs(2462) <= not(layer2_outputs(6344)) or (layer2_outputs(1655));
    outputs(2463) <= not(layer2_outputs(12168));
    outputs(2464) <= layer2_outputs(775);
    outputs(2465) <= (layer2_outputs(12725)) and (layer2_outputs(6161));
    outputs(2466) <= layer2_outputs(2569);
    outputs(2467) <= layer2_outputs(6469);
    outputs(2468) <= not(layer2_outputs(10176));
    outputs(2469) <= layer2_outputs(3173);
    outputs(2470) <= not((layer2_outputs(3834)) or (layer2_outputs(2456)));
    outputs(2471) <= (layer2_outputs(10656)) and not (layer2_outputs(4080));
    outputs(2472) <= (layer2_outputs(6866)) and not (layer2_outputs(8620));
    outputs(2473) <= not(layer2_outputs(9886));
    outputs(2474) <= layer2_outputs(5374);
    outputs(2475) <= layer2_outputs(3043);
    outputs(2476) <= (layer2_outputs(5944)) and not (layer2_outputs(8967));
    outputs(2477) <= not(layer2_outputs(695));
    outputs(2478) <= not(layer2_outputs(12006));
    outputs(2479) <= not((layer2_outputs(361)) xor (layer2_outputs(3435)));
    outputs(2480) <= (layer2_outputs(1009)) and not (layer2_outputs(7186));
    outputs(2481) <= not(layer2_outputs(10387));
    outputs(2482) <= (layer2_outputs(12281)) xor (layer2_outputs(12104));
    outputs(2483) <= (layer2_outputs(3092)) xor (layer2_outputs(12447));
    outputs(2484) <= (layer2_outputs(11444)) xor (layer2_outputs(9105));
    outputs(2485) <= (layer2_outputs(8652)) and not (layer2_outputs(8153));
    outputs(2486) <= (layer2_outputs(6113)) xor (layer2_outputs(9899));
    outputs(2487) <= (layer2_outputs(3738)) and not (layer2_outputs(3756));
    outputs(2488) <= (layer2_outputs(11020)) xor (layer2_outputs(6892));
    outputs(2489) <= not((layer2_outputs(2792)) xor (layer2_outputs(4947)));
    outputs(2490) <= (layer2_outputs(1644)) and not (layer2_outputs(8058));
    outputs(2491) <= (layer2_outputs(8811)) and not (layer2_outputs(11935));
    outputs(2492) <= (layer2_outputs(11969)) xor (layer2_outputs(1739));
    outputs(2493) <= not(layer2_outputs(11711));
    outputs(2494) <= not(layer2_outputs(4142));
    outputs(2495) <= (layer2_outputs(10706)) and (layer2_outputs(3889));
    outputs(2496) <= not((layer2_outputs(9949)) xor (layer2_outputs(991)));
    outputs(2497) <= not((layer2_outputs(11594)) xor (layer2_outputs(8077)));
    outputs(2498) <= not((layer2_outputs(11325)) or (layer2_outputs(5030)));
    outputs(2499) <= (layer2_outputs(2725)) xor (layer2_outputs(2245));
    outputs(2500) <= (layer2_outputs(6838)) and not (layer2_outputs(5136));
    outputs(2501) <= not((layer2_outputs(7682)) xor (layer2_outputs(8896)));
    outputs(2502) <= layer2_outputs(8948);
    outputs(2503) <= not(layer2_outputs(9351));
    outputs(2504) <= not((layer2_outputs(5197)) xor (layer2_outputs(11339)));
    outputs(2505) <= not(layer2_outputs(10955));
    outputs(2506) <= not(layer2_outputs(2487));
    outputs(2507) <= layer2_outputs(6772);
    outputs(2508) <= not((layer2_outputs(3054)) xor (layer2_outputs(1845)));
    outputs(2509) <= not((layer2_outputs(7902)) or (layer2_outputs(6904)));
    outputs(2510) <= (layer2_outputs(6406)) and not (layer2_outputs(7178));
    outputs(2511) <= not((layer2_outputs(12278)) xor (layer2_outputs(7074)));
    outputs(2512) <= not((layer2_outputs(2124)) xor (layer2_outputs(1104)));
    outputs(2513) <= (layer2_outputs(2149)) and not (layer2_outputs(4809));
    outputs(2514) <= not((layer2_outputs(3010)) or (layer2_outputs(4502)));
    outputs(2515) <= not(layer2_outputs(9424));
    outputs(2516) <= (layer2_outputs(7085)) and (layer2_outputs(4076));
    outputs(2517) <= layer2_outputs(7703);
    outputs(2518) <= (layer2_outputs(10074)) and not (layer2_outputs(1171));
    outputs(2519) <= not((layer2_outputs(4523)) xor (layer2_outputs(6510)));
    outputs(2520) <= layer2_outputs(12613);
    outputs(2521) <= not((layer2_outputs(2291)) xor (layer2_outputs(3746)));
    outputs(2522) <= not(layer2_outputs(2206));
    outputs(2523) <= (layer2_outputs(6506)) xor (layer2_outputs(705));
    outputs(2524) <= layer2_outputs(10238);
    outputs(2525) <= not((layer2_outputs(2899)) xor (layer2_outputs(6935)));
    outputs(2526) <= layer2_outputs(38);
    outputs(2527) <= not(layer2_outputs(10277));
    outputs(2528) <= (layer2_outputs(8169)) and not (layer2_outputs(11612));
    outputs(2529) <= (layer2_outputs(8075)) xor (layer2_outputs(6937));
    outputs(2530) <= layer2_outputs(8739);
    outputs(2531) <= (layer2_outputs(8562)) xor (layer2_outputs(2708));
    outputs(2532) <= layer2_outputs(7698);
    outputs(2533) <= (layer2_outputs(1745)) xor (layer2_outputs(3938));
    outputs(2534) <= not((layer2_outputs(3912)) xor (layer2_outputs(8818)));
    outputs(2535) <= layer2_outputs(4689);
    outputs(2536) <= layer2_outputs(203);
    outputs(2537) <= not((layer2_outputs(2350)) and (layer2_outputs(3470)));
    outputs(2538) <= not((layer2_outputs(2173)) or (layer2_outputs(8158)));
    outputs(2539) <= (layer2_outputs(4412)) and not (layer2_outputs(9699));
    outputs(2540) <= not((layer2_outputs(470)) and (layer2_outputs(1070)));
    outputs(2541) <= layer2_outputs(6751);
    outputs(2542) <= not((layer2_outputs(4022)) xor (layer2_outputs(9719)));
    outputs(2543) <= (layer2_outputs(9879)) xor (layer2_outputs(3494));
    outputs(2544) <= layer2_outputs(5242);
    outputs(2545) <= not((layer2_outputs(503)) xor (layer2_outputs(10460)));
    outputs(2546) <= layer2_outputs(3942);
    outputs(2547) <= not(layer2_outputs(3715)) or (layer2_outputs(7527));
    outputs(2548) <= not((layer2_outputs(1817)) xor (layer2_outputs(5753)));
    outputs(2549) <= (layer2_outputs(4246)) xor (layer2_outputs(10992));
    outputs(2550) <= not((layer2_outputs(11282)) or (layer2_outputs(748)));
    outputs(2551) <= not((layer2_outputs(1088)) xor (layer2_outputs(3187)));
    outputs(2552) <= (layer2_outputs(5149)) xor (layer2_outputs(36));
    outputs(2553) <= not((layer2_outputs(9363)) xor (layer2_outputs(4608)));
    outputs(2554) <= layer2_outputs(5112);
    outputs(2555) <= not((layer2_outputs(6447)) xor (layer2_outputs(10487)));
    outputs(2556) <= not((layer2_outputs(2369)) xor (layer2_outputs(10162)));
    outputs(2557) <= not(layer2_outputs(11382));
    outputs(2558) <= layer2_outputs(7509);
    outputs(2559) <= not(layer2_outputs(11620));
    outputs(2560) <= not(layer2_outputs(7056));
    outputs(2561) <= layer2_outputs(9161);
    outputs(2562) <= not((layer2_outputs(11194)) xor (layer2_outputs(4170)));
    outputs(2563) <= (layer2_outputs(4406)) and (layer2_outputs(10265));
    outputs(2564) <= not(layer2_outputs(7807)) or (layer2_outputs(491));
    outputs(2565) <= not(layer2_outputs(11094));
    outputs(2566) <= layer2_outputs(3000);
    outputs(2567) <= not((layer2_outputs(7395)) xor (layer2_outputs(11946)));
    outputs(2568) <= (layer2_outputs(1167)) xor (layer2_outputs(2732));
    outputs(2569) <= not(layer2_outputs(6594));
    outputs(2570) <= layer2_outputs(3925);
    outputs(2571) <= not(layer2_outputs(1206)) or (layer2_outputs(10447));
    outputs(2572) <= not(layer2_outputs(1653));
    outputs(2573) <= layer2_outputs(1172);
    outputs(2574) <= not((layer2_outputs(11950)) and (layer2_outputs(1532)));
    outputs(2575) <= (layer2_outputs(886)) and (layer2_outputs(7852));
    outputs(2576) <= not((layer2_outputs(1474)) xor (layer2_outputs(5973)));
    outputs(2577) <= not((layer2_outputs(3491)) xor (layer2_outputs(3242)));
    outputs(2578) <= not(layer2_outputs(11106));
    outputs(2579) <= not(layer2_outputs(9156)) or (layer2_outputs(2052));
    outputs(2580) <= not(layer2_outputs(1179));
    outputs(2581) <= (layer2_outputs(8239)) or (layer2_outputs(9753));
    outputs(2582) <= layer2_outputs(6353);
    outputs(2583) <= (layer2_outputs(1841)) or (layer2_outputs(732));
    outputs(2584) <= not(layer2_outputs(6157));
    outputs(2585) <= not((layer2_outputs(3443)) xor (layer2_outputs(2788)));
    outputs(2586) <= not(layer2_outputs(2851));
    outputs(2587) <= not(layer2_outputs(10835)) or (layer2_outputs(2714));
    outputs(2588) <= (layer2_outputs(12412)) xor (layer2_outputs(7994));
    outputs(2589) <= not((layer2_outputs(5966)) xor (layer2_outputs(3595)));
    outputs(2590) <= layer2_outputs(7174);
    outputs(2591) <= not(layer2_outputs(10458));
    outputs(2592) <= not(layer2_outputs(9084));
    outputs(2593) <= not(layer2_outputs(2870));
    outputs(2594) <= not(layer2_outputs(5338)) or (layer2_outputs(6552));
    outputs(2595) <= not(layer2_outputs(2586));
    outputs(2596) <= layer2_outputs(648);
    outputs(2597) <= layer2_outputs(4808);
    outputs(2598) <= (layer2_outputs(12121)) and not (layer2_outputs(10040));
    outputs(2599) <= not(layer2_outputs(1937));
    outputs(2600) <= not(layer2_outputs(7124));
    outputs(2601) <= not((layer2_outputs(7960)) or (layer2_outputs(1338)));
    outputs(2602) <= not((layer2_outputs(7184)) xor (layer2_outputs(6809)));
    outputs(2603) <= not(layer2_outputs(8291));
    outputs(2604) <= not((layer2_outputs(9174)) xor (layer2_outputs(3052)));
    outputs(2605) <= (layer2_outputs(7454)) xor (layer2_outputs(1712));
    outputs(2606) <= not(layer2_outputs(8077)) or (layer2_outputs(5602));
    outputs(2607) <= layer2_outputs(3222);
    outputs(2608) <= not(layer2_outputs(4455));
    outputs(2609) <= layer2_outputs(8638);
    outputs(2610) <= not(layer2_outputs(3713)) or (layer2_outputs(519));
    outputs(2611) <= (layer2_outputs(354)) xor (layer2_outputs(3933));
    outputs(2612) <= (layer2_outputs(9510)) and (layer2_outputs(9973));
    outputs(2613) <= not((layer2_outputs(6828)) xor (layer2_outputs(2887)));
    outputs(2614) <= (layer2_outputs(10820)) and not (layer2_outputs(1292));
    outputs(2615) <= not((layer2_outputs(8771)) xor (layer2_outputs(12491)));
    outputs(2616) <= not(layer2_outputs(53));
    outputs(2617) <= layer2_outputs(7556);
    outputs(2618) <= not((layer2_outputs(6160)) or (layer2_outputs(9583)));
    outputs(2619) <= not(layer2_outputs(9538));
    outputs(2620) <= not((layer2_outputs(3402)) xor (layer2_outputs(618)));
    outputs(2621) <= layer2_outputs(6523);
    outputs(2622) <= layer2_outputs(1868);
    outputs(2623) <= (layer2_outputs(6154)) xor (layer2_outputs(5548));
    outputs(2624) <= not((layer2_outputs(3304)) xor (layer2_outputs(7394)));
    outputs(2625) <= layer2_outputs(5004);
    outputs(2626) <= (layer2_outputs(3151)) or (layer2_outputs(2217));
    outputs(2627) <= not(layer2_outputs(1229));
    outputs(2628) <= not(layer2_outputs(7558));
    outputs(2629) <= (layer2_outputs(10657)) xor (layer2_outputs(11267));
    outputs(2630) <= layer2_outputs(4483);
    outputs(2631) <= not(layer2_outputs(2481));
    outputs(2632) <= not(layer2_outputs(4231));
    outputs(2633) <= layer2_outputs(4592);
    outputs(2634) <= (layer2_outputs(11867)) xor (layer2_outputs(9659));
    outputs(2635) <= not(layer2_outputs(4258));
    outputs(2636) <= layer2_outputs(12587);
    outputs(2637) <= not((layer2_outputs(12683)) xor (layer2_outputs(6701)));
    outputs(2638) <= layer2_outputs(6041);
    outputs(2639) <= not(layer2_outputs(2253));
    outputs(2640) <= not(layer2_outputs(11265));
    outputs(2641) <= not((layer2_outputs(12312)) xor (layer2_outputs(7853)));
    outputs(2642) <= layer2_outputs(9195);
    outputs(2643) <= not((layer2_outputs(3600)) xor (layer2_outputs(7020)));
    outputs(2644) <= not(layer2_outputs(12578));
    outputs(2645) <= not(layer2_outputs(3265)) or (layer2_outputs(2131));
    outputs(2646) <= layer2_outputs(12146);
    outputs(2647) <= not((layer2_outputs(558)) xor (layer2_outputs(9436)));
    outputs(2648) <= not(layer2_outputs(1726));
    outputs(2649) <= not(layer2_outputs(5990));
    outputs(2650) <= (layer2_outputs(8195)) and not (layer2_outputs(2068));
    outputs(2651) <= not(layer2_outputs(6734));
    outputs(2652) <= not((layer2_outputs(6569)) xor (layer2_outputs(7943)));
    outputs(2653) <= not(layer2_outputs(8060)) or (layer2_outputs(3487));
    outputs(2654) <= not(layer2_outputs(9340)) or (layer2_outputs(11566));
    outputs(2655) <= layer2_outputs(11915);
    outputs(2656) <= (layer2_outputs(9964)) or (layer2_outputs(10941));
    outputs(2657) <= not(layer2_outputs(8824));
    outputs(2658) <= not(layer2_outputs(9766));
    outputs(2659) <= not(layer2_outputs(11418));
    outputs(2660) <= not(layer2_outputs(11992));
    outputs(2661) <= (layer2_outputs(1511)) and not (layer2_outputs(146));
    outputs(2662) <= not((layer2_outputs(3076)) xor (layer2_outputs(11383)));
    outputs(2663) <= not((layer2_outputs(2192)) xor (layer2_outputs(11272)));
    outputs(2664) <= not((layer2_outputs(1286)) xor (layer2_outputs(723)));
    outputs(2665) <= (layer2_outputs(918)) or (layer2_outputs(2480));
    outputs(2666) <= (layer2_outputs(3245)) xor (layer2_outputs(2211));
    outputs(2667) <= layer2_outputs(11386);
    outputs(2668) <= layer2_outputs(5002);
    outputs(2669) <= not(layer2_outputs(7088));
    outputs(2670) <= not(layer2_outputs(2136));
    outputs(2671) <= not(layer2_outputs(10531));
    outputs(2672) <= (layer2_outputs(5938)) xor (layer2_outputs(6321));
    outputs(2673) <= layer2_outputs(4698);
    outputs(2674) <= not(layer2_outputs(1600));
    outputs(2675) <= layer2_outputs(7793);
    outputs(2676) <= not(layer2_outputs(3851));
    outputs(2677) <= (layer2_outputs(6662)) xor (layer2_outputs(12644));
    outputs(2678) <= not((layer2_outputs(1154)) xor (layer2_outputs(8960)));
    outputs(2679) <= not(layer2_outputs(4714)) or (layer2_outputs(8822));
    outputs(2680) <= not(layer2_outputs(8284)) or (layer2_outputs(3496));
    outputs(2681) <= (layer2_outputs(2805)) xor (layer2_outputs(566));
    outputs(2682) <= layer2_outputs(12518);
    outputs(2683) <= not((layer2_outputs(12706)) xor (layer2_outputs(7059)));
    outputs(2684) <= not(layer2_outputs(6111));
    outputs(2685) <= not(layer2_outputs(10961));
    outputs(2686) <= not(layer2_outputs(11564));
    outputs(2687) <= (layer2_outputs(1445)) and (layer2_outputs(6968));
    outputs(2688) <= layer2_outputs(9294);
    outputs(2689) <= not(layer2_outputs(6571));
    outputs(2690) <= layer2_outputs(4188);
    outputs(2691) <= (layer2_outputs(2973)) xor (layer2_outputs(2559));
    outputs(2692) <= not(layer2_outputs(7796));
    outputs(2693) <= (layer2_outputs(6807)) xor (layer2_outputs(750));
    outputs(2694) <= layer2_outputs(2032);
    outputs(2695) <= layer2_outputs(9421);
    outputs(2696) <= not((layer2_outputs(10692)) and (layer2_outputs(7637)));
    outputs(2697) <= not(layer2_outputs(9723));
    outputs(2698) <= not((layer2_outputs(8891)) and (layer2_outputs(12486)));
    outputs(2699) <= layer2_outputs(10332);
    outputs(2700) <= (layer2_outputs(3164)) or (layer2_outputs(10454));
    outputs(2701) <= (layer2_outputs(8334)) and (layer2_outputs(10580));
    outputs(2702) <= not(layer2_outputs(4292)) or (layer2_outputs(11530));
    outputs(2703) <= (layer2_outputs(1003)) and (layer2_outputs(9198));
    outputs(2704) <= not((layer2_outputs(10605)) xor (layer2_outputs(3810)));
    outputs(2705) <= layer2_outputs(4663);
    outputs(2706) <= layer2_outputs(11607);
    outputs(2707) <= not(layer2_outputs(2308));
    outputs(2708) <= (layer2_outputs(11239)) or (layer2_outputs(10190));
    outputs(2709) <= not(layer2_outputs(9863)) or (layer2_outputs(604));
    outputs(2710) <= not(layer2_outputs(7733));
    outputs(2711) <= not(layer2_outputs(5639));
    outputs(2712) <= not(layer2_outputs(2615));
    outputs(2713) <= not(layer2_outputs(7182));
    outputs(2714) <= not(layer2_outputs(8482));
    outputs(2715) <= layer2_outputs(11405);
    outputs(2716) <= layer2_outputs(3967);
    outputs(2717) <= not((layer2_outputs(1756)) xor (layer2_outputs(7549)));
    outputs(2718) <= (layer2_outputs(3532)) or (layer2_outputs(4811));
    outputs(2719) <= (layer2_outputs(8118)) and not (layer2_outputs(11488));
    outputs(2720) <= not(layer2_outputs(7464));
    outputs(2721) <= not((layer2_outputs(11390)) and (layer2_outputs(1994)));
    outputs(2722) <= layer2_outputs(4616);
    outputs(2723) <= layer2_outputs(12660);
    outputs(2724) <= not((layer2_outputs(6271)) xor (layer2_outputs(3704)));
    outputs(2725) <= layer2_outputs(7422);
    outputs(2726) <= not(layer2_outputs(9486));
    outputs(2727) <= layer2_outputs(2553);
    outputs(2728) <= not(layer2_outputs(1189));
    outputs(2729) <= not((layer2_outputs(2380)) xor (layer2_outputs(3325)));
    outputs(2730) <= layer2_outputs(2043);
    outputs(2731) <= layer2_outputs(9166);
    outputs(2732) <= layer2_outputs(12099);
    outputs(2733) <= not(layer2_outputs(12206));
    outputs(2734) <= not(layer2_outputs(3065));
    outputs(2735) <= (layer2_outputs(6086)) xor (layer2_outputs(12242));
    outputs(2736) <= not(layer2_outputs(889));
    outputs(2737) <= not(layer2_outputs(6943));
    outputs(2738) <= not((layer2_outputs(2408)) or (layer2_outputs(3678)));
    outputs(2739) <= (layer2_outputs(3844)) and (layer2_outputs(8113));
    outputs(2740) <= layer2_outputs(12398);
    outputs(2741) <= (layer2_outputs(476)) xor (layer2_outputs(10599));
    outputs(2742) <= not(layer2_outputs(6538));
    outputs(2743) <= layer2_outputs(1964);
    outputs(2744) <= not((layer2_outputs(8938)) xor (layer2_outputs(11858)));
    outputs(2745) <= (layer2_outputs(5325)) xor (layer2_outputs(10529));
    outputs(2746) <= layer2_outputs(3550);
    outputs(2747) <= not(layer2_outputs(4831));
    outputs(2748) <= not((layer2_outputs(3971)) or (layer2_outputs(874)));
    outputs(2749) <= layer2_outputs(7704);
    outputs(2750) <= not((layer2_outputs(12157)) and (layer2_outputs(23)));
    outputs(2751) <= not((layer2_outputs(11965)) xor (layer2_outputs(8930)));
    outputs(2752) <= layer2_outputs(5428);
    outputs(2753) <= not((layer2_outputs(6865)) xor (layer2_outputs(5403)));
    outputs(2754) <= layer2_outputs(3744);
    outputs(2755) <= not(layer2_outputs(381));
    outputs(2756) <= not(layer2_outputs(4276));
    outputs(2757) <= not(layer2_outputs(7469));
    outputs(2758) <= (layer2_outputs(12077)) and (layer2_outputs(6797));
    outputs(2759) <= (layer2_outputs(3011)) or (layer2_outputs(1829));
    outputs(2760) <= layer2_outputs(4005);
    outputs(2761) <= layer2_outputs(7188);
    outputs(2762) <= not(layer2_outputs(12520)) or (layer2_outputs(11633));
    outputs(2763) <= (layer2_outputs(11765)) and not (layer2_outputs(4574));
    outputs(2764) <= layer2_outputs(1638);
    outputs(2765) <= layer2_outputs(5766);
    outputs(2766) <= not((layer2_outputs(5036)) xor (layer2_outputs(12404)));
    outputs(2767) <= not((layer2_outputs(8867)) and (layer2_outputs(10132)));
    outputs(2768) <= (layer2_outputs(9808)) and not (layer2_outputs(1303));
    outputs(2769) <= not(layer2_outputs(2906)) or (layer2_outputs(3559));
    outputs(2770) <= not((layer2_outputs(175)) or (layer2_outputs(8829)));
    outputs(2771) <= not(layer2_outputs(3225));
    outputs(2772) <= (layer2_outputs(4404)) and not (layer2_outputs(6154));
    outputs(2773) <= not(layer2_outputs(6551));
    outputs(2774) <= not((layer2_outputs(4657)) xor (layer2_outputs(10837)));
    outputs(2775) <= not(layer2_outputs(5510)) or (layer2_outputs(4187));
    outputs(2776) <= (layer2_outputs(6574)) and not (layer2_outputs(10156));
    outputs(2777) <= not(layer2_outputs(4495));
    outputs(2778) <= not(layer2_outputs(1244));
    outputs(2779) <= (layer2_outputs(1155)) xor (layer2_outputs(9764));
    outputs(2780) <= not(layer2_outputs(8703)) or (layer2_outputs(9211));
    outputs(2781) <= not((layer2_outputs(5492)) xor (layer2_outputs(62)));
    outputs(2782) <= not((layer2_outputs(3169)) xor (layer2_outputs(3446)));
    outputs(2783) <= not((layer2_outputs(10376)) xor (layer2_outputs(2958)));
    outputs(2784) <= not(layer2_outputs(5661));
    outputs(2785) <= not(layer2_outputs(8918)) or (layer2_outputs(6531));
    outputs(2786) <= not(layer2_outputs(5374));
    outputs(2787) <= (layer2_outputs(5808)) xor (layer2_outputs(9811));
    outputs(2788) <= layer2_outputs(5393);
    outputs(2789) <= layer2_outputs(8500);
    outputs(2790) <= layer2_outputs(7955);
    outputs(2791) <= (layer2_outputs(5041)) and (layer2_outputs(7738));
    outputs(2792) <= (layer2_outputs(7547)) or (layer2_outputs(4786));
    outputs(2793) <= not(layer2_outputs(7678));
    outputs(2794) <= layer2_outputs(3306);
    outputs(2795) <= not((layer2_outputs(4482)) xor (layer2_outputs(9732)));
    outputs(2796) <= layer2_outputs(380);
    outputs(2797) <= layer2_outputs(6287);
    outputs(2798) <= layer2_outputs(1470);
    outputs(2799) <= layer2_outputs(9590);
    outputs(2800) <= layer2_outputs(5714);
    outputs(2801) <= not(layer2_outputs(6498));
    outputs(2802) <= (layer2_outputs(8302)) and not (layer2_outputs(2376));
    outputs(2803) <= layer2_outputs(9592);
    outputs(2804) <= not(layer2_outputs(4561));
    outputs(2805) <= (layer2_outputs(1364)) xor (layer2_outputs(3249));
    outputs(2806) <= not(layer2_outputs(10944)) or (layer2_outputs(6290));
    outputs(2807) <= layer2_outputs(8032);
    outputs(2808) <= not(layer2_outputs(12057));
    outputs(2809) <= (layer2_outputs(2635)) and (layer2_outputs(11585));
    outputs(2810) <= not(layer2_outputs(5069));
    outputs(2811) <= not((layer2_outputs(197)) xor (layer2_outputs(9746)));
    outputs(2812) <= not(layer2_outputs(2688));
    outputs(2813) <= not(layer2_outputs(6042)) or (layer2_outputs(8725));
    outputs(2814) <= (layer2_outputs(8332)) xor (layer2_outputs(7312));
    outputs(2815) <= layer2_outputs(7823);
    outputs(2816) <= not(layer2_outputs(230));
    outputs(2817) <= not(layer2_outputs(759)) or (layer2_outputs(6027));
    outputs(2818) <= not((layer2_outputs(1375)) xor (layer2_outputs(2723)));
    outputs(2819) <= (layer2_outputs(10204)) or (layer2_outputs(6826));
    outputs(2820) <= (layer2_outputs(7890)) xor (layer2_outputs(11930));
    outputs(2821) <= (layer2_outputs(11146)) and not (layer2_outputs(8238));
    outputs(2822) <= layer2_outputs(4394);
    outputs(2823) <= (layer2_outputs(5579)) xor (layer2_outputs(2841));
    outputs(2824) <= (layer2_outputs(9251)) or (layer2_outputs(11738));
    outputs(2825) <= layer2_outputs(3178);
    outputs(2826) <= not(layer2_outputs(9766));
    outputs(2827) <= not((layer2_outputs(11395)) and (layer2_outputs(5676)));
    outputs(2828) <= (layer2_outputs(12631)) and not (layer2_outputs(9399));
    outputs(2829) <= not((layer2_outputs(12079)) and (layer2_outputs(8160)));
    outputs(2830) <= not(layer2_outputs(2637));
    outputs(2831) <= not(layer2_outputs(2280));
    outputs(2832) <= not((layer2_outputs(6452)) xor (layer2_outputs(1624)));
    outputs(2833) <= not(layer2_outputs(12491));
    outputs(2834) <= not(layer2_outputs(5200));
    outputs(2835) <= not(layer2_outputs(9341));
    outputs(2836) <= (layer2_outputs(3969)) xor (layer2_outputs(3417));
    outputs(2837) <= not(layer2_outputs(7531)) or (layer2_outputs(3976));
    outputs(2838) <= (layer2_outputs(1774)) or (layer2_outputs(5690));
    outputs(2839) <= (layer2_outputs(861)) or (layer2_outputs(6619));
    outputs(2840) <= layer2_outputs(6849);
    outputs(2841) <= not((layer2_outputs(320)) xor (layer2_outputs(4378)));
    outputs(2842) <= not(layer2_outputs(3602));
    outputs(2843) <= not(layer2_outputs(6352));
    outputs(2844) <= not(layer2_outputs(833));
    outputs(2845) <= not(layer2_outputs(5868));
    outputs(2846) <= layer2_outputs(11739);
    outputs(2847) <= not(layer2_outputs(3048)) or (layer2_outputs(9768));
    outputs(2848) <= not(layer2_outputs(1285));
    outputs(2849) <= layer2_outputs(1547);
    outputs(2850) <= not(layer2_outputs(1466));
    outputs(2851) <= (layer2_outputs(12306)) xor (layer2_outputs(3620));
    outputs(2852) <= layer2_outputs(9566);
    outputs(2853) <= not(layer2_outputs(11999));
    outputs(2854) <= layer2_outputs(7863);
    outputs(2855) <= not((layer2_outputs(7185)) xor (layer2_outputs(9452)));
    outputs(2856) <= layer2_outputs(9235);
    outputs(2857) <= layer2_outputs(320);
    outputs(2858) <= (layer2_outputs(4000)) and (layer2_outputs(4052));
    outputs(2859) <= not((layer2_outputs(5302)) xor (layer2_outputs(11294)));
    outputs(2860) <= not((layer2_outputs(7158)) xor (layer2_outputs(8846)));
    outputs(2861) <= not((layer2_outputs(10757)) xor (layer2_outputs(3614)));
    outputs(2862) <= not((layer2_outputs(5972)) xor (layer2_outputs(12571)));
    outputs(2863) <= layer2_outputs(5859);
    outputs(2864) <= not((layer2_outputs(6149)) xor (layer2_outputs(10230)));
    outputs(2865) <= not(layer2_outputs(6318));
    outputs(2866) <= not(layer2_outputs(854));
    outputs(2867) <= not((layer2_outputs(1386)) xor (layer2_outputs(8265)));
    outputs(2868) <= layer2_outputs(9122);
    outputs(2869) <= not((layer2_outputs(11698)) xor (layer2_outputs(8033)));
    outputs(2870) <= (layer2_outputs(8234)) and not (layer2_outputs(9094));
    outputs(2871) <= layer2_outputs(8024);
    outputs(2872) <= (layer2_outputs(3587)) and not (layer2_outputs(10021));
    outputs(2873) <= layer2_outputs(1294);
    outputs(2874) <= (layer2_outputs(9773)) xor (layer2_outputs(11910));
    outputs(2875) <= not(layer2_outputs(2659));
    outputs(2876) <= not(layer2_outputs(6003));
    outputs(2877) <= not(layer2_outputs(12575)) or (layer2_outputs(794));
    outputs(2878) <= not((layer2_outputs(10973)) and (layer2_outputs(7148)));
    outputs(2879) <= layer2_outputs(11711);
    outputs(2880) <= layer2_outputs(3294);
    outputs(2881) <= layer2_outputs(9448);
    outputs(2882) <= (layer2_outputs(4356)) or (layer2_outputs(4616));
    outputs(2883) <= layer2_outputs(4869);
    outputs(2884) <= layer2_outputs(11823);
    outputs(2885) <= layer2_outputs(12087);
    outputs(2886) <= (layer2_outputs(7583)) xor (layer2_outputs(4921));
    outputs(2887) <= not((layer2_outputs(3421)) xor (layer2_outputs(4998)));
    outputs(2888) <= not((layer2_outputs(2725)) xor (layer2_outputs(6528)));
    outputs(2889) <= not(layer2_outputs(1330));
    outputs(2890) <= not((layer2_outputs(896)) and (layer2_outputs(8273)));
    outputs(2891) <= not(layer2_outputs(12293));
    outputs(2892) <= not(layer2_outputs(9930)) or (layer2_outputs(480));
    outputs(2893) <= layer2_outputs(1687);
    outputs(2894) <= layer2_outputs(11208);
    outputs(2895) <= not((layer2_outputs(10952)) and (layer2_outputs(10360)));
    outputs(2896) <= (layer2_outputs(7314)) and not (layer2_outputs(6320));
    outputs(2897) <= (layer2_outputs(9536)) and not (layer2_outputs(1265));
    outputs(2898) <= (layer2_outputs(11154)) xor (layer2_outputs(1607));
    outputs(2899) <= layer2_outputs(3396);
    outputs(2900) <= not(layer2_outputs(2951));
    outputs(2901) <= (layer2_outputs(9269)) xor (layer2_outputs(12562));
    outputs(2902) <= not(layer2_outputs(7858));
    outputs(2903) <= layer2_outputs(610);
    outputs(2904) <= layer2_outputs(4059);
    outputs(2905) <= not((layer2_outputs(1673)) xor (layer2_outputs(2128)));
    outputs(2906) <= not(layer2_outputs(10335));
    outputs(2907) <= not(layer2_outputs(3857));
    outputs(2908) <= (layer2_outputs(1082)) xor (layer2_outputs(10027));
    outputs(2909) <= (layer2_outputs(8185)) xor (layer2_outputs(11431));
    outputs(2910) <= (layer2_outputs(8905)) xor (layer2_outputs(4918));
    outputs(2911) <= not((layer2_outputs(9835)) xor (layer2_outputs(11374)));
    outputs(2912) <= not((layer2_outputs(9746)) or (layer2_outputs(4199)));
    outputs(2913) <= not(layer2_outputs(10426)) or (layer2_outputs(7842));
    outputs(2914) <= not(layer2_outputs(3689));
    outputs(2915) <= layer2_outputs(10683);
    outputs(2916) <= not(layer2_outputs(8508));
    outputs(2917) <= (layer2_outputs(8070)) and not (layer2_outputs(11497));
    outputs(2918) <= not(layer2_outputs(1838));
    outputs(2919) <= (layer2_outputs(3681)) xor (layer2_outputs(3877));
    outputs(2920) <= layer2_outputs(4585);
    outputs(2921) <= layer2_outputs(9325);
    outputs(2922) <= layer2_outputs(8012);
    outputs(2923) <= (layer2_outputs(5455)) xor (layer2_outputs(3788));
    outputs(2924) <= layer2_outputs(6900);
    outputs(2925) <= not((layer2_outputs(2979)) xor (layer2_outputs(7571)));
    outputs(2926) <= layer2_outputs(11042);
    outputs(2927) <= not(layer2_outputs(12544));
    outputs(2928) <= not((layer2_outputs(3846)) xor (layer2_outputs(8331)));
    outputs(2929) <= not((layer2_outputs(6454)) or (layer2_outputs(9278)));
    outputs(2930) <= layer2_outputs(6278);
    outputs(2931) <= not((layer2_outputs(4650)) xor (layer2_outputs(2215)));
    outputs(2932) <= not(layer2_outputs(12655));
    outputs(2933) <= not(layer2_outputs(6966));
    outputs(2934) <= layer2_outputs(1758);
    outputs(2935) <= not(layer2_outputs(8927));
    outputs(2936) <= not(layer2_outputs(912));
    outputs(2937) <= (layer2_outputs(1747)) and not (layer2_outputs(11285));
    outputs(2938) <= (layer2_outputs(9219)) xor (layer2_outputs(5628));
    outputs(2939) <= layer2_outputs(10984);
    outputs(2940) <= layer2_outputs(6189);
    outputs(2941) <= not((layer2_outputs(10118)) xor (layer2_outputs(6796)));
    outputs(2942) <= not(layer2_outputs(1418));
    outputs(2943) <= not(layer2_outputs(9022));
    outputs(2944) <= layer2_outputs(1044);
    outputs(2945) <= not(layer2_outputs(4665));
    outputs(2946) <= layer2_outputs(1694);
    outputs(2947) <= not((layer2_outputs(11884)) xor (layer2_outputs(2019)));
    outputs(2948) <= layer2_outputs(1735);
    outputs(2949) <= not(layer2_outputs(11107));
    outputs(2950) <= not(layer2_outputs(1209));
    outputs(2951) <= not(layer2_outputs(12580));
    outputs(2952) <= not(layer2_outputs(8351));
    outputs(2953) <= not(layer2_outputs(10348));
    outputs(2954) <= not(layer2_outputs(3439));
    outputs(2955) <= layer2_outputs(6999);
    outputs(2956) <= not(layer2_outputs(12037));
    outputs(2957) <= layer2_outputs(2633);
    outputs(2958) <= not(layer2_outputs(11992));
    outputs(2959) <= not(layer2_outputs(10821));
    outputs(2960) <= layer2_outputs(909);
    outputs(2961) <= (layer2_outputs(8401)) xor (layer2_outputs(1357));
    outputs(2962) <= not((layer2_outputs(8771)) xor (layer2_outputs(316)));
    outputs(2963) <= layer2_outputs(6341);
    outputs(2964) <= layer2_outputs(10776);
    outputs(2965) <= layer2_outputs(513);
    outputs(2966) <= layer2_outputs(7537);
    outputs(2967) <= not(layer2_outputs(2351));
    outputs(2968) <= (layer2_outputs(2676)) and (layer2_outputs(7938));
    outputs(2969) <= (layer2_outputs(240)) xor (layer2_outputs(6718));
    outputs(2970) <= layer2_outputs(11348);
    outputs(2971) <= layer2_outputs(7422);
    outputs(2972) <= not(layer2_outputs(588));
    outputs(2973) <= not(layer2_outputs(1726));
    outputs(2974) <= not((layer2_outputs(10484)) xor (layer2_outputs(9442)));
    outputs(2975) <= (layer2_outputs(8968)) xor (layer2_outputs(9771));
    outputs(2976) <= not(layer2_outputs(4521));
    outputs(2977) <= not(layer2_outputs(7971));
    outputs(2978) <= not(layer2_outputs(7876));
    outputs(2979) <= not((layer2_outputs(10472)) xor (layer2_outputs(9964)));
    outputs(2980) <= not(layer2_outputs(7466));
    outputs(2981) <= not(layer2_outputs(11872));
    outputs(2982) <= not(layer2_outputs(4750));
    outputs(2983) <= not(layer2_outputs(12770));
    outputs(2984) <= not(layer2_outputs(2357));
    outputs(2985) <= not(layer2_outputs(11127));
    outputs(2986) <= layer2_outputs(1510);
    outputs(2987) <= layer2_outputs(939);
    outputs(2988) <= layer2_outputs(11334);
    outputs(2989) <= not(layer2_outputs(3986));
    outputs(2990) <= layer2_outputs(10256);
    outputs(2991) <= layer2_outputs(3519);
    outputs(2992) <= layer2_outputs(4269);
    outputs(2993) <= not((layer2_outputs(3643)) xor (layer2_outputs(1134)));
    outputs(2994) <= layer2_outputs(12382);
    outputs(2995) <= not(layer2_outputs(10397)) or (layer2_outputs(4548));
    outputs(2996) <= not((layer2_outputs(11054)) xor (layer2_outputs(6105)));
    outputs(2997) <= not(layer2_outputs(8835));
    outputs(2998) <= (layer2_outputs(5970)) xor (layer2_outputs(1056));
    outputs(2999) <= not(layer2_outputs(9928));
    outputs(3000) <= layer2_outputs(3906);
    outputs(3001) <= not((layer2_outputs(8049)) xor (layer2_outputs(7675)));
    outputs(3002) <= not((layer2_outputs(9814)) and (layer2_outputs(1280)));
    outputs(3003) <= not(layer2_outputs(3426));
    outputs(3004) <= (layer2_outputs(8903)) and not (layer2_outputs(5369));
    outputs(3005) <= not(layer2_outputs(1112));
    outputs(3006) <= not(layer2_outputs(11508));
    outputs(3007) <= not((layer2_outputs(33)) xor (layer2_outputs(1801)));
    outputs(3008) <= (layer2_outputs(816)) xor (layer2_outputs(10924));
    outputs(3009) <= (layer2_outputs(8335)) and not (layer2_outputs(1304));
    outputs(3010) <= layer2_outputs(4959);
    outputs(3011) <= not(layer2_outputs(3776));
    outputs(3012) <= not(layer2_outputs(1466));
    outputs(3013) <= not(layer2_outputs(12138));
    outputs(3014) <= not(layer2_outputs(9981));
    outputs(3015) <= not(layer2_outputs(11884));
    outputs(3016) <= (layer2_outputs(10875)) xor (layer2_outputs(4350));
    outputs(3017) <= (layer2_outputs(362)) or (layer2_outputs(6451));
    outputs(3018) <= layer2_outputs(8445);
    outputs(3019) <= layer2_outputs(1662);
    outputs(3020) <= not(layer2_outputs(8227));
    outputs(3021) <= not((layer2_outputs(637)) xor (layer2_outputs(7263)));
    outputs(3022) <= (layer2_outputs(11395)) xor (layer2_outputs(1432));
    outputs(3023) <= layer2_outputs(11302);
    outputs(3024) <= (layer2_outputs(12297)) or (layer2_outputs(12733));
    outputs(3025) <= (layer2_outputs(10322)) xor (layer2_outputs(4295));
    outputs(3026) <= layer2_outputs(5208);
    outputs(3027) <= not(layer2_outputs(1490));
    outputs(3028) <= not(layer2_outputs(5807));
    outputs(3029) <= not(layer2_outputs(10358)) or (layer2_outputs(6895));
    outputs(3030) <= layer2_outputs(3720);
    outputs(3031) <= layer2_outputs(11648);
    outputs(3032) <= (layer2_outputs(7236)) and not (layer2_outputs(2827));
    outputs(3033) <= not(layer2_outputs(10165)) or (layer2_outputs(6094));
    outputs(3034) <= not(layer2_outputs(9450)) or (layer2_outputs(4537));
    outputs(3035) <= layer2_outputs(11090);
    outputs(3036) <= not((layer2_outputs(5452)) xor (layer2_outputs(5219)));
    outputs(3037) <= layer2_outputs(5508);
    outputs(3038) <= not(layer2_outputs(5604));
    outputs(3039) <= layer2_outputs(8377);
    outputs(3040) <= not(layer2_outputs(4420));
    outputs(3041) <= not(layer2_outputs(10489));
    outputs(3042) <= (layer2_outputs(7378)) and not (layer2_outputs(11267));
    outputs(3043) <= not(layer2_outputs(8416)) or (layer2_outputs(6680));
    outputs(3044) <= layer2_outputs(12664);
    outputs(3045) <= (layer2_outputs(5790)) and (layer2_outputs(5914));
    outputs(3046) <= layer2_outputs(9494);
    outputs(3047) <= layer2_outputs(8172);
    outputs(3048) <= layer2_outputs(11818);
    outputs(3049) <= layer2_outputs(7514);
    outputs(3050) <= not(layer2_outputs(8484));
    outputs(3051) <= not(layer2_outputs(10821));
    outputs(3052) <= not(layer2_outputs(11109));
    outputs(3053) <= layer2_outputs(4049);
    outputs(3054) <= not(layer2_outputs(10923));
    outputs(3055) <= not(layer2_outputs(9761));
    outputs(3056) <= (layer2_outputs(3640)) and not (layer2_outputs(11394));
    outputs(3057) <= layer2_outputs(10977);
    outputs(3058) <= not((layer2_outputs(9148)) xor (layer2_outputs(12299)));
    outputs(3059) <= (layer2_outputs(11367)) xor (layer2_outputs(1096));
    outputs(3060) <= not(layer2_outputs(7459));
    outputs(3061) <= layer2_outputs(703);
    outputs(3062) <= (layer2_outputs(2902)) xor (layer2_outputs(1367));
    outputs(3063) <= not((layer2_outputs(4456)) xor (layer2_outputs(10398)));
    outputs(3064) <= (layer2_outputs(378)) xor (layer2_outputs(8002));
    outputs(3065) <= layer2_outputs(457);
    outputs(3066) <= not(layer2_outputs(10600));
    outputs(3067) <= not((layer2_outputs(12296)) xor (layer2_outputs(9080)));
    outputs(3068) <= (layer2_outputs(4431)) and (layer2_outputs(9808));
    outputs(3069) <= (layer2_outputs(9035)) or (layer2_outputs(7632));
    outputs(3070) <= not(layer2_outputs(11521));
    outputs(3071) <= layer2_outputs(5812);
    outputs(3072) <= layer2_outputs(337);
    outputs(3073) <= layer2_outputs(10317);
    outputs(3074) <= not(layer2_outputs(8957));
    outputs(3075) <= (layer2_outputs(2322)) and not (layer2_outputs(8927));
    outputs(3076) <= (layer2_outputs(3319)) or (layer2_outputs(6239));
    outputs(3077) <= not(layer2_outputs(6269));
    outputs(3078) <= layer2_outputs(7388);
    outputs(3079) <= (layer2_outputs(2693)) xor (layer2_outputs(5065));
    outputs(3080) <= not(layer2_outputs(3833));
    outputs(3081) <= layer2_outputs(9977);
    outputs(3082) <= not(layer2_outputs(5811)) or (layer2_outputs(4002));
    outputs(3083) <= layer2_outputs(11370);
    outputs(3084) <= (layer2_outputs(8868)) xor (layer2_outputs(4725));
    outputs(3085) <= (layer2_outputs(5786)) xor (layer2_outputs(7705));
    outputs(3086) <= (layer2_outputs(5325)) or (layer2_outputs(7962));
    outputs(3087) <= layer2_outputs(3119);
    outputs(3088) <= not(layer2_outputs(6002));
    outputs(3089) <= not(layer2_outputs(8000));
    outputs(3090) <= layer2_outputs(5364);
    outputs(3091) <= not(layer2_outputs(3094));
    outputs(3092) <= not(layer2_outputs(6696));
    outputs(3093) <= not((layer2_outputs(3159)) and (layer2_outputs(1334)));
    outputs(3094) <= layer2_outputs(3949);
    outputs(3095) <= (layer2_outputs(2779)) and (layer2_outputs(3995));
    outputs(3096) <= not(layer2_outputs(10859));
    outputs(3097) <= not(layer2_outputs(8542));
    outputs(3098) <= not(layer2_outputs(3354));
    outputs(3099) <= layer2_outputs(2552);
    outputs(3100) <= not(layer2_outputs(3040));
    outputs(3101) <= (layer2_outputs(7575)) or (layer2_outputs(968));
    outputs(3102) <= not(layer2_outputs(11662));
    outputs(3103) <= not(layer2_outputs(6709));
    outputs(3104) <= (layer2_outputs(9762)) or (layer2_outputs(6968));
    outputs(3105) <= (layer2_outputs(7635)) or (layer2_outputs(6741));
    outputs(3106) <= (layer2_outputs(11602)) and not (layer2_outputs(1797));
    outputs(3107) <= not(layer2_outputs(7371));
    outputs(3108) <= not(layer2_outputs(3118)) or (layer2_outputs(3947));
    outputs(3109) <= not((layer2_outputs(6803)) xor (layer2_outputs(5897)));
    outputs(3110) <= layer2_outputs(1882);
    outputs(3111) <= not(layer2_outputs(1377));
    outputs(3112) <= (layer2_outputs(2708)) xor (layer2_outputs(11439));
    outputs(3113) <= not((layer2_outputs(990)) xor (layer2_outputs(6187)));
    outputs(3114) <= (layer2_outputs(2016)) or (layer2_outputs(5029));
    outputs(3115) <= (layer2_outputs(2121)) xor (layer2_outputs(2710));
    outputs(3116) <= (layer2_outputs(8604)) and not (layer2_outputs(11949));
    outputs(3117) <= layer2_outputs(5571);
    outputs(3118) <= not(layer2_outputs(11554));
    outputs(3119) <= (layer2_outputs(1412)) and not (layer2_outputs(1518));
    outputs(3120) <= layer2_outputs(8789);
    outputs(3121) <= layer2_outputs(12144);
    outputs(3122) <= not(layer2_outputs(11787));
    outputs(3123) <= not(layer2_outputs(9807));
    outputs(3124) <= not(layer2_outputs(8350));
    outputs(3125) <= not(layer2_outputs(9169));
    outputs(3126) <= not((layer2_outputs(5232)) or (layer2_outputs(9381)));
    outputs(3127) <= not(layer2_outputs(4223));
    outputs(3128) <= not(layer2_outputs(5102)) or (layer2_outputs(1701));
    outputs(3129) <= (layer2_outputs(5221)) xor (layer2_outputs(5800));
    outputs(3130) <= (layer2_outputs(582)) xor (layer2_outputs(6470));
    outputs(3131) <= not((layer2_outputs(4122)) and (layer2_outputs(2600)));
    outputs(3132) <= layer2_outputs(3955);
    outputs(3133) <= layer2_outputs(1856);
    outputs(3134) <= layer2_outputs(5844);
    outputs(3135) <= not(layer2_outputs(5494)) or (layer2_outputs(10732));
    outputs(3136) <= layer2_outputs(1655);
    outputs(3137) <= not((layer2_outputs(11821)) or (layer2_outputs(7089)));
    outputs(3138) <= layer2_outputs(2217);
    outputs(3139) <= layer2_outputs(11888);
    outputs(3140) <= not(layer2_outputs(4929));
    outputs(3141) <= layer2_outputs(4797);
    outputs(3142) <= not(layer2_outputs(8949));
    outputs(3143) <= not(layer2_outputs(2892));
    outputs(3144) <= not(layer2_outputs(11421)) or (layer2_outputs(10317));
    outputs(3145) <= not(layer2_outputs(962));
    outputs(3146) <= not(layer2_outputs(9832));
    outputs(3147) <= not((layer2_outputs(646)) xor (layer2_outputs(7611)));
    outputs(3148) <= layer2_outputs(12310);
    outputs(3149) <= layer2_outputs(1459);
    outputs(3150) <= not(layer2_outputs(3520));
    outputs(3151) <= layer2_outputs(9523);
    outputs(3152) <= (layer2_outputs(2362)) and not (layer2_outputs(5793));
    outputs(3153) <= not(layer2_outputs(1106));
    outputs(3154) <= not(layer2_outputs(9993));
    outputs(3155) <= layer2_outputs(2022);
    outputs(3156) <= (layer2_outputs(3411)) xor (layer2_outputs(12136));
    outputs(3157) <= layer2_outputs(3549);
    outputs(3158) <= layer2_outputs(9989);
    outputs(3159) <= not((layer2_outputs(2628)) and (layer2_outputs(8598)));
    outputs(3160) <= not((layer2_outputs(1341)) xor (layer2_outputs(8580)));
    outputs(3161) <= layer2_outputs(5452);
    outputs(3162) <= layer2_outputs(909);
    outputs(3163) <= layer2_outputs(7585);
    outputs(3164) <= (layer2_outputs(11473)) and (layer2_outputs(1429));
    outputs(3165) <= (layer2_outputs(5672)) and not (layer2_outputs(12039));
    outputs(3166) <= layer2_outputs(10768);
    outputs(3167) <= not(layer2_outputs(4780));
    outputs(3168) <= layer2_outputs(5654);
    outputs(3169) <= not((layer2_outputs(8328)) xor (layer2_outputs(11714)));
    outputs(3170) <= (layer2_outputs(1330)) xor (layer2_outputs(7934));
    outputs(3171) <= not(layer2_outputs(29)) or (layer2_outputs(9787));
    outputs(3172) <= (layer2_outputs(2956)) xor (layer2_outputs(6801));
    outputs(3173) <= not((layer2_outputs(802)) and (layer2_outputs(7215)));
    outputs(3174) <= not(layer2_outputs(4235));
    outputs(3175) <= layer2_outputs(5253);
    outputs(3176) <= (layer2_outputs(8139)) xor (layer2_outputs(10042));
    outputs(3177) <= not((layer2_outputs(11003)) or (layer2_outputs(370)));
    outputs(3178) <= not((layer2_outputs(3960)) xor (layer2_outputs(12708)));
    outputs(3179) <= not(layer2_outputs(10066));
    outputs(3180) <= not((layer2_outputs(9930)) and (layer2_outputs(12263)));
    outputs(3181) <= not((layer2_outputs(1526)) xor (layer2_outputs(11917)));
    outputs(3182) <= layer2_outputs(2472);
    outputs(3183) <= layer2_outputs(7375);
    outputs(3184) <= not(layer2_outputs(9241));
    outputs(3185) <= layer2_outputs(694);
    outputs(3186) <= layer2_outputs(2299);
    outputs(3187) <= not((layer2_outputs(3427)) xor (layer2_outputs(2434)));
    outputs(3188) <= not(layer2_outputs(4444));
    outputs(3189) <= not(layer2_outputs(5726)) or (layer2_outputs(11475));
    outputs(3190) <= not(layer2_outputs(4594)) or (layer2_outputs(355));
    outputs(3191) <= not((layer2_outputs(7151)) or (layer2_outputs(4867)));
    outputs(3192) <= layer2_outputs(720);
    outputs(3193) <= not(layer2_outputs(260));
    outputs(3194) <= not(layer2_outputs(7872));
    outputs(3195) <= not(layer2_outputs(8683)) or (layer2_outputs(3045));
    outputs(3196) <= not(layer2_outputs(1313));
    outputs(3197) <= layer2_outputs(10175);
    outputs(3198) <= not(layer2_outputs(5857));
    outputs(3199) <= layer2_outputs(737);
    outputs(3200) <= layer2_outputs(7261);
    outputs(3201) <= not(layer2_outputs(1921));
    outputs(3202) <= layer2_outputs(1282);
    outputs(3203) <= not(layer2_outputs(10146));
    outputs(3204) <= layer2_outputs(7882);
    outputs(3205) <= not(layer2_outputs(2261));
    outputs(3206) <= not((layer2_outputs(10134)) and (layer2_outputs(1629)));
    outputs(3207) <= not(layer2_outputs(3216));
    outputs(3208) <= not(layer2_outputs(5034));
    outputs(3209) <= layer2_outputs(2946);
    outputs(3210) <= (layer2_outputs(8314)) xor (layer2_outputs(11471));
    outputs(3211) <= (layer2_outputs(1727)) and not (layer2_outputs(8223));
    outputs(3212) <= layer2_outputs(9603);
    outputs(3213) <= not((layer2_outputs(4194)) xor (layer2_outputs(8144)));
    outputs(3214) <= not(layer2_outputs(32));
    outputs(3215) <= not((layer2_outputs(2918)) xor (layer2_outputs(1763)));
    outputs(3216) <= not(layer2_outputs(3568));
    outputs(3217) <= not(layer2_outputs(200));
    outputs(3218) <= (layer2_outputs(5924)) xor (layer2_outputs(2167));
    outputs(3219) <= layer2_outputs(10379);
    outputs(3220) <= (layer2_outputs(1484)) xor (layer2_outputs(8713));
    outputs(3221) <= not(layer2_outputs(4160)) or (layer2_outputs(11396));
    outputs(3222) <= layer2_outputs(11713);
    outputs(3223) <= (layer2_outputs(7865)) or (layer2_outputs(3148));
    outputs(3224) <= not(layer2_outputs(2248));
    outputs(3225) <= not(layer2_outputs(2443));
    outputs(3226) <= not(layer2_outputs(5828)) or (layer2_outputs(10621));
    outputs(3227) <= not((layer2_outputs(6208)) and (layer2_outputs(5005)));
    outputs(3228) <= not((layer2_outputs(6683)) xor (layer2_outputs(8431)));
    outputs(3229) <= layer2_outputs(11900);
    outputs(3230) <= (layer2_outputs(12738)) and not (layer2_outputs(1133));
    outputs(3231) <= not(layer2_outputs(95));
    outputs(3232) <= not(layer2_outputs(7647));
    outputs(3233) <= not(layer2_outputs(4365)) or (layer2_outputs(3731));
    outputs(3234) <= not(layer2_outputs(12130));
    outputs(3235) <= layer2_outputs(275);
    outputs(3236) <= not(layer2_outputs(2802));
    outputs(3237) <= layer2_outputs(2778);
    outputs(3238) <= layer2_outputs(4363);
    outputs(3239) <= layer2_outputs(7168);
    outputs(3240) <= layer2_outputs(10693);
    outputs(3241) <= not(layer2_outputs(3264)) or (layer2_outputs(3522));
    outputs(3242) <= layer2_outputs(696);
    outputs(3243) <= not(layer2_outputs(2241));
    outputs(3244) <= not((layer2_outputs(4900)) or (layer2_outputs(9774)));
    outputs(3245) <= not((layer2_outputs(3978)) xor (layer2_outputs(9676)));
    outputs(3246) <= layer2_outputs(6102);
    outputs(3247) <= not(layer2_outputs(2323));
    outputs(3248) <= (layer2_outputs(7183)) and not (layer2_outputs(11682));
    outputs(3249) <= not(layer2_outputs(1135));
    outputs(3250) <= layer2_outputs(8823);
    outputs(3251) <= layer2_outputs(10128);
    outputs(3252) <= not((layer2_outputs(4402)) and (layer2_outputs(10755)));
    outputs(3253) <= not((layer2_outputs(9301)) and (layer2_outputs(7292)));
    outputs(3254) <= not((layer2_outputs(12003)) xor (layer2_outputs(6763)));
    outputs(3255) <= not(layer2_outputs(2611)) or (layer2_outputs(10966));
    outputs(3256) <= not(layer2_outputs(831)) or (layer2_outputs(6795));
    outputs(3257) <= (layer2_outputs(4962)) xor (layer2_outputs(4108));
    outputs(3258) <= not(layer2_outputs(1421));
    outputs(3259) <= layer2_outputs(10948);
    outputs(3260) <= not((layer2_outputs(11852)) or (layer2_outputs(5880)));
    outputs(3261) <= not((layer2_outputs(7763)) and (layer2_outputs(6630)));
    outputs(3262) <= layer2_outputs(11848);
    outputs(3263) <= layer2_outputs(9564);
    outputs(3264) <= (layer2_outputs(3563)) xor (layer2_outputs(6197));
    outputs(3265) <= (layer2_outputs(3707)) or (layer2_outputs(3532));
    outputs(3266) <= not(layer2_outputs(7517)) or (layer2_outputs(140));
    outputs(3267) <= layer2_outputs(3283);
    outputs(3268) <= not(layer2_outputs(1438));
    outputs(3269) <= layer2_outputs(8399);
    outputs(3270) <= not(layer2_outputs(7866));
    outputs(3271) <= not(layer2_outputs(6688));
    outputs(3272) <= layer2_outputs(4631);
    outputs(3273) <= not(layer2_outputs(1594));
    outputs(3274) <= not(layer2_outputs(11528));
    outputs(3275) <= not(layer2_outputs(8014));
    outputs(3276) <= not((layer2_outputs(7487)) and (layer2_outputs(12164)));
    outputs(3277) <= not((layer2_outputs(11790)) or (layer2_outputs(3392)));
    outputs(3278) <= layer2_outputs(8337);
    outputs(3279) <= not((layer2_outputs(8511)) xor (layer2_outputs(8602)));
    outputs(3280) <= not((layer2_outputs(135)) xor (layer2_outputs(6475)));
    outputs(3281) <= layer2_outputs(1584);
    outputs(3282) <= layer2_outputs(1296);
    outputs(3283) <= layer2_outputs(6302);
    outputs(3284) <= not(layer2_outputs(1088));
    outputs(3285) <= (layer2_outputs(5313)) or (layer2_outputs(6054));
    outputs(3286) <= layer2_outputs(4278);
    outputs(3287) <= not(layer2_outputs(4227));
    outputs(3288) <= layer2_outputs(3538);
    outputs(3289) <= (layer2_outputs(6098)) and (layer2_outputs(484));
    outputs(3290) <= layer2_outputs(5667);
    outputs(3291) <= (layer2_outputs(9005)) xor (layer2_outputs(6757));
    outputs(3292) <= layer2_outputs(484);
    outputs(3293) <= not(layer2_outputs(6581)) or (layer2_outputs(12054));
    outputs(3294) <= not((layer2_outputs(12172)) or (layer2_outputs(856)));
    outputs(3295) <= (layer2_outputs(5559)) xor (layer2_outputs(9822));
    outputs(3296) <= not(layer2_outputs(4596));
    outputs(3297) <= not(layer2_outputs(3002));
    outputs(3298) <= not(layer2_outputs(7173));
    outputs(3299) <= not(layer2_outputs(6926));
    outputs(3300) <= layer2_outputs(2184);
    outputs(3301) <= (layer2_outputs(1873)) and not (layer2_outputs(3700));
    outputs(3302) <= not(layer2_outputs(10200));
    outputs(3303) <= not(layer2_outputs(8649));
    outputs(3304) <= not(layer2_outputs(1669));
    outputs(3305) <= not(layer2_outputs(1483));
    outputs(3306) <= (layer2_outputs(1515)) xor (layer2_outputs(7651));
    outputs(3307) <= (layer2_outputs(9296)) xor (layer2_outputs(937));
    outputs(3308) <= (layer2_outputs(4461)) xor (layer2_outputs(11926));
    outputs(3309) <= layer2_outputs(5113);
    outputs(3310) <= not((layer2_outputs(4011)) and (layer2_outputs(9646)));
    outputs(3311) <= not((layer2_outputs(298)) xor (layer2_outputs(12192)));
    outputs(3312) <= layer2_outputs(8656);
    outputs(3313) <= not(layer2_outputs(11230)) or (layer2_outputs(9631));
    outputs(3314) <= not(layer2_outputs(9914)) or (layer2_outputs(4902));
    outputs(3315) <= layer2_outputs(634);
    outputs(3316) <= layer2_outputs(9128);
    outputs(3317) <= (layer2_outputs(9207)) xor (layer2_outputs(10930));
    outputs(3318) <= not(layer2_outputs(10396)) or (layer2_outputs(2428));
    outputs(3319) <= not(layer2_outputs(2854));
    outputs(3320) <= (layer2_outputs(4502)) and not (layer2_outputs(4872));
    outputs(3321) <= not(layer2_outputs(739));
    outputs(3322) <= layer2_outputs(7019);
    outputs(3323) <= (layer2_outputs(6066)) xor (layer2_outputs(11275));
    outputs(3324) <= (layer2_outputs(11356)) and not (layer2_outputs(12487));
    outputs(3325) <= layer2_outputs(2817);
    outputs(3326) <= not(layer2_outputs(8473));
    outputs(3327) <= not(layer2_outputs(11158));
    outputs(3328) <= layer2_outputs(1459);
    outputs(3329) <= not(layer2_outputs(3431));
    outputs(3330) <= layer2_outputs(3539);
    outputs(3331) <= not((layer2_outputs(487)) and (layer2_outputs(6247)));
    outputs(3332) <= (layer2_outputs(9456)) xor (layer2_outputs(3769));
    outputs(3333) <= layer2_outputs(3230);
    outputs(3334) <= not((layer2_outputs(1743)) xor (layer2_outputs(3205)));
    outputs(3335) <= not(layer2_outputs(11745));
    outputs(3336) <= layer2_outputs(2150);
    outputs(3337) <= layer2_outputs(7625);
    outputs(3338) <= not(layer2_outputs(6286)) or (layer2_outputs(5177));
    outputs(3339) <= not(layer2_outputs(1982));
    outputs(3340) <= not(layer2_outputs(5151)) or (layer2_outputs(2476));
    outputs(3341) <= layer2_outputs(420);
    outputs(3342) <= not((layer2_outputs(193)) xor (layer2_outputs(5556)));
    outputs(3343) <= layer2_outputs(4099);
    outputs(3344) <= not(layer2_outputs(8523));
    outputs(3345) <= not(layer2_outputs(9897));
    outputs(3346) <= layer2_outputs(903);
    outputs(3347) <= not((layer2_outputs(4802)) or (layer2_outputs(2926)));
    outputs(3348) <= not((layer2_outputs(1173)) xor (layer2_outputs(6533)));
    outputs(3349) <= not(layer2_outputs(10777));
    outputs(3350) <= (layer2_outputs(7389)) xor (layer2_outputs(5758));
    outputs(3351) <= layer2_outputs(2272);
    outputs(3352) <= (layer2_outputs(2252)) xor (layer2_outputs(4396));
    outputs(3353) <= layer2_outputs(11304);
    outputs(3354) <= not((layer2_outputs(3979)) xor (layer2_outputs(8654)));
    outputs(3355) <= not(layer2_outputs(11508));
    outputs(3356) <= layer2_outputs(4183);
    outputs(3357) <= not(layer2_outputs(7765));
    outputs(3358) <= not(layer2_outputs(7006)) or (layer2_outputs(2480));
    outputs(3359) <= (layer2_outputs(5465)) and not (layer2_outputs(2657));
    outputs(3360) <= not((layer2_outputs(795)) and (layer2_outputs(11452)));
    outputs(3361) <= layer2_outputs(4983);
    outputs(3362) <= not(layer2_outputs(11109));
    outputs(3363) <= layer2_outputs(6057);
    outputs(3364) <= not(layer2_outputs(8130));
    outputs(3365) <= not(layer2_outputs(9912)) or (layer2_outputs(7136));
    outputs(3366) <= layer2_outputs(3876);
    outputs(3367) <= (layer2_outputs(11056)) xor (layer2_outputs(5322));
    outputs(3368) <= (layer2_outputs(1516)) and (layer2_outputs(3027));
    outputs(3369) <= not(layer2_outputs(3894));
    outputs(3370) <= not(layer2_outputs(6615));
    outputs(3371) <= layer2_outputs(7416);
    outputs(3372) <= layer2_outputs(11901);
    outputs(3373) <= layer2_outputs(5919);
    outputs(3374) <= layer2_outputs(9003);
    outputs(3375) <= layer2_outputs(3881);
    outputs(3376) <= (layer2_outputs(5936)) xor (layer2_outputs(445));
    outputs(3377) <= not((layer2_outputs(9840)) xor (layer2_outputs(1343)));
    outputs(3378) <= layer2_outputs(10542);
    outputs(3379) <= not(layer2_outputs(310));
    outputs(3380) <= (layer2_outputs(4302)) xor (layer2_outputs(3307));
    outputs(3381) <= not((layer2_outputs(7267)) and (layer2_outputs(9539)));
    outputs(3382) <= layer2_outputs(5606);
    outputs(3383) <= not((layer2_outputs(12634)) or (layer2_outputs(4682)));
    outputs(3384) <= not(layer2_outputs(2695)) or (layer2_outputs(4498));
    outputs(3385) <= layer2_outputs(8204);
    outputs(3386) <= not((layer2_outputs(6936)) xor (layer2_outputs(2333)));
    outputs(3387) <= (layer2_outputs(12641)) and not (layer2_outputs(2989));
    outputs(3388) <= layer2_outputs(4966);
    outputs(3389) <= not(layer2_outputs(4539));
    outputs(3390) <= not((layer2_outputs(3334)) xor (layer2_outputs(6149)));
    outputs(3391) <= not(layer2_outputs(8944)) or (layer2_outputs(3745));
    outputs(3392) <= (layer2_outputs(4233)) xor (layer2_outputs(9256));
    outputs(3393) <= (layer2_outputs(5044)) and not (layer2_outputs(7550));
    outputs(3394) <= layer2_outputs(10673);
    outputs(3395) <= layer2_outputs(12730);
    outputs(3396) <= not(layer2_outputs(5263));
    outputs(3397) <= not(layer2_outputs(4353)) or (layer2_outputs(2986));
    outputs(3398) <= layer2_outputs(4483);
    outputs(3399) <= layer2_outputs(1358);
    outputs(3400) <= (layer2_outputs(2119)) xor (layer2_outputs(6717));
    outputs(3401) <= not(layer2_outputs(10056));
    outputs(3402) <= not(layer2_outputs(2695));
    outputs(3403) <= not(layer2_outputs(1054));
    outputs(3404) <= not(layer2_outputs(8772));
    outputs(3405) <= not(layer2_outputs(7744));
    outputs(3406) <= (layer2_outputs(7072)) and (layer2_outputs(9707));
    outputs(3407) <= layer2_outputs(9488);
    outputs(3408) <= not(layer2_outputs(2535));
    outputs(3409) <= (layer2_outputs(9707)) and not (layer2_outputs(11444));
    outputs(3410) <= not(layer2_outputs(10424));
    outputs(3411) <= not(layer2_outputs(6216));
    outputs(3412) <= not(layer2_outputs(1331));
    outputs(3413) <= not(layer2_outputs(5008)) or (layer2_outputs(9472));
    outputs(3414) <= layer2_outputs(10295);
    outputs(3415) <= not(layer2_outputs(659));
    outputs(3416) <= (layer2_outputs(8681)) xor (layer2_outputs(10136));
    outputs(3417) <= layer2_outputs(4338);
    outputs(3418) <= (layer2_outputs(7051)) xor (layer2_outputs(11709));
    outputs(3419) <= not(layer2_outputs(6627));
    outputs(3420) <= (layer2_outputs(1546)) xor (layer2_outputs(2937));
    outputs(3421) <= layer2_outputs(4454);
    outputs(3422) <= layer2_outputs(4345);
    outputs(3423) <= not(layer2_outputs(7590));
    outputs(3424) <= layer2_outputs(4416);
    outputs(3425) <= not(layer2_outputs(4276));
    outputs(3426) <= (layer2_outputs(6451)) or (layer2_outputs(3810));
    outputs(3427) <= not(layer2_outputs(5721)) or (layer2_outputs(8047));
    outputs(3428) <= not((layer2_outputs(11712)) xor (layer2_outputs(5422)));
    outputs(3429) <= not(layer2_outputs(7368));
    outputs(3430) <= (layer2_outputs(1609)) xor (layer2_outputs(7393));
    outputs(3431) <= layer2_outputs(6545);
    outputs(3432) <= layer2_outputs(7084);
    outputs(3433) <= not(layer2_outputs(820));
    outputs(3434) <= not((layer2_outputs(11169)) and (layer2_outputs(12337)));
    outputs(3435) <= not(layer2_outputs(392));
    outputs(3436) <= not(layer2_outputs(5407));
    outputs(3437) <= not((layer2_outputs(11245)) xor (layer2_outputs(7434)));
    outputs(3438) <= (layer2_outputs(3674)) xor (layer2_outputs(8014));
    outputs(3439) <= (layer2_outputs(130)) xor (layer2_outputs(9756));
    outputs(3440) <= not(layer2_outputs(8145));
    outputs(3441) <= layer2_outputs(11234);
    outputs(3442) <= layer2_outputs(10731);
    outputs(3443) <= not(layer2_outputs(6409));
    outputs(3444) <= not(layer2_outputs(1717));
    outputs(3445) <= not(layer2_outputs(5306)) or (layer2_outputs(12381));
    outputs(3446) <= layer2_outputs(1419);
    outputs(3447) <= (layer2_outputs(2691)) xor (layer2_outputs(7915));
    outputs(3448) <= not(layer2_outputs(10515)) or (layer2_outputs(12712));
    outputs(3449) <= (layer2_outputs(5501)) or (layer2_outputs(3792));
    outputs(3450) <= not(layer2_outputs(10159));
    outputs(3451) <= not(layer2_outputs(11479));
    outputs(3452) <= not(layer2_outputs(7301));
    outputs(3453) <= (layer2_outputs(2842)) xor (layer2_outputs(6610));
    outputs(3454) <= layer2_outputs(9224);
    outputs(3455) <= not(layer2_outputs(8412));
    outputs(3456) <= (layer2_outputs(11565)) xor (layer2_outputs(7552));
    outputs(3457) <= layer2_outputs(8612);
    outputs(3458) <= layer2_outputs(6942);
    outputs(3459) <= not(layer2_outputs(3569));
    outputs(3460) <= not((layer2_outputs(11459)) xor (layer2_outputs(6314)));
    outputs(3461) <= not(layer2_outputs(11761));
    outputs(3462) <= (layer2_outputs(11368)) xor (layer2_outputs(8139));
    outputs(3463) <= layer2_outputs(6273);
    outputs(3464) <= (layer2_outputs(8166)) and not (layer2_outputs(8637));
    outputs(3465) <= layer2_outputs(2580);
    outputs(3466) <= not(layer2_outputs(63));
    outputs(3467) <= layer2_outputs(4806);
    outputs(3468) <= not((layer2_outputs(10680)) or (layer2_outputs(860)));
    outputs(3469) <= layer2_outputs(5035);
    outputs(3470) <= not(layer2_outputs(10593)) or (layer2_outputs(9048));
    outputs(3471) <= not(layer2_outputs(6333));
    outputs(3472) <= not(layer2_outputs(10891));
    outputs(3473) <= not((layer2_outputs(8787)) and (layer2_outputs(8099)));
    outputs(3474) <= not(layer2_outputs(6311));
    outputs(3475) <= not(layer2_outputs(5701));
    outputs(3476) <= layer2_outputs(3088);
    outputs(3477) <= (layer2_outputs(5791)) xor (layer2_outputs(9555));
    outputs(3478) <= layer2_outputs(9721);
    outputs(3479) <= (layer2_outputs(7430)) and not (layer2_outputs(3197));
    outputs(3480) <= not((layer2_outputs(3453)) or (layer2_outputs(9285)));
    outputs(3481) <= not(layer2_outputs(12269)) or (layer2_outputs(1723));
    outputs(3482) <= not(layer2_outputs(4087));
    outputs(3483) <= not((layer2_outputs(8208)) and (layer2_outputs(11586)));
    outputs(3484) <= layer2_outputs(585);
    outputs(3485) <= not(layer2_outputs(4840));
    outputs(3486) <= (layer2_outputs(587)) and (layer2_outputs(4924));
    outputs(3487) <= not((layer2_outputs(8131)) xor (layer2_outputs(11423)));
    outputs(3488) <= layer2_outputs(9320);
    outputs(3489) <= not(layer2_outputs(12748));
    outputs(3490) <= layer2_outputs(9144);
    outputs(3491) <= not(layer2_outputs(12578)) or (layer2_outputs(10170));
    outputs(3492) <= layer2_outputs(10754);
    outputs(3493) <= not(layer2_outputs(9457));
    outputs(3494) <= (layer2_outputs(11224)) or (layer2_outputs(5422));
    outputs(3495) <= layer2_outputs(9321);
    outputs(3496) <= not((layer2_outputs(4975)) xor (layer2_outputs(10445)));
    outputs(3497) <= not((layer2_outputs(7648)) and (layer2_outputs(369)));
    outputs(3498) <= layer2_outputs(1671);
    outputs(3499) <= not(layer2_outputs(6632));
    outputs(3500) <= not(layer2_outputs(7610));
    outputs(3501) <= layer2_outputs(4742);
    outputs(3502) <= layer2_outputs(4163);
    outputs(3503) <= not(layer2_outputs(12774)) or (layer2_outputs(9090));
    outputs(3504) <= (layer2_outputs(6263)) xor (layer2_outputs(10533));
    outputs(3505) <= layer2_outputs(1635);
    outputs(3506) <= layer2_outputs(8001);
    outputs(3507) <= (layer2_outputs(12256)) xor (layer2_outputs(4249));
    outputs(3508) <= not(layer2_outputs(5706));
    outputs(3509) <= layer2_outputs(1346);
    outputs(3510) <= (layer2_outputs(8366)) xor (layer2_outputs(33));
    outputs(3511) <= (layer2_outputs(10508)) and not (layer2_outputs(221));
    outputs(3512) <= not(layer2_outputs(2138));
    outputs(3513) <= not(layer2_outputs(1575));
    outputs(3514) <= not((layer2_outputs(2894)) xor (layer2_outputs(5215)));
    outputs(3515) <= layer2_outputs(8191);
    outputs(3516) <= layer2_outputs(12637);
    outputs(3517) <= (layer2_outputs(8875)) or (layer2_outputs(4065));
    outputs(3518) <= (layer2_outputs(6323)) and not (layer2_outputs(7313));
    outputs(3519) <= layer2_outputs(1777);
    outputs(3520) <= not((layer2_outputs(1259)) xor (layer2_outputs(4898)));
    outputs(3521) <= (layer2_outputs(10689)) and not (layer2_outputs(2656));
    outputs(3522) <= not((layer2_outputs(219)) and (layer2_outputs(100)));
    outputs(3523) <= not((layer2_outputs(556)) xor (layer2_outputs(5558)));
    outputs(3524) <= layer2_outputs(2622);
    outputs(3525) <= not((layer2_outputs(603)) xor (layer2_outputs(4812)));
    outputs(3526) <= not(layer2_outputs(11425));
    outputs(3527) <= (layer2_outputs(8079)) xor (layer2_outputs(1325));
    outputs(3528) <= layer2_outputs(8167);
    outputs(3529) <= (layer2_outputs(3655)) or (layer2_outputs(4952));
    outputs(3530) <= not(layer2_outputs(12298));
    outputs(3531) <= layer2_outputs(8876);
    outputs(3532) <= not(layer2_outputs(6345));
    outputs(3533) <= layer2_outputs(7852);
    outputs(3534) <= layer2_outputs(11652);
    outputs(3535) <= not(layer2_outputs(6661));
    outputs(3536) <= layer2_outputs(11296);
    outputs(3537) <= not((layer2_outputs(4818)) and (layer2_outputs(2885)));
    outputs(3538) <= layer2_outputs(610);
    outputs(3539) <= not(layer2_outputs(11029));
    outputs(3540) <= not(layer2_outputs(2463));
    outputs(3541) <= layer2_outputs(8309);
    outputs(3542) <= layer2_outputs(4623);
    outputs(3543) <= (layer2_outputs(9790)) and not (layer2_outputs(6163));
    outputs(3544) <= (layer2_outputs(2934)) xor (layer2_outputs(1369));
    outputs(3545) <= not((layer2_outputs(4934)) and (layer2_outputs(12400)));
    outputs(3546) <= not(layer2_outputs(2233));
    outputs(3547) <= (layer2_outputs(10429)) xor (layer2_outputs(12012));
    outputs(3548) <= not(layer2_outputs(7160));
    outputs(3549) <= (layer2_outputs(10316)) or (layer2_outputs(10153));
    outputs(3550) <= (layer2_outputs(5207)) xor (layer2_outputs(3859));
    outputs(3551) <= (layer2_outputs(5023)) or (layer2_outputs(5753));
    outputs(3552) <= layer2_outputs(11731);
    outputs(3553) <= (layer2_outputs(2316)) xor (layer2_outputs(11926));
    outputs(3554) <= (layer2_outputs(5074)) xor (layer2_outputs(46));
    outputs(3555) <= layer2_outputs(8718);
    outputs(3556) <= not(layer2_outputs(6526));
    outputs(3557) <= not((layer2_outputs(5433)) and (layer2_outputs(911)));
    outputs(3558) <= (layer2_outputs(5397)) and (layer2_outputs(4019));
    outputs(3559) <= not((layer2_outputs(6237)) xor (layer2_outputs(9878)));
    outputs(3560) <= (layer2_outputs(2700)) and (layer2_outputs(8687));
    outputs(3561) <= not(layer2_outputs(4207));
    outputs(3562) <= layer2_outputs(4830);
    outputs(3563) <= not(layer2_outputs(1674));
    outputs(3564) <= layer2_outputs(3667);
    outputs(3565) <= layer2_outputs(8525);
    outputs(3566) <= not(layer2_outputs(11948));
    outputs(3567) <= (layer2_outputs(918)) xor (layer2_outputs(12567));
    outputs(3568) <= layer2_outputs(8541);
    outputs(3569) <= (layer2_outputs(4358)) xor (layer2_outputs(11877));
    outputs(3570) <= layer2_outputs(12183);
    outputs(3571) <= layer2_outputs(10970);
    outputs(3572) <= not(layer2_outputs(4153));
    outputs(3573) <= not(layer2_outputs(615));
    outputs(3574) <= not(layer2_outputs(11150)) or (layer2_outputs(1971));
    outputs(3575) <= layer2_outputs(11346);
    outputs(3576) <= (layer2_outputs(5555)) and (layer2_outputs(7036));
    outputs(3577) <= not(layer2_outputs(7896));
    outputs(3578) <= layer2_outputs(11547);
    outputs(3579) <= not(layer2_outputs(6906));
    outputs(3580) <= (layer2_outputs(8126)) and not (layer2_outputs(665));
    outputs(3581) <= layer2_outputs(8086);
    outputs(3582) <= not(layer2_outputs(6522));
    outputs(3583) <= layer2_outputs(1328);
    outputs(3584) <= layer2_outputs(10553);
    outputs(3585) <= not((layer2_outputs(4593)) xor (layer2_outputs(7120)));
    outputs(3586) <= (layer2_outputs(2796)) xor (layer2_outputs(7669));
    outputs(3587) <= not(layer2_outputs(1703));
    outputs(3588) <= not(layer2_outputs(10009));
    outputs(3589) <= layer2_outputs(11137);
    outputs(3590) <= (layer2_outputs(9813)) xor (layer2_outputs(12720));
    outputs(3591) <= not(layer2_outputs(11209));
    outputs(3592) <= not(layer2_outputs(2713)) or (layer2_outputs(4530));
    outputs(3593) <= (layer2_outputs(10120)) or (layer2_outputs(7514));
    outputs(3594) <= layer2_outputs(2890);
    outputs(3595) <= (layer2_outputs(11476)) xor (layer2_outputs(2302));
    outputs(3596) <= (layer2_outputs(1733)) xor (layer2_outputs(567));
    outputs(3597) <= layer2_outputs(8823);
    outputs(3598) <= not((layer2_outputs(5525)) and (layer2_outputs(3980)));
    outputs(3599) <= layer2_outputs(5395);
    outputs(3600) <= not((layer2_outputs(12548)) or (layer2_outputs(9484)));
    outputs(3601) <= layer2_outputs(11235);
    outputs(3602) <= layer2_outputs(6246);
    outputs(3603) <= (layer2_outputs(3198)) and (layer2_outputs(4814));
    outputs(3604) <= not(layer2_outputs(11091));
    outputs(3605) <= (layer2_outputs(594)) xor (layer2_outputs(9726));
    outputs(3606) <= (layer2_outputs(9470)) xor (layer2_outputs(5188));
    outputs(3607) <= layer2_outputs(6123);
    outputs(3608) <= layer2_outputs(11277);
    outputs(3609) <= (layer2_outputs(6392)) xor (layer2_outputs(10522));
    outputs(3610) <= not(layer2_outputs(2396));
    outputs(3611) <= not(layer2_outputs(9307));
    outputs(3612) <= not(layer2_outputs(2016));
    outputs(3613) <= not((layer2_outputs(3866)) and (layer2_outputs(7771)));
    outputs(3614) <= (layer2_outputs(11893)) xor (layer2_outputs(4571));
    outputs(3615) <= (layer2_outputs(5034)) xor (layer2_outputs(8836));
    outputs(3616) <= (layer2_outputs(2021)) or (layer2_outputs(6606));
    outputs(3617) <= not(layer2_outputs(11397));
    outputs(3618) <= layer2_outputs(1232);
    outputs(3619) <= layer2_outputs(10031);
    outputs(3620) <= layer2_outputs(2483);
    outputs(3621) <= (layer2_outputs(10657)) xor (layer2_outputs(4218));
    outputs(3622) <= (layer2_outputs(11007)) and not (layer2_outputs(11280));
    outputs(3623) <= not(layer2_outputs(6889));
    outputs(3624) <= (layer2_outputs(11084)) xor (layer2_outputs(4072));
    outputs(3625) <= layer2_outputs(12643);
    outputs(3626) <= (layer2_outputs(11376)) xor (layer2_outputs(932));
    outputs(3627) <= layer2_outputs(7473);
    outputs(3628) <= layer2_outputs(5657);
    outputs(3629) <= (layer2_outputs(6365)) and not (layer2_outputs(4331));
    outputs(3630) <= not(layer2_outputs(1518));
    outputs(3631) <= not(layer2_outputs(9254));
    outputs(3632) <= not(layer2_outputs(2108));
    outputs(3633) <= not(layer2_outputs(5431));
    outputs(3634) <= not((layer2_outputs(10675)) and (layer2_outputs(2967)));
    outputs(3635) <= layer2_outputs(10609);
    outputs(3636) <= not((layer2_outputs(6953)) xor (layer2_outputs(2359)));
    outputs(3637) <= not(layer2_outputs(8393));
    outputs(3638) <= not(layer2_outputs(7529)) or (layer2_outputs(2719));
    outputs(3639) <= not(layer2_outputs(9955)) or (layer2_outputs(6112));
    outputs(3640) <= layer2_outputs(12769);
    outputs(3641) <= (layer2_outputs(11255)) or (layer2_outputs(7506));
    outputs(3642) <= (layer2_outputs(10476)) xor (layer2_outputs(11716));
    outputs(3643) <= (layer2_outputs(803)) and (layer2_outputs(12064));
    outputs(3644) <= not((layer2_outputs(9333)) and (layer2_outputs(10232)));
    outputs(3645) <= not(layer2_outputs(3936));
    outputs(3646) <= (layer2_outputs(3283)) or (layer2_outputs(1142));
    outputs(3647) <= not(layer2_outputs(8548));
    outputs(3648) <= layer2_outputs(9295);
    outputs(3649) <= layer2_outputs(287);
    outputs(3650) <= not((layer2_outputs(11343)) xor (layer2_outputs(7801)));
    outputs(3651) <= (layer2_outputs(3778)) and (layer2_outputs(7325));
    outputs(3652) <= layer2_outputs(11600);
    outputs(3653) <= not(layer2_outputs(7719));
    outputs(3654) <= not(layer2_outputs(7944));
    outputs(3655) <= (layer2_outputs(9910)) xor (layer2_outputs(7460));
    outputs(3656) <= not((layer2_outputs(7954)) xor (layer2_outputs(3365)));
    outputs(3657) <= layer2_outputs(9444);
    outputs(3658) <= not(layer2_outputs(10182));
    outputs(3659) <= (layer2_outputs(8392)) xor (layer2_outputs(3724));
    outputs(3660) <= not(layer2_outputs(597));
    outputs(3661) <= not(layer2_outputs(6725)) or (layer2_outputs(5922));
    outputs(3662) <= not(layer2_outputs(6448));
    outputs(3663) <= not(layer2_outputs(4539));
    outputs(3664) <= not(layer2_outputs(2742));
    outputs(3665) <= layer2_outputs(3719);
    outputs(3666) <= not(layer2_outputs(3332));
    outputs(3667) <= layer2_outputs(7320);
    outputs(3668) <= layer2_outputs(4440);
    outputs(3669) <= not(layer2_outputs(920)) or (layer2_outputs(11447));
    outputs(3670) <= (layer2_outputs(12125)) xor (layer2_outputs(7911));
    outputs(3671) <= not(layer2_outputs(621));
    outputs(3672) <= (layer2_outputs(2188)) and (layer2_outputs(1362));
    outputs(3673) <= layer2_outputs(10718);
    outputs(3674) <= not(layer2_outputs(12745));
    outputs(3675) <= layer2_outputs(883);
    outputs(3676) <= not(layer2_outputs(786)) or (layer2_outputs(7635));
    outputs(3677) <= not(layer2_outputs(612));
    outputs(3678) <= (layer2_outputs(1165)) xor (layer2_outputs(8063));
    outputs(3679) <= not(layer2_outputs(6835));
    outputs(3680) <= layer2_outputs(9651);
    outputs(3681) <= (layer2_outputs(9288)) xor (layer2_outputs(7296));
    outputs(3682) <= layer2_outputs(2673);
    outputs(3683) <= layer2_outputs(9536);
    outputs(3684) <= layer2_outputs(1766);
    outputs(3685) <= (layer2_outputs(4987)) and not (layer2_outputs(955));
    outputs(3686) <= (layer2_outputs(12722)) xor (layer2_outputs(5972));
    outputs(3687) <= not(layer2_outputs(11023));
    outputs(3688) <= layer2_outputs(4056);
    outputs(3689) <= not(layer2_outputs(12380)) or (layer2_outputs(780));
    outputs(3690) <= layer2_outputs(3210);
    outputs(3691) <= not(layer2_outputs(7087)) or (layer2_outputs(10965));
    outputs(3692) <= (layer2_outputs(4592)) and not (layer2_outputs(2595));
    outputs(3693) <= not(layer2_outputs(8248));
    outputs(3694) <= layer2_outputs(2872);
    outputs(3695) <= (layer2_outputs(1278)) and (layer2_outputs(11807));
    outputs(3696) <= (layer2_outputs(2807)) xor (layer2_outputs(6299));
    outputs(3697) <= not((layer2_outputs(1531)) and (layer2_outputs(1444)));
    outputs(3698) <= layer2_outputs(6798);
    outputs(3699) <= (layer2_outputs(9087)) xor (layer2_outputs(3292));
    outputs(3700) <= not(layer2_outputs(3537));
    outputs(3701) <= not(layer2_outputs(5110));
    outputs(3702) <= layer2_outputs(11144);
    outputs(3703) <= (layer2_outputs(8630)) or (layer2_outputs(3091));
    outputs(3704) <= not((layer2_outputs(5076)) xor (layer2_outputs(3772)));
    outputs(3705) <= not(layer2_outputs(3869));
    outputs(3706) <= layer2_outputs(4220);
    outputs(3707) <= (layer2_outputs(967)) xor (layer2_outputs(2036));
    outputs(3708) <= not(layer2_outputs(3553));
    outputs(3709) <= layer2_outputs(2919);
    outputs(3710) <= (layer2_outputs(4969)) xor (layer2_outputs(5237));
    outputs(3711) <= layer2_outputs(4341);
    outputs(3712) <= not((layer2_outputs(9394)) xor (layer2_outputs(3919)));
    outputs(3713) <= not(layer2_outputs(9666));
    outputs(3714) <= layer2_outputs(11188);
    outputs(3715) <= layer2_outputs(10571);
    outputs(3716) <= layer2_outputs(9977);
    outputs(3717) <= layer2_outputs(2352);
    outputs(3718) <= layer2_outputs(9268);
    outputs(3719) <= not(layer2_outputs(7344));
    outputs(3720) <= not((layer2_outputs(2029)) xor (layer2_outputs(5522)));
    outputs(3721) <= layer2_outputs(1713);
    outputs(3722) <= not(layer2_outputs(7598));
    outputs(3723) <= (layer2_outputs(5692)) xor (layer2_outputs(3762));
    outputs(3724) <= (layer2_outputs(2134)) or (layer2_outputs(5961));
    outputs(3725) <= not(layer2_outputs(11913));
    outputs(3726) <= not((layer2_outputs(2430)) and (layer2_outputs(4528)));
    outputs(3727) <= not(layer2_outputs(4776));
    outputs(3728) <= (layer2_outputs(4547)) xor (layer2_outputs(3513));
    outputs(3729) <= (layer2_outputs(1648)) or (layer2_outputs(8023));
    outputs(3730) <= layer2_outputs(959);
    outputs(3731) <= layer2_outputs(11776);
    outputs(3732) <= layer2_outputs(4971);
    outputs(3733) <= (layer2_outputs(7136)) and not (layer2_outputs(9040));
    outputs(3734) <= not(layer2_outputs(12458));
    outputs(3735) <= not(layer2_outputs(8773));
    outputs(3736) <= layer2_outputs(6487);
    outputs(3737) <= layer2_outputs(2971);
    outputs(3738) <= not((layer2_outputs(10665)) xor (layer2_outputs(7043)));
    outputs(3739) <= (layer2_outputs(2263)) and not (layer2_outputs(2265));
    outputs(3740) <= (layer2_outputs(6974)) xor (layer2_outputs(6794));
    outputs(3741) <= not(layer2_outputs(10011));
    outputs(3742) <= layer2_outputs(4876);
    outputs(3743) <= not(layer2_outputs(4584));
    outputs(3744) <= (layer2_outputs(7197)) xor (layer2_outputs(7030));
    outputs(3745) <= not(layer2_outputs(9794));
    outputs(3746) <= layer2_outputs(5472);
    outputs(3747) <= not(layer2_outputs(11705));
    outputs(3748) <= not(layer2_outputs(9482));
    outputs(3749) <= layer2_outputs(6672);
    outputs(3750) <= not(layer2_outputs(6623));
    outputs(3751) <= (layer2_outputs(9974)) xor (layer2_outputs(10682));
    outputs(3752) <= not(layer2_outputs(8405));
    outputs(3753) <= not((layer2_outputs(7609)) xor (layer2_outputs(1294)));
    outputs(3754) <= (layer2_outputs(11626)) xor (layer2_outputs(3401));
    outputs(3755) <= not(layer2_outputs(987));
    outputs(3756) <= not((layer2_outputs(3679)) or (layer2_outputs(1513)));
    outputs(3757) <= not(layer2_outputs(9825));
    outputs(3758) <= layer2_outputs(9722);
    outputs(3759) <= not(layer2_outputs(11814)) or (layer2_outputs(12059));
    outputs(3760) <= not((layer2_outputs(2896)) xor (layer2_outputs(10496)));
    outputs(3761) <= layer2_outputs(7519);
    outputs(3762) <= layer2_outputs(12356);
    outputs(3763) <= layer2_outputs(2569);
    outputs(3764) <= not((layer2_outputs(295)) xor (layer2_outputs(1808)));
    outputs(3765) <= not(layer2_outputs(11461));
    outputs(3766) <= not(layer2_outputs(7469)) or (layer2_outputs(774));
    outputs(3767) <= not(layer2_outputs(5923));
    outputs(3768) <= not(layer2_outputs(5795));
    outputs(3769) <= not((layer2_outputs(3023)) xor (layer2_outputs(12584)));
    outputs(3770) <= layer2_outputs(12651);
    outputs(3771) <= (layer2_outputs(1484)) xor (layer2_outputs(6867));
    outputs(3772) <= not((layer2_outputs(9670)) xor (layer2_outputs(11222)));
    outputs(3773) <= not((layer2_outputs(12000)) and (layer2_outputs(4030)));
    outputs(3774) <= layer2_outputs(12279);
    outputs(3775) <= (layer2_outputs(1884)) xor (layer2_outputs(11180));
    outputs(3776) <= layer2_outputs(8466);
    outputs(3777) <= layer2_outputs(8212);
    outputs(3778) <= not(layer2_outputs(4479));
    outputs(3779) <= not(layer2_outputs(3872));
    outputs(3780) <= layer2_outputs(7276);
    outputs(3781) <= not(layer2_outputs(2755));
    outputs(3782) <= layer2_outputs(11096);
    outputs(3783) <= layer2_outputs(4655);
    outputs(3784) <= not(layer2_outputs(12181)) or (layer2_outputs(5754));
    outputs(3785) <= not((layer2_outputs(11156)) xor (layer2_outputs(2306)));
    outputs(3786) <= not(layer2_outputs(4426));
    outputs(3787) <= not(layer2_outputs(4432));
    outputs(3788) <= not(layer2_outputs(1573));
    outputs(3789) <= not(layer2_outputs(4161));
    outputs(3790) <= not(layer2_outputs(7229)) or (layer2_outputs(1666));
    outputs(3791) <= (layer2_outputs(9543)) and not (layer2_outputs(6398));
    outputs(3792) <= not(layer2_outputs(1263));
    outputs(3793) <= layer2_outputs(505);
    outputs(3794) <= (layer2_outputs(2644)) and not (layer2_outputs(5071));
    outputs(3795) <= not(layer2_outputs(11202));
    outputs(3796) <= layer2_outputs(2163);
    outputs(3797) <= not(layer2_outputs(2865));
    outputs(3798) <= (layer2_outputs(3208)) xor (layer2_outputs(10694));
    outputs(3799) <= (layer2_outputs(8337)) and not (layer2_outputs(6932));
    outputs(3800) <= layer2_outputs(2763);
    outputs(3801) <= not((layer2_outputs(2234)) xor (layer2_outputs(10421)));
    outputs(3802) <= layer2_outputs(5928);
    outputs(3803) <= not((layer2_outputs(3087)) xor (layer2_outputs(4572)));
    outputs(3804) <= not(layer2_outputs(486)) or (layer2_outputs(12259));
    outputs(3805) <= not((layer2_outputs(3815)) xor (layer2_outputs(12473)));
    outputs(3806) <= not(layer2_outputs(3786));
    outputs(3807) <= not(layer2_outputs(3104));
    outputs(3808) <= not((layer2_outputs(6821)) xor (layer2_outputs(8170)));
    outputs(3809) <= not(layer2_outputs(9286));
    outputs(3810) <= (layer2_outputs(7166)) xor (layer2_outputs(7038));
    outputs(3811) <= not(layer2_outputs(5040)) or (layer2_outputs(10964));
    outputs(3812) <= not(layer2_outputs(9469));
    outputs(3813) <= layer2_outputs(3670);
    outputs(3814) <= layer2_outputs(10063);
    outputs(3815) <= not(layer2_outputs(10887)) or (layer2_outputs(4412));
    outputs(3816) <= not((layer2_outputs(2212)) xor (layer2_outputs(8251)));
    outputs(3817) <= not((layer2_outputs(5077)) xor (layer2_outputs(249)));
    outputs(3818) <= not(layer2_outputs(5829)) or (layer2_outputs(8650));
    outputs(3819) <= not(layer2_outputs(7008));
    outputs(3820) <= not((layer2_outputs(10277)) and (layer2_outputs(3362)));
    outputs(3821) <= not(layer2_outputs(6318));
    outputs(3822) <= not(layer2_outputs(8148));
    outputs(3823) <= layer2_outputs(48);
    outputs(3824) <= (layer2_outputs(4859)) xor (layer2_outputs(2195));
    outputs(3825) <= not(layer2_outputs(4443));
    outputs(3826) <= not(layer2_outputs(12036));
    outputs(3827) <= (layer2_outputs(2080)) xor (layer2_outputs(8050));
    outputs(3828) <= not(layer2_outputs(4529));
    outputs(3829) <= (layer2_outputs(5341)) xor (layer2_outputs(1109));
    outputs(3830) <= not(layer2_outputs(943));
    outputs(3831) <= layer2_outputs(1782);
    outputs(3832) <= not(layer2_outputs(10737)) or (layer2_outputs(3047));
    outputs(3833) <= not(layer2_outputs(7132));
    outputs(3834) <= (layer2_outputs(3068)) or (layer2_outputs(411));
    outputs(3835) <= layer2_outputs(7958);
    outputs(3836) <= not(layer2_outputs(6593)) or (layer2_outputs(9554));
    outputs(3837) <= not(layer2_outputs(7996));
    outputs(3838) <= layer2_outputs(2242);
    outputs(3839) <= not(layer2_outputs(12313));
    outputs(3840) <= (layer2_outputs(5056)) and (layer2_outputs(618));
    outputs(3841) <= not(layer2_outputs(12313));
    outputs(3842) <= layer2_outputs(4737);
    outputs(3843) <= layer2_outputs(4175);
    outputs(3844) <= not((layer2_outputs(5984)) and (layer2_outputs(12703)));
    outputs(3845) <= layer2_outputs(12194);
    outputs(3846) <= not((layer2_outputs(8315)) xor (layer2_outputs(6397)));
    outputs(3847) <= not((layer2_outputs(3893)) xor (layer2_outputs(3853)));
    outputs(3848) <= (layer2_outputs(3145)) xor (layer2_outputs(10092));
    outputs(3849) <= not((layer2_outputs(4687)) xor (layer2_outputs(7932)));
    outputs(3850) <= layer2_outputs(7080);
    outputs(3851) <= not(layer2_outputs(6201));
    outputs(3852) <= layer2_outputs(2057);
    outputs(3853) <= not(layer2_outputs(11895));
    outputs(3854) <= not((layer2_outputs(9174)) xor (layer2_outputs(6041)));
    outputs(3855) <= layer2_outputs(11311);
    outputs(3856) <= (layer2_outputs(6605)) and (layer2_outputs(8811));
    outputs(3857) <= not(layer2_outputs(5135));
    outputs(3858) <= layer2_outputs(2691);
    outputs(3859) <= layer2_outputs(7);
    outputs(3860) <= not(layer2_outputs(1262));
    outputs(3861) <= layer2_outputs(7033);
    outputs(3862) <= not((layer2_outputs(6964)) xor (layer2_outputs(3829)));
    outputs(3863) <= layer2_outputs(7330);
    outputs(3864) <= not(layer2_outputs(11975));
    outputs(3865) <= layer2_outputs(1296);
    outputs(3866) <= not((layer2_outputs(7799)) xor (layer2_outputs(4401)));
    outputs(3867) <= not(layer2_outputs(9982));
    outputs(3868) <= (layer2_outputs(6169)) xor (layer2_outputs(6221));
    outputs(3869) <= layer2_outputs(3506);
    outputs(3870) <= layer2_outputs(7098);
    outputs(3871) <= not(layer2_outputs(4371));
    outputs(3872) <= layer2_outputs(5651);
    outputs(3873) <= layer2_outputs(10880);
    outputs(3874) <= (layer2_outputs(6766)) xor (layer2_outputs(1184));
    outputs(3875) <= layer2_outputs(4970);
    outputs(3876) <= not(layer2_outputs(12504));
    outputs(3877) <= not(layer2_outputs(11776));
    outputs(3878) <= not((layer2_outputs(6103)) or (layer2_outputs(5723)));
    outputs(3879) <= not(layer2_outputs(3126));
    outputs(3880) <= not(layer2_outputs(10329)) or (layer2_outputs(7800));
    outputs(3881) <= (layer2_outputs(10818)) xor (layer2_outputs(11919));
    outputs(3882) <= not(layer2_outputs(3380)) or (layer2_outputs(6307));
    outputs(3883) <= not(layer2_outputs(8375));
    outputs(3884) <= not(layer2_outputs(10883));
    outputs(3885) <= (layer2_outputs(12244)) or (layer2_outputs(11747));
    outputs(3886) <= layer2_outputs(11020);
    outputs(3887) <= not(layer2_outputs(6978));
    outputs(3888) <= not((layer2_outputs(6194)) or (layer2_outputs(7251)));
    outputs(3889) <= layer2_outputs(3165);
    outputs(3890) <= not((layer2_outputs(4427)) xor (layer2_outputs(12568)));
    outputs(3891) <= (layer2_outputs(9797)) xor (layer2_outputs(8958));
    outputs(3892) <= (layer2_outputs(11316)) and not (layer2_outputs(4856));
    outputs(3893) <= not((layer2_outputs(2721)) xor (layer2_outputs(11596)));
    outputs(3894) <= layer2_outputs(12705);
    outputs(3895) <= (layer2_outputs(2141)) and not (layer2_outputs(5921));
    outputs(3896) <= layer2_outputs(5284);
    outputs(3897) <= not((layer2_outputs(2709)) xor (layer2_outputs(2193)));
    outputs(3898) <= not(layer2_outputs(7060));
    outputs(3899) <= layer2_outputs(1041);
    outputs(3900) <= not(layer2_outputs(9839));
    outputs(3901) <= (layer2_outputs(9820)) xor (layer2_outputs(5471));
    outputs(3902) <= layer2_outputs(5965);
    outputs(3903) <= not(layer2_outputs(5653));
    outputs(3904) <= layer2_outputs(3331);
    outputs(3905) <= not(layer2_outputs(9193));
    outputs(3906) <= layer2_outputs(12659);
    outputs(3907) <= not((layer2_outputs(12487)) xor (layer2_outputs(1103)));
    outputs(3908) <= layer2_outputs(3347);
    outputs(3909) <= not((layer2_outputs(6876)) xor (layer2_outputs(10412)));
    outputs(3910) <= layer2_outputs(11157);
    outputs(3911) <= (layer2_outputs(1589)) and (layer2_outputs(4315));
    outputs(3912) <= (layer2_outputs(740)) xor (layer2_outputs(3159));
    outputs(3913) <= (layer2_outputs(7639)) or (layer2_outputs(11918));
    outputs(3914) <= not(layer2_outputs(313));
    outputs(3915) <= (layer2_outputs(9209)) xor (layer2_outputs(11042));
    outputs(3916) <= layer2_outputs(4327);
    outputs(3917) <= (layer2_outputs(12099)) and not (layer2_outputs(6220));
    outputs(3918) <= (layer2_outputs(5333)) and not (layer2_outputs(8482));
    outputs(3919) <= not(layer2_outputs(10394));
    outputs(3920) <= layer2_outputs(8572);
    outputs(3921) <= layer2_outputs(10722);
    outputs(3922) <= not(layer2_outputs(2385));
    outputs(3923) <= not(layer2_outputs(3086));
    outputs(3924) <= not(layer2_outputs(3468));
    outputs(3925) <= not(layer2_outputs(7408));
    outputs(3926) <= layer2_outputs(9132);
    outputs(3927) <= layer2_outputs(2200);
    outputs(3928) <= not(layer2_outputs(2336));
    outputs(3929) <= layer2_outputs(10557);
    outputs(3930) <= not((layer2_outputs(6019)) xor (layer2_outputs(10532)));
    outputs(3931) <= (layer2_outputs(5120)) xor (layer2_outputs(8098));
    outputs(3932) <= not((layer2_outputs(3956)) xor (layer2_outputs(11916)));
    outputs(3933) <= (layer2_outputs(6400)) xor (layer2_outputs(11310));
    outputs(3934) <= not((layer2_outputs(7830)) xor (layer2_outputs(6134)));
    outputs(3935) <= (layer2_outputs(11558)) xor (layer2_outputs(1711));
    outputs(3936) <= not(layer2_outputs(7983));
    outputs(3937) <= (layer2_outputs(1558)) xor (layer2_outputs(5220));
    outputs(3938) <= not(layer2_outputs(5600));
    outputs(3939) <= not((layer2_outputs(6559)) xor (layer2_outputs(12361)));
    outputs(3940) <= not(layer2_outputs(2919));
    outputs(3941) <= (layer2_outputs(8354)) xor (layer2_outputs(1399));
    outputs(3942) <= layer2_outputs(6537);
    outputs(3943) <= not((layer2_outputs(9950)) xor (layer2_outputs(440)));
    outputs(3944) <= (layer2_outputs(7284)) xor (layer2_outputs(3397));
    outputs(3945) <= not((layer2_outputs(12482)) xor (layer2_outputs(8473)));
    outputs(3946) <= (layer2_outputs(1319)) and not (layer2_outputs(12765));
    outputs(3947) <= (layer2_outputs(12038)) and not (layer2_outputs(8404));
    outputs(3948) <= layer2_outputs(5704);
    outputs(3949) <= not((layer2_outputs(7665)) xor (layer2_outputs(6491)));
    outputs(3950) <= not(layer2_outputs(6523));
    outputs(3951) <= not(layer2_outputs(12717));
    outputs(3952) <= not((layer2_outputs(12102)) xor (layer2_outputs(9278)));
    outputs(3953) <= not(layer2_outputs(9659));
    outputs(3954) <= layer2_outputs(5519);
    outputs(3955) <= not(layer2_outputs(8246));
    outputs(3956) <= not((layer2_outputs(10575)) or (layer2_outputs(1527)));
    outputs(3957) <= not(layer2_outputs(2686));
    outputs(3958) <= layer2_outputs(10388);
    outputs(3959) <= not(layer2_outputs(12488)) or (layer2_outputs(10123));
    outputs(3960) <= layer2_outputs(791);
    outputs(3961) <= not(layer2_outputs(537)) or (layer2_outputs(235));
    outputs(3962) <= layer2_outputs(11531);
    outputs(3963) <= not(layer2_outputs(12536));
    outputs(3964) <= not((layer2_outputs(4330)) or (layer2_outputs(10855)));
    outputs(3965) <= not((layer2_outputs(442)) xor (layer2_outputs(11009)));
    outputs(3966) <= not(layer2_outputs(6794));
    outputs(3967) <= not(layer2_outputs(5695));
    outputs(3968) <= not((layer2_outputs(11290)) xor (layer2_outputs(6980)));
    outputs(3969) <= not((layer2_outputs(4787)) xor (layer2_outputs(2884)));
    outputs(3970) <= layer2_outputs(12013);
    outputs(3971) <= not(layer2_outputs(4309));
    outputs(3972) <= (layer2_outputs(3266)) xor (layer2_outputs(7486));
    outputs(3973) <= layer2_outputs(9459);
    outputs(3974) <= not(layer2_outputs(8936)) or (layer2_outputs(11469));
    outputs(3975) <= layer2_outputs(10885);
    outputs(3976) <= not((layer2_outputs(4841)) and (layer2_outputs(10073)));
    outputs(3977) <= not(layer2_outputs(9599)) or (layer2_outputs(8506));
    outputs(3978) <= not(layer2_outputs(7470));
    outputs(3979) <= not(layer2_outputs(97));
    outputs(3980) <= (layer2_outputs(8780)) and not (layer2_outputs(2026));
    outputs(3981) <= layer2_outputs(301);
    outputs(3982) <= layer2_outputs(6644);
    outputs(3983) <= not(layer2_outputs(3896));
    outputs(3984) <= layer2_outputs(3623);
    outputs(3985) <= layer2_outputs(11844);
    outputs(3986) <= layer2_outputs(11897);
    outputs(3987) <= not((layer2_outputs(10931)) xor (layer2_outputs(11934)));
    outputs(3988) <= (layer2_outputs(866)) and (layer2_outputs(6068));
    outputs(3989) <= not((layer2_outputs(4508)) or (layer2_outputs(2324)));
    outputs(3990) <= (layer2_outputs(11768)) xor (layer2_outputs(2495));
    outputs(3991) <= not((layer2_outputs(8973)) xor (layer2_outputs(6547)));
    outputs(3992) <= not(layer2_outputs(12165));
    outputs(3993) <= layer2_outputs(12507);
    outputs(3994) <= (layer2_outputs(9983)) and not (layer2_outputs(6288));
    outputs(3995) <= layer2_outputs(2605);
    outputs(3996) <= not(layer2_outputs(8554));
    outputs(3997) <= not(layer2_outputs(4490));
    outputs(3998) <= (layer2_outputs(4426)) or (layer2_outputs(12754));
    outputs(3999) <= (layer2_outputs(3218)) and (layer2_outputs(8492));
    outputs(4000) <= (layer2_outputs(12171)) and (layer2_outputs(12747));
    outputs(4001) <= not(layer2_outputs(1635));
    outputs(4002) <= layer2_outputs(9393);
    outputs(4003) <= (layer2_outputs(7595)) xor (layer2_outputs(9735));
    outputs(4004) <= (layer2_outputs(3865)) and (layer2_outputs(3844));
    outputs(4005) <= (layer2_outputs(1581)) xor (layer2_outputs(10854));
    outputs(4006) <= not(layer2_outputs(6241));
    outputs(4007) <= layer2_outputs(3815);
    outputs(4008) <= not(layer2_outputs(7465));
    outputs(4009) <= layer2_outputs(10957);
    outputs(4010) <= not(layer2_outputs(6886));
    outputs(4011) <= not(layer2_outputs(10474)) or (layer2_outputs(672));
    outputs(4012) <= layer2_outputs(5828);
    outputs(4013) <= not(layer2_outputs(10202));
    outputs(4014) <= (layer2_outputs(7330)) and not (layer2_outputs(112));
    outputs(4015) <= layer2_outputs(10089);
    outputs(4016) <= layer2_outputs(8925);
    outputs(4017) <= layer2_outputs(9844);
    outputs(4018) <= layer2_outputs(2757);
    outputs(4019) <= (layer2_outputs(421)) xor (layer2_outputs(8203));
    outputs(4020) <= (layer2_outputs(7872)) xor (layer2_outputs(8494));
    outputs(4021) <= (layer2_outputs(4944)) xor (layer2_outputs(8322));
    outputs(4022) <= (layer2_outputs(8839)) and not (layer2_outputs(1659));
    outputs(4023) <= not(layer2_outputs(9411));
    outputs(4024) <= not(layer2_outputs(10217));
    outputs(4025) <= not(layer2_outputs(8988));
    outputs(4026) <= not(layer2_outputs(10995));
    outputs(4027) <= not(layer2_outputs(450));
    outputs(4028) <= (layer2_outputs(3508)) xor (layer2_outputs(8267));
    outputs(4029) <= not((layer2_outputs(1678)) xor (layer2_outputs(3593)));
    outputs(4030) <= (layer2_outputs(3511)) xor (layer2_outputs(492));
    outputs(4031) <= layer2_outputs(8837);
    outputs(4032) <= not(layer2_outputs(2292));
    outputs(4033) <= not(layer2_outputs(3793));
    outputs(4034) <= (layer2_outputs(6498)) or (layer2_outputs(311));
    outputs(4035) <= layer2_outputs(2714);
    outputs(4036) <= layer2_outputs(12735);
    outputs(4037) <= (layer2_outputs(10366)) and not (layer2_outputs(10631));
    outputs(4038) <= not(layer2_outputs(4136));
    outputs(4039) <= not((layer2_outputs(7907)) xor (layer2_outputs(12066)));
    outputs(4040) <= (layer2_outputs(3570)) and (layer2_outputs(5336));
    outputs(4041) <= (layer2_outputs(10116)) and not (layer2_outputs(2823));
    outputs(4042) <= not((layer2_outputs(493)) xor (layer2_outputs(80)));
    outputs(4043) <= layer2_outputs(164);
    outputs(4044) <= not(layer2_outputs(4898));
    outputs(4045) <= not(layer2_outputs(8736)) or (layer2_outputs(4740));
    outputs(4046) <= not((layer2_outputs(8841)) xor (layer2_outputs(6842)));
    outputs(4047) <= layer2_outputs(7714);
    outputs(4048) <= (layer2_outputs(2444)) xor (layer2_outputs(4903));
    outputs(4049) <= layer2_outputs(5955);
    outputs(4050) <= (layer2_outputs(3082)) xor (layer2_outputs(3628));
    outputs(4051) <= not(layer2_outputs(692));
    outputs(4052) <= (layer2_outputs(7753)) xor (layer2_outputs(6332));
    outputs(4053) <= not(layer2_outputs(1002));
    outputs(4054) <= (layer2_outputs(370)) or (layer2_outputs(436));
    outputs(4055) <= (layer2_outputs(1040)) xor (layer2_outputs(12379));
    outputs(4056) <= not(layer2_outputs(12185)) or (layer2_outputs(9140));
    outputs(4057) <= layer2_outputs(9302);
    outputs(4058) <= not(layer2_outputs(5652));
    outputs(4059) <= layer2_outputs(3673);
    outputs(4060) <= not(layer2_outputs(8640));
    outputs(4061) <= (layer2_outputs(1989)) xor (layer2_outputs(8306));
    outputs(4062) <= layer2_outputs(10574);
    outputs(4063) <= not(layer2_outputs(5107));
    outputs(4064) <= not((layer2_outputs(8576)) or (layer2_outputs(1914)));
    outputs(4065) <= (layer2_outputs(9902)) and not (layer2_outputs(2950));
    outputs(4066) <= not(layer2_outputs(2529));
    outputs(4067) <= layer2_outputs(5565);
    outputs(4068) <= layer2_outputs(1799);
    outputs(4069) <= not((layer2_outputs(4348)) xor (layer2_outputs(9167)));
    outputs(4070) <= not((layer2_outputs(8733)) xor (layer2_outputs(6987)));
    outputs(4071) <= not((layer2_outputs(11688)) xor (layer2_outputs(10803)));
    outputs(4072) <= (layer2_outputs(2273)) xor (layer2_outputs(9786));
    outputs(4073) <= (layer2_outputs(12320)) and not (layer2_outputs(9500));
    outputs(4074) <= layer2_outputs(2314);
    outputs(4075) <= not((layer2_outputs(9202)) xor (layer2_outputs(9715)));
    outputs(4076) <= (layer2_outputs(1787)) xor (layer2_outputs(2340));
    outputs(4077) <= (layer2_outputs(10034)) and not (layer2_outputs(10143));
    outputs(4078) <= (layer2_outputs(12062)) xor (layer2_outputs(3848));
    outputs(4079) <= (layer2_outputs(7105)) xor (layer2_outputs(982));
    outputs(4080) <= (layer2_outputs(7897)) and not (layer2_outputs(11837));
    outputs(4081) <= not(layer2_outputs(1759));
    outputs(4082) <= layer2_outputs(5124);
    outputs(4083) <= (layer2_outputs(4457)) and not (layer2_outputs(2432));
    outputs(4084) <= not((layer2_outputs(2694)) and (layer2_outputs(991)));
    outputs(4085) <= layer2_outputs(2804);
    outputs(4086) <= (layer2_outputs(1327)) xor (layer2_outputs(11435));
    outputs(4087) <= not((layer2_outputs(6380)) and (layer2_outputs(2696)));
    outputs(4088) <= not((layer2_outputs(72)) xor (layer2_outputs(1701)));
    outputs(4089) <= not(layer2_outputs(12198));
    outputs(4090) <= not(layer2_outputs(9581));
    outputs(4091) <= not(layer2_outputs(1676));
    outputs(4092) <= (layer2_outputs(12552)) or (layer2_outputs(557));
    outputs(4093) <= (layer2_outputs(7493)) xor (layer2_outputs(10655));
    outputs(4094) <= (layer2_outputs(9153)) and not (layer2_outputs(12474));
    outputs(4095) <= (layer2_outputs(2903)) and (layer2_outputs(2328));
    outputs(4096) <= (layer2_outputs(1198)) xor (layer2_outputs(10753));
    outputs(4097) <= (layer2_outputs(9369)) and (layer2_outputs(11996));
    outputs(4098) <= not((layer2_outputs(8919)) and (layer2_outputs(6383)));
    outputs(4099) <= not((layer2_outputs(4533)) xor (layer2_outputs(3744)));
    outputs(4100) <= not(layer2_outputs(12399)) or (layer2_outputs(5359));
    outputs(4101) <= not((layer2_outputs(11829)) xor (layer2_outputs(9378)));
    outputs(4102) <= layer2_outputs(8426);
    outputs(4103) <= layer2_outputs(6933);
    outputs(4104) <= (layer2_outputs(4897)) xor (layer2_outputs(6180));
    outputs(4105) <= not(layer2_outputs(3890));
    outputs(4106) <= not(layer2_outputs(5414));
    outputs(4107) <= not(layer2_outputs(3962));
    outputs(4108) <= not((layer2_outputs(5349)) xor (layer2_outputs(5129)));
    outputs(4109) <= layer2_outputs(7505);
    outputs(4110) <= (layer2_outputs(5395)) and not (layer2_outputs(1876));
    outputs(4111) <= not(layer2_outputs(4047));
    outputs(4112) <= not(layer2_outputs(10792));
    outputs(4113) <= not((layer2_outputs(4174)) xor (layer2_outputs(10590)));
    outputs(4114) <= layer2_outputs(8950);
    outputs(4115) <= not(layer2_outputs(1147));
    outputs(4116) <= (layer2_outputs(12774)) and (layer2_outputs(11028));
    outputs(4117) <= layer2_outputs(5713);
    outputs(4118) <= not((layer2_outputs(5629)) xor (layer2_outputs(2196)));
    outputs(4119) <= (layer2_outputs(274)) xor (layer2_outputs(6476));
    outputs(4120) <= (layer2_outputs(1734)) xor (layer2_outputs(5768));
    outputs(4121) <= layer2_outputs(12716);
    outputs(4122) <= layer2_outputs(5111);
    outputs(4123) <= not(layer2_outputs(8712)) or (layer2_outputs(3738));
    outputs(4124) <= layer2_outputs(6403);
    outputs(4125) <= layer2_outputs(7002);
    outputs(4126) <= layer2_outputs(9183);
    outputs(4127) <= (layer2_outputs(10919)) xor (layer2_outputs(11955));
    outputs(4128) <= (layer2_outputs(10105)) xor (layer2_outputs(12532));
    outputs(4129) <= (layer2_outputs(8034)) and (layer2_outputs(471));
    outputs(4130) <= not(layer2_outputs(1874));
    outputs(4131) <= not(layer2_outputs(8199));
    outputs(4132) <= (layer2_outputs(10513)) xor (layer2_outputs(6473));
    outputs(4133) <= (layer2_outputs(11071)) and not (layer2_outputs(3425));
    outputs(4134) <= layer2_outputs(2528);
    outputs(4135) <= layer2_outputs(7064);
    outputs(4136) <= not((layer2_outputs(12387)) or (layer2_outputs(2515)));
    outputs(4137) <= layer2_outputs(12680);
    outputs(4138) <= (layer2_outputs(8541)) and (layer2_outputs(2964));
    outputs(4139) <= layer2_outputs(5977);
    outputs(4140) <= (layer2_outputs(10090)) xor (layer2_outputs(7786));
    outputs(4141) <= (layer2_outputs(3611)) or (layer2_outputs(11496));
    outputs(4142) <= layer2_outputs(10111);
    outputs(4143) <= layer2_outputs(7053);
    outputs(4144) <= not(layer2_outputs(9036));
    outputs(4145) <= not((layer2_outputs(8930)) xor (layer2_outputs(6665)));
    outputs(4146) <= (layer2_outputs(3321)) xor (layer2_outputs(11023));
    outputs(4147) <= layer2_outputs(1592);
    outputs(4148) <= not(layer2_outputs(5311));
    outputs(4149) <= layer2_outputs(10877);
    outputs(4150) <= layer2_outputs(5350);
    outputs(4151) <= (layer2_outputs(12246)) xor (layer2_outputs(12220));
    outputs(4152) <= not(layer2_outputs(7235)) or (layer2_outputs(188));
    outputs(4153) <= not(layer2_outputs(12462));
    outputs(4154) <= not(layer2_outputs(2207));
    outputs(4155) <= (layer2_outputs(3681)) and not (layer2_outputs(5367));
    outputs(4156) <= layer2_outputs(7026);
    outputs(4157) <= not((layer2_outputs(10362)) xor (layer2_outputs(8686)));
    outputs(4158) <= not(layer2_outputs(8009));
    outputs(4159) <= not(layer2_outputs(8010));
    outputs(4160) <= layer2_outputs(594);
    outputs(4161) <= (layer2_outputs(117)) xor (layer2_outputs(1258));
    outputs(4162) <= (layer2_outputs(549)) and (layer2_outputs(1476));
    outputs(4163) <= not(layer2_outputs(2140));
    outputs(4164) <= layer2_outputs(12445);
    outputs(4165) <= not(layer2_outputs(6165)) or (layer2_outputs(5234));
    outputs(4166) <= (layer2_outputs(1670)) and not (layer2_outputs(12464));
    outputs(4167) <= layer2_outputs(4434);
    outputs(4168) <= (layer2_outputs(11279)) xor (layer2_outputs(10270));
    outputs(4169) <= (layer2_outputs(6299)) xor (layer2_outputs(446));
    outputs(4170) <= not(layer2_outputs(4063));
    outputs(4171) <= layer2_outputs(9789);
    outputs(4172) <= (layer2_outputs(7807)) xor (layer2_outputs(10556));
    outputs(4173) <= layer2_outputs(2943);
    outputs(4174) <= not(layer2_outputs(7776));
    outputs(4175) <= not((layer2_outputs(89)) xor (layer2_outputs(2709)));
    outputs(4176) <= not(layer2_outputs(6113));
    outputs(4177) <= not((layer2_outputs(3860)) and (layer2_outputs(5980)));
    outputs(4178) <= not(layer2_outputs(4729)) or (layer2_outputs(2001));
    outputs(4179) <= layer2_outputs(549);
    outputs(4180) <= layer2_outputs(7040);
    outputs(4181) <= (layer2_outputs(3921)) xor (layer2_outputs(4205));
    outputs(4182) <= not(layer2_outputs(2044));
    outputs(4183) <= not(layer2_outputs(3905));
    outputs(4184) <= not(layer2_outputs(3895));
    outputs(4185) <= layer2_outputs(10639);
    outputs(4186) <= (layer2_outputs(6744)) xor (layer2_outputs(3511));
    outputs(4187) <= not(layer2_outputs(7204)) or (layer2_outputs(7813));
    outputs(4188) <= layer2_outputs(3104);
    outputs(4189) <= not(layer2_outputs(233));
    outputs(4190) <= layer2_outputs(12616);
    outputs(4191) <= not(layer2_outputs(9625));
    outputs(4192) <= not((layer2_outputs(11968)) or (layer2_outputs(11026)));
    outputs(4193) <= layer2_outputs(1483);
    outputs(4194) <= (layer2_outputs(500)) xor (layer2_outputs(251));
    outputs(4195) <= layer2_outputs(10983);
    outputs(4196) <= not(layer2_outputs(4680));
    outputs(4197) <= (layer2_outputs(125)) and not (layer2_outputs(3655));
    outputs(4198) <= not(layer2_outputs(6471));
    outputs(4199) <= layer2_outputs(8065);
    outputs(4200) <= layer2_outputs(5122);
    outputs(4201) <= (layer2_outputs(12467)) and (layer2_outputs(3110));
    outputs(4202) <= layer2_outputs(232);
    outputs(4203) <= not((layer2_outputs(4551)) xor (layer2_outputs(8232)));
    outputs(4204) <= not((layer2_outputs(11972)) xor (layer2_outputs(4621)));
    outputs(4205) <= layer2_outputs(6816);
    outputs(4206) <= not((layer2_outputs(5257)) or (layer2_outputs(9222)));
    outputs(4207) <= not(layer2_outputs(10103));
    outputs(4208) <= layer2_outputs(1631);
    outputs(4209) <= layer2_outputs(8975);
    outputs(4210) <= layer2_outputs(7373);
    outputs(4211) <= not((layer2_outputs(3108)) or (layer2_outputs(7634)));
    outputs(4212) <= (layer2_outputs(12255)) xor (layer2_outputs(10124));
    outputs(4213) <= layer2_outputs(10839);
    outputs(4214) <= not(layer2_outputs(10687)) or (layer2_outputs(1223));
    outputs(4215) <= layer2_outputs(8102);
    outputs(4216) <= (layer2_outputs(3204)) xor (layer2_outputs(5696));
    outputs(4217) <= not((layer2_outputs(3856)) or (layer2_outputs(7671)));
    outputs(4218) <= layer2_outputs(2969);
    outputs(4219) <= not((layer2_outputs(7857)) xor (layer2_outputs(4810)));
    outputs(4220) <= not(layer2_outputs(7412));
    outputs(4221) <= not(layer2_outputs(80));
    outputs(4222) <= layer2_outputs(5852);
    outputs(4223) <= not((layer2_outputs(7889)) xor (layer2_outputs(3648)));
    outputs(4224) <= (layer2_outputs(11256)) and (layer2_outputs(8153));
    outputs(4225) <= layer2_outputs(9078);
    outputs(4226) <= layer2_outputs(9668);
    outputs(4227) <= layer2_outputs(4626);
    outputs(4228) <= (layer2_outputs(7987)) xor (layer2_outputs(11506));
    outputs(4229) <= (layer2_outputs(8882)) xor (layer2_outputs(8635));
    outputs(4230) <= layer2_outputs(10711);
    outputs(4231) <= not(layer2_outputs(12336));
    outputs(4232) <= layer2_outputs(2341);
    outputs(4233) <= layer2_outputs(280);
    outputs(4234) <= not((layer2_outputs(9795)) xor (layer2_outputs(6898)));
    outputs(4235) <= (layer2_outputs(4074)) xor (layer2_outputs(8184));
    outputs(4236) <= layer2_outputs(3213);
    outputs(4237) <= not(layer2_outputs(9806));
    outputs(4238) <= (layer2_outputs(3767)) xor (layer2_outputs(6864));
    outputs(4239) <= not(layer2_outputs(8785));
    outputs(4240) <= (layer2_outputs(7450)) xor (layer2_outputs(5106));
    outputs(4241) <= not((layer2_outputs(4050)) xor (layer2_outputs(9687)));
    outputs(4242) <= (layer2_outputs(10110)) xor (layer2_outputs(20));
    outputs(4243) <= layer2_outputs(11266);
    outputs(4244) <= layer2_outputs(11778);
    outputs(4245) <= (layer2_outputs(10096)) xor (layer2_outputs(6320));
    outputs(4246) <= not(layer2_outputs(10276));
    outputs(4247) <= not(layer2_outputs(7181));
    outputs(4248) <= (layer2_outputs(708)) xor (layer2_outputs(1394));
    outputs(4249) <= not(layer2_outputs(7106));
    outputs(4250) <= layer2_outputs(5305);
    outputs(4251) <= not(layer2_outputs(1933));
    outputs(4252) <= not((layer2_outputs(11719)) xor (layer2_outputs(4743)));
    outputs(4253) <= layer2_outputs(6913);
    outputs(4254) <= not(layer2_outputs(11792));
    outputs(4255) <= (layer2_outputs(897)) xor (layer2_outputs(4743));
    outputs(4256) <= not(layer2_outputs(7847));
    outputs(4257) <= (layer2_outputs(7900)) and not (layer2_outputs(12526));
    outputs(4258) <= not(layer2_outputs(6453));
    outputs(4259) <= not(layer2_outputs(12105));
    outputs(4260) <= layer2_outputs(4393);
    outputs(4261) <= layer2_outputs(2707);
    outputs(4262) <= not(layer2_outputs(11514));
    outputs(4263) <= not((layer2_outputs(4534)) xor (layer2_outputs(3774)));
    outputs(4264) <= not(layer2_outputs(10879));
    outputs(4265) <= (layer2_outputs(11371)) xor (layer2_outputs(1806));
    outputs(4266) <= not((layer2_outputs(10652)) xor (layer2_outputs(2972)));
    outputs(4267) <= not((layer2_outputs(6080)) or (layer2_outputs(9129)));
    outputs(4268) <= layer2_outputs(11628);
    outputs(4269) <= not((layer2_outputs(3690)) xor (layer2_outputs(12317)));
    outputs(4270) <= layer2_outputs(1664);
    outputs(4271) <= layer2_outputs(11047);
    outputs(4272) <= layer2_outputs(606);
    outputs(4273) <= (layer2_outputs(11608)) xor (layer2_outputs(2583));
    outputs(4274) <= layer2_outputs(10071);
    outputs(4275) <= not((layer2_outputs(4415)) xor (layer2_outputs(4191)));
    outputs(4276) <= layer2_outputs(3871);
    outputs(4277) <= (layer2_outputs(5053)) and not (layer2_outputs(5538));
    outputs(4278) <= not(layer2_outputs(2609));
    outputs(4279) <= (layer2_outputs(4012)) and (layer2_outputs(7438));
    outputs(4280) <= (layer2_outputs(7681)) xor (layer2_outputs(4687));
    outputs(4281) <= not(layer2_outputs(4920));
    outputs(4282) <= (layer2_outputs(2486)) or (layer2_outputs(583));
    outputs(4283) <= not((layer2_outputs(11859)) xor (layer2_outputs(4353)));
    outputs(4284) <= not((layer2_outputs(1602)) xor (layer2_outputs(2360)));
    outputs(4285) <= layer2_outputs(8407);
    outputs(4286) <= (layer2_outputs(6074)) xor (layer2_outputs(9711));
    outputs(4287) <= not(layer2_outputs(11159));
    outputs(4288) <= layer2_outputs(8162);
    outputs(4289) <= (layer2_outputs(9657)) xor (layer2_outputs(10783));
    outputs(4290) <= (layer2_outputs(12200)) xor (layer2_outputs(5218));
    outputs(4291) <= layer2_outputs(9618);
    outputs(4292) <= layer2_outputs(9349);
    outputs(4293) <= not(layer2_outputs(10338));
    outputs(4294) <= not((layer2_outputs(2772)) xor (layer2_outputs(4219)));
    outputs(4295) <= (layer2_outputs(10212)) or (layer2_outputs(8727));
    outputs(4296) <= (layer2_outputs(5720)) xor (layer2_outputs(1579));
    outputs(4297) <= layer2_outputs(6859);
    outputs(4298) <= layer2_outputs(1017);
    outputs(4299) <= layer2_outputs(12514);
    outputs(4300) <= (layer2_outputs(6133)) and not (layer2_outputs(2923));
    outputs(4301) <= not(layer2_outputs(7355));
    outputs(4302) <= (layer2_outputs(4400)) xor (layer2_outputs(5098));
    outputs(4303) <= not(layer2_outputs(11578));
    outputs(4304) <= not((layer2_outputs(2704)) and (layer2_outputs(11851)));
    outputs(4305) <= not(layer2_outputs(10488));
    outputs(4306) <= (layer2_outputs(10876)) xor (layer2_outputs(1364));
    outputs(4307) <= (layer2_outputs(1808)) xor (layer2_outputs(8519));
    outputs(4308) <= (layer2_outputs(9635)) or (layer2_outputs(5708));
    outputs(4309) <= layer2_outputs(6722);
    outputs(4310) <= not(layer2_outputs(2553));
    outputs(4311) <= layer2_outputs(2151);
    outputs(4312) <= (layer2_outputs(2204)) xor (layer2_outputs(4167));
    outputs(4313) <= not(layer2_outputs(1297));
    outputs(4314) <= not(layer2_outputs(1904)) or (layer2_outputs(4249));
    outputs(4315) <= not(layer2_outputs(713));
    outputs(4316) <= not(layer2_outputs(5483));
    outputs(4317) <= (layer2_outputs(11407)) or (layer2_outputs(5507));
    outputs(4318) <= layer2_outputs(8933);
    outputs(4319) <= not(layer2_outputs(1920));
    outputs(4320) <= not(layer2_outputs(11999));
    outputs(4321) <= not((layer2_outputs(8893)) xor (layer2_outputs(5804)));
    outputs(4322) <= (layer2_outputs(2681)) and not (layer2_outputs(12613));
    outputs(4323) <= layer2_outputs(1021);
    outputs(4324) <= not(layer2_outputs(8135));
    outputs(4325) <= not(layer2_outputs(3173));
    outputs(4326) <= layer2_outputs(893);
    outputs(4327) <= layer2_outputs(5021);
    outputs(4328) <= layer2_outputs(4627);
    outputs(4329) <= not(layer2_outputs(12481));
    outputs(4330) <= layer2_outputs(587);
    outputs(4331) <= (layer2_outputs(6854)) and not (layer2_outputs(930));
    outputs(4332) <= not((layer2_outputs(3071)) xor (layer2_outputs(8632)));
    outputs(4333) <= layer2_outputs(7262);
    outputs(4334) <= not((layer2_outputs(12082)) xor (layer2_outputs(8061)));
    outputs(4335) <= not(layer2_outputs(4590));
    outputs(4336) <= not((layer2_outputs(9259)) xor (layer2_outputs(10304)));
    outputs(4337) <= layer2_outputs(3418);
    outputs(4338) <= (layer2_outputs(8678)) and not (layer2_outputs(5821));
    outputs(4339) <= not((layer2_outputs(7064)) xor (layer2_outputs(7281)));
    outputs(4340) <= layer2_outputs(6698);
    outputs(4341) <= (layer2_outputs(4510)) xor (layer2_outputs(8299));
    outputs(4342) <= layer2_outputs(12583);
    outputs(4343) <= not(layer2_outputs(2722));
    outputs(4344) <= not(layer2_outputs(5532));
    outputs(4345) <= not((layer2_outputs(9310)) xor (layer2_outputs(2816)));
    outputs(4346) <= (layer2_outputs(5179)) xor (layer2_outputs(2464));
    outputs(4347) <= not(layer2_outputs(1064));
    outputs(4348) <= layer2_outputs(4121);
    outputs(4349) <= (layer2_outputs(10986)) xor (layer2_outputs(4340));
    outputs(4350) <= (layer2_outputs(1745)) or (layer2_outputs(9450));
    outputs(4351) <= not(layer2_outputs(11603));
    outputs(4352) <= layer2_outputs(7155);
    outputs(4353) <= (layer2_outputs(6810)) xor (layer2_outputs(11242));
    outputs(4354) <= (layer2_outputs(12675)) and not (layer2_outputs(4666));
    outputs(4355) <= layer2_outputs(7757);
    outputs(4356) <= layer2_outputs(8142);
    outputs(4357) <= not(layer2_outputs(8078));
    outputs(4358) <= layer2_outputs(8016);
    outputs(4359) <= (layer2_outputs(12552)) or (layer2_outputs(9936));
    outputs(4360) <= not(layer2_outputs(10678)) or (layer2_outputs(10439));
    outputs(4361) <= (layer2_outputs(6869)) xor (layer2_outputs(1658));
    outputs(4362) <= not(layer2_outputs(4333)) or (layer2_outputs(8235));
    outputs(4363) <= layer2_outputs(8549);
    outputs(4364) <= not((layer2_outputs(5326)) xor (layer2_outputs(7629)));
    outputs(4365) <= not((layer2_outputs(12228)) xor (layer2_outputs(2518)));
    outputs(4366) <= not(layer2_outputs(9803));
    outputs(4367) <= (layer2_outputs(5875)) xor (layer2_outputs(8788));
    outputs(4368) <= (layer2_outputs(12736)) xor (layer2_outputs(3485));
    outputs(4369) <= not((layer2_outputs(11240)) xor (layer2_outputs(109)));
    outputs(4370) <= not(layer2_outputs(293));
    outputs(4371) <= not(layer2_outputs(3433)) or (layer2_outputs(4879));
    outputs(4372) <= not(layer2_outputs(6233));
    outputs(4373) <= not((layer2_outputs(1545)) xor (layer2_outputs(846)));
    outputs(4374) <= not(layer2_outputs(1011));
    outputs(4375) <= layer2_outputs(11113);
    outputs(4376) <= (layer2_outputs(1085)) xor (layer2_outputs(11595));
    outputs(4377) <= layer2_outputs(10727);
    outputs(4378) <= layer2_outputs(7411);
    outputs(4379) <= not((layer2_outputs(7556)) and (layer2_outputs(10431)));
    outputs(4380) <= not(layer2_outputs(7250));
    outputs(4381) <= (layer2_outputs(5849)) or (layer2_outputs(333));
    outputs(4382) <= (layer2_outputs(4926)) xor (layer2_outputs(2841));
    outputs(4383) <= not((layer2_outputs(7346)) xor (layer2_outputs(9160)));
    outputs(4384) <= not(layer2_outputs(5154));
    outputs(4385) <= layer2_outputs(933);
    outputs(4386) <= (layer2_outputs(11247)) xor (layer2_outputs(5610));
    outputs(4387) <= not(layer2_outputs(4410));
    outputs(4388) <= not((layer2_outputs(4473)) xor (layer2_outputs(10361)));
    outputs(4389) <= not(layer2_outputs(12597));
    outputs(4390) <= not(layer2_outputs(7614));
    outputs(4391) <= layer2_outputs(728);
    outputs(4392) <= not((layer2_outputs(1612)) xor (layer2_outputs(6938)));
    outputs(4393) <= (layer2_outputs(5396)) xor (layer2_outputs(12205));
    outputs(4394) <= (layer2_outputs(8481)) and not (layer2_outputs(11968));
    outputs(4395) <= layer2_outputs(10804);
    outputs(4396) <= not(layer2_outputs(4224));
    outputs(4397) <= (layer2_outputs(4360)) and not (layer2_outputs(4783));
    outputs(4398) <= not(layer2_outputs(1366)) or (layer2_outputs(623));
    outputs(4399) <= (layer2_outputs(5347)) xor (layer2_outputs(6535));
    outputs(4400) <= layer2_outputs(3200);
    outputs(4401) <= not((layer2_outputs(3728)) and (layer2_outputs(10661)));
    outputs(4402) <= not(layer2_outputs(10548));
    outputs(4403) <= not((layer2_outputs(8269)) or (layer2_outputs(5592)));
    outputs(4404) <= not(layer2_outputs(538));
    outputs(4405) <= (layer2_outputs(3743)) and not (layer2_outputs(635));
    outputs(4406) <= not((layer2_outputs(8890)) xor (layer2_outputs(4425)));
    outputs(4407) <= layer2_outputs(6789);
    outputs(4408) <= layer2_outputs(7920);
    outputs(4409) <= layer2_outputs(11413);
    outputs(4410) <= not(layer2_outputs(6667));
    outputs(4411) <= layer2_outputs(600);
    outputs(4412) <= layer2_outputs(11736);
    outputs(4413) <= not(layer2_outputs(6538));
    outputs(4414) <= layer2_outputs(7824);
    outputs(4415) <= (layer2_outputs(10287)) xor (layer2_outputs(5727));
    outputs(4416) <= not(layer2_outputs(8674));
    outputs(4417) <= (layer2_outputs(10896)) xor (layer2_outputs(6070));
    outputs(4418) <= not(layer2_outputs(10280));
    outputs(4419) <= layer2_outputs(11916);
    outputs(4420) <= not((layer2_outputs(7837)) xor (layer2_outputs(2564)));
    outputs(4421) <= not((layer2_outputs(1668)) xor (layer2_outputs(10796)));
    outputs(4422) <= not(layer2_outputs(12533));
    outputs(4423) <= (layer2_outputs(2174)) and (layer2_outputs(5198));
    outputs(4424) <= layer2_outputs(7666);
    outputs(4425) <= layer2_outputs(11463);
    outputs(4426) <= not(layer2_outputs(5798));
    outputs(4427) <= layer2_outputs(9535);
    outputs(4428) <= not(layer2_outputs(8906));
    outputs(4429) <= (layer2_outputs(2536)) and (layer2_outputs(3997));
    outputs(4430) <= (layer2_outputs(9454)) and (layer2_outputs(988));
    outputs(4431) <= layer2_outputs(3500);
    outputs(4432) <= not(layer2_outputs(7429));
    outputs(4433) <= not(layer2_outputs(4768));
    outputs(4434) <= (layer2_outputs(7714)) and (layer2_outputs(11844));
    outputs(4435) <= (layer2_outputs(9927)) and not (layer2_outputs(11692));
    outputs(4436) <= not((layer2_outputs(2830)) xor (layer2_outputs(373)));
    outputs(4437) <= (layer2_outputs(4491)) xor (layer2_outputs(4880));
    outputs(4438) <= layer2_outputs(679);
    outputs(4439) <= not((layer2_outputs(3595)) xor (layer2_outputs(11637)));
    outputs(4440) <= layer2_outputs(12411);
    outputs(4441) <= not((layer2_outputs(3637)) or (layer2_outputs(10559)));
    outputs(4442) <= not(layer2_outputs(10076));
    outputs(4443) <= not(layer2_outputs(7021)) or (layer2_outputs(9273));
    outputs(4444) <= not(layer2_outputs(2390)) or (layer2_outputs(607));
    outputs(4445) <= layer2_outputs(7729);
    outputs(4446) <= not(layer2_outputs(6844)) or (layer2_outputs(215));
    outputs(4447) <= (layer2_outputs(500)) and (layer2_outputs(2784));
    outputs(4448) <= not(layer2_outputs(4319));
    outputs(4449) <= not(layer2_outputs(5534));
    outputs(4450) <= not(layer2_outputs(3324));
    outputs(4451) <= layer2_outputs(12448);
    outputs(4452) <= not(layer2_outputs(6893));
    outputs(4453) <= layer2_outputs(8308);
    outputs(4454) <= not((layer2_outputs(3415)) xor (layer2_outputs(11725)));
    outputs(4455) <= layer2_outputs(3549);
    outputs(4456) <= not(layer2_outputs(5233));
    outputs(4457) <= (layer2_outputs(12670)) and (layer2_outputs(2067));
    outputs(4458) <= not(layer2_outputs(48));
    outputs(4459) <= layer2_outputs(6588);
    outputs(4460) <= (layer2_outputs(7035)) xor (layer2_outputs(11749));
    outputs(4461) <= not((layer2_outputs(6306)) xor (layer2_outputs(1619)));
    outputs(4462) <= (layer2_outputs(8)) xor (layer2_outputs(3201));
    outputs(4463) <= (layer2_outputs(1212)) and not (layer2_outputs(2264));
    outputs(4464) <= (layer2_outputs(2965)) xor (layer2_outputs(7581));
    outputs(4465) <= not((layer2_outputs(12060)) xor (layer2_outputs(10259)));
    outputs(4466) <= layer2_outputs(1706);
    outputs(4467) <= layer2_outputs(10070);
    outputs(4468) <= not((layer2_outputs(3044)) xor (layer2_outputs(3586)));
    outputs(4469) <= not((layer2_outputs(4741)) xor (layer2_outputs(1458)));
    outputs(4470) <= layer2_outputs(4417);
    outputs(4471) <= (layer2_outputs(5045)) and not (layer2_outputs(11942));
    outputs(4472) <= (layer2_outputs(9194)) and (layer2_outputs(7383));
    outputs(4473) <= (layer2_outputs(1522)) and not (layer2_outputs(1569));
    outputs(4474) <= not((layer2_outputs(3097)) xor (layer2_outputs(1718)));
    outputs(4475) <= not(layer2_outputs(10297));
    outputs(4476) <= not(layer2_outputs(2718));
    outputs(4477) <= (layer2_outputs(356)) xor (layer2_outputs(10697));
    outputs(4478) <= not((layer2_outputs(11745)) xor (layer2_outputs(2386)));
    outputs(4479) <= layer2_outputs(12161);
    outputs(4480) <= not(layer2_outputs(5667));
    outputs(4481) <= (layer2_outputs(9541)) and (layer2_outputs(6502));
    outputs(4482) <= layer2_outputs(3656);
    outputs(4483) <= not(layer2_outputs(9770)) or (layer2_outputs(1125));
    outputs(4484) <= not(layer2_outputs(5113));
    outputs(4485) <= not((layer2_outputs(6441)) xor (layer2_outputs(8788)));
    outputs(4486) <= layer2_outputs(329);
    outputs(4487) <= not(layer2_outputs(12103));
    outputs(4488) <= not(layer2_outputs(8566));
    outputs(4489) <= not(layer2_outputs(8728));
    outputs(4490) <= (layer2_outputs(3037)) xor (layer2_outputs(11923));
    outputs(4491) <= (layer2_outputs(11840)) xor (layer2_outputs(9390));
    outputs(4492) <= not(layer2_outputs(10210));
    outputs(4493) <= layer2_outputs(3469);
    outputs(4494) <= (layer2_outputs(3165)) xor (layer2_outputs(7003));
    outputs(4495) <= layer2_outputs(10566);
    outputs(4496) <= (layer2_outputs(942)) xor (layer2_outputs(940));
    outputs(4497) <= layer2_outputs(1257);
    outputs(4498) <= (layer2_outputs(11212)) xor (layer2_outputs(4959));
    outputs(4499) <= not((layer2_outputs(765)) xor (layer2_outputs(9060)));
    outputs(4500) <= layer2_outputs(927);
    outputs(4501) <= not((layer2_outputs(3358)) xor (layer2_outputs(7218)));
    outputs(4502) <= (layer2_outputs(2753)) and not (layer2_outputs(11969));
    outputs(4503) <= layer2_outputs(6783);
    outputs(4504) <= (layer2_outputs(6867)) or (layer2_outputs(7667));
    outputs(4505) <= (layer2_outputs(1288)) xor (layer2_outputs(5645));
    outputs(4506) <= not(layer2_outputs(8123));
    outputs(4507) <= not(layer2_outputs(12046));
    outputs(4508) <= not((layer2_outputs(11779)) and (layer2_outputs(138)));
    outputs(4509) <= not(layer2_outputs(11551));
    outputs(4510) <= not((layer2_outputs(1025)) or (layer2_outputs(9999)));
    outputs(4511) <= (layer2_outputs(7663)) or (layer2_outputs(10495));
    outputs(4512) <= not(layer2_outputs(5832));
    outputs(4513) <= not(layer2_outputs(4181));
    outputs(4514) <= (layer2_outputs(8228)) and not (layer2_outputs(4990));
    outputs(4515) <= not((layer2_outputs(4961)) or (layer2_outputs(2284)));
    outputs(4516) <= not(layer2_outputs(12526));
    outputs(4517) <= layer2_outputs(7918);
    outputs(4518) <= not(layer2_outputs(11936));
    outputs(4519) <= not(layer2_outputs(10521)) or (layer2_outputs(12312));
    outputs(4520) <= not(layer2_outputs(4089));
    outputs(4521) <= not(layer2_outputs(10530));
    outputs(4522) <= not((layer2_outputs(2950)) or (layer2_outputs(956)));
    outputs(4523) <= layer2_outputs(5816);
    outputs(4524) <= not(layer2_outputs(10641));
    outputs(4525) <= not((layer2_outputs(32)) xor (layer2_outputs(9887)));
    outputs(4526) <= (layer2_outputs(10180)) and not (layer2_outputs(6758));
    outputs(4527) <= not(layer2_outputs(6612));
    outputs(4528) <= not(layer2_outputs(6108));
    outputs(4529) <= (layer2_outputs(1469)) xor (layer2_outputs(5970));
    outputs(4530) <= (layer2_outputs(418)) xor (layer2_outputs(2800));
    outputs(4531) <= not(layer2_outputs(10697)) or (layer2_outputs(2675));
    outputs(4532) <= not((layer2_outputs(9470)) xor (layer2_outputs(12266)));
    outputs(4533) <= not(layer2_outputs(483));
    outputs(4534) <= layer2_outputs(5732);
    outputs(4535) <= (layer2_outputs(1816)) and (layer2_outputs(4627));
    outputs(4536) <= not(layer2_outputs(6678));
    outputs(4537) <= (layer2_outputs(6000)) and (layer2_outputs(12795));
    outputs(4538) <= layer2_outputs(12078);
    outputs(4539) <= not(layer2_outputs(1636));
    outputs(4540) <= (layer2_outputs(4398)) or (layer2_outputs(10244));
    outputs(4541) <= layer2_outputs(9366);
    outputs(4542) <= (layer2_outputs(5134)) and not (layer2_outputs(12080));
    outputs(4543) <= layer2_outputs(646);
    outputs(4544) <= not(layer2_outputs(8359));
    outputs(4545) <= (layer2_outputs(6245)) xor (layer2_outputs(2478));
    outputs(4546) <= not(layer2_outputs(4635));
    outputs(4547) <= layer2_outputs(8757);
    outputs(4548) <= not((layer2_outputs(11782)) xor (layer2_outputs(811)));
    outputs(4549) <= not(layer2_outputs(7646));
    outputs(4550) <= (layer2_outputs(4598)) xor (layer2_outputs(8425));
    outputs(4551) <= not((layer2_outputs(672)) xor (layer2_outputs(2885)));
    outputs(4552) <= not(layer2_outputs(7646));
    outputs(4553) <= not(layer2_outputs(2065));
    outputs(4554) <= (layer2_outputs(9589)) xor (layer2_outputs(10197));
    outputs(4555) <= (layer2_outputs(2487)) xor (layer2_outputs(2442));
    outputs(4556) <= (layer2_outputs(10962)) and not (layer2_outputs(7742));
    outputs(4557) <= not(layer2_outputs(1998));
    outputs(4558) <= (layer2_outputs(2704)) xor (layer2_outputs(2653));
    outputs(4559) <= not(layer2_outputs(12015));
    outputs(4560) <= (layer2_outputs(1219)) and not (layer2_outputs(4148));
    outputs(4561) <= layer2_outputs(855);
    outputs(4562) <= layer2_outputs(6890);
    outputs(4563) <= not((layer2_outputs(1354)) xor (layer2_outputs(815)));
    outputs(4564) <= (layer2_outputs(12445)) and not (layer2_outputs(10771));
    outputs(4565) <= not(layer2_outputs(1207));
    outputs(4566) <= not(layer2_outputs(11568));
    outputs(4567) <= layer2_outputs(12365);
    outputs(4568) <= not((layer2_outputs(1759)) xor (layer2_outputs(10608)));
    outputs(4569) <= layer2_outputs(6177);
    outputs(4570) <= layer2_outputs(7845);
    outputs(4571) <= (layer2_outputs(8705)) xor (layer2_outputs(2809));
    outputs(4572) <= not(layer2_outputs(11087));
    outputs(4573) <= not(layer2_outputs(7171));
    outputs(4574) <= not(layer2_outputs(1935));
    outputs(4575) <= layer2_outputs(3448);
    outputs(4576) <= not((layer2_outputs(2377)) xor (layer2_outputs(5900)));
    outputs(4577) <= not((layer2_outputs(8254)) xor (layer2_outputs(747)));
    outputs(4578) <= not(layer2_outputs(2671)) or (layer2_outputs(1742));
    outputs(4579) <= layer2_outputs(7168);
    outputs(4580) <= (layer2_outputs(4294)) xor (layer2_outputs(9879));
    outputs(4581) <= not(layer2_outputs(4450)) or (layer2_outputs(2811));
    outputs(4582) <= not(layer2_outputs(9291));
    outputs(4583) <= not((layer2_outputs(12034)) xor (layer2_outputs(3495)));
    outputs(4584) <= not((layer2_outputs(7600)) and (layer2_outputs(5546)));
    outputs(4585) <= not(layer2_outputs(10876));
    outputs(4586) <= not(layer2_outputs(12428));
    outputs(4587) <= not(layer2_outputs(2076));
    outputs(4588) <= not((layer2_outputs(9890)) xor (layer2_outputs(1863)));
    outputs(4589) <= not(layer2_outputs(8992));
    outputs(4590) <= layer2_outputs(5184);
    outputs(4591) <= (layer2_outputs(6777)) xor (layer2_outputs(1142));
    outputs(4592) <= not((layer2_outputs(9649)) or (layer2_outputs(9134)));
    outputs(4593) <= (layer2_outputs(8411)) xor (layer2_outputs(12494));
    outputs(4594) <= (layer2_outputs(4836)) and not (layer2_outputs(6346));
    outputs(4595) <= layer2_outputs(9330);
    outputs(4596) <= not((layer2_outputs(10206)) xor (layer2_outputs(4717)));
    outputs(4597) <= (layer2_outputs(2280)) or (layer2_outputs(894));
    outputs(4598) <= (layer2_outputs(9922)) and (layer2_outputs(3221));
    outputs(4599) <= not(layer2_outputs(2793));
    outputs(4600) <= (layer2_outputs(10119)) and not (layer2_outputs(1668));
    outputs(4601) <= layer2_outputs(600);
    outputs(4602) <= not(layer2_outputs(8501));
    outputs(4603) <= (layer2_outputs(4733)) xor (layer2_outputs(6222));
    outputs(4604) <= layer2_outputs(11978);
    outputs(4605) <= (layer2_outputs(11237)) and not (layer2_outputs(11062));
    outputs(4606) <= not((layer2_outputs(1309)) xor (layer2_outputs(4765)));
    outputs(4607) <= layer2_outputs(4814);
    outputs(4608) <= not((layer2_outputs(2515)) xor (layer2_outputs(6151)));
    outputs(4609) <= layer2_outputs(5163);
    outputs(4610) <= not((layer2_outputs(5626)) xor (layer2_outputs(9640)));
    outputs(4611) <= not(layer2_outputs(11568));
    outputs(4612) <= (layer2_outputs(4655)) and not (layer2_outputs(3515));
    outputs(4613) <= not(layer2_outputs(3583));
    outputs(4614) <= (layer2_outputs(9479)) xor (layer2_outputs(11932));
    outputs(4615) <= layer2_outputs(6859);
    outputs(4616) <= (layer2_outputs(2304)) xor (layer2_outputs(5824));
    outputs(4617) <= layer2_outputs(8649);
    outputs(4618) <= layer2_outputs(6945);
    outputs(4619) <= not((layer2_outputs(10395)) xor (layer2_outputs(810)));
    outputs(4620) <= (layer2_outputs(3663)) xor (layer2_outputs(7028));
    outputs(4621) <= not(layer2_outputs(5846));
    outputs(4622) <= not((layer2_outputs(5950)) xor (layer2_outputs(8201)));
    outputs(4623) <= (layer2_outputs(2092)) and not (layer2_outputs(3695));
    outputs(4624) <= layer2_outputs(495);
    outputs(4625) <= (layer2_outputs(4217)) xor (layer2_outputs(9192));
    outputs(4626) <= not((layer2_outputs(11073)) xor (layer2_outputs(4577)));
    outputs(4627) <= layer2_outputs(7449);
    outputs(4628) <= not(layer2_outputs(4449));
    outputs(4629) <= (layer2_outputs(10357)) xor (layer2_outputs(1182));
    outputs(4630) <= not((layer2_outputs(6691)) xor (layer2_outputs(1729)));
    outputs(4631) <= layer2_outputs(4310);
    outputs(4632) <= not((layer2_outputs(8646)) xor (layer2_outputs(756)));
    outputs(4633) <= not(layer2_outputs(1573));
    outputs(4634) <= not(layer2_outputs(1251)) or (layer2_outputs(3293));
    outputs(4635) <= (layer2_outputs(6005)) and not (layer2_outputs(11761));
    outputs(4636) <= not((layer2_outputs(6922)) xor (layer2_outputs(3271)));
    outputs(4637) <= not(layer2_outputs(2630));
    outputs(4638) <= not(layer2_outputs(7923));
    outputs(4639) <= not(layer2_outputs(4807));
    outputs(4640) <= layer2_outputs(4579);
    outputs(4641) <= not(layer2_outputs(7758));
    outputs(4642) <= not(layer2_outputs(11529));
    outputs(4643) <= layer2_outputs(12229);
    outputs(4644) <= not(layer2_outputs(11574));
    outputs(4645) <= not(layer2_outputs(2060));
    outputs(4646) <= (layer2_outputs(2756)) xor (layer2_outputs(7949));
    outputs(4647) <= layer2_outputs(11449);
    outputs(4648) <= layer2_outputs(9784);
    outputs(4649) <= not((layer2_outputs(4542)) or (layer2_outputs(10691)));
    outputs(4650) <= not((layer2_outputs(4210)) xor (layer2_outputs(8414)));
    outputs(4651) <= not((layer2_outputs(4451)) or (layer2_outputs(4159)));
    outputs(4652) <= not(layer2_outputs(10135)) or (layer2_outputs(12732));
    outputs(4653) <= not((layer2_outputs(7832)) xor (layer2_outputs(11464)));
    outputs(4654) <= not(layer2_outputs(5795));
    outputs(4655) <= layer2_outputs(2233);
    outputs(4656) <= layer2_outputs(8590);
    outputs(4657) <= layer2_outputs(7623);
    outputs(4658) <= not(layer2_outputs(4200));
    outputs(4659) <= not(layer2_outputs(1945));
    outputs(4660) <= not((layer2_outputs(4475)) xor (layer2_outputs(7854)));
    outputs(4661) <= not(layer2_outputs(12048)) or (layer2_outputs(9123));
    outputs(4662) <= layer2_outputs(6028);
    outputs(4663) <= not((layer2_outputs(11900)) xor (layer2_outputs(7685)));
    outputs(4664) <= layer2_outputs(9073);
    outputs(4665) <= layer2_outputs(6733);
    outputs(4666) <= not(layer2_outputs(10314));
    outputs(4667) <= not(layer2_outputs(9085));
    outputs(4668) <= not((layer2_outputs(6230)) xor (layer2_outputs(4999)));
    outputs(4669) <= (layer2_outputs(5036)) xor (layer2_outputs(3334));
    outputs(4670) <= (layer2_outputs(5564)) or (layer2_outputs(7033));
    outputs(4671) <= layer2_outputs(5372);
    outputs(4672) <= not(layer2_outputs(11707));
    outputs(4673) <= layer2_outputs(11297);
    outputs(4674) <= not((layer2_outputs(9348)) xor (layer2_outputs(7175)));
    outputs(4675) <= not((layer2_outputs(10433)) xor (layer2_outputs(11796)));
    outputs(4676) <= not(layer2_outputs(2074));
    outputs(4677) <= (layer2_outputs(12370)) xor (layer2_outputs(11116));
    outputs(4678) <= (layer2_outputs(10539)) xor (layer2_outputs(145));
    outputs(4679) <= not(layer2_outputs(2436)) or (layer2_outputs(10561));
    outputs(4680) <= layer2_outputs(10004);
    outputs(4681) <= not((layer2_outputs(12780)) xor (layer2_outputs(2307)));
    outputs(4682) <= not(layer2_outputs(2469)) or (layer2_outputs(10491));
    outputs(4683) <= layer2_outputs(4553);
    outputs(4684) <= not(layer2_outputs(9742)) or (layer2_outputs(3964));
    outputs(4685) <= (layer2_outputs(1034)) xor (layer2_outputs(7107));
    outputs(4686) <= (layer2_outputs(2988)) and not (layer2_outputs(6607));
    outputs(4687) <= not(layer2_outputs(4830));
    outputs(4688) <= not(layer2_outputs(7811));
    outputs(4689) <= not(layer2_outputs(3069)) or (layer2_outputs(10888));
    outputs(4690) <= not(layer2_outputs(8836));
    outputs(4691) <= (layer2_outputs(4500)) xor (layer2_outputs(9391));
    outputs(4692) <= not(layer2_outputs(2952)) or (layer2_outputs(4435));
    outputs(4693) <= not(layer2_outputs(6357)) or (layer2_outputs(12635));
    outputs(4694) <= not(layer2_outputs(3585));
    outputs(4695) <= not(layer2_outputs(5490));
    outputs(4696) <= (layer2_outputs(1491)) xor (layer2_outputs(11813));
    outputs(4697) <= not(layer2_outputs(10947));
    outputs(4698) <= layer2_outputs(8330);
    outputs(4699) <= not(layer2_outputs(10528));
    outputs(4700) <= not((layer2_outputs(1818)) xor (layer2_outputs(4789)));
    outputs(4701) <= not((layer2_outputs(425)) xor (layer2_outputs(11634)));
    outputs(4702) <= (layer2_outputs(12646)) and not (layer2_outputs(7621));
    outputs(4703) <= layer2_outputs(3483);
    outputs(4704) <= not(layer2_outputs(8011));
    outputs(4705) <= not(layer2_outputs(3965));
    outputs(4706) <= layer2_outputs(4795);
    outputs(4707) <= not(layer2_outputs(2169));
    outputs(4708) <= layer2_outputs(10949);
    outputs(4709) <= layer2_outputs(5222);
    outputs(4710) <= layer2_outputs(10596);
    outputs(4711) <= not(layer2_outputs(5963));
    outputs(4712) <= layer2_outputs(4256);
    outputs(4713) <= not((layer2_outputs(3886)) xor (layer2_outputs(9583)));
    outputs(4714) <= layer2_outputs(6396);
    outputs(4715) <= not(layer2_outputs(10225));
    outputs(4716) <= layer2_outputs(1021);
    outputs(4717) <= not((layer2_outputs(7492)) xor (layer2_outputs(9229)));
    outputs(4718) <= not(layer2_outputs(10644));
    outputs(4719) <= not(layer2_outputs(1542));
    outputs(4720) <= not(layer2_outputs(4948));
    outputs(4721) <= (layer2_outputs(188)) and not (layer2_outputs(4023));
    outputs(4722) <= not(layer2_outputs(9579)) or (layer2_outputs(3074));
    outputs(4723) <= layer2_outputs(9332);
    outputs(4724) <= not(layer2_outputs(11353)) or (layer2_outputs(3297));
    outputs(4725) <= not(layer2_outputs(8257));
    outputs(4726) <= not(layer2_outputs(5664)) or (layer2_outputs(4925));
    outputs(4727) <= (layer2_outputs(1958)) xor (layer2_outputs(7378));
    outputs(4728) <= not((layer2_outputs(11817)) xor (layer2_outputs(1055)));
    outputs(4729) <= (layer2_outputs(2724)) and not (layer2_outputs(4433));
    outputs(4730) <= not(layer2_outputs(4953));
    outputs(4731) <= (layer2_outputs(8677)) and (layer2_outputs(96));
    outputs(4732) <= not(layer2_outputs(5594));
    outputs(4733) <= not((layer2_outputs(540)) xor (layer2_outputs(9461)));
    outputs(4734) <= layer2_outputs(327);
    outputs(4735) <= layer2_outputs(674);
    outputs(4736) <= layer2_outputs(5557);
    outputs(4737) <= not(layer2_outputs(3854));
    outputs(4738) <= layer2_outputs(10753);
    outputs(4739) <= not(layer2_outputs(6061));
    outputs(4740) <= layer2_outputs(2786);
    outputs(4741) <= layer2_outputs(12253);
    outputs(4742) <= not((layer2_outputs(6507)) xor (layer2_outputs(7207)));
    outputs(4743) <= layer2_outputs(1100);
    outputs(4744) <= not((layer2_outputs(7909)) xor (layer2_outputs(11114)));
    outputs(4745) <= not(layer2_outputs(4198)) or (layer2_outputs(1478));
    outputs(4746) <= layer2_outputs(981);
    outputs(4747) <= (layer2_outputs(3116)) xor (layer2_outputs(4307));
    outputs(4748) <= not(layer2_outputs(2618));
    outputs(4749) <= (layer2_outputs(1208)) xor (layer2_outputs(722));
    outputs(4750) <= (layer2_outputs(8266)) xor (layer2_outputs(3642));
    outputs(4751) <= (layer2_outputs(4038)) and not (layer2_outputs(11100));
    outputs(4752) <= not((layer2_outputs(4503)) xor (layer2_outputs(1173)));
    outputs(4753) <= not(layer2_outputs(1151)) or (layer2_outputs(1960));
    outputs(4754) <= layer2_outputs(12786);
    outputs(4755) <= layer2_outputs(12755);
    outputs(4756) <= not((layer2_outputs(9693)) xor (layer2_outputs(10432)));
    outputs(4757) <= not(layer2_outputs(11975));
    outputs(4758) <= not(layer2_outputs(7958));
    outputs(4759) <= layer2_outputs(1822);
    outputs(4760) <= layer2_outputs(3434);
    outputs(4761) <= (layer2_outputs(10906)) and not (layer2_outputs(3087));
    outputs(4762) <= not(layer2_outputs(5307));
    outputs(4763) <= not(layer2_outputs(5838));
    outputs(4764) <= not((layer2_outputs(9956)) xor (layer2_outputs(557)));
    outputs(4765) <= (layer2_outputs(5518)) and (layer2_outputs(11963));
    outputs(4766) <= layer2_outputs(3175);
    outputs(4767) <= not(layer2_outputs(3515));
    outputs(4768) <= not(layer2_outputs(8056));
    outputs(4769) <= not((layer2_outputs(12790)) and (layer2_outputs(473)));
    outputs(4770) <= not((layer2_outputs(8642)) xor (layer2_outputs(7778)));
    outputs(4771) <= layer2_outputs(2525);
    outputs(4772) <= layer2_outputs(7633);
    outputs(4773) <= (layer2_outputs(4279)) xor (layer2_outputs(12359));
    outputs(4774) <= layer2_outputs(6914);
    outputs(4775) <= not((layer2_outputs(1371)) xor (layer2_outputs(4735)));
    outputs(4776) <= layer2_outputs(5707);
    outputs(4777) <= layer2_outputs(8252);
    outputs(4778) <= not((layer2_outputs(4532)) xor (layer2_outputs(8808)));
    outputs(4779) <= not(layer2_outputs(7381));
    outputs(4780) <= not(layer2_outputs(8858));
    outputs(4781) <= layer2_outputs(8054);
    outputs(4782) <= (layer2_outputs(10715)) and (layer2_outputs(6102));
    outputs(4783) <= not(layer2_outputs(5380));
    outputs(4784) <= (layer2_outputs(11486)) and not (layer2_outputs(5746));
    outputs(4785) <= (layer2_outputs(8161)) xor (layer2_outputs(9230));
    outputs(4786) <= layer2_outputs(10326);
    outputs(4787) <= layer2_outputs(9225);
    outputs(4788) <= not(layer2_outputs(12348));
    outputs(4789) <= layer2_outputs(4821);
    outputs(4790) <= (layer2_outputs(5445)) xor (layer2_outputs(1181));
    outputs(4791) <= not(layer2_outputs(3854));
    outputs(4792) <= (layer2_outputs(4749)) and (layer2_outputs(10804));
    outputs(4793) <= not(layer2_outputs(5192));
    outputs(4794) <= not((layer2_outputs(12222)) and (layer2_outputs(7654)));
    outputs(4795) <= not((layer2_outputs(1647)) xor (layer2_outputs(1755)));
    outputs(4796) <= layer2_outputs(4205);
    outputs(4797) <= not(layer2_outputs(6051));
    outputs(4798) <= (layer2_outputs(10208)) xor (layer2_outputs(3475));
    outputs(4799) <= layer2_outputs(10971);
    outputs(4800) <= (layer2_outputs(9072)) xor (layer2_outputs(162));
    outputs(4801) <= layer2_outputs(7873);
    outputs(4802) <= layer2_outputs(12675);
    outputs(4803) <= not(layer2_outputs(6282));
    outputs(4804) <= layer2_outputs(11937);
    outputs(4805) <= layer2_outputs(6329);
    outputs(4806) <= not((layer2_outputs(10834)) xor (layer2_outputs(7264)));
    outputs(4807) <= not(layer2_outputs(7265));
    outputs(4808) <= layer2_outputs(5320);
    outputs(4809) <= (layer2_outputs(11443)) xor (layer2_outputs(11907));
    outputs(4810) <= (layer2_outputs(11468)) xor (layer2_outputs(2908));
    outputs(4811) <= not((layer2_outputs(12667)) xor (layer2_outputs(11522)));
    outputs(4812) <= (layer2_outputs(8118)) and (layer2_outputs(12220));
    outputs(4813) <= layer2_outputs(6182);
    outputs(4814) <= layer2_outputs(10068);
    outputs(4815) <= layer2_outputs(1886);
    outputs(4816) <= (layer2_outputs(9921)) and not (layer2_outputs(118));
    outputs(4817) <= not(layer2_outputs(7279));
    outputs(4818) <= layer2_outputs(8463);
    outputs(4819) <= (layer2_outputs(1557)) xor (layer2_outputs(4756));
    outputs(4820) <= (layer2_outputs(9449)) xor (layer2_outputs(9516));
    outputs(4821) <= not((layer2_outputs(286)) or (layer2_outputs(6127)));
    outputs(4822) <= not(layer2_outputs(1436));
    outputs(4823) <= layer2_outputs(2451);
    outputs(4824) <= (layer2_outputs(11843)) xor (layer2_outputs(2925));
    outputs(4825) <= not(layer2_outputs(11724)) or (layer2_outputs(2220));
    outputs(4826) <= layer2_outputs(5968);
    outputs(4827) <= layer2_outputs(12679);
    outputs(4828) <= not(layer2_outputs(3327));
    outputs(4829) <= layer2_outputs(11756);
    outputs(4830) <= not(layer2_outputs(9381));
    outputs(4831) <= layer2_outputs(5412);
    outputs(4832) <= not(layer2_outputs(1857));
    outputs(4833) <= layer2_outputs(3157);
    outputs(4834) <= layer2_outputs(5495);
    outputs(4835) <= not((layer2_outputs(7244)) or (layer2_outputs(7783)));
    outputs(4836) <= (layer2_outputs(543)) and (layer2_outputs(5528));
    outputs(4837) <= not((layer2_outputs(11895)) xor (layer2_outputs(5788)));
    outputs(4838) <= (layer2_outputs(5255)) or (layer2_outputs(2983));
    outputs(4839) <= layer2_outputs(4349);
    outputs(4840) <= layer2_outputs(5924);
    outputs(4841) <= layer2_outputs(2025);
    outputs(4842) <= not(layer2_outputs(2612));
    outputs(4843) <= not((layer2_outputs(4118)) and (layer2_outputs(8581)));
    outputs(4844) <= (layer2_outputs(2442)) and (layer2_outputs(2333));
    outputs(4845) <= not((layer2_outputs(1985)) or (layer2_outputs(300)));
    outputs(4846) <= not(layer2_outputs(2071));
    outputs(4847) <= (layer2_outputs(9736)) xor (layer2_outputs(4397));
    outputs(4848) <= (layer2_outputs(8416)) xor (layer2_outputs(9471));
    outputs(4849) <= not(layer2_outputs(11335));
    outputs(4850) <= not((layer2_outputs(2863)) xor (layer2_outputs(6112)));
    outputs(4851) <= layer2_outputs(1617);
    outputs(4852) <= not(layer2_outputs(10154));
    outputs(4853) <= not((layer2_outputs(11710)) and (layer2_outputs(2432)));
    outputs(4854) <= layer2_outputs(8737);
    outputs(4855) <= not((layer2_outputs(5400)) xor (layer2_outputs(10309)));
    outputs(4856) <= layer2_outputs(5058);
    outputs(4857) <= not(layer2_outputs(9563));
    outputs(4858) <= (layer2_outputs(7697)) and (layer2_outputs(7420));
    outputs(4859) <= not(layer2_outputs(8660)) or (layer2_outputs(4842));
    outputs(4860) <= (layer2_outputs(3273)) xor (layer2_outputs(338));
    outputs(4861) <= not(layer2_outputs(2088));
    outputs(4862) <= (layer2_outputs(9693)) or (layer2_outputs(7180));
    outputs(4863) <= (layer2_outputs(668)) xor (layer2_outputs(10686));
    outputs(4864) <= layer2_outputs(2308);
    outputs(4865) <= layer2_outputs(10751);
    outputs(4866) <= not((layer2_outputs(4203)) xor (layer2_outputs(3944)));
    outputs(4867) <= (layer2_outputs(11408)) or (layer2_outputs(11140));
    outputs(4868) <= layer2_outputs(11281);
    outputs(4869) <= layer2_outputs(6682);
    outputs(4870) <= not(layer2_outputs(7737));
    outputs(4871) <= layer2_outputs(9643);
    outputs(4872) <= not(layer2_outputs(6638));
    outputs(4873) <= layer2_outputs(3768);
    outputs(4874) <= not(layer2_outputs(4177));
    outputs(4875) <= not((layer2_outputs(4642)) xor (layer2_outputs(841)));
    outputs(4876) <= layer2_outputs(4586);
    outputs(4877) <= not(layer2_outputs(6640));
    outputs(4878) <= not((layer2_outputs(9546)) xor (layer2_outputs(7603)));
    outputs(4879) <= (layer2_outputs(9465)) xor (layer2_outputs(5287));
    outputs(4880) <= not((layer2_outputs(10834)) and (layer2_outputs(10629)));
    outputs(4881) <= not(layer2_outputs(12439)) or (layer2_outputs(10004));
    outputs(4882) <= not(layer2_outputs(8447));
    outputs(4883) <= (layer2_outputs(5801)) and not (layer2_outputs(12257));
    outputs(4884) <= not((layer2_outputs(5523)) xor (layer2_outputs(7560)));
    outputs(4885) <= not(layer2_outputs(795));
    outputs(4886) <= (layer2_outputs(6741)) xor (layer2_outputs(1119));
    outputs(4887) <= (layer2_outputs(7532)) or (layer2_outputs(4515));
    outputs(4888) <= not(layer2_outputs(779));
    outputs(4889) <= not(layer2_outputs(6463));
    outputs(4890) <= (layer2_outputs(9794)) and not (layer2_outputs(11453));
    outputs(4891) <= layer2_outputs(11642);
    outputs(4892) <= not(layer2_outputs(5926)) or (layer2_outputs(10047));
    outputs(4893) <= not(layer2_outputs(6065));
    outputs(4894) <= not((layer2_outputs(8638)) xor (layer2_outputs(7965)));
    outputs(4895) <= not(layer2_outputs(2387));
    outputs(4896) <= layer2_outputs(220);
    outputs(4897) <= not(layer2_outputs(6875));
    outputs(4898) <= layer2_outputs(6);
    outputs(4899) <= (layer2_outputs(5821)) xor (layer2_outputs(6998));
    outputs(4900) <= layer2_outputs(8280);
    outputs(4901) <= layer2_outputs(5528);
    outputs(4902) <= (layer2_outputs(5919)) xor (layer2_outputs(12186));
    outputs(4903) <= layer2_outputs(9368);
    outputs(4904) <= layer2_outputs(2978);
    outputs(4905) <= not(layer2_outputs(1089));
    outputs(4906) <= (layer2_outputs(5788)) xor (layer2_outputs(3444));
    outputs(4907) <= not((layer2_outputs(12517)) and (layer2_outputs(5180)));
    outputs(4908) <= layer2_outputs(9884);
    outputs(4909) <= layer2_outputs(4234);
    outputs(4910) <= not((layer2_outputs(2976)) xor (layer2_outputs(6304)));
    outputs(4911) <= layer2_outputs(1199);
    outputs(4912) <= not(layer2_outputs(12335));
    outputs(4913) <= (layer2_outputs(949)) or (layer2_outputs(4411));
    outputs(4914) <= (layer2_outputs(3064)) or (layer2_outputs(7495));
    outputs(4915) <= (layer2_outputs(5454)) and (layer2_outputs(5234));
    outputs(4916) <= not(layer2_outputs(1460));
    outputs(4917) <= layer2_outputs(5197);
    outputs(4918) <= not((layer2_outputs(4675)) xor (layer2_outputs(2593)));
    outputs(4919) <= not(layer2_outputs(5467));
    outputs(4920) <= (layer2_outputs(26)) xor (layer2_outputs(1837));
    outputs(4921) <= (layer2_outputs(1032)) and (layer2_outputs(2692));
    outputs(4922) <= not(layer2_outputs(9688)) or (layer2_outputs(10169));
    outputs(4923) <= (layer2_outputs(4282)) xor (layer2_outputs(7042));
    outputs(4924) <= (layer2_outputs(2374)) and not (layer2_outputs(12402));
    outputs(4925) <= not((layer2_outputs(12573)) xor (layer2_outputs(10017)));
    outputs(4926) <= not(layer2_outputs(11646));
    outputs(4927) <= (layer2_outputs(2602)) and not (layer2_outputs(2665));
    outputs(4928) <= not(layer2_outputs(5204));
    outputs(4929) <= layer2_outputs(4626);
    outputs(4930) <= layer2_outputs(9631);
    outputs(4931) <= (layer2_outputs(11413)) and (layer2_outputs(1283));
    outputs(4932) <= (layer2_outputs(66)) and not (layer2_outputs(9567));
    outputs(4933) <= (layer2_outputs(8675)) xor (layer2_outputs(7268));
    outputs(4934) <= layer2_outputs(5125);
    outputs(4935) <= not(layer2_outputs(8706));
    outputs(4936) <= (layer2_outputs(1267)) xor (layer2_outputs(816));
    outputs(4937) <= layer2_outputs(11881);
    outputs(4938) <= not(layer2_outputs(651)) or (layer2_outputs(2));
    outputs(4939) <= not(layer2_outputs(8807));
    outputs(4940) <= (layer2_outputs(4218)) xor (layer2_outputs(2528));
    outputs(4941) <= (layer2_outputs(432)) xor (layer2_outputs(4978));
    outputs(4942) <= not((layer2_outputs(1819)) xor (layer2_outputs(6889)));
    outputs(4943) <= not((layer2_outputs(12779)) xor (layer2_outputs(10781)));
    outputs(4944) <= layer2_outputs(11324);
    outputs(4945) <= not(layer2_outputs(11346));
    outputs(4946) <= layer2_outputs(9139);
    outputs(4947) <= layer2_outputs(12756);
    outputs(4948) <= layer2_outputs(4057);
    outputs(4949) <= (layer2_outputs(5636)) xor (layer2_outputs(1704));
    outputs(4950) <= layer2_outputs(10649);
    outputs(4951) <= not((layer2_outputs(7072)) and (layer2_outputs(7576)));
    outputs(4952) <= not(layer2_outputs(6901));
    outputs(4953) <= not(layer2_outputs(3687));
    outputs(4954) <= not(layer2_outputs(3720));
    outputs(4955) <= layer2_outputs(430);
    outputs(4956) <= layer2_outputs(6217);
    outputs(4957) <= (layer2_outputs(5346)) xor (layer2_outputs(12057));
    outputs(4958) <= not((layer2_outputs(11076)) and (layer2_outputs(9462)));
    outputs(4959) <= (layer2_outputs(4672)) and not (layer2_outputs(3733));
    outputs(4960) <= (layer2_outputs(8952)) xor (layer2_outputs(10892));
    outputs(4961) <= not(layer2_outputs(12290));
    outputs(4962) <= (layer2_outputs(3035)) and not (layer2_outputs(7726));
    outputs(4963) <= (layer2_outputs(2052)) and not (layer2_outputs(6670));
    outputs(4964) <= not(layer2_outputs(1245));
    outputs(4965) <= not((layer2_outputs(7414)) xor (layer2_outputs(10945)));
    outputs(4966) <= not(layer2_outputs(7102));
    outputs(4967) <= not(layer2_outputs(2989));
    outputs(4968) <= not(layer2_outputs(8226));
    outputs(4969) <= (layer2_outputs(8019)) xor (layer2_outputs(551));
    outputs(4970) <= not(layer2_outputs(421));
    outputs(4971) <= not(layer2_outputs(8986)) or (layer2_outputs(5663));
    outputs(4972) <= layer2_outputs(1333);
    outputs(4973) <= not((layer2_outputs(7759)) or (layer2_outputs(6071)));
    outputs(4974) <= not(layer2_outputs(11562));
    outputs(4975) <= (layer2_outputs(1387)) and not (layer2_outputs(12628));
    outputs(4976) <= (layer2_outputs(4845)) and not (layer2_outputs(407));
    outputs(4977) <= layer2_outputs(5338);
    outputs(4978) <= layer2_outputs(6423);
    outputs(4979) <= (layer2_outputs(5134)) and (layer2_outputs(7487));
    outputs(4980) <= not(layer2_outputs(10716));
    outputs(4981) <= layer2_outputs(792);
    outputs(4982) <= not((layer2_outputs(7826)) xor (layer2_outputs(2347)));
    outputs(4983) <= layer2_outputs(4027);
    outputs(4984) <= not((layer2_outputs(772)) or (layer2_outputs(10513)));
    outputs(4985) <= not((layer2_outputs(359)) or (layer2_outputs(6224)));
    outputs(4986) <= (layer2_outputs(5943)) xor (layer2_outputs(12543));
    outputs(4987) <= not(layer2_outputs(7509));
    outputs(4988) <= layer2_outputs(3367);
    outputs(4989) <= layer2_outputs(11971);
    outputs(4990) <= not(layer2_outputs(268)) or (layer2_outputs(9021));
    outputs(4991) <= not(layer2_outputs(9376));
    outputs(4992) <= layer2_outputs(8810);
    outputs(4993) <= not(layer2_outputs(3802));
    outputs(4994) <= layer2_outputs(2980);
    outputs(4995) <= layer2_outputs(5506);
    outputs(4996) <= layer2_outputs(2544);
    outputs(4997) <= layer2_outputs(3440);
    outputs(4998) <= not((layer2_outputs(10497)) xor (layer2_outputs(199)));
    outputs(4999) <= not(layer2_outputs(3453));
    outputs(5000) <= (layer2_outputs(1236)) and not (layer2_outputs(11550));
    outputs(5001) <= layer2_outputs(3132);
    outputs(5002) <= not((layer2_outputs(12761)) or (layer2_outputs(7256)));
    outputs(5003) <= (layer2_outputs(149)) xor (layer2_outputs(2311));
    outputs(5004) <= not(layer2_outputs(9697)) or (layer2_outputs(12720));
    outputs(5005) <= layer2_outputs(8417);
    outputs(5006) <= layer2_outputs(3017);
    outputs(5007) <= layer2_outputs(4150);
    outputs(5008) <= layer2_outputs(12273);
    outputs(5009) <= (layer2_outputs(201)) xor (layer2_outputs(5746));
    outputs(5010) <= not((layer2_outputs(9772)) xor (layer2_outputs(5908)));
    outputs(5011) <= (layer2_outputs(4480)) xor (layer2_outputs(8288));
    outputs(5012) <= layer2_outputs(6104);
    outputs(5013) <= layer2_outputs(10382);
    outputs(5014) <= not((layer2_outputs(857)) xor (layer2_outputs(10235)));
    outputs(5015) <= not(layer2_outputs(905));
    outputs(5016) <= not(layer2_outputs(6082));
    outputs(5017) <= (layer2_outputs(10623)) and not (layer2_outputs(5204));
    outputs(5018) <= not(layer2_outputs(727));
    outputs(5019) <= (layer2_outputs(1677)) xor (layer2_outputs(5427));
    outputs(5020) <= (layer2_outputs(7548)) and not (layer2_outputs(5516));
    outputs(5021) <= (layer2_outputs(7277)) xor (layer2_outputs(3540));
    outputs(5022) <= (layer2_outputs(265)) and (layer2_outputs(3391));
    outputs(5023) <= layer2_outputs(5584);
    outputs(5024) <= not(layer2_outputs(3792));
    outputs(5025) <= not((layer2_outputs(12164)) or (layer2_outputs(881)));
    outputs(5026) <= (layer2_outputs(11051)) xor (layer2_outputs(455));
    outputs(5027) <= layer2_outputs(1250);
    outputs(5028) <= not(layer2_outputs(9489));
    outputs(5029) <= not(layer2_outputs(2083));
    outputs(5030) <= (layer2_outputs(9040)) xor (layer2_outputs(8378));
    outputs(5031) <= (layer2_outputs(11522)) xor (layer2_outputs(2234));
    outputs(5032) <= (layer2_outputs(254)) xor (layer2_outputs(7510));
    outputs(5033) <= layer2_outputs(10646);
    outputs(5034) <= layer2_outputs(9239);
    outputs(5035) <= layer2_outputs(1480);
    outputs(5036) <= (layer2_outputs(6385)) and not (layer2_outputs(5096));
    outputs(5037) <= not(layer2_outputs(12233));
    outputs(5038) <= layer2_outputs(612);
    outputs(5039) <= layer2_outputs(12268);
    outputs(5040) <= (layer2_outputs(4014)) xor (layer2_outputs(7972));
    outputs(5041) <= layer2_outputs(8507);
    outputs(5042) <= (layer2_outputs(7407)) and not (layer2_outputs(5470));
    outputs(5043) <= layer2_outputs(10983);
    outputs(5044) <= (layer2_outputs(12298)) xor (layer2_outputs(7498));
    outputs(5045) <= not(layer2_outputs(1876));
    outputs(5046) <= (layer2_outputs(7766)) and not (layer2_outputs(7280));
    outputs(5047) <= not((layer2_outputs(5022)) xor (layer2_outputs(3698)));
    outputs(5048) <= not(layer2_outputs(7385));
    outputs(5049) <= layer2_outputs(5596);
    outputs(5050) <= not(layer2_outputs(1901));
    outputs(5051) <= layer2_outputs(12053);
    outputs(5052) <= layer2_outputs(7402);
    outputs(5053) <= (layer2_outputs(11985)) or (layer2_outputs(3710));
    outputs(5054) <= not(layer2_outputs(9096));
    outputs(5055) <= not((layer2_outputs(7152)) xor (layer2_outputs(9888)));
    outputs(5056) <= not(layer2_outputs(10534));
    outputs(5057) <= not((layer2_outputs(9082)) or (layer2_outputs(2909)));
    outputs(5058) <= layer2_outputs(8810);
    outputs(5059) <= layer2_outputs(4079);
    outputs(5060) <= layer2_outputs(10253);
    outputs(5061) <= layer2_outputs(10447);
    outputs(5062) <= (layer2_outputs(9813)) xor (layer2_outputs(1166));
    outputs(5063) <= not((layer2_outputs(12340)) or (layer2_outputs(6512)));
    outputs(5064) <= layer2_outputs(9855);
    outputs(5065) <= not(layer2_outputs(8332));
    outputs(5066) <= layer2_outputs(10745);
    outputs(5067) <= layer2_outputs(2984);
    outputs(5068) <= layer2_outputs(8398);
    outputs(5069) <= layer2_outputs(6336);
    outputs(5070) <= layer2_outputs(10714);
    outputs(5071) <= not(layer2_outputs(12080));
    outputs(5072) <= layer2_outputs(4602);
    outputs(5073) <= not(layer2_outputs(9090));
    outputs(5074) <= not(layer2_outputs(5430));
    outputs(5075) <= not((layer2_outputs(7772)) xor (layer2_outputs(1529)));
    outputs(5076) <= layer2_outputs(10340);
    outputs(5077) <= not(layer2_outputs(12309));
    outputs(5078) <= (layer2_outputs(12019)) xor (layer2_outputs(3612));
    outputs(5079) <= layer2_outputs(10199);
    outputs(5080) <= (layer2_outputs(7031)) and (layer2_outputs(2649));
    outputs(5081) <= not(layer2_outputs(250));
    outputs(5082) <= not(layer2_outputs(9136));
    outputs(5083) <= (layer2_outputs(8642)) and (layer2_outputs(7352));
    outputs(5084) <= layer2_outputs(201);
    outputs(5085) <= (layer2_outputs(2149)) xor (layer2_outputs(2591));
    outputs(5086) <= not((layer2_outputs(3155)) xor (layer2_outputs(5241)));
    outputs(5087) <= not(layer2_outputs(579));
    outputs(5088) <= (layer2_outputs(11316)) and not (layer2_outputs(5896));
    outputs(5089) <= not((layer2_outputs(3682)) xor (layer2_outputs(7779)));
    outputs(5090) <= not(layer2_outputs(9307));
    outputs(5091) <= (layer2_outputs(11983)) xor (layer2_outputs(11273));
    outputs(5092) <= not(layer2_outputs(12346));
    outputs(5093) <= layer2_outputs(11666);
    outputs(5094) <= not(layer2_outputs(8163));
    outputs(5095) <= (layer2_outputs(2133)) and not (layer2_outputs(8662));
    outputs(5096) <= not((layer2_outputs(8174)) xor (layer2_outputs(11980)));
    outputs(5097) <= (layer2_outputs(2087)) and not (layer2_outputs(9781));
    outputs(5098) <= not(layer2_outputs(9217));
    outputs(5099) <= layer2_outputs(1713);
    outputs(5100) <= not(layer2_outputs(11967)) or (layer2_outputs(7790));
    outputs(5101) <= not(layer2_outputs(3488));
    outputs(5102) <= layer2_outputs(7160);
    outputs(5103) <= (layer2_outputs(3433)) xor (layer2_outputs(1159));
    outputs(5104) <= layer2_outputs(6328);
    outputs(5105) <= (layer2_outputs(7081)) xor (layer2_outputs(7835));
    outputs(5106) <= not(layer2_outputs(9035));
    outputs(5107) <= not(layer2_outputs(10091));
    outputs(5108) <= not((layer2_outputs(12360)) xor (layer2_outputs(8892)));
    outputs(5109) <= layer2_outputs(4828);
    outputs(5110) <= not((layer2_outputs(10057)) xor (layer2_outputs(6851)));
    outputs(5111) <= not(layer2_outputs(2664));
    outputs(5112) <= not(layer2_outputs(11773));
    outputs(5113) <= layer2_outputs(7009);
    outputs(5114) <= layer2_outputs(5831);
    outputs(5115) <= not(layer2_outputs(6616));
    outputs(5116) <= layer2_outputs(12723);
    outputs(5117) <= not(layer2_outputs(204));
    outputs(5118) <= not(layer2_outputs(3134));
    outputs(5119) <= (layer2_outputs(6508)) xor (layer2_outputs(8545));
    outputs(5120) <= not((layer2_outputs(12238)) or (layer2_outputs(8886)));
    outputs(5121) <= (layer2_outputs(6668)) xor (layer2_outputs(7295));
    outputs(5122) <= layer2_outputs(4767);
    outputs(5123) <= layer2_outputs(3229);
    outputs(5124) <= not(layer2_outputs(10517));
    outputs(5125) <= layer2_outputs(10225);
    outputs(5126) <= layer2_outputs(1033);
    outputs(5127) <= not(layer2_outputs(261));
    outputs(5128) <= not(layer2_outputs(5061));
    outputs(5129) <= not(layer2_outputs(3113));
    outputs(5130) <= not((layer2_outputs(4152)) xor (layer2_outputs(3958)));
    outputs(5131) <= (layer2_outputs(8924)) or (layer2_outputs(1072));
    outputs(5132) <= (layer2_outputs(10943)) xor (layer2_outputs(6265));
    outputs(5133) <= not(layer2_outputs(1368));
    outputs(5134) <= (layer2_outputs(6276)) xor (layer2_outputs(6520));
    outputs(5135) <= layer2_outputs(9749);
    outputs(5136) <= not(layer2_outputs(9149)) or (layer2_outputs(6490));
    outputs(5137) <= (layer2_outputs(8058)) xor (layer2_outputs(3933));
    outputs(5138) <= not((layer2_outputs(9377)) xor (layer2_outputs(648)));
    outputs(5139) <= layer2_outputs(1750);
    outputs(5140) <= (layer2_outputs(3342)) xor (layer2_outputs(7097));
    outputs(5141) <= (layer2_outputs(5922)) xor (layer2_outputs(11401));
    outputs(5142) <= layer2_outputs(8633);
    outputs(5143) <= not((layer2_outputs(12531)) xor (layer2_outputs(4188)));
    outputs(5144) <= (layer2_outputs(6032)) and (layer2_outputs(11190));
    outputs(5145) <= (layer2_outputs(11511)) and not (layer2_outputs(11633));
    outputs(5146) <= layer2_outputs(12609);
    outputs(5147) <= layer2_outputs(6038);
    outputs(5148) <= (layer2_outputs(3546)) xor (layer2_outputs(3361));
    outputs(5149) <= not((layer2_outputs(694)) or (layer2_outputs(12269)));
    outputs(5150) <= not((layer2_outputs(4588)) xor (layer2_outputs(819)));
    outputs(5151) <= (layer2_outputs(3228)) xor (layer2_outputs(3624));
    outputs(5152) <= (layer2_outputs(12767)) xor (layer2_outputs(7320));
    outputs(5153) <= (layer2_outputs(11044)) xor (layer2_outputs(5044));
    outputs(5154) <= not(layer2_outputs(5890));
    outputs(5155) <= not(layer2_outputs(5699)) or (layer2_outputs(12765));
    outputs(5156) <= (layer2_outputs(11171)) xor (layer2_outputs(5093));
    outputs(5157) <= (layer2_outputs(5649)) xor (layer2_outputs(7640));
    outputs(5158) <= layer2_outputs(10855);
    outputs(5159) <= not((layer2_outputs(11201)) or (layer2_outputs(8312)));
    outputs(5160) <= not(layer2_outputs(850));
    outputs(5161) <= (layer2_outputs(10505)) xor (layer2_outputs(2624));
    outputs(5162) <= (layer2_outputs(12749)) xor (layer2_outputs(3829));
    outputs(5163) <= not(layer2_outputs(8453)) or (layer2_outputs(8361));
    outputs(5164) <= not(layer2_outputs(5440));
    outputs(5165) <= (layer2_outputs(1196)) xor (layer2_outputs(3573));
    outputs(5166) <= not((layer2_outputs(5081)) and (layer2_outputs(7046)));
    outputs(5167) <= not(layer2_outputs(517));
    outputs(5168) <= not((layer2_outputs(7702)) or (layer2_outputs(4884)));
    outputs(5169) <= not(layer2_outputs(4953));
    outputs(5170) <= layer2_outputs(474);
    outputs(5171) <= (layer2_outputs(8573)) xor (layer2_outputs(5194));
    outputs(5172) <= (layer2_outputs(5001)) xor (layer2_outputs(6592));
    outputs(5173) <= not(layer2_outputs(10477));
    outputs(5174) <= not(layer2_outputs(2138));
    outputs(5175) <= not((layer2_outputs(10833)) or (layer2_outputs(7695)));
    outputs(5176) <= layer2_outputs(10812);
    outputs(5177) <= not(layer2_outputs(7019));
    outputs(5178) <= not(layer2_outputs(6912));
    outputs(5179) <= not(layer2_outputs(7724));
    outputs(5180) <= layer2_outputs(5451);
    outputs(5181) <= layer2_outputs(2258);
    outputs(5182) <= (layer2_outputs(11211)) xor (layer2_outputs(5796));
    outputs(5183) <= (layer2_outputs(6936)) xor (layer2_outputs(10042));
    outputs(5184) <= layer2_outputs(10993);
    outputs(5185) <= not((layer2_outputs(9441)) xor (layer2_outputs(6031)));
    outputs(5186) <= not(layer2_outputs(3864));
    outputs(5187) <= (layer2_outputs(11696)) xor (layer2_outputs(3233));
    outputs(5188) <= layer2_outputs(12753);
    outputs(5189) <= not(layer2_outputs(3716));
    outputs(5190) <= layer2_outputs(6995);
    outputs(5191) <= (layer2_outputs(8619)) and (layer2_outputs(12598));
    outputs(5192) <= layer2_outputs(7701);
    outputs(5193) <= not(layer2_outputs(5156));
    outputs(5194) <= layer2_outputs(10022);
    outputs(5195) <= (layer2_outputs(3613)) xor (layer2_outputs(1961));
    outputs(5196) <= (layer2_outputs(5334)) xor (layer2_outputs(7592));
    outputs(5197) <= (layer2_outputs(757)) xor (layer2_outputs(2098));
    outputs(5198) <= not(layer2_outputs(4575));
    outputs(5199) <= not(layer2_outputs(5291));
    outputs(5200) <= not(layer2_outputs(1516));
    outputs(5201) <= not(layer2_outputs(510));
    outputs(5202) <= not(layer2_outputs(8419));
    outputs(5203) <= layer2_outputs(5778);
    outputs(5204) <= layer2_outputs(8943);
    outputs(5205) <= not(layer2_outputs(7568));
    outputs(5206) <= (layer2_outputs(12544)) xor (layer2_outputs(10274));
    outputs(5207) <= not(layer2_outputs(52));
    outputs(5208) <= not(layer2_outputs(602)) or (layer2_outputs(9686));
    outputs(5209) <= not(layer2_outputs(7137));
    outputs(5210) <= not(layer2_outputs(3754));
    outputs(5211) <= layer2_outputs(9101);
    outputs(5212) <= not(layer2_outputs(6447));
    outputs(5213) <= not(layer2_outputs(12038));
    outputs(5214) <= not((layer2_outputs(7246)) xor (layer2_outputs(3908)));
    outputs(5215) <= layer2_outputs(12454);
    outputs(5216) <= not((layer2_outputs(5330)) xor (layer2_outputs(1380)));
    outputs(5217) <= not(layer2_outputs(8173)) or (layer2_outputs(9456));
    outputs(5218) <= (layer2_outputs(5925)) xor (layer2_outputs(10598));
    outputs(5219) <= not(layer2_outputs(2702));
    outputs(5220) <= not(layer2_outputs(378));
    outputs(5221) <= layer2_outputs(946);
    outputs(5222) <= (layer2_outputs(7425)) or (layer2_outputs(10174));
    outputs(5223) <= not((layer2_outputs(7232)) xor (layer2_outputs(4271)));
    outputs(5224) <= layer2_outputs(3838);
    outputs(5225) <= layer2_outputs(8326);
    outputs(5226) <= not((layer2_outputs(11200)) xor (layer2_outputs(8546)));
    outputs(5227) <= not((layer2_outputs(1914)) xor (layer2_outputs(8304)));
    outputs(5228) <= layer2_outputs(7650);
    outputs(5229) <= not(layer2_outputs(4172));
    outputs(5230) <= layer2_outputs(12652);
    outputs(5231) <= layer2_outputs(7408);
    outputs(5232) <= not(layer2_outputs(12650));
    outputs(5233) <= not(layer2_outputs(3006));
    outputs(5234) <= not((layer2_outputs(8466)) and (layer2_outputs(1062)));
    outputs(5235) <= (layer2_outputs(7)) and not (layer2_outputs(10169));
    outputs(5236) <= (layer2_outputs(10721)) and not (layer2_outputs(319));
    outputs(5237) <= not((layer2_outputs(1019)) and (layer2_outputs(997)));
    outputs(5238) <= layer2_outputs(7249);
    outputs(5239) <= not((layer2_outputs(8015)) xor (layer2_outputs(6089)));
    outputs(5240) <= not((layer2_outputs(1554)) xor (layer2_outputs(8883)));
    outputs(5241) <= layer2_outputs(7957);
    outputs(5242) <= not(layer2_outputs(3861));
    outputs(5243) <= not(layer2_outputs(8920)) or (layer2_outputs(661));
    outputs(5244) <= layer2_outputs(3690);
    outputs(5245) <= not(layer2_outputs(4736)) or (layer2_outputs(3659));
    outputs(5246) <= not(layer2_outputs(10747));
    outputs(5247) <= layer2_outputs(7922);
    outputs(5248) <= not(layer2_outputs(1967));
    outputs(5249) <= not(layer2_outputs(8129)) or (layer2_outputs(7237));
    outputs(5250) <= (layer2_outputs(1633)) and (layer2_outputs(12459));
    outputs(5251) <= layer2_outputs(2499);
    outputs(5252) <= layer2_outputs(7927);
    outputs(5253) <= not(layer2_outputs(10746));
    outputs(5254) <= not(layer2_outputs(12440)) or (layer2_outputs(6728));
    outputs(5255) <= layer2_outputs(2398);
    outputs(5256) <= not((layer2_outputs(4025)) and (layer2_outputs(8467)));
    outputs(5257) <= layer2_outputs(116);
    outputs(5258) <= layer2_outputs(12235);
    outputs(5259) <= not(layer2_outputs(2473)) or (layer2_outputs(7370));
    outputs(5260) <= (layer2_outputs(10122)) or (layer2_outputs(5923));
    outputs(5261) <= layer2_outputs(2721);
    outputs(5262) <= not(layer2_outputs(9719));
    outputs(5263) <= not(layer2_outputs(8769));
    outputs(5264) <= not(layer2_outputs(11078));
    outputs(5265) <= layer2_outputs(9314);
    outputs(5266) <= not(layer2_outputs(11223)) or (layer2_outputs(724));
    outputs(5267) <= layer2_outputs(7409);
    outputs(5268) <= not(layer2_outputs(9016));
    outputs(5269) <= not((layer2_outputs(101)) xor (layer2_outputs(5058)));
    outputs(5270) <= (layer2_outputs(8516)) and (layer2_outputs(325));
    outputs(5271) <= not(layer2_outputs(6342));
    outputs(5272) <= not((layer2_outputs(12400)) xor (layer2_outputs(1495)));
    outputs(5273) <= layer2_outputs(376);
    outputs(5274) <= (layer2_outputs(4652)) xor (layer2_outputs(11584));
    outputs(5275) <= not(layer2_outputs(10312)) or (layer2_outputs(1785));
    outputs(5276) <= layer2_outputs(9545);
    outputs(5277) <= not(layer2_outputs(4342));
    outputs(5278) <= (layer2_outputs(4659)) or (layer2_outputs(10922));
    outputs(5279) <= not(layer2_outputs(7683)) or (layer2_outputs(8913));
    outputs(5280) <= not(layer2_outputs(9172));
    outputs(5281) <= (layer2_outputs(183)) xor (layer2_outputs(3179));
    outputs(5282) <= not(layer2_outputs(7638));
    outputs(5283) <= not((layer2_outputs(4557)) xor (layer2_outputs(8288)));
    outputs(5284) <= (layer2_outputs(6384)) xor (layer2_outputs(5931));
    outputs(5285) <= layer2_outputs(5764);
    outputs(5286) <= (layer2_outputs(6703)) and (layer2_outputs(7087));
    outputs(5287) <= not(layer2_outputs(8453));
    outputs(5288) <= (layer2_outputs(4470)) xor (layer2_outputs(6873));
    outputs(5289) <= not((layer2_outputs(7751)) xor (layer2_outputs(232)));
    outputs(5290) <= layer2_outputs(8439);
    outputs(5291) <= not(layer2_outputs(6294));
    outputs(5292) <= not((layer2_outputs(2957)) xor (layer2_outputs(3215)));
    outputs(5293) <= layer2_outputs(11130);
    outputs(5294) <= (layer2_outputs(11065)) xor (layer2_outputs(6225));
    outputs(5295) <= not(layer2_outputs(12752));
    outputs(5296) <= not(layer2_outputs(5008));
    outputs(5297) <= not(layer2_outputs(8813));
    outputs(5298) <= not(layer2_outputs(283));
    outputs(5299) <= not(layer2_outputs(7063));
    outputs(5300) <= not(layer2_outputs(3835));
    outputs(5301) <= not((layer2_outputs(8151)) xor (layer2_outputs(5760)));
    outputs(5302) <= not(layer2_outputs(3077));
    outputs(5303) <= layer2_outputs(10062);
    outputs(5304) <= layer2_outputs(1273);
    outputs(5305) <= (layer2_outputs(11012)) or (layer2_outputs(5068));
    outputs(5306) <= not((layer2_outputs(8035)) xor (layer2_outputs(1315)));
    outputs(5307) <= (layer2_outputs(11856)) xor (layer2_outputs(4924));
    outputs(5308) <= layer2_outputs(2290);
    outputs(5309) <= layer2_outputs(2664);
    outputs(5310) <= layer2_outputs(3653);
    outputs(5311) <= not((layer2_outputs(6425)) xor (layer2_outputs(7894)));
    outputs(5312) <= (layer2_outputs(1942)) and not (layer2_outputs(2143));
    outputs(5313) <= (layer2_outputs(11004)) xor (layer2_outputs(9313));
    outputs(5314) <= (layer2_outputs(4567)) and (layer2_outputs(11147));
    outputs(5315) <= not((layer2_outputs(1493)) or (layer2_outputs(548)));
    outputs(5316) <= layer2_outputs(10422);
    outputs(5317) <= layer2_outputs(11175);
    outputs(5318) <= layer2_outputs(4090);
    outputs(5319) <= not(layer2_outputs(8520));
    outputs(5320) <= layer2_outputs(718);
    outputs(5321) <= (layer2_outputs(8611)) and not (layer2_outputs(3840));
    outputs(5322) <= (layer2_outputs(10819)) xor (layer2_outputs(9965));
    outputs(5323) <= not(layer2_outputs(9696));
    outputs(5324) <= (layer2_outputs(4565)) xor (layer2_outputs(3571));
    outputs(5325) <= layer2_outputs(9627);
    outputs(5326) <= layer2_outputs(10978);
    outputs(5327) <= not(layer2_outputs(11547));
    outputs(5328) <= layer2_outputs(8634);
    outputs(5329) <= (layer2_outputs(6338)) xor (layer2_outputs(561));
    outputs(5330) <= not(layer2_outputs(4104));
    outputs(5331) <= not(layer2_outputs(645));
    outputs(5332) <= (layer2_outputs(1404)) xor (layer2_outputs(1620));
    outputs(5333) <= not((layer2_outputs(227)) xor (layer2_outputs(8825)));
    outputs(5334) <= (layer2_outputs(11414)) or (layer2_outputs(1334));
    outputs(5335) <= layer2_outputs(4897);
    outputs(5336) <= layer2_outputs(9629);
    outputs(5337) <= (layer2_outputs(5598)) and (layer2_outputs(7243));
    outputs(5338) <= layer2_outputs(10484);
    outputs(5339) <= (layer2_outputs(7756)) xor (layer2_outputs(1328));
    outputs(5340) <= not(layer2_outputs(10081));
    outputs(5341) <= (layer2_outputs(8632)) xor (layer2_outputs(2202));
    outputs(5342) <= layer2_outputs(5187);
    outputs(5343) <= not((layer2_outputs(2927)) xor (layer2_outputs(9345)));
    outputs(5344) <= not((layer2_outputs(8002)) or (layer2_outputs(2712)));
    outputs(5345) <= (layer2_outputs(3650)) and not (layer2_outputs(8133));
    outputs(5346) <= not(layer2_outputs(2220));
    outputs(5347) <= layer2_outputs(6438);
    outputs(5348) <= not((layer2_outputs(4730)) xor (layer2_outputs(2837)));
    outputs(5349) <= not(layer2_outputs(6305));
    outputs(5350) <= layer2_outputs(5989);
    outputs(5351) <= not(layer2_outputs(5699));
    outputs(5352) <= not(layer2_outputs(8859));
    outputs(5353) <= (layer2_outputs(1952)) and not (layer2_outputs(8000));
    outputs(5354) <= layer2_outputs(7906);
    outputs(5355) <= not(layer2_outputs(1326));
    outputs(5356) <= layer2_outputs(11378);
    outputs(5357) <= layer2_outputs(5730);
    outputs(5358) <= not(layer2_outputs(2384));
    outputs(5359) <= not(layer2_outputs(12602));
    outputs(5360) <= not(layer2_outputs(3333)) or (layer2_outputs(1469));
    outputs(5361) <= layer2_outputs(2382);
    outputs(5362) <= not(layer2_outputs(3317));
    outputs(5363) <= (layer2_outputs(11289)) xor (layer2_outputs(46));
    outputs(5364) <= not(layer2_outputs(1268));
    outputs(5365) <= not(layer2_outputs(9600)) or (layer2_outputs(8346));
    outputs(5366) <= not(layer2_outputs(8372));
    outputs(5367) <= (layer2_outputs(12506)) and not (layer2_outputs(191));
    outputs(5368) <= not((layer2_outputs(9331)) xor (layer2_outputs(7300)));
    outputs(5369) <= layer2_outputs(2358);
    outputs(5370) <= layer2_outputs(11111);
    outputs(5371) <= not(layer2_outputs(904));
    outputs(5372) <= not(layer2_outputs(3374));
    outputs(5373) <= not((layer2_outputs(9480)) xor (layer2_outputs(10167)));
    outputs(5374) <= not((layer2_outputs(2770)) xor (layer2_outputs(1059)));
    outputs(5375) <= (layer2_outputs(8805)) and not (layer2_outputs(9426));
    outputs(5376) <= not(layer2_outputs(5962));
    outputs(5377) <= not((layer2_outputs(7012)) or (layer2_outputs(5662)));
    outputs(5378) <= (layer2_outputs(885)) xor (layer2_outputs(5913));
    outputs(5379) <= (layer2_outputs(2987)) and (layer2_outputs(1070));
    outputs(5380) <= layer2_outputs(3082);
    outputs(5381) <= layer2_outputs(8190);
    outputs(5382) <= not(layer2_outputs(6110));
    outputs(5383) <= layer2_outputs(6137);
    outputs(5384) <= not(layer2_outputs(4357));
    outputs(5385) <= layer2_outputs(5632);
    outputs(5386) <= layer2_outputs(4870);
    outputs(5387) <= layer2_outputs(6199);
    outputs(5388) <= (layer2_outputs(6181)) and not (layer2_outputs(8229));
    outputs(5389) <= not(layer2_outputs(5859));
    outputs(5390) <= not(layer2_outputs(725));
    outputs(5391) <= not((layer2_outputs(9602)) xor (layer2_outputs(5841)));
    outputs(5392) <= not((layer2_outputs(8833)) and (layer2_outputs(10766)));
    outputs(5393) <= layer2_outputs(5932);
    outputs(5394) <= (layer2_outputs(539)) or (layer2_outputs(7725));
    outputs(5395) <= (layer2_outputs(8273)) xor (layer2_outputs(10710));
    outputs(5396) <= (layer2_outputs(11344)) xor (layer2_outputs(4607));
    outputs(5397) <= not(layer2_outputs(12284));
    outputs(5398) <= not(layer2_outputs(5324));
    outputs(5399) <= not(layer2_outputs(11)) or (layer2_outputs(11950));
    outputs(5400) <= layer2_outputs(6425);
    outputs(5401) <= not(layer2_outputs(2496));
    outputs(5402) <= not(layer2_outputs(9106));
    outputs(5403) <= not(layer2_outputs(8802)) or (layer2_outputs(6225));
    outputs(5404) <= (layer2_outputs(5770)) and not (layer2_outputs(12353));
    outputs(5405) <= not((layer2_outputs(10182)) or (layer2_outputs(9500)));
    outputs(5406) <= (layer2_outputs(5253)) xor (layer2_outputs(5199));
    outputs(5407) <= not(layer2_outputs(10321));
    outputs(5408) <= not((layer2_outputs(11086)) xor (layer2_outputs(810)));
    outputs(5409) <= not(layer2_outputs(11314));
    outputs(5410) <= (layer2_outputs(10048)) xor (layer2_outputs(10642));
    outputs(5411) <= not((layer2_outputs(7451)) xor (layer2_outputs(2438)));
    outputs(5412) <= (layer2_outputs(223)) xor (layer2_outputs(5344));
    outputs(5413) <= not(layer2_outputs(12660));
    outputs(5414) <= not(layer2_outputs(2039));
    outputs(5415) <= not(layer2_outputs(2734));
    outputs(5416) <= layer2_outputs(2825);
    outputs(5417) <= layer2_outputs(7963);
    outputs(5418) <= (layer2_outputs(295)) xor (layer2_outputs(12337));
    outputs(5419) <= not(layer2_outputs(343));
    outputs(5420) <= not(layer2_outputs(3345));
    outputs(5421) <= not((layer2_outputs(6625)) and (layer2_outputs(2999)));
    outputs(5422) <= not(layer2_outputs(7662));
    outputs(5423) <= (layer2_outputs(10867)) xor (layer2_outputs(8112));
    outputs(5424) <= not(layer2_outputs(1302)) or (layer2_outputs(598));
    outputs(5425) <= not((layer2_outputs(9990)) xor (layer2_outputs(5589)));
    outputs(5426) <= not(layer2_outputs(5777)) or (layer2_outputs(11080));
    outputs(5427) <= (layer2_outputs(6486)) or (layer2_outputs(12472));
    outputs(5428) <= layer2_outputs(12296);
    outputs(5429) <= not(layer2_outputs(3139));
    outputs(5430) <= layer2_outputs(11763);
    outputs(5431) <= (layer2_outputs(4739)) and not (layer2_outputs(2509));
    outputs(5432) <= not(layer2_outputs(4558));
    outputs(5433) <= layer2_outputs(2647);
    outputs(5434) <= layer2_outputs(12174);
    outputs(5435) <= not((layer2_outputs(7627)) or (layer2_outputs(2193)));
    outputs(5436) <= layer2_outputs(6381);
    outputs(5437) <= (layer2_outputs(4194)) or (layer2_outputs(7162));
    outputs(5438) <= not(layer2_outputs(12444));
    outputs(5439) <= (layer2_outputs(8859)) xor (layer2_outputs(11303));
    outputs(5440) <= (layer2_outputs(797)) and not (layer2_outputs(4169));
    outputs(5441) <= layer2_outputs(3393);
    outputs(5442) <= not(layer2_outputs(3016));
    outputs(5443) <= (layer2_outputs(1186)) and (layer2_outputs(9586));
    outputs(5444) <= (layer2_outputs(12332)) and not (layer2_outputs(4594));
    outputs(5445) <= not(layer2_outputs(5215));
    outputs(5446) <= layer2_outputs(12143);
    outputs(5447) <= layer2_outputs(1421);
    outputs(5448) <= layer2_outputs(10807);
    outputs(5449) <= not(layer2_outputs(11096));
    outputs(5450) <= layer2_outputs(3760);
    outputs(5451) <= (layer2_outputs(4387)) xor (layer2_outputs(10685));
    outputs(5452) <= layer2_outputs(1260);
    outputs(5453) <= layer2_outputs(6325);
    outputs(5454) <= layer2_outputs(2453);
    outputs(5455) <= (layer2_outputs(2402)) xor (layer2_outputs(4746));
    outputs(5456) <= not(layer2_outputs(8847)) or (layer2_outputs(1090));
    outputs(5457) <= not(layer2_outputs(6496));
    outputs(5458) <= layer2_outputs(12410);
    outputs(5459) <= layer2_outputs(10109);
    outputs(5460) <= not(layer2_outputs(4251)) or (layer2_outputs(7372));
    outputs(5461) <= layer2_outputs(4477);
    outputs(5462) <= not(layer2_outputs(10216));
    outputs(5463) <= not((layer2_outputs(11642)) and (layer2_outputs(4986)));
    outputs(5464) <= not(layer2_outputs(4466));
    outputs(5465) <= not((layer2_outputs(6426)) or (layer2_outputs(4906)));
    outputs(5466) <= (layer2_outputs(12760)) and not (layer2_outputs(1986));
    outputs(5467) <= not(layer2_outputs(10811));
    outputs(5468) <= layer2_outputs(7976);
    outputs(5469) <= (layer2_outputs(622)) xor (layer2_outputs(3800));
    outputs(5470) <= not((layer2_outputs(103)) xor (layer2_outputs(12762)));
    outputs(5471) <= not((layer2_outputs(1045)) xor (layer2_outputs(2421)));
    outputs(5472) <= not(layer2_outputs(5527));
    outputs(5473) <= not(layer2_outputs(10231));
    outputs(5474) <= not(layer2_outputs(11771));
    outputs(5475) <= layer2_outputs(3556);
    outputs(5476) <= layer2_outputs(11364);
    outputs(5477) <= (layer2_outputs(6124)) and (layer2_outputs(2062));
    outputs(5478) <= not(layer2_outputs(3112));
    outputs(5479) <= not(layer2_outputs(4951));
    outputs(5480) <= not((layer2_outputs(5665)) xor (layer2_outputs(6454)));
    outputs(5481) <= not(layer2_outputs(6860));
    outputs(5482) <= (layer2_outputs(9542)) and not (layer2_outputs(11226));
    outputs(5483) <= layer2_outputs(10603);
    outputs(5484) <= layer2_outputs(5601);
    outputs(5485) <= layer2_outputs(12474);
    outputs(5486) <= not(layer2_outputs(8386)) or (layer2_outputs(4173));
    outputs(5487) <= not((layer2_outputs(9116)) xor (layer2_outputs(10291)));
    outputs(5488) <= not(layer2_outputs(4256));
    outputs(5489) <= layer2_outputs(2981);
    outputs(5490) <= not(layer2_outputs(4189));
    outputs(5491) <= layer2_outputs(10849);
    outputs(5492) <= not(layer2_outputs(9721));
    outputs(5493) <= not((layer2_outputs(9358)) xor (layer2_outputs(5855)));
    outputs(5494) <= (layer2_outputs(9115)) and not (layer2_outputs(10219));
    outputs(5495) <= not(layer2_outputs(10165)) or (layer2_outputs(1802));
    outputs(5496) <= not(layer2_outputs(11521));
    outputs(5497) <= not((layer2_outputs(265)) xor (layer2_outputs(6014)));
    outputs(5498) <= not(layer2_outputs(3618));
    outputs(5499) <= not(layer2_outputs(799));
    outputs(5500) <= (layer2_outputs(5893)) xor (layer2_outputs(9850));
    outputs(5501) <= not(layer2_outputs(374));
    outputs(5502) <= (layer2_outputs(7100)) xor (layer2_outputs(6058));
    outputs(5503) <= layer2_outputs(12300);
    outputs(5504) <= not((layer2_outputs(8025)) xor (layer2_outputs(1742)));
    outputs(5505) <= (layer2_outputs(5833)) xor (layer2_outputs(5550));
    outputs(5506) <= (layer2_outputs(5767)) xor (layer2_outputs(9432));
    outputs(5507) <= not((layer2_outputs(10742)) xor (layer2_outputs(7014)));
    outputs(5508) <= (layer2_outputs(4080)) or (layer2_outputs(10577));
    outputs(5509) <= layer2_outputs(11372);
    outputs(5510) <= (layer2_outputs(9093)) xor (layer2_outputs(10310));
    outputs(5511) <= (layer2_outputs(7803)) and (layer2_outputs(11119));
    outputs(5512) <= not(layer2_outputs(10700));
    outputs(5513) <= layer2_outputs(3730);
    outputs(5514) <= (layer2_outputs(7390)) and not (layer2_outputs(5137));
    outputs(5515) <= (layer2_outputs(11055)) and (layer2_outputs(122));
    outputs(5516) <= not(layer2_outputs(5588)) or (layer2_outputs(1862));
    outputs(5517) <= layer2_outputs(8021);
    outputs(5518) <= (layer2_outputs(390)) xor (layer2_outputs(6133));
    outputs(5519) <= layer2_outputs(9645);
    outputs(5520) <= not(layer2_outputs(11174));
    outputs(5521) <= layer2_outputs(8230);
    outputs(5522) <= layer2_outputs(2122);
    outputs(5523) <= not(layer2_outputs(512));
    outputs(5524) <= not((layer2_outputs(11665)) xor (layer2_outputs(3747)));
    outputs(5525) <= not(layer2_outputs(1461));
    outputs(5526) <= (layer2_outputs(3758)) xor (layer2_outputs(10770));
    outputs(5527) <= (layer2_outputs(10303)) xor (layer2_outputs(6837));
    outputs(5528) <= (layer2_outputs(3960)) and (layer2_outputs(12388));
    outputs(5529) <= layer2_outputs(1616);
    outputs(5530) <= layer2_outputs(6418);
    outputs(5531) <= not((layer2_outputs(12252)) or (layer2_outputs(10113)));
    outputs(5532) <= (layer2_outputs(2849)) and (layer2_outputs(2293));
    outputs(5533) <= not((layer2_outputs(2671)) and (layer2_outputs(12190)));
    outputs(5534) <= not((layer2_outputs(2352)) xor (layer2_outputs(12549)));
    outputs(5535) <= not(layer2_outputs(11324));
    outputs(5536) <= layer2_outputs(4911);
    outputs(5537) <= (layer2_outputs(3335)) and (layer2_outputs(8358));
    outputs(5538) <= not(layer2_outputs(23));
    outputs(5539) <= layer2_outputs(1642);
    outputs(5540) <= not(layer2_outputs(3146));
    outputs(5541) <= (layer2_outputs(1623)) xor (layer2_outputs(6134));
    outputs(5542) <= not((layer2_outputs(1405)) and (layer2_outputs(11014)));
    outputs(5543) <= (layer2_outputs(4214)) xor (layer2_outputs(8985));
    outputs(5544) <= not(layer2_outputs(988));
    outputs(5545) <= layer2_outputs(775);
    outputs(5546) <= not((layer2_outputs(8169)) xor (layer2_outputs(2272)));
    outputs(5547) <= not(layer2_outputs(1747)) or (layer2_outputs(11638));
    outputs(5548) <= (layer2_outputs(10073)) or (layer2_outputs(8257));
    outputs(5549) <= layer2_outputs(6132);
    outputs(5550) <= not(layer2_outputs(3321));
    outputs(5551) <= layer2_outputs(3723);
    outputs(5552) <= not(layer2_outputs(8530));
    outputs(5553) <= not(layer2_outputs(5553));
    outputs(5554) <= layer2_outputs(10143);
    outputs(5555) <= not((layer2_outputs(2105)) xor (layer2_outputs(12095)));
    outputs(5556) <= not(layer2_outputs(4670)) or (layer2_outputs(11172));
    outputs(5557) <= layer2_outputs(1575);
    outputs(5558) <= not(layer2_outputs(627));
    outputs(5559) <= not(layer2_outputs(11585));
    outputs(5560) <= layer2_outputs(5054);
    outputs(5561) <= (layer2_outputs(208)) xor (layer2_outputs(1149));
    outputs(5562) <= not(layer2_outputs(4403));
    outputs(5563) <= layer2_outputs(11801);
    outputs(5564) <= not(layer2_outputs(2316));
    outputs(5565) <= (layer2_outputs(6802)) and not (layer2_outputs(1793));
    outputs(5566) <= (layer2_outputs(6337)) xor (layer2_outputs(6673));
    outputs(5567) <= layer2_outputs(10524);
    outputs(5568) <= (layer2_outputs(1654)) xor (layer2_outputs(7711));
    outputs(5569) <= not(layer2_outputs(2384));
    outputs(5570) <= layer2_outputs(11922);
    outputs(5571) <= layer2_outputs(6685);
    outputs(5572) <= not(layer2_outputs(1841));
    outputs(5573) <= layer2_outputs(8580);
    outputs(5574) <= layer2_outputs(4561);
    outputs(5575) <= not((layer2_outputs(206)) xor (layer2_outputs(472)));
    outputs(5576) <= not(layer2_outputs(12075));
    outputs(5577) <= not(layer2_outputs(8770));
    outputs(5578) <= not((layer2_outputs(2635)) xor (layer2_outputs(6139)));
    outputs(5579) <= not(layer2_outputs(3820));
    outputs(5580) <= layer2_outputs(6107);
    outputs(5581) <= not((layer2_outputs(8197)) xor (layer2_outputs(6762)));
    outputs(5582) <= (layer2_outputs(185)) xor (layer2_outputs(4024));
    outputs(5583) <= not(layer2_outputs(7738)) or (layer2_outputs(5246));
    outputs(5584) <= (layer2_outputs(8619)) and (layer2_outputs(688));
    outputs(5585) <= not(layer2_outputs(7369));
    outputs(5586) <= (layer2_outputs(1126)) xor (layer2_outputs(4086));
    outputs(5587) <= not((layer2_outputs(8442)) xor (layer2_outputs(8727)));
    outputs(5588) <= not(layer2_outputs(9954));
    outputs(5589) <= not(layer2_outputs(5536));
    outputs(5590) <= layer2_outputs(4933);
    outputs(5591) <= layer2_outputs(5818);
    outputs(5592) <= layer2_outputs(1719);
    outputs(5593) <= not((layer2_outputs(8776)) or (layer2_outputs(1191)));
    outputs(5594) <= not(layer2_outputs(7309));
    outputs(5595) <= not((layer2_outputs(3268)) xor (layer2_outputs(8752)));
    outputs(5596) <= (layer2_outputs(8380)) xor (layer2_outputs(1384));
    outputs(5597) <= not(layer2_outputs(12568));
    outputs(5598) <= not(layer2_outputs(7227));
    outputs(5599) <= layer2_outputs(1941);
    outputs(5600) <= (layer2_outputs(4976)) and not (layer2_outputs(2077));
    outputs(5601) <= not((layer2_outputs(2505)) xor (layer2_outputs(10695)));
    outputs(5602) <= not(layer2_outputs(8088));
    outputs(5603) <= not((layer2_outputs(11466)) xor (layer2_outputs(363)));
    outputs(5604) <= (layer2_outputs(5988)) xor (layer2_outputs(8713));
    outputs(5605) <= not((layer2_outputs(3847)) xor (layer2_outputs(10736)));
    outputs(5606) <= layer2_outputs(6886);
    outputs(5607) <= layer2_outputs(3318);
    outputs(5608) <= (layer2_outputs(1570)) xor (layer2_outputs(2312));
    outputs(5609) <= layer2_outputs(5187);
    outputs(5610) <= not(layer2_outputs(2839)) or (layer2_outputs(1856));
    outputs(5611) <= not(layer2_outputs(3180));
    outputs(5612) <= not(layer2_outputs(9958));
    outputs(5613) <= not((layer2_outputs(4526)) xor (layer2_outputs(1619)));
    outputs(5614) <= not(layer2_outputs(7986));
    outputs(5615) <= (layer2_outputs(4118)) xor (layer2_outputs(11218));
    outputs(5616) <= layer2_outputs(10881);
    outputs(5617) <= (layer2_outputs(3409)) xor (layer2_outputs(3094));
    outputs(5618) <= not(layer2_outputs(2345));
    outputs(5619) <= not(layer2_outputs(274)) or (layer2_outputs(5752));
    outputs(5620) <= not(layer2_outputs(6779));
    outputs(5621) <= layer2_outputs(12342);
    outputs(5622) <= (layer2_outputs(10087)) xor (layer2_outputs(1320));
    outputs(5623) <= not((layer2_outputs(84)) and (layer2_outputs(8955)));
    outputs(5624) <= (layer2_outputs(524)) xor (layer2_outputs(613));
    outputs(5625) <= layer2_outputs(4440);
    outputs(5626) <= (layer2_outputs(5935)) xor (layer2_outputs(9372));
    outputs(5627) <= (layer2_outputs(1229)) and (layer2_outputs(461));
    outputs(5628) <= not((layer2_outputs(4021)) xor (layer2_outputs(8556)));
    outputs(5629) <= not(layer2_outputs(1751));
    outputs(5630) <= not(layer2_outputs(10985));
    outputs(5631) <= not((layer2_outputs(11209)) xor (layer2_outputs(1016)));
    outputs(5632) <= (layer2_outputs(3378)) xor (layer2_outputs(9234));
    outputs(5633) <= (layer2_outputs(12170)) xor (layer2_outputs(12742));
    outputs(5634) <= layer2_outputs(10129);
    outputs(5635) <= not((layer2_outputs(6390)) xor (layer2_outputs(301)));
    outputs(5636) <= (layer2_outputs(1231)) xor (layer2_outputs(10684));
    outputs(5637) <= layer2_outputs(10183);
    outputs(5638) <= not(layer2_outputs(8391));
    outputs(5639) <= not(layer2_outputs(2171));
    outputs(5640) <= not(layer2_outputs(4494));
    outputs(5641) <= (layer2_outputs(9759)) and not (layer2_outputs(9432));
    outputs(5642) <= not(layer2_outputs(11939));
    outputs(5643) <= not((layer2_outputs(11613)) or (layer2_outputs(2959)));
    outputs(5644) <= not((layer2_outputs(1810)) xor (layer2_outputs(9611)));
    outputs(5645) <= not(layer2_outputs(6512));
    outputs(5646) <= not((layer2_outputs(7154)) xor (layer2_outputs(7377)));
    outputs(5647) <= not(layer2_outputs(1391));
    outputs(5648) <= (layer2_outputs(2889)) xor (layer2_outputs(10140));
    outputs(5649) <= not(layer2_outputs(3180));
    outputs(5650) <= (layer2_outputs(6736)) and (layer2_outputs(5304));
    outputs(5651) <= layer2_outputs(7083);
    outputs(5652) <= not((layer2_outputs(5442)) xor (layer2_outputs(309)));
    outputs(5653) <= (layer2_outputs(6787)) xor (layer2_outputs(11035));
    outputs(5654) <= not(layer2_outputs(259));
    outputs(5655) <= layer2_outputs(3669);
    outputs(5656) <= not(layer2_outputs(108));
    outputs(5657) <= not(layer2_outputs(1975));
    outputs(5658) <= not(layer2_outputs(9110));
    outputs(5659) <= not(layer2_outputs(9076));
    outputs(5660) <= layer2_outputs(4861);
    outputs(5661) <= layer2_outputs(195);
    outputs(5662) <= layer2_outputs(10910);
    outputs(5663) <= layer2_outputs(11330);
    outputs(5664) <= not((layer2_outputs(3790)) and (layer2_outputs(10824)));
    outputs(5665) <= (layer2_outputs(3590)) and not (layer2_outputs(8299));
    outputs(5666) <= layer2_outputs(8960);
    outputs(5667) <= not((layer2_outputs(10209)) xor (layer2_outputs(10016)));
    outputs(5668) <= layer2_outputs(5329);
    outputs(5669) <= layer2_outputs(8041);
    outputs(5670) <= not((layer2_outputs(12090)) xor (layer2_outputs(1811)));
    outputs(5671) <= layer2_outputs(4496);
    outputs(5672) <= layer2_outputs(3730);
    outputs(5673) <= (layer2_outputs(9395)) xor (layer2_outputs(5227));
    outputs(5674) <= not(layer2_outputs(577));
    outputs(5675) <= layer2_outputs(1288);
    outputs(5676) <= not(layer2_outputs(4728));
    outputs(5677) <= layer2_outputs(5559);
    outputs(5678) <= not(layer2_outputs(7819));
    outputs(5679) <= (layer2_outputs(11117)) and not (layer2_outputs(6729));
    outputs(5680) <= (layer2_outputs(3215)) and (layer2_outputs(12433));
    outputs(5681) <= not(layer2_outputs(2754));
    outputs(5682) <= not(layer2_outputs(7069));
    outputs(5683) <= (layer2_outputs(11350)) and (layer2_outputs(72));
    outputs(5684) <= (layer2_outputs(12421)) xor (layer2_outputs(6822));
    outputs(5685) <= not((layer2_outputs(8177)) xor (layer2_outputs(11536)));
    outputs(5686) <= not(layer2_outputs(9206));
    outputs(5687) <= not((layer2_outputs(9041)) or (layer2_outputs(3429)));
    outputs(5688) <= layer2_outputs(2064);
    outputs(5689) <= not(layer2_outputs(4157));
    outputs(5690) <= not(layer2_outputs(3966));
    outputs(5691) <= (layer2_outputs(2195)) xor (layer2_outputs(10851));
    outputs(5692) <= not((layer2_outputs(5199)) xor (layer2_outputs(11673)));
    outputs(5693) <= not(layer2_outputs(2538)) or (layer2_outputs(12681));
    outputs(5694) <= not(layer2_outputs(544));
    outputs(5695) <= not(layer2_outputs(4512));
    outputs(5696) <= not(layer2_outputs(7473));
    outputs(5697) <= layer2_outputs(1590);
    outputs(5698) <= not((layer2_outputs(11891)) xor (layer2_outputs(4263)));
    outputs(5699) <= (layer2_outputs(7756)) xor (layer2_outputs(3884));
    outputs(5700) <= layer2_outputs(6051);
    outputs(5701) <= not(layer2_outputs(9896));
    outputs(5702) <= layer2_outputs(11249);
    outputs(5703) <= (layer2_outputs(6879)) xor (layer2_outputs(7125));
    outputs(5704) <= (layer2_outputs(7006)) xor (layer2_outputs(4863));
    outputs(5705) <= layer2_outputs(8721);
    outputs(5706) <= not(layer2_outputs(2812));
    outputs(5707) <= not(layer2_outputs(9504));
    outputs(5708) <= not((layer2_outputs(5819)) or (layer2_outputs(6848)));
    outputs(5709) <= not(layer2_outputs(3350));
    outputs(5710) <= not((layer2_outputs(11271)) xor (layer2_outputs(3205)));
    outputs(5711) <= layer2_outputs(7305);
    outputs(5712) <= not(layer2_outputs(3371));
    outputs(5713) <= not(layer2_outputs(2971));
    outputs(5714) <= layer2_outputs(2396);
    outputs(5715) <= not(layer2_outputs(4782));
    outputs(5716) <= not(layer2_outputs(7694));
    outputs(5717) <= not(layer2_outputs(8683));
    outputs(5718) <= layer2_outputs(11658);
    outputs(5719) <= layer2_outputs(1435);
    outputs(5720) <= not(layer2_outputs(7975));
    outputs(5721) <= not((layer2_outputs(1968)) xor (layer2_outputs(176)));
    outputs(5722) <= not(layer2_outputs(3128));
    outputs(5723) <= not(layer2_outputs(5021));
    outputs(5724) <= (layer2_outputs(12706)) or (layer2_outputs(1262));
    outputs(5725) <= layer2_outputs(11063);
    outputs(5726) <= not(layer2_outputs(60));
    outputs(5727) <= not(layer2_outputs(1185));
    outputs(5728) <= layer2_outputs(5280);
    outputs(5729) <= not(layer2_outputs(9375));
    outputs(5730) <= (layer2_outputs(8048)) or (layer2_outputs(5931));
    outputs(5731) <= layer2_outputs(8828);
    outputs(5732) <= (layer2_outputs(11402)) xor (layer2_outputs(4063));
    outputs(5733) <= layer2_outputs(5558);
    outputs(5734) <= not(layer2_outputs(1617));
    outputs(5735) <= (layer2_outputs(3639)) xor (layer2_outputs(7273));
    outputs(5736) <= not(layer2_outputs(11747));
    outputs(5737) <= not(layer2_outputs(6913));
    outputs(5738) <= not(layer2_outputs(9527));
    outputs(5739) <= not((layer2_outputs(2899)) xor (layer2_outputs(5205)));
    outputs(5740) <= not(layer2_outputs(5250));
    outputs(5741) <= layer2_outputs(4219);
    outputs(5742) <= not(layer2_outputs(11091));
    outputs(5743) <= (layer2_outputs(10886)) xor (layer2_outputs(1303));
    outputs(5744) <= not(layer2_outputs(12377));
    outputs(5745) <= not(layer2_outputs(11032));
    outputs(5746) <= not((layer2_outputs(7243)) xor (layer2_outputs(11388)));
    outputs(5747) <= not(layer2_outputs(4610));
    outputs(5748) <= layer2_outputs(4132);
    outputs(5749) <= layer2_outputs(12058);
    outputs(5750) <= (layer2_outputs(8937)) and not (layer2_outputs(1597));
    outputs(5751) <= layer2_outputs(3675);
    outputs(5752) <= layer2_outputs(6411);
    outputs(5753) <= not(layer2_outputs(6303));
    outputs(5754) <= not((layer2_outputs(1908)) or (layer2_outputs(11367)));
    outputs(5755) <= not((layer2_outputs(7745)) xor (layer2_outputs(5637)));
    outputs(5756) <= (layer2_outputs(6405)) or (layer2_outputs(1336));
    outputs(5757) <= not(layer2_outputs(12305));
    outputs(5758) <= layer2_outputs(11410);
    outputs(5759) <= layer2_outputs(1973);
    outputs(5760) <= not((layer2_outputs(11941)) or (layer2_outputs(8871)));
    outputs(5761) <= (layer2_outputs(6300)) xor (layer2_outputs(8734));
    outputs(5762) <= not((layer2_outputs(7655)) and (layer2_outputs(7192)));
    outputs(5763) <= (layer2_outputs(5532)) and not (layer2_outputs(8797));
    outputs(5764) <= layer2_outputs(6777);
    outputs(5765) <= not(layer2_outputs(1276));
    outputs(5766) <= layer2_outputs(11511);
    outputs(5767) <= (layer2_outputs(4947)) xor (layer2_outputs(6297));
    outputs(5768) <= not((layer2_outputs(4731)) xor (layer2_outputs(11309)));
    outputs(5769) <= not(layer2_outputs(5620));
    outputs(5770) <= (layer2_outputs(10820)) xor (layer2_outputs(6248));
    outputs(5771) <= (layer2_outputs(10874)) xor (layer2_outputs(2136));
    outputs(5772) <= not((layer2_outputs(7115)) xor (layer2_outputs(6714)));
    outputs(5773) <= layer2_outputs(9761);
    outputs(5774) <= (layer2_outputs(10650)) and (layer2_outputs(3416));
    outputs(5775) <= not(layer2_outputs(6731));
    outputs(5776) <= layer2_outputs(8639);
    outputs(5777) <= not(layer2_outputs(7668));
    outputs(5778) <= not(layer2_outputs(7393)) or (layer2_outputs(6293));
    outputs(5779) <= not((layer2_outputs(8174)) xor (layer2_outputs(8151)));
    outputs(5780) <= (layer2_outputs(3819)) xor (layer2_outputs(12355));
    outputs(5781) <= layer2_outputs(1890);
    outputs(5782) <= not((layer2_outputs(9592)) or (layer2_outputs(5259)));
    outputs(5783) <= layer2_outputs(323);
    outputs(5784) <= (layer2_outputs(3007)) xor (layer2_outputs(7548));
    outputs(5785) <= (layer2_outputs(4965)) xor (layer2_outputs(669));
    outputs(5786) <= not(layer2_outputs(9202)) or (layer2_outputs(10544));
    outputs(5787) <= not(layer2_outputs(8621));
    outputs(5788) <= not(layer2_outputs(11555)) or (layer2_outputs(8271));
    outputs(5789) <= layer2_outputs(11351);
    outputs(5790) <= layer2_outputs(7362);
    outputs(5791) <= layer2_outputs(2690);
    outputs(5792) <= not(layer2_outputs(4736)) or (layer2_outputs(1632));
    outputs(5793) <= layer2_outputs(3387);
    outputs(5794) <= layer2_outputs(6148);
    outputs(5795) <= (layer2_outputs(3999)) or (layer2_outputs(2837));
    outputs(5796) <= not(layer2_outputs(1212));
    outputs(5797) <= (layer2_outputs(12372)) xor (layer2_outputs(10178));
    outputs(5798) <= layer2_outputs(9939);
    outputs(5799) <= not(layer2_outputs(12135));
    outputs(5800) <= layer2_outputs(713);
    outputs(5801) <= (layer2_outputs(11549)) xor (layer2_outputs(10927));
    outputs(5802) <= (layer2_outputs(11902)) xor (layer2_outputs(6142));
    outputs(5803) <= layer2_outputs(8287);
    outputs(5804) <= (layer2_outputs(2833)) and (layer2_outputs(5867));
    outputs(5805) <= layer2_outputs(3753);
    outputs(5806) <= layer2_outputs(3057);
    outputs(5807) <= (layer2_outputs(10009)) and not (layer2_outputs(3049));
    outputs(5808) <= not(layer2_outputs(4078));
    outputs(5809) <= (layer2_outputs(6332)) xor (layer2_outputs(9913));
    outputs(5810) <= not(layer2_outputs(9246)) or (layer2_outputs(1226));
    outputs(5811) <= layer2_outputs(7237);
    outputs(5812) <= layer2_outputs(8221);
    outputs(5813) <= layer2_outputs(8154);
    outputs(5814) <= layer2_outputs(8790);
    outputs(5815) <= not((layer2_outputs(4184)) xor (layer2_outputs(7690)));
    outputs(5816) <= not((layer2_outputs(12004)) and (layer2_outputs(4991)));
    outputs(5817) <= not((layer2_outputs(2102)) xor (layer2_outputs(7194)));
    outputs(5818) <= not(layer2_outputs(3151));
    outputs(5819) <= (layer2_outputs(4103)) and not (layer2_outputs(3817));
    outputs(5820) <= not((layer2_outputs(10696)) xor (layer2_outputs(10998)));
    outputs(5821) <= (layer2_outputs(8344)) xor (layer2_outputs(1413));
    outputs(5822) <= not(layer2_outputs(302));
    outputs(5823) <= layer2_outputs(9972);
    outputs(5824) <= layer2_outputs(9472);
    outputs(5825) <= layer2_outputs(4703);
    outputs(5826) <= not((layer2_outputs(384)) xor (layer2_outputs(2494)));
    outputs(5827) <= not(layer2_outputs(9279));
    outputs(5828) <= not(layer2_outputs(8068));
    outputs(5829) <= (layer2_outputs(2449)) xor (layer2_outputs(4166));
    outputs(5830) <= not(layer2_outputs(2674));
    outputs(5831) <= not(layer2_outputs(9004));
    outputs(5832) <= (layer2_outputs(2844)) xor (layer2_outputs(12243));
    outputs(5833) <= not(layer2_outputs(5521));
    outputs(5834) <= (layer2_outputs(6965)) xor (layer2_outputs(6947));
    outputs(5835) <= (layer2_outputs(10012)) or (layer2_outputs(907));
    outputs(5836) <= not((layer2_outputs(60)) xor (layer2_outputs(2355)));
    outputs(5837) <= not((layer2_outputs(2262)) or (layer2_outputs(8138)));
    outputs(5838) <= (layer2_outputs(790)) and not (layer2_outputs(1523));
    outputs(5839) <= not(layer2_outputs(598)) or (layer2_outputs(3236));
    outputs(5840) <= layer2_outputs(5288);
    outputs(5841) <= (layer2_outputs(9947)) and (layer2_outputs(1238));
    outputs(5842) <= not(layer2_outputs(10749));
    outputs(5843) <= layer2_outputs(4832);
    outputs(5844) <= not(layer2_outputs(6764));
    outputs(5845) <= not(layer2_outputs(6742));
    outputs(5846) <= layer2_outputs(7464);
    outputs(5847) <= not(layer2_outputs(1503));
    outputs(5848) <= not(layer2_outputs(12420));
    outputs(5849) <= not(layer2_outputs(8039));
    outputs(5850) <= not(layer2_outputs(10841));
    outputs(5851) <= layer2_outputs(2103);
    outputs(5852) <= layer2_outputs(535);
    outputs(5853) <= layer2_outputs(6938);
    outputs(5854) <= (layer2_outputs(12663)) xor (layer2_outputs(6989));
    outputs(5855) <= not(layer2_outputs(12413));
    outputs(5856) <= not((layer2_outputs(3765)) xor (layer2_outputs(895)));
    outputs(5857) <= layer2_outputs(3545);
    outputs(5858) <= not(layer2_outputs(2200));
    outputs(5859) <= (layer2_outputs(5310)) or (layer2_outputs(10779));
    outputs(5860) <= not(layer2_outputs(6833));
    outputs(5861) <= not(layer2_outputs(3928));
    outputs(5862) <= layer2_outputs(8024);
    outputs(5863) <= not(layer2_outputs(3422));
    outputs(5864) <= not(layer2_outputs(6170));
    outputs(5865) <= not((layer2_outputs(8083)) xor (layer2_outputs(12658)));
    outputs(5866) <= not(layer2_outputs(4631)) or (layer2_outputs(8749));
    outputs(5867) <= (layer2_outputs(8794)) xor (layer2_outputs(3091));
    outputs(5868) <= not((layer2_outputs(1178)) xor (layer2_outputs(9701)));
    outputs(5869) <= layer2_outputs(3473);
    outputs(5870) <= not((layer2_outputs(2142)) and (layer2_outputs(6564)));
    outputs(5871) <= not(layer2_outputs(564));
    outputs(5872) <= layer2_outputs(2294);
    outputs(5873) <= (layer2_outputs(166)) or (layer2_outputs(2783));
    outputs(5874) <= (layer2_outputs(4005)) xor (layer2_outputs(12453));
    outputs(5875) <= layer2_outputs(3562);
    outputs(5876) <= not(layer2_outputs(9515));
    outputs(5877) <= layer2_outputs(3);
    outputs(5878) <= layer2_outputs(5806);
    outputs(5879) <= not(layer2_outputs(6950)) or (layer2_outputs(8543));
    outputs(5880) <= not(layer2_outputs(8464));
    outputs(5881) <= not(layer2_outputs(5579)) or (layer2_outputs(8673));
    outputs(5882) <= layer2_outputs(4745);
    outputs(5883) <= not(layer2_outputs(11520));
    outputs(5884) <= not(layer2_outputs(3284));
    outputs(5885) <= not(layer2_outputs(5769));
    outputs(5886) <= not(layer2_outputs(12698));
    outputs(5887) <= layer2_outputs(12515);
    outputs(5888) <= (layer2_outputs(6080)) and not (layer2_outputs(2565));
    outputs(5889) <= not((layer2_outputs(11471)) xor (layer2_outputs(9978)));
    outputs(5890) <= not((layer2_outputs(12074)) xor (layer2_outputs(2570)));
    outputs(5891) <= not((layer2_outputs(8644)) xor (layer2_outputs(584)));
    outputs(5892) <= not((layer2_outputs(6147)) xor (layer2_outputs(4151)));
    outputs(5893) <= not((layer2_outputs(12572)) xor (layer2_outputs(11234)));
    outputs(5894) <= not(layer2_outputs(9249)) or (layer2_outputs(6501));
    outputs(5895) <= not(layer2_outputs(10696));
    outputs(5896) <= not(layer2_outputs(12670));
    outputs(5897) <= (layer2_outputs(9007)) and not (layer2_outputs(2277));
    outputs(5898) <= (layer2_outputs(7171)) or (layer2_outputs(1724));
    outputs(5899) <= not(layer2_outputs(1318)) or (layer2_outputs(381));
    outputs(5900) <= layer2_outputs(11341);
    outputs(5901) <= layer2_outputs(7030);
    outputs(5902) <= not((layer2_outputs(7817)) or (layer2_outputs(6363)));
    outputs(5903) <= layer2_outputs(6418);
    outputs(5904) <= not(layer2_outputs(10763));
    outputs(5905) <= (layer2_outputs(5854)) xor (layer2_outputs(7140));
    outputs(5906) <= layer2_outputs(662);
    outputs(5907) <= not(layer2_outputs(12311));
    outputs(5908) <= layer2_outputs(9750);
    outputs(5909) <= (layer2_outputs(8196)) xor (layer2_outputs(12508));
    outputs(5910) <= (layer2_outputs(5000)) and not (layer2_outputs(6153));
    outputs(5911) <= layer2_outputs(277);
    outputs(5912) <= (layer2_outputs(9754)) and not (layer2_outputs(2925));
    outputs(5913) <= (layer2_outputs(1)) xor (layer2_outputs(10838));
    outputs(5914) <= layer2_outputs(1178);
    outputs(5915) <= (layer2_outputs(9756)) and not (layer2_outputs(1643));
    outputs(5916) <= layer2_outputs(5435);
    outputs(5917) <= not((layer2_outputs(443)) xor (layer2_outputs(1253)));
    outputs(5918) <= (layer2_outputs(3412)) xor (layer2_outputs(6662));
    outputs(5919) <= layer2_outputs(35);
    outputs(5920) <= layer2_outputs(2479);
    outputs(5921) <= layer2_outputs(6652);
    outputs(5922) <= layer2_outputs(5214);
    outputs(5923) <= (layer2_outputs(7974)) xor (layer2_outputs(2588));
    outputs(5924) <= not(layer2_outputs(494));
    outputs(5925) <= not(layer2_outputs(3594));
    outputs(5926) <= not(layer2_outputs(271)) or (layer2_outputs(2146));
    outputs(5927) <= layer2_outputs(6760);
    outputs(5928) <= not(layer2_outputs(8170));
    outputs(5929) <= not((layer2_outputs(10451)) xor (layer2_outputs(11181)));
    outputs(5930) <= not(layer2_outputs(8253)) or (layer2_outputs(3445));
    outputs(5931) <= layer2_outputs(11726);
    outputs(5932) <= not(layer2_outputs(12657));
    outputs(5933) <= layer2_outputs(12124);
    outputs(5934) <= layer2_outputs(9094);
    outputs(5935) <= layer2_outputs(5494);
    outputs(5936) <= (layer2_outputs(6399)) or (layer2_outputs(9437));
    outputs(5937) <= layer2_outputs(9411);
    outputs(5938) <= not(layer2_outputs(367)) or (layer2_outputs(4752));
    outputs(5939) <= not((layer2_outputs(4146)) xor (layer2_outputs(3356)));
    outputs(5940) <= not((layer2_outputs(9416)) xor (layer2_outputs(10454)));
    outputs(5941) <= (layer2_outputs(6462)) and not (layer2_outputs(4527));
    outputs(5942) <= not(layer2_outputs(1132));
    outputs(5943) <= not((layer2_outputs(10318)) xor (layer2_outputs(3867)));
    outputs(5944) <= not(layer2_outputs(2342));
    outputs(5945) <= not(layer2_outputs(4748));
    outputs(5946) <= layer2_outputs(7132);
    outputs(5947) <= layer2_outputs(2956);
    outputs(5948) <= layer2_outputs(6549);
    outputs(5949) <= not((layer2_outputs(93)) or (layer2_outputs(8485)));
    outputs(5950) <= not((layer2_outputs(6366)) xor (layer2_outputs(7870)));
    outputs(5951) <= layer2_outputs(10918);
    outputs(5952) <= (layer2_outputs(228)) and not (layer2_outputs(7137));
    outputs(5953) <= not(layer2_outputs(7928));
    outputs(5954) <= (layer2_outputs(2424)) and not (layer2_outputs(957));
    outputs(5955) <= not((layer2_outputs(9309)) xor (layer2_outputs(3404)));
    outputs(5956) <= not(layer2_outputs(2675));
    outputs(5957) <= (layer2_outputs(606)) or (layer2_outputs(12360));
    outputs(5958) <= not(layer2_outputs(340));
    outputs(5959) <= not(layer2_outputs(7543));
    outputs(5960) <= not(layer2_outputs(4131));
    outputs(5961) <= layer2_outputs(794);
    outputs(5962) <= (layer2_outputs(832)) xor (layer2_outputs(10830));
    outputs(5963) <= layer2_outputs(10466);
    outputs(5964) <= layer2_outputs(9893);
    outputs(5965) <= not((layer2_outputs(1219)) xor (layer2_outputs(9669)));
    outputs(5966) <= not((layer2_outputs(10861)) xor (layer2_outputs(9549)));
    outputs(5967) <= layer2_outputs(9915);
    outputs(5968) <= not((layer2_outputs(12145)) xor (layer2_outputs(7327)));
    outputs(5969) <= (layer2_outputs(205)) xor (layer2_outputs(7238));
    outputs(5970) <= layer2_outputs(7215);
    outputs(5971) <= not((layer2_outputs(5502)) and (layer2_outputs(10878)));
    outputs(5972) <= (layer2_outputs(4298)) xor (layer2_outputs(7564));
    outputs(5973) <= layer2_outputs(11584);
    outputs(5974) <= not((layer2_outputs(4129)) xor (layer2_outputs(4967)));
    outputs(5975) <= layer2_outputs(6782);
    outputs(5976) <= not(layer2_outputs(9403));
    outputs(5977) <= not(layer2_outputs(2017));
    outputs(5978) <= not(layer2_outputs(1964));
    outputs(5979) <= not((layer2_outputs(12059)) xor (layer2_outputs(1534)));
    outputs(5980) <= not(layer2_outputs(10267));
    outputs(5981) <= not(layer2_outputs(11402));
    outputs(5982) <= not(layer2_outputs(8750));
    outputs(5983) <= not(layer2_outputs(4033));
    outputs(5984) <= layer2_outputs(11693);
    outputs(5985) <= not(layer2_outputs(8974)) or (layer2_outputs(5001));
    outputs(5986) <= not((layer2_outputs(4428)) xor (layer2_outputs(5582)));
    outputs(5987) <= (layer2_outputs(4921)) xor (layer2_outputs(9525));
    outputs(5988) <= layer2_outputs(11349);
    outputs(5989) <= (layer2_outputs(1087)) xor (layer2_outputs(158));
    outputs(5990) <= layer2_outputs(6878);
    outputs(5991) <= not((layer2_outputs(9304)) xor (layer2_outputs(9588)));
    outputs(5992) <= (layer2_outputs(10146)) and not (layer2_outputs(8488));
    outputs(5993) <= (layer2_outputs(4004)) and not (layer2_outputs(4642));
    outputs(5994) <= not(layer2_outputs(5173));
    outputs(5995) <= layer2_outputs(8135);
    outputs(5996) <= not(layer2_outputs(9946));
    outputs(5997) <= not(layer2_outputs(9728)) or (layer2_outputs(429));
    outputs(5998) <= layer2_outputs(6361);
    outputs(5999) <= not(layer2_outputs(6811));
    outputs(6000) <= layer2_outputs(9467);
    outputs(6001) <= not(layer2_outputs(7708));
    outputs(6002) <= layer2_outputs(6148);
    outputs(6003) <= layer2_outputs(6771);
    outputs(6004) <= (layer2_outputs(913)) and not (layer2_outputs(7791));
    outputs(6005) <= (layer2_outputs(2506)) xor (layer2_outputs(10103));
    outputs(6006) <= not(layer2_outputs(5264));
    outputs(6007) <= not((layer2_outputs(3189)) xor (layer2_outputs(4638)));
    outputs(6008) <= layer2_outputs(4855);
    outputs(6009) <= layer2_outputs(12488);
    outputs(6010) <= not(layer2_outputs(1001));
    outputs(6011) <= layer2_outputs(49);
    outputs(6012) <= not(layer2_outputs(1093));
    outputs(6013) <= layer2_outputs(6458);
    outputs(6014) <= (layer2_outputs(12258)) and not (layer2_outputs(10478));
    outputs(6015) <= (layer2_outputs(3887)) xor (layer2_outputs(547));
    outputs(6016) <= not(layer2_outputs(886));
    outputs(6017) <= not(layer2_outputs(8947)) or (layer2_outputs(2941));
    outputs(6018) <= not(layer2_outputs(9823));
    outputs(6019) <= layer2_outputs(12047);
    outputs(6020) <= not((layer2_outputs(10969)) xor (layer2_outputs(8668)));
    outputs(6021) <= not(layer2_outputs(10986));
    outputs(6022) <= layer2_outputs(7045);
    outputs(6023) <= layer2_outputs(4956);
    outputs(6024) <= not((layer2_outputs(10071)) xor (layer2_outputs(712)));
    outputs(6025) <= (layer2_outputs(11313)) xor (layer2_outputs(10852));
    outputs(6026) <= not(layer2_outputs(3195));
    outputs(6027) <= not(layer2_outputs(3213));
    outputs(6028) <= not(layer2_outputs(1007));
    outputs(6029) <= not(layer2_outputs(10652));
    outputs(6030) <= (layer2_outputs(6427)) xor (layer2_outputs(11732));
    outputs(6031) <= not((layer2_outputs(6020)) or (layer2_outputs(12334)));
    outputs(6032) <= not(layer2_outputs(1006));
    outputs(6033) <= not(layer2_outputs(11611));
    outputs(6034) <= not((layer2_outputs(8167)) xor (layer2_outputs(9907)));
    outputs(6035) <= layer2_outputs(6589);
    outputs(6036) <= not(layer2_outputs(1807));
    outputs(6037) <= not(layer2_outputs(4652));
    outputs(6038) <= not((layer2_outputs(4608)) xor (layer2_outputs(5555)));
    outputs(6039) <= layer2_outputs(9380);
    outputs(6040) <= not(layer2_outputs(3906));
    outputs(6041) <= layer2_outputs(3669);
    outputs(6042) <= not(layer2_outputs(8467));
    outputs(6043) <= not((layer2_outputs(4154)) xor (layer2_outputs(4116)));
    outputs(6044) <= layer2_outputs(7927);
    outputs(6045) <= not((layer2_outputs(7427)) or (layer2_outputs(1570)));
    outputs(6046) <= not(layer2_outputs(11771)) or (layer2_outputs(3671));
    outputs(6047) <= not(layer2_outputs(7658));
    outputs(6048) <= not(layer2_outputs(11017));
    outputs(6049) <= not((layer2_outputs(7579)) xor (layer2_outputs(3913)));
    outputs(6050) <= (layer2_outputs(11529)) and (layer2_outputs(10520));
    outputs(6051) <= not(layer2_outputs(11133));
    outputs(6052) <= layer2_outputs(263);
    outputs(6053) <= layer2_outputs(7437);
    outputs(6054) <= layer2_outputs(1982);
    outputs(6055) <= layer2_outputs(6851);
    outputs(6056) <= (layer2_outputs(5883)) and (layer2_outputs(9283));
    outputs(6057) <= layer2_outputs(12597);
    outputs(6058) <= not(layer2_outputs(5032));
    outputs(6059) <= (layer2_outputs(145)) xor (layer2_outputs(12270));
    outputs(6060) <= not((layer2_outputs(1282)) xor (layer2_outputs(1280)));
    outputs(6061) <= not(layer2_outputs(590));
    outputs(6062) <= not(layer2_outputs(12716));
    outputs(6063) <= (layer2_outputs(10052)) and not (layer2_outputs(12041));
    outputs(6064) <= not(layer2_outputs(3090));
    outputs(6065) <= layer2_outputs(3896);
    outputs(6066) <= not(layer2_outputs(1370));
    outputs(6067) <= (layer2_outputs(10847)) xor (layer2_outputs(994));
    outputs(6068) <= not((layer2_outputs(2745)) xor (layer2_outputs(9549)));
    outputs(6069) <= not((layer2_outputs(8931)) xor (layer2_outputs(7244)));
    outputs(6070) <= not((layer2_outputs(9895)) xor (layer2_outputs(11705)));
    outputs(6071) <= not(layer2_outputs(3140));
    outputs(6072) <= layer2_outputs(2126);
    outputs(6073) <= not(layer2_outputs(2510));
    outputs(6074) <= (layer2_outputs(6441)) and not (layer2_outputs(6814));
    outputs(6075) <= layer2_outputs(914);
    outputs(6076) <= not((layer2_outputs(6719)) or (layer2_outputs(5682)));
    outputs(6077) <= not((layer2_outputs(10939)) xor (layer2_outputs(11472)));
    outputs(6078) <= layer2_outputs(388);
    outputs(6079) <= layer2_outputs(236);
    outputs(6080) <= not((layer2_outputs(9883)) xor (layer2_outputs(7791)));
    outputs(6081) <= (layer2_outputs(11073)) xor (layer2_outputs(11068));
    outputs(6082) <= layer2_outputs(12288);
    outputs(6083) <= (layer2_outputs(5554)) xor (layer2_outputs(154));
    outputs(6084) <= not(layer2_outputs(6090));
    outputs(6085) <= (layer2_outputs(5063)) or (layer2_outputs(7350));
    outputs(6086) <= not(layer2_outputs(4646));
    outputs(6087) <= (layer2_outputs(741)) xor (layer2_outputs(7169));
    outputs(6088) <= layer2_outputs(3761);
    outputs(6089) <= layer2_outputs(4333);
    outputs(6090) <= (layer2_outputs(7360)) xor (layer2_outputs(12525));
    outputs(6091) <= not(layer2_outputs(6205));
    outputs(6092) <= not(layer2_outputs(845));
    outputs(6093) <= layer2_outputs(9315);
    outputs(6094) <= not(layer2_outputs(788));
    outputs(6095) <= not((layer2_outputs(5498)) xor (layer2_outputs(12314)));
    outputs(6096) <= layer2_outputs(8767);
    outputs(6097) <= layer2_outputs(5778);
    outputs(6098) <= not(layer2_outputs(12271));
    outputs(6099) <= layer2_outputs(1565);
    outputs(6100) <= not(layer2_outputs(3263));
    outputs(6101) <= layer2_outputs(11080);
    outputs(6102) <= not(layer2_outputs(68));
    outputs(6103) <= layer2_outputs(394);
    outputs(6104) <= not(layer2_outputs(7079));
    outputs(6105) <= not(layer2_outputs(4845));
    outputs(6106) <= not(layer2_outputs(499));
    outputs(6107) <= not((layer2_outputs(3526)) xor (layer2_outputs(10628)));
    outputs(6108) <= not(layer2_outputs(1843));
    outputs(6109) <= layer2_outputs(8575);
    outputs(6110) <= (layer2_outputs(3276)) xor (layer2_outputs(6296));
    outputs(6111) <= layer2_outputs(10415);
    outputs(6112) <= layer2_outputs(12369);
    outputs(6113) <= not(layer2_outputs(9309));
    outputs(6114) <= not(layer2_outputs(12682));
    outputs(6115) <= not((layer2_outputs(565)) or (layer2_outputs(515)));
    outputs(6116) <= not((layer2_outputs(1994)) xor (layer2_outputs(1572)));
    outputs(6117) <= (layer2_outputs(6349)) and not (layer2_outputs(9223));
    outputs(6118) <= not((layer2_outputs(5117)) xor (layer2_outputs(5887)));
    outputs(6119) <= not((layer2_outputs(5771)) xor (layer2_outputs(5299)));
    outputs(6120) <= layer2_outputs(1127);
    outputs(6121) <= layer2_outputs(8091);
    outputs(6122) <= (layer2_outputs(8317)) or (layer2_outputs(6434));
    outputs(6123) <= not(layer2_outputs(8594));
    outputs(6124) <= (layer2_outputs(7952)) and (layer2_outputs(11679));
    outputs(6125) <= not(layer2_outputs(5927)) or (layer2_outputs(4848));
    outputs(6126) <= not((layer2_outputs(1117)) xor (layer2_outputs(8614)));
    outputs(6127) <= not(layer2_outputs(7446));
    outputs(6128) <= layer2_outputs(9370);
    outputs(6129) <= not(layer2_outputs(396));
    outputs(6130) <= (layer2_outputs(12500)) xor (layer2_outputs(8071));
    outputs(6131) <= not(layer2_outputs(52));
    outputs(6132) <= (layer2_outputs(189)) and (layer2_outputs(9282));
    outputs(6133) <= (layer2_outputs(10650)) and not (layer2_outputs(11603));
    outputs(6134) <= (layer2_outputs(4381)) xor (layer2_outputs(2163));
    outputs(6135) <= layer2_outputs(1804);
    outputs(6136) <= layer2_outputs(3693);
    outputs(6137) <= not(layer2_outputs(3330));
    outputs(6138) <= not((layer2_outputs(2039)) and (layer2_outputs(11043)));
    outputs(6139) <= layer2_outputs(964);
    outputs(6140) <= (layer2_outputs(321)) and (layer2_outputs(9552));
    outputs(6141) <= (layer2_outputs(3783)) xor (layer2_outputs(9126));
    outputs(6142) <= layer2_outputs(6349);
    outputs(6143) <= (layer2_outputs(5787)) xor (layer2_outputs(1024));
    outputs(6144) <= not((layer2_outputs(9142)) or (layer2_outputs(6788)));
    outputs(6145) <= (layer2_outputs(6174)) or (layer2_outputs(567));
    outputs(6146) <= not((layer2_outputs(12037)) or (layer2_outputs(3993)));
    outputs(6147) <= not(layer2_outputs(8338));
    outputs(6148) <= not((layer2_outputs(44)) xor (layer2_outputs(4395)));
    outputs(6149) <= (layer2_outputs(12208)) xor (layer2_outputs(209));
    outputs(6150) <= not(layer2_outputs(4108));
    outputs(6151) <= (layer2_outputs(4359)) xor (layer2_outputs(2009));
    outputs(6152) <= not((layer2_outputs(2375)) xor (layer2_outputs(824)));
    outputs(6153) <= not(layer2_outputs(512));
    outputs(6154) <= layer2_outputs(6865);
    outputs(6155) <= (layer2_outputs(3553)) or (layer2_outputs(9049));
    outputs(6156) <= not(layer2_outputs(10526));
    outputs(6157) <= layer2_outputs(2571);
    outputs(6158) <= not((layer2_outputs(6053)) xor (layer2_outputs(11142)));
    outputs(6159) <= not((layer2_outputs(8419)) or (layer2_outputs(7457)));
    outputs(6160) <= layer2_outputs(615);
    outputs(6161) <= not(layer2_outputs(1431));
    outputs(6162) <= layer2_outputs(10299);
    outputs(6163) <= not((layer2_outputs(11727)) and (layer2_outputs(12179)));
    outputs(6164) <= (layer2_outputs(8963)) xor (layer2_outputs(1660));
    outputs(6165) <= not((layer2_outputs(2547)) xor (layer2_outputs(7492)));
    outputs(6166) <= not(layer2_outputs(673)) or (layer2_outputs(515));
    outputs(6167) <= layer2_outputs(4927);
    outputs(6168) <= not(layer2_outputs(11979));
    outputs(6169) <= (layer2_outputs(12692)) xor (layer2_outputs(6516));
    outputs(6170) <= not(layer2_outputs(8396));
    outputs(6171) <= (layer2_outputs(640)) xor (layer2_outputs(9831));
    outputs(6172) <= not((layer2_outputs(9931)) and (layer2_outputs(6176)));
    outputs(6173) <= layer2_outputs(6702);
    outputs(6174) <= (layer2_outputs(11120)) xor (layer2_outputs(9776));
    outputs(6175) <= not(layer2_outputs(12477));
    outputs(6176) <= (layer2_outputs(1885)) xor (layer2_outputs(852));
    outputs(6177) <= (layer2_outputs(5798)) xor (layer2_outputs(1149));
    outputs(6178) <= not(layer2_outputs(11281));
    outputs(6179) <= (layer2_outputs(1624)) and not (layer2_outputs(9317));
    outputs(6180) <= not(layer2_outputs(4038));
    outputs(6181) <= not(layer2_outputs(12338));
    outputs(6182) <= layer2_outputs(7447);
    outputs(6183) <= not(layer2_outputs(2279));
    outputs(6184) <= layer2_outputs(9181);
    outputs(6185) <= (layer2_outputs(12566)) xor (layer2_outputs(9952));
    outputs(6186) <= (layer2_outputs(8168)) and (layer2_outputs(450));
    outputs(6187) <= layer2_outputs(4549);
    outputs(6188) <= not(layer2_outputs(8570));
    outputs(6189) <= layer2_outputs(6132);
    outputs(6190) <= not(layer2_outputs(5145)) or (layer2_outputs(2343));
    outputs(6191) <= layer2_outputs(5166);
    outputs(6192) <= not((layer2_outputs(4801)) xor (layer2_outputs(8509)));
    outputs(6193) <= not(layer2_outputs(3998));
    outputs(6194) <= not((layer2_outputs(6824)) xor (layer2_outputs(54)));
    outputs(6195) <= not((layer2_outputs(4678)) xor (layer2_outputs(1233)));
    outputs(6196) <= not(layer2_outputs(4865));
    outputs(6197) <= not(layer2_outputs(2454));
    outputs(6198) <= not((layer2_outputs(7751)) or (layer2_outputs(7090)));
    outputs(6199) <= not(layer2_outputs(6715));
    outputs(6200) <= not(layer2_outputs(11661));
    outputs(6201) <= not(layer2_outputs(5519));
    outputs(6202) <= not(layer2_outputs(5444)) or (layer2_outputs(5358));
    outputs(6203) <= (layer2_outputs(11331)) xor (layer2_outputs(8805));
    outputs(6204) <= not(layer2_outputs(1249));
    outputs(6205) <= not(layer2_outputs(3724));
    outputs(6206) <= layer2_outputs(7275);
    outputs(6207) <= not(layer2_outputs(4321));
    outputs(6208) <= (layer2_outputs(8661)) and (layer2_outputs(8957));
    outputs(6209) <= not((layer2_outputs(561)) xor (layer2_outputs(5772)));
    outputs(6210) <= not(layer2_outputs(652));
    outputs(6211) <= layer2_outputs(1206);
    outputs(6212) <= (layer2_outputs(2125)) xor (layer2_outputs(12674));
    outputs(6213) <= layer2_outputs(11989);
    outputs(6214) <= layer2_outputs(806);
    outputs(6215) <= not(layer2_outputs(11967));
    outputs(6216) <= not(layer2_outputs(847));
    outputs(6217) <= not(layer2_outputs(5565));
    outputs(6218) <= (layer2_outputs(8605)) xor (layer2_outputs(7049));
    outputs(6219) <= (layer2_outputs(4813)) xor (layer2_outputs(4062));
    outputs(6220) <= not(layer2_outputs(6586));
    outputs(6221) <= not((layer2_outputs(4615)) xor (layer2_outputs(9728)));
    outputs(6222) <= not(layer2_outputs(11706));
    outputs(6223) <= layer2_outputs(12218);
    outputs(6224) <= not(layer2_outputs(6357));
    outputs(6225) <= (layer2_outputs(11239)) xor (layer2_outputs(8178));
    outputs(6226) <= layer2_outputs(9353);
    outputs(6227) <= layer2_outputs(9265);
    outputs(6228) <= not(layer2_outputs(6431));
    outputs(6229) <= layer2_outputs(4111);
    outputs(6230) <= layer2_outputs(6203);
    outputs(6231) <= not((layer2_outputs(10575)) and (layer2_outputs(4241)));
    outputs(6232) <= (layer2_outputs(9503)) or (layer2_outputs(3653));
    outputs(6233) <= not(layer2_outputs(4254));
    outputs(6234) <= not(layer2_outputs(11233));
    outputs(6235) <= not(layer2_outputs(11125));
    outputs(6236) <= layer2_outputs(1439);
    outputs(6237) <= not(layer2_outputs(8063));
    outputs(6238) <= not(layer2_outputs(5418)) or (layer2_outputs(1911));
    outputs(6239) <= layer2_outputs(9857);
    outputs(6240) <= not((layer2_outputs(10100)) xor (layer2_outputs(12562)));
    outputs(6241) <= not(layer2_outputs(3186));
    outputs(6242) <= not(layer2_outputs(11000)) or (layer2_outputs(2900));
    outputs(6243) <= not(layer2_outputs(10160));
    outputs(6244) <= not((layer2_outputs(160)) or (layer2_outputs(9776)));
    outputs(6245) <= not((layer2_outputs(10343)) or (layer2_outputs(4098)));
    outputs(6246) <= not(layer2_outputs(8228));
    outputs(6247) <= not(layer2_outputs(6284));
    outputs(6248) <= (layer2_outputs(12044)) xor (layer2_outputs(4489));
    outputs(6249) <= (layer2_outputs(5037)) xor (layer2_outputs(4879));
    outputs(6250) <= not(layer2_outputs(2816));
    outputs(6251) <= not((layer2_outputs(9158)) and (layer2_outputs(6792)));
    outputs(6252) <= layer2_outputs(2005);
    outputs(6253) <= layer2_outputs(7587);
    outputs(6254) <= not((layer2_outputs(3658)) xor (layer2_outputs(7946)));
    outputs(6255) <= (layer2_outputs(5857)) xor (layer2_outputs(6578));
    outputs(6256) <= layer2_outputs(8759);
    outputs(6257) <= (layer2_outputs(2144)) or (layer2_outputs(6260));
    outputs(6258) <= layer2_outputs(7933);
    outputs(6259) <= not((layer2_outputs(7436)) xor (layer2_outputs(410)));
    outputs(6260) <= not(layer2_outputs(7359));
    outputs(6261) <= not(layer2_outputs(6326));
    outputs(6262) <= layer2_outputs(9457);
    outputs(6263) <= (layer2_outputs(2558)) xor (layer2_outputs(10562));
    outputs(6264) <= not((layer2_outputs(4914)) xor (layer2_outputs(141)));
    outputs(6265) <= not(layer2_outputs(4940));
    outputs(6266) <= not((layer2_outputs(968)) xor (layer2_outputs(5955)));
    outputs(6267) <= not(layer2_outputs(10934));
    outputs(6268) <= not(layer2_outputs(8396));
    outputs(6269) <= layer2_outputs(6107);
    outputs(6270) <= layer2_outputs(9057);
    outputs(6271) <= layer2_outputs(8831);
    outputs(6272) <= not(layer2_outputs(6419)) or (layer2_outputs(11675));
    outputs(6273) <= (layer2_outputs(2517)) xor (layer2_outputs(3580));
    outputs(6274) <= not(layer2_outputs(7538));
    outputs(6275) <= (layer2_outputs(631)) and not (layer2_outputs(9626));
    outputs(6276) <= not((layer2_outputs(9258)) xor (layer2_outputs(11446)));
    outputs(6277) <= layer2_outputs(11567);
    outputs(6278) <= not((layer2_outputs(9612)) and (layer2_outputs(11397)));
    outputs(6279) <= not(layer2_outputs(11168));
    outputs(6280) <= (layer2_outputs(8953)) and not (layer2_outputs(11236));
    outputs(6281) <= not(layer2_outputs(5331));
    outputs(6282) <= not(layer2_outputs(9284));
    outputs(6283) <= (layer2_outputs(3009)) xor (layer2_outputs(5712));
    outputs(6284) <= layer2_outputs(6770);
    outputs(6285) <= not((layer2_outputs(6449)) xor (layer2_outputs(8592)));
    outputs(6286) <= layer2_outputs(1108);
    outputs(6287) <= (layer2_outputs(8435)) xor (layer2_outputs(552));
    outputs(6288) <= (layer2_outputs(10873)) xor (layer2_outputs(5158));
    outputs(6289) <= not((layer2_outputs(5864)) or (layer2_outputs(2889)));
    outputs(6290) <= (layer2_outputs(8881)) xor (layer2_outputs(10063));
    outputs(6291) <= not(layer2_outputs(11286));
    outputs(6292) <= layer2_outputs(7673);
    outputs(6293) <= (layer2_outputs(5600)) xor (layer2_outputs(3454));
    outputs(6294) <= layer2_outputs(2887);
    outputs(6295) <= not((layer2_outputs(9663)) xor (layer2_outputs(10061)));
    outputs(6296) <= (layer2_outputs(9714)) or (layer2_outputs(3766));
    outputs(6297) <= layer2_outputs(10423);
    outputs(6298) <= (layer2_outputs(12361)) xor (layer2_outputs(9039));
    outputs(6299) <= layer2_outputs(5063);
    outputs(6300) <= not(layer2_outputs(5236));
    outputs(6301) <= layer2_outputs(6961);
    outputs(6302) <= (layer2_outputs(11381)) xor (layer2_outputs(6533));
    outputs(6303) <= layer2_outputs(5176);
    outputs(6304) <= not(layer2_outputs(3517));
    outputs(6305) <= not(layer2_outputs(11890));
    outputs(6306) <= not(layer2_outputs(9635));
    outputs(6307) <= not(layer2_outputs(1445));
    outputs(6308) <= not(layer2_outputs(47));
    outputs(6309) <= (layer2_outputs(12272)) or (layer2_outputs(7315));
    outputs(6310) <= not((layer2_outputs(6657)) xor (layer2_outputs(6747)));
    outputs(6311) <= layer2_outputs(9716);
    outputs(6312) <= not(layer2_outputs(9295));
    outputs(6313) <= layer2_outputs(3992);
    outputs(6314) <= not((layer2_outputs(11697)) xor (layer2_outputs(5825)));
    outputs(6315) <= not((layer2_outputs(1950)) xor (layer2_outputs(2864)));
    outputs(6316) <= not(layer2_outputs(1036));
    outputs(6317) <= layer2_outputs(11954);
    outputs(6318) <= not((layer2_outputs(10352)) xor (layer2_outputs(6122)));
    outputs(6319) <= not(layer2_outputs(8353));
    outputs(6320) <= not((layer2_outputs(7455)) or (layer2_outputs(9025)));
    outputs(6321) <= (layer2_outputs(3084)) xor (layer2_outputs(10653));
    outputs(6322) <= (layer2_outputs(5945)) xor (layer2_outputs(3042));
    outputs(6323) <= layer2_outputs(5438);
    outputs(6324) <= not(layer2_outputs(5488)) or (layer2_outputs(8978));
    outputs(6325) <= layer2_outputs(5633);
    outputs(6326) <= not(layer2_outputs(644));
    outputs(6327) <= layer2_outputs(8037);
    outputs(6328) <= layer2_outputs(5352);
    outputs(6329) <= layer2_outputs(12489);
    outputs(6330) <= (layer2_outputs(5092)) and not (layer2_outputs(11659));
    outputs(6331) <= not((layer2_outputs(7401)) xor (layer2_outputs(7011)));
    outputs(6332) <= not((layer2_outputs(893)) xor (layer2_outputs(8592)));
    outputs(6333) <= not((layer2_outputs(4165)) xor (layer2_outputs(2766)));
    outputs(6334) <= not(layer2_outputs(4764));
    outputs(6335) <= not(layer2_outputs(3339));
    outputs(6336) <= not(layer2_outputs(9163));
    outputs(6337) <= (layer2_outputs(2311)) xor (layer2_outputs(2028));
    outputs(6338) <= not(layer2_outputs(4355));
    outputs(6339) <= not(layer2_outputs(10956));
    outputs(6340) <= (layer2_outputs(7667)) and not (layer2_outputs(1657));
    outputs(6341) <= layer2_outputs(1818);
    outputs(6342) <= not((layer2_outputs(5569)) xor (layer2_outputs(4291)));
    outputs(6343) <= not(layer2_outputs(66));
    outputs(6344) <= not(layer2_outputs(1015));
    outputs(6345) <= not((layer2_outputs(10030)) xor (layer2_outputs(7622)));
    outputs(6346) <= (layer2_outputs(3413)) xor (layer2_outputs(2304));
    outputs(6347) <= not(layer2_outputs(1014));
    outputs(6348) <= (layer2_outputs(5608)) xor (layer2_outputs(2433));
    outputs(6349) <= not(layer2_outputs(6765));
    outputs(6350) <= layer2_outputs(7338);
    outputs(6351) <= (layer2_outputs(4335)) and (layer2_outputs(8646));
    outputs(6352) <= not(layer2_outputs(1934));
    outputs(6353) <= not(layer2_outputs(5623));
    outputs(6354) <= not(layer2_outputs(12438));
    outputs(6355) <= (layer2_outputs(4690)) xor (layer2_outputs(11368));
    outputs(6356) <= not((layer2_outputs(6663)) xor (layer2_outputs(5516)));
    outputs(6357) <= not(layer2_outputs(10963));
    outputs(6358) <= (layer2_outputs(12134)) xor (layer2_outputs(9091));
    outputs(6359) <= not(layer2_outputs(5613)) or (layer2_outputs(3233));
    outputs(6360) <= layer2_outputs(4710);
    outputs(6361) <= layer2_outputs(6660);
    outputs(6362) <= not(layer2_outputs(4068));
    outputs(6363) <= layer2_outputs(7804);
    outputs(6364) <= layer2_outputs(5748);
    outputs(6365) <= not((layer2_outputs(11408)) xor (layer2_outputs(11172)));
    outputs(6366) <= not(layer2_outputs(10464));
    outputs(6367) <= layer2_outputs(2425);
    outputs(6368) <= not(layer2_outputs(6731));
    outputs(6369) <= not(layer2_outputs(6276));
    outputs(6370) <= not(layer2_outputs(1081));
    outputs(6371) <= (layer2_outputs(835)) and not (layer2_outputs(1783));
    outputs(6372) <= layer2_outputs(400);
    outputs(6373) <= layer2_outputs(6485);
    outputs(6374) <= layer2_outputs(8900);
    outputs(6375) <= not(layer2_outputs(8827));
    outputs(6376) <= not(layer2_outputs(1536));
    outputs(6377) <= (layer2_outputs(12734)) xor (layer2_outputs(7276));
    outputs(6378) <= not(layer2_outputs(1158));
    outputs(6379) <= layer2_outputs(4495);
    outputs(6380) <= (layer2_outputs(9875)) xor (layer2_outputs(12154));
    outputs(6381) <= layer2_outputs(2246);
    outputs(6382) <= (layer2_outputs(4753)) or (layer2_outputs(12647));
    outputs(6383) <= not((layer2_outputs(10564)) xor (layer2_outputs(11296)));
    outputs(6384) <= layer2_outputs(3803);
    outputs(6385) <= layer2_outputs(7061);
    outputs(6386) <= layer2_outputs(1169);
    outputs(6387) <= not((layer2_outputs(9484)) xor (layer2_outputs(3930)));
    outputs(6388) <= not(layer2_outputs(2991));
    outputs(6389) <= layer2_outputs(10913);
    outputs(6390) <= layer2_outputs(8832);
    outputs(6391) <= layer2_outputs(5103);
    outputs(6392) <= not(layer2_outputs(12184)) or (layer2_outputs(12270));
    outputs(6393) <= not(layer2_outputs(1308));
    outputs(6394) <= not((layer2_outputs(7853)) xor (layer2_outputs(3869)));
    outputs(6395) <= layer2_outputs(11826);
    outputs(6396) <= (layer2_outputs(11448)) and not (layer2_outputs(5837));
    outputs(6397) <= not(layer2_outputs(6840));
    outputs(6398) <= not((layer2_outputs(9559)) or (layer2_outputs(5252)));
    outputs(6399) <= not((layer2_outputs(1763)) xor (layer2_outputs(1450)));
    outputs(6400) <= layer2_outputs(2104);
    outputs(6401) <= (layer2_outputs(9557)) or (layer2_outputs(105));
    outputs(6402) <= not(layer2_outputs(12415));
    outputs(6403) <= layer2_outputs(8565);
    outputs(6404) <= layer2_outputs(4686);
    outputs(6405) <= layer2_outputs(9317);
    outputs(6406) <= not((layer2_outputs(11857)) and (layer2_outputs(7050)));
    outputs(6407) <= (layer2_outputs(4325)) xor (layer2_outputs(5371));
    outputs(6408) <= not(layer2_outputs(7410));
    outputs(6409) <= layer2_outputs(1382);
    outputs(6410) <= not((layer2_outputs(10852)) xor (layer2_outputs(11970)));
    outputs(6411) <= not(layer2_outputs(2054));
    outputs(6412) <= layer2_outputs(8161);
    outputs(6413) <= not(layer2_outputs(12226));
    outputs(6414) <= not((layer2_outputs(12340)) xor (layer2_outputs(7630)));
    outputs(6415) <= not(layer2_outputs(11192));
    outputs(6416) <= not((layer2_outputs(12189)) xor (layer2_outputs(4408)));
    outputs(6417) <= not(layer2_outputs(3385));
    outputs(6418) <= not(layer2_outputs(11225));
    outputs(6419) <= not(layer2_outputs(9444));
    outputs(6420) <= (layer2_outputs(8006)) xor (layer2_outputs(8547));
    outputs(6421) <= (layer2_outputs(8882)) xor (layer2_outputs(5386));
    outputs(6422) <= not(layer2_outputs(7467));
    outputs(6423) <= layer2_outputs(8990);
    outputs(6424) <= not(layer2_outputs(3170));
    outputs(6425) <= layer2_outputs(4764);
    outputs(6426) <= not((layer2_outputs(873)) or (layer2_outputs(11970)));
    outputs(6427) <= not(layer2_outputs(10390)) or (layer2_outputs(8216));
    outputs(6428) <= layer2_outputs(974);
    outputs(6429) <= not(layer2_outputs(3743));
    outputs(6430) <= layer2_outputs(6827);
    outputs(6431) <= not(layer2_outputs(10543));
    outputs(6432) <= layer2_outputs(11742);
    outputs(6433) <= not(layer2_outputs(10800));
    outputs(6434) <= not((layer2_outputs(107)) xor (layer2_outputs(3160)));
    outputs(6435) <= layer2_outputs(6796);
    outputs(6436) <= (layer2_outputs(3592)) and not (layer2_outputs(3664));
    outputs(6437) <= not((layer2_outputs(1402)) xor (layer2_outputs(1956)));
    outputs(6438) <= not((layer2_outputs(8107)) xor (layer2_outputs(7450)));
    outputs(6439) <= not(layer2_outputs(5822)) or (layer2_outputs(9633));
    outputs(6440) <= not(layer2_outputs(8495));
    outputs(6441) <= (layer2_outputs(9114)) and not (layer2_outputs(1750));
    outputs(6442) <= layer2_outputs(9280);
    outputs(6443) <= not((layer2_outputs(7500)) and (layer2_outputs(1124)));
    outputs(6444) <= not(layer2_outputs(2051)) or (layer2_outputs(3522));
    outputs(6445) <= not(layer2_outputs(2003));
    outputs(6446) <= (layer2_outputs(10653)) xor (layer2_outputs(10457));
    outputs(6447) <= not(layer2_outputs(4632));
    outputs(6448) <= (layer2_outputs(5811)) xor (layer2_outputs(11332));
    outputs(6449) <= layer2_outputs(12103);
    outputs(6450) <= not((layer2_outputs(8194)) xor (layer2_outputs(6249)));
    outputs(6451) <= layer2_outputs(9418);
    outputs(6452) <= not(layer2_outputs(9537));
    outputs(6453) <= not(layer2_outputs(11116));
    outputs(6454) <= not(layer2_outputs(2774));
    outputs(6455) <= layer2_outputs(8820);
    outputs(6456) <= layer2_outputs(8321);
    outputs(6457) <= not((layer2_outputs(12354)) xor (layer2_outputs(2617)));
    outputs(6458) <= layer2_outputs(486);
    outputs(6459) <= layer2_outputs(7010);
    outputs(6460) <= (layer2_outputs(5381)) xor (layer2_outputs(8083));
    outputs(6461) <= layer2_outputs(11959);
    outputs(6462) <= not(layer2_outputs(4920));
    outputs(6463) <= layer2_outputs(2229);
    outputs(6464) <= layer2_outputs(5279);
    outputs(6465) <= not(layer2_outputs(9971)) or (layer2_outputs(10325));
    outputs(6466) <= not((layer2_outputs(2143)) xor (layer2_outputs(1099)));
    outputs(6467) <= (layer2_outputs(1416)) and (layer2_outputs(1429));
    outputs(6468) <= not((layer2_outputs(6811)) xor (layer2_outputs(11868)));
    outputs(6469) <= not(layer2_outputs(9575));
    outputs(6470) <= layer2_outputs(5892);
    outputs(6471) <= (layer2_outputs(4417)) xor (layer2_outputs(501));
    outputs(6472) <= not(layer2_outputs(1494));
    outputs(6473) <= (layer2_outputs(6156)) and (layer2_outputs(8313));
    outputs(6474) <= not(layer2_outputs(3779));
    outputs(6475) <= not((layer2_outputs(9162)) xor (layer2_outputs(10502)));
    outputs(6476) <= layer2_outputs(5423);
    outputs(6477) <= (layer2_outputs(9574)) xor (layer2_outputs(10604));
    outputs(6478) <= (layer2_outputs(8379)) xor (layer2_outputs(12702));
    outputs(6479) <= layer2_outputs(908);
    outputs(6480) <= not(layer2_outputs(12126));
    outputs(6481) <= layer2_outputs(669);
    outputs(6482) <= not(layer2_outputs(2514));
    outputs(6483) <= not((layer2_outputs(3830)) xor (layer2_outputs(11925)));
    outputs(6484) <= (layer2_outputs(10869)) or (layer2_outputs(5478));
    outputs(6485) <= (layer2_outputs(6617)) xor (layer2_outputs(7716));
    outputs(6486) <= not(layer2_outputs(281)) or (layer2_outputs(11389));
    outputs(6487) <= layer2_outputs(11490);
    outputs(6488) <= not(layer2_outputs(10379));
    outputs(6489) <= layer2_outputs(9043);
    outputs(6490) <= not((layer2_outputs(2274)) xor (layer2_outputs(2)));
    outputs(6491) <= not(layer2_outputs(11252));
    outputs(6492) <= layer2_outputs(3382);
    outputs(6493) <= not(layer2_outputs(12040));
    outputs(6494) <= layer2_outputs(1628);
    outputs(6495) <= not((layer2_outputs(2392)) xor (layer2_outputs(1817)));
    outputs(6496) <= layer2_outputs(9274);
    outputs(6497) <= not((layer2_outputs(8021)) and (layer2_outputs(6925)));
    outputs(6498) <= not(layer2_outputs(12586));
    outputs(6499) <= (layer2_outputs(11781)) and not (layer2_outputs(5911));
    outputs(6500) <= not(layer2_outputs(3795));
    outputs(6501) <= not(layer2_outputs(8686));
    outputs(6502) <= layer2_outputs(1512);
    outputs(6503) <= not((layer2_outputs(12170)) xor (layer2_outputs(1468)));
    outputs(6504) <= (layer2_outputs(3777)) and not (layer2_outputs(5130));
    outputs(6505) <= layer2_outputs(4936);
    outputs(6506) <= not((layer2_outputs(1605)) xor (layer2_outputs(9545)));
    outputs(6507) <= layer2_outputs(7190);
    outputs(6508) <= layer2_outputs(2199);
    outputs(6509) <= layer2_outputs(1661);
    outputs(6510) <= layer2_outputs(315);
    outputs(6511) <= layer2_outputs(6823);
    outputs(6512) <= layer2_outputs(4313);
    outputs(6513) <= (layer2_outputs(3299)) xor (layer2_outputs(2040));
    outputs(6514) <= (layer2_outputs(7903)) and not (layer2_outputs(7329));
    outputs(6515) <= not((layer2_outputs(4996)) and (layer2_outputs(9665)));
    outputs(6516) <= layer2_outputs(11095);
    outputs(6517) <= layer2_outputs(6316);
    outputs(6518) <= not((layer2_outputs(10622)) xor (layer2_outputs(1456)));
    outputs(6519) <= not(layer2_outputs(6382));
    outputs(6520) <= not((layer2_outputs(8390)) xor (layer2_outputs(5027)));
    outputs(6521) <= not(layer2_outputs(7329));
    outputs(6522) <= layer2_outputs(6833);
    outputs(6523) <= not(layer2_outputs(11164));
    outputs(6524) <= not((layer2_outputs(5148)) xor (layer2_outputs(7181)));
    outputs(6525) <= not((layer2_outputs(4146)) xor (layer2_outputs(1000)));
    outputs(6526) <= layer2_outputs(6223);
    outputs(6527) <= (layer2_outputs(10364)) or (layer2_outputs(8094));
    outputs(6528) <= not(layer2_outputs(10507));
    outputs(6529) <= not(layer2_outputs(10025)) or (layer2_outputs(4391));
    outputs(6530) <= not(layer2_outputs(8817)) or (layer2_outputs(11251));
    outputs(6531) <= not((layer2_outputs(10829)) xor (layer2_outputs(3769)));
    outputs(6532) <= not(layer2_outputs(9167));
    outputs(6533) <= not((layer2_outputs(3855)) xor (layer2_outputs(9852)));
    outputs(6534) <= layer2_outputs(3241);
    outputs(6535) <= (layer2_outputs(2063)) and (layer2_outputs(10932));
    outputs(6536) <= not((layer2_outputs(3450)) xor (layer2_outputs(4402)));
    outputs(6537) <= not((layer2_outputs(4487)) xor (layer2_outputs(845)));
    outputs(6538) <= not(layer2_outputs(5012));
    outputs(6539) <= layer2_outputs(1102);
    outputs(6540) <= (layer2_outputs(5697)) xor (layer2_outputs(4046));
    outputs(6541) <= layer2_outputs(8889);
    outputs(6542) <= not(layer2_outputs(2027));
    outputs(6543) <= (layer2_outputs(3288)) xor (layer2_outputs(5813));
    outputs(6544) <= (layer2_outputs(3836)) and not (layer2_outputs(6071));
    outputs(6545) <= not(layer2_outputs(11869)) or (layer2_outputs(7058));
    outputs(6546) <= layer2_outputs(7367);
    outputs(6547) <= layer2_outputs(245);
    outputs(6548) <= not(layer2_outputs(2774));
    outputs(6549) <= (layer2_outputs(1027)) xor (layer2_outputs(12721));
    outputs(6550) <= layer2_outputs(654);
    outputs(6551) <= not(layer2_outputs(1910));
    outputs(6552) <= (layer2_outputs(2238)) xor (layer2_outputs(12484));
    outputs(6553) <= layer2_outputs(1121);
    outputs(6554) <= not(layer2_outputs(7341));
    outputs(6555) <= (layer2_outputs(5747)) and not (layer2_outputs(1417));
    outputs(6556) <= not(layer2_outputs(10343)) or (layer2_outputs(9315));
    outputs(6557) <= (layer2_outputs(640)) xor (layer2_outputs(9059));
    outputs(6558) <= layer2_outputs(9671);
    outputs(6559) <= not(layer2_outputs(8954));
    outputs(6560) <= not(layer2_outputs(11482));
    outputs(6561) <= not(layer2_outputs(6327));
    outputs(6562) <= not(layer2_outputs(12024));
    outputs(6563) <= not(layer2_outputs(950));
    outputs(6564) <= layer2_outputs(7665);
    outputs(6565) <= not(layer2_outputs(1322));
    outputs(6566) <= not(layer2_outputs(3675));
    outputs(6567) <= (layer2_outputs(229)) xor (layer2_outputs(3781));
    outputs(6568) <= not(layer2_outputs(134));
    outputs(6569) <= not(layer2_outputs(9352)) or (layer2_outputs(11114));
    outputs(6570) <= layer2_outputs(7232);
    outputs(6571) <= not((layer2_outputs(1923)) xor (layer2_outputs(9227)));
    outputs(6572) <= not(layer2_outputs(987));
    outputs(6573) <= layer2_outputs(11800);
    outputs(6574) <= layer2_outputs(10761);
    outputs(6575) <= not((layer2_outputs(8547)) xor (layer2_outputs(10064)));
    outputs(6576) <= not(layer2_outputs(1153)) or (layer2_outputs(10310));
    outputs(6577) <= layer2_outputs(4262);
    outputs(6578) <= layer2_outputs(10164);
    outputs(6579) <= (layer2_outputs(9851)) xor (layer2_outputs(755));
    outputs(6580) <= layer2_outputs(1245);
    outputs(6581) <= not(layer2_outputs(1577));
    outputs(6582) <= not((layer2_outputs(5421)) xor (layer2_outputs(2856)));
    outputs(6583) <= layer2_outputs(5640);
    outputs(6584) <= layer2_outputs(5275);
    outputs(6585) <= (layer2_outputs(1579)) xor (layer2_outputs(6764));
    outputs(6586) <= not(layer2_outputs(2832));
    outputs(6587) <= (layer2_outputs(12737)) xor (layer2_outputs(9254));
    outputs(6588) <= (layer2_outputs(7479)) xor (layer2_outputs(9396));
    outputs(6589) <= layer2_outputs(5301);
    outputs(6590) <= not(layer2_outputs(11833));
    outputs(6591) <= (layer2_outputs(10094)) and not (layer2_outputs(4996));
    outputs(6592) <= (layer2_outputs(9386)) xor (layer2_outputs(6734));
    outputs(6593) <= (layer2_outputs(7978)) xor (layer2_outputs(5363));
    outputs(6594) <= not((layer2_outputs(10756)) xor (layer2_outputs(2144)));
    outputs(6595) <= not((layer2_outputs(3126)) xor (layer2_outputs(605)));
    outputs(6596) <= layer2_outputs(5738);
    outputs(6597) <= layer2_outputs(2378);
    outputs(6598) <= not(layer2_outputs(10507));
    outputs(6599) <= (layer2_outputs(8895)) xor (layer2_outputs(50));
    outputs(6600) <= not(layer2_outputs(11817));
    outputs(6601) <= (layer2_outputs(9113)) xor (layer2_outputs(3060));
    outputs(6602) <= (layer2_outputs(1948)) and not (layer2_outputs(12159));
    outputs(6603) <= layer2_outputs(3472);
    outputs(6604) <= (layer2_outputs(3347)) xor (layer2_outputs(868));
    outputs(6605) <= (layer2_outputs(5889)) xor (layer2_outputs(4366));
    outputs(6606) <= (layer2_outputs(8424)) and (layer2_outputs(8149));
    outputs(6607) <= (layer2_outputs(7206)) xor (layer2_outputs(1413));
    outputs(6608) <= layer2_outputs(4466);
    outputs(6609) <= layer2_outputs(8425);
    outputs(6610) <= (layer2_outputs(10108)) xor (layer2_outputs(3722));
    outputs(6611) <= not(layer2_outputs(6073));
    outputs(6612) <= not(layer2_outputs(12061));
    outputs(6613) <= layer2_outputs(10394);
    outputs(6614) <= layer2_outputs(7001);
    outputs(6615) <= layer2_outputs(7015);
    outputs(6616) <= not(layer2_outputs(6970));
    outputs(6617) <= not((layer2_outputs(10664)) or (layer2_outputs(6075)));
    outputs(6618) <= layer2_outputs(9532);
    outputs(6619) <= (layer2_outputs(128)) xor (layer2_outputs(6260));
    outputs(6620) <= not((layer2_outputs(5535)) or (layer2_outputs(5635)));
    outputs(6621) <= (layer2_outputs(11919)) or (layer2_outputs(2815));
    outputs(6622) <= (layer2_outputs(3370)) and (layer2_outputs(12122));
    outputs(6623) <= not(layer2_outputs(2768));
    outputs(6624) <= not(layer2_outputs(3668));
    outputs(6625) <= (layer2_outputs(3460)) xor (layer2_outputs(6949));
    outputs(6626) <= (layer2_outputs(9200)) or (layer2_outputs(11777));
    outputs(6627) <= not(layer2_outputs(4884));
    outputs(6628) <= layer2_outputs(9155);
    outputs(6629) <= (layer2_outputs(12364)) xor (layer2_outputs(7660));
    outputs(6630) <= not(layer2_outputs(2064));
    outputs(6631) <= layer2_outputs(7687);
    outputs(6632) <= layer2_outputs(9551);
    outputs(6633) <= not(layer2_outputs(17));
    outputs(6634) <= layer2_outputs(7037);
    outputs(6635) <= layer2_outputs(11943);
    outputs(6636) <= (layer2_outputs(7792)) and not (layer2_outputs(8382));
    outputs(6637) <= layer2_outputs(8484);
    outputs(6638) <= not(layer2_outputs(3210)) or (layer2_outputs(0));
    outputs(6639) <= (layer2_outputs(4506)) and (layer2_outputs(7153));
    outputs(6640) <= not((layer2_outputs(3541)) and (layer2_outputs(2520)));
    outputs(6641) <= not((layer2_outputs(9099)) or (layer2_outputs(3289)));
    outputs(6642) <= layer2_outputs(10860);
    outputs(6643) <= (layer2_outputs(2595)) xor (layer2_outputs(7195));
    outputs(6644) <= (layer2_outputs(11754)) xor (layer2_outputs(8993));
    outputs(6645) <= not((layer2_outputs(1135)) xor (layer2_outputs(6957)));
    outputs(6646) <= (layer2_outputs(7380)) xor (layer2_outputs(5390));
    outputs(6647) <= not(layer2_outputs(5416)) or (layer2_outputs(9483));
    outputs(6648) <= layer2_outputs(10843);
    outputs(6649) <= not(layer2_outputs(1035));
    outputs(6650) <= layer2_outputs(4691);
    outputs(6651) <= not(layer2_outputs(10033));
    outputs(6652) <= not((layer2_outputs(4485)) and (layer2_outputs(10894)));
    outputs(6653) <= not(layer2_outputs(4275));
    outputs(6654) <= not((layer2_outputs(6613)) xor (layer2_outputs(1360)));
    outputs(6655) <= layer2_outputs(10223);
    outputs(6656) <= layer2_outputs(2415);
    outputs(6657) <= not(layer2_outputs(10664));
    outputs(6658) <= not(layer2_outputs(2951));
    outputs(6659) <= not(layer2_outputs(3437));
    outputs(6660) <= layer2_outputs(7741);
    outputs(6661) <= not(layer2_outputs(2643));
    outputs(6662) <= layer2_outputs(3904);
    outputs(6663) <= layer2_outputs(10339);
    outputs(6664) <= (layer2_outputs(9243)) and (layer2_outputs(5874));
    outputs(6665) <= (layer2_outputs(4158)) xor (layer2_outputs(9173));
    outputs(6666) <= not(layer2_outputs(9849)) or (layer2_outputs(6002));
    outputs(6667) <= layer2_outputs(11352);
    outputs(6668) <= layer2_outputs(867);
    outputs(6669) <= (layer2_outputs(11718)) xor (layer2_outputs(6146));
    outputs(6670) <= layer2_outputs(9191);
    outputs(6671) <= layer2_outputs(11451);
    outputs(6672) <= not((layer2_outputs(5224)) xor (layer2_outputs(12305)));
    outputs(6673) <= not((layer2_outputs(4183)) or (layer2_outputs(9541)));
    outputs(6674) <= (layer2_outputs(11536)) xor (layer2_outputs(3013));
    outputs(6675) <= (layer2_outputs(3061)) and not (layer2_outputs(9294));
    outputs(6676) <= (layer2_outputs(11729)) xor (layer2_outputs(1286));
    outputs(6677) <= layer2_outputs(10611);
    outputs(6678) <= layer2_outputs(2677);
    outputs(6679) <= layer2_outputs(7862);
    outputs(6680) <= not((layer2_outputs(1076)) xor (layer2_outputs(12707)));
    outputs(6681) <= not(layer2_outputs(5228));
    outputs(6682) <= not(layer2_outputs(625)) or (layer2_outputs(9400));
    outputs(6683) <= layer2_outputs(3610);
    outputs(6684) <= (layer2_outputs(7433)) xor (layer2_outputs(2596));
    outputs(6685) <= (layer2_outputs(1983)) and (layer2_outputs(1476));
    outputs(6686) <= not(layer2_outputs(4437));
    outputs(6687) <= not(layer2_outputs(2916));
    outputs(6688) <= layer2_outputs(4257);
    outputs(6689) <= not((layer2_outputs(15)) xor (layer2_outputs(3945)));
    outputs(6690) <= (layer2_outputs(10706)) xor (layer2_outputs(6901));
    outputs(6691) <= not(layer2_outputs(3400));
    outputs(6692) <= not(layer2_outputs(844));
    outputs(6693) <= not(layer2_outputs(1738));
    outputs(6694) <= (layer2_outputs(1711)) and not (layer2_outputs(12083));
    outputs(6695) <= not(layer2_outputs(5887));
    outputs(6696) <= not((layer2_outputs(12240)) or (layer2_outputs(5477)));
    outputs(6697) <= layer2_outputs(4229);
    outputs(6698) <= (layer2_outputs(12436)) and not (layer2_outputs(9708));
    outputs(6699) <= not(layer2_outputs(12388));
    outputs(6700) <= (layer2_outputs(4051)) xor (layer2_outputs(2941));
    outputs(6701) <= (layer2_outputs(6495)) xor (layer2_outputs(2814));
    outputs(6702) <= (layer2_outputs(5789)) xor (layer2_outputs(3245));
    outputs(6703) <= layer2_outputs(4578);
    outputs(6704) <= not((layer2_outputs(4836)) xor (layer2_outputs(1018)));
    outputs(6705) <= not(layer2_outputs(5410));
    outputs(6706) <= not(layer2_outputs(2294));
    outputs(6707) <= layer2_outputs(9520);
    outputs(6708) <= not((layer2_outputs(11071)) and (layer2_outputs(1180)));
    outputs(6709) <= (layer2_outputs(6152)) xor (layer2_outputs(11349));
    outputs(6710) <= layer2_outputs(9940);
    outputs(6711) <= (layer2_outputs(6959)) and not (layer2_outputs(3697));
    outputs(6712) <= (layer2_outputs(4342)) xor (layer2_outputs(4900));
    outputs(6713) <= not((layer2_outputs(4297)) xor (layer2_outputs(4574)));
    outputs(6714) <= not((layer2_outputs(3008)) xor (layer2_outputs(12350)));
    outputs(6715) <= not(layer2_outputs(5475));
    outputs(6716) <= (layer2_outputs(3168)) xor (layer2_outputs(12010));
    outputs(6717) <= layer2_outputs(4089);
    outputs(6718) <= (layer2_outputs(1878)) and not (layer2_outputs(526));
    outputs(6719) <= layer2_outputs(1901);
    outputs(6720) <= not((layer2_outputs(8512)) xor (layer2_outputs(9262)));
    outputs(6721) <= layer2_outputs(2065);
    outputs(6722) <= not(layer2_outputs(10571));
    outputs(6723) <= not((layer2_outputs(3363)) xor (layer2_outputs(1133)));
    outputs(6724) <= not(layer2_outputs(1492));
    outputs(6725) <= not(layer2_outputs(10567));
    outputs(6726) <= not(layer2_outputs(4865));
    outputs(6727) <= (layer2_outputs(3338)) or (layer2_outputs(1653));
    outputs(6728) <= layer2_outputs(9968);
    outputs(6729) <= not((layer2_outputs(11680)) xor (layer2_outputs(3447)));
    outputs(6730) <= not(layer2_outputs(3166));
    outputs(6731) <= not(layer2_outputs(2423));
    outputs(6732) <= (layer2_outputs(5882)) and not (layer2_outputs(12724));
    outputs(6733) <= (layer2_outputs(11947)) xor (layer2_outputs(9726));
    outputs(6734) <= layer2_outputs(7892);
    outputs(6735) <= not(layer2_outputs(1920)) or (layer2_outputs(5864));
    outputs(6736) <= layer2_outputs(3493);
    outputs(6737) <= (layer2_outputs(1793)) or (layer2_outputs(1281));
    outputs(6738) <= layer2_outputs(11206);
    outputs(6739) <= layer2_outputs(11592);
    outputs(6740) <= not(layer2_outputs(7093));
    outputs(6741) <= (layer2_outputs(12168)) and not (layer2_outputs(9565));
    outputs(6742) <= not(layer2_outputs(7533)) or (layer2_outputs(3230));
    outputs(6743) <= not((layer2_outputs(12791)) xor (layer2_outputs(5132)));
    outputs(6744) <= not(layer2_outputs(5471));
    outputs(6745) <= layer2_outputs(10420);
    outputs(6746) <= layer2_outputs(3073);
    outputs(6747) <= layer2_outputs(1502);
    outputs(6748) <= (layer2_outputs(3819)) xor (layer2_outputs(5866));
    outputs(6749) <= not(layer2_outputs(11517));
    outputs(6750) <= not(layer2_outputs(10280));
    outputs(6751) <= not((layer2_outputs(10774)) and (layer2_outputs(7907)));
    outputs(6752) <= not(layer2_outputs(6623));
    outputs(6753) <= layer2_outputs(3877);
    outputs(6754) <= not((layer2_outputs(7028)) xor (layer2_outputs(9826)));
    outputs(6755) <= layer2_outputs(2199);
    outputs(6756) <= not(layer2_outputs(3323));
    outputs(6757) <= layer2_outputs(3017);
    outputs(6758) <= layer2_outputs(6542);
    outputs(6759) <= not(layer2_outputs(333));
    outputs(6760) <= (layer2_outputs(2716)) xor (layer2_outputs(5331));
    outputs(6761) <= not(layer2_outputs(5950)) or (layer2_outputs(7216));
    outputs(6762) <= not((layer2_outputs(329)) xor (layer2_outputs(5673)));
    outputs(6763) <= layer2_outputs(8399);
    outputs(6764) <= (layer2_outputs(1502)) and not (layer2_outputs(3036));
    outputs(6765) <= not(layer2_outputs(8535));
    outputs(6766) <= (layer2_outputs(10082)) or (layer2_outputs(5982));
    outputs(6767) <= not(layer2_outputs(9530));
    outputs(6768) <= (layer2_outputs(1737)) xor (layer2_outputs(3696));
    outputs(6769) <= layer2_outputs(5771);
    outputs(6770) <= not((layer2_outputs(257)) xor (layer2_outputs(9909)));
    outputs(6771) <= (layer2_outputs(3420)) xor (layer2_outputs(2730));
    outputs(6772) <= not(layer2_outputs(9316));
    outputs(6773) <= not(layer2_outputs(917));
    outputs(6774) <= (layer2_outputs(6758)) xor (layer2_outputs(5378));
    outputs(6775) <= not(layer2_outputs(6695));
    outputs(6776) <= not(layer2_outputs(6574));
    outputs(6777) <= (layer2_outputs(9654)) and not (layer2_outputs(1104));
    outputs(6778) <= not(layer2_outputs(1947));
    outputs(6779) <= not((layer2_outputs(2672)) and (layer2_outputs(2017)));
    outputs(6780) <= layer2_outputs(10135);
    outputs(6781) <= (layer2_outputs(8919)) and not (layer2_outputs(11366));
    outputs(6782) <= not(layer2_outputs(5384)) or (layer2_outputs(3527));
    outputs(6783) <= layer2_outputs(9392);
    outputs(6784) <= (layer2_outputs(10334)) xor (layer2_outputs(819));
    outputs(6785) <= not(layer2_outputs(7542));
    outputs(6786) <= layer2_outputs(6401);
    outputs(6787) <= not(layer2_outputs(7952));
    outputs(6788) <= not(layer2_outputs(156));
    outputs(6789) <= not(layer2_outputs(1116));
    outputs(6790) <= (layer2_outputs(3883)) xor (layer2_outputs(11822));
    outputs(6791) <= not(layer2_outputs(6916));
    outputs(6792) <= (layer2_outputs(4330)) and not (layer2_outputs(10329));
    outputs(6793) <= (layer2_outputs(12171)) and (layer2_outputs(2879));
    outputs(6794) <= not((layer2_outputs(3956)) xor (layer2_outputs(1422)));
    outputs(6795) <= (layer2_outputs(8456)) xor (layer2_outputs(4030));
    outputs(6796) <= (layer2_outputs(8207)) and not (layer2_outputs(7289));
    outputs(6797) <= not(layer2_outputs(7213));
    outputs(6798) <= not(layer2_outputs(760));
    outputs(6799) <= layer2_outputs(4738);
    outputs(6800) <= layer2_outputs(10788);
    outputs(6801) <= (layer2_outputs(10591)) and (layer2_outputs(3389));
    outputs(6802) <= not(layer2_outputs(5016));
    outputs(6803) <= not(layer2_outputs(10242));
    outputs(6804) <= layer2_outputs(5722);
    outputs(6805) <= not(layer2_outputs(7021)) or (layer2_outputs(9735));
    outputs(6806) <= layer2_outputs(10483);
    outputs(6807) <= not(layer2_outputs(1825));
    outputs(6808) <= layer2_outputs(10810);
    outputs(6809) <= (layer2_outputs(4852)) xor (layer2_outputs(8745));
    outputs(6810) <= not((layer2_outputs(5848)) xor (layer2_outputs(3567)));
    outputs(6811) <= (layer2_outputs(1488)) xor (layer2_outputs(3500));
    outputs(6812) <= not(layer2_outputs(11842));
    outputs(6813) <= (layer2_outputs(2931)) and not (layer2_outputs(6707));
    outputs(6814) <= not(layer2_outputs(4981));
    outputs(6815) <= not(layer2_outputs(3096));
    outputs(6816) <= layer2_outputs(768);
    outputs(6817) <= not(layer2_outputs(10751));
    outputs(6818) <= not(layer2_outputs(10939)) or (layer2_outputs(2106));
    outputs(6819) <= not(layer2_outputs(7546));
    outputs(6820) <= layer2_outputs(11935);
    outputs(6821) <= not((layer2_outputs(6537)) and (layer2_outputs(5637)));
    outputs(6822) <= (layer2_outputs(11208)) xor (layer2_outputs(5895));
    outputs(6823) <= layer2_outputs(5164);
    outputs(6824) <= not(layer2_outputs(10724)) or (layer2_outputs(1208));
    outputs(6825) <= layer2_outputs(9351);
    outputs(6826) <= layer2_outputs(7015);
    outputs(6827) <= (layer2_outputs(2381)) xor (layer2_outputs(9306));
    outputs(6828) <= not(layer2_outputs(9460)) or (layer2_outputs(9153));
    outputs(6829) <= layer2_outputs(1751);
    outputs(6830) <= not((layer2_outputs(6804)) and (layer2_outputs(7979)));
    outputs(6831) <= not(layer2_outputs(1378));
    outputs(6832) <= (layer2_outputs(3193)) xor (layer2_outputs(6159));
    outputs(6833) <= not(layer2_outputs(3083));
    outputs(6834) <= layer2_outputs(10368);
    outputs(6835) <= not((layer2_outputs(1430)) xor (layer2_outputs(10563)));
    outputs(6836) <= layer2_outputs(1767);
    outputs(6837) <= not(layer2_outputs(9339)) or (layer2_outputs(4784));
    outputs(6838) <= not((layer2_outputs(11432)) xor (layer2_outputs(1839)));
    outputs(6839) <= not(layer2_outputs(12766));
    outputs(6840) <= layer2_outputs(10870);
    outputs(6841) <= not(layer2_outputs(2204));
    outputs(6842) <= layer2_outputs(7944);
    outputs(6843) <= (layer2_outputs(8994)) xor (layer2_outputs(7025));
    outputs(6844) <= (layer2_outputs(7594)) and not (layer2_outputs(9237));
    outputs(6845) <= not((layer2_outputs(789)) and (layer2_outputs(1205)));
    outputs(6846) <= (layer2_outputs(8253)) xor (layer2_outputs(1789));
    outputs(6847) <= (layer2_outputs(5638)) and not (layer2_outputs(1316));
    outputs(6848) <= not((layer2_outputs(11793)) xor (layer2_outputs(146)));
    outputs(6849) <= not((layer2_outputs(1773)) xor (layer2_outputs(9159)));
    outputs(6850) <= not((layer2_outputs(3101)) and (layer2_outputs(6045)));
    outputs(6851) <= not((layer2_outputs(9877)) or (layer2_outputs(1339)));
    outputs(6852) <= (layer2_outputs(3892)) or (layer2_outputs(6969));
    outputs(6853) <= not(layer2_outputs(10897));
    outputs(6854) <= layer2_outputs(4428);
    outputs(6855) <= not(layer2_outputs(2441));
    outputs(6856) <= layer2_outputs(1017);
    outputs(6857) <= not(layer2_outputs(1980));
    outputs(6858) <= not((layer2_outputs(7929)) xor (layer2_outputs(127)));
    outputs(6859) <= layer2_outputs(10057);
    outputs(6860) <= not((layer2_outputs(5091)) or (layer2_outputs(12068)));
    outputs(6861) <= layer2_outputs(2162);
    outputs(6862) <= not((layer2_outputs(1571)) xor (layer2_outputs(9412)));
    outputs(6863) <= not(layer2_outputs(2514));
    outputs(6864) <= not(layer2_outputs(8609));
    outputs(6865) <= (layer2_outputs(7338)) xor (layer2_outputs(3640));
    outputs(6866) <= not(layer2_outputs(2046));
    outputs(6867) <= (layer2_outputs(2105)) and not (layer2_outputs(1482));
    outputs(6868) <= layer2_outputs(12372);
    outputs(6869) <= not(layer2_outputs(5418));
    outputs(6870) <= not((layer2_outputs(10338)) xor (layer2_outputs(839)));
    outputs(6871) <= not((layer2_outputs(5361)) xor (layer2_outputs(4390)));
    outputs(6872) <= (layer2_outputs(2318)) xor (layer2_outputs(8720));
    outputs(6873) <= not(layer2_outputs(8979));
    outputs(6874) <= (layer2_outputs(8875)) or (layer2_outputs(12511));
    outputs(6875) <= (layer2_outputs(4895)) xor (layer2_outputs(11059));
    outputs(6876) <= not((layer2_outputs(10501)) xor (layer2_outputs(6034)));
    outputs(6877) <= not(layer2_outputs(3541));
    outputs(6878) <= not((layer2_outputs(12684)) xor (layer2_outputs(9144)));
    outputs(6879) <= not(layer2_outputs(10013));
    outputs(6880) <= (layer2_outputs(11871)) xor (layer2_outputs(6872));
    outputs(6881) <= layer2_outputs(6556);
    outputs(6882) <= not(layer2_outputs(10514));
    outputs(6883) <= (layer2_outputs(1698)) xor (layer2_outputs(8224));
    outputs(6884) <= (layer2_outputs(7792)) and not (layer2_outputs(7719));
    outputs(6885) <= not(layer2_outputs(4543));
    outputs(6886) <= not(layer2_outputs(6799));
    outputs(6887) <= (layer2_outputs(11103)) or (layer2_outputs(6175));
    outputs(6888) <= (layer2_outputs(6762)) and (layer2_outputs(1532));
    outputs(6889) <= layer2_outputs(4600);
    outputs(6890) <= not((layer2_outputs(9082)) xor (layer2_outputs(4581)));
    outputs(6891) <= not(layer2_outputs(4973));
    outputs(6892) <= not((layer2_outputs(8137)) xor (layer2_outputs(8685)));
    outputs(6893) <= not((layer2_outputs(5709)) and (layer2_outputs(1157)));
    outputs(6894) <= not(layer2_outputs(3562));
    outputs(6895) <= layer2_outputs(3275);
    outputs(6896) <= not(layer2_outputs(3992));
    outputs(6897) <= not((layer2_outputs(1359)) xor (layer2_outputs(4963)));
    outputs(6898) <= layer2_outputs(2228);
    outputs(6899) <= not((layer2_outputs(11820)) xor (layer2_outputs(6568)));
    outputs(6900) <= not(layer2_outputs(10581));
    outputs(6901) <= not(layer2_outputs(8188));
    outputs(6902) <= layer2_outputs(9679);
    outputs(6903) <= (layer2_outputs(4126)) xor (layer2_outputs(12017));
    outputs(6904) <= layer2_outputs(1279);
    outputs(6905) <= (layer2_outputs(5074)) xor (layer2_outputs(5170));
    outputs(6906) <= layer2_outputs(10646);
    outputs(6907) <= not((layer2_outputs(715)) xor (layer2_outputs(1544)));
    outputs(6908) <= layer2_outputs(8129);
    outputs(6909) <= layer2_outputs(10786);
    outputs(6910) <= layer2_outputs(2165);
    outputs(6911) <= not(layer2_outputs(9620));
    outputs(6912) <= layer2_outputs(9355);
    outputs(6913) <= layer2_outputs(5684);
    outputs(6914) <= not(layer2_outputs(10487));
    outputs(6915) <= (layer2_outputs(8141)) and not (layer2_outputs(5755));
    outputs(6916) <= layer2_outputs(6836);
    outputs(6917) <= (layer2_outputs(1689)) xor (layer2_outputs(9680));
    outputs(6918) <= (layer2_outputs(7412)) xor (layer2_outputs(10813));
    outputs(6919) <= not((layer2_outputs(6267)) xor (layer2_outputs(11002)));
    outputs(6920) <= not((layer2_outputs(7731)) or (layer2_outputs(522)));
    outputs(6921) <= not(layer2_outputs(1639));
    outputs(6922) <= not(layer2_outputs(6482));
    outputs(6923) <= not(layer2_outputs(4943));
    outputs(6924) <= (layer2_outputs(3863)) xor (layer2_outputs(8490));
    outputs(6925) <= (layer2_outputs(8112)) and not (layer2_outputs(6450));
    outputs(6926) <= not((layer2_outputs(827)) and (layer2_outputs(8628)));
    outputs(6927) <= not(layer2_outputs(5050));
    outputs(6928) <= not(layer2_outputs(641));
    outputs(6929) <= not((layer2_outputs(1962)) xor (layer2_outputs(5151)));
    outputs(6930) <= (layer2_outputs(10730)) xor (layer2_outputs(9577));
    outputs(6931) <= (layer2_outputs(2535)) xor (layer2_outputs(1477));
    outputs(6932) <= layer2_outputs(958);
    outputs(6933) <= not(layer2_outputs(1268));
    outputs(6934) <= layer2_outputs(3069);
    outputs(6935) <= (layer2_outputs(12144)) and not (layer2_outputs(7366));
    outputs(6936) <= not(layer2_outputs(12776));
    outputs(6937) <= (layer2_outputs(570)) xor (layer2_outputs(7660));
    outputs(6938) <= layer2_outputs(5985);
    outputs(6939) <= layer2_outputs(9527);
    outputs(6940) <= (layer2_outputs(1693)) xor (layer2_outputs(7102));
    outputs(6941) <= (layer2_outputs(61)) xor (layer2_outputs(2375));
    outputs(6942) <= layer2_outputs(8985);
    outputs(6943) <= layer2_outputs(2344);
    outputs(6944) <= (layer2_outputs(1249)) or (layer2_outputs(11838));
    outputs(6945) <= (layer2_outputs(695)) xor (layer2_outputs(699));
    outputs(6946) <= layer2_outputs(6046);
    outputs(6947) <= layer2_outputs(2560);
    outputs(6948) <= layer2_outputs(5305);
    outputs(6949) <= layer2_outputs(5783);
    outputs(6950) <= not((layer2_outputs(4651)) xor (layer2_outputs(7504)));
    outputs(6951) <= (layer2_outputs(6021)) or (layer2_outputs(6919));
    outputs(6952) <= layer2_outputs(12545);
    outputs(6953) <= not(layer2_outputs(2061)) or (layer2_outputs(6664));
    outputs(6954) <= not(layer2_outputs(5181));
    outputs(6955) <= layer2_outputs(6223);
    outputs(6956) <= (layer2_outputs(3376)) xor (layer2_outputs(1981));
    outputs(6957) <= (layer2_outputs(9165)) and not (layer2_outputs(11525));
    outputs(6958) <= not(layer2_outputs(6312));
    outputs(6959) <= layer2_outputs(2315);
    outputs(6960) <= layer2_outputs(5476);
    outputs(6961) <= not(layer2_outputs(2213));
    outputs(6962) <= not(layer2_outputs(2235));
    outputs(6963) <= layer2_outputs(11943);
    outputs(6964) <= not((layer2_outputs(1119)) xor (layer2_outputs(3045)));
    outputs(6965) <= not(layer2_outputs(3490));
    outputs(6966) <= (layer2_outputs(435)) xor (layer2_outputs(1600));
    outputs(6967) <= layer2_outputs(8754);
    outputs(6968) <= not(layer2_outputs(7650));
    outputs(6969) <= layer2_outputs(4826);
    outputs(6970) <= not(layer2_outputs(5295));
    outputs(6971) <= layer2_outputs(11428);
    outputs(6972) <= not(layer2_outputs(11848));
    outputs(6973) <= not((layer2_outputs(1055)) xor (layer2_outputs(9028)));
    outputs(6974) <= layer2_outputs(6468);
    outputs(6975) <= (layer2_outputs(7717)) xor (layer2_outputs(1016));
    outputs(6976) <= layer2_outputs(8413);
    outputs(6977) <= not(layer2_outputs(3295));
    outputs(6978) <= not(layer2_outputs(10479));
    outputs(6979) <= not((layer2_outputs(2129)) and (layer2_outputs(7086)));
    outputs(6980) <= not((layer2_outputs(4033)) or (layer2_outputs(12126)));
    outputs(6981) <= (layer2_outputs(2798)) xor (layer2_outputs(1917));
    outputs(6982) <= not((layer2_outputs(3001)) or (layer2_outputs(9369)));
    outputs(6983) <= not(layer2_outputs(1569));
    outputs(6984) <= not(layer2_outputs(6278));
    outputs(6985) <= not((layer2_outputs(4907)) xor (layer2_outputs(8705)));
    outputs(6986) <= not((layer2_outputs(5038)) and (layer2_outputs(11211)));
    outputs(6987) <= not((layer2_outputs(5067)) xor (layer2_outputs(4511)));
    outputs(6988) <= layer2_outputs(863);
    outputs(6989) <= not((layer2_outputs(11765)) xor (layer2_outputs(3474)));
    outputs(6990) <= (layer2_outputs(7670)) and not (layer2_outputs(979));
    outputs(6991) <= not((layer2_outputs(7166)) xor (layer2_outputs(6863)));
    outputs(6992) <= layer2_outputs(2164);
    outputs(6993) <= layer2_outputs(3564);
    outputs(6994) <= (layer2_outputs(8180)) xor (layer2_outputs(7812));
    outputs(6995) <= layer2_outputs(2908);
    outputs(6996) <= layer2_outputs(5404);
    outputs(6997) <= layer2_outputs(199);
    outputs(6998) <= not(layer2_outputs(11041));
    outputs(6999) <= not(layer2_outputs(11869)) or (layer2_outputs(4300));
    outputs(7000) <= not(layer2_outputs(3893));
    outputs(7001) <= not(layer2_outputs(2546));
    outputs(7002) <= not(layer2_outputs(6070));
    outputs(7003) <= not((layer2_outputs(8311)) xor (layer2_outputs(10211)));
    outputs(7004) <= not(layer2_outputs(12056));
    outputs(7005) <= (layer2_outputs(8187)) xor (layer2_outputs(626));
    outputs(7006) <= not((layer2_outputs(10594)) xor (layer2_outputs(11151)));
    outputs(7007) <= not((layer2_outputs(11986)) xor (layer2_outputs(2106)));
    outputs(7008) <= not((layer2_outputs(3466)) and (layer2_outputs(10392)));
    outputs(7009) <= (layer2_outputs(5300)) and (layer2_outputs(6861));
    outputs(7010) <= (layer2_outputs(2735)) or (layer2_outputs(8643));
    outputs(7011) <= layer2_outputs(6857);
    outputs(7012) <= layer2_outputs(7278);
    outputs(7013) <= (layer2_outputs(7633)) xor (layer2_outputs(11436));
    outputs(7014) <= not((layer2_outputs(5737)) xor (layer2_outputs(7486)));
    outputs(7015) <= layer2_outputs(5262);
    outputs(7016) <= layer2_outputs(7482);
    outputs(7017) <= (layer2_outputs(236)) and not (layer2_outputs(11532));
    outputs(7018) <= not(layer2_outputs(11081));
    outputs(7019) <= layer2_outputs(2702);
    outputs(7020) <= (layer2_outputs(3682)) xor (layer2_outputs(1712));
    outputs(7021) <= not(layer2_outputs(1284)) or (layer2_outputs(3337));
    outputs(7022) <= (layer2_outputs(588)) xor (layer2_outputs(8799));
    outputs(7023) <= not((layer2_outputs(11075)) or (layer2_outputs(1253)));
    outputs(7024) <= not(layer2_outputs(3773)) or (layer2_outputs(11036));
    outputs(7025) <= layer2_outputs(6331);
    outputs(7026) <= layer2_outputs(6325);
    outputs(7027) <= (layer2_outputs(1769)) or (layer2_outputs(955));
    outputs(7028) <= not(layer2_outputs(10136));
    outputs(7029) <= layer2_outputs(5463);
    outputs(7030) <= layer2_outputs(12591);
    outputs(7031) <= layer2_outputs(10991);
    outputs(7032) <= layer2_outputs(12678);
    outputs(7033) <= (layer2_outputs(3342)) xor (layer2_outputs(10404));
    outputs(7034) <= layer2_outputs(2115);
    outputs(7035) <= (layer2_outputs(11677)) and not (layer2_outputs(763));
    outputs(7036) <= not(layer2_outputs(12000));
    outputs(7037) <= layer2_outputs(9177);
    outputs(7038) <= not((layer2_outputs(11034)) xor (layer2_outputs(1482)));
    outputs(7039) <= not(layer2_outputs(3833));
    outputs(7040) <= layer2_outputs(5102);
    outputs(7041) <= not(layer2_outputs(9531));
    outputs(7042) <= not(layer2_outputs(3850));
    outputs(7043) <= (layer2_outputs(7805)) and not (layer2_outputs(8690));
    outputs(7044) <= layer2_outputs(1383);
    outputs(7045) <= not(layer2_outputs(7133)) or (layer2_outputs(9860));
    outputs(7046) <= not((layer2_outputs(6029)) xor (layer2_outputs(10782)));
    outputs(7047) <= (layer2_outputs(12346)) xor (layer2_outputs(1379));
    outputs(7048) <= layer2_outputs(2612);
    outputs(7049) <= layer2_outputs(10792);
    outputs(7050) <= not(layer2_outputs(8863));
    outputs(7051) <= not((layer2_outputs(10593)) or (layer2_outputs(11512)));
    outputs(7052) <= not((layer2_outputs(5878)) or (layer2_outputs(11436)));
    outputs(7053) <= (layer2_outputs(1959)) or (layer2_outputs(4963));
    outputs(7054) <= not(layer2_outputs(12542));
    outputs(7055) <= not(layer2_outputs(5899));
    outputs(7056) <= layer2_outputs(12396);
    outputs(7057) <= not(layer2_outputs(2107));
    outputs(7058) <= layer2_outputs(9366);
    outputs(7059) <= layer2_outputs(4558);
    outputs(7060) <= layer2_outputs(2237);
    outputs(7061) <= (layer2_outputs(5053)) and not (layer2_outputs(10927));
    outputs(7062) <= not((layer2_outputs(5617)) xor (layer2_outputs(1403)));
    outputs(7063) <= layer2_outputs(11430);
    outputs(7064) <= not(layer2_outputs(1114));
    outputs(7065) <= (layer2_outputs(5258)) and (layer2_outputs(12322));
    outputs(7066) <= not((layer2_outputs(9159)) xor (layer2_outputs(12588)));
    outputs(7067) <= layer2_outputs(10996);
    outputs(7068) <= not((layer2_outputs(11815)) xor (layer2_outputs(6793)));
    outputs(7069) <= not(layer2_outputs(10921));
    outputs(7070) <= (layer2_outputs(3525)) and not (layer2_outputs(11655));
    outputs(7071) <= not(layer2_outputs(12040));
    outputs(7072) <= (layer2_outputs(11708)) or (layer2_outputs(5953));
    outputs(7073) <= (layer2_outputs(5085)) xor (layer2_outputs(6739));
    outputs(7074) <= (layer2_outputs(3527)) xor (layer2_outputs(5759));
    outputs(7075) <= not(layer2_outputs(2522));
    outputs(7076) <= (layer2_outputs(3282)) xor (layer2_outputs(9562));
    outputs(7077) <= not(layer2_outputs(4145));
    outputs(7078) <= layer2_outputs(9891);
    outputs(7079) <= layer2_outputs(8689);
    outputs(7080) <= not(layer2_outputs(8264)) or (layer2_outputs(9446));
    outputs(7081) <= not(layer2_outputs(9401));
    outputs(7082) <= (layer2_outputs(5264)) and (layer2_outputs(2843));
    outputs(7083) <= layer2_outputs(4101);
    outputs(7084) <= not((layer2_outputs(9802)) xor (layer2_outputs(2245)));
    outputs(7085) <= (layer2_outputs(5728)) xor (layer2_outputs(931));
    outputs(7086) <= not((layer2_outputs(5232)) or (layer2_outputs(11297)));
    outputs(7087) <= not(layer2_outputs(10316));
    outputs(7088) <= (layer2_outputs(210)) and not (layer2_outputs(2226));
    outputs(7089) <= (layer2_outputs(11433)) xor (layer2_outputs(10608));
    outputs(7090) <= not(layer2_outputs(2650));
    outputs(7091) <= (layer2_outputs(8432)) or (layer2_outputs(8647));
    outputs(7092) <= not(layer2_outputs(270));
    outputs(7093) <= not((layer2_outputs(11183)) xor (layer2_outputs(1652)));
    outputs(7094) <= layer2_outputs(3298);
    outputs(7095) <= layer2_outputs(10857);
    outputs(7096) <= not((layer2_outputs(2282)) xor (layer2_outputs(4248)));
    outputs(7097) <= not(layer2_outputs(38));
    outputs(7098) <= not((layer2_outputs(12608)) xor (layer2_outputs(5902)));
    outputs(7099) <= not(layer2_outputs(8731));
    outputs(7100) <= not((layer2_outputs(203)) xor (layer2_outputs(10361)));
    outputs(7101) <= not(layer2_outputs(5160));
    outputs(7102) <= (layer2_outputs(3261)) xor (layer2_outputs(12525));
    outputs(7103) <= (layer2_outputs(12537)) xor (layer2_outputs(7606));
    outputs(7104) <= not((layer2_outputs(1274)) xor (layer2_outputs(2706)));
    outputs(7105) <= not(layer2_outputs(3383));
    outputs(7106) <= not(layer2_outputs(4238));
    outputs(7107) <= not(layer2_outputs(3491));
    outputs(7108) <= layer2_outputs(1976);
    outputs(7109) <= layer2_outputs(7483);
    outputs(7110) <= (layer2_outputs(751)) xor (layer2_outputs(4788));
    outputs(7111) <= (layer2_outputs(8493)) and (layer2_outputs(10420));
    outputs(7112) <= layer2_outputs(10319);
    outputs(7113) <= (layer2_outputs(10911)) xor (layer2_outputs(1704));
    outputs(7114) <= not((layer2_outputs(3507)) and (layer2_outputs(10908)));
    outputs(7115) <= not((layer2_outputs(7208)) xor (layer2_outputs(5011)));
    outputs(7116) <= not((layer2_outputs(4400)) xor (layer2_outputs(3285)));
    outputs(7117) <= not((layer2_outputs(4628)) xor (layer2_outputs(10943)));
    outputs(7118) <= (layer2_outputs(1559)) xor (layer2_outputs(7574));
    outputs(7119) <= (layer2_outputs(3029)) xor (layer2_outputs(11362));
    outputs(7120) <= not(layer2_outputs(2669));
    outputs(7121) <= layer2_outputs(12799);
    outputs(7122) <= layer2_outputs(12450);
    outputs(7123) <= not((layer2_outputs(6309)) xor (layer2_outputs(5480)));
    outputs(7124) <= (layer2_outputs(7780)) or (layer2_outputs(523));
    outputs(7125) <= not(layer2_outputs(7981));
    outputs(7126) <= not((layer2_outputs(12469)) xor (layer2_outputs(10868)));
    outputs(7127) <= not(layer2_outputs(6273));
    outputs(7128) <= layer2_outputs(1112);
    outputs(7129) <= layer2_outputs(10798);
    outputs(7130) <= layer2_outputs(4047);
    outputs(7131) <= not(layer2_outputs(2917));
    outputs(7132) <= not((layer2_outputs(4066)) xor (layer2_outputs(2554)));
    outputs(7133) <= layer2_outputs(4864);
    outputs(7134) <= (layer2_outputs(11570)) or (layer2_outputs(6334));
    outputs(7135) <= not(layer2_outputs(5939));
    outputs(7136) <= not(layer2_outputs(10643));
    outputs(7137) <= not(layer2_outputs(10174));
    outputs(7138) <= (layer2_outputs(9720)) and not (layer2_outputs(12626));
    outputs(7139) <= not(layer2_outputs(10126));
    outputs(7140) <= layer2_outputs(117);
    outputs(7141) <= not((layer2_outputs(9906)) xor (layer2_outputs(9629)));
    outputs(7142) <= not(layer2_outputs(534));
    outputs(7143) <= not((layer2_outputs(3596)) xor (layer2_outputs(2795)));
    outputs(7144) <= (layer2_outputs(8795)) and not (layer2_outputs(12795));
    outputs(7145) <= (layer2_outputs(2869)) xor (layer2_outputs(879));
    outputs(7146) <= layer2_outputs(3529);
    outputs(7147) <= not(layer2_outputs(9261));
    outputs(7148) <= (layer2_outputs(1201)) or (layer2_outputs(1320));
    outputs(7149) <= layer2_outputs(7073);
    outputs(7150) <= (layer2_outputs(595)) and (layer2_outputs(3103));
    outputs(7151) <= (layer2_outputs(12285)) and (layer2_outputs(12560));
    outputs(7152) <= not((layer2_outputs(1972)) xor (layer2_outputs(879)));
    outputs(7153) <= layer2_outputs(994);
    outputs(7154) <= (layer2_outputs(4012)) and (layer2_outputs(1925));
    outputs(7155) <= not(layer2_outputs(6115)) or (layer2_outputs(11144));
    outputs(7156) <= layer2_outputs(2557);
    outputs(7157) <= not(layer2_outputs(9647));
    outputs(7158) <= layer2_outputs(773);
    outputs(7159) <= not(layer2_outputs(11318));
    outputs(7160) <= not((layer2_outputs(3194)) xor (layer2_outputs(6504)));
    outputs(7161) <= layer2_outputs(9429);
    outputs(7162) <= not((layer2_outputs(1265)) xor (layer2_outputs(5624)));
    outputs(7163) <= layer2_outputs(6021);
    outputs(7164) <= layer2_outputs(1007);
    outputs(7165) <= (layer2_outputs(10495)) xor (layer2_outputs(5419));
    outputs(7166) <= layer2_outputs(10028);
    outputs(7167) <= layer2_outputs(1414);
    outputs(7168) <= (layer2_outputs(4184)) xor (layer2_outputs(3943));
    outputs(7169) <= not((layer2_outputs(3394)) xor (layer2_outputs(5574)));
    outputs(7170) <= not(layer2_outputs(681));
    outputs(7171) <= layer2_outputs(12617);
    outputs(7172) <= not((layer2_outputs(12744)) xor (layer2_outputs(3278)));
    outputs(7173) <= not((layer2_outputs(12262)) and (layer2_outputs(1379)));
    outputs(7174) <= (layer2_outputs(2486)) or (layer2_outputs(12466));
    outputs(7175) <= not((layer2_outputs(6632)) xor (layer2_outputs(10678)));
    outputs(7176) <= not(layer2_outputs(3437)) or (layer2_outputs(10796));
    outputs(7177) <= (layer2_outputs(8976)) xor (layer2_outputs(12222));
    outputs(7178) <= not(layer2_outputs(6810));
    outputs(7179) <= layer2_outputs(5656);
    outputs(7180) <= not(layer2_outputs(39));
    outputs(7181) <= not((layer2_outputs(11264)) xor (layer2_outputs(9595)));
    outputs(7182) <= layer2_outputs(2915);
    outputs(7183) <= not(layer2_outputs(11594));
    outputs(7184) <= not(layer2_outputs(1961));
    outputs(7185) <= not(layer2_outputs(136));
    outputs(7186) <= not((layer2_outputs(7413)) xor (layer2_outputs(1266)));
    outputs(7187) <= (layer2_outputs(7200)) xor (layer2_outputs(2773));
    outputs(7188) <= (layer2_outputs(5669)) xor (layer2_outputs(6689));
    outputs(7189) <= layer2_outputs(7541);
    outputs(7190) <= layer2_outputs(6352);
    outputs(7191) <= (layer2_outputs(8143)) xor (layer2_outputs(12250));
    outputs(7192) <= not(layer2_outputs(5350));
    outputs(7193) <= (layer2_outputs(5115)) xor (layer2_outputs(12739));
    outputs(7194) <= not(layer2_outputs(3516));
    outputs(7195) <= (layer2_outputs(1272)) xor (layer2_outputs(7567));
    outputs(7196) <= not((layer2_outputs(11560)) xor (layer2_outputs(5457)));
    outputs(7197) <= not((layer2_outputs(12275)) xor (layer2_outputs(5585)));
    outputs(7198) <= layer2_outputs(11248);
    outputs(7199) <= layer2_outputs(6286);
    outputs(7200) <= layer2_outputs(2317);
    outputs(7201) <= not((layer2_outputs(57)) xor (layer2_outputs(2594)));
    outputs(7202) <= (layer2_outputs(8091)) or (layer2_outputs(8082));
    outputs(7203) <= layer2_outputs(9903);
    outputs(7204) <= not((layer2_outputs(9227)) or (layer2_outputs(11255)));
    outputs(7205) <= not(layer2_outputs(1344));
    outputs(7206) <= (layer2_outputs(2965)) xor (layer2_outputs(5544));
    outputs(7207) <= not((layer2_outputs(11880)) or (layer2_outputs(8617)));
    outputs(7208) <= not((layer2_outputs(1078)) xor (layer2_outputs(10199)));
    outputs(7209) <= not(layer2_outputs(6928));
    outputs(7210) <= (layer2_outputs(11067)) or (layer2_outputs(3929));
    outputs(7211) <= layer2_outputs(171);
    outputs(7212) <= not(layer2_outputs(12243));
    outputs(7213) <= (layer2_outputs(5706)) and not (layer2_outputs(182));
    outputs(7214) <= layer2_outputs(10114);
    outputs(7215) <= not(layer2_outputs(4478));
    outputs(7216) <= not(layer2_outputs(1923));
    outputs(7217) <= not(layer2_outputs(2777));
    outputs(7218) <= not(layer2_outputs(10294));
    outputs(7219) <= not(layer2_outputs(5619)) or (layer2_outputs(12685));
    outputs(7220) <= not(layer2_outputs(9038));
    outputs(7221) <= (layer2_outputs(11685)) xor (layer2_outputs(4204));
    outputs(7222) <= layer2_outputs(6675);
    outputs(7223) <= not((layer2_outputs(2185)) xor (layer2_outputs(8934)));
    outputs(7224) <= not(layer2_outputs(4781));
    outputs(7225) <= not(layer2_outputs(8389));
    outputs(7226) <= (layer2_outputs(1360)) xor (layer2_outputs(6838));
    outputs(7227) <= layer2_outputs(8724);
    outputs(7228) <= not((layer2_outputs(9512)) and (layer2_outputs(1140)));
    outputs(7229) <= (layer2_outputs(1727)) xor (layer2_outputs(9179));
    outputs(7230) <= (layer2_outputs(2994)) xor (layer2_outputs(4676));
    outputs(7231) <= layer2_outputs(12072);
    outputs(7232) <= (layer2_outputs(5714)) xor (layer2_outputs(1443));
    outputs(7233) <= (layer2_outputs(2542)) xor (layer2_outputs(11201));
    outputs(7234) <= layer2_outputs(4817);
    outputs(7235) <= (layer2_outputs(1629)) and (layer2_outputs(2378));
    outputs(7236) <= layer2_outputs(6412);
    outputs(7237) <= (layer2_outputs(7869)) and not (layer2_outputs(2101));
    outputs(7238) <= (layer2_outputs(4840)) xor (layer2_outputs(2485));
    outputs(7239) <= not((layer2_outputs(5321)) xor (layer2_outputs(4210)));
    outputs(7240) <= not(layer2_outputs(4683));
    outputs(7241) <= layer2_outputs(4905);
    outputs(7242) <= (layer2_outputs(856)) xor (layer2_outputs(3684));
    outputs(7243) <= layer2_outputs(7007);
    outputs(7244) <= not(layer2_outputs(6417));
    outputs(7245) <= not(layer2_outputs(9792));
    outputs(7246) <= layer2_outputs(9809);
    outputs(7247) <= (layer2_outputs(1717)) or (layer2_outputs(10660));
    outputs(7248) <= (layer2_outputs(506)) xor (layer2_outputs(3063));
    outputs(7249) <= not(layer2_outputs(1784));
    outputs(7250) <= not(layer2_outputs(2207));
    outputs(7251) <= (layer2_outputs(29)) xor (layer2_outputs(12160));
    outputs(7252) <= (layer2_outputs(1761)) xor (layer2_outputs(8961));
    outputs(7253) <= not(layer2_outputs(2978));
    outputs(7254) <= (layer2_outputs(9886)) xor (layer2_outputs(7593));
    outputs(7255) <= layer2_outputs(8216);
    outputs(7256) <= layer2_outputs(9538);
    outputs(7257) <= not(layer2_outputs(4531));
    outputs(7258) <= not(layer2_outputs(7275));
    outputs(7259) <= (layer2_outputs(8732)) and (layer2_outputs(10386));
    outputs(7260) <= layer2_outputs(6990);
    outputs(7261) <= (layer2_outputs(6106)) and (layer2_outputs(4965));
    outputs(7262) <= layer2_outputs(3973);
    outputs(7263) <= layer2_outputs(7937);
    outputs(7264) <= (layer2_outputs(1667)) xor (layer2_outputs(4305));
    outputs(7265) <= layer2_outputs(12228);
    outputs(7266) <= not((layer2_outputs(5561)) and (layer2_outputs(5613)));
    outputs(7267) <= not(layer2_outputs(7542));
    outputs(7268) <= (layer2_outputs(6116)) and not (layer2_outputs(6620));
    outputs(7269) <= (layer2_outputs(11984)) xor (layer2_outputs(7567));
    outputs(7270) <= layer2_outputs(11227);
    outputs(7271) <= (layer2_outputs(2263)) or (layer2_outputs(3346));
    outputs(7272) <= not(layer2_outputs(6916));
    outputs(7273) <= (layer2_outputs(10268)) xor (layer2_outputs(8284));
    outputs(7274) <= not(layer2_outputs(10228));
    outputs(7275) <= (layer2_outputs(5742)) xor (layer2_outputs(7999));
    outputs(7276) <= not(layer2_outputs(12331));
    outputs(7277) <= layer2_outputs(630);
    outputs(7278) <= not(layer2_outputs(485)) or (layer2_outputs(850));
    outputs(7279) <= layer2_outputs(3652);
    outputs(7280) <= not((layer2_outputs(4311)) xor (layer2_outputs(749)));
    outputs(7281) <= not((layer2_outputs(5707)) xor (layer2_outputs(11283)));
    outputs(7282) <= not((layer2_outputs(9276)) or (layer2_outputs(5329)));
    outputs(7283) <= not((layer2_outputs(2132)) or (layer2_outputs(678)));
    outputs(7284) <= not(layer2_outputs(11640));
    outputs(7285) <= not(layer2_outputs(2647));
    outputs(7286) <= not(layer2_outputs(1097));
    outputs(7287) <= layer2_outputs(9561);
    outputs(7288) <= (layer2_outputs(2733)) xor (layer2_outputs(8263));
    outputs(7289) <= not(layer2_outputs(11743));
    outputs(7290) <= not(layer2_outputs(1023));
    outputs(7291) <= not((layer2_outputs(12191)) xor (layer2_outputs(8331)));
    outputs(7292) <= (layer2_outputs(11982)) xor (layer2_outputs(9407));
    outputs(7293) <= layer2_outputs(7222);
    outputs(7294) <= not((layer2_outputs(792)) xor (layer2_outputs(12516)));
    outputs(7295) <= layer2_outputs(12732);
    outputs(7296) <= layer2_outputs(12358);
    outputs(7297) <= not((layer2_outputs(4693)) xor (layer2_outputs(8961)));
    outputs(7298) <= (layer2_outputs(539)) xor (layer2_outputs(6251));
    outputs(7299) <= (layer2_outputs(3296)) xor (layer2_outputs(8125));
    outputs(7300) <= not(layer2_outputs(7082));
    outputs(7301) <= (layer2_outputs(4647)) and not (layer2_outputs(4820));
    outputs(7302) <= layer2_outputs(1240);
    outputs(7303) <= not((layer2_outputs(9189)) xor (layer2_outputs(299)));
    outputs(7304) <= (layer2_outputs(5781)) xor (layer2_outputs(5115));
    outputs(7305) <= not(layer2_outputs(8533));
    outputs(7306) <= not((layer2_outputs(4018)) and (layer2_outputs(12627)));
    outputs(7307) <= layer2_outputs(7392);
    outputs(7308) <= not((layer2_outputs(10144)) xor (layer2_outputs(11484)));
    outputs(7309) <= layer2_outputs(3863);
    outputs(7310) <= (layer2_outputs(9182)) xor (layer2_outputs(1576));
    outputs(7311) <= not((layer2_outputs(8637)) xor (layer2_outputs(12496)));
    outputs(7312) <= (layer2_outputs(10526)) xor (layer2_outputs(3621));
    outputs(7313) <= (layer2_outputs(5314)) xor (layer2_outputs(5185));
    outputs(7314) <= (layer2_outputs(6006)) or (layer2_outputs(530));
    outputs(7315) <= not((layer2_outputs(6317)) and (layer2_outputs(2033)));
    outputs(7316) <= (layer2_outputs(11920)) or (layer2_outputs(9713));
    outputs(7317) <= layer2_outputs(9077);
    outputs(7318) <= not(layer2_outputs(8336));
    outputs(7319) <= layer2_outputs(187);
    outputs(7320) <= (layer2_outputs(12435)) xor (layer2_outputs(12385));
    outputs(7321) <= (layer2_outputs(2680)) and not (layer2_outputs(4525));
    outputs(7322) <= (layer2_outputs(2259)) xor (layer2_outputs(5202));
    outputs(7323) <= (layer2_outputs(10247)) and not (layer2_outputs(11480));
    outputs(7324) <= (layer2_outputs(3868)) xor (layer2_outputs(3032));
    outputs(7325) <= not(layer2_outputs(5055));
    outputs(7326) <= layer2_outputs(11866);
    outputs(7327) <= layer2_outputs(4131);
    outputs(7328) <= layer2_outputs(8040);
    outputs(7329) <= layer2_outputs(7067);
    outputs(7330) <= (layer2_outputs(2437)) xor (layer2_outputs(2648));
    outputs(7331) <= (layer2_outputs(614)) and not (layer2_outputs(5856));
    outputs(7332) <= not(layer2_outputs(4839));
    outputs(7333) <= layer2_outputs(9737);
    outputs(7334) <= not((layer2_outputs(12148)) xor (layer2_outputs(3073)));
    outputs(7335) <= (layer2_outputs(4015)) xor (layer2_outputs(11488));
    outputs(7336) <= layer2_outputs(12403);
    outputs(7337) <= not((layer2_outputs(1409)) and (layer2_outputs(4496)));
    outputs(7338) <= layer2_outputs(5313);
    outputs(7339) <= layer2_outputs(7016);
    outputs(7340) <= (layer2_outputs(3120)) xor (layer2_outputs(7881));
    outputs(7341) <= not(layer2_outputs(4363));
    outputs(7342) <= not(layer2_outputs(5971));
    outputs(7343) <= not((layer2_outputs(5663)) xor (layer2_outputs(566)));
    outputs(7344) <= layer2_outputs(7471);
    outputs(7345) <= not(layer2_outputs(11870));
    outputs(7346) <= layer2_outputs(5099);
    outputs(7347) <= (layer2_outputs(9896)) xor (layer2_outputs(4972));
    outputs(7348) <= not(layer2_outputs(11081));
    outputs(7349) <= not(layer2_outputs(10173));
    outputs(7350) <= not(layer2_outputs(12710));
    outputs(7351) <= not(layer2_outputs(7631));
    outputs(7352) <= not(layer2_outputs(6367));
    outputs(7353) <= not((layer2_outputs(5144)) xor (layer2_outputs(5047)));
    outputs(7354) <= not(layer2_outputs(4555));
    outputs(7355) <= not((layer2_outputs(1601)) xor (layer2_outputs(6442)));
    outputs(7356) <= layer2_outputs(5510);
    outputs(7357) <= not((layer2_outputs(12533)) xor (layer2_outputs(5142)));
    outputs(7358) <= not(layer2_outputs(11292));
    outputs(7359) <= layer2_outputs(2993);
    outputs(7360) <= not(layer2_outputs(3442));
    outputs(7361) <= layer2_outputs(11478);
    outputs(7362) <= not((layer2_outputs(10455)) xor (layer2_outputs(3358)));
    outputs(7363) <= not((layer2_outputs(11146)) and (layer2_outputs(6484)));
    outputs(7364) <= layer2_outputs(10344);
    outputs(7365) <= layer2_outputs(12260);
    outputs(7366) <= layer2_outputs(4990);
    outputs(7367) <= (layer2_outputs(818)) xor (layer2_outputs(977));
    outputs(7368) <= not(layer2_outputs(6534));
    outputs(7369) <= (layer2_outputs(9797)) xor (layer2_outputs(12107));
    outputs(7370) <= (layer2_outputs(3106)) and not (layer2_outputs(3752));
    outputs(7371) <= layer2_outputs(7385);
    outputs(7372) <= (layer2_outputs(4237)) and not (layer2_outputs(639));
    outputs(7373) <= not(layer2_outputs(12539));
    outputs(7374) <= layer2_outputs(10288);
    outputs(7375) <= layer2_outputs(6499);
    outputs(7376) <= not((layer2_outputs(11827)) or (layer2_outputs(3332)));
    outputs(7377) <= (layer2_outputs(10995)) xor (layer2_outputs(3067));
    outputs(7378) <= layer2_outputs(4411);
    outputs(7379) <= layer2_outputs(3880);
    outputs(7380) <= not((layer2_outputs(2954)) xor (layer2_outputs(5960)));
    outputs(7381) <= not((layer2_outputs(3482)) xor (layer2_outputs(7143)));
    outputs(7382) <= layer2_outputs(4654);
    outputs(7383) <= (layer2_outputs(9945)) xor (layer2_outputs(12639));
    outputs(7384) <= not(layer2_outputs(11616));
    outputs(7385) <= not(layer2_outputs(9427));
    outputs(7386) <= not((layer2_outputs(7511)) xor (layer2_outputs(864)));
    outputs(7387) <= (layer2_outputs(2507)) xor (layer2_outputs(3534));
    outputs(7388) <= layer2_outputs(7968);
    outputs(7389) <= not(layer2_outputs(11785));
    outputs(7390) <= not(layer2_outputs(12255));
    outputs(7391) <= (layer2_outputs(1821)) and not (layer2_outputs(3664));
    outputs(7392) <= not(layer2_outputs(10890)) or (layer2_outputs(4668));
    outputs(7393) <= (layer2_outputs(9957)) xor (layer2_outputs(7503));
    outputs(7394) <= not(layer2_outputs(9748));
    outputs(7395) <= (layer2_outputs(6909)) xor (layer2_outputs(711));
    outputs(7396) <= layer2_outputs(10198);
    outputs(7397) <= not(layer2_outputs(5195)) or (layer2_outputs(1657));
    outputs(7398) <= (layer2_outputs(2743)) and (layer2_outputs(11690));
    outputs(7399) <= not((layer2_outputs(7091)) xor (layer2_outputs(9924)));
    outputs(7400) <= (layer2_outputs(10815)) xor (layer2_outputs(11515));
    outputs(7401) <= not((layer2_outputs(7321)) xor (layer2_outputs(4422)));
    outputs(7402) <= layer2_outputs(1485);
    outputs(7403) <= layer2_outputs(10980);
    outputs(7404) <= not(layer2_outputs(6771));
    outputs(7405) <= layer2_outputs(5382);
    outputs(7406) <= layer2_outputs(9988);
    outputs(7407) <= layer2_outputs(6372);
    outputs(7408) <= not(layer2_outputs(3096));
    outputs(7409) <= not(layer2_outputs(10773));
    outputs(7410) <= not(layer2_outputs(6808));
    outputs(7411) <= not((layer2_outputs(6850)) xor (layer2_outputs(11834)));
    outputs(7412) <= (layer2_outputs(4785)) xor (layer2_outputs(9421));
    outputs(7413) <= not(layer2_outputs(8962));
    outputs(7414) <= not(layer2_outputs(1555)) or (layer2_outputs(7697));
    outputs(7415) <= not((layer2_outputs(9534)) and (layer2_outputs(5946)));
    outputs(7416) <= not(layer2_outputs(10795));
    outputs(7417) <= not(layer2_outputs(4969)) or (layer2_outputs(8301));
    outputs(7418) <= not(layer2_outputs(8422));
    outputs(7419) <= not(layer2_outputs(2764));
    outputs(7420) <= (layer2_outputs(7075)) and not (layer2_outputs(699));
    outputs(7421) <= (layer2_outputs(9025)) xor (layer2_outputs(7876));
    outputs(7422) <= not(layer2_outputs(2266));
    outputs(7423) <= layer2_outputs(10887);
    outputs(7424) <= (layer2_outputs(11833)) xor (layer2_outputs(3477));
    outputs(7425) <= layer2_outputs(62);
    outputs(7426) <= not(layer2_outputs(5244));
    outputs(7427) <= layer2_outputs(5250);
    outputs(7428) <= not(layer2_outputs(2209));
    outputs(7429) <= layer2_outputs(245);
    outputs(7430) <= (layer2_outputs(3305)) or (layer2_outputs(6644));
    outputs(7431) <= (layer2_outputs(2392)) xor (layer2_outputs(8742));
    outputs(7432) <= not(layer2_outputs(11905));
    outputs(7433) <= layer2_outputs(11622);
    outputs(7434) <= (layer2_outputs(4739)) and not (layer2_outputs(1715));
    outputs(7435) <= not(layer2_outputs(1929));
    outputs(7436) <= not((layer2_outputs(9226)) and (layer2_outputs(11052)));
    outputs(7437) <= layer2_outputs(6170);
    outputs(7438) <= layer2_outputs(11390);
    outputs(7439) <= layer2_outputs(10046);
    outputs(7440) <= (layer2_outputs(8189)) xor (layer2_outputs(12219));
    outputs(7441) <= (layer2_outputs(3313)) or (layer2_outputs(912));
    outputs(7442) <= (layer2_outputs(3763)) xor (layer2_outputs(3317));
    outputs(7443) <= (layer2_outputs(2244)) xor (layer2_outputs(5794));
    outputs(7444) <= (layer2_outputs(7340)) and (layer2_outputs(7724));
    outputs(7445) <= (layer2_outputs(10041)) or (layer2_outputs(4797));
    outputs(7446) <= not(layer2_outputs(6461));
    outputs(7447) <= not(layer2_outputs(8657));
    outputs(7448) <= not(layer2_outputs(4292)) or (layer2_outputs(10569));
    outputs(7449) <= not(layer2_outputs(10897));
    outputs(7450) <= not((layer2_outputs(9359)) xor (layer2_outputs(2416)));
    outputs(7451) <= layer2_outputs(7318);
    outputs(7452) <= not(layer2_outputs(5230));
    outputs(7453) <= not((layer2_outputs(8576)) xor (layer2_outputs(5357)));
    outputs(7454) <= not(layer2_outputs(8962));
    outputs(7455) <= not(layer2_outputs(9993));
    outputs(7456) <= (layer2_outputs(6711)) xor (layer2_outputs(9653));
    outputs(7457) <= not(layer2_outputs(5231));
    outputs(7458) <= not(layer2_outputs(3721));
    outputs(7459) <= not((layer2_outputs(5214)) and (layer2_outputs(10144)));
    outputs(7460) <= not(layer2_outputs(3927));
    outputs(7461) <= layer2_outputs(4360);
    outputs(7462) <= not((layer2_outputs(8524)) xor (layer2_outputs(798)));
    outputs(7463) <= (layer2_outputs(2583)) xor (layer2_outputs(2711));
    outputs(7464) <= not(layer2_outputs(12432));
    outputs(7465) <= not(layer2_outputs(8286));
    outputs(7466) <= (layer2_outputs(4591)) and not (layer2_outputs(3979));
    outputs(7467) <= (layer2_outputs(6749)) xor (layer2_outputs(3641));
    outputs(7468) <= (layer2_outputs(514)) xor (layer2_outputs(424));
    outputs(7469) <= layer2_outputs(5692);
    outputs(7470) <= (layer2_outputs(8036)) xor (layer2_outputs(5824));
    outputs(7471) <= not((layer2_outputs(11995)) or (layer2_outputs(2556)));
    outputs(7472) <= layer2_outputs(37);
    outputs(7473) <= not(layer2_outputs(10762)) or (layer2_outputs(3186));
    outputs(7474) <= not((layer2_outputs(12344)) xor (layer2_outputs(2621)));
    outputs(7475) <= layer2_outputs(6637);
    outputs(7476) <= (layer2_outputs(5245)) xor (layer2_outputs(842));
    outputs(7477) <= (layer2_outputs(2880)) and (layer2_outputs(4319));
    outputs(7478) <= not((layer2_outputs(8171)) and (layer2_outputs(10823)));
    outputs(7479) <= layer2_outputs(3248);
    outputs(7480) <= layer2_outputs(11032);
    outputs(7481) <= not(layer2_outputs(4794));
    outputs(7482) <= layer2_outputs(8444);
    outputs(7483) <= (layer2_outputs(5631)) and not (layer2_outputs(11503));
    outputs(7484) <= not((layer2_outputs(8585)) xor (layer2_outputs(12753)));
    outputs(7485) <= not(layer2_outputs(5126));
    outputs(7486) <= not((layer2_outputs(5273)) xor (layer2_outputs(12151)));
    outputs(7487) <= not(layer2_outputs(913)) or (layer2_outputs(11715));
    outputs(7488) <= not(layer2_outputs(9616));
    outputs(7489) <= (layer2_outputs(11892)) xor (layer2_outputs(8983));
    outputs(7490) <= not(layer2_outputs(6695));
    outputs(7491) <= layer2_outputs(453);
    outputs(7492) <= layer2_outputs(4878);
    outputs(7493) <= layer2_outputs(12606);
    outputs(7494) <= (layer2_outputs(11347)) xor (layer2_outputs(7964));
    outputs(7495) <= layer2_outputs(9738);
    outputs(7496) <= not((layer2_outputs(5490)) or (layer2_outputs(4968)));
    outputs(7497) <= layer2_outputs(4444);
    outputs(7498) <= layer2_outputs(8115);
    outputs(7499) <= (layer2_outputs(7399)) xor (layer2_outputs(3398));
    outputs(7500) <= (layer2_outputs(4100)) and not (layer2_outputs(9343));
    outputs(7501) <= not(layer2_outputs(6899));
    outputs(7502) <= not((layer2_outputs(5025)) xor (layer2_outputs(3050)));
    outputs(7503) <= not((layer2_outputs(5110)) xor (layer2_outputs(3221)));
    outputs(7504) <= not((layer2_outputs(9650)) xor (layer2_outputs(3401)));
    outputs(7505) <= layer2_outputs(4035);
    outputs(7506) <= not(layer2_outputs(10179)) or (layer2_outputs(6716));
    outputs(7507) <= layer2_outputs(11764);
    outputs(7508) <= not(layer2_outputs(253));
    outputs(7509) <= layer2_outputs(3860);
    outputs(7510) <= layer2_outputs(6819);
    outputs(7511) <= not((layer2_outputs(10813)) xor (layer2_outputs(8448)));
    outputs(7512) <= not(layer2_outputs(12407));
    outputs(7513) <= not((layer2_outputs(3997)) xor (layer2_outputs(6081)));
    outputs(7514) <= not((layer2_outputs(1311)) xor (layer2_outputs(4667)));
    outputs(7515) <= layer2_outputs(11987);
    outputs(7516) <= layer2_outputs(710);
    outputs(7517) <= (layer2_outputs(4414)) xor (layer2_outputs(8201));
    outputs(7518) <= (layer2_outputs(1508)) xor (layer2_outputs(3981));
    outputs(7519) <= not((layer2_outputs(2814)) and (layer2_outputs(6301)));
    outputs(7520) <= not((layer2_outputs(11630)) xor (layer2_outputs(690)));
    outputs(7521) <= not(layer2_outputs(5457));
    outputs(7522) <= not(layer2_outputs(4178));
    outputs(7523) <= (layer2_outputs(11980)) xor (layer2_outputs(231));
    outputs(7524) <= layer2_outputs(12036);
    outputs(7525) <= (layer2_outputs(607)) and not (layer2_outputs(12051));
    outputs(7526) <= layer2_outputs(532);
    outputs(7527) <= (layer2_outputs(8352)) xor (layer2_outputs(1049));
    outputs(7528) <= layer2_outputs(12663);
    outputs(7529) <= (layer2_outputs(12794)) xor (layer2_outputs(7901));
    outputs(7530) <= not(layer2_outputs(6131));
    outputs(7531) <= not(layer2_outputs(5840)) or (layer2_outputs(11484));
    outputs(7532) <= layer2_outputs(8321);
    outputs(7533) <= not((layer2_outputs(7916)) xor (layer2_outputs(2495)));
    outputs(7534) <= not(layer2_outputs(5524));
    outputs(7535) <= not((layer2_outputs(741)) xor (layer2_outputs(9443)));
    outputs(7536) <= layer2_outputs(649);
    outputs(7537) <= not((layer2_outputs(10545)) xor (layer2_outputs(5412)));
    outputs(7538) <= (layer2_outputs(6227)) and not (layer2_outputs(3639));
    outputs(7539) <= not(layer2_outputs(3878));
    outputs(7540) <= not(layer2_outputs(8276));
    outputs(7541) <= not((layer2_outputs(1510)) xor (layer2_outputs(2361)));
    outputs(7542) <= layer2_outputs(444);
    outputs(7543) <= not(layer2_outputs(3523));
    outputs(7544) <= not((layer2_outputs(11131)) xor (layer2_outputs(7799)));
    outputs(7545) <= not(layer2_outputs(11347)) or (layer2_outputs(54));
    outputs(7546) <= (layer2_outputs(10806)) xor (layer2_outputs(8993));
    outputs(7547) <= not(layer2_outputs(10107));
    outputs(7548) <= not((layer2_outputs(1018)) xor (layer2_outputs(12224)));
    outputs(7549) <= not(layer2_outputs(4844));
    outputs(7550) <= layer2_outputs(4621);
    outputs(7551) <= layer2_outputs(6969);
    outputs(7552) <= layer2_outputs(4429);
    outputs(7553) <= layer2_outputs(2344);
    outputs(7554) <= (layer2_outputs(3775)) xor (layer2_outputs(545));
    outputs(7555) <= not(layer2_outputs(8116));
    outputs(7556) <= layer2_outputs(6759);
    outputs(7557) <= (layer2_outputs(1167)) xor (layer2_outputs(4125));
    outputs(7558) <= not(layer2_outputs(10658)) or (layer2_outputs(1427));
    outputs(7559) <= not(layer2_outputs(8534));
    outputs(7560) <= not(layer2_outputs(5265));
    outputs(7561) <= not((layer2_outputs(11153)) xor (layer2_outputs(7335)));
    outputs(7562) <= (layer2_outputs(418)) xor (layer2_outputs(1443));
    outputs(7563) <= (layer2_outputs(1905)) xor (layer2_outputs(9465));
    outputs(7564) <= not(layer2_outputs(7536));
    outputs(7565) <= not(layer2_outputs(3797));
    outputs(7566) <= (layer2_outputs(9242)) and not (layer2_outputs(11519));
    outputs(7567) <= layer2_outputs(2737);
    outputs(7568) <= not(layer2_outputs(9618));
    outputs(7569) <= layer2_outputs(12681);
    outputs(7570) <= not((layer2_outputs(5396)) xor (layer2_outputs(2098)));
    outputs(7571) <= not(layer2_outputs(8400));
    outputs(7572) <= (layer2_outputs(7308)) xor (layer2_outputs(3022));
    outputs(7573) <= not(layer2_outputs(9387));
    outputs(7574) <= not(layer2_outputs(1024)) or (layer2_outputs(10219));
    outputs(7575) <= layer2_outputs(9968);
    outputs(7576) <= not(layer2_outputs(8055));
    outputs(7577) <= (layer2_outputs(3501)) xor (layer2_outputs(7228));
    outputs(7578) <= not(layer2_outputs(10002)) or (layer2_outputs(4668));
    outputs(7579) <= (layer2_outputs(7333)) xor (layer2_outputs(12722));
    outputs(7580) <= layer2_outputs(11336);
    outputs(7581) <= not(layer2_outputs(11187));
    outputs(7582) <= layer2_outputs(11443);
    outputs(7583) <= not(layer2_outputs(8812));
    outputs(7584) <= layer2_outputs(8851);
    outputs(7585) <= not(layer2_outputs(12785));
    outputs(7586) <= (layer2_outputs(8403)) xor (layer2_outputs(948));
    outputs(7587) <= layer2_outputs(4288);
    outputs(7588) <= not((layer2_outputs(10735)) and (layer2_outputs(5878)));
    outputs(7589) <= not((layer2_outputs(11489)) xor (layer2_outputs(3740)));
    outputs(7590) <= not(layer2_outputs(9581));
    outputs(7591) <= layer2_outputs(11082);
    outputs(7592) <= not((layer2_outputs(6509)) and (layer2_outputs(7887)));
    outputs(7593) <= not((layer2_outputs(1372)) and (layer2_outputs(9911)));
    outputs(7594) <= not(layer2_outputs(1493)) or (layer2_outputs(6587));
    outputs(7595) <= not((layer2_outputs(10950)) and (layer2_outputs(2012)));
    outputs(7596) <= not(layer2_outputs(6977)) or (layer2_outputs(12132));
    outputs(7597) <= layer2_outputs(7435);
    outputs(7598) <= layer2_outputs(12092);
    outputs(7599) <= not(layer2_outputs(4901));
    outputs(7600) <= not(layer2_outputs(8517));
    outputs(7601) <= not(layer2_outputs(8037));
    outputs(7602) <= (layer2_outputs(9383)) xor (layer2_outputs(4699));
    outputs(7603) <= not(layer2_outputs(6951));
    outputs(7604) <= (layer2_outputs(7865)) and (layer2_outputs(9591));
    outputs(7605) <= not(layer2_outputs(10956));
    outputs(7606) <= layer2_outputs(3959);
    outputs(7607) <= layer2_outputs(12005);
    outputs(7608) <= layer2_outputs(12789);
    outputs(7609) <= layer2_outputs(11904);
    outputs(7610) <= (layer2_outputs(6967)) xor (layer2_outputs(2205));
    outputs(7611) <= (layer2_outputs(8792)) and not (layer2_outputs(5697));
    outputs(7612) <= not((layer2_outputs(3853)) or (layer2_outputs(6832)));
    outputs(7613) <= (layer2_outputs(8084)) xor (layer2_outputs(1634));
    outputs(7614) <= not(layer2_outputs(6927));
    outputs(7615) <= not(layer2_outputs(11170));
    outputs(7616) <= not(layer2_outputs(7426));
    outputs(7617) <= layer2_outputs(9034);
    outputs(7618) <= (layer2_outputs(7083)) xor (layer2_outputs(8542));
    outputs(7619) <= not((layer2_outputs(1813)) xor (layer2_outputs(6907)));
    outputs(7620) <= not(layer2_outputs(11746));
    outputs(7621) <= (layer2_outputs(5853)) xor (layer2_outputs(10043));
    outputs(7622) <= not((layer2_outputs(7537)) and (layer2_outputs(10503)));
    outputs(7623) <= not((layer2_outputs(5568)) xor (layer2_outputs(4084)));
    outputs(7624) <= layer2_outputs(10798);
    outputs(7625) <= not(layer2_outputs(8670));
    outputs(7626) <= layer2_outputs(4997);
    outputs(7627) <= (layer2_outputs(9605)) xor (layer2_outputs(9634));
    outputs(7628) <= (layer2_outputs(6704)) xor (layer2_outputs(4250));
    outputs(7629) <= layer2_outputs(1053);
    outputs(7630) <= layer2_outputs(732);
    outputs(7631) <= layer2_outputs(577);
    outputs(7632) <= (layer2_outputs(1501)) xor (layer2_outputs(5093));
    outputs(7633) <= (layer2_outputs(11593)) and not (layer2_outputs(3750));
    outputs(7634) <= (layer2_outputs(5018)) xor (layer2_outputs(430));
    outputs(7635) <= not(layer2_outputs(3924));
    outputs(7636) <= layer2_outputs(673);
    outputs(7637) <= (layer2_outputs(10400)) xor (layer2_outputs(9166));
    outputs(7638) <= not(layer2_outputs(2389));
    outputs(7639) <= (layer2_outputs(5458)) xor (layer2_outputs(10026));
    outputs(7640) <= (layer2_outputs(9992)) and not (layer2_outputs(4771));
    outputs(7641) <= (layer2_outputs(6295)) xor (layer2_outputs(1820));
    outputs(7642) <= (layer2_outputs(4401)) xor (layer2_outputs(10474));
    outputs(7643) <= (layer2_outputs(11700)) xor (layer2_outputs(11149));
    outputs(7644) <= not(layer2_outputs(4670));
    outputs(7645) <= (layer2_outputs(7721)) and not (layer2_outputs(1732));
    outputs(7646) <= layer2_outputs(3430);
    outputs(7647) <= layer2_outputs(9206);
    outputs(7648) <= (layer2_outputs(10072)) xor (layer2_outputs(9012));
    outputs(7649) <= layer2_outputs(2510);
    outputs(7650) <= (layer2_outputs(1863)) xor (layer2_outputs(11780));
    outputs(7651) <= not((layer2_outputs(10845)) or (layer2_outputs(1188)));
    outputs(7652) <= not((layer2_outputs(9327)) xor (layer2_outputs(4491)));
    outputs(7653) <= layer2_outputs(3354);
    outputs(7654) <= (layer2_outputs(5710)) and not (layer2_outputs(1729));
    outputs(7655) <= not(layer2_outputs(8353));
    outputs(7656) <= (layer2_outputs(1626)) and not (layer2_outputs(4544));
    outputs(7657) <= layer2_outputs(11526);
    outputs(7658) <= not((layer2_outputs(6909)) xor (layer2_outputs(12202)));
    outputs(7659) <= layer2_outputs(7849);
    outputs(7660) <= not((layer2_outputs(3088)) xor (layer2_outputs(9214)));
    outputs(7661) <= (layer2_outputs(5281)) xor (layer2_outputs(10121));
    outputs(7662) <= not((layer2_outputs(1256)) xor (layer2_outputs(5734)));
    outputs(7663) <= not(layer2_outputs(2485));
    outputs(7664) <= not(layer2_outputs(8349));
    outputs(7665) <= layer2_outputs(8763);
    outputs(7666) <= layer2_outputs(8813);
    outputs(7667) <= layer2_outputs(11703);
    outputs(7668) <= layer2_outputs(12501);
    outputs(7669) <= layer2_outputs(1659);
    outputs(7670) <= not(layer2_outputs(11261)) or (layer2_outputs(6868));
    outputs(7671) <= not((layer2_outputs(1560)) xor (layer2_outputs(2232)));
    outputs(7672) <= (layer2_outputs(7943)) and not (layer2_outputs(6306));
    outputs(7673) <= not(layer2_outputs(10051)) or (layer2_outputs(11903));
    outputs(7674) <= layer2_outputs(12216);
    outputs(7675) <= not((layer2_outputs(4445)) xor (layer2_outputs(5059)));
    outputs(7676) <= not(layer2_outputs(11384));
    outputs(7677) <= layer2_outputs(10889);
    outputs(7678) <= layer2_outputs(9898);
    outputs(7679) <= not(layer2_outputs(7703));
    outputs(7680) <= layer2_outputs(9212);
    outputs(7681) <= layer2_outputs(10775);
    outputs(7682) <= not(layer2_outputs(1933));
    outputs(7683) <= (layer2_outputs(2928)) xor (layer2_outputs(6847));
    outputs(7684) <= layer2_outputs(11767);
    outputs(7685) <= layer2_outputs(5029);
    outputs(7686) <= layer2_outputs(6376);
    outputs(7687) <= not(layer2_outputs(6178));
    outputs(7688) <= layer2_outputs(5152);
    outputs(7689) <= not(layer2_outputs(10130));
    outputs(7690) <= not(layer2_outputs(413));
    outputs(7691) <= not(layer2_outputs(7908));
    outputs(7692) <= not(layer2_outputs(2239));
    outputs(7693) <= not(layer2_outputs(9286)) or (layer2_outputs(7248));
    outputs(7694) <= not(layer2_outputs(7511)) or (layer2_outputs(551));
    outputs(7695) <= (layer2_outputs(7419)) xor (layer2_outputs(5895));
    outputs(7696) <= not((layer2_outputs(12385)) and (layer2_outputs(823)));
    outputs(7697) <= layer2_outputs(6487);
    outputs(7698) <= layer2_outputs(12509);
    outputs(7699) <= (layer2_outputs(1939)) and (layer2_outputs(100));
    outputs(7700) <= not(layer2_outputs(11962));
    outputs(7701) <= (layer2_outputs(1452)) xor (layer2_outputs(3911));
    outputs(7702) <= (layer2_outputs(6872)) and not (layer2_outputs(4563));
    outputs(7703) <= not(layer2_outputs(4421));
    outputs(7704) <= layer2_outputs(4281);
    outputs(7705) <= not(layer2_outputs(5710));
    outputs(7706) <= (layer2_outputs(4039)) and not (layer2_outputs(4082));
    outputs(7707) <= layer2_outputs(4405);
    outputs(7708) <= not(layer2_outputs(3156));
    outputs(7709) <= layer2_outputs(10610);
    outputs(7710) <= layer2_outputs(10952);
    outputs(7711) <= layer2_outputs(4791);
    outputs(7712) <= layer2_outputs(12530);
    outputs(7713) <= (layer2_outputs(1213)) and not (layer2_outputs(5092));
    outputs(7714) <= (layer2_outputs(9934)) xor (layer2_outputs(218));
    outputs(7715) <= not(layer2_outputs(2331));
    outputs(7716) <= layer2_outputs(6334);
    outputs(7717) <= layer2_outputs(1972);
    outputs(7718) <= layer2_outputs(2354);
    outputs(7719) <= not(layer2_outputs(4766));
    outputs(7720) <= layer2_outputs(6846);
    outputs(7721) <= not((layer2_outputs(11750)) and (layer2_outputs(2668)));
    outputs(7722) <= not(layer2_outputs(5729)) or (layer2_outputs(12467));
    outputs(7723) <= not((layer2_outputs(36)) xor (layer2_outputs(6437)));
    outputs(7724) <= not(layer2_outputs(12519));
    outputs(7725) <= (layer2_outputs(11623)) and not (layer2_outputs(11743));
    outputs(7726) <= not((layer2_outputs(8890)) xor (layer2_outputs(4298)));
    outputs(7727) <= layer2_outputs(12219);
    outputs(7728) <= (layer2_outputs(6391)) and (layer2_outputs(10619));
    outputs(7729) <= layer2_outputs(7365);
    outputs(7730) <= not(layer2_outputs(12455));
    outputs(7731) <= not(layer2_outputs(8831));
    outputs(7732) <= not((layer2_outputs(3257)) xor (layer2_outputs(12152)));
    outputs(7733) <= layer2_outputs(4169);
    outputs(7734) <= not(layer2_outputs(8558));
    outputs(7735) <= (layer2_outputs(8535)) and not (layer2_outputs(8371));
    outputs(7736) <= not(layer2_outputs(6549));
    outputs(7737) <= not(layer2_outputs(11161));
    outputs(7738) <= not(layer2_outputs(10248));
    outputs(7739) <= layer2_outputs(7271);
    outputs(7740) <= not(layer2_outputs(4112));
    outputs(7741) <= not(layer2_outputs(3577));
    outputs(7742) <= not((layer2_outputs(5615)) xor (layer2_outputs(6168)));
    outputs(7743) <= layer2_outputs(7784);
    outputs(7744) <= (layer2_outputs(12710)) and (layer2_outputs(267));
    outputs(7745) <= not(layer2_outputs(2858)) or (layer2_outputs(8980));
    outputs(7746) <= layer2_outputs(702);
    outputs(7747) <= layer2_outputs(1029);
    outputs(7748) <= layer2_outputs(4912);
    outputs(7749) <= layer2_outputs(590);
    outputs(7750) <= (layer2_outputs(11773)) and (layer2_outputs(4995));
    outputs(7751) <= not(layer2_outputs(11537));
    outputs(7752) <= not((layer2_outputs(3528)) xor (layer2_outputs(4633)));
    outputs(7753) <= not(layer2_outputs(6848));
    outputs(7754) <= layer2_outputs(11688);
    outputs(7755) <= (layer2_outputs(414)) xor (layer2_outputs(4945));
    outputs(7756) <= not(layer2_outputs(9805));
    outputs(7757) <= layer2_outputs(4821);
    outputs(7758) <= not(layer2_outputs(4480));
    outputs(7759) <= not((layer2_outputs(9575)) or (layer2_outputs(3124)));
    outputs(7760) <= layer2_outputs(6536);
    outputs(7761) <= not(layer2_outputs(11400)) or (layer2_outputs(1848));
    outputs(7762) <= not(layer2_outputs(10853));
    outputs(7763) <= not((layer2_outputs(9347)) xor (layer2_outputs(11836)));
    outputs(7764) <= layer2_outputs(8057);
    outputs(7765) <= layer2_outputs(10370);
    outputs(7766) <= layer2_outputs(10418);
    outputs(7767) <= layer2_outputs(3647);
    outputs(7768) <= layer2_outputs(8685);
    outputs(7769) <= layer2_outputs(3921);
    outputs(7770) <= layer2_outputs(6440);
    outputs(7771) <= not((layer2_outputs(219)) xor (layer2_outputs(4514)));
    outputs(7772) <= (layer2_outputs(1061)) and not (layer2_outputs(9758));
    outputs(7773) <= not(layer2_outputs(8318));
    outputs(7774) <= not(layer2_outputs(6263)) or (layer2_outputs(3740));
    outputs(7775) <= (layer2_outputs(10380)) and not (layer2_outputs(12610));
    outputs(7776) <= not((layer2_outputs(2370)) and (layer2_outputs(6275)));
    outputs(7777) <= (layer2_outputs(10824)) and not (layer2_outputs(4982));
    outputs(7778) <= layer2_outputs(3767);
    outputs(7779) <= not(layer2_outputs(6587));
    outputs(7780) <= layer2_outputs(6780);
    outputs(7781) <= (layer2_outputs(94)) xor (layer2_outputs(483));
    outputs(7782) <= layer2_outputs(6613);
    outputs(7783) <= not(layer2_outputs(5437));
    outputs(7784) <= not((layer2_outputs(7796)) xor (layer2_outputs(4530)));
    outputs(7785) <= not(layer2_outputs(1002));
    outputs(7786) <= not(layer2_outputs(4503));
    outputs(7787) <= not(layer2_outputs(10431));
    outputs(7788) <= not(layer2_outputs(11602));
    outputs(7789) <= not(layer2_outputs(11556));
    outputs(7790) <= not(layer2_outputs(10536));
    outputs(7791) <= layer2_outputs(330);
    outputs(7792) <= not(layer2_outputs(12294));
    outputs(7793) <= not(layer2_outputs(8013)) or (layer2_outputs(2186));
    outputs(7794) <= not(layer2_outputs(9825));
    outputs(7795) <= layer2_outputs(12404);
    outputs(7796) <= layer2_outputs(6460);
    outputs(7797) <= not(layer2_outputs(11944));
    outputs(7798) <= layer2_outputs(12391);
    outputs(7799) <= (layer2_outputs(11921)) xor (layer2_outputs(9253));
    outputs(7800) <= (layer2_outputs(1069)) xor (layer2_outputs(305));
    outputs(7801) <= layer2_outputs(9523);
    outputs(7802) <= layer2_outputs(8365);
    outputs(7803) <= (layer2_outputs(4769)) xor (layer2_outputs(8838));
    outputs(7804) <= (layer2_outputs(3365)) xor (layer2_outputs(5283));
    outputs(7805) <= (layer2_outputs(10190)) and not (layer2_outputs(3887));
    outputs(7806) <= not(layer2_outputs(12394));
    outputs(7807) <= not(layer2_outputs(884));
    outputs(7808) <= layer2_outputs(12427);
    outputs(7809) <= not(layer2_outputs(4147));
    outputs(7810) <= (layer2_outputs(11027)) and not (layer2_outputs(9736));
    outputs(7811) <= layer2_outputs(5967);
    outputs(7812) <= not((layer2_outputs(8682)) or (layer2_outputs(6167)));
    outputs(7813) <= (layer2_outputs(3222)) and (layer2_outputs(8857));
    outputs(7814) <= layer2_outputs(1561);
    outputs(7815) <= (layer2_outputs(2379)) xor (layer2_outputs(1362));
    outputs(7816) <= not((layer2_outputs(3051)) xor (layer2_outputs(3277)));
    outputs(7817) <= (layer2_outputs(9419)) and not (layer2_outputs(752));
    outputs(7818) <= not((layer2_outputs(2666)) and (layer2_outputs(1367)));
    outputs(7819) <= (layer2_outputs(6931)) and not (layer2_outputs(2115));
    outputs(7820) <= (layer2_outputs(1587)) and not (layer2_outputs(12555));
    outputs(7821) <= not((layer2_outputs(7510)) xor (layer2_outputs(7561)));
    outputs(7822) <= not(layer2_outputs(7468));
    outputs(7823) <= layer2_outputs(7418);
    outputs(7824) <= not(layer2_outputs(12638));
    outputs(7825) <= not(layer2_outputs(5726));
    outputs(7826) <= not(layer2_outputs(437)) or (layer2_outputs(11741));
    outputs(7827) <= not(layer2_outputs(5192));
    outputs(7828) <= layer2_outputs(3351);
    outputs(7829) <= not(layer2_outputs(6141));
    outputs(7830) <= (layer2_outputs(9763)) and not (layer2_outputs(2226));
    outputs(7831) <= layer2_outputs(12120);
    outputs(7832) <= not(layer2_outputs(12111));
    outputs(7833) <= not((layer2_outputs(4284)) and (layer2_outputs(7298)));
    outputs(7834) <= not((layer2_outputs(12755)) xor (layer2_outputs(8559)));
    outputs(7835) <= layer2_outputs(9293);
    outputs(7836) <= not((layer2_outputs(5340)) or (layer2_outputs(12289)));
    outputs(7837) <= (layer2_outputs(11805)) and (layer2_outputs(2470));
    outputs(7838) <= layer2_outputs(19);
    outputs(7839) <= (layer2_outputs(1195)) or (layer2_outputs(2825));
    outputs(7840) <= (layer2_outputs(11898)) and (layer2_outputs(7346));
    outputs(7841) <= (layer2_outputs(6670)) xor (layer2_outputs(6063));
    outputs(7842) <= not(layer2_outputs(1725));
    outputs(7843) <= (layer2_outputs(8456)) xor (layer2_outputs(8061));
    outputs(7844) <= not((layer2_outputs(12106)) xor (layer2_outputs(9559)));
    outputs(7845) <= not(layer2_outputs(1588));
    outputs(7846) <= layer2_outputs(7299);
    outputs(7847) <= not((layer2_outputs(10761)) xor (layer2_outputs(194)));
    outputs(7848) <= not(layer2_outputs(7924));
    outputs(7849) <= layer2_outputs(1561);
    outputs(7850) <= not(layer2_outputs(5687));
    outputs(7851) <= (layer2_outputs(2579)) xor (layer2_outputs(858));
    outputs(7852) <= layer2_outputs(336);
    outputs(7853) <= not(layer2_outputs(5998));
    outputs(7854) <= not((layer2_outputs(4949)) xor (layer2_outputs(5995)));
    outputs(7855) <= layer2_outputs(11613);
    outputs(7856) <= (layer2_outputs(1424)) and not (layer2_outputs(1152));
    outputs(7857) <= layer2_outputs(4719);
    outputs(7858) <= not((layer2_outputs(9184)) xor (layer2_outputs(12674)));
    outputs(7859) <= not((layer2_outputs(8767)) and (layer2_outputs(6768)));
    outputs(7860) <= layer2_outputs(11483);
    outputs(7861) <= not(layer2_outputs(738)) or (layer2_outputs(2354));
    outputs(7862) <= (layer2_outputs(5370)) and not (layer2_outputs(9507));
    outputs(7863) <= layer2_outputs(4028);
    outputs(7864) <= layer2_outputs(6788);
    outputs(7865) <= layer2_outputs(11333);
    outputs(7866) <= layer2_outputs(7129);
    outputs(7867) <= (layer2_outputs(12530)) or (layer2_outputs(11577));
    outputs(7868) <= not((layer2_outputs(3331)) xor (layer2_outputs(3249)));
    outputs(7869) <= layer2_outputs(591);
    outputs(7870) <= layer2_outputs(9584);
    outputs(7871) <= layer2_outputs(3037);
    outputs(7872) <= not(layer2_outputs(8335));
    outputs(7873) <= layer2_outputs(899);
    outputs(7874) <= not(layer2_outputs(7380));
    outputs(7875) <= (layer2_outputs(8519)) and (layer2_outputs(11972));
    outputs(7876) <= not(layer2_outputs(7755));
    outputs(7877) <= not(layer2_outputs(11850));
    outputs(7878) <= layer2_outputs(1834);
    outputs(7879) <= (layer2_outputs(8422)) or (layer2_outputs(4346));
    outputs(7880) <= not(layer2_outputs(6793));
    outputs(7881) <= layer2_outputs(6823);
    outputs(7882) <= not((layer2_outputs(11503)) xor (layer2_outputs(11078)));
    outputs(7883) <= not(layer2_outputs(2422));
    outputs(7884) <= layer2_outputs(2533);
    outputs(7885) <= (layer2_outputs(2824)) xor (layer2_outputs(8043));
    outputs(7886) <= (layer2_outputs(9718)) and not (layer2_outputs(7620));
    outputs(7887) <= layer2_outputs(193);
    outputs(7888) <= layer2_outputs(11759);
    outputs(7889) <= (layer2_outputs(9558)) and (layer2_outputs(11181));
    outputs(7890) <= not(layer2_outputs(6564));
    outputs(7891) <= not(layer2_outputs(4448));
    outputs(7892) <= not((layer2_outputs(12676)) xor (layer2_outputs(4915)));
    outputs(7893) <= (layer2_outputs(11513)) and not (layer2_outputs(8564));
    outputs(7894) <= (layer2_outputs(1528)) xor (layer2_outputs(1216));
    outputs(7895) <= not((layer2_outputs(10721)) xor (layer2_outputs(5871)));
    outputs(7896) <= not(layer2_outputs(2279));
    outputs(7897) <= not((layer2_outputs(10831)) or (layer2_outputs(9395)));
    outputs(7898) <= not((layer2_outputs(1028)) xor (layer2_outputs(1300)));
    outputs(7899) <= not(layer2_outputs(2130)) or (layer2_outputs(2298));
    outputs(7900) <= not(layer2_outputs(6664));
    outputs(7901) <= not(layer2_outputs(9458));
    outputs(7902) <= not(layer2_outputs(7386));
    outputs(7903) <= not(layer2_outputs(1236));
    outputs(7904) <= layer2_outputs(700);
    outputs(7905) <= not(layer2_outputs(2617));
    outputs(7906) <= (layer2_outputs(8857)) and (layer2_outputs(7405));
    outputs(7907) <= not(layer2_outputs(12612));
    outputs(7908) <= (layer2_outputs(12216)) xor (layer2_outputs(11050));
    outputs(7909) <= not((layer2_outputs(3054)) or (layer2_outputs(4525)));
    outputs(7910) <= not(layer2_outputs(7187));
    outputs(7911) <= not((layer2_outputs(5780)) xor (layer2_outputs(1488)));
    outputs(7912) <= not(layer2_outputs(9218));
    outputs(7913) <= not(layer2_outputs(4559));
    outputs(7914) <= not(layer2_outputs(11270));
    outputs(7915) <= not(layer2_outputs(8499));
    outputs(7916) <= layer2_outputs(9244);
    outputs(7917) <= layer2_outputs(6440);
    outputs(7918) <= layer2_outputs(6014);
    outputs(7919) <= not(layer2_outputs(12539));
    outputs(7920) <= not(layer2_outputs(3798));
    outputs(7921) <= not(layer2_outputs(5992));
    outputs(7922) <= layer2_outputs(3174);
    outputs(7923) <= not(layer2_outputs(8171)) or (layer2_outputs(9045));
    outputs(7924) <= layer2_outputs(1217);
    outputs(7925) <= not(layer2_outputs(4520));
    outputs(7926) <= not(layer2_outputs(5462));
    outputs(7927) <= not(layer2_outputs(8897));
    outputs(7928) <= not(layer2_outputs(4372));
    outputs(7929) <= layer2_outputs(5118);
    outputs(7930) <= (layer2_outputs(11927)) and not (layer2_outputs(9120));
    outputs(7931) <= not((layer2_outputs(6236)) xor (layer2_outputs(11728)));
    outputs(7932) <= not(layer2_outputs(10756));
    outputs(7933) <= not(layer2_outputs(9504));
    outputs(7934) <= layer2_outputs(11305);
    outputs(7935) <= not(layer2_outputs(6439));
    outputs(7936) <= not((layer2_outputs(7134)) and (layer2_outputs(8259)));
    outputs(7937) <= not(layer2_outputs(1465));
    outputs(7938) <= not(layer2_outputs(8915)) or (layer2_outputs(837));
    outputs(7939) <= layer2_outputs(11572);
    outputs(7940) <= not((layer2_outputs(9948)) or (layer2_outputs(5190)));
    outputs(7941) <= layer2_outputs(6687);
    outputs(7942) <= not(layer2_outputs(5185)) or (layer2_outputs(12503));
    outputs(7943) <= (layer2_outputs(10263)) and not (layer2_outputs(7969));
    outputs(7944) <= layer2_outputs(5858);
    outputs(7945) <= not(layer2_outputs(7707));
    outputs(7946) <= layer2_outputs(10271);
    outputs(7947) <= not((layer2_outputs(12)) xor (layer2_outputs(11977)));
    outputs(7948) <= layer2_outputs(7316);
    outputs(7949) <= layer2_outputs(1139);
    outputs(7950) <= (layer2_outputs(954)) and not (layer2_outputs(6118));
    outputs(7951) <= layer2_outputs(12649);
    outputs(7952) <= layer2_outputs(9283);
    outputs(7953) <= not(layer2_outputs(4919));
    outputs(7954) <= (layer2_outputs(11572)) and not (layer2_outputs(9880));
    outputs(7955) <= not(layer2_outputs(10951));
    outputs(7956) <= (layer2_outputs(12521)) xor (layer2_outputs(6576));
    outputs(7957) <= layer2_outputs(3481);
    outputs(7958) <= not(layer2_outputs(11010));
    outputs(7959) <= not((layer2_outputs(3385)) xor (layer2_outputs(1138)));
    outputs(7960) <= not(layer2_outputs(11129)) or (layer2_outputs(1129));
    outputs(7961) <= not(layer2_outputs(4109));
    outputs(7962) <= layer2_outputs(2258);
    outputs(7963) <= (layer2_outputs(12760)) and (layer2_outputs(5590));
    outputs(7964) <= not(layer2_outputs(4613));
    outputs(7965) <= not(layer2_outputs(5965));
    outputs(7966) <= (layer2_outputs(10920)) xor (layer2_outputs(9913));
    outputs(7967) <= not((layer2_outputs(11506)) xor (layer2_outputs(4980)));
    outputs(7968) <= not(layer2_outputs(7967));
    outputs(7969) <= (layer2_outputs(6803)) and (layer2_outputs(5777));
    outputs(7970) <= not((layer2_outputs(5190)) or (layer2_outputs(2048)));
    outputs(7971) <= not(layer2_outputs(2404));
    outputs(7972) <= layer2_outputs(2067);
    outputs(7973) <= not(layer2_outputs(1487));
    outputs(7974) <= layer2_outputs(10333);
    outputs(7975) <= layer2_outputs(8858);
    outputs(7976) <= '0';
    outputs(7977) <= not(layer2_outputs(10766));
    outputs(7978) <= layer2_outputs(8661);
    outputs(7979) <= layer2_outputs(12336);
    outputs(7980) <= not(layer2_outputs(8243));
    outputs(7981) <= layer2_outputs(4892);
    outputs(7982) <= (layer2_outputs(10592)) xor (layer2_outputs(7074));
    outputs(7983) <= not(layer2_outputs(11978));
    outputs(7984) <= not(layer2_outputs(6544));
    outputs(7985) <= not(layer2_outputs(2777));
    outputs(7986) <= layer2_outputs(7601);
    outputs(7987) <= layer2_outputs(10066);
    outputs(7988) <= not(layer2_outputs(9194));
    outputs(7989) <= (layer2_outputs(8854)) xor (layer2_outputs(8028));
    outputs(7990) <= (layer2_outputs(11450)) and not (layer2_outputs(5282));
    outputs(7991) <= (layer2_outputs(285)) and (layer2_outputs(8465));
    outputs(7992) <= not(layer2_outputs(9847));
    outputs(7993) <= not((layer2_outputs(3600)) and (layer2_outputs(855)));
    outputs(7994) <= not((layer2_outputs(8510)) xor (layer2_outputs(8433)));
    outputs(7995) <= layer2_outputs(10257);
    outputs(7996) <= layer2_outputs(589);
    outputs(7997) <= (layer2_outputs(11811)) or (layer2_outputs(9065));
    outputs(7998) <= (layer2_outputs(10471)) and not (layer2_outputs(8244));
    outputs(7999) <= not(layer2_outputs(5431));
    outputs(8000) <= (layer2_outputs(3651)) xor (layer2_outputs(8656));
    outputs(8001) <= layer2_outputs(12574);
    outputs(8002) <= layer2_outputs(11447);
    outputs(8003) <= not((layer2_outputs(3280)) xor (layer2_outputs(7355)));
    outputs(8004) <= not(layer2_outputs(537)) or (layer2_outputs(11587));
    outputs(8005) <= not(layer2_outputs(5937));
    outputs(8006) <= layer2_outputs(939);
    outputs(8007) <= layer2_outputs(12044);
    outputs(8008) <= layer2_outputs(950);
    outputs(8009) <= (layer2_outputs(7770)) and not (layer2_outputs(5803));
    outputs(8010) <= layer2_outputs(332);
    outputs(8011) <= not((layer2_outputs(5260)) xor (layer2_outputs(2114)));
    outputs(8012) <= not((layer2_outputs(517)) or (layer2_outputs(8623)));
    outputs(8013) <= not(layer2_outputs(132));
    outputs(8014) <= not(layer2_outputs(310));
    outputs(8015) <= layer2_outputs(1184);
    outputs(8016) <= not(layer2_outputs(2512));
    outputs(8017) <= layer2_outputs(4780);
    outputs(8018) <= not(layer2_outputs(224));
    outputs(8019) <= not(layer2_outputs(746));
    outputs(8020) <= not(layer2_outputs(5651)) or (layer2_outputs(6622));
    outputs(8021) <= not((layer2_outputs(11481)) xor (layer2_outputs(1993)));
    outputs(8022) <= layer2_outputs(5293);
    outputs(8023) <= not(layer2_outputs(11598));
    outputs(8024) <= (layer2_outputs(11273)) xor (layer2_outputs(1441));
    outputs(8025) <= not(layer2_outputs(2751)) or (layer2_outputs(11063));
    outputs(8026) <= not(layer2_outputs(663));
    outputs(8027) <= not((layer2_outputs(4541)) xor (layer2_outputs(5545)));
    outputs(8028) <= layer2_outputs(6188);
    outputs(8029) <= not(layer2_outputs(5780)) or (layer2_outputs(9297));
    outputs(8030) <= not(layer2_outputs(7671));
    outputs(8031) <= not(layer2_outputs(12609));
    outputs(8032) <= not(layer2_outputs(1943));
    outputs(8033) <= not((layer2_outputs(7452)) xor (layer2_outputs(3913)));
    outputs(8034) <= not(layer2_outputs(3451));
    outputs(8035) <= layer2_outputs(2910);
    outputs(8036) <= not(layer2_outputs(7652));
    outputs(8037) <= layer2_outputs(8027);
    outputs(8038) <= not((layer2_outputs(263)) or (layer2_outputs(12431)));
    outputs(8039) <= layer2_outputs(11639);
    outputs(8040) <= not(layer2_outputs(5469));
    outputs(8041) <= not(layer2_outputs(8039));
    outputs(8042) <= not(layer2_outputs(8255));
    outputs(8043) <= (layer2_outputs(5483)) and not (layer2_outputs(502));
    outputs(8044) <= layer2_outputs(8210);
    outputs(8045) <= not(layer2_outputs(9335));
    outputs(8046) <= not(layer2_outputs(8988));
    outputs(8047) <= not((layer2_outputs(7349)) or (layer2_outputs(3846)));
    outputs(8048) <= not(layer2_outputs(9054));
    outputs(8049) <= not(layer2_outputs(1823));
    outputs(8050) <= layer2_outputs(1495);
    outputs(8051) <= layer2_outputs(1311);
    outputs(8052) <= not(layer2_outputs(6264));
    outputs(8053) <= layer2_outputs(3622);
    outputs(8054) <= not((layer2_outputs(8271)) xor (layer2_outputs(781)));
    outputs(8055) <= (layer2_outputs(10077)) and not (layer2_outputs(11379));
    outputs(8056) <= not(layer2_outputs(12292));
    outputs(8057) <= not(layer2_outputs(11233));
    outputs(8058) <= not(layer2_outputs(6364));
    outputs(8059) <= (layer2_outputs(10298)) and (layer2_outputs(2018));
    outputs(8060) <= layer2_outputs(9740);
    outputs(8061) <= (layer2_outputs(2534)) xor (layer2_outputs(5425));
    outputs(8062) <= (layer2_outputs(7000)) and not (layer2_outputs(2256));
    outputs(8063) <= not(layer2_outputs(9121));
    outputs(8064) <= not(layer2_outputs(2112));
    outputs(8065) <= layer2_outputs(675);
    outputs(8066) <= not((layer2_outputs(10365)) xor (layer2_outputs(348)));
    outputs(8067) <= not(layer2_outputs(1692));
    outputs(8068) <= layer2_outputs(2954);
    outputs(8069) <= not(layer2_outputs(8998));
    outputs(8070) <= not(layer2_outputs(524));
    outputs(8071) <= not((layer2_outputs(9953)) and (layer2_outputs(2502)));
    outputs(8072) <= (layer2_outputs(3944)) and (layer2_outputs(10163));
    outputs(8073) <= (layer2_outputs(12008)) xor (layer2_outputs(8555));
    outputs(8074) <= layer2_outputs(1708);
    outputs(8075) <= not(layer2_outputs(7788));
    outputs(8076) <= (layer2_outputs(4212)) and not (layer2_outputs(6007));
    outputs(8077) <= not(layer2_outputs(5701));
    outputs(8078) <= layer2_outputs(4004);
    outputs(8079) <= not((layer2_outputs(770)) or (layer2_outputs(7259)));
    outputs(8080) <= (layer2_outputs(8636)) xor (layer2_outputs(7286));
    outputs(8081) <= not(layer2_outputs(1949));
    outputs(8082) <= not(layer2_outputs(9557));
    outputs(8083) <= not(layer2_outputs(4591));
    outputs(8084) <= layer2_outputs(490);
    outputs(8085) <= not((layer2_outputs(4154)) or (layer2_outputs(3264)));
    outputs(8086) <= layer2_outputs(10958);
    outputs(8087) <= layer2_outputs(7470);
    outputs(8088) <= not(layer2_outputs(9066));
    outputs(8089) <= layer2_outputs(5533);
    outputs(8090) <= (layer2_outputs(6655)) xor (layer2_outputs(11359));
    outputs(8091) <= not(layer2_outputs(9139));
    outputs(8092) <= (layer2_outputs(4162)) and not (layer2_outputs(6754));
    outputs(8093) <= (layer2_outputs(2770)) and (layer2_outputs(3262));
    outputs(8094) <= not(layer2_outputs(5822));
    outputs(8095) <= layer2_outputs(8903);
    outputs(8096) <= (layer2_outputs(11220)) and not (layer2_outputs(7455));
    outputs(8097) <= layer2_outputs(9961);
    outputs(8098) <= not((layer2_outputs(8994)) xor (layer2_outputs(9220)));
    outputs(8099) <= layer2_outputs(2599);
    outputs(8100) <= not(layer2_outputs(11462));
    outputs(8101) <= layer2_outputs(9240);
    outputs(8102) <= layer2_outputs(1300);
    outputs(8103) <= layer2_outputs(6048);
    outputs(8104) <= not((layer2_outputs(7518)) xor (layer2_outputs(11976)));
    outputs(8105) <= layer2_outputs(9158);
    outputs(8106) <= layer2_outputs(6469);
    outputs(8107) <= not(layer2_outputs(12577));
    outputs(8108) <= not((layer2_outputs(7604)) xor (layer2_outputs(2731)));
    outputs(8109) <= (layer2_outputs(12077)) xor (layer2_outputs(6707));
    outputs(8110) <= layer2_outputs(779);
    outputs(8111) <= (layer2_outputs(2862)) and (layer2_outputs(2436));
    outputs(8112) <= layer2_outputs(11445);
    outputs(8113) <= not(layer2_outputs(7761));
    outputs(8114) <= (layer2_outputs(7353)) and (layer2_outputs(7989));
    outputs(8115) <= not((layer2_outputs(1353)) xor (layer2_outputs(8320)));
    outputs(8116) <= layer2_outputs(11778);
    outputs(8117) <= layer2_outputs(2892);
    outputs(8118) <= layer2_outputs(2577);
    outputs(8119) <= layer2_outputs(8183);
    outputs(8120) <= not(layer2_outputs(2444)) or (layer2_outputs(2281));
    outputs(8121) <= not(layer2_outputs(12289));
    outputs(8122) <= not((layer2_outputs(4199)) xor (layer2_outputs(12047)));
    outputs(8123) <= not(layer2_outputs(5229));
    outputs(8124) <= (layer2_outputs(6213)) xor (layer2_outputs(7476));
    outputs(8125) <= (layer2_outputs(7302)) and not (layer2_outputs(10723));
    outputs(8126) <= not(layer2_outputs(1081));
    outputs(8127) <= not((layer2_outputs(2967)) xor (layer2_outputs(5314)));
    outputs(8128) <= not(layer2_outputs(9875));
    outputs(8129) <= not(layer2_outputs(2632));
    outputs(8130) <= layer2_outputs(12694);
    outputs(8131) <= layer2_outputs(6144);
    outputs(8132) <= (layer2_outputs(10619)) and not (layer2_outputs(10778));
    outputs(8133) <= (layer2_outputs(8147)) and (layer2_outputs(8691));
    outputs(8134) <= (layer2_outputs(629)) and not (layer2_outputs(4549));
    outputs(8135) <= not((layer2_outputs(3314)) or (layer2_outputs(111)));
    outputs(8136) <= not(layer2_outputs(1406));
    outputs(8137) <= not(layer2_outputs(10567));
    outputs(8138) <= not(layer2_outputs(5087));
    outputs(8139) <= not(layer2_outputs(7972));
    outputs(8140) <= not(layer2_outputs(8293));
    outputs(8141) <= layer2_outputs(4832);
    outputs(8142) <= not((layer2_outputs(6388)) xor (layer2_outputs(1271)));
    outputs(8143) <= (layer2_outputs(9723)) and not (layer2_outputs(11341));
    outputs(8144) <= not(layer2_outputs(3599));
    outputs(8145) <= (layer2_outputs(1061)) and not (layer2_outputs(12383));
    outputs(8146) <= layer2_outputs(4569);
    outputs(8147) <= not(layer2_outputs(4049));
    outputs(8148) <= not(layer2_outputs(10516));
    outputs(8149) <= layer2_outputs(3488);
    outputs(8150) <= layer2_outputs(8948);
    outputs(8151) <= not(layer2_outputs(3269));
    outputs(8152) <= layer2_outputs(6887);
    outputs(8153) <= not(layer2_outputs(11537));
    outputs(8154) <= (layer2_outputs(1625)) and not (layer2_outputs(5));
    outputs(8155) <= not(layer2_outputs(5484));
    outputs(8156) <= not(layer2_outputs(4545));
    outputs(8157) <= layer2_outputs(2440);
    outputs(8158) <= not((layer2_outputs(9984)) xor (layer2_outputs(1350)));
    outputs(8159) <= not(layer2_outputs(7167));
    outputs(8160) <= (layer2_outputs(10289)) or (layer2_outputs(8562));
    outputs(8161) <= not(layer2_outputs(4605));
    outputs(8162) <= not(layer2_outputs(942));
    outputs(8163) <= not(layer2_outputs(823));
    outputs(8164) <= (layer2_outputs(5912)) and not (layer2_outputs(12416));
    outputs(8165) <= not(layer2_outputs(7438));
    outputs(8166) <= not(layer2_outputs(454));
    outputs(8167) <= not((layer2_outputs(9213)) or (layer2_outputs(3494)));
    outputs(8168) <= not(layer2_outputs(7810));
    outputs(8169) <= not(layer2_outputs(10555)) or (layer2_outputs(3288));
    outputs(8170) <= not(layer2_outputs(4149));
    outputs(8171) <= layer2_outputs(5529);
    outputs(8172) <= not((layer2_outputs(2519)) and (layer2_outputs(12748)));
    outputs(8173) <= layer2_outputs(9474);
    outputs(8174) <= layer2_outputs(8157);
    outputs(8175) <= not(layer2_outputs(10673));
    outputs(8176) <= (layer2_outputs(3485)) and not (layer2_outputs(2366));
    outputs(8177) <= not(layer2_outputs(212));
    outputs(8178) <= layer2_outputs(4748);
    outputs(8179) <= (layer2_outputs(9306)) xor (layer2_outputs(10399));
    outputs(8180) <= not(layer2_outputs(6230));
    outputs(8181) <= (layer2_outputs(3779)) xor (layer2_outputs(12431));
    outputs(8182) <= not(layer2_outputs(12192));
    outputs(8183) <= not(layer2_outputs(6885)) or (layer2_outputs(12375));
    outputs(8184) <= not((layer2_outputs(1415)) or (layer2_outputs(2209)));
    outputs(8185) <= not(layer2_outputs(4766));
    outputs(8186) <= layer2_outputs(3635);
    outputs(8187) <= layer2_outputs(7080);
    outputs(8188) <= (layer2_outputs(1852)) and not (layer2_outputs(11730));
    outputs(8189) <= not((layer2_outputs(1197)) xor (layer2_outputs(7785)));
    outputs(8190) <= not(layer2_outputs(1663));
    outputs(8191) <= layer2_outputs(1067);
    outputs(8192) <= not(layer2_outputs(511));
    outputs(8193) <= (layer2_outputs(6923)) and (layer2_outputs(7058));
    outputs(8194) <= layer2_outputs(1622);
    outputs(8195) <= (layer2_outputs(12570)) xor (layer2_outputs(10538));
    outputs(8196) <= not(layer2_outputs(8707));
    outputs(8197) <= layer2_outputs(2645);
    outputs(8198) <= not((layer2_outputs(3803)) xor (layer2_outputs(11008)));
    outputs(8199) <= not(layer2_outputs(605));
    outputs(8200) <= layer2_outputs(8134);
    outputs(8201) <= not(layer2_outputs(4419));
    outputs(8202) <= (layer2_outputs(2332)) xor (layer2_outputs(11240));
    outputs(8203) <= not(layer2_outputs(6222));
    outputs(8204) <= not((layer2_outputs(3629)) xor (layer2_outputs(2037)));
    outputs(8205) <= (layer2_outputs(7104)) and not (layer2_outputs(10723));
    outputs(8206) <= not(layer2_outputs(5691));
    outputs(8207) <= not((layer2_outputs(978)) xor (layer2_outputs(1230)));
    outputs(8208) <= layer2_outputs(10330);
    outputs(8209) <= layer2_outputs(9830);
    outputs(8210) <= not((layer2_outputs(4541)) xor (layer2_outputs(1307)));
    outputs(8211) <= not((layer2_outputs(12110)) xor (layer2_outputs(887)));
    outputs(8212) <= (layer2_outputs(7383)) and not (layer2_outputs(8430));
    outputs(8213) <= layer2_outputs(11740);
    outputs(8214) <= (layer2_outputs(12308)) or (layer2_outputs(1829));
    outputs(8215) <= (layer2_outputs(1938)) xor (layer2_outputs(5013));
    outputs(8216) <= layer2_outputs(1472);
    outputs(8217) <= not(layer2_outputs(5736));
    outputs(8218) <= (layer2_outputs(3864)) xor (layer2_outputs(5702));
    outputs(8219) <= layer2_outputs(4815);
    outputs(8220) <= not(layer2_outputs(7448));
    outputs(8221) <= not((layer2_outputs(10699)) xor (layer2_outputs(2810)));
    outputs(8222) <= not(layer2_outputs(2657));
    outputs(8223) <= not(layer2_outputs(10999));
    outputs(8224) <= layer2_outputs(11697);
    outputs(8225) <= layer2_outputs(5660);
    outputs(8226) <= not(layer2_outputs(1182));
    outputs(8227) <= not(layer2_outputs(8991));
    outputs(8228) <= not((layer2_outputs(8737)) xor (layer2_outputs(768)));
    outputs(8229) <= not(layer2_outputs(5244));
    outputs(8230) <= (layer2_outputs(4976)) and (layer2_outputs(6016));
    outputs(8231) <= layer2_outputs(3172);
    outputs(8232) <= not(layer2_outputs(10518));
    outputs(8233) <= layer2_outputs(6262);
    outputs(8234) <= layer2_outputs(9021);
    outputs(8235) <= not((layer2_outputs(6503)) and (layer2_outputs(8154)));
    outputs(8236) <= layer2_outputs(2044);
    outputs(8237) <= (layer2_outputs(5213)) or (layer2_outputs(12182));
    outputs(8238) <= layer2_outputs(6189);
    outputs(8239) <= not(layer2_outputs(10349));
    outputs(8240) <= not(layer2_outputs(4796));
    outputs(8241) <= not(layer2_outputs(3619));
    outputs(8242) <= not(layer2_outputs(1778));
    outputs(8243) <= layer2_outputs(9208);
    outputs(8244) <= (layer2_outputs(2531)) and (layer2_outputs(3645));
    outputs(8245) <= layer2_outputs(9175);
    outputs(8246) <= not((layer2_outputs(880)) xor (layer2_outputs(1693)));
    outputs(8247) <= not(layer2_outputs(7769));
    outputs(8248) <= not(layer2_outputs(4035));
    outputs(8249) <= (layer2_outputs(7471)) and (layer2_outputs(10373));
    outputs(8250) <= not(layer2_outputs(2794));
    outputs(8251) <= not(layer2_outputs(12607));
    outputs(8252) <= not(layer2_outputs(2030));
    outputs(8253) <= not(layer2_outputs(4123));
    outputs(8254) <= not(layer2_outputs(4542));
    outputs(8255) <= not(layer2_outputs(10765));
    outputs(8256) <= layer2_outputs(2580);
    outputs(8257) <= (layer2_outputs(12010)) or (layer2_outputs(1084));
    outputs(8258) <= layer2_outputs(1988);
    outputs(8259) <= not((layer2_outputs(12323)) and (layer2_outputs(8777)));
    outputs(8260) <= not((layer2_outputs(1705)) xor (layer2_outputs(5120)));
    outputs(8261) <= not(layer2_outputs(7315));
    outputs(8262) <= layer2_outputs(1449);
    outputs(8263) <= not(layer2_outputs(2906));
    outputs(8264) <= layer2_outputs(10266);
    outputs(8265) <= not(layer2_outputs(12088));
    outputs(8266) <= layer2_outputs(4576);
    outputs(8267) <= not(layer2_outputs(5560));
    outputs(8268) <= layer2_outputs(3882);
    outputs(8269) <= not((layer2_outputs(2446)) xor (layer2_outputs(12362)));
    outputs(8270) <= (layer2_outputs(6524)) and (layer2_outputs(6573));
    outputs(8271) <= not(layer2_outputs(9458));
    outputs(8272) <= not(layer2_outputs(2521));
    outputs(8273) <= not((layer2_outputs(5562)) or (layer2_outputs(9009)));
    outputs(8274) <= (layer2_outputs(6155)) xor (layer2_outputs(1193));
    outputs(8275) <= not(layer2_outputs(6353));
    outputs(8276) <= not((layer2_outputs(11000)) xor (layer2_outputs(9180)));
    outputs(8277) <= not(layer2_outputs(7821));
    outputs(8278) <= layer2_outputs(589);
    outputs(8279) <= (layer2_outputs(4127)) and not (layer2_outputs(3714));
    outputs(8280) <= not(layer2_outputs(5254));
    outputs(8281) <= (layer2_outputs(10293)) xor (layer2_outputs(2457));
    outputs(8282) <= layer2_outputs(2962);
    outputs(8283) <= layer2_outputs(4681);
    outputs(8284) <= (layer2_outputs(651)) and not (layer2_outputs(2660));
    outputs(8285) <= not(layer2_outputs(6860));
    outputs(8286) <= (layer2_outputs(476)) xor (layer2_outputs(10886));
    outputs(8287) <= layer2_outputs(6330);
    outputs(8288) <= layer2_outputs(11931);
    outputs(8289) <= layer2_outputs(11578);
    outputs(8290) <= not(layer2_outputs(5910));
    outputs(8291) <= not(layer2_outputs(6883));
    outputs(8292) <= not(layer2_outputs(1060));
    outputs(8293) <= not((layer2_outputs(2604)) xor (layer2_outputs(3885)));
    outputs(8294) <= (layer2_outputs(6359)) and not (layer2_outputs(4820));
    outputs(8295) <= (layer2_outputs(1064)) xor (layer2_outputs(10554));
    outputs(8296) <= not(layer2_outputs(8478));
    outputs(8297) <= layer2_outputs(351);
    outputs(8298) <= (layer2_outputs(7135)) and not (layer2_outputs(6494));
    outputs(8299) <= not(layer2_outputs(1238));
    outputs(8300) <= layer2_outputs(8283);
    outputs(8301) <= (layer2_outputs(4357)) and not (layer2_outputs(5316));
    outputs(8302) <= (layer2_outputs(2876)) xor (layer2_outputs(3931));
    outputs(8303) <= not(layer2_outputs(7716)) or (layer2_outputs(11038));
    outputs(8304) <= not((layer2_outputs(2289)) xor (layer2_outputs(8743)));
    outputs(8305) <= layer2_outputs(7095);
    outputs(8306) <= not(layer2_outputs(5276));
    outputs(8307) <= not((layer2_outputs(3031)) xor (layer2_outputs(8316)));
    outputs(8308) <= layer2_outputs(11516);
    outputs(8309) <= not(layer2_outputs(2148));
    outputs(8310) <= not(layer2_outputs(5562));
    outputs(8311) <= not(layer2_outputs(9910));
    outputs(8312) <= layer2_outputs(3839);
    outputs(8313) <= (layer2_outputs(782)) and (layer2_outputs(9739));
    outputs(8314) <= not(layer2_outputs(4647));
    outputs(8315) <= not(layer2_outputs(7569));
    outputs(8316) <= not((layer2_outputs(10674)) xor (layer2_outputs(12640)));
    outputs(8317) <= not(layer2_outputs(7057));
    outputs(8318) <= (layer2_outputs(10086)) xor (layer2_outputs(77));
    outputs(8319) <= not(layer2_outputs(9344));
    outputs(8320) <= not(layer2_outputs(5917));
    outputs(8321) <= layer2_outputs(9675);
    outputs(8322) <= (layer2_outputs(5886)) and not (layer2_outputs(4793));
    outputs(8323) <= layer2_outputs(5606);
    outputs(8324) <= not(layer2_outputs(10780));
    outputs(8325) <= layer2_outputs(6818);
    outputs(8326) <= (layer2_outputs(1)) xor (layer2_outputs(6829));
    outputs(8327) <= not(layer2_outputs(8023));
    outputs(8328) <= not((layer2_outputs(12341)) xor (layer2_outputs(1039)));
    outputs(8329) <= (layer2_outputs(5207)) and not (layer2_outputs(3557));
    outputs(8330) <= not(layer2_outputs(3085));
    outputs(8331) <= layer2_outputs(6047);
    outputs(8332) <= not((layer2_outputs(194)) xor (layer2_outputs(6147)));
    outputs(8333) <= (layer2_outputs(1902)) xor (layer2_outputs(5020));
    outputs(8334) <= layer2_outputs(5679);
    outputs(8335) <= not(layer2_outputs(5080));
    outputs(8336) <= not(layer2_outputs(553));
    outputs(8337) <= not(layer2_outputs(3415));
    outputs(8338) <= not(layer2_outputs(2450)) or (layer2_outputs(10547));
    outputs(8339) <= layer2_outputs(9812);
    outputs(8340) <= not(layer2_outputs(10479));
    outputs(8341) <= not((layer2_outputs(12394)) or (layer2_outputs(8015)));
    outputs(8342) <= layer2_outputs(9790);
    outputs(8343) <= layer2_outputs(7642);
    outputs(8344) <= not((layer2_outputs(12175)) or (layer2_outputs(172)));
    outputs(8345) <= not(layer2_outputs(8652));
    outputs(8346) <= (layer2_outputs(10693)) and not (layer2_outputs(7800));
    outputs(8347) <= not(layer2_outputs(8208));
    outputs(8348) <= not((layer2_outputs(6656)) or (layer2_outputs(7559)));
    outputs(8349) <= (layer2_outputs(8180)) and not (layer2_outputs(3145));
    outputs(8350) <= not(layer2_outputs(2385));
    outputs(8351) <= (layer2_outputs(6194)) xor (layer2_outputs(3142));
    outputs(8352) <= not(layer2_outputs(12363)) or (layer2_outputs(10005));
    outputs(8353) <= not(layer2_outputs(411));
    outputs(8354) <= not((layer2_outputs(2490)) xor (layer2_outputs(8202)));
    outputs(8355) <= not(layer2_outputs(7121));
    outputs(8356) <= (layer2_outputs(499)) and (layer2_outputs(3258));
    outputs(8357) <= not(layer2_outputs(9670));
    outputs(8358) <= layer2_outputs(6428);
    outputs(8359) <= layer2_outputs(10738);
    outputs(8360) <= not(layer2_outputs(1109));
    outputs(8361) <= not(layer2_outputs(4128));
    outputs(8362) <= not(layer2_outputs(5172));
    outputs(8363) <= layer2_outputs(451);
    outputs(8364) <= layer2_outputs(7709);
    outputs(8365) <= not(layer2_outputs(98));
    outputs(8366) <= not(layer2_outputs(2652));
    outputs(8367) <= layer2_outputs(9894);
    outputs(8368) <= (layer2_outputs(8198)) and (layer2_outputs(2996));
    outputs(8369) <= (layer2_outputs(11683)) and not (layer2_outputs(11808));
    outputs(8370) <= layer2_outputs(7809);
    outputs(8371) <= (layer2_outputs(7407)) and not (layer2_outputs(5183));
    outputs(8372) <= (layer2_outputs(632)) xor (layer2_outputs(12237));
    outputs(8373) <= not(layer2_outputs(6185));
    outputs(8374) <= not(layer2_outputs(2738));
    outputs(8375) <= layer2_outputs(10636);
    outputs(8376) <= (layer2_outputs(7672)) and not (layer2_outputs(2551));
    outputs(8377) <= (layer2_outputs(17)) and not (layer2_outputs(5007));
    outputs(8378) <= not(layer2_outputs(10837));
    outputs(8379) <= (layer2_outputs(641)) and not (layer2_outputs(11810));
    outputs(8380) <= (layer2_outputs(1651)) and not (layer2_outputs(8276));
    outputs(8381) <= layer2_outputs(11540);
    outputs(8382) <= not(layer2_outputs(3118));
    outputs(8383) <= not(layer2_outputs(2758));
    outputs(8384) <= layer2_outputs(3862);
    outputs(8385) <= not(layer2_outputs(10167));
    outputs(8386) <= (layer2_outputs(3530)) xor (layer2_outputs(8402));
    outputs(8387) <= (layer2_outputs(11804)) and not (layer2_outputs(10850));
    outputs(8388) <= (layer2_outputs(8830)) and not (layer2_outputs(1892));
    outputs(8389) <= not((layer2_outputs(10315)) and (layer2_outputs(9018)));
    outputs(8390) <= (layer2_outputs(1225)) xor (layer2_outputs(3110));
    outputs(8391) <= layer2_outputs(1390);
    outputs(8392) <= not(layer2_outputs(7158));
    outputs(8393) <= not(layer2_outputs(8471));
    outputs(8394) <= layer2_outputs(9621);
    outputs(8395) <= (layer2_outputs(5749)) and (layer2_outputs(6215));
    outputs(8396) <= (layer2_outputs(2190)) xor (layer2_outputs(1467));
    outputs(8397) <= layer2_outputs(11289);
    outputs(8398) <= not(layer2_outputs(1116));
    outputs(8399) <= not(layer2_outputs(383));
    outputs(8400) <= not(layer2_outputs(1631));
    outputs(8401) <= not(layer2_outputs(2328));
    outputs(8402) <= not(layer2_outputs(7204)) or (layer2_outputs(3660));
    outputs(8403) <= (layer2_outputs(6354)) xor (layer2_outputs(9705));
    outputs(8404) <= (layer2_outputs(10471)) and not (layer2_outputs(5624));
    outputs(8405) <= (layer2_outputs(12028)) and not (layer2_outputs(6705));
    outputs(8406) <= not(layer2_outputs(12443));
    outputs(8407) <= (layer2_outputs(8267)) xor (layer2_outputs(12236));
    outputs(8408) <= not(layer2_outputs(10305));
    outputs(8409) <= (layer2_outputs(12279)) and (layer2_outputs(5391));
    outputs(8410) <= layer2_outputs(2401);
    outputs(8411) <= not((layer2_outputs(2638)) xor (layer2_outputs(11224)));
    outputs(8412) <= not(layer2_outputs(11553));
    outputs(8413) <= not(layer2_outputs(7860));
    outputs(8414) <= layer2_outputs(10634);
    outputs(8415) <= not((layer2_outputs(9547)) xor (layer2_outputs(532)));
    outputs(8416) <= not((layer2_outputs(5466)) xor (layer2_outputs(6718)));
    outputs(8417) <= layer2_outputs(7065);
    outputs(8418) <= not((layer2_outputs(9092)) xor (layer2_outputs(7515)));
    outputs(8419) <= not((layer2_outputs(8322)) and (layer2_outputs(8272)));
    outputs(8420) <= layer2_outputs(259);
    outputs(8421) <= not(layer2_outputs(7157));
    outputs(8422) <= (layer2_outputs(3395)) xor (layer2_outputs(734));
    outputs(8423) <= layer2_outputs(10734);
    outputs(8424) <= (layer2_outputs(337)) and not (layer2_outputs(11165));
    outputs(8425) <= not(layer2_outputs(8496)) or (layer2_outputs(1148));
    outputs(8426) <= layer2_outputs(4903);
    outputs(8427) <= not(layer2_outputs(10224)) or (layer2_outputs(1058));
    outputs(8428) <= layer2_outputs(12784);
    outputs(8429) <= not(layer2_outputs(1663)) or (layer2_outputs(6028));
    outputs(8430) <= not((layer2_outputs(6594)) xor (layer2_outputs(345)));
    outputs(8431) <= (layer2_outputs(578)) and not (layer2_outputs(11107));
    outputs(8432) <= (layer2_outputs(4858)) and (layer2_outputs(11509));
    outputs(8433) <= not(layer2_outputs(2613));
    outputs(8434) <= (layer2_outputs(8434)) and not (layer2_outputs(5926));
    outputs(8435) <= not(layer2_outputs(5056));
    outputs(8436) <= layer2_outputs(4479);
    outputs(8437) <= (layer2_outputs(4925)) or (layer2_outputs(6800));
    outputs(8438) <= (layer2_outputs(3256)) and (layer2_outputs(2541));
    outputs(8439) <= (layer2_outputs(6776)) and (layer2_outputs(3946));
    outputs(8440) <= layer2_outputs(11118);
    outputs(8441) <= (layer2_outputs(12319)) xor (layer2_outputs(6322));
    outputs(8442) <= not(layer2_outputs(12401)) or (layer2_outputs(12614));
    outputs(8443) <= not((layer2_outputs(12266)) xor (layer2_outputs(2213)));
    outputs(8444) <= not(layer2_outputs(6394));
    outputs(8445) <= layer2_outputs(10353);
    outputs(8446) <= not(layer2_outputs(9689));
    outputs(8447) <= (layer2_outputs(8664)) and (layer2_outputs(2698));
    outputs(8448) <= layer2_outputs(9889);
    outputs(8449) <= not((layer2_outputs(5038)) xor (layer2_outputs(11934)));
    outputs(8450) <= not(layer2_outputs(9323));
    outputs(8451) <= (layer2_outputs(5577)) xor (layer2_outputs(9300));
    outputs(8452) <= (layer2_outputs(6596)) and (layer2_outputs(7768));
    outputs(8453) <= layer2_outputs(7534);
    outputs(8454) <= (layer2_outputs(7522)) and not (layer2_outputs(9235));
    outputs(8455) <= not(layer2_outputs(4657));
    outputs(8456) <= not(layer2_outputs(5223)) or (layer2_outputs(1610));
    outputs(8457) <= not(layer2_outputs(6641)) or (layer2_outputs(10674));
    outputs(8458) <= (layer2_outputs(12628)) xor (layer2_outputs(7684));
    outputs(8459) <= not(layer2_outputs(776));
    outputs(8460) <= not(layer2_outputs(12719));
    outputs(8461) <= layer2_outputs(5191);
    outputs(8462) <= not((layer2_outputs(1210)) xor (layer2_outputs(11210)));
    outputs(8463) <= layer2_outputs(1080);
    outputs(8464) <= (layer2_outputs(3994)) and (layer2_outputs(9476));
    outputs(8465) <= layer2_outputs(6330);
    outputs(8466) <= not(layer2_outputs(4851));
    outputs(8467) <= not(layer2_outputs(7563));
    outputs(8468) <= (layer2_outputs(9354)) and not (layer2_outputs(10568));
    outputs(8469) <= layer2_outputs(5203);
    outputs(8470) <= layer2_outputs(2577);
    outputs(8471) <= (layer2_outputs(12515)) and not (layer2_outputs(999));
    outputs(8472) <= not(layer2_outputs(12392));
    outputs(8473) <= layer2_outputs(2670);
    outputs(8474) <= (layer2_outputs(2170)) xor (layer2_outputs(4337));
    outputs(8475) <= not(layer2_outputs(5595));
    outputs(8476) <= layer2_outputs(5967);
    outputs(8477) <= not(layer2_outputs(6015));
    outputs(8478) <= layer2_outputs(4459);
    outputs(8479) <= layer2_outputs(3192);
    outputs(8480) <= not(layer2_outputs(1335));
    outputs(8481) <= (layer2_outputs(5877)) xor (layer2_outputs(8881));
    outputs(8482) <= (layer2_outputs(6880)) xor (layer2_outputs(4509));
    outputs(8483) <= layer2_outputs(9119);
    outputs(8484) <= layer2_outputs(3535);
    outputs(8485) <= not(layer2_outputs(6456));
    outputs(8486) <= not(layer2_outputs(11246));
    outputs(8487) <= not(layer2_outputs(2407)) or (layer2_outputs(12174));
    outputs(8488) <= (layer2_outputs(609)) xor (layer2_outputs(10324));
    outputs(8489) <= layer2_outputs(2812);
    outputs(8490) <= not(layer2_outputs(6862));
    outputs(8491) <= not(layer2_outputs(770));
    outputs(8492) <= layer2_outputs(2498);
    outputs(8493) <= not((layer2_outputs(2668)) xor (layer2_outputs(10911)));
    outputs(8494) <= not((layer2_outputs(1944)) xor (layer2_outputs(10287)));
    outputs(8495) <= not((layer2_outputs(12136)) or (layer2_outputs(993)));
    outputs(8496) <= not(layer2_outputs(543));
    outputs(8497) <= (layer2_outputs(1416)) xor (layer2_outputs(4589));
    outputs(8498) <= not(layer2_outputs(4478));
    outputs(8499) <= (layer2_outputs(10257)) xor (layer2_outputs(9438));
    outputs(8500) <= (layer2_outputs(5466)) and (layer2_outputs(4116));
    outputs(8501) <= not(layer2_outputs(9436));
    outputs(8502) <= (layer2_outputs(1630)) or (layer2_outputs(5602));
    outputs(8503) <= not(layer2_outputs(2159));
    outputs(8504) <= (layer2_outputs(69)) and not (layer2_outputs(10131));
    outputs(8505) <= not(layer2_outputs(11403));
    outputs(8506) <= (layer2_outputs(683)) and (layer2_outputs(155));
    outputs(8507) <= not((layer2_outputs(6598)) xor (layer2_outputs(7259)));
    outputs(8508) <= not((layer2_outputs(5511)) xor (layer2_outputs(1650)));
    outputs(8509) <= not(layer2_outputs(11535));
    outputs(8510) <= layer2_outputs(2560);
    outputs(8511) <= (layer2_outputs(5833)) xor (layer2_outputs(3652));
    outputs(8512) <= not(layer2_outputs(3254));
    outputs(8513) <= layer2_outputs(8677);
    outputs(8514) <= not((layer2_outputs(719)) xor (layer2_outputs(1305)));
    outputs(8515) <= layer2_outputs(3561);
    outputs(8516) <= layer2_outputs(7285);
    outputs(8517) <= layer2_outputs(3839);
    outputs(8518) <= not((layer2_outputs(5665)) xor (layer2_outputs(3388)));
    outputs(8519) <= (layer2_outputs(3867)) xor (layer2_outputs(11726));
    outputs(8520) <= not((layer2_outputs(6674)) xor (layer2_outputs(11775)));
    outputs(8521) <= layer2_outputs(10928);
    outputs(8522) <= (layer2_outputs(6087)) and not (layer2_outputs(9971));
    outputs(8523) <= not(layer2_outputs(7795));
    outputs(8524) <= not(layer2_outputs(2488));
    outputs(8525) <= not(layer2_outputs(7368));
    outputs(8526) <= (layer2_outputs(2327)) xor (layer2_outputs(3284));
    outputs(8527) <= layer2_outputs(11427);
    outputs(8528) <= layer2_outputs(11931);
    outputs(8529) <= layer2_outputs(5094);
    outputs(8530) <= (layer2_outputs(12435)) xor (layer2_outputs(6324));
    outputs(8531) <= not(layer2_outputs(9350)) or (layer2_outputs(11333));
    outputs(8532) <= layer2_outputs(4705);
    outputs(8533) <= not(layer2_outputs(12693));
    outputs(8534) <= (layer2_outputs(9697)) xor (layer2_outputs(8904));
    outputs(8535) <= layer2_outputs(1689);
    outputs(8536) <= not(layer2_outputs(6703)) or (layer2_outputs(7395));
    outputs(8537) <= layer2_outputs(3308);
    outputs(8538) <= layer2_outputs(853);
    outputs(8539) <= layer2_outputs(4705);
    outputs(8540) <= (layer2_outputs(10501)) and (layer2_outputs(7875));
    outputs(8541) <= not((layer2_outputs(12615)) xor (layer2_outputs(8630)));
    outputs(8542) <= (layer2_outputs(867)) and (layer2_outputs(8934));
    outputs(8543) <= layer2_outputs(9091);
    outputs(8544) <= not(layer2_outputs(10189));
    outputs(8545) <= layer2_outputs(7196);
    outputs(8546) <= not((layer2_outputs(11161)) or (layer2_outputs(10391)));
    outputs(8547) <= not(layer2_outputs(1152));
    outputs(8548) <= (layer2_outputs(12214)) and not (layer2_outputs(9975));
    outputs(8549) <= not((layer2_outputs(929)) xor (layer2_outputs(6784)));
    outputs(8550) <= layer2_outputs(8843);
    outputs(8551) <= not(layer2_outputs(10659));
    outputs(8552) <= layer2_outputs(427);
    outputs(8553) <= not(layer2_outputs(10623));
    outputs(8554) <= layer2_outputs(7078);
    outputs(8555) <= not(layer2_outputs(4434));
    outputs(8556) <= (layer2_outputs(3757)) xor (layer2_outputs(7955));
    outputs(8557) <= not(layer2_outputs(3609));
    outputs(8558) <= (layer2_outputs(39)) and not (layer2_outputs(3450));
    outputs(8559) <= (layer2_outputs(5070)) and (layer2_outputs(11301));
    outputs(8560) <= not((layer2_outputs(10592)) xor (layer2_outputs(2589)));
    outputs(8561) <= not((layer2_outputs(1215)) xor (layer2_outputs(6888)));
    outputs(8562) <= layer2_outputs(2212);
    outputs(8563) <= not(layer2_outputs(11260));
    outputs(8564) <= not(layer2_outputs(7288));
    outputs(8565) <= (layer2_outputs(6024)) and (layer2_outputs(12739));
    outputs(8566) <= (layer2_outputs(11479)) xor (layer2_outputs(10462));
    outputs(8567) <= layer2_outputs(3231);
    outputs(8568) <= layer2_outputs(11274);
    outputs(8569) <= not(layer2_outputs(5459));
    outputs(8570) <= not((layer2_outputs(12510)) or (layer2_outputs(5914)));
    outputs(8571) <= layer2_outputs(764);
    outputs(8572) <= not((layer2_outputs(2614)) and (layer2_outputs(8387)));
    outputs(8573) <= not(layer2_outputs(7553)) or (layer2_outputs(10473));
    outputs(8574) <= (layer2_outputs(1566)) and not (layer2_outputs(6475));
    outputs(8575) <= not(layer2_outputs(7235)) or (layer2_outputs(5905));
    outputs(8576) <= not(layer2_outputs(8558));
    outputs(8577) <= (layer2_outputs(5803)) xor (layer2_outputs(687));
    outputs(8578) <= not(layer2_outputs(168)) or (layer2_outputs(34));
    outputs(8579) <= not(layer2_outputs(6840));
    outputs(8580) <= not(layer2_outputs(10552));
    outputs(8581) <= (layer2_outputs(9)) and (layer2_outputs(5979));
    outputs(8582) <= (layer2_outputs(12142)) xor (layer2_outputs(1481));
    outputs(8583) <= (layer2_outputs(1939)) or (layer2_outputs(9597));
    outputs(8584) <= (layer2_outputs(8604)) and not (layer2_outputs(1543));
    outputs(8585) <= (layer2_outputs(9068)) and (layer2_outputs(12117));
    outputs(8586) <= layer2_outputs(11583);
    outputs(8587) <= not(layer2_outputs(7916));
    outputs(8588) <= (layer2_outputs(1187)) xor (layer2_outputs(11687));
    outputs(8589) <= not(layer2_outputs(1191));
    outputs(8590) <= not(layer2_outputs(3801));
    outputs(8591) <= not(layer2_outputs(10068));
    outputs(8592) <= layer2_outputs(11118);
    outputs(8593) <= not(layer2_outputs(575));
    outputs(8594) <= layer2_outputs(3400);
    outputs(8595) <= layer2_outputs(5449);
    outputs(8596) <= (layer2_outputs(4280)) and (layer2_outputs(3459));
    outputs(8597) <= layer2_outputs(2933);
    outputs(8598) <= not(layer2_outputs(5482));
    outputs(8599) <= layer2_outputs(5958);
    outputs(8600) <= layer2_outputs(11302);
    outputs(8601) <= layer2_outputs(9602);
    outputs(8602) <= not(layer2_outputs(7998));
    outputs(8603) <= not((layer2_outputs(8928)) xor (layer2_outputs(10625)));
    outputs(8604) <= layer2_outputs(12364);
    outputs(8605) <= (layer2_outputs(9682)) and not (layer2_outputs(9053));
    outputs(8606) <= not(layer2_outputs(1554));
    outputs(8607) <= not((layer2_outputs(2291)) xor (layer2_outputs(8824)));
    outputs(8608) <= layer2_outputs(6025);
    outputs(8609) <= (layer2_outputs(11092)) xor (layer2_outputs(12633));
    outputs(8610) <= not((layer2_outputs(9942)) and (layer2_outputs(1838)));
    outputs(8611) <= layer2_outputs(187);
    outputs(8612) <= layer2_outputs(9160);
    outputs(8613) <= layer2_outputs(5830);
    outputs(8614) <= not((layer2_outputs(4003)) or (layer2_outputs(9610)));
    outputs(8615) <= not(layer2_outputs(3970));
    outputs(8616) <= layer2_outputs(6374);
    outputs(8617) <= not(layer2_outputs(3542));
    outputs(8618) <= not((layer2_outputs(4449)) xor (layer2_outputs(1275)));
    outputs(8619) <= layer2_outputs(9419);
    outputs(8620) <= (layer2_outputs(6106)) and not (layer2_outputs(8146));
    outputs(8621) <= not((layer2_outputs(4695)) xor (layer2_outputs(10335)));
    outputs(8622) <= not(layer2_outputs(12647));
    outputs(8623) <= not((layer2_outputs(6617)) or (layer2_outputs(6210)));
    outputs(8624) <= (layer2_outputs(1113)) xor (layer2_outputs(5975));
    outputs(8625) <= not(layer2_outputs(1324));
    outputs(8626) <= not(layer2_outputs(12619)) or (layer2_outputs(276));
    outputs(8627) <= not(layer2_outputs(9232));
    outputs(8628) <= layer2_outputs(11376);
    outputs(8629) <= not(layer2_outputs(2773));
    outputs(8630) <= not(layer2_outputs(6439));
    outputs(8631) <= layer2_outputs(3191);
    outputs(8632) <= not((layer2_outputs(4803)) xor (layer2_outputs(4023)));
    outputs(8633) <= layer2_outputs(12061);
    outputs(8634) <= (layer2_outputs(6200)) and not (layer2_outputs(8106));
    outputs(8635) <= not(layer2_outputs(4351));
    outputs(8636) <= not(layer2_outputs(3149)) or (layer2_outputs(10270));
    outputs(8637) <= not((layer2_outputs(11796)) or (layer2_outputs(459)));
    outputs(8638) <= layer2_outputs(2181);
    outputs(8639) <= layer2_outputs(9729);
    outputs(8640) <= not(layer2_outputs(7748));
    outputs(8641) <= layer2_outputs(5650);
    outputs(8642) <= not(layer2_outputs(10570));
    outputs(8643) <= not((layer2_outputs(10171)) and (layer2_outputs(2563)));
    outputs(8644) <= not((layer2_outputs(2399)) and (layer2_outputs(2538)));
    outputs(8645) <= not((layer2_outputs(4387)) xor (layer2_outputs(12498)));
    outputs(8646) <= layer2_outputs(4130);
    outputs(8647) <= not(layer2_outputs(2679));
    outputs(8648) <= (layer2_outputs(2069)) xor (layer2_outputs(5718));
    outputs(8649) <= layer2_outputs(2483);
    outputs(8650) <= not(layer2_outputs(3139));
    outputs(8651) <= not(layer2_outputs(8584));
    outputs(8652) <= layer2_outputs(3552);
    outputs(8653) <= layer2_outputs(10015);
    outputs(8654) <= not(layer2_outputs(2471));
    outputs(8655) <= not(layer2_outputs(8833));
    outputs(8656) <= not(layer2_outputs(5106));
    outputs(8657) <= not(layer2_outputs(11643)) or (layer2_outputs(2746));
    outputs(8658) <= layer2_outputs(3601);
    outputs(8659) <= not((layer2_outputs(12348)) xor (layer2_outputs(99)));
    outputs(8660) <= (layer2_outputs(11295)) xor (layer2_outputs(10455));
    outputs(8661) <= not(layer2_outputs(6684));
    outputs(8662) <= not(layer2_outputs(3438));
    outputs(8663) <= layer2_outputs(5235);
    outputs(8664) <= not(layer2_outputs(1295));
    outputs(8665) <= not(layer2_outputs(12589));
    outputs(8666) <= (layer2_outputs(10331)) and not (layer2_outputs(9232));
    outputs(8667) <= not(layer2_outputs(4849));
    outputs(8668) <= layer2_outputs(3499);
    outputs(8669) <= not(layer2_outputs(5694)) or (layer2_outputs(11753));
    outputs(8670) <= (layer2_outputs(12786)) or (layer2_outputs(12387));
    outputs(8671) <= layer2_outputs(9771);
    outputs(8672) <= layer2_outputs(6052);
    outputs(8673) <= not((layer2_outputs(10532)) xor (layer2_outputs(8514)));
    outputs(8674) <= layer2_outputs(8250);
    outputs(8675) <= not(layer2_outputs(8523));
    outputs(8676) <= not(layer2_outputs(8816));
    outputs(8677) <= not((layer2_outputs(3778)) xor (layer2_outputs(10758)));
    outputs(8678) <= (layer2_outputs(1147)) xor (layer2_outputs(8110));
    outputs(8679) <= (layer2_outputs(10735)) and not (layer2_outputs(1588));
    outputs(8680) <= not(layer2_outputs(2590));
    outputs(8681) <= layer2_outputs(4815);
    outputs(8682) <= not(layer2_outputs(8437));
    outputs(8683) <= layer2_outputs(2575);
    outputs(8684) <= layer2_outputs(4971);
    outputs(8685) <= layer2_outputs(3948);
    outputs(8686) <= not((layer2_outputs(4778)) xor (layer2_outputs(1879)));
    outputs(8687) <= not(layer2_outputs(10236));
    outputs(8688) <= not(layer2_outputs(9769));
    outputs(8689) <= (layer2_outputs(12104)) xor (layer2_outputs(12073));
    outputs(8690) <= (layer2_outputs(632)) and (layer2_outputs(5354));
    outputs(8691) <= not(layer2_outputs(4301));
    outputs(8692) <= (layer2_outputs(3026)) and not (layer2_outputs(12188));
    outputs(8693) <= not((layer2_outputs(5901)) or (layer2_outputs(1122)));
    outputs(8694) <= layer2_outputs(2981);
    outputs(8695) <= layer2_outputs(9281);
    outputs(8696) <= layer2_outputs(527);
    outputs(8697) <= not(layer2_outputs(8508));
    outputs(8698) <= not((layer2_outputs(1228)) xor (layer2_outputs(7427)));
    outputs(8699) <= not(layer2_outputs(12311));
    outputs(8700) <= (layer2_outputs(12652)) and (layer2_outputs(10550));
    outputs(8701) <= layer2_outputs(10527);
    outputs(8702) <= not((layer2_outputs(9744)) or (layer2_outputs(8489)));
    outputs(8703) <= (layer2_outputs(3765)) and not (layer2_outputs(8844));
    outputs(8704) <= not(layer2_outputs(2459));
    outputs(8705) <= not(layer2_outputs(1912));
    outputs(8706) <= layer2_outputs(8064);
    outputs(8707) <= layer2_outputs(7240);
    outputs(8708) <= layer2_outputs(7798);
    outputs(8709) <= not(layer2_outputs(8398)) or (layer2_outputs(10938));
    outputs(8710) <= layer2_outputs(6653);
    outputs(8711) <= not(layer2_outputs(12455));
    outputs(8712) <= (layer2_outputs(863)) and (layer2_outputs(6696));
    outputs(8713) <= layer2_outputs(8917);
    outputs(8714) <= layer2_outputs(4974);
    outputs(8715) <= not((layer2_outputs(7636)) or (layer2_outputs(6238)));
    outputs(8716) <= (layer2_outputs(1377)) xor (layer2_outputs(3024));
    outputs(8717) <= (layer2_outputs(2031)) and not (layer2_outputs(4398));
    outputs(8718) <= layer2_outputs(6994);
    outputs(8719) <= not((layer2_outputs(1246)) xor (layer2_outputs(1969)));
    outputs(8720) <= layer2_outputs(3097);
    outputs(8721) <= layer2_outputs(12173);
    outputs(8722) <= not(layer2_outputs(841));
    outputs(8723) <= layer2_outputs(10741);
    outputs(8724) <= not(layer2_outputs(7825));
    outputs(8725) <= not(layer2_outputs(1821));
    outputs(8726) <= (layer2_outputs(8540)) xor (layer2_outputs(3193));
    outputs(8727) <= not((layer2_outputs(464)) xor (layer2_outputs(12191)));
    outputs(8728) <= (layer2_outputs(8914)) and (layer2_outputs(2435));
    outputs(8729) <= layer2_outputs(12787);
    outputs(8730) <= not(layer2_outputs(6924));
    outputs(8731) <= layer2_outputs(4159);
    outputs(8732) <= layer2_outputs(5518);
    outputs(8733) <= layer2_outputs(4685);
    outputs(8734) <= not(layer2_outputs(2230));
    outputs(8735) <= not(layer2_outputs(2249));
    outputs(8736) <= not(layer2_outputs(6502));
    outputs(8737) <= layer2_outputs(5474);
    outputs(8738) <= layer2_outputs(3457);
    outputs(8739) <= (layer2_outputs(8800)) xor (layer2_outputs(1150));
    outputs(8740) <= (layer2_outputs(8395)) and not (layer2_outputs(1647));
    outputs(8741) <= (layer2_outputs(9279)) and not (layer2_outputs(6971));
    outputs(8742) <= (layer2_outputs(8092)) or (layer2_outputs(8579));
    outputs(8743) <= layer2_outputs(693);
    outputs(8744) <= not(layer2_outputs(3711));
    outputs(8745) <= layer2_outputs(6040);
    outputs(8746) <= layer2_outputs(1065);
    outputs(8747) <= layer2_outputs(10075);
    outputs(8748) <= (layer2_outputs(12058)) and (layer2_outputs(12071));
    outputs(8749) <= not(layer2_outputs(4453));
    outputs(8750) <= (layer2_outputs(11738)) or (layer2_outputs(3680));
    outputs(8751) <= not(layer2_outputs(5266));
    outputs(8752) <= not((layer2_outputs(3201)) or (layer2_outputs(7055)));
    outputs(8753) <= not((layer2_outputs(2606)) xor (layer2_outputs(6472)));
    outputs(8754) <= not((layer2_outputs(2893)) xor (layer2_outputs(7192)));
    outputs(8755) <= (layer2_outputs(1369)) and not (layer2_outputs(9623));
    outputs(8756) <= not(layer2_outputs(2808));
    outputs(8757) <= not(layer2_outputs(1503));
    outputs(8758) <= (layer2_outputs(90)) xor (layer2_outputs(11544));
    outputs(8759) <= not(layer2_outputs(239));
    outputs(8760) <= layer2_outputs(7753);
    outputs(8761) <= layer2_outputs(7522);
    outputs(8762) <= not(layer2_outputs(3923)) or (layer2_outputs(4804));
    outputs(8763) <= not((layer2_outputs(2883)) xor (layer2_outputs(9453)));
    outputs(8764) <= layer2_outputs(4952);
    outputs(8765) <= not(layer2_outputs(12217));
    outputs(8766) <= not((layer2_outputs(11832)) xor (layer2_outputs(7138)));
    outputs(8767) <= not(layer2_outputs(216));
    outputs(8768) <= not(layer2_outputs(9711));
    outputs(8769) <= (layer2_outputs(4989)) and not (layer2_outputs(9881));
    outputs(8770) <= not(layer2_outputs(8684));
    outputs(8771) <= layer2_outputs(944);
    outputs(8772) <= not((layer2_outputs(1123)) xor (layer2_outputs(12147)));
    outputs(8773) <= layer2_outputs(9997);
    outputs(8774) <= layer2_outputs(11799);
    outputs(8775) <= not((layer2_outputs(6571)) xor (layer2_outputs(6813)));
    outputs(8776) <= (layer2_outputs(520)) xor (layer2_outputs(12250));
    outputs(8777) <= layer2_outputs(4887);
    outputs(8778) <= not(layer2_outputs(5765));
    outputs(8779) <= (layer2_outputs(5290)) and not (layer2_outputs(8408));
    outputs(8780) <= (layer2_outputs(11283)) xor (layer2_outputs(9267));
    outputs(8781) <= (layer2_outputs(1596)) xor (layer2_outputs(4837));
    outputs(8782) <= not(layer2_outputs(11971));
    outputs(8783) <= not(layer2_outputs(3301));
    outputs(8784) <= not(layer2_outputs(324));
    outputs(8785) <= (layer2_outputs(3926)) xor (layer2_outputs(10433));
    outputs(8786) <= not(layer2_outputs(10836));
    outputs(8787) <= layer2_outputs(12002);
    outputs(8788) <= not((layer2_outputs(11933)) xor (layer2_outputs(12645)));
    outputs(8789) <= (layer2_outputs(7031)) xor (layer2_outputs(7140));
    outputs(8790) <= not((layer2_outputs(12195)) or (layer2_outputs(10011)));
    outputs(8791) <= layer2_outputs(7303);
    outputs(8792) <= not(layer2_outputs(6489));
    outputs(8793) <= not((layer2_outputs(1860)) xor (layer2_outputs(2191)));
    outputs(8794) <= layer2_outputs(9648);
    outputs(8795) <= (layer2_outputs(7012)) xor (layer2_outputs(9757));
    outputs(8796) <= not((layer2_outputs(2230)) xor (layer2_outputs(9787)));
    outputs(8797) <= (layer2_outputs(7827)) and not (layer2_outputs(592));
    outputs(8798) <= not(layer2_outputs(7956));
    outputs(8799) <= layer2_outputs(12505);
    outputs(8800) <= (layer2_outputs(7356)) xor (layer2_outputs(2974));
    outputs(8801) <= layer2_outputs(9124);
    outputs(8802) <= not(layer2_outputs(4904)) or (layer2_outputs(371));
    outputs(8803) <= not((layer2_outputs(9493)) xor (layer2_outputs(2194)));
    outputs(8804) <= not((layer2_outputs(12306)) xor (layer2_outputs(12384)));
    outputs(8805) <= not((layer2_outputs(12232)) xor (layer2_outputs(9147)));
    outputs(8806) <= layer2_outputs(12101);
    outputs(8807) <= layer2_outputs(5402);
    outputs(8808) <= not(layer2_outputs(383));
    outputs(8809) <= not(layer2_outputs(8334));
    outputs(8810) <= layer2_outputs(6187);
    outputs(8811) <= (layer2_outputs(10980)) and not (layer2_outputs(7591));
    outputs(8812) <= not(layer2_outputs(3556));
    outputs(8813) <= layer2_outputs(6162);
    outputs(8814) <= not(layer2_outputs(7351));
    outputs(8815) <= layer2_outputs(1792);
    outputs(8816) <= layer2_outputs(2888);
    outputs(8817) <= (layer2_outputs(2830)) and (layer2_outputs(4991));
    outputs(8818) <= not(layer2_outputs(12460));
    outputs(8819) <= (layer2_outputs(8847)) xor (layer2_outputs(6540));
    outputs(8820) <= not(layer2_outputs(5540));
    outputs(8821) <= layer2_outputs(7905);
    outputs(8822) <= (layer2_outputs(12408)) xor (layer2_outputs(10791));
    outputs(8823) <= not(layer2_outputs(3550));
    outputs(8824) <= not(layer2_outputs(11084));
    outputs(8825) <= layer2_outputs(645);
    outputs(8826) <= not(layer2_outputs(4493));
    outputs(8827) <= layer2_outputs(690);
    outputs(8828) <= layer2_outputs(1641);
    outputs(8829) <= not(layer2_outputs(7163));
    outputs(8830) <= not(layer2_outputs(678));
    outputs(8831) <= not((layer2_outputs(2424)) xor (layer2_outputs(10881)));
    outputs(8832) <= (layer2_outputs(6156)) and not (layer2_outputs(773));
    outputs(8833) <= not(layer2_outputs(6975));
    outputs(8834) <= not(layer2_outputs(9424));
    outputs(8835) <= layer2_outputs(5165);
    outputs(8836) <= not(layer2_outputs(8877));
    outputs(8837) <= layer2_outputs(3386);
    outputs(8838) <= not(layer2_outputs(2942));
    outputs(8839) <= (layer2_outputs(6874)) and (layer2_outputs(3758));
    outputs(8840) <= not((layer2_outputs(2061)) or (layer2_outputs(8966)));
    outputs(8841) <= layer2_outputs(4148);
    outputs(8842) <= layer2_outputs(11720);
    outputs(8843) <= (layer2_outputs(8613)) xor (layer2_outputs(830));
    outputs(8844) <= not(layer2_outputs(7296)) or (layer2_outputs(11657));
    outputs(8845) <= not(layer2_outputs(9141)) or (layer2_outputs(3086));
    outputs(8846) <= not((layer2_outputs(4603)) xor (layer2_outputs(8518)));
    outputs(8847) <= layer2_outputs(6712);
    outputs(8848) <= layer2_outputs(1467);
    outputs(8849) <= not((layer2_outputs(7428)) xor (layer2_outputs(2567)));
    outputs(8850) <= not(layer2_outputs(11962));
    outputs(8851) <= layer2_outputs(4883);
    outputs(8852) <= (layer2_outputs(5641)) xor (layer2_outputs(3868));
    outputs(8853) <= layer2_outputs(11317);
    outputs(8854) <= not(layer2_outputs(7253)) or (layer2_outputs(4212));
    outputs(8855) <= not(layer2_outputs(731));
    outputs(8856) <= layer2_outputs(11742);
    outputs(8857) <= (layer2_outputs(3766)) xor (layer2_outputs(4995));
    outputs(8858) <= not((layer2_outputs(11329)) xor (layer2_outputs(2736)));
    outputs(8859) <= not((layer2_outputs(6829)) or (layer2_outputs(809)));
    outputs(8860) <= (layer2_outputs(7433)) xor (layer2_outputs(7444));
    outputs(8861) <= not(layer2_outputs(12032));
    outputs(8862) <= layer2_outputs(6595);
    outputs(8863) <= layer2_outputs(2381);
    outputs(8864) <= (layer2_outputs(12617)) xor (layer2_outputs(10647));
    outputs(8865) <= not((layer2_outputs(825)) xor (layer2_outputs(2955)));
    outputs(8866) <= layer2_outputs(5612);
    outputs(8867) <= (layer2_outputs(6049)) xor (layer2_outputs(11426));
    outputs(8868) <= layer2_outputs(10296);
    outputs(8869) <= not(layer2_outputs(1455));
    outputs(8870) <= layer2_outputs(6488);
    outputs(8871) <= not(layer2_outputs(12447));
    outputs(8872) <= not(layer2_outputs(7481));
    outputs(8873) <= not((layer2_outputs(3759)) xor (layer2_outputs(2765)));
    outputs(8874) <= not((layer2_outputs(4361)) xor (layer2_outputs(5702)));
    outputs(8875) <= not(layer2_outputs(10148));
    outputs(8876) <= layer2_outputs(8373);
    outputs(8877) <= layer2_outputs(4653);
    outputs(8878) <= (layer2_outputs(3636)) and not (layer2_outputs(11246));
    outputs(8879) <= layer2_outputs(292);
    outputs(8880) <= not(layer2_outputs(546));
    outputs(8881) <= not(layer2_outputs(5999));
    outputs(8882) <= layer2_outputs(11470);
    outputs(8883) <= layer2_outputs(6040);
    outputs(8884) <= layer2_outputs(8030);
    outputs(8885) <= layer2_outputs(9185);
    outputs(8886) <= layer2_outputs(9972);
    outputs(8887) <= not((layer2_outputs(2390)) xor (layer2_outputs(8498)));
    outputs(8888) <= (layer2_outputs(8101)) and (layer2_outputs(7699));
    outputs(8889) <= (layer2_outputs(2530)) xor (layer2_outputs(3704));
    outputs(8890) <= not(layer2_outputs(7210));
    outputs(8891) <= not(layer2_outputs(11998));
    outputs(8892) <= layer2_outputs(6676);
    outputs(8893) <= not(layer2_outputs(11655));
    outputs(8894) <= layer2_outputs(7300);
    outputs(8895) <= not((layer2_outputs(12511)) or (layer2_outputs(115)));
    outputs(8896) <= (layer2_outputs(9528)) and (layer2_outputs(5851));
    outputs(8897) <= not(layer2_outputs(616));
    outputs(8898) <= not(layer2_outputs(7996));
    outputs(8899) <= not(layer2_outputs(7448));
    outputs(8900) <= (layer2_outputs(8512)) and not (layer2_outputs(6390));
    outputs(8901) <= not(layer2_outputs(3808));
    outputs(8902) <= (layer2_outputs(7415)) xor (layer2_outputs(8104));
    outputs(8903) <= (layer2_outputs(6980)) xor (layer2_outputs(5407));
    outputs(8904) <= layer2_outputs(5847);
    outputs(8905) <= (layer2_outputs(2550)) and not (layer2_outputs(3735));
    outputs(8906) <= not(layer2_outputs(6828)) or (layer2_outputs(6463));
    outputs(8907) <= not((layer2_outputs(12278)) xor (layer2_outputs(6520)));
    outputs(8908) <= (layer2_outputs(10777)) or (layer2_outputs(3594));
    outputs(8909) <= not(layer2_outputs(4460)) or (layer2_outputs(8032));
    outputs(8910) <= not(layer2_outputs(111));
    outputs(8911) <= not(layer2_outputs(12457));
    outputs(8912) <= not(layer2_outputs(10375));
    outputs(8913) <= not((layer2_outputs(2222)) or (layer2_outputs(120)));
    outputs(8914) <= layer2_outputs(9704);
    outputs(8915) <= not((layer2_outputs(5153)) xor (layer2_outputs(3929)));
    outputs(8916) <= not(layer2_outputs(3850));
    outputs(8917) <= (layer2_outputs(278)) and not (layer2_outputs(554));
    outputs(8918) <= not(layer2_outputs(6477));
    outputs(8919) <= not(layer2_outputs(12100));
    outputs(8920) <= not((layer2_outputs(10282)) xor (layer2_outputs(207)));
    outputs(8921) <= layer2_outputs(4241);
    outputs(8922) <= not(layer2_outputs(12042));
    outputs(8923) <= not(layer2_outputs(2642));
    outputs(8924) <= not(layer2_outputs(5124));
    outputs(8925) <= not(layer2_outputs(7277)) or (layer2_outputs(434));
    outputs(8926) <= (layer2_outputs(11231)) xor (layer2_outputs(7840));
    outputs(8927) <= not(layer2_outputs(11263));
    outputs(8928) <= not(layer2_outputs(3103));
    outputs(8929) <= layer2_outputs(10842);
    outputs(8930) <= not((layer2_outputs(6442)) xor (layer2_outputs(1909)));
    outputs(8931) <= not(layer2_outputs(9507));
    outputs(8932) <= not(layer2_outputs(5384));
    outputs(8933) <= not(layer2_outputs(3303));
    outputs(8934) <= not(layer2_outputs(1997));
    outputs(8935) <= not((layer2_outputs(6122)) or (layer2_outputs(1787)));
    outputs(8936) <= layer2_outputs(1957);
    outputs(8937) <= not(layer2_outputs(7456));
    outputs(8938) <= not(layer2_outputs(6403));
    outputs(8939) <= layer2_outputs(8784);
    outputs(8940) <= not(layer2_outputs(2011));
    outputs(8941) <= not(layer2_outputs(2761));
    outputs(8942) <= (layer2_outputs(6033)) xor (layer2_outputs(5738));
    outputs(8943) <= (layer2_outputs(6536)) and not (layer2_outputs(2421));
    outputs(8944) <= not((layer2_outputs(4888)) or (layer2_outputs(9487)));
    outputs(8945) <= not(layer2_outputs(8146));
    outputs(8946) <= (layer2_outputs(8764)) and not (layer2_outputs(10640));
    outputs(8947) <= not(layer2_outputs(4166));
    outputs(8948) <= (layer2_outputs(339)) and not (layer2_outputs(3279));
    outputs(8949) <= not(layer2_outputs(6500));
    outputs(8950) <= not((layer2_outputs(3526)) or (layer2_outputs(8865)));
    outputs(8951) <= layer2_outputs(6142);
    outputs(8952) <= not(layer2_outputs(10780));
    outputs(8953) <= not((layer2_outputs(8260)) xor (layer2_outputs(7467)));
    outputs(8954) <= layer2_outputs(8347);
    outputs(8955) <= not(layer2_outputs(7032));
    outputs(8956) <= (layer2_outputs(11287)) and (layer2_outputs(2982));
    outputs(8957) <= layer2_outputs(1946);
    outputs(8958) <= (layer2_outputs(10364)) or (layer2_outputs(3558));
    outputs(8959) <= not(layer2_outputs(12703));
    outputs(8960) <= (layer2_outputs(3520)) xor (layer2_outputs(3371));
    outputs(8961) <= layer2_outputs(508);
    outputs(8962) <= layer2_outputs(9060);
    outputs(8963) <= layer2_outputs(7765);
    outputs(8964) <= (layer2_outputs(11523)) xor (layer2_outputs(10825));
    outputs(8965) <= not(layer2_outputs(11486)) or (layer2_outputs(6335));
    outputs(8966) <= not(layer2_outputs(697));
    outputs(8967) <= not((layer2_outputs(1140)) xor (layer2_outputs(7358)));
    outputs(8968) <= (layer2_outputs(12757)) and not (layer2_outputs(9621));
    outputs(8969) <= (layer2_outputs(11354)) and not (layer2_outputs(11802));
    outputs(8970) <= not(layer2_outputs(1940));
    outputs(8971) <= not((layer2_outputs(7649)) xor (layer2_outputs(1538)));
    outputs(8972) <= (layer2_outputs(11684)) xor (layer2_outputs(3963));
    outputs(8973) <= (layer2_outputs(8537)) xor (layer2_outputs(10246));
    outputs(8974) <= layer2_outputs(965);
    outputs(8975) <= not((layer2_outputs(198)) and (layer2_outputs(3939)));
    outputs(8976) <= (layer2_outputs(3083)) xor (layer2_outputs(8680));
    outputs(8977) <= layer2_outputs(8888);
    outputs(8978) <= layer2_outputs(7299);
    outputs(8979) <= (layer2_outputs(11595)) and not (layer2_outputs(7984));
    outputs(8980) <= not(layer2_outputs(5869));
    outputs(8981) <= (layer2_outputs(3048)) xor (layer2_outputs(11115));
    outputs(8982) <= layer2_outputs(9118);
    outputs(8983) <= (layer2_outputs(2315)) and not (layer2_outputs(2497));
    outputs(8984) <= layer2_outputs(2198);
    outputs(8985) <= layer2_outputs(11991);
    outputs(8986) <= not(layer2_outputs(3587));
    outputs(8987) <= (layer2_outputs(8793)) and not (layer2_outputs(10157));
    outputs(8988) <= (layer2_outputs(5552)) xor (layer2_outputs(5786));
    outputs(8989) <= layer2_outputs(12020);
    outputs(8990) <= not(layer2_outputs(8339));
    outputs(8991) <= not(layer2_outputs(9498)) or (layer2_outputs(5127));
    outputs(8992) <= (layer2_outputs(474)) or (layer2_outputs(1372));
    outputs(8993) <= (layer2_outputs(3650)) xor (layer2_outputs(12218));
    outputs(8994) <= not(layer2_outputs(1716));
    outputs(8995) <= layer2_outputs(9344);
    outputs(8996) <= not(layer2_outputs(4296));
    outputs(8997) <= (layer2_outputs(6745)) and (layer2_outputs(925));
    outputs(8998) <= not((layer2_outputs(9155)) xor (layer2_outputs(2069)));
    outputs(8999) <= layer2_outputs(9442);
    outputs(9000) <= not(layer2_outputs(6253)) or (layer2_outputs(1386));
    outputs(9001) <= not((layer2_outputs(6233)) xor (layer2_outputs(9383)));
    outputs(9002) <= not(layer2_outputs(8912));
    outputs(9003) <= layer2_outputs(3399);
    outputs(9004) <= not((layer2_outputs(5762)) or (layer2_outputs(10726)));
    outputs(9005) <= layer2_outputs(10975);
    outputs(9006) <= not(layer2_outputs(801));
    outputs(9007) <= not((layer2_outputs(10218)) xor (layer2_outputs(8615)));
    outputs(9008) <= layer2_outputs(8577);
    outputs(9009) <= (layer2_outputs(6847)) xor (layer2_outputs(1562));
    outputs(9010) <= (layer2_outputs(4546)) and not (layer2_outputs(5883));
    outputs(9011) <= not(layer2_outputs(3959));
    outputs(9012) <= layer2_outputs(10882);
    outputs(9013) <= layer2_outputs(3806);
    outputs(9014) <= not((layer2_outputs(2244)) and (layer2_outputs(2933)));
    outputs(9015) <= (layer2_outputs(12013)) and not (layer2_outputs(11619));
    outputs(9016) <= layer2_outputs(9255);
    outputs(9017) <= not(layer2_outputs(1519));
    outputs(9018) <= (layer2_outputs(11202)) and not (layer2_outputs(1601));
    outputs(9019) <= not(layer2_outputs(10031));
    outputs(9020) <= (layer2_outputs(6982)) and not (layer2_outputs(4102));
    outputs(9021) <= (layer2_outputs(1313)) and not (layer2_outputs(5398));
    outputs(9022) <= not(layer2_outputs(10083));
    outputs(9023) <= layer2_outputs(3495);
    outputs(9024) <= layer2_outputs(7766);
    outputs(9025) <= not(layer2_outputs(10611));
    outputs(9026) <= not(layer2_outputs(12276));
    outputs(9027) <= not(layer2_outputs(1571));
    outputs(9028) <= not(layer2_outputs(8976));
    outputs(9029) <= not(layer2_outputs(3691));
    outputs(9030) <= not((layer2_outputs(2594)) or (layer2_outputs(9209)));
    outputs(9031) <= not(layer2_outputs(8780));
    outputs(9032) <= not((layer2_outputs(1115)) xor (layer2_outputs(2460)));
    outputs(9033) <= layer2_outputs(7797);
    outputs(9034) <= not(layer2_outputs(7245));
    outputs(9035) <= not(layer2_outputs(6093));
    outputs(9036) <= not(layer2_outputs(9796));
    outputs(9037) <= (layer2_outputs(1627)) xor (layer2_outputs(10286));
    outputs(9038) <= not(layer2_outputs(6496));
    outputs(9039) <= (layer2_outputs(9066)) or (layer2_outputs(1603));
    outputs(9040) <= not((layer2_outputs(8367)) xor (layer2_outputs(12527)));
    outputs(9041) <= not((layer2_outputs(6290)) xor (layer2_outputs(4465)));
    outputs(9042) <= layer2_outputs(2687);
    outputs(9043) <= not(layer2_outputs(3117));
    outputs(9044) <= not(layer2_outputs(12169));
    outputs(9045) <= not(layer2_outputs(9818)) or (layer2_outputs(2140));
    outputs(9046) <= (layer2_outputs(6083)) and (layer2_outputs(9106));
    outputs(9047) <= layer2_outputs(3974);
    outputs(9048) <= (layer2_outputs(5523)) xor (layer2_outputs(2884));
    outputs(9049) <= (layer2_outputs(9970)) xor (layer2_outputs(553));
    outputs(9050) <= not(layer2_outputs(6783));
    outputs(9051) <= not(layer2_outputs(11509));
    outputs(9052) <= not(layer2_outputs(4535));
    outputs(9053) <= not(layer2_outputs(9032));
    outputs(9054) <= not(layer2_outputs(2501));
    outputs(9055) <= layer2_outputs(8657);
    outputs(9056) <= (layer2_outputs(5891)) xor (layer2_outputs(6732));
    outputs(9057) <= (layer2_outputs(1223)) and not (layer2_outputs(6633));
    outputs(9058) <= not(layer2_outputs(1359));
    outputs(9059) <= not((layer2_outputs(2476)) xor (layer2_outputs(1535)));
    outputs(9060) <= not(layer2_outputs(4582));
    outputs(9061) <= not(layer2_outputs(2722));
    outputs(9062) <= not((layer2_outputs(4986)) xor (layer2_outputs(6618)));
    outputs(9063) <= not(layer2_outputs(8200));
    outputs(9064) <= not((layer2_outputs(7245)) xor (layer2_outputs(12261)));
    outputs(9065) <= (layer2_outputs(12777)) xor (layer2_outputs(5472));
    outputs(9066) <= layer2_outputs(8327);
    outputs(9067) <= not(layer2_outputs(10101));
    outputs(9068) <= (layer2_outputs(4988)) and not (layer2_outputs(10341));
    outputs(9069) <= not((layer2_outputs(7005)) xor (layer2_outputs(11340)));
    outputs(9070) <= layer2_outputs(9694);
    outputs(9071) <= layer2_outputs(1978);
    outputs(9072) <= layer2_outputs(8451);
    outputs(9073) <= not((layer2_outputs(7054)) and (layer2_outputs(209)));
    outputs(9074) <= layer2_outputs(6787);
    outputs(9075) <= (layer2_outputs(9386)) and not (layer2_outputs(5337));
    outputs(9076) <= not(layer2_outputs(6573));
    outputs(9077) <= layer2_outputs(3312);
    outputs(9078) <= not((layer2_outputs(10663)) or (layer2_outputs(3490)));
    outputs(9079) <= layer2_outputs(986);
    outputs(9080) <= not(layer2_outputs(10559)) or (layer2_outputs(8563));
    outputs(9081) <= (layer2_outputs(4040)) xor (layer2_outputs(6991));
    outputs(9082) <= (layer2_outputs(7723)) and not (layer2_outputs(5286));
    outputs(9083) <= layer2_outputs(1033);
    outputs(9084) <= not(layer2_outputs(1013));
    outputs(9085) <= not(layer2_outputs(11907));
    outputs(9086) <= not(layer2_outputs(478));
    outputs(9087) <= not(layer2_outputs(9402));
    outputs(9088) <= (layer2_outputs(9019)) xor (layer2_outputs(91));
    outputs(9089) <= not(layer2_outputs(10533));
    outputs(9090) <= layer2_outputs(2637);
    outputs(9091) <= (layer2_outputs(10372)) and not (layer2_outputs(7733));
    outputs(9092) <= not(layer2_outputs(3319));
    outputs(9093) <= layer2_outputs(10375);
    outputs(9094) <= not(layer2_outputs(12309));
    outputs(9095) <= not(layer2_outputs(12762)) or (layer2_outputs(11097));
    outputs(9096) <= not(layer2_outputs(1259));
    outputs(9097) <= layer2_outputs(9904);
    outputs(9098) <= not(layer2_outputs(1218));
    outputs(9099) <= not(layer2_outputs(11044));
    outputs(9100) <= layer2_outputs(7410);
    outputs(9101) <= not(layer2_outputs(3328));
    outputs(9102) <= not(layer2_outputs(5582));
    outputs(9103) <= not(layer2_outputs(12247));
    outputs(9104) <= not(layer2_outputs(2992));
    outputs(9105) <= layer2_outputs(2875);
    outputs(9106) <= (layer2_outputs(813)) and not (layer2_outputs(314));
    outputs(9107) <= (layer2_outputs(1748)) and not (layer2_outputs(6685));
    outputs(9108) <= not((layer2_outputs(7293)) xor (layer2_outputs(4811)));
    outputs(9109) <= layer2_outputs(6934);
    outputs(9110) <= not(layer2_outputs(10020));
    outputs(9111) <= layer2_outputs(1927);
    outputs(9112) <= (layer2_outputs(5432)) xor (layer2_outputs(8560));
    outputs(9113) <= not(layer2_outputs(262));
    outputs(9114) <= (layer2_outputs(5560)) xor (layer2_outputs(8019));
    outputs(9115) <= not((layer2_outputs(12107)) or (layer2_outputs(6983)));
    outputs(9116) <= (layer2_outputs(7309)) or (layer2_outputs(2408));
    outputs(9117) <= not(layer2_outputs(1431));
    outputs(9118) <= layer2_outputs(7797);
    outputs(9119) <= (layer2_outputs(4105)) or (layer2_outputs(3831));
    outputs(9120) <= not(layer2_outputs(10128));
    outputs(9121) <= (layer2_outputs(8765)) and (layer2_outputs(6445));
    outputs(9122) <= not((layer2_outputs(4436)) or (layer2_outputs(307)));
    outputs(9123) <= layer2_outputs(11222);
    outputs(9124) <= not(layer2_outputs(3171));
    outputs(9125) <= not((layer2_outputs(4458)) xor (layer2_outputs(11452)));
    outputs(9126) <= not((layer2_outputs(5415)) xor (layer2_outputs(7879)));
    outputs(9127) <= layer2_outputs(10442);
    outputs(9128) <= (layer2_outputs(12540)) xor (layer2_outputs(11217));
    outputs(9129) <= not((layer2_outputs(3059)) xor (layer2_outputs(5298)));
    outputs(9130) <= not(layer2_outputs(891));
    outputs(9131) <= not((layer2_outputs(4202)) xor (layer2_outputs(11454)));
    outputs(9132) <= layer2_outputs(4658);
    outputs(9133) <= layer2_outputs(6259);
    outputs(9134) <= not((layer2_outputs(7694)) xor (layer2_outputs(7995)));
    outputs(9135) <= not(layer2_outputs(2002));
    outputs(9136) <= not(layer2_outputs(7026));
    outputs(9137) <= (layer2_outputs(2667)) xor (layer2_outputs(7750));
    outputs(9138) <= not(layer2_outputs(4992));
    outputs(9139) <= not(layer2_outputs(4383));
    outputs(9140) <= not((layer2_outputs(8814)) xor (layer2_outputs(11393)));
    outputs(9141) <= not((layer2_outputs(12267)) xor (layer2_outputs(1186)));
    outputs(9142) <= not(layer2_outputs(9293));
    outputs(9143) <= layer2_outputs(6284);
    outputs(9144) <= not((layer2_outputs(8475)) xor (layer2_outputs(4557)));
    outputs(9145) <= not(layer2_outputs(5343));
    outputs(9146) <= not(layer2_outputs(5075));
    outputs(9147) <= layer2_outputs(8111);
    outputs(9148) <= layer2_outputs(4465);
    outputs(9149) <= not(layer2_outputs(5556));
    outputs(9150) <= not(layer2_outputs(12271)) or (layer2_outputs(8186));
    outputs(9151) <= layer2_outputs(5670);
    outputs(9152) <= (layer2_outputs(6781)) xor (layer2_outputs(9055));
    outputs(9153) <= not(layer2_outputs(12287));
    outputs(9154) <= not((layer2_outputs(9176)) xor (layer2_outputs(10104)));
    outputs(9155) <= not(layer2_outputs(8488));
    outputs(9156) <= layer2_outputs(12323);
    outputs(9157) <= (layer2_outputs(6235)) xor (layer2_outputs(1672));
    outputs(9158) <= not(layer2_outputs(10346));
    outputs(9159) <= not(layer2_outputs(8397));
    outputs(9160) <= not(layer2_outputs(10534));
    outputs(9161) <= not(layer2_outputs(599)) or (layer2_outputs(5575));
    outputs(9162) <= not(layer2_outputs(192));
    outputs(9163) <= (layer2_outputs(12689)) and (layer2_outputs(857));
    outputs(9164) <= not(layer2_outputs(4026)) or (layer2_outputs(10355));
    outputs(9165) <= not(layer2_outputs(5238));
    outputs(9166) <= not((layer2_outputs(5346)) xor (layer2_outputs(1099)));
    outputs(9167) <= not((layer2_outputs(3336)) xor (layer2_outputs(5023)));
    outputs(9168) <= layer2_outputs(10383);
    outputs(9169) <= layer2_outputs(11111);
    outputs(9170) <= not(layer2_outputs(2570));
    outputs(9171) <= (layer2_outputs(5517)) xor (layer2_outputs(11005));
    outputs(9172) <= not(layer2_outputs(8701));
    outputs(9173) <= (layer2_outputs(3489)) and not (layer2_outputs(9412));
    outputs(9174) <= not(layer2_outputs(908));
    outputs(9175) <= not(layer2_outputs(8794));
    outputs(9176) <= layer2_outputs(6435);
    outputs(9177) <= layer2_outputs(296);
    outputs(9178) <= not(layer2_outputs(1402));
    outputs(9179) <= (layer2_outputs(12673)) xor (layer2_outputs(10451));
    outputs(9180) <= (layer2_outputs(2859)) and (layer2_outputs(2473));
    outputs(9181) <= not(layer2_outputs(11474));
    outputs(9182) <= not(layer2_outputs(9793));
    outputs(9183) <= not(layer2_outputs(11327));
    outputs(9184) <= not((layer2_outputs(6715)) xor (layer2_outputs(4822)));
    outputs(9185) <= layer2_outputs(2847);
    outputs(9186) <= not((layer2_outputs(11624)) xor (layer2_outputs(3909)));
    outputs(9187) <= (layer2_outputs(8798)) and not (layer2_outputs(946));
    outputs(9188) <= (layer2_outputs(9044)) xor (layer2_outputs(3644));
    outputs(9189) <= layer2_outputs(3270);
    outputs(9190) <= layer2_outputs(2118);
    outputs(9191) <= (layer2_outputs(10504)) xor (layer2_outputs(11795));
    outputs(9192) <= (layer2_outputs(4358)) and not (layer2_outputs(5256));
    outputs(9193) <= layer2_outputs(1312);
    outputs(9194) <= (layer2_outputs(12480)) and not (layer2_outputs(306));
    outputs(9195) <= (layer2_outputs(7094)) and (layer2_outputs(4160));
    outputs(9196) <= not(layer2_outputs(3814));
    outputs(9197) <= not(layer2_outputs(1951));
    outputs(9198) <= layer2_outputs(1110);
    outputs(9199) <= not(layer2_outputs(8434));
    outputs(9200) <= (layer2_outputs(9943)) and not (layer2_outputs(10449));
    outputs(9201) <= (layer2_outputs(1335)) and (layer2_outputs(6947));
    outputs(9202) <= not((layer2_outputs(8319)) xor (layer2_outputs(7969)));
    outputs(9203) <= layer2_outputs(3375);
    outputs(9204) <= (layer2_outputs(3218)) and not (layer2_outputs(7988));
    outputs(9205) <= layer2_outputs(11269);
    outputs(9206) <= not(layer2_outputs(5022));
    outputs(9207) <= (layer2_outputs(8789)) and not (layer2_outputs(8540));
    outputs(9208) <= layer2_outputs(12624);
    outputs(9209) <= not((layer2_outputs(11626)) xor (layer2_outputs(504)));
    outputs(9210) <= not(layer2_outputs(4069));
    outputs(9211) <= not(layer2_outputs(3953));
    outputs(9212) <= not((layer2_outputs(1513)) or (layer2_outputs(9423)));
    outputs(9213) <= layer2_outputs(230);
    outputs(9214) <= layer2_outputs(1978);
    outputs(9215) <= not(layer2_outputs(2071));
    outputs(9216) <= (layer2_outputs(898)) or (layer2_outputs(4910));
    outputs(9217) <= layer2_outputs(12767);
    outputs(9218) <= not(layer2_outputs(3171));
    outputs(9219) <= (layer2_outputs(10242)) xor (layer2_outputs(10125));
    outputs(9220) <= (layer2_outputs(5913)) xor (layer2_outputs(2593));
    outputs(9221) <= (layer2_outputs(670)) or (layer2_outputs(10809));
    outputs(9222) <= layer2_outputs(9370);
    outputs(9223) <= layer2_outputs(10709);
    outputs(9224) <= not(layer2_outputs(6584));
    outputs(9225) <= not(layer2_outputs(6018));
    outputs(9226) <= not((layer2_outputs(3206)) and (layer2_outputs(3302)));
    outputs(9227) <= not((layer2_outputs(6219)) xor (layer2_outputs(12492)));
    outputs(9228) <= (layer2_outputs(5784)) and not (layer2_outputs(5800));
    outputs(9229) <= not(layer2_outputs(8333));
    outputs(9230) <= layer2_outputs(1291);
    outputs(9231) <= layer2_outputs(7055);
    outputs(9232) <= not((layer2_outputs(1246)) xor (layer2_outputs(7896)));
    outputs(9233) <= not(layer2_outputs(865));
    outputs(9234) <= layer2_outputs(2757);
    outputs(9235) <= not(layer2_outputs(328));
    outputs(9236) <= not(layer2_outputs(3305));
    outputs(9237) <= not((layer2_outputs(11614)) or (layer2_outputs(10216)));
    outputs(9238) <= not(layer2_outputs(8116)) or (layer2_outputs(5368));
    outputs(9239) <= not(layer2_outputs(1388));
    outputs(9240) <= not(layer2_outputs(8210)) or (layer2_outputs(1397));
    outputs(9241) <= (layer2_outputs(2654)) or (layer2_outputs(106));
    outputs(9242) <= not(layer2_outputs(9271));
    outputs(9243) <= not((layer2_outputs(1598)) xor (layer2_outputs(11162)));
    outputs(9244) <= (layer2_outputs(2070)) and not (layer2_outputs(7802));
    outputs(9245) <= not(layer2_outputs(6939));
    outputs(9246) <= not(layer2_outputs(12752));
    outputs(9247) <= not(layer2_outputs(5317)) or (layer2_outputs(4134));
    outputs(9248) <= layer2_outputs(5277);
    outputs(9249) <= layer2_outputs(9962);
    outputs(9250) <= not((layer2_outputs(8226)) or (layer2_outputs(11045)));
    outputs(9251) <= layer2_outputs(7535);
    outputs(9252) <= not(layer2_outputs(4492));
    outputs(9253) <= layer2_outputs(10771);
    outputs(9254) <= layer2_outputs(3897);
    outputs(9255) <= not(layer2_outputs(4977));
    outputs(9256) <= not(layer2_outputs(8098));
    outputs(9257) <= not(layer2_outputs(7664));
    outputs(9258) <= layer2_outputs(7523);
    outputs(9259) <= (layer2_outputs(4917)) xor (layer2_outputs(8997));
    outputs(9260) <= not((layer2_outputs(7625)) or (layer2_outputs(11482)));
    outputs(9261) <= (layer2_outputs(11565)) xor (layer2_outputs(4649));
    outputs(9262) <= (layer2_outputs(7763)) xor (layer2_outputs(11812));
    outputs(9263) <= not(layer2_outputs(8840));
    outputs(9264) <= not((layer2_outputs(3579)) xor (layer2_outputs(5983)));
    outputs(9265) <= not((layer2_outputs(2574)) xor (layer2_outputs(5576)));
    outputs(9266) <= (layer2_outputs(8319)) xor (layer2_outputs(10994));
    outputs(9267) <= (layer2_outputs(11540)) xor (layer2_outputs(4233));
    outputs(9268) <= (layer2_outputs(494)) and (layer2_outputs(8213));
    outputs(9269) <= (layer2_outputs(6121)) xor (layer2_outputs(3219));
    outputs(9270) <= not(layer2_outputs(11965));
    outputs(9271) <= not((layer2_outputs(6344)) or (layer2_outputs(4712)));
    outputs(9272) <= not(layer2_outputs(8631)) or (layer2_outputs(6585));
    outputs(9273) <= (layer2_outputs(397)) xor (layer2_outputs(373));
    outputs(9274) <= layer2_outputs(2278);
    outputs(9275) <= not((layer2_outputs(5790)) xor (layer2_outputs(1272)));
    outputs(9276) <= not(layer2_outputs(3077));
    outputs(9277) <= (layer2_outputs(3207)) xor (layer2_outputs(5928));
    outputs(9278) <= not(layer2_outputs(5161));
    outputs(9279) <= (layer2_outputs(5932)) and not (layer2_outputs(4688));
    outputs(9280) <= not((layer2_outputs(8490)) xor (layer2_outputs(8711)));
    outputs(9281) <= (layer2_outputs(848)) xor (layer2_outputs(10727));
    outputs(9282) <= layer2_outputs(12583);
    outputs(9283) <= not(layer2_outputs(509));
    outputs(9284) <= not((layer2_outputs(7034)) xor (layer2_outputs(969)));
    outputs(9285) <= (layer2_outputs(1457)) and (layer2_outputs(11103));
    outputs(9286) <= layer2_outputs(7727);
    outputs(9287) <= not((layer2_outputs(6450)) xor (layer2_outputs(5724)));
    outputs(9288) <= not(layer2_outputs(10052));
    outputs(9289) <= not((layer2_outputs(2419)) xor (layer2_outputs(11762)));
    outputs(9290) <= layer2_outputs(3240);
    outputs(9291) <= layer2_outputs(12003);
    outputs(9292) <= not((layer2_outputs(12156)) xor (layer2_outputs(11863)));
    outputs(9293) <= not(layer2_outputs(5150));
    outputs(9294) <= (layer2_outputs(5035)) and not (layer2_outputs(2562));
    outputs(9295) <= layer2_outputs(7773);
    outputs(9296) <= layer2_outputs(9000);
    outputs(9297) <= not(layer2_outputs(9703));
    outputs(9298) <= layer2_outputs(9314);
    outputs(9299) <= (layer2_outputs(2361)) and (layer2_outputs(2452));
    outputs(9300) <= layer2_outputs(10793);
    outputs(9301) <= not(layer2_outputs(745)) or (layer2_outputs(5949));
    outputs(9302) <= not(layer2_outputs(7476));
    outputs(9303) <= layer2_outputs(11710);
    outputs(9304) <= layer2_outputs(8235);
    outputs(9305) <= (layer2_outputs(12441)) xor (layer2_outputs(11849));
    outputs(9306) <= not(layer2_outputs(246));
    outputs(9307) <= not(layer2_outputs(490));
    outputs(9308) <= not(layer2_outputs(2835));
    outputs(9309) <= layer2_outputs(5157);
    outputs(9310) <= not(layer2_outputs(9853));
    outputs(9311) <= not((layer2_outputs(6527)) xor (layer2_outputs(6408)));
    outputs(9312) <= not(layer2_outputs(6586));
    outputs(9313) <= layer2_outputs(1602);
    outputs(9314) <= (layer2_outputs(6812)) xor (layer2_outputs(12197));
    outputs(9315) <= (layer2_outputs(11085)) xor (layer2_outputs(2139));
    outputs(9316) <= not((layer2_outputs(2928)) xor (layer2_outputs(8038)));
    outputs(9317) <= (layer2_outputs(11204)) xor (layer2_outputs(9262));
    outputs(9318) <= not((layer2_outputs(11589)) xor (layer2_outputs(11816)));
    outputs(9319) <= not((layer2_outputs(438)) and (layer2_outputs(2502)));
    outputs(9320) <= not(layer2_outputs(6773));
    outputs(9321) <= not(layer2_outputs(2484));
    outputs(9322) <= not((layer2_outputs(1548)) xor (layer2_outputs(5563)));
    outputs(9323) <= (layer2_outputs(3324)) or (layer2_outputs(11956));
    outputs(9324) <= layer2_outputs(11414);
    outputs(9325) <= not(layer2_outputs(9550));
    outputs(9326) <= layer2_outputs(9502);
    outputs(9327) <= layer2_outputs(2468);
    outputs(9328) <= layer2_outputs(6389);
    outputs(9329) <= (layer2_outputs(10312)) xor (layer2_outputs(604));
    outputs(9330) <= not(layer2_outputs(3117));
    outputs(9331) <= not((layer2_outputs(5940)) and (layer2_outputs(8908)));
    outputs(9332) <= (layer2_outputs(7712)) xor (layer2_outputs(6184));
    outputs(9333) <= (layer2_outputs(2913)) xor (layer2_outputs(9760));
    outputs(9334) <= not((layer2_outputs(8130)) xor (layer2_outputs(3028)));
    outputs(9335) <= not((layer2_outputs(11828)) xor (layer2_outputs(3728)));
    outputs(9336) <= not((layer2_outputs(4009)) xor (layer2_outputs(10425)));
    outputs(9337) <= (layer2_outputs(12444)) xor (layer2_outputs(2758));
    outputs(9338) <= not((layer2_outputs(5101)) and (layer2_outputs(8119)));
    outputs(9339) <= (layer2_outputs(10498)) and not (layer2_outputs(2780));
    outputs(9340) <= not((layer2_outputs(5441)) xor (layer2_outputs(5918)));
    outputs(9341) <= not(layer2_outputs(368));
    outputs(9342) <= layer2_outputs(286);
    outputs(9343) <= layer2_outputs(3357);
    outputs(9344) <= not((layer2_outputs(9300)) xor (layer2_outputs(3447)));
    outputs(9345) <= layer2_outputs(4141);
    outputs(9346) <= layer2_outputs(5789);
    outputs(9347) <= not(layer2_outputs(4482));
    outputs(9348) <= not(layer2_outputs(4964));
    outputs(9349) <= not(layer2_outputs(9062));
    outputs(9350) <= not((layer2_outputs(181)) xor (layer2_outputs(3359)));
    outputs(9351) <= (layer2_outputs(11952)) and not (layer2_outputs(5813));
    outputs(9352) <= not((layer2_outputs(2610)) xor (layer2_outputs(1052)));
    outputs(9353) <= not((layer2_outputs(5424)) or (layer2_outputs(1993)));
    outputs(9354) <= (layer2_outputs(2606)) xor (layer2_outputs(2944));
    outputs(9355) <= not((layer2_outputs(12143)) xor (layer2_outputs(9108)));
    outputs(9356) <= not(layer2_outputs(9571));
    outputs(9357) <= (layer2_outputs(1800)) and not (layer2_outputs(4833));
    outputs(9358) <= not(layer2_outputs(10094));
    outputs(9359) <= not(layer2_outputs(3337));
    outputs(9360) <= layer2_outputs(2632);
    outputs(9361) <= not((layer2_outputs(3122)) xor (layer2_outputs(8128)));
    outputs(9362) <= not(layer2_outputs(9892));
    outputs(9363) <= layer2_outputs(5537);
    outputs(9364) <= layer2_outputs(2329);
    outputs(9365) <= not((layer2_outputs(2073)) xor (layer2_outputs(6414)));
    outputs(9366) <= (layer2_outputs(12671)) and not (layer2_outputs(6414));
    outputs(9367) <= layer2_outputs(1756);
    outputs(9368) <= layer2_outputs(8258);
    outputs(9369) <= layer2_outputs(297);
    outputs(9370) <= layer2_outputs(10443);
    outputs(9371) <= not(layer2_outputs(4829)) or (layer2_outputs(5622));
    outputs(9372) <= layer2_outputs(1652);
    outputs(9373) <= layer2_outputs(6264);
    outputs(9374) <= layer2_outputs(6105);
    outputs(9375) <= (layer2_outputs(3654)) and not (layer2_outputs(3465));
    outputs(9376) <= not(layer2_outputs(6688));
    outputs(9377) <= (layer2_outputs(11355)) xor (layer2_outputs(9065));
    outputs(9378) <= (layer2_outputs(7521)) xor (layer2_outputs(2296));
    outputs(9379) <= not(layer2_outputs(3761));
    outputs(9380) <= not(layer2_outputs(4418));
    outputs(9381) <= layer2_outputs(2639);
    outputs(9382) <= layer2_outputs(1342);
    outputs(9383) <= not(layer2_outputs(8931));
    outputs(9384) <= not((layer2_outputs(8115)) xor (layer2_outputs(2683)));
    outputs(9385) <= not((layer2_outputs(8137)) xor (layer2_outputs(3309)));
    outputs(9386) <= not((layer2_outputs(6553)) or (layer2_outputs(12096)));
    outputs(9387) <= not((layer2_outputs(12429)) or (layer2_outputs(6382)));
    outputs(9388) <= not(layer2_outputs(11027));
    outputs(9389) <= layer2_outputs(6634);
    outputs(9390) <= not((layer2_outputs(12293)) xor (layer2_outputs(2863)));
    outputs(9391) <= (layer2_outputs(4723)) xor (layer2_outputs(7939));
    outputs(9392) <= layer2_outputs(2475);
    outputs(9393) <= not((layer2_outputs(9010)) or (layer2_outputs(12395)));
    outputs(9394) <= (layer2_outputs(2653)) and (layer2_outputs(5222));
    outputs(9395) <= layer2_outputs(798);
    outputs(9396) <= layer2_outputs(10119);
    outputs(9397) <= (layer2_outputs(11652)) xor (layer2_outputs(4629));
    outputs(9398) <= not(layer2_outputs(2111));
    outputs(9399) <= not(layer2_outputs(6649));
    outputs(9400) <= (layer2_outputs(2558)) xor (layer2_outputs(2661));
    outputs(9401) <= not((layer2_outputs(11979)) xor (layer2_outputs(3746)));
    outputs(9402) <= not((layer2_outputs(4283)) xor (layer2_outputs(3247)));
    outputs(9403) <= (layer2_outputs(6971)) or (layer2_outputs(7528));
    outputs(9404) <= not((layer2_outputs(5496)) xor (layer2_outputs(10617)));
    outputs(9405) <= not(layer2_outputs(1831));
    outputs(9406) <= (layer2_outputs(6084)) xor (layer2_outputs(3583));
    outputs(9407) <= not((layer2_outputs(174)) or (layer2_outputs(2192)));
    outputs(9408) <= layer2_outputs(7222);
    outputs(9409) <= not((layer2_outputs(11657)) or (layer2_outputs(764)));
    outputs(9410) <= layer2_outputs(6024);
    outputs(9411) <= (layer2_outputs(3954)) and not (layer2_outputs(9900));
    outputs(9412) <= (layer2_outputs(2636)) xor (layer2_outputs(1475));
    outputs(9413) <= not((layer2_outputs(11809)) xor (layer2_outputs(3561)));
    outputs(9414) <= not(layer2_outputs(9552));
    outputs(9415) <= not((layer2_outputs(972)) or (layer2_outputs(3703)));
    outputs(9416) <= not((layer2_outputs(138)) xor (layer2_outputs(9207)));
    outputs(9417) <= layer2_outputs(10700);
    outputs(9418) <= layer2_outputs(10909);
    outputs(9419) <= not(layer2_outputs(5045));
    outputs(9420) <= layer2_outputs(11941);
    outputs(9421) <= layer2_outputs(12424);
    outputs(9422) <= not((layer2_outputs(786)) xor (layer2_outputs(8910)));
    outputs(9423) <= (layer2_outputs(5026)) or (layer2_outputs(12330));
    outputs(9424) <= not(layer2_outputs(3512));
    outputs(9425) <= not((layer2_outputs(1336)) xor (layer2_outputs(1802)));
    outputs(9426) <= (layer2_outputs(7600)) xor (layer2_outputs(872));
    outputs(9427) <= layer2_outputs(11351);
    outputs(9428) <= not(layer2_outputs(5143));
    outputs(9429) <= not(layer2_outputs(1539));
    outputs(9430) <= not((layer2_outputs(1342)) xor (layer2_outputs(757)));
    outputs(9431) <= not(layer2_outputs(1640));
    outputs(9432) <= (layer2_outputs(7468)) and not (layer2_outputs(5817));
    outputs(9433) <= not(layer2_outputs(11946));
    outputs(9434) <= (layer2_outputs(2268)) and not (layer2_outputs(7461));
    outputs(9435) <= not(layer2_outputs(9929));
    outputs(9436) <= layer2_outputs(6570);
    outputs(9437) <= (layer2_outputs(9940)) xor (layer2_outputs(5997));
    outputs(9438) <= layer2_outputs(5666);
    outputs(9439) <= (layer2_outputs(3154)) and not (layer2_outputs(9475));
    outputs(9440) <= layer2_outputs(12499);
    outputs(9441) <= not(layer2_outputs(9737));
    outputs(9442) <= (layer2_outputs(10039)) and (layer2_outputs(2804));
    outputs(9443) <= layer2_outputs(2082);
    outputs(9444) <= not(layer2_outputs(9673));
    outputs(9445) <= layer2_outputs(2007);
    outputs(9446) <= not(layer2_outputs(10616));
    outputs(9447) <= (layer2_outputs(1642)) or (layer2_outputs(5247));
    outputs(9448) <= not((layer2_outputs(8982)) xor (layer2_outputs(609)));
    outputs(9449) <= (layer2_outputs(3914)) and not (layer2_outputs(4760));
    outputs(9450) <= not((layer2_outputs(1398)) xor (layer2_outputs(11974)));
    outputs(9451) <= layer2_outputs(12282);
    outputs(9452) <= not(layer2_outputs(6596));
    outputs(9453) <= (layer2_outputs(901)) or (layer2_outputs(11515));
    outputs(9454) <= not(layer2_outputs(11474));
    outputs(9455) <= not(layer2_outputs(1867));
    outputs(9456) <= not(layer2_outputs(12690));
    outputs(9457) <= layer2_outputs(4625);
    outputs(9458) <= not(layer2_outputs(11656));
    outputs(9459) <= not(layer2_outputs(7284));
    outputs(9460) <= not(layer2_outputs(11501));
    outputs(9461) <= not(layer2_outputs(6918));
    outputs(9462) <= not(layer2_outputs(1137));
    outputs(9463) <= not((layer2_outputs(9291)) xor (layer2_outputs(3783)));
    outputs(9464) <= layer2_outputs(2307);
    outputs(9465) <= layer2_outputs(182);
    outputs(9466) <= layer2_outputs(4819);
    outputs(9467) <= not(layer2_outputs(2537));
    outputs(9468) <= not((layer2_outputs(1931)) xor (layer2_outputs(5349)));
    outputs(9469) <= (layer2_outputs(8114)) xor (layer2_outputs(3918));
    outputs(9470) <= (layer2_outputs(1572)) and (layer2_outputs(6358));
    outputs(9471) <= (layer2_outputs(3174)) xor (layer2_outputs(8854));
    outputs(9472) <= layer2_outputs(7139);
    outputs(9473) <= (layer2_outputs(2846)) and (layer2_outputs(1179));
    outputs(9474) <= not(layer2_outputs(3903));
    outputs(9475) <= not(layer2_outputs(11940));
    outputs(9476) <= not(layer2_outputs(12141));
    outputs(9477) <= layer2_outputs(11453);
    outputs(9478) <= layer2_outputs(8802);
    outputs(9479) <= not(layer2_outputs(1791));
    outputs(9480) <= layer2_outputs(6468);
    outputs(9481) <= layer2_outputs(2198);
    outputs(9482) <= layer2_outputs(1748);
    outputs(9483) <= (layer2_outputs(4799)) and not (layer2_outputs(8561));
    outputs(9484) <= (layer2_outputs(6562)) xor (layer2_outputs(5460));
    outputs(9485) <= not(layer2_outputs(1137));
    outputs(9486) <= layer2_outputs(3493);
    outputs(9487) <= not((layer2_outputs(1946)) or (layer2_outputs(6287)));
    outputs(9488) <= layer2_outputs(10372);
    outputs(9489) <= (layer2_outputs(2218)) or (layer2_outputs(7762));
    outputs(9490) <= (layer2_outputs(12119)) xor (layer2_outputs(10848));
    outputs(9491) <= not(layer2_outputs(9931));
    outputs(9492) <= layer2_outputs(5089);
    outputs(9493) <= not(layer2_outputs(4171));
    outputs(9494) <= (layer2_outputs(4083)) xor (layer2_outputs(10131));
    outputs(9495) <= layer2_outputs(8162);
    outputs(9496) <= layer2_outputs(12109);
    outputs(9497) <= not(layer2_outputs(12114)) or (layer2_outputs(7230));
    outputs(9498) <= not(layer2_outputs(3143));
    outputs(9499) <= not(layer2_outputs(1278));
    outputs(9500) <= not((layer2_outputs(2997)) xor (layer2_outputs(6339)));
    outputs(9501) <= not((layer2_outputs(8938)) and (layer2_outputs(7363)));
    outputs(9502) <= not(layer2_outputs(8754));
    outputs(9503) <= not(layer2_outputs(2674));
    outputs(9504) <= (layer2_outputs(8045)) and not (layer2_outputs(11854));
    outputs(9505) <= not(layer2_outputs(7023));
    outputs(9506) <= not((layer2_outputs(9870)) and (layer2_outputs(2831)));
    outputs(9507) <= layer2_outputs(8567);
    outputs(9508) <= not(layer2_outputs(1521));
    outputs(9509) <= layer2_outputs(3462);
    outputs(9510) <= (layer2_outputs(10637)) xor (layer2_outputs(224));
    outputs(9511) <= layer2_outputs(4032);
    outputs(9512) <= layer2_outputs(9983);
    outputs(9513) <= not(layer2_outputs(7530));
    outputs(9514) <= layer2_outputs(4018);
    outputs(9515) <= not(layer2_outputs(10613));
    outputs(9516) <= layer2_outputs(2118);
    outputs(9517) <= not(layer2_outputs(4175));
    outputs(9518) <= not(layer2_outputs(3670));
    outputs(9519) <= layer2_outputs(8297);
    outputs(9520) <= (layer2_outputs(2216)) xor (layer2_outputs(12069));
    outputs(9521) <= not(layer2_outputs(7394)) or (layer2_outputs(12619));
    outputs(9522) <= not((layer2_outputs(10393)) or (layer2_outputs(1638)));
    outputs(9523) <= layer2_outputs(4583);
    outputs(9524) <= not(layer2_outputs(6350));
    outputs(9525) <= (layer2_outputs(12553)) xor (layer2_outputs(8806));
    outputs(9526) <= not((layer2_outputs(5484)) xor (layer2_outputs(7409)));
    outputs(9527) <= layer2_outputs(6996);
    outputs(9528) <= not(layer2_outputs(8553));
    outputs(9529) <= not(layer2_outputs(9667));
    outputs(9530) <= layer2_outputs(766);
    outputs(9531) <= not(layer2_outputs(11450));
    outputs(9532) <= layer2_outputs(412);
    outputs(9533) <= not((layer2_outputs(8573)) xor (layer2_outputs(5870)));
    outputs(9534) <= layer2_outputs(9792);
    outputs(9535) <= not((layer2_outputs(10467)) xor (layer2_outputs(8314)));
    outputs(9536) <= not(layer2_outputs(6245));
    outputs(9537) <= not(layer2_outputs(4515));
    outputs(9538) <= not(layer2_outputs(8373));
    outputs(9539) <= not(layer2_outputs(1555));
    outputs(9540) <= layer2_outputs(12167);
    outputs(9541) <= not(layer2_outputs(3256));
    outputs(9542) <= not(layer2_outputs(9838));
    outputs(9543) <= not(layer2_outputs(7779));
    outputs(9544) <= not(layer2_outputs(10588));
    outputs(9545) <= layer2_outputs(10097);
    outputs(9546) <= not((layer2_outputs(6946)) xor (layer2_outputs(2066)));
    outputs(9547) <= not(layer2_outputs(10565));
    outputs(9548) <= not(layer2_outputs(5646));
    outputs(9549) <= not(layer2_outputs(11147));
    outputs(9550) <= not(layer2_outputs(10916));
    outputs(9551) <= (layer2_outputs(8369)) and not (layer2_outputs(2203));
    outputs(9552) <= not(layer2_outputs(4702));
    outputs(9553) <= not(layer2_outputs(7954));
    outputs(9554) <= (layer2_outputs(6743)) and not (layer2_outputs(10741));
    outputs(9555) <= not(layer2_outputs(10880));
    outputs(9556) <= not(layer2_outputs(4016)) or (layer2_outputs(10304));
    outputs(9557) <= not((layer2_outputs(5860)) xor (layer2_outputs(6597)));
    outputs(9558) <= layer2_outputs(10838);
    outputs(9559) <= not((layer2_outputs(344)) xor (layer2_outputs(3957)));
    outputs(9560) <= not(layer2_outputs(6490)) or (layer2_outputs(8298));
    outputs(9561) <= (layer2_outputs(4661)) xor (layer2_outputs(1107));
    outputs(9562) <= not(layer2_outputs(4777));
    outputs(9563) <= (layer2_outputs(6566)) or (layer2_outputs(10914));
    outputs(9564) <= not(layer2_outputs(2621));
    outputs(9565) <= layer2_outputs(3780);
    outputs(9566) <= layer2_outputs(4421);
    outputs(9567) <= (layer2_outputs(4679)) xor (layer2_outputs(9577));
    outputs(9568) <= layer2_outputs(7197);
    outputs(9569) <= (layer2_outputs(2554)) xor (layer2_outputs(3157));
    outputs(9570) <= layer2_outputs(10133);
    outputs(9571) <= not(layer2_outputs(131));
    outputs(9572) <= not(layer2_outputs(6039));
    outputs(9573) <= layer2_outputs(11415);
    outputs(9574) <= layer2_outputs(7913);
    outputs(9575) <= (layer2_outputs(2351)) and not (layer2_outputs(12301));
    outputs(9576) <= layer2_outputs(5836);
    outputs(9577) <= (layer2_outputs(10830)) xor (layer2_outputs(5142));
    outputs(9578) <= layer2_outputs(2880);
    outputs(9579) <= (layer2_outputs(6668)) and (layer2_outputs(6483));
    outputs(9580) <= not(layer2_outputs(151));
    outputs(9581) <= layer2_outputs(11901);
    outputs(9582) <= not(layer2_outputs(3163)) or (layer2_outputs(3706));
    outputs(9583) <= (layer2_outputs(5946)) and not (layer2_outputs(6321));
    outputs(9584) <= layer2_outputs(6307);
    outputs(9585) <= not((layer2_outputs(12783)) or (layer2_outputs(12761)));
    outputs(9586) <= layer2_outputs(11085);
    outputs(9587) <= not(layer2_outputs(7302)) or (layer2_outputs(12492));
    outputs(9588) <= not(layer2_outputs(9378));
    outputs(9589) <= layer2_outputs(7376);
    outputs(9590) <= layer2_outputs(4114);
    outputs(9591) <= layer2_outputs(8818);
    outputs(9592) <= layer2_outputs(10800);
    outputs(9593) <= (layer2_outputs(930)) xor (layer2_outputs(7126));
    outputs(9594) <= not((layer2_outputs(9985)) or (layer2_outputs(10622)));
    outputs(9595) <= layer2_outputs(9716);
    outputs(9596) <= layer2_outputs(4997);
    outputs(9597) <= not((layer2_outputs(4860)) xor (layer2_outputs(9017)));
    outputs(9598) <= layer2_outputs(8308);
    outputs(9599) <= layer2_outputs(7516);
    outputs(9600) <= layer2_outputs(5545);
    outputs(9601) <= layer2_outputs(5478);
    outputs(9602) <= (layer2_outputs(1128)) xor (layer2_outputs(6131));
    outputs(9603) <= not((layer2_outputs(9434)) xor (layer2_outputs(721)));
    outputs(9604) <= not(layer2_outputs(4155));
    outputs(9605) <= layer2_outputs(4875);
    outputs(9606) <= (layer2_outputs(4790)) xor (layer2_outputs(10150));
    outputs(9607) <= not(layer2_outputs(6972));
    outputs(9608) <= layer2_outputs(11695);
    outputs(9609) <= not(layer2_outputs(4801));
    outputs(9610) <= layer2_outputs(10871);
    outputs(9611) <= not(layer2_outputs(1867));
    outputs(9612) <= layer2_outputs(1220);
    outputs(9613) <= layer2_outputs(12451);
    outputs(9614) <= layer2_outputs(3606);
    outputs(9615) <= not(layer2_outputs(5119));
    outputs(9616) <= not(layer2_outputs(5512));
    outputs(9617) <= (layer2_outputs(897)) xor (layer2_outputs(1875));
    outputs(9618) <= not(layer2_outputs(7829));
    outputs(9619) <= (layer2_outputs(6816)) xor (layer2_outputs(8979));
    outputs(9620) <= not((layer2_outputs(5892)) or (layer2_outputs(5978)));
    outputs(9621) <= not(layer2_outputs(8809));
    outputs(9622) <= not(layer2_outputs(4810));
    outputs(9623) <= (layer2_outputs(4347)) xor (layer2_outputs(2561));
    outputs(9624) <= not(layer2_outputs(11961));
    outputs(9625) <= layer2_outputs(1739);
    outputs(9626) <= layer2_outputs(10444);
    outputs(9627) <= (layer2_outputs(2537)) xor (layer2_outputs(2174));
    outputs(9628) <= (layer2_outputs(996)) xor (layer2_outputs(3388));
    outputs(9629) <= layer2_outputs(6478);
    outputs(9630) <= (layer2_outputs(12233)) and (layer2_outputs(6292));
    outputs(9631) <= not(layer2_outputs(9893));
    outputs(9632) <= layer2_outputs(9962);
    outputs(9633) <= (layer2_outputs(2572)) xor (layer2_outputs(1884));
    outputs(9634) <= (layer2_outputs(6529)) or (layer2_outputs(12529));
    outputs(9635) <= not(layer2_outputs(2752));
    outputs(9636) <= not(layer2_outputs(2796));
    outputs(9637) <= layer2_outputs(6513);
    outputs(9638) <= layer2_outputs(3542);
    outputs(9639) <= not(layer2_outputs(5573));
    outputs(9640) <= (layer2_outputs(2093)) xor (layer2_outputs(5987));
    outputs(9641) <= layer2_outputs(12547);
    outputs(9642) <= layer2_outputs(9422);
    outputs(9643) <= layer2_outputs(10645);
    outputs(9644) <= layer2_outputs(2133);
    outputs(9645) <= not(layer2_outputs(7078));
    outputs(9646) <= layer2_outputs(9163);
    outputs(9647) <= layer2_outputs(9277);
    outputs(9648) <= layer2_outputs(12414);
    outputs(9649) <= (layer2_outputs(7206)) xor (layer2_outputs(244));
    outputs(9650) <= not(layer2_outputs(8826));
    outputs(9651) <= not(layer2_outputs(2953));
    outputs(9652) <= not(layer2_outputs(1831));
    outputs(9653) <= layer2_outputs(2081);
    outputs(9654) <= (layer2_outputs(489)) and (layer2_outputs(2371));
    outputs(9655) <= (layer2_outputs(4467)) xor (layer2_outputs(4325));
    outputs(9656) <= layer2_outputs(5096);
    outputs(9657) <= layer2_outputs(12596);
    outputs(9658) <= not(layer2_outputs(7490));
    outputs(9659) <= layer2_outputs(4568);
    outputs(9660) <= (layer2_outputs(9157)) xor (layer2_outputs(11325));
    outputs(9661) <= not((layer2_outputs(9734)) xor (layer2_outputs(6634)));
    outputs(9662) <= not(layer2_outputs(8826));
    outputs(9663) <= layer2_outputs(9594);
    outputs(9664) <= not(layer2_outputs(1811));
    outputs(9665) <= not(layer2_outputs(12690));
    outputs(9666) <= not(layer2_outputs(938));
    outputs(9667) <= (layer2_outputs(75)) xor (layer2_outputs(8447));
    outputs(9668) <= not(layer2_outputs(4772));
    outputs(9669) <= (layer2_outputs(6017)) xor (layer2_outputs(10403));
    outputs(9670) <= not(layer2_outputs(5417));
    outputs(9671) <= not((layer2_outputs(10699)) or (layer2_outputs(11305)));
    outputs(9672) <= not(layer2_outputs(4463));
    outputs(9673) <= layer2_outputs(304);
    outputs(9674) <= not((layer2_outputs(1479)) xor (layer2_outputs(3812)));
    outputs(9675) <= (layer2_outputs(6532)) xor (layer2_outputs(7497));
    outputs(9676) <= (layer2_outputs(2656)) xor (layer2_outputs(7398));
    outputs(9677) <= not((layer2_outputs(2145)) xor (layer2_outputs(3486)));
    outputs(9678) <= not((layer2_outputs(1632)) and (layer2_outputs(1332)));
    outputs(9679) <= (layer2_outputs(7993)) and not (layer2_outputs(6854));
    outputs(9680) <= (layer2_outputs(1801)) xor (layer2_outputs(2413));
    outputs(9681) <= not(layer2_outputs(8999));
    outputs(9682) <= not(layer2_outputs(916));
    outputs(9683) <= not(layer2_outputs(2496)) or (layer2_outputs(10822));
    outputs(9684) <= (layer2_outputs(2526)) xor (layer2_outputs(3202));
    outputs(9685) <= layer2_outputs(9661);
    outputs(9686) <= not((layer2_outputs(217)) xor (layer2_outputs(4550)));
    outputs(9687) <= layer2_outputs(139);
    outputs(9688) <= layer2_outputs(10722);
    outputs(9689) <= not(layer2_outputs(7246)) or (layer2_outputs(624));
    outputs(9690) <= not(layer2_outputs(12620));
    outputs(9691) <= not(layer2_outputs(10784));
    outputs(9692) <= (layer2_outputs(12715)) xor (layer2_outputs(2260));
    outputs(9693) <= (layer2_outputs(7069)) and not (layer2_outputs(8587));
    outputs(9694) <= not((layer2_outputs(11634)) xor (layer2_outputs(1094)));
    outputs(9695) <= layer2_outputs(12055);
    outputs(9696) <= layer2_outputs(5228);
    outputs(9697) <= layer2_outputs(2072);
    outputs(9698) <= not(layer2_outputs(10448));
    outputs(9699) <= layer2_outputs(3250);
    outputs(9700) <= (layer2_outputs(4253)) xor (layer2_outputs(2726));
    outputs(9701) <= not(layer2_outputs(3699));
    outputs(9702) <= not(layer2_outputs(1650)) or (layer2_outputs(10909));
    outputs(9703) <= not((layer2_outputs(3535)) or (layer2_outputs(6795)));
    outputs(9704) <= (layer2_outputs(11069)) xor (layer2_outputs(6824));
    outputs(9705) <= layer2_outputs(8290);
    outputs(9706) <= not((layer2_outputs(5514)) xor (layer2_outputs(9980)));
    outputs(9707) <= not((layer2_outputs(9639)) xor (layer2_outputs(7177)));
    outputs(9708) <= not(layer2_outputs(12717));
    outputs(9709) <= (layer2_outputs(8522)) xor (layer2_outputs(10789));
    outputs(9710) <= not(layer2_outputs(1667));
    outputs(9711) <= (layer2_outputs(10728)) and not (layer2_outputs(1707));
    outputs(9712) <= not((layer2_outputs(9352)) or (layer2_outputs(1699)));
    outputs(9713) <= not((layer2_outputs(5956)) xor (layer2_outputs(4633)));
    outputs(9714) <= layer2_outputs(4545);
    outputs(9715) <= layer2_outputs(9004);
    outputs(9716) <= not(layer2_outputs(4320));
    outputs(9717) <= not(layer2_outputs(11656));
    outputs(9718) <= (layer2_outputs(8491)) and not (layer2_outputs(8766));
    outputs(9719) <= (layer2_outputs(2101)) and not (layer2_outputs(2314));
    outputs(9720) <= not((layer2_outputs(4941)) or (layer2_outputs(7507)));
    outputs(9721) <= layer2_outputs(9857);
    outputs(9722) <= layer2_outputs(12593);
    outputs(9723) <= not((layer2_outputs(1974)) and (layer2_outputs(8681)));
    outputs(9724) <= layer2_outputs(8775);
    outputs(9725) <= not(layer2_outputs(11139)) or (layer2_outputs(7700));
    outputs(9726) <= not(layer2_outputs(5290));
    outputs(9727) <= layer2_outputs(9358);
    outputs(9728) <= (layer2_outputs(8577)) and not (layer2_outputs(6763));
    outputs(9729) <= layer2_outputs(452);
    outputs(9730) <= not((layer2_outputs(8122)) or (layer2_outputs(12442)));
    outputs(9731) <= layer2_outputs(1580);
    outputs(9732) <= layer2_outputs(98);
    outputs(9733) <= (layer2_outputs(12379)) or (layer2_outputs(6157));
    outputs(9734) <= (layer2_outputs(4486)) xor (layer2_outputs(11369));
    outputs(9735) <= not((layer2_outputs(6241)) or (layer2_outputs(8554)));
    outputs(9736) <= layer2_outputs(3323);
    outputs(9737) <= (layer2_outputs(2007)) and (layer2_outputs(9955));
    outputs(9738) <= (layer2_outputs(934)) and not (layer2_outputs(2191));
    outputs(9739) <= not(layer2_outputs(10110));
    outputs(9740) <= not((layer2_outputs(5898)) xor (layer2_outputs(3665)));
    outputs(9741) <= layer2_outputs(11093);
    outputs(9742) <= layer2_outputs(3089);
    outputs(9743) <= not(layer2_outputs(9580));
    outputs(9744) <= not(layer2_outputs(6362));
    outputs(9745) <= layer2_outputs(11651);
    outputs(9746) <= layer2_outputs(7063);
    outputs(9747) <= not(layer2_outputs(9338));
    outputs(9748) <= not(layer2_outputs(6753));
    outputs(9749) <= not((layer2_outputs(4554)) or (layer2_outputs(11064)));
    outputs(9750) <= layer2_outputs(7607);
    outputs(9751) <= layer2_outputs(10195);
    outputs(9752) <= layer2_outputs(9102);
    outputs(9753) <= layer2_outputs(4967);
    outputs(9754) <= not(layer2_outputs(7082));
    outputs(9755) <= not(layer2_outputs(12253));
    outputs(9756) <= not(layer2_outputs(7589)) or (layer2_outputs(293));
    outputs(9757) <= not(layer2_outputs(2116));
    outputs(9758) <= not((layer2_outputs(7841)) or (layer2_outputs(8887)));
    outputs(9759) <= (layer2_outputs(104)) xor (layer2_outputs(4506));
    outputs(9760) <= not((layer2_outputs(5627)) or (layer2_outputs(3742)));
    outputs(9761) <= not(layer2_outputs(10920));
    outputs(9762) <= not((layer2_outputs(9901)) or (layer2_outputs(6939)));
    outputs(9763) <= (layer2_outputs(5360)) xor (layer2_outputs(3794));
    outputs(9764) <= (layer2_outputs(5357)) xor (layer2_outputs(11770));
    outputs(9765) <= not((layer2_outputs(4364)) or (layer2_outputs(91)));
    outputs(9766) <= (layer2_outputs(3223)) and not (layer2_outputs(5033));
    outputs(9767) <= (layer2_outputs(9396)) xor (layer2_outputs(12727));
    outputs(9768) <= layer2_outputs(2288);
    outputs(9769) <= (layer2_outputs(2158)) xor (layer2_outputs(11155));
    outputs(9770) <= not(layer2_outputs(8047));
    outputs(9771) <= not(layer2_outputs(1889));
    outputs(9772) <= not(layer2_outputs(1895));
    outputs(9773) <= not(layer2_outputs(8804));
    outputs(9774) <= layer2_outputs(4179);
    outputs(9775) <= not((layer2_outputs(8894)) xor (layer2_outputs(191)));
    outputs(9776) <= not((layer2_outputs(2214)) xor (layer2_outputs(8977)));
    outputs(9777) <= not(layer2_outputs(9522));
    outputs(9778) <= (layer2_outputs(550)) xor (layer2_outputs(8214));
    outputs(9779) <= layer2_outputs(8018);
    outputs(9780) <= layer2_outputs(6291);
    outputs(9781) <= (layer2_outputs(3124)) or (layer2_outputs(7194));
    outputs(9782) <= not(layer2_outputs(10424));
    outputs(9783) <= (layer2_outputs(6645)) and (layer2_outputs(4563));
    outputs(9784) <= not(layer2_outputs(1539));
    outputs(9785) <= (layer2_outputs(11299)) and not (layer2_outputs(6055));
    outputs(9786) <= not(layer2_outputs(9807));
    outputs(9787) <= layer2_outputs(61);
    outputs(9788) <= not(layer2_outputs(3328));
    outputs(9789) <= not(layer2_outputs(1390));
    outputs(9790) <= not(layer2_outputs(971));
    outputs(9791) <= (layer2_outputs(843)) and not (layer2_outputs(7491));
    outputs(9792) <= (layer2_outputs(10552)) and not (layer2_outputs(7859));
    outputs(9793) <= layer2_outputs(1565);
    outputs(9794) <= not(layer2_outputs(7783));
    outputs(9795) <= not((layer2_outputs(5907)) xor (layer2_outputs(12437)));
    outputs(9796) <= not(layer2_outputs(6643));
    outputs(9797) <= (layer2_outputs(6023)) and (layer2_outputs(3158));
    outputs(9798) <= layer2_outputs(9322);
    outputs(9799) <= not((layer2_outputs(9428)) xor (layer2_outputs(5630)));
    outputs(9800) <= (layer2_outputs(7496)) xor (layer2_outputs(7146));
    outputs(9801) <= layer2_outputs(2803);
    outputs(9802) <= not(layer2_outputs(3521)) or (layer2_outputs(7612));
    outputs(9803) <= not(layer2_outputs(1979));
    outputs(9804) <= (layer2_outputs(7769)) and not (layer2_outputs(7973));
    outputs(9805) <= layer2_outputs(3297);
    outputs(9806) <= not(layer2_outputs(78));
    outputs(9807) <= (layer2_outputs(12152)) or (layer2_outputs(3970));
    outputs(9808) <= not(layer2_outputs(1984));
    outputs(9809) <= layer2_outputs(4638);
    outputs(9810) <= (layer2_outputs(10668)) xor (layer2_outputs(6858));
    outputs(9811) <= layer2_outputs(7843);
    outputs(9812) <= layer2_outputs(10382);
    outputs(9813) <= layer2_outputs(3891);
    outputs(9814) <= layer2_outputs(9744);
    outputs(9815) <= not(layer2_outputs(7176)) or (layer2_outputs(11653));
    outputs(9816) <= (layer2_outputs(10327)) or (layer2_outputs(8873));
    outputs(9817) <= (layer2_outputs(10059)) and (layer2_outputs(12742));
    outputs(9818) <= not((layer2_outputs(4343)) or (layer2_outputs(7381)));
    outputs(9819) <= not(layer2_outputs(5226));
    outputs(9820) <= (layer2_outputs(4046)) and not (layer2_outputs(6191));
    outputs(9821) <= not(layer2_outputs(6351));
    outputs(9822) <= not(layer2_outputs(1009));
    outputs(9823) <= layer2_outputs(8274);
    outputs(9824) <= layer2_outputs(6963);
    outputs(9825) <= not(layer2_outputs(5392));
    outputs(9826) <= not(layer2_outputs(5889));
    outputs(9827) <= layer2_outputs(11612);
    outputs(9828) <= layer2_outputs(12089);
    outputs(9829) <= not((layer2_outputs(10092)) or (layer2_outputs(5826)));
    outputs(9830) <= not((layer2_outputs(3634)) and (layer2_outputs(8078)));
    outputs(9831) <= layer2_outputs(11945);
    outputs(9832) <= not(layer2_outputs(3310));
    outputs(9833) <= layer2_outputs(11518);
    outputs(9834) <= layer2_outputs(173);
    outputs(9835) <= not(layer2_outputs(8289));
    outputs(9836) <= layer2_outputs(5212);
    outputs(9837) <= not((layer2_outputs(7904)) xor (layer2_outputs(9410)));
    outputs(9838) <= not(layer2_outputs(2703));
    outputs(9839) <= (layer2_outputs(1089)) and (layer2_outputs(3149));
    outputs(9840) <= not(layer2_outputs(351));
    outputs(9841) <= not(layer2_outputs(9800));
    outputs(9842) <= (layer2_outputs(3449)) xor (layer2_outputs(1963));
    outputs(9843) <= (layer2_outputs(1522)) xor (layer2_outputs(3727));
    outputs(9844) <= (layer2_outputs(9505)) xor (layer2_outputs(5166));
    outputs(9845) <= (layer2_outputs(8142)) and not (layer2_outputs(5850));
    outputs(9846) <= (layer2_outputs(8729)) and not (layer2_outputs(10328));
    outputs(9847) <= (layer2_outputs(8717)) and not (layer2_outputs(4037));
    outputs(9848) <= layer2_outputs(8973);
    outputs(9849) <= (layer2_outputs(11672)) and not (layer2_outputs(6937));
    outputs(9850) <= not(layer2_outputs(12483));
    outputs(9851) <= layer2_outputs(785);
    outputs(9852) <= not((layer2_outputs(3207)) or (layer2_outputs(7875)));
    outputs(9853) <= layer2_outputs(3429);
    outputs(9854) <= not(layer2_outputs(8254)) or (layer2_outputs(8343));
    outputs(9855) <= not(layer2_outputs(3858));
    outputs(9856) <= not(layer2_outputs(11323));
    outputs(9857) <= layer2_outputs(1455);
    outputs(9858) <= not(layer2_outputs(9722));
    outputs(9859) <= not(layer2_outputs(1509));
    outputs(9860) <= not(layer2_outputs(5512));
    outputs(9861) <= (layer2_outputs(6164)) and (layer2_outputs(5152));
    outputs(9862) <= not(layer2_outputs(8659)) or (layer2_outputs(12798));
    outputs(9863) <= not((layer2_outputs(5465)) and (layer2_outputs(4873)));
    outputs(9864) <= not(layer2_outputs(9999));
    outputs(9865) <= not(layer2_outputs(10734));
    outputs(9866) <= (layer2_outputs(1894)) and (layer2_outputs(10581));
    outputs(9867) <= not(layer2_outputs(2697)) or (layer2_outputs(8940));
    outputs(9868) <= layer2_outputs(5844);
    outputs(9869) <= layer2_outputs(5024);
    outputs(9870) <= not((layer2_outputs(7985)) xor (layer2_outputs(7925)));
    outputs(9871) <= not(layer2_outputs(7357));
    outputs(9872) <= not((layer2_outputs(1446)) xor (layer2_outputs(11416)));
    outputs(9873) <= layer2_outputs(7727);
    outputs(9874) <= not((layer2_outputs(9543)) xor (layer2_outputs(172)));
    outputs(9875) <= (layer2_outputs(2452)) xor (layer2_outputs(79));
    outputs(9876) <= not(layer2_outputs(7895));
    outputs(9877) <= not((layer2_outputs(2909)) and (layer2_outputs(3138)));
    outputs(9878) <= not((layer2_outputs(2225)) xor (layer2_outputs(5775)));
    outputs(9879) <= (layer2_outputs(560)) xor (layer2_outputs(9063));
    outputs(9880) <= (layer2_outputs(7951)) and not (layer2_outputs(7628));
    outputs(9881) <= not(layer2_outputs(7613));
    outputs(9882) <= layer2_outputs(6083);
    outputs(9883) <= not(layer2_outputs(828));
    outputs(9884) <= not(layer2_outputs(5683));
    outputs(9885) <= layer2_outputs(4324);
    outputs(9886) <= layer2_outputs(5105);
    outputs(9887) <= not((layer2_outputs(714)) xor (layer2_outputs(10237)));
    outputs(9888) <= layer2_outputs(3686);
    outputs(9889) <= (layer2_outputs(5064)) xor (layer2_outputs(1567));
    outputs(9890) <= not(layer2_outputs(2783));
    outputs(9891) <= layer2_outputs(10234);
    outputs(9892) <= (layer2_outputs(2429)) xor (layer2_outputs(9133));
    outputs(9893) <= layer2_outputs(2120);
    outputs(9894) <= (layer2_outputs(11669)) xor (layer2_outputs(12203));
    outputs(9895) <= layer2_outputs(7526);
    outputs(9896) <= not(layer2_outputs(8595));
    outputs(9897) <= layer2_outputs(6517);
    outputs(9898) <= layer2_outputs(108);
    outputs(9899) <= layer2_outputs(1504);
    outputs(9900) <= (layer2_outputs(12185)) xor (layer2_outputs(10831));
    outputs(9901) <= not(layer2_outputs(6360)) or (layer2_outputs(10672));
    outputs(9902) <= not((layer2_outputs(9843)) xor (layer2_outputs(12073)));
    outputs(9903) <= layer2_outputs(8886);
    outputs(9904) <= (layer2_outputs(7114)) or (layer2_outputs(7421));
    outputs(9905) <= (layer2_outputs(11701)) xor (layer2_outputs(7452));
    outputs(9906) <= (layer2_outputs(7910)) and not (layer2_outputs(7106));
    outputs(9907) <= not(layer2_outputs(5581));
    outputs(9908) <= (layer2_outputs(619)) xor (layer2_outputs(9685));
    outputs(9909) <= not((layer2_outputs(4117)) xor (layer2_outputs(3162)));
    outputs(9910) <= layer2_outputs(3974);
    outputs(9911) <= layer2_outputs(11704);
    outputs(9912) <= not(layer2_outputs(7255));
    outputs(9913) <= layer2_outputs(11257);
    outputs(9914) <= not(layer2_outputs(4752));
    outputs(9915) <= not((layer2_outputs(469)) xor (layer2_outputs(929)));
    outputs(9916) <= (layer2_outputs(1953)) and (layer2_outputs(7402));
    outputs(9917) <= layer2_outputs(7258);
    outputs(9918) <= not((layer2_outputs(6202)) xor (layer2_outputs(12463)));
    outputs(9919) <= not(layer2_outputs(4512));
    outputs(9920) <= (layer2_outputs(7975)) or (layer2_outputs(4625));
    outputs(9921) <= not(layer2_outputs(8753));
    outputs(9922) <= not(layer2_outputs(8773));
    outputs(9923) <= not(layer2_outputs(9911));
    outputs(9924) <= not(layer2_outputs(7530));
    outputs(9925) <= layer2_outputs(9587);
    outputs(9926) <= layer2_outputs(2741);
    outputs(9927) <= layer2_outputs(11964);
    outputs(9928) <= not(layer2_outputs(6686));
    outputs(9929) <= (layer2_outputs(10594)) xor (layer2_outputs(8778));
    outputs(9930) <= not((layer2_outputs(4439)) or (layer2_outputs(2838)));
    outputs(9931) <= layer2_outputs(9829);
    outputs(9932) <= layer2_outputs(7607);
    outputs(9933) <= layer2_outputs(11400);
    outputs(9934) <= not(layer2_outputs(2181));
    outputs(9935) <= not(layer2_outputs(2947));
    outputs(9936) <= layer2_outputs(1111);
    outputs(9937) <= not((layer2_outputs(9011)) xor (layer2_outputs(10987)));
    outputs(9938) <= (layer2_outputs(5868)) xor (layer2_outputs(10617));
    outputs(9939) <= not((layer2_outputs(1096)) and (layer2_outputs(9408)));
    outputs(9940) <= not((layer2_outputs(5409)) xor (layer2_outputs(7144)));
    outputs(9941) <= not(layer2_outputs(6706)) or (layer2_outputs(1844));
    outputs(9942) <= (layer2_outputs(11045)) xor (layer2_outputs(8744));
    outputs(9943) <= layer2_outputs(8148);
    outputs(9944) <= layer2_outputs(9048);
    outputs(9945) <= layer2_outputs(4032);
    outputs(9946) <= layer2_outputs(10519);
    outputs(9947) <= not(layer2_outputs(3917));
    outputs(9948) <= (layer2_outputs(12093)) and (layer2_outputs(10412));
    outputs(9949) <= not((layer2_outputs(5405)) and (layer2_outputs(8900)));
    outputs(9950) <= not((layer2_outputs(12730)) xor (layer2_outputs(3617)));
    outputs(9951) <= layer2_outputs(8302);
    outputs(9952) <= not(layer2_outputs(386));
    outputs(9953) <= not(layer2_outputs(2912));
    outputs(9954) <= layer2_outputs(8729);
    outputs(9955) <= layer2_outputs(12257);
    outputs(9956) <= not(layer2_outputs(2300));
    outputs(9957) <= layer2_outputs(1074);
    outputs(9958) <= (layer2_outputs(11523)) xor (layer2_outputs(261));
    outputs(9959) <= layer2_outputs(3188);
    outputs(9960) <= (layer2_outputs(6393)) and not (layer2_outputs(2186));
    outputs(9961) <= not((layer2_outputs(7945)) and (layer2_outputs(5884)));
    outputs(9962) <= not(layer2_outputs(4601)) or (layer2_outputs(4507));
    outputs(9963) <= (layer2_outputs(10266)) xor (layer2_outputs(6648));
    outputs(9964) <= (layer2_outputs(8548)) and not (layer2_outputs(322));
    outputs(9965) <= layer2_outputs(5158);
    outputs(9966) <= not(layer2_outputs(12213));
    outputs(9967) <= not(layer2_outputs(7022));
    outputs(9968) <= not((layer2_outputs(10872)) xor (layer2_outputs(5461)));
    outputs(9969) <= (layer2_outputs(2289)) and not (layer2_outputs(8725));
    outputs(9970) <= not(layer2_outputs(8029));
    outputs(9971) <= not((layer2_outputs(11847)) xor (layer2_outputs(6986)));
    outputs(9972) <= not(layer2_outputs(6591));
    outputs(9973) <= not(layer2_outputs(10453)) or (layer2_outputs(12225));
    outputs(9974) <= layer2_outputs(10767);
    outputs(9975) <= layer2_outputs(7588);
    outputs(9976) <= not(layer2_outputs(4458));
    outputs(9977) <= layer2_outputs(8534);
    outputs(9978) <= layer2_outputs(5447);
    outputs(9979) <= not(layer2_outputs(10815));
    outputs(9980) <= not((layer2_outputs(11360)) xor (layer2_outputs(9841)));
    outputs(9981) <= layer2_outputs(275);
    outputs(9982) <= not((layer2_outputs(9789)) xor (layer2_outputs(5776)));
    outputs(9983) <= (layer2_outputs(5441)) and not (layer2_outputs(427));
    outputs(9984) <= (layer2_outputs(3348)) xor (layer2_outputs(7270));
    outputs(9985) <= not(layer2_outputs(12030));
    outputs(9986) <= not(layer2_outputs(4727));
    outputs(9987) <= not(layer2_outputs(1879));
    outputs(9988) <= not((layer2_outputs(1592)) xor (layer2_outputs(11477)));
    outputs(9989) <= (layer2_outputs(5716)) xor (layer2_outputs(4091));
    outputs(9990) <= layer2_outputs(3197);
    outputs(9991) <= not(layer2_outputs(10859)) or (layer2_outputs(11377));
    outputs(9992) <= not((layer2_outputs(10423)) xor (layer2_outputs(10325)));
    outputs(9993) <= not((layer2_outputs(5271)) xor (layer2_outputs(9878)));
    outputs(9994) <= layer2_outputs(3095);
    outputs(9995) <= not((layer2_outputs(3152)) xor (layer2_outputs(2574)));
    outputs(9996) <= not(layer2_outputs(185));
    outputs(9997) <= not(layer2_outputs(10997));
    outputs(9998) <= layer2_outputs(4798);
    outputs(9999) <= not(layer2_outputs(8004));
    outputs(10000) <= layer2_outputs(8127);
    outputs(10001) <= (layer2_outputs(772)) xor (layer2_outputs(4094));
    outputs(10002) <= (layer2_outputs(10153)) xor (layer2_outputs(10856));
    outputs(10003) <= not((layer2_outputs(6530)) xor (layer2_outputs(11836)));
    outputs(10004) <= not(layer2_outputs(4394));
    outputs(10005) <= layer2_outputs(7773);
    outputs(10006) <= not(layer2_outputs(5730));
    outputs(10007) <= (layer2_outputs(5918)) xor (layer2_outputs(11839));
    outputs(10008) <= not(layer2_outputs(7119));
    outputs(10009) <= (layer2_outputs(12110)) and not (layer2_outputs(3518));
    outputs(10010) <= layer2_outputs(10647);
    outputs(10011) <= not(layer2_outputs(12027));
    outputs(10012) <= (layer2_outputs(11673)) and not (layer2_outputs(10904));
    outputs(10013) <= (layer2_outputs(10041)) xor (layer2_outputs(5217));
    outputs(10014) <= not(layer2_outputs(7728));
    outputs(10015) <= (layer2_outputs(1757)) xor (layer2_outputs(9330));
    outputs(10016) <= layer2_outputs(5694);
    outputs(10017) <= layer2_outputs(6289);
    outputs(10018) <= layer2_outputs(4696);
    outputs(10019) <= not(layer2_outputs(7572));
    outputs(10020) <= not((layer2_outputs(4883)) xor (layer2_outputs(9098)));
    outputs(10021) <= (layer2_outputs(12653)) xor (layer2_outputs(11618));
    outputs(10022) <= not(layer2_outputs(9918));
    outputs(10023) <= not(layer2_outputs(9086));
    outputs(10024) <= not(layer2_outputs(4418));
    outputs(10025) <= not(layer2_outputs(11789));
    outputs(10026) <= not((layer2_outputs(9323)) xor (layer2_outputs(6462)));
    outputs(10027) <= (layer2_outputs(9989)) xor (layer2_outputs(6550));
    outputs(10028) <= not(layer2_outputs(2935));
    outputs(10029) <= (layer2_outputs(4385)) and not (layer2_outputs(4805));
    outputs(10030) <= (layer2_outputs(9001)) or (layer2_outputs(12229));
    outputs(10031) <= (layer2_outputs(8692)) xor (layer2_outputs(4344));
    outputs(10032) <= layer2_outputs(7830);
    outputs(10033) <= not(layer2_outputs(10249));
    outputs(10034) <= not(layer2_outputs(9188));
    outputs(10035) <= (layer2_outputs(5781)) xor (layer2_outputs(8689));
    outputs(10036) <= not((layer2_outputs(1987)) xor (layer2_outputs(2701)));
    outputs(10037) <= not(layer2_outputs(4267)) or (layer2_outputs(4255));
    outputs(10038) <= not((layer2_outputs(8593)) xor (layer2_outputs(2835)));
    outputs(10039) <= not(layer2_outputs(4656));
    outputs(10040) <= not(layer2_outputs(2723));
    outputs(10041) <= not(layer2_outputs(5088));
    outputs(10042) <= layer2_outputs(11083);
    outputs(10043) <= layer2_outputs(9164);
    outputs(10044) <= not((layer2_outputs(12334)) xor (layer2_outputs(6159)));
    outputs(10045) <= not((layer2_outputs(2618)) xor (layer2_outputs(9799)));
    outputs(10046) <= not((layer2_outputs(12076)) xor (layer2_outputs(2740)));
    outputs(10047) <= not((layer2_outputs(6868)) or (layer2_outputs(6813)));
    outputs(10048) <= not(layer2_outputs(3416));
    outputs(10049) <= not((layer2_outputs(11582)) xor (layer2_outputs(466)));
    outputs(10050) <= not(layer2_outputs(87));
    outputs(10051) <= layer2_outputs(6254);
    outputs(10052) <= layer2_outputs(1205);
    outputs(10053) <= layer2_outputs(8653);
    outputs(10054) <= (layer2_outputs(12538)) xor (layer2_outputs(8225));
    outputs(10055) <= (layer2_outputs(6906)) and not (layer2_outputs(10459));
    outputs(10056) <= layer2_outputs(7757);
    outputs(10057) <= layer2_outputs(3915);
    outputs(10058) <= not(layer2_outputs(4527));
    outputs(10059) <= layer2_outputs(572);
    outputs(10060) <= (layer2_outputs(292)) and not (layer2_outputs(10177));
    outputs(10061) <= not(layer2_outputs(5743));
    outputs(10062) <= layer2_outputs(6434);
    outputs(10063) <= (layer2_outputs(8150)) and not (layer2_outputs(6600));
    outputs(10064) <= not((layer2_outputs(1696)) or (layer2_outputs(10435)));
    outputs(10065) <= not((layer2_outputs(11374)) and (layer2_outputs(750)));
    outputs(10066) <= not(layer2_outputs(6839)) or (layer2_outputs(1111));
    outputs(10067) <= (layer2_outputs(5272)) xor (layer2_outputs(6433));
    outputs(10068) <= layer2_outputs(424);
    outputs(10069) <= layer2_outputs(10035);
    outputs(10070) <= not((layer2_outputs(7603)) or (layer2_outputs(11492)));
    outputs(10071) <= layer2_outputs(791);
    outputs(10072) <= layer2_outputs(4369);
    outputs(10073) <= not(layer2_outputs(5445));
    outputs(10074) <= not(layer2_outputs(4712));
    outputs(10075) <= layer2_outputs(4788);
    outputs(10076) <= (layer2_outputs(1465)) and (layer2_outputs(9204));
    outputs(10077) <= not(layer2_outputs(9652));
    outputs(10078) <= not((layer2_outputs(1289)) xor (layer2_outputs(5223)));
    outputs(10079) <= layer2_outputs(4197);
    outputs(10080) <= not(layer2_outputs(6519));
    outputs(10081) <= layer2_outputs(9245);
    outputs(10082) <= layer2_outputs(8439);
    outputs(10083) <= layer2_outputs(12101);
    outputs(10084) <= layer2_outputs(4041);
    outputs(10085) <= not(layer2_outputs(9548));
    outputs(10086) <= (layer2_outputs(12523)) and not (layer2_outputs(119));
    outputs(10087) <= not((layer2_outputs(2534)) xor (layer2_outputs(11580)));
    outputs(10088) <= not(layer2_outputs(8325));
    outputs(10089) <= (layer2_outputs(9685)) xor (layer2_outputs(6130));
    outputs(10090) <= layer2_outputs(6311);
    outputs(10091) <= (layer2_outputs(8521)) and not (layer2_outputs(5311));
    outputs(10092) <= not((layer2_outputs(10126)) xor (layer2_outputs(8247)));
    outputs(10093) <= (layer2_outputs(290)) xor (layer2_outputs(357));
    outputs(10094) <= not(layer2_outputs(1530));
    outputs(10095) <= not(layer2_outputs(10702));
    outputs(10096) <= not(layer2_outputs(6905));
    outputs(10097) <= (layer2_outputs(9448)) xor (layer2_outputs(1749));
    outputs(10098) <= not(layer2_outputs(5389));
    outputs(10099) <= layer2_outputs(10645);
    outputs(10100) <= not((layer2_outputs(3953)) xor (layer2_outputs(1910)));
    outputs(10101) <= not(layer2_outputs(1381));
    outputs(10102) <= not(layer2_outputs(5593));
    outputs(10103) <= (layer2_outputs(12517)) and not (layer2_outputs(8152));
    outputs(10104) <= layer2_outputs(1097);
    outputs(10105) <= layer2_outputs(12140);
    outputs(10106) <= not(layer2_outputs(9271)) or (layer2_outputs(4618));
    outputs(10107) <= (layer2_outputs(7584)) and (layer2_outputs(10354));
    outputs(10108) <= layer2_outputs(9342);
    outputs(10109) <= layer2_outputs(2937);
    outputs(10110) <= (layer2_outputs(7680)) xor (layer2_outputs(10333));
    outputs(10111) <= not(layer2_outputs(1531));
    outputs(10112) <= layer2_outputs(4009);
    outputs(10113) <= not(layer2_outputs(5387));
    outputs(10114) <= not(layer2_outputs(5549));
    outputs(10115) <= not(layer2_outputs(9573));
    outputs(10116) <= not(layer2_outputs(7387));
    outputs(10117) <= not(layer2_outputs(10198));
    outputs(10118) <= layer2_outputs(11774);
    outputs(10119) <= layer2_outputs(7998);
    outputs(10120) <= layer2_outputs(6066);
    outputs(10121) <= (layer2_outputs(5303)) and not (layer2_outputs(6582));
    outputs(10122) <= not(layer2_outputs(5128));
    outputs(10123) <= (layer2_outputs(8801)) or (layer2_outputs(9477));
    outputs(10124) <= not((layer2_outputs(8246)) and (layer2_outputs(12591)));
    outputs(10125) <= layer2_outputs(9324);
    outputs(10126) <= (layer2_outputs(3214)) xor (layer2_outputs(9734));
    outputs(10127) <= layer2_outputs(642);
    outputs(10128) <= not((layer2_outputs(1774)) xor (layer2_outputs(10502)));
    outputs(10129) <= not(layer2_outputs(12335));
    outputs(10130) <= not(layer2_outputs(6026));
    outputs(10131) <= not((layer2_outputs(9867)) or (layer2_outputs(3)));
    outputs(10132) <= (layer2_outputs(2363)) and not (layer2_outputs(1365));
    outputs(10133) <= (layer2_outputs(8127)) xor (layer2_outputs(1423));
    outputs(10134) <= layer2_outputs(5641);
    outputs(10135) <= not(layer2_outputs(10625)) or (layer2_outputs(11519));
    outputs(10136) <= (layer2_outputs(10573)) xor (layer2_outputs(11219));
    outputs(10137) <= (layer2_outputs(10544)) xor (layer2_outputs(10016));
    outputs(10138) <= not(layer2_outputs(5908));
    outputs(10139) <= layer2_outputs(8440);
    outputs(10140) <= not(layer2_outputs(12290));
    outputs(10141) <= not((layer2_outputs(10914)) xor (layer2_outputs(1775)));
    outputs(10142) <= not(layer2_outputs(460));
    outputs(10143) <= layer2_outputs(11207);
    outputs(10144) <= (layer2_outputs(9939)) xor (layer2_outputs(1789));
    outputs(10145) <= not(layer2_outputs(8884));
    outputs(10146) <= (layer2_outputs(8544)) xor (layer2_outputs(12071));
    outputs(10147) <= (layer2_outputs(10620)) and not (layer2_outputs(528));
    outputs(10148) <= not(layer2_outputs(4501)) or (layer2_outputs(331));
    outputs(10149) <= not(layer2_outputs(11824));
    outputs(10150) <= not((layer2_outputs(11496)) xor (layer2_outputs(7088)));
    outputs(10151) <= layer2_outputs(2511);
    outputs(10152) <= layer2_outputs(2833);
    outputs(10153) <= not(layer2_outputs(941));
    outputs(10154) <= not(layer2_outputs(8724));
    outputs(10155) <= (layer2_outputs(2787)) xor (layer2_outputs(9641));
    outputs(10156) <= not((layer2_outputs(9037)) xor (layer2_outputs(7565)));
    outputs(10157) <= not((layer2_outputs(9415)) xor (layer2_outputs(9783)));
    outputs(10158) <= not((layer2_outputs(3623)) xor (layer2_outputs(4834)));
    outputs(10159) <= not((layer2_outputs(4928)) and (layer2_outputs(7717)));
    outputs(10160) <= layer2_outputs(4385);
    outputs(10161) <= (layer2_outputs(3802)) and (layer2_outputs(5542));
    outputs(10162) <= layer2_outputs(11631);
    outputs(10163) <= not(layer2_outputs(9561));
    outputs(10164) <= not((layer2_outputs(5167)) xor (layer2_outputs(10294)));
    outputs(10165) <= not((layer2_outputs(1665)) or (layer2_outputs(6323)));
    outputs(10166) <= layer2_outputs(1227);
    outputs(10167) <= (layer2_outputs(11957)) and (layer2_outputs(469));
    outputs(10168) <= not(layer2_outputs(5981));
    outputs(10169) <= not((layer2_outputs(1922)) xor (layer2_outputs(3300)));
    outputs(10170) <= (layer2_outputs(5903)) xor (layer2_outputs(2097));
    outputs(10171) <= not(layer2_outputs(7598));
    outputs(10172) <= layer2_outputs(4488);
    outputs(10173) <= layer2_outputs(3533);
    outputs(10174) <= layer2_outputs(1095);
    outputs(10175) <= layer2_outputs(6602);
    outputs(10176) <= not(layer2_outputs(151));
    outputs(10177) <= layer2_outputs(3973);
    outputs(10178) <= not((layer2_outputs(1277)) or (layer2_outputs(9015)));
    outputs(10179) <= (layer2_outputs(1916)) and (layer2_outputs(5711));
    outputs(10180) <= not(layer2_outputs(3410)) or (layer2_outputs(4636));
    outputs(10181) <= layer2_outputs(12718);
    outputs(10182) <= layer2_outputs(8159);
    outputs(10183) <= not((layer2_outputs(10973)) xor (layer2_outputs(8536)));
    outputs(10184) <= layer2_outputs(7024);
    outputs(10185) <= not(layer2_outputs(1578));
    outputs(10186) <= not(layer2_outputs(4389));
    outputs(10187) <= layer2_outputs(1169);
    outputs(10188) <= layer2_outputs(1227);
    outputs(10189) <= layer2_outputs(11330);
    outputs(10190) <= layer2_outputs(4208);
    outputs(10191) <= layer2_outputs(9769);
    outputs(10192) <= layer2_outputs(11798);
    outputs(10193) <= layer2_outputs(8414);
    outputs(10194) <= not(layer2_outputs(12622));
    outputs(10195) <= not(layer2_outputs(2031));
    outputs(10196) <= not((layer2_outputs(10490)) or (layer2_outputs(6607)));
    outputs(10197) <= not(layer2_outputs(2771));
    outputs(10198) <= not((layer2_outputs(9928)) xor (layer2_outputs(8690)));
    outputs(10199) <= not(layer2_outputs(1614));
    outputs(10200) <= not(layer2_outputs(9433));
    outputs(10201) <= (layer2_outputs(12409)) xor (layer2_outputs(12687));
    outputs(10202) <= layer2_outputs(3637);
    outputs(10203) <= layer2_outputs(2836);
    outputs(10204) <= not(layer2_outputs(2539)) or (layer2_outputs(2348));
    outputs(10205) <= layer2_outputs(9246);
    outputs(10206) <= not(layer2_outputs(763));
    outputs(10207) <= not(layer2_outputs(9338));
    outputs(10208) <= layer2_outputs(7564);
    outputs(10209) <= (layer2_outputs(10442)) and not (layer2_outputs(7701));
    outputs(10210) <= (layer2_outputs(11897)) or (layer2_outputs(2448));
    outputs(10211) <= layer2_outputs(8726);
    outputs(10212) <= not(layer2_outputs(5740));
    outputs(10213) <= layer2_outputs(8363);
    outputs(10214) <= layer2_outputs(2477);
    outputs(10215) <= not((layer2_outputs(11358)) or (layer2_outputs(8221)));
    outputs(10216) <= (layer2_outputs(8593)) xor (layer2_outputs(9023));
    outputs(10217) <= (layer2_outputs(10356)) and (layer2_outputs(11398));
    outputs(10218) <= (layer2_outputs(9743)) and not (layer2_outputs(1685));
    outputs(10219) <= not(layer2_outputs(314));
    outputs(10220) <= not(layer2_outputs(2117));
    outputs(10221) <= not(layer2_outputs(3874));
    outputs(10222) <= (layer2_outputs(10390)) and not (layer2_outputs(7423));
    outputs(10223) <= not(layer2_outputs(8583));
    outputs(10224) <= not((layer2_outputs(8781)) xor (layer2_outputs(6855)));
    outputs(10225) <= (layer2_outputs(1105)) xor (layer2_outputs(3406));
    outputs(10226) <= (layer2_outputs(3794)) xor (layer2_outputs(2388));
    outputs(10227) <= not((layer2_outputs(6244)) xor (layer2_outputs(5979)));
    outputs(10228) <= layer2_outputs(7062);
    outputs(10229) <= layer2_outputs(81);
    outputs(10230) <= not(layer2_outputs(5353));
    outputs(10231) <= not(layer2_outputs(3642));
    outputs(10232) <= (layer2_outputs(902)) xor (layer2_outputs(1395));
    outputs(10233) <= layer2_outputs(8082);
    outputs(10234) <= not(layer2_outputs(2911));
    outputs(10235) <= not((layer2_outputs(4176)) xor (layer2_outputs(7743)));
    outputs(10236) <= layer2_outputs(5070);
    outputs(10237) <= not(layer2_outputs(3198));
    outputs(10238) <= (layer2_outputs(11575)) xor (layer2_outputs(793));
    outputs(10239) <= not(layer2_outputs(4129));
    outputs(10240) <= layer2_outputs(9755);
    outputs(10241) <= (layer2_outputs(6815)) or (layer2_outputs(10147));
    outputs(10242) <= layer2_outputs(10117);
    outputs(10243) <= not((layer2_outputs(11370)) xor (layer2_outputs(11391)));
    outputs(10244) <= layer2_outputs(10540);
    outputs(10245) <= layer2_outputs(10614);
    outputs(10246) <= not(layer2_outputs(7147));
    outputs(10247) <= not(layer2_outputs(4701)) or (layer2_outputs(10353));
    outputs(10248) <= not(layer2_outputs(11030));
    outputs(10249) <= (layer2_outputs(4163)) and (layer2_outputs(9006));
    outputs(10250) <= not(layer2_outputs(682));
    outputs(10251) <= (layer2_outputs(3700)) xor (layer2_outputs(12230));
    outputs(10252) <= layer2_outputs(522);
    outputs(10253) <= not(layer2_outputs(12239)) or (layer2_outputs(10725));
    outputs(10254) <= not((layer2_outputs(1404)) xor (layer2_outputs(6135)));
    outputs(10255) <= not(layer2_outputs(6769));
    outputs(10256) <= (layer2_outputs(10819)) xor (layer2_outputs(1700));
    outputs(10257) <= not((layer2_outputs(3911)) xor (layer2_outputs(3098)));
    outputs(10258) <= not(layer2_outputs(1353));
    outputs(10259) <= not(layer2_outputs(8658));
    outputs(10260) <= (layer2_outputs(6506)) xor (layer2_outputs(6770));
    outputs(10261) <= (layer2_outputs(1609)) xor (layer2_outputs(3364));
    outputs(10262) <= layer2_outputs(8992);
    outputs(10263) <= (layer2_outputs(947)) or (layer2_outputs(1309));
    outputs(10264) <= (layer2_outputs(9682)) xor (layer2_outputs(2058));
    outputs(10265) <= not(layer2_outputs(1005));
    outputs(10266) <= layer2_outputs(11243);
    outputs(10267) <= layer2_outputs(4153);
    outputs(10268) <= not(layer2_outputs(4456));
    outputs(10269) <= not(layer2_outputs(1568));
    outputs(10270) <= (layer2_outputs(3857)) and (layer2_outputs(7095));
    outputs(10271) <= layer2_outputs(12314);
    outputs(10272) <= not(layer2_outputs(5080)) or (layer2_outputs(10631));
    outputs(10273) <= not(layer2_outputs(3694)) or (layer2_outputs(527));
    outputs(10274) <= (layer2_outputs(9570)) xor (layer2_outputs(9811));
    outputs(10275) <= (layer2_outputs(2362)) xor (layer2_outputs(4584));
    outputs(10276) <= layer2_outputs(9223);
    outputs(10277) <= not(layer2_outputs(7690));
    outputs(10278) <= (layer2_outputs(4889)) xor (layer2_outputs(12793));
    outputs(10279) <= not((layer2_outputs(487)) xor (layer2_outputs(8606)));
    outputs(10280) <= layer2_outputs(10374);
    outputs(10281) <= not(layer2_outputs(3191));
    outputs(10282) <= not((layer2_outputs(12129)) xor (layer2_outputs(4488)));
    outputs(10283) <= not(layer2_outputs(11177));
    outputs(10284) <= layer2_outputs(9187);
    outputs(10285) <= (layer2_outputs(2949)) and not (layer2_outputs(8964));
    outputs(10286) <= not((layer2_outputs(377)) xor (layer2_outputs(2178)));
    outputs(10287) <= not(layer2_outputs(3737));
    outputs(10288) <= (layer2_outputs(5716)) xor (layer2_outputs(2100));
    outputs(10289) <= not(layer2_outputs(4606));
    outputs(10290) <= layer2_outputs(7507);
    outputs(10291) <= layer2_outputs(3248);
    outputs(10292) <= layer2_outputs(11001);
    outputs(10293) <= not((layer2_outputs(10305)) xor (layer2_outputs(10509)));
    outputs(10294) <= (layer2_outputs(9292)) xor (layer2_outputs(12116));
    outputs(10295) <= (layer2_outputs(3340)) xor (layer2_outputs(8655));
    outputs(10296) <= (layer2_outputs(4422)) xor (layer2_outputs(7228));
    outputs(10297) <= layer2_outputs(12625);
    outputs(10298) <= not(layer2_outputs(11553));
    outputs(10299) <= layer2_outputs(1779);
    outputs(10300) <= not((layer2_outputs(12345)) xor (layer2_outputs(8792)));
    outputs(10301) <= layer2_outputs(5817);
    outputs(10302) <= layer2_outputs(6283);
    outputs(10303) <= not(layer2_outputs(1014));
    outputs(10304) <= not(layer2_outputs(9845));
    outputs(10305) <= not(layer2_outputs(7419));
    outputs(10306) <= (layer2_outputs(11604)) xor (layer2_outputs(1132));
    outputs(10307) <= not(layer2_outputs(5535));
    outputs(10308) <= layer2_outputs(12788);
    outputs(10309) <= not((layer2_outputs(168)) xor (layer2_outputs(10303)));
    outputs(10310) <= not(layer2_outputs(3147));
    outputs(10311) <= not(layer2_outputs(5836));
    outputs(10312) <= layer2_outputs(9747);
    outputs(10313) <= layer2_outputs(195);
    outputs(10314) <= not(layer2_outputs(5362));
    outputs(10315) <= not(layer2_outputs(5131));
    outputs(10316) <= not(layer2_outputs(10255));
    outputs(10317) <= layer2_outputs(12215);
    outputs(10318) <= not((layer2_outputs(4862)) or (layer2_outputs(4696)));
    outputs(10319) <= layer2_outputs(1436);
    outputs(10320) <= (layer2_outputs(10449)) or (layer2_outputs(434));
    outputs(10321) <= not(layer2_outputs(8964)) or (layer2_outputs(5400));
    outputs(10322) <= not((layer2_outputs(8064)) xor (layer2_outputs(1951)));
    outputs(10323) <= not(layer2_outputs(919));
    outputs(10324) <= (layer2_outputs(6044)) xor (layer2_outputs(11319));
    outputs(10325) <= not((layer2_outputs(11772)) xor (layer2_outputs(10854)));
    outputs(10326) <= not((layer2_outputs(8109)) xor (layer2_outputs(1496)));
    outputs(10327) <= not((layer2_outputs(12432)) xor (layer2_outputs(7233)));
    outputs(10328) <= (layer2_outputs(8128)) xor (layer2_outputs(9243));
    outputs(10329) <= not(layer2_outputs(2433)) or (layer2_outputs(6120));
    outputs(10330) <= (layer2_outputs(12601)) xor (layer2_outputs(5088));
    outputs(10331) <= not(layer2_outputs(8708));
    outputs(10332) <= not(layer2_outputs(8631)) or (layer2_outputs(468));
    outputs(10333) <= (layer2_outputs(4352)) xor (layer2_outputs(10243));
    outputs(10334) <= layer2_outputs(6359);
    outputs(10335) <= layer2_outputs(12728);
    outputs(10336) <= not((layer2_outputs(3465)) xor (layer2_outputs(10411)));
    outputs(10337) <= (layer2_outputs(173)) and not (layer2_outputs(9447));
    outputs(10338) <= (layer2_outputs(1836)) xor (layer2_outputs(5287));
    outputs(10339) <= layer2_outputs(10351);
    outputs(10340) <= not(layer2_outputs(11293));
    outputs(10341) <= layer2_outputs(1669);
    outputs(10342) <= not(layer2_outputs(11690)) or (layer2_outputs(5976));
    outputs(10343) <= not(layer2_outputs(6313));
    outputs(10344) <= layer2_outputs(2008);
    outputs(10345) <= not(layer2_outputs(10511));
    outputs(10346) <= layer2_outputs(4128);
    outputs(10347) <= not((layer2_outputs(1326)) xor (layer2_outputs(4471)));
    outputs(10348) <= not(layer2_outputs(5138));
    outputs(10349) <= (layer2_outputs(10245)) xor (layer2_outputs(9146));
    outputs(10350) <= not((layer2_outputs(3044)) and (layer2_outputs(7903)));
    outputs(10351) <= not((layer2_outputs(8744)) xor (layer2_outputs(12366)));
    outputs(10352) <= not(layer2_outputs(8438));
    outputs(10353) <= not(layer2_outputs(6585)) or (layer2_outputs(10898));
    outputs(10354) <= not(layer2_outputs(10313)) or (layer2_outputs(686));
    outputs(10355) <= not(layer2_outputs(5481));
    outputs(10356) <= not((layer2_outputs(4892)) xor (layer2_outputs(10628)));
    outputs(10357) <= not(layer2_outputs(4645));
    outputs(10358) <= layer2_outputs(9550);
    outputs(10359) <= layer2_outputs(12193);
    outputs(10360) <= not((layer2_outputs(1348)) xor (layer2_outputs(2008)));
    outputs(10361) <= not(layer2_outputs(4331));
    outputs(10362) <= not(layer2_outputs(6954));
    outputs(10363) <= layer2_outputs(2748);
    outputs(10364) <= not(layer2_outputs(2109));
    outputs(10365) <= (layer2_outputs(8634)) xor (layer2_outputs(11352));
    outputs(10366) <= layer2_outputs(8552);
    outputs(10367) <= layer2_outputs(280);
    outputs(10368) <= not((layer2_outputs(4022)) xor (layer2_outputs(10417)));
    outputs(10369) <= not(layer2_outputs(9134)) or (layer2_outputs(4634));
    outputs(10370) <= (layer2_outputs(8461)) xor (layer2_outputs(3299));
    outputs(10371) <= (layer2_outputs(9123)) xor (layer2_outputs(7214));
    outputs(10372) <= layer2_outputs(4442);
    outputs(10373) <= layer2_outputs(2196);
    outputs(10374) <= not(layer2_outputs(11681));
    outputs(10375) <= not(layer2_outputs(3066)) or (layer2_outputs(10776));
    outputs(10376) <= not(layer2_outputs(2904));
    outputs(10377) <= layer2_outputs(11877);
    outputs(10378) <= not((layer2_outputs(9433)) xor (layer2_outputs(10790)));
    outputs(10379) <= layer2_outputs(4277);
    outputs(10380) <= not(layer2_outputs(12065));
    outputs(10381) <= not(layer2_outputs(7966));
    outputs(10382) <= (layer2_outputs(7176)) xor (layer2_outputs(11504));
    outputs(10383) <= not((layer2_outputs(5301)) or (layer2_outputs(5875)));
    outputs(10384) <= not(layer2_outputs(6525));
    outputs(10385) <= layer2_outputs(8901);
    outputs(10386) <= not((layer2_outputs(9143)) xor (layer2_outputs(6699)));
    outputs(10387) <= not((layer2_outputs(4734)) xor (layer2_outputs(210)));
    outputs(10388) <= (layer2_outputs(2549)) xor (layer2_outputs(1827));
    outputs(10389) <= not(layer2_outputs(9214)) or (layer2_outputs(10510));
    outputs(10390) <= (layer2_outputs(4659)) and not (layer2_outputs(11551));
    outputs(10391) <= not(layer2_outputs(433));
    outputs(10392) <= (layer2_outputs(2030)) xor (layer2_outputs(2772));
    outputs(10393) <= (layer2_outputs(1389)) and not (layer2_outputs(1284));
    outputs(10394) <= layer2_outputs(9228);
    outputs(10395) <= not((layer2_outputs(10179)) xor (layer2_outputs(9445)));
    outputs(10396) <= not(layer2_outputs(1155));
    outputs(10397) <= not((layer2_outputs(6117)) or (layer2_outputs(8522)));
    outputs(10398) <= not(layer2_outputs(4468)) or (layer2_outputs(5724));
    outputs(10399) <= not(layer2_outputs(8515));
    outputs(10400) <= not(layer2_outputs(6422));
    outputs(10401) <= layer2_outputs(6076);
    outputs(10402) <= (layer2_outputs(12735)) or (layer2_outputs(3034));
    outputs(10403) <= not(layer2_outputs(6004)) or (layer2_outputs(12034));
    outputs(10404) <= (layer2_outputs(10281)) or (layer2_outputs(12575));
    outputs(10405) <= layer2_outputs(6229);
    outputs(10406) <= not(layer2_outputs(585));
    outputs(10407) <= (layer2_outputs(4189)) and (layer2_outputs(9854));
    outputs(10408) <= not((layer2_outputs(10194)) xor (layer2_outputs(7406)));
    outputs(10409) <= not(layer2_outputs(1963));
    outputs(10410) <= not(layer2_outputs(6846));
    outputs(10411) <= not(layer2_outputs(10149)) or (layer2_outputs(10607));
    outputs(10412) <= (layer2_outputs(8340)) xor (layer2_outputs(3329));
    outputs(10413) <= layer2_outputs(10056);
    outputs(10414) <= layer2_outputs(2640);
    outputs(10415) <= (layer2_outputs(7657)) xor (layer2_outputs(2817));
    outputs(10416) <= (layer2_outputs(1656)) or (layer2_outputs(4908));
    outputs(10417) <= not((layer2_outputs(12709)) xor (layer2_outputs(11407)));
    outputs(10418) <= not(layer2_outputs(8797)) or (layer2_outputs(12601));
    outputs(10419) <= not(layer2_outputs(12433));
    outputs(10420) <= not(layer2_outputs(10709));
    outputs(10421) <= layer2_outputs(1547);
    outputs(10422) <= not(layer2_outputs(1118)) or (layer2_outputs(7208));
    outputs(10423) <= not((layer2_outputs(4158)) xor (layer2_outputs(8031)));
    outputs(10424) <= (layer2_outputs(462)) xor (layer2_outputs(8559));
    outputs(10425) <= layer2_outputs(3316);
    outputs(10426) <= (layer2_outputs(4922)) or (layer2_outputs(6929));
    outputs(10427) <= layer2_outputs(7085);
    outputs(10428) <= layer2_outputs(3981);
    outputs(10429) <= layer2_outputs(10508);
    outputs(10430) <= (layer2_outputs(12441)) xor (layer2_outputs(10214));
    outputs(10431) <= not((layer2_outputs(12557)) xor (layer2_outputs(11337)));
    outputs(10432) <= (layer2_outputs(9089)) or (layer2_outputs(10850));
    outputs(10433) <= not(layer2_outputs(5050));
    outputs(10434) <= (layer2_outputs(7730)) xor (layer2_outputs(753));
    outputs(10435) <= layer2_outputs(1710);
    outputs(10436) <= not(layer2_outputs(9008)) or (layer2_outputs(1329));
    outputs(10437) <= not(layer2_outputs(177));
    outputs(10438) <= layer2_outputs(6258);
    outputs(10439) <= (layer2_outputs(9328)) xor (layer2_outputs(6740));
    outputs(10440) <= (layer2_outputs(1999)) xor (layer2_outputs(12778));
    outputs(10441) <= (layer2_outputs(3825)) xor (layer2_outputs(2999));
    outputs(10442) <= not((layer2_outputs(8277)) xor (layer2_outputs(960)));
    outputs(10443) <= (layer2_outputs(8561)) xor (layer2_outputs(3926));
    outputs(10444) <= (layer2_outputs(1980)) xor (layer2_outputs(4008));
    outputs(10445) <= not((layer2_outputs(2868)) xor (layer2_outputs(5051)));
    outputs(10446) <= layer2_outputs(13);
    outputs(10447) <= not(layer2_outputs(8874)) or (layer2_outputs(5285));
    outputs(10448) <= not(layer2_outputs(11883)) or (layer2_outputs(597));
    outputs(10449) <= (layer2_outputs(4733)) xor (layer2_outputs(10275));
    outputs(10450) <= (layer2_outputs(4408)) xor (layer2_outputs(1765));
    outputs(10451) <= (layer2_outputs(3811)) xor (layer2_outputs(4142));
    outputs(10452) <= not(layer2_outputs(12283)) or (layer2_outputs(6061));
    outputs(10453) <= (layer2_outputs(11449)) and not (layer2_outputs(8513));
    outputs(10454) <= (layer2_outputs(4290)) xor (layer2_outputs(8028));
    outputs(10455) <= (layer2_outputs(11387)) xor (layer2_outputs(7931));
    outputs(10456) <= not(layer2_outputs(6474));
    outputs(10457) <= not((layer2_outputs(7732)) xor (layer2_outputs(10083)));
    outputs(10458) <= layer2_outputs(9250);
    outputs(10459) <= layer2_outputs(510);
    outputs(10460) <= not((layer2_outputs(3983)) xor (layer2_outputs(11497)));
    outputs(10461) <= layer2_outputs(9871);
    outputs(10462) <= (layer2_outputs(3874)) xor (layer2_outputs(8012));
    outputs(10463) <= not(layer2_outputs(9751)) or (layer2_outputs(2990));
    outputs(10464) <= not((layer2_outputs(3046)) xor (layer2_outputs(1777)));
    outputs(10465) <= (layer2_outputs(3940)) xor (layer2_outputs(873));
    outputs(10466) <= not(layer2_outputs(8164));
    outputs(10467) <= (layer2_outputs(7743)) xor (layer2_outputs(10085));
    outputs(10468) <= not(layer2_outputs(11682));
    outputs(10469) <= (layer2_outputs(238)) and not (layer2_outputs(1026));
    outputs(10470) <= layer2_outputs(2604);
    outputs(10471) <= not(layer2_outputs(6006)) or (layer2_outputs(7348));
    outputs(10472) <= layer2_outputs(11803);
    outputs(10473) <= (layer2_outputs(3914)) xor (layer2_outputs(10512));
    outputs(10474) <= layer2_outputs(10576);
    outputs(10475) <= (layer2_outputs(2276)) xor (layer2_outputs(2592));
    outputs(10476) <= not((layer2_outputs(4634)) xor (layer2_outputs(11323)));
    outputs(10477) <= not((layer2_outputs(7051)) and (layer2_outputs(11845)));
    outputs(10478) <= layer2_outputs(11487);
    outputs(10479) <= layer2_outputs(5713);
    outputs(10480) <= (layer2_outputs(1163)) xor (layer2_outputs(10281));
    outputs(10481) <= layer2_outputs(477);
    outputs(10482) <= layer2_outputs(9031);
    outputs(10483) <= not(layer2_outputs(7961)) or (layer2_outputs(7110));
    outputs(10484) <= layer2_outputs(1557);
    outputs(10485) <= not(layer2_outputs(1008));
    outputs(10486) <= not(layer2_outputs(9199));
    outputs(10487) <= not((layer2_outputs(12214)) xor (layer2_outputs(3142)));
    outputs(10488) <= layer2_outputs(2900);
    outputs(10489) <= not(layer2_outputs(2536));
    outputs(10490) <= (layer2_outputs(1114)) xor (layer2_outputs(12251));
    outputs(10491) <= (layer2_outputs(4809)) xor (layer2_outputs(8436));
    outputs(10492) <= not((layer2_outputs(3820)) and (layer2_outputs(2993)));
    outputs(10493) <= not((layer2_outputs(744)) xor (layer2_outputs(2584)));
    outputs(10494) <= layer2_outputs(12299);
    outputs(10495) <= not((layer2_outputs(11539)) xor (layer2_outputs(6515)));
    outputs(10496) <= not((layer2_outputs(113)) xor (layer2_outputs(6552)));
    outputs(10497) <= (layer2_outputs(5577)) and not (layer2_outputs(7558));
    outputs(10498) <= (layer2_outputs(2646)) or (layer2_outputs(3053));
    outputs(10499) <= layer2_outputs(2335);
    outputs(10500) <= not(layer2_outputs(8285));
    outputs(10501) <= layer2_outputs(10239);
    outputs(10502) <= not(layer2_outputs(8602));
    outputs(10503) <= layer2_outputs(11674);
    outputs(10504) <= not((layer2_outputs(7431)) xor (layer2_outputs(11182)));
    outputs(10505) <= not((layer2_outputs(8520)) and (layer2_outputs(9555)));
    outputs(10506) <= not((layer2_outputs(8296)) xor (layer2_outputs(2099)));
    outputs(10507) <= not(layer2_outputs(8479));
    outputs(10508) <= not((layer2_outputs(6993)) xor (layer2_outputs(8472)));
    outputs(10509) <= layer2_outputs(2886);
    outputs(10510) <= not(layer2_outputs(7535));
    outputs(10511) <= not(layer2_outputs(2083));
    outputs(10512) <= not(layer2_outputs(3988)) or (layer2_outputs(9691));
    outputs(10513) <= layer2_outputs(5448);
    outputs(10514) <= (layer2_outputs(8199)) xor (layer2_outputs(2603));
    outputs(10515) <= not((layer2_outputs(5446)) xor (layer2_outputs(5752)));
    outputs(10516) <= not((layer2_outputs(3463)) and (layer2_outputs(6198)));
    outputs(10517) <= layer2_outputs(10115);
    outputs(10518) <= (layer2_outputs(1348)) xor (layer2_outputs(6046));
    outputs(10519) <= not(layer2_outputs(4236)) or (layer2_outputs(10557));
    outputs(10520) <= not(layer2_outputs(2090));
    outputs(10521) <= (layer2_outputs(8760)) xor (layer2_outputs(11719));
    outputs(10522) <= (layer2_outputs(11831)) xor (layer2_outputs(4119));
    outputs(10523) <= layer2_outputs(11859);
    outputs(10524) <= layer2_outputs(2914);
    outputs(10525) <= layer2_outputs(4559);
    outputs(10526) <= not(layer2_outputs(4170));
    outputs(10527) <= not((layer2_outputs(8549)) xor (layer2_outputs(4145)));
    outputs(10528) <= (layer2_outputs(5141)) xor (layer2_outputs(10137));
    outputs(10529) <= not(layer2_outputs(11392));
    outputs(10530) <= not(layer2_outputs(3302));
    outputs(10531) <= (layer2_outputs(4438)) xor (layer2_outputs(4505));
    outputs(10532) <= not(layer2_outputs(10406));
    outputs(10533) <= layer2_outputs(565);
    outputs(10534) <= layer2_outputs(9755);
    outputs(10535) <= not(layer2_outputs(4870));
    outputs(10536) <= not(layer2_outputs(11891));
    outputs(10537) <= not(layer2_outputs(4209));
    outputs(10538) <= not(layer2_outputs(536));
    outputs(10539) <= not(layer2_outputs(4216));
    outputs(10540) <= layer2_outputs(9088);
    outputs(10541) <= not(layer2_outputs(11878));
    outputs(10542) <= not(layer2_outputs(12049)) or (layer2_outputs(2092));
    outputs(10543) <= not(layer2_outputs(9891));
    outputs(10544) <= not((layer2_outputs(6304)) xor (layer2_outputs(3042)));
    outputs(10545) <= not((layer2_outputs(8096)) xor (layer2_outputs(4467)));
    outputs(10546) <= (layer2_outputs(6485)) xor (layer2_outputs(7036));
    outputs(10547) <= not(layer2_outputs(5135)) or (layer2_outputs(7138));
    outputs(10548) <= layer2_outputs(4973);
    outputs(10549) <= not((layer2_outputs(12451)) or (layer2_outputs(10669)));
    outputs(10550) <= not((layer2_outputs(1690)) and (layer2_outputs(5147)));
    outputs(10551) <= not((layer2_outputs(2208)) xor (layer2_outputs(3355)));
    outputs(10552) <= layer2_outputs(3111);
    outputs(10553) <= not(layer2_outputs(47));
    outputs(10554) <= not(layer2_outputs(3079));
    outputs(10555) <= not(layer2_outputs(4663));
    outputs(10556) <= not((layer2_outputs(11757)) xor (layer2_outputs(8101)));
    outputs(10557) <= (layer2_outputs(10537)) and (layer2_outputs(11748));
    outputs(10558) <= not(layer2_outputs(9151)) or (layer2_outputs(10941));
    outputs(10559) <= not((layer2_outputs(12264)) xor (layer2_outputs(214)));
    outputs(10560) <= (layer2_outputs(10825)) xor (layer2_outputs(6404));
    outputs(10561) <= layer2_outputs(6292);
    outputs(10562) <= not(layer2_outputs(6965));
    outputs(10563) <= layer2_outputs(9373);
    outputs(10564) <= (layer2_outputs(6884)) and (layer2_outputs(2546));
    outputs(10565) <= (layer2_outputs(2509)) xor (layer2_outputs(4106));
    outputs(10566) <= not((layer2_outputs(4610)) xor (layer2_outputs(3022)));
    outputs(10567) <= not((layer2_outputs(398)) and (layer2_outputs(8658)));
    outputs(10568) <= (layer2_outputs(7018)) xor (layer2_outputs(9322));
    outputs(10569) <= (layer2_outputs(11359)) and (layer2_outputs(9704));
    outputs(10570) <= not(layer2_outputs(3464));
    outputs(10571) <= not(layer2_outputs(9833));
    outputs(10572) <= not((layer2_outputs(11668)) xor (layer2_outputs(4701)));
    outputs(10573) <= layer2_outputs(6897);
    outputs(10574) <= not(layer2_outputs(9273));
    outputs(10575) <= not((layer2_outputs(7413)) xor (layer2_outputs(6343)));
    outputs(10576) <= (layer2_outputs(4152)) xor (layer2_outputs(8342));
    outputs(10577) <= not((layer2_outputs(1043)) xor (layer2_outputs(12757)));
    outputs(10578) <= not(layer2_outputs(2267));
    outputs(10579) <= not((layer2_outputs(8622)) xor (layer2_outputs(12411)));
    outputs(10580) <= not((layer2_outputs(1853)) xor (layer2_outputs(4336)));
    outputs(10581) <= not(layer2_outputs(6540));
    outputs(10582) <= not(layer2_outputs(11793));
    outputs(10583) <= (layer2_outputs(11582)) xor (layer2_outputs(997));
    outputs(10584) <= not((layer2_outputs(1931)) and (layer2_outputs(5079)));
    outputs(10585) <= layer2_outputs(365);
    outputs(10586) <= layer2_outputs(6274);
    outputs(10587) <= layer2_outputs(8793);
    outputs(10588) <= layer2_outputs(1989);
    outputs(10589) <= not((layer2_outputs(9374)) and (layer2_outputs(11699)));
    outputs(10590) <= not((layer2_outputs(4747)) xor (layer2_outputs(11006)));
    outputs(10591) <= not(layer2_outputs(5799)) or (layer2_outputs(7100));
    outputs(10592) <= not(layer2_outputs(9833));
    outputs(10593) <= layer2_outputs(8165);
    outputs(10594) <= layer2_outputs(317);
    outputs(10595) <= not(layer2_outputs(9493));
    outputs(10596) <= not(layer2_outputs(9607)) or (layer2_outputs(10019));
    outputs(10597) <= not((layer2_outputs(1267)) xor (layer2_outputs(3866)));
    outputs(10598) <= (layer2_outputs(11533)) xor (layer2_outputs(3346));
    outputs(10599) <= (layer2_outputs(2269)) and not (layer2_outputs(2561));
    outputs(10600) <= layer2_outputs(4931);
    outputs(10601) <= layer2_outputs(10434);
    outputs(10602) <= not((layer2_outputs(8939)) xor (layer2_outputs(5761)));
    outputs(10603) <= layer2_outputs(5401);
    outputs(10604) <= not((layer2_outputs(9445)) and (layer2_outputs(959)));
    outputs(10605) <= layer2_outputs(282);
    outputs(10606) <= not(layer2_outputs(2959)) or (layer2_outputs(10811));
    outputs(10607) <= (layer2_outputs(9379)) xor (layer2_outputs(12550));
    outputs(10608) <= (layer2_outputs(6492)) or (layer2_outputs(4255));
    outputs(10609) <= layer2_outputs(7462);
    outputs(10610) <= layer2_outputs(3722);
    outputs(10611) <= not((layer2_outputs(5066)) xor (layer2_outputs(9261)));
    outputs(10612) <= (layer2_outputs(7529)) xor (layer2_outputs(10572));
    outputs(10613) <= layer2_outputs(9591);
    outputs(10614) <= (layer2_outputs(4105)) xor (layer2_outputs(8956));
    outputs(10615) <= layer2_outputs(12729);
    outputs(10616) <= (layer2_outputs(11199)) xor (layer2_outputs(599));
    outputs(10617) <= not(layer2_outputs(6048)) or (layer2_outputs(1855));
    outputs(10618) <= (layer2_outputs(1709)) xor (layer2_outputs(12599));
    outputs(10619) <= (layer2_outputs(6992)) xor (layer2_outputs(1144));
    outputs(10620) <= layer2_outputs(8094);
    outputs(10621) <= layer2_outputs(1529);
    outputs(10622) <= (layer2_outputs(3242)) xor (layer2_outputs(8862));
    outputs(10623) <= layer2_outputs(4192);
    outputs(10624) <= not((layer2_outputs(981)) xor (layer2_outputs(11994)));
    outputs(10625) <= not(layer2_outputs(3046)) or (layer2_outputs(6075));
    outputs(10626) <= not((layer2_outputs(2866)) xor (layer2_outputs(9590)));
    outputs(10627) <= layer2_outputs(391);
    outputs(10628) <= (layer2_outputs(4322)) and not (layer2_outputs(4979));
    outputs(10629) <= not(layer2_outputs(5590));
    outputs(10630) <= (layer2_outputs(11225)) xor (layer2_outputs(11888));
    outputs(10631) <= not(layer2_outputs(2852));
    outputs(10632) <= (layer2_outputs(11099)) or (layer2_outputs(5731));
    outputs(10633) <= not((layer2_outputs(7017)) xor (layer2_outputs(5957)));
    outputs(10634) <= not((layer2_outputs(4901)) and (layer2_outputs(742)));
    outputs(10635) <= layer2_outputs(8860);
    outputs(10636) <= not((layer2_outputs(8292)) xor (layer2_outputs(6653)));
    outputs(10637) <= not(layer2_outputs(9185)) or (layer2_outputs(4551));
    outputs(10638) <= layer2_outputs(3613);
    outputs(10639) <= not(layer2_outputs(3622));
    outputs(10640) <= (layer2_outputs(3580)) and not (layer2_outputs(5239));
    outputs(10641) <= not((layer2_outputs(9702)) or (layer2_outputs(2730)));
    outputs(10642) <= not(layer2_outputs(10313)) or (layer2_outputs(9109));
    outputs(10643) <= (layer2_outputs(12635)) xor (layer2_outputs(5019));
    outputs(10644) <= layer2_outputs(1174);
    outputs(10645) <= not(layer2_outputs(8616));
    outputs(10646) <= not((layer2_outputs(7494)) xor (layer2_outputs(7398)));
    outputs(10647) <= not((layer2_outputs(5652)) xor (layer2_outputs(529)));
    outputs(10648) <= not(layer2_outputs(7894));
    outputs(10649) <= not(layer2_outputs(9385));
    outputs(10650) <= layer2_outputs(11433);
    outputs(10651) <= not(layer2_outputs(8697)) or (layer2_outputs(2782));
    outputs(10652) <= layer2_outputs(350);
    outputs(10653) <= (layer2_outputs(5078)) xor (layer2_outputs(2672));
    outputs(10654) <= (layer2_outputs(858)) and not (layer2_outputs(8982));
    outputs(10655) <= not(layer2_outputs(1731)) or (layer2_outputs(1790));
    outputs(10656) <= not(layer2_outputs(9311));
    outputs(10657) <= not((layer2_outputs(7940)) xor (layer2_outputs(12128)));
    outputs(10658) <= (layer2_outputs(8950)) and not (layer2_outputs(11355));
    outputs(10659) <= not(layer2_outputs(5534)) or (layer2_outputs(7364));
    outputs(10660) <= not(layer2_outputs(3648));
    outputs(10661) <= not((layer2_outputs(9100)) xor (layer2_outputs(2864)));
    outputs(10662) <= (layer2_outputs(9340)) and not (layer2_outputs(1648));
    outputs(10663) <= (layer2_outputs(11028)) xor (layer2_outputs(3975));
    outputs(10664) <= not((layer2_outputs(184)) and (layer2_outputs(8173)));
    outputs(10665) <= (layer2_outputs(5057)) xor (layer2_outputs(347));
    outputs(10666) <= not(layer2_outputs(1608)) or (layer2_outputs(7307));
    outputs(10667) <= not((layer2_outputs(11495)) xor (layer2_outputs(5954)));
    outputs(10668) <= not((layer2_outputs(4560)) xor (layer2_outputs(8719)));
    outputs(10669) <= not(layer2_outputs(12437));
    outputs(10670) <= layer2_outputs(4727);
    outputs(10671) <= not((layer2_outputs(12672)) or (layer2_outputs(3871)));
    outputs(10672) <= (layer2_outputs(5446)) xor (layer2_outputs(11571));
    outputs(10673) <= not((layer2_outputs(4232)) xor (layer2_outputs(7196)));
    outputs(10674) <= layer2_outputs(8510);
    outputs(10675) <= not((layer2_outputs(10359)) xor (layer2_outputs(7150)));
    outputs(10676) <= (layer2_outputs(12020)) xor (layer2_outputs(4270));
    outputs(10677) <= layer2_outputs(7696);
    outputs(10678) <= not(layer2_outputs(5186));
    outputs(10679) <= (layer2_outputs(9556)) xor (layer2_outputs(3253));
    outputs(10680) <= not(layer2_outputs(11215));
    outputs(10681) <= layer2_outputs(3143);
    outputs(10682) <= (layer2_outputs(8261)) or (layer2_outputs(6576));
    outputs(10683) <= (layer2_outputs(3721)) xor (layer2_outputs(129));
    outputs(10684) <= not(layer2_outputs(1414));
    outputs(10685) <= not(layer2_outputs(10595)) or (layer2_outputs(4));
    outputs(10686) <= not(layer2_outputs(572));
    outputs(10687) <= not((layer2_outputs(2518)) xor (layer2_outputs(1703)));
    outputs(10688) <= not((layer2_outputs(11182)) xor (layer2_outputs(7404)));
    outputs(10689) <= layer2_outputs(1351);
    outputs(10690) <= (layer2_outputs(6694)) and not (layer2_outputs(6601));
    outputs(10691) <= (layer2_outputs(153)) or (layer2_outputs(3809));
    outputs(10692) <= not((layer2_outputs(6972)) or (layer2_outputs(504)));
    outputs(10693) <= (layer2_outputs(11676)) xor (layer2_outputs(5299));
    outputs(10694) <= not(layer2_outputs(3760));
    outputs(10695) <= not((layer2_outputs(8443)) and (layer2_outputs(5433)));
    outputs(10696) <= (layer2_outputs(341)) xor (layer2_outputs(3449));
    outputs(10697) <= (layer2_outputs(2372)) xor (layer2_outputs(6249));
    outputs(10698) <= not((layer2_outputs(9914)) xor (layer2_outputs(2890)));
    outputs(10699) <= layer2_outputs(11153);
    outputs(10700) <= (layer2_outputs(2582)) xor (layer2_outputs(3012));
    outputs(10701) <= not(layer2_outputs(10070)) or (layer2_outputs(9574));
    outputs(10702) <= layer2_outputs(6250);
    outputs(10703) <= (layer2_outputs(9354)) and not (layer2_outputs(10867));
    outputs(10704) <= not(layer2_outputs(4875));
    outputs(10705) <= not(layer2_outputs(10256)) or (layer2_outputs(7764));
    outputs(10706) <= (layer2_outputs(11770)) and (layer2_outputs(2127));
    outputs(10707) <= not((layer2_outputs(11317)) xor (layer2_outputs(4528)));
    outputs(10708) <= (layer2_outputs(1881)) xor (layer2_outputs(6127));
    outputs(10709) <= (layer2_outputs(869)) xor (layer2_outputs(4472));
    outputs(10710) <= layer2_outputs(431);
    outputs(10711) <= layer2_outputs(11686);
    outputs(10712) <= layer2_outputs(10272);
    outputs(10713) <= not(layer2_outputs(4854));
    outputs(10714) <= layer2_outputs(8933);
    outputs(10715) <= not((layer2_outputs(10717)) xor (layer2_outputs(8059)));
    outputs(10716) <= layer2_outputs(11438);
    outputs(10717) <= layer2_outputs(12473);
    outputs(10718) <= not((layer2_outputs(1068)) and (layer2_outputs(5840)));
    outputs(10719) <= layer2_outputs(9818);
    outputs(10720) <= layer2_outputs(1411);
    outputs(10721) <= not(layer2_outputs(9483));
    outputs(10722) <= not(layer2_outputs(4366));
    outputs(10723) <= (layer2_outputs(12196)) and not (layer2_outputs(9478));
    outputs(10724) <= layer2_outputs(934);
    outputs(10725) <= not(layer2_outputs(3514));
    outputs(10726) <= layer2_outputs(11623);
    outputs(10727) <= layer2_outputs(558);
    outputs(10728) <= not(layer2_outputs(3843));
    outputs(10729) <= not((layer2_outputs(10856)) xor (layer2_outputs(8379)));
    outputs(10730) <= (layer2_outputs(10480)) and (layer2_outputs(9324));
    outputs(10731) <= (layer2_outputs(8908)) xor (layer2_outputs(8233));
    outputs(10732) <= not(layer2_outputs(3105)) or (layer2_outputs(1327));
    outputs(10733) <= not(layer2_outputs(4524));
    outputs(10734) <= not(layer2_outputs(9600));
    outputs(10735) <= not(layer2_outputs(6830));
    outputs(10736) <= layer2_outputs(2271);
    outputs(10737) <= not((layer2_outputs(488)) xor (layer2_outputs(2180)));
    outputs(10738) <= not(layer2_outputs(11520));
    outputs(10739) <= not((layer2_outputs(12648)) or (layer2_outputs(4258)));
    outputs(10740) <= layer2_outputs(12098);
    outputs(10741) <= not((layer2_outputs(395)) and (layer2_outputs(5127)));
    outputs(10742) <= not(layer2_outputs(3939));
    outputs(10743) <= layer2_outputs(12402);
    outputs(10744) <= not(layer2_outputs(7400));
    outputs(10745) <= not(layer2_outputs(7108));
    outputs(10746) <= not((layer2_outputs(8016)) xor (layer2_outputs(1605)));
    outputs(10747) <= (layer2_outputs(11166)) xor (layer2_outputs(2601));
    outputs(10748) <= (layer2_outputs(10843)) xor (layer2_outputs(3823));
    outputs(10749) <= layer2_outputs(9154);
    outputs(10750) <= layer2_outputs(1639);
    outputs(10751) <= not((layer2_outputs(4058)) and (layer2_outputs(3475)));
    outputs(10752) <= not((layer2_outputs(5097)) and (layer2_outputs(1046)));
    outputs(10753) <= not((layer2_outputs(10808)) and (layer2_outputs(12577)));
    outputs(10754) <= not(layer2_outputs(6885));
    outputs(10755) <= not(layer2_outputs(10779));
    outputs(10756) <= not((layer2_outputs(10511)) xor (layer2_outputs(4064)));
    outputs(10757) <= not((layer2_outputs(12027)) xor (layer2_outputs(1204)));
    outputs(10758) <= not(layer2_outputs(10400)) or (layer2_outputs(413));
    outputs(10759) <= not(layer2_outputs(10752));
    outputs(10760) <= layer2_outputs(4304);
    outputs(10761) <= (layer2_outputs(6167)) xor (layer2_outputs(1188));
    outputs(10762) <= not(layer2_outputs(10962));
    outputs(10763) <= not(layer2_outputs(12055)) or (layer2_outputs(2063));
    outputs(10764) <= not(layer2_outputs(394)) or (layer2_outputs(1540));
    outputs(10765) <= layer2_outputs(4185);
    outputs(10766) <= not(layer2_outputs(3596)) or (layer2_outputs(2185));
    outputs(10767) <= not((layer2_outputs(2878)) xor (layer2_outputs(1474)));
    outputs(10768) <= (layer2_outputs(6058)) xor (layer2_outputs(8999));
    outputs(10769) <= layer2_outputs(12084);
    outputs(10770) <= layer2_outputs(3525);
    outputs(10771) <= layer2_outputs(9513);
    outputs(10772) <= not((layer2_outputs(6366)) xor (layer2_outputs(9033)));
    outputs(10773) <= (layer2_outputs(9546)) and not (layer2_outputs(12284));
    outputs(10774) <= not((layer2_outputs(9403)) xor (layer2_outputs(2075)));
    outputs(10775) <= not(layer2_outputs(8605));
    outputs(10776) <= not(layer2_outputs(9478));
    outputs(10777) <= layer2_outputs(11258);
    outputs(10778) <= layer2_outputs(11587);
    outputs(10779) <= not((layer2_outputs(12798)) or (layer2_outputs(5766)));
    outputs(10780) <= not((layer2_outputs(12486)) and (layer2_outputs(6177)));
    outputs(10781) <= layer2_outputs(2493);
    outputs(10782) <= layer2_outputs(9192);
    outputs(10783) <= not((layer2_outputs(6460)) xor (layer2_outputs(11977)));
    outputs(10784) <= not((layer2_outputs(10262)) xor (layer2_outputs(422)));
    outputs(10785) <= not(layer2_outputs(8758)) or (layer2_outputs(8156));
    outputs(10786) <= not((layer2_outputs(10356)) xor (layer2_outputs(3260)));
    outputs(10787) <= (layer2_outputs(10258)) and not (layer2_outputs(7475));
    outputs(10788) <= not(layer2_outputs(10038)) or (layer2_outputs(6850));
    outputs(10789) <= not(layer2_outputs(8584));
    outputs(10790) <= not(layer2_outputs(1499));
    outputs(10791) <= not((layer2_outputs(399)) xor (layer2_outputs(4719)));
    outputs(10792) <= layer2_outputs(1705);
    outputs(10793) <= (layer2_outputs(9843)) or (layer2_outputs(5527));
    outputs(10794) <= not(layer2_outputs(9817));
    outputs(10795) <= not(layer2_outputs(11178)) or (layer2_outputs(2417));
    outputs(10796) <= layer2_outputs(6258);
    outputs(10797) <= layer2_outputs(3752);
    outputs(10798) <= not((layer2_outputs(4597)) and (layer2_outputs(9073)));
    outputs(10799) <= not(layer2_outputs(9509));
    outputs(10800) <= (layer2_outputs(1842)) xor (layer2_outputs(3660));
    outputs(10801) <= layer2_outputs(10306);
    outputs(10802) <= layer2_outputs(7787);
    outputs(10803) <= not(layer2_outputs(1675));
    outputs(10804) <= not((layer2_outputs(2285)) xor (layer2_outputs(7098)));
    outputs(10805) <= not(layer2_outputs(8861)) or (layer2_outputs(3706));
    outputs(10806) <= not((layer2_outputs(4755)) xor (layer2_outputs(150)));
    outputs(10807) <= layer2_outputs(12723);
    outputs(10808) <= (layer2_outputs(10633)) xor (layer2_outputs(12551));
    outputs(10809) <= (layer2_outputs(12759)) xor (layer2_outputs(5156));
    outputs(10810) <= not((layer2_outputs(3426)) xor (layer2_outputs(6410)));
    outputs(10811) <= not(layer2_outputs(1446));
    outputs(10812) <= not(layer2_outputs(3418));
    outputs(10813) <= layer2_outputs(2168);
    outputs(10814) <= (layer2_outputs(12117)) and (layer2_outputs(7904));
    outputs(10815) <= layer2_outputs(5894);
    outputs(10816) <= not((layer2_outputs(3368)) xor (layer2_outputs(4598)));
    outputs(10817) <= (layer2_outputs(11380)) xor (layer2_outputs(10809));
    outputs(10818) <= not(layer2_outputs(4731));
    outputs(10819) <= layer2_outputs(12091);
    outputs(10820) <= not((layer2_outputs(505)) xor (layer2_outputs(7728)));
    outputs(10821) <= layer2_outputs(11621);
    outputs(10822) <= not((layer2_outputs(10536)) xor (layer2_outputs(10787)));
    outputs(10823) <= not(layer2_outputs(12436));
    outputs(10824) <= (layer2_outputs(7551)) or (layer2_outputs(12783));
    outputs(10825) <= (layer2_outputs(9252)) and (layer2_outputs(7213));
    outputs(10826) <= not(layer2_outputs(760));
    outputs(10827) <= layer2_outputs(6897);
    outputs(10828) <= not(layer2_outputs(5481));
    outputs(10829) <= not(layer2_outputs(12796));
    outputs(10830) <= not((layer2_outputs(6834)) and (layer2_outputs(7539)));
    outputs(10831) <= layer2_outputs(11378);
    outputs(10832) <= layer2_outputs(12089);
    outputs(10833) <= not(layer2_outputs(2441));
    outputs(10834) <= not(layer2_outputs(8231));
    outputs(10835) <= layer2_outputs(2321);
    outputs(10836) <= layer2_outputs(1900);
    outputs(10837) <= not((layer2_outputs(11424)) xor (layer2_outputs(375)));
    outputs(10838) <= not(layer2_outputs(6677));
    outputs(10839) <= layer2_outputs(11007);
    outputs(10840) <= not(layer2_outputs(4225));
    outputs(10841) <= (layer2_outputs(8769)) and (layer2_outputs(6808));
    outputs(10842) <= not(layer2_outputs(992));
    outputs(10843) <= not(layer2_outputs(300));
    outputs(10844) <= not(layer2_outputs(11241));
    outputs(10845) <= not(layer2_outputs(2055)) or (layer2_outputs(2678));
    outputs(10846) <= layer2_outputs(4016);
    outputs(10847) <= not(layer2_outputs(6254));
    outputs(10848) <= not(layer2_outputs(11412));
    outputs(10849) <= layer2_outputs(8224);
    outputs(10850) <= layer2_outputs(10883);
    outputs(10851) <= layer2_outputs(6033);
    outputs(10852) <= (layer2_outputs(12698)) xor (layer2_outputs(2491));
    outputs(10853) <= not((layer2_outputs(11622)) xor (layer2_outputs(4375)));
    outputs(10854) <= (layer2_outputs(11207)) xor (layer2_outputs(3512));
    outputs(10855) <= (layer2_outputs(8870)) and not (layer2_outputs(12231));
    outputs(10856) <= not((layer2_outputs(5509)) xor (layer2_outputs(3572)));
    outputs(10857) <= (layer2_outputs(5211)) and (layer2_outputs(11734));
    outputs(10858) <= not(layer2_outputs(2931)) or (layer2_outputs(7764));
    outputs(10859) <= not((layer2_outputs(11310)) xor (layer2_outputs(319)));
    outputs(10860) <= not((layer2_outputs(11266)) xor (layer2_outputs(7334)));
    outputs(10861) <= (layer2_outputs(5174)) xor (layer2_outputs(7882));
    outputs(10862) <= (layer2_outputs(5189)) xor (layer2_outputs(8030));
    outputs(10863) <= layer2_outputs(4239);
    outputs(10864) <= (layer2_outputs(11575)) or (layer2_outputs(8898));
    outputs(10865) <= (layer2_outputs(9190)) xor (layer2_outputs(9529));
    outputs(10866) <= (layer2_outputs(3759)) xor (layer2_outputs(7101));
    outputs(10867) <= layer2_outputs(3701);
    outputs(10868) <= layer2_outputs(7096);
    outputs(10869) <= layer2_outputs(10827);
    outputs(10870) <= (layer2_outputs(5307)) or (layer2_outputs(2273));
    outputs(10871) <= not(layer2_outputs(4045));
    outputs(10872) <= (layer2_outputs(9967)) xor (layer2_outputs(196));
    outputs(10873) <= not(layer2_outputs(12518)) or (layer2_outputs(3628));
    outputs(10874) <= not((layer2_outputs(8743)) and (layer2_outputs(1054)));
    outputs(10875) <= (layer2_outputs(2177)) xor (layer2_outputs(2359));
    outputs(10876) <= layer2_outputs(1314);
    outputs(10877) <= not(layer2_outputs(10849));
    outputs(10878) <= not(layer2_outputs(12796));
    outputs(10879) <= (layer2_outputs(10548)) xor (layer2_outputs(1907));
    outputs(10880) <= layer2_outputs(12715);
    outputs(10881) <= not((layer2_outputs(11788)) and (layer2_outputs(6140)));
    outputs(10882) <= (layer2_outputs(4181)) xor (layer2_outputs(9263));
    outputs(10883) <= layer2_outputs(9640);
    outputs(10884) <= layer2_outputs(9475);
    outputs(10885) <= not(layer2_outputs(4446));
    outputs(10886) <= layer2_outputs(8227);
    outputs(10887) <= not(layer2_outputs(8290));
    outputs(10888) <= not(layer2_outputs(11868));
    outputs(10889) <= not(layer2_outputs(12307)) or (layer2_outputs(1781));
    outputs(10890) <= not((layer2_outputs(5873)) xor (layer2_outputs(8845)));
    outputs(10891) <= layer2_outputs(4168);
    outputs(10892) <= not((layer2_outputs(6894)) xor (layer2_outputs(1889)));
    outputs(10893) <= not((layer2_outputs(9328)) and (layer2_outputs(12792)));
    outputs(10894) <= (layer2_outputs(542)) or (layer2_outputs(1460));
    outputs(10895) <= layer2_outputs(2265);
    outputs(10896) <= layer2_outputs(11571);
    outputs(10897) <= (layer2_outputs(3920)) or (layer2_outputs(2629));
    outputs(10898) <= (layer2_outputs(6096)) xor (layer2_outputs(4604));
    outputs(10899) <= layer2_outputs(924);
    outputs(10900) <= layer2_outputs(8383);
    outputs(10901) <= layer2_outputs(3903);
    outputs(10902) <= layer2_outputs(11342);
    outputs(10903) <= layer2_outputs(2676);
    outputs(10904) <= not((layer2_outputs(2455)) xor (layer2_outputs(10452)));
    outputs(10905) <= not((layer2_outputs(335)) xor (layer2_outputs(1788)));
    outputs(10906) <= layer2_outputs(10405);
    outputs(10907) <= layer2_outputs(675);
    outputs(10908) <= not(layer2_outputs(2474));
    outputs(10909) <= (layer2_outputs(12282)) and (layer2_outputs(4262));
    outputs(10910) <= not(layer2_outputs(3800)) or (layer2_outputs(4056));
    outputs(10911) <= not(layer2_outputs(4135));
    outputs(10912) <= not(layer2_outputs(11025));
    outputs(10913) <= layer2_outputs(12559);
    outputs(10914) <= (layer2_outputs(2129)) xor (layer2_outputs(4881));
    outputs(10915) <= (layer2_outputs(3252)) xor (layer2_outputs(11717));
    outputs(10916) <= (layer2_outputs(11142)) xor (layer2_outputs(9496));
    outputs(10917) <= not(layer2_outputs(2372));
    outputs(10918) <= not((layer2_outputs(5515)) xor (layer2_outputs(8259)));
    outputs(10919) <= layer2_outputs(6921);
    outputs(10920) <= not(layer2_outputs(5274));
    outputs(10921) <= (layer2_outputs(3209)) xor (layer2_outputs(9346));
    outputs(10922) <= (layer2_outputs(3128)) xor (layer2_outputs(712));
    outputs(10923) <= (layer2_outputs(1352)) or (layer2_outputs(10089));
    outputs(10924) <= layer2_outputs(9876);
    outputs(10925) <= not((layer2_outputs(3954)) xor (layer2_outputs(3791)));
    outputs(10926) <= layer2_outputs(1389);
    outputs(10927) <= not((layer2_outputs(3271)) xor (layer2_outputs(11921)));
    outputs(10928) <= (layer2_outputs(11722)) and (layer2_outputs(2727));
    outputs(10929) <= not(layer2_outputs(3617));
    outputs(10930) <= layer2_outputs(2379);
    outputs(10931) <= layer2_outputs(391);
    outputs(10932) <= not((layer2_outputs(6609)) xor (layer2_outputs(2410)));
    outputs(10933) <= layer2_outputs(1828);
    outputs(10934) <= layer2_outputs(5176);
    outputs(10935) <= not(layer2_outputs(1550));
    outputs(10936) <= not(layer2_outputs(9700)) or (layer2_outputs(2364));
    outputs(10937) <= not((layer2_outputs(1840)) xor (layer2_outputs(6493)));
    outputs(10938) <= (layer2_outputs(5181)) xor (layer2_outputs(7553));
    outputs(10939) <= not(layer2_outputs(1580));
    outputs(10940) <= not(layer2_outputs(11649));
    outputs(10941) <= (layer2_outputs(2498)) xor (layer2_outputs(4664));
    outputs(10942) <= not((layer2_outputs(184)) and (layer2_outputs(1008)));
    outputs(10943) <= (layer2_outputs(2851)) and (layer2_outputs(9586));
    outputs(10944) <= not(layer2_outputs(12615));
    outputs(10945) <= (layer2_outputs(6671)) or (layer2_outputs(8282));
    outputs(10946) <= not((layer2_outputs(5874)) xor (layer2_outputs(2223)));
    outputs(10947) <= not(layer2_outputs(7327));
    outputs(10948) <= (layer2_outputs(1645)) xor (layer2_outputs(1958));
    outputs(10949) <= not((layer2_outputs(2347)) xor (layer2_outputs(7130)));
    outputs(10950) <= layer2_outputs(10748);
    outputs(10951) <= not((layer2_outputs(1217)) xor (layer2_outputs(3478)));
    outputs(10952) <= layer2_outputs(11804);
    outputs(10953) <= not(layer2_outputs(4588)) or (layer2_outputs(5054));
    outputs(10954) <= (layer2_outputs(387)) or (layer2_outputs(2464));
    outputs(10955) <= layer2_outputs(7110);
    outputs(10956) <= layer2_outputs(1066);
    outputs(10957) <= layer2_outputs(2665);
    outputs(10958) <= not((layer2_outputs(7142)) xor (layer2_outputs(3828)));
    outputs(10959) <= not((layer2_outputs(11899)) xor (layer2_outputs(6853)));
    outputs(10960) <= (layer2_outputs(11670)) xor (layer2_outputs(9055));
    outputs(10961) <= not(layer2_outputs(10588)) or (layer2_outputs(3615));
    outputs(10962) <= not(layer2_outputs(1719));
    outputs(10963) <= not(layer2_outputs(11291));
    outputs(10964) <= (layer2_outputs(9229)) xor (layer2_outputs(6023));
    outputs(10965) <= (layer2_outputs(6505)) xor (layer2_outputs(788));
    outputs(10966) <= not((layer2_outputs(2545)) and (layer2_outputs(6298)));
    outputs(10967) <= not(layer2_outputs(6372)) or (layer2_outputs(4715));
    outputs(10968) <= not((layer2_outputs(6472)) xor (layer2_outputs(7022)));
    outputs(10969) <= layer2_outputs(7081);
    outputs(10970) <= not(layer2_outputs(453));
    outputs(10971) <= layer2_outputs(11660);
    outputs(10972) <= (layer2_outputs(312)) and (layer2_outputs(6908));
    outputs(10973) <= (layer2_outputs(6120)) xor (layer2_outputs(3084));
    outputs(10974) <= layer2_outputs(8423);
    outputs(10975) <= not((layer2_outputs(4713)) and (layer2_outputs(4392)));
    outputs(10976) <= (layer2_outputs(89)) xor (layer2_outputs(697));
    outputs(10977) <= not(layer2_outputs(4423));
    outputs(10978) <= layer2_outputs(2912);
    outputs(10979) <= not((layer2_outputs(1974)) xor (layer2_outputs(170)));
    outputs(10980) <= layer2_outputs(2194);
    outputs(10981) <= not(layer2_outputs(8357)) or (layer2_outputs(7752));
    outputs(10982) <= layer2_outputs(3671);
    outputs(10983) <= not(layer2_outputs(11513)) or (layer2_outputs(3119));
    outputs(10984) <= not((layer2_outputs(10907)) xor (layer2_outputs(3055)));
    outputs(10985) <= not(layer2_outputs(10535));
    outputs(10986) <= not(layer2_outputs(9509));
    outputs(10987) <= (layer2_outputs(6413)) xor (layer2_outputs(2929));
    outputs(10988) <= not((layer2_outputs(7760)) xor (layer2_outputs(8281)));
    outputs(10989) <= (layer2_outputs(3131)) xor (layer2_outputs(1740));
    outputs(10990) <= not((layer2_outputs(6368)) and (layer2_outputs(7736)));
    outputs(10991) <= (layer2_outputs(4253)) and not (layer2_outputs(2651));
    outputs(10992) <= not(layer2_outputs(12629));
    outputs(10993) <= not(layer2_outputs(12687));
    outputs(10994) <= (layer2_outputs(4685)) or (layer2_outputs(10323));
    outputs(10995) <= not((layer2_outputs(3856)) and (layer2_outputs(9937)));
    outputs(10996) <= not(layer2_outputs(10587));
    outputs(10997) <= not(layer2_outputs(4125));
    outputs(10998) <= not(layer2_outputs(7392));
    outputs(10999) <= '1';
    outputs(11000) <= not(layer2_outputs(5557));
    outputs(11001) <= layer2_outputs(3247);
    outputs(11002) <= not(layer2_outputs(7560));
    outputs(11003) <= not((layer2_outputs(12097)) xor (layer2_outputs(10842)));
    outputs(11004) <= not((layer2_outputs(5470)) xor (layer2_outputs(9121)));
    outputs(11005) <= not(layer2_outputs(12775));
    outputs(11006) <= not((layer2_outputs(6049)) xor (layer2_outputs(6319)));
    outputs(11007) <= (layer2_outputs(11165)) xor (layer2_outputs(3750));
    outputs(11008) <= not(layer2_outputs(7770));
    outputs(11009) <= (layer2_outputs(11386)) xor (layer2_outputs(7478));
    outputs(11010) <= not(layer2_outputs(3725));
    outputs(11011) <= not((layer2_outputs(2091)) xor (layer2_outputs(3360)));
    outputs(11012) <= (layer2_outputs(7389)) xor (layer2_outputs(2746));
    outputs(11013) <= (layer2_outputs(12240)) xor (layer2_outputs(8382));
    outputs(11014) <= not(layer2_outputs(10028)) or (layer2_outputs(5193));
    outputs(11015) <= layer2_outputs(1411);
    outputs(11016) <= not(layer2_outputs(9312));
    outputs(11017) <= not((layer2_outputs(6944)) xor (layer2_outputs(5921)));
    outputs(11018) <= not(layer2_outputs(12618));
    outputs(11019) <= not(layer2_outputs(11364));
    outputs(11020) <= layer2_outputs(12032);
    outputs(11021) <= not(layer2_outputs(5177));
    outputs(11022) <= (layer2_outputs(11227)) and (layer2_outputs(10979));
    outputs(11023) <= not((layer2_outputs(11251)) xor (layer2_outputs(3492)));
    outputs(11024) <= layer2_outputs(9029);
    outputs(11025) <= not(layer2_outputs(5784));
    outputs(11026) <= (layer2_outputs(4994)) xor (layer2_outputs(11841));
    outputs(11027) <= layer2_outputs(7251);
    outputs(11028) <= (layer2_outputs(136)) and not (layer2_outputs(8845));
    outputs(11029) <= (layer2_outputs(11851)) xor (layer2_outputs(10161));
    outputs(11030) <= not((layer2_outputs(7460)) xor (layer2_outputs(531)));
    outputs(11031) <= not(layer2_outputs(3461));
    outputs(11032) <= not(layer2_outputs(9608));
    outputs(11033) <= (layer2_outputs(10598)) xor (layer2_outputs(4890));
    outputs(11034) <= (layer2_outputs(4716)) xor (layer2_outputs(12746));
    outputs(11035) <= not(layer2_outputs(1878));
    outputs(11036) <= not((layer2_outputs(10589)) xor (layer2_outputs(4992)));
    outputs(11037) <= layer2_outputs(7787);
    outputs(11038) <= layer2_outputs(6291);
    outputs(11039) <= not((layer2_outputs(1628)) and (layer2_outputs(12699)));
    outputs(11040) <= (layer2_outputs(4348)) and (layer2_outputs(6446));
    outputs(11041) <= (layer2_outputs(11546)) or (layer2_outputs(4540));
    outputs(11042) <= (layer2_outputs(1896)) or (layer2_outputs(12371));
    outputs(11043) <= layer2_outputs(8878);
    outputs(11044) <= (layer2_outputs(10175)) and not (layer2_outputs(2425));
    outputs(11045) <= not(layer2_outputs(11998));
    outputs(11046) <= not(layer2_outputs(9957)) or (layer2_outputs(2219));
    outputs(11047) <= layer2_outputs(617);
    outputs(11048) <= (layer2_outputs(6997)) xor (layer2_outputs(251));
    outputs(11049) <= not(layer2_outputs(3805));
    outputs(11050) <= not((layer2_outputs(6479)) or (layer2_outputs(6072)));
    outputs(11051) <= layer2_outputs(11621);
    outputs(11052) <= layer2_outputs(238);
    outputs(11053) <= not(layer2_outputs(3464)) or (layer2_outputs(2492));
    outputs(11054) <= (layer2_outputs(3448)) xor (layer2_outputs(11806));
    outputs(11055) <= not(layer2_outputs(9861));
    outputs(11056) <= layer2_outputs(282);
    outputs(11057) <= not((layer2_outputs(4926)) and (layer2_outputs(1341)));
    outputs(11058) <= (layer2_outputs(4697)) xor (layer2_outputs(2309));
    outputs(11059) <= not(layer2_outputs(7892));
    outputs(11060) <= (layer2_outputs(1953)) xor (layer2_outputs(4837));
    outputs(11061) <= not(layer2_outputs(9495));
    outputs(11062) <= layer2_outputs(8232);
    outputs(11063) <= layer2_outputs(3841);
    outputs(11064) <= layer2_outputs(12221);
    outputs(11065) <= not((layer2_outputs(2559)) xor (layer2_outputs(3243)));
    outputs(11066) <= (layer2_outputs(9326)) or (layer2_outputs(41));
    outputs(11067) <= not(layer2_outputs(1006));
    outputs(11068) <= layer2_outputs(4941);
    outputs(11069) <= not(layer2_outputs(6990));
    outputs(11070) <= layer2_outputs(10351);
    outputs(11071) <= not(layer2_outputs(65));
    outputs(11072) <= not(layer2_outputs(7426));
    outputs(11073) <= (layer2_outputs(4043)) xor (layer2_outputs(11059));
    outputs(11074) <= layer2_outputs(9301);
    outputs(11075) <= (layer2_outputs(5649)) xor (layer2_outputs(3018));
    outputs(11076) <= not(layer2_outputs(12512));
    outputs(11077) <= layer2_outputs(4612);
    outputs(11078) <= layer2_outputs(4490);
    outputs(11079) <= (layer2_outputs(2966)) and not (layer2_outputs(9661));
    outputs(11080) <= layer2_outputs(1984);
    outputs(11081) <= not(layer2_outputs(6786)) or (layer2_outputs(10221));
    outputs(11082) <= not(layer2_outputs(7211));
    outputs(11083) <= not(layer2_outputs(10340));
    outputs(11084) <= not(layer2_outputs(5741));
    outputs(11085) <= not(layer2_outputs(5681));
    outputs(11086) <= not(layer2_outputs(11338));
    outputs(11087) <= (layer2_outputs(7841)) or (layer2_outputs(2419));
    outputs(11088) <= not(layer2_outputs(12395)) or (layer2_outputs(4604));
    outputs(11089) <= not(layer2_outputs(724));
    outputs(11090) <= layer2_outputs(3223);
    outputs(11091) <= layer2_outputs(5618);
    outputs(11092) <= (layer2_outputs(426)) xor (layer2_outputs(1091));
    outputs(11093) <= (layer2_outputs(7947)) xor (layer2_outputs(5266));
    outputs(11094) <= (layer2_outputs(5200)) xor (layer2_outputs(10355));
    outputs(11095) <= not(layer2_outputs(76));
    outputs(11096) <= not((layer2_outputs(9039)) xor (layer2_outputs(4570)));
    outputs(11097) <= layer2_outputs(3009);
    outputs(11098) <= (layer2_outputs(12508)) or (layer2_outputs(4523));
    outputs(11099) <= layer2_outputs(3187);
    outputs(11100) <= (layer2_outputs(2187)) or (layer2_outputs(3133));
    outputs(11101) <= layer2_outputs(2467);
    outputs(11102) <= not((layer2_outputs(7692)) xor (layer2_outputs(9319)));
    outputs(11103) <= not((layer2_outputs(9186)) xor (layer2_outputs(11394)));
    outputs(11104) <= not(layer2_outputs(4020));
    outputs(11105) <= not(layer2_outputs(11681));
    outputs(11106) <= not(layer2_outputs(5751)) or (layer2_outputs(8073));
    outputs(11107) <= not(layer2_outputs(4761)) or (layer2_outputs(5495));
    outputs(11108) <= (layer2_outputs(11105)) xor (layer2_outputs(7844));
    outputs(11109) <= layer2_outputs(1363);
    outputs(11110) <= not(layer2_outputs(10370));
    outputs(11111) <= layer2_outputs(2469);
    outputs(11112) <= not(layer2_outputs(4433));
    outputs(11113) <= not((layer2_outputs(439)) xor (layer2_outputs(2658)));
    outputs(11114) <= layer2_outputs(2780);
    outputs(11115) <= layer2_outputs(6958);
    outputs(11116) <= not(layer2_outputs(390)) or (layer2_outputs(12209));
    outputs(11117) <= not(layer2_outputs(3445)) or (layer2_outputs(8025));
    outputs(11118) <= (layer2_outputs(10354)) xor (layer2_outputs(11675));
    outputs(11119) <= not(layer2_outputs(603)) or (layer2_outputs(1509));
    outputs(11120) <= layer2_outputs(10405);
    outputs(11121) <= (layer2_outputs(11371)) xor (layer2_outputs(12460));
    outputs(11122) <= layer2_outputs(1412);
    outputs(11123) <= not(layer2_outputs(6195));
    outputs(11124) <= layer2_outputs(2753);
    outputs(11125) <= not((layer2_outputs(11632)) xor (layer2_outputs(1749)));
    outputs(11126) <= not(layer2_outputs(6699)) or (layer2_outputs(148));
    outputs(11127) <= layer2_outputs(4464);
    outputs(11128) <= not((layer2_outputs(388)) and (layer2_outputs(8141)));
    outputs(11129) <= layer2_outputs(2264);
    outputs(11130) <= (layer2_outputs(10227)) xor (layer2_outputs(12149));
    outputs(11131) <= layer2_outputs(2694);
    outputs(11132) <= not(layer2_outputs(9312));
    outputs(11133) <= not((layer2_outputs(808)) xor (layer2_outputs(11790)));
    outputs(11134) <= layer2_outputs(8795);
    outputs(11135) <= (layer2_outputs(9933)) or (layer2_outputs(8458));
    outputs(11136) <= (layer2_outputs(1338)) or (layer2_outputs(7109));
    outputs(11137) <= not(layer2_outputs(3990)) or (layer2_outputs(4794));
    outputs(11138) <= (layer2_outputs(2440)) xor (layer2_outputs(5491));
    outputs(11139) <= not((layer2_outputs(7941)) xor (layer2_outputs(4611)));
    outputs(11140) <= not(layer2_outputs(10468));
    outputs(11141) <= not(layer2_outputs(10826)) or (layer2_outputs(3686));
    outputs(11142) <= layer2_outputs(2697);
    outputs(11143) <= (layer2_outputs(6973)) and (layer2_outputs(2947));
    outputs(11144) <= layer2_outputs(2155);
    outputs(11145) <= layer2_outputs(7953);
    outputs(11146) <= not((layer2_outputs(1141)) xor (layer2_outputs(12389)));
    outputs(11147) <= not((layer2_outputs(4382)) or (layer2_outputs(7442)));
    outputs(11148) <= layer2_outputs(8869);
    outputs(11149) <= layer2_outputs(12195);
    outputs(11150) <= not(layer2_outputs(5999));
    outputs(11151) <= layer2_outputs(8163);
    outputs(11152) <= (layer2_outputs(114)) or (layer2_outputs(4121));
    outputs(11153) <= not(layer2_outputs(735));
    outputs(11154) <= not(layer2_outputs(4250)) or (layer2_outputs(1970));
    outputs(11155) <= not(layer2_outputs(4988));
    outputs(11156) <= not((layer2_outputs(11912)) or (layer2_outputs(3571)));
    outputs(11157) <= (layer2_outputs(10864)) xor (layer2_outputs(4287));
    outputs(11158) <= layer2_outputs(493);
    outputs(11159) <= (layer2_outputs(2556)) and not (layer2_outputs(10861));
    outputs(11160) <= layer2_outputs(7077);
    outputs(11161) <= (layer2_outputs(9437)) xor (layer2_outputs(8871));
    outputs(11162) <= layer2_outputs(13);
    outputs(11163) <= layer2_outputs(10739);
    outputs(11164) <= (layer2_outputs(8851)) xor (layer2_outputs(1700));
    outputs(11165) <= not((layer2_outputs(4374)) and (layer2_outputs(10288)));
    outputs(11166) <= layer2_outputs(1420);
    outputs(11167) <= (layer2_outputs(12319)) and not (layer2_outputs(143));
    outputs(11168) <= not((layer2_outputs(2945)) xor (layer2_outputs(7540)));
    outputs(11169) <= not(layer2_outputs(8106));
    outputs(11170) <= layer2_outputs(2153);
    outputs(11171) <= not(layer2_outputs(7294));
    outputs(11172) <= layer2_outputs(10720);
    outputs(11173) <= (layer2_outputs(4494)) or (layer2_outputs(6560));
    outputs(11174) <= not(layer2_outputs(3399));
    outputs(11175) <= layer2_outputs(10466);
    outputs(11176) <= (layer2_outputs(3757)) xor (layer2_outputs(3260));
    outputs(11177) <= not((layer2_outputs(938)) xor (layer2_outputs(11163)));
    outputs(11178) <= (layer2_outputs(5043)) xor (layer2_outputs(5947));
    outputs(11179) <= layer2_outputs(5865);
    outputs(11180) <= layer2_outputs(4380);
    outputs(11181) <= (layer2_outputs(8431)) xor (layer2_outputs(6128));
    outputs(11182) <= not(layer2_outputs(12285));
    outputs(11183) <= (layer2_outputs(7497)) and not (layer2_outputs(11672));
    outputs(11184) <= (layer2_outputs(1670)) and not (layer2_outputs(5815));
    outputs(11185) <= (layer2_outputs(5968)) or (layer2_outputs(9521));
    outputs(11186) <= not((layer2_outputs(8693)) xor (layer2_outputs(12563)));
    outputs(11187) <= not((layer2_outputs(3806)) or (layer2_outputs(2240)));
    outputs(11188) <= not((layer2_outputs(118)) or (layer2_outputs(4791)));
    outputs(11189) <= not(layer2_outputs(11046));
    outputs(11190) <= not(layer2_outputs(7221)) or (layer2_outputs(2597));
    outputs(11191) <= layer2_outputs(7693);
    outputs(11192) <= (layer2_outputs(10793)) xor (layer2_outputs(6376));
    outputs(11193) <= (layer2_outputs(6738)) and not (layer2_outputs(12239));
    outputs(11194) <= not(layer2_outputs(807)) or (layer2_outputs(11555));
    outputs(11195) <= (layer2_outputs(7578)) and (layer2_outputs(2717));
    outputs(11196) <= not(layer2_outputs(4275));
    outputs(11197) <= (layer2_outputs(6459)) or (layer2_outputs(7145));
    outputs(11198) <= not(layer2_outputs(666));
    outputs(11199) <= layer2_outputs(3647);
    outputs(11200) <= (layer2_outputs(1321)) or (layer2_outputs(2785));
    outputs(11201) <= not(layer2_outputs(11576)) or (layer2_outputs(12308));
    outputs(11202) <= not((layer2_outputs(8441)) xor (layer2_outputs(4165)));
    outputs(11203) <= (layer2_outputs(7313)) xor (layer2_outputs(6087));
    outputs(11204) <= not((layer2_outputs(1498)) and (layer2_outputs(8085)));
    outputs(11205) <= not((layer2_outputs(10794)) xor (layer2_outputs(2705)));
    outputs(11206) <= (layer2_outputs(4247)) xor (layer2_outputs(12295));
    outputs(11207) <= not(layer2_outputs(249));
    outputs(11208) <= not((layer2_outputs(12423)) xor (layer2_outputs(1199)));
    outputs(11209) <= layer2_outputs(1524);
    outputs(11210) <= not(layer2_outputs(8787));
    outputs(11211) <= not((layer2_outputs(8429)) or (layer2_outputs(3352)));
    outputs(11212) <= not((layer2_outputs(11268)) xor (layer2_outputs(258)));
    outputs(11213) <= layer2_outputs(2151);
    outputs(11214) <= not(layer2_outputs(1322));
    outputs(11215) <= not(layer2_outputs(6227));
    outputs(11216) <= not((layer2_outputs(9882)) xor (layer2_outputs(9221)));
    outputs(11217) <= not(layer2_outputs(384));
    outputs(11218) <= not((layer2_outputs(12246)) or (layer2_outputs(12699)));
    outputs(11219) <= not(layer2_outputs(656));
    outputs(11220) <= not(layer2_outputs(10597));
    outputs(11221) <= not((layer2_outputs(5685)) xor (layer2_outputs(12118)));
    outputs(11222) <= '1';
    outputs(11223) <= not(layer2_outputs(12173));
    outputs(11224) <= (layer2_outputs(7248)) or (layer2_outputs(663));
    outputs(11225) <= not(layer2_outputs(10445)) or (layer2_outputs(37));
    outputs(11226) <= not((layer2_outputs(2028)) and (layer2_outputs(5937)));
    outputs(11227) <= not((layer2_outputs(544)) xor (layer2_outputs(7611)));
    outputs(11228) <= layer2_outputs(1003);
    outputs(11229) <= layer2_outputs(10940);
    outputs(11230) <= not((layer2_outputs(4073)) xor (layer2_outputs(703)));
    outputs(11231) <= (layer2_outputs(12535)) xor (layer2_outputs(1595));
    outputs(11232) <= not(layer2_outputs(9376));
    outputs(11233) <= (layer2_outputs(7122)) xor (layer2_outputs(3011));
    outputs(11234) <= layer2_outputs(5930);
    outputs(11235) <= not(layer2_outputs(3784));
    outputs(11236) <= (layer2_outputs(6055)) xor (layer2_outputs(4569));
    outputs(11237) <= layer2_outputs(1708);
    outputs(11238) <= layer2_outputs(10654);
    outputs(11239) <= not((layer2_outputs(848)) and (layer2_outputs(11669)));
    outputs(11240) <= not((layer2_outputs(6430)) and (layer2_outputs(8198)));
    outputs(11241) <= layer2_outputs(7165);
    outputs(11242) <= layer2_outputs(12417);
    outputs(11243) <= not((layer2_outputs(9276)) or (layer2_outputs(2940)));
    outputs(11244) <= not((layer2_outputs(12700)) or (layer2_outputs(1888)));
    outputs(11245) <= (layer2_outputs(12401)) xor (layer2_outputs(3167));
    outputs(11246) <= not(layer2_outputs(5757));
    outputs(11247) <= (layer2_outputs(3836)) xor (layer2_outputs(4316));
    outputs(11248) <= (layer2_outputs(4859)) xor (layer2_outputs(4648));
    outputs(11249) <= layer2_outputs(9867);
    outputs(11250) <= (layer2_outputs(4168)) and not (layer2_outputs(1769));
    outputs(11251) <= (layer2_outputs(11885)) or (layer2_outputs(10743));
    outputs(11252) <= layer2_outputs(9404);
    outputs(11253) <= not(layer2_outputs(2805)) or (layer2_outputs(3591));
    outputs(11254) <= not((layer2_outputs(10456)) xor (layer2_outputs(9486)));
    outputs(11255) <= layer2_outputs(2682);
    outputs(11256) <= not(layer2_outputs(4680));
    outputs(11257) <= not(layer2_outputs(7722));
    outputs(11258) <= (layer2_outputs(6908)) and (layer2_outputs(12534));
    outputs(11259) <= '0';
    outputs(11260) <= layer2_outputs(2882);
    outputs(11261) <= not((layer2_outputs(9487)) xor (layer2_outputs(12558)));
    outputs(11262) <= not(layer2_outputs(1192));
    outputs(11263) <= (layer2_outputs(1433)) or (layer2_outputs(110));
    outputs(11264) <= layer2_outputs(6012);
    outputs(11265) <= not(layer2_outputs(3030));
    outputs(11266) <= (layer2_outputs(7677)) and not (layer2_outputs(680));
    outputs(11267) <= not((layer2_outputs(9748)) xor (layer2_outputs(6896)));
    outputs(11268) <= not(layer2_outputs(12499));
    outputs(11269) <= not((layer2_outputs(1235)) xor (layer2_outputs(7440)));
    outputs(11270) <= not(layer2_outputs(10671));
    outputs(11271) <= not((layer2_outputs(4956)) xor (layer2_outputs(11874)));
    outputs(11272) <= not((layer2_outputs(11353)) xor (layer2_outputs(12303)));
    outputs(11273) <= layer2_outputs(9353);
    outputs(11274) <= (layer2_outputs(11701)) xor (layer2_outputs(10058));
    outputs(11275) <= (layer2_outputs(4362)) and not (layer2_outputs(6368));
    outputs(11276) <= layer2_outputs(6592);
    outputs(11277) <= (layer2_outputs(8105)) xor (layer2_outputs(9720));
    outputs(11278) <= layer2_outputs(4609);
    outputs(11279) <= not(layer2_outputs(9519)) or (layer2_outputs(12324));
    outputs(11280) <= (layer2_outputs(6992)) and (layer2_outputs(4055));
    outputs(11281) <= not((layer2_outputs(4565)) xor (layer2_outputs(8755)));
    outputs(11282) <= (layer2_outputs(8581)) xor (layer2_outputs(5066));
    outputs(11283) <= not(layer2_outputs(10261));
    outputs(11284) <= not(layer2_outputs(294));
    outputs(11285) <= not((layer2_outputs(7699)) and (layer2_outputs(4776)));
    outputs(11286) <= not(layer2_outputs(12679));
    outputs(11287) <= layer2_outputs(4922);
    outputs(11288) <= not(layer2_outputs(11058));
    outputs(11289) <= not((layer2_outputs(9782)) xor (layer2_outputs(10478)));
    outputs(11290) <= not(layer2_outputs(10807));
    outputs(11291) <= not((layer2_outputs(12029)) xor (layer2_outputs(903)));
    outputs(11292) <= not((layer2_outputs(1714)) xor (layer2_outputs(11128)));
    outputs(11293) <= not(layer2_outputs(9401));
    outputs(11294) <= layer2_outputs(6772);
    outputs(11295) <= layer2_outputs(4730);
    outputs(11296) <= not(layer2_outputs(4036));
    outputs(11297) <= (layer2_outputs(4102)) xor (layer2_outputs(231));
    outputs(11298) <= layer2_outputs(389);
    outputs(11299) <= layer2_outputs(11597);
    outputs(11300) <= layer2_outputs(6092);
    outputs(11301) <= not((layer2_outputs(5031)) xor (layer2_outputs(9005)));
    outputs(11302) <= layer2_outputs(7798);
    outputs(11303) <= not((layer2_outputs(10418)) and (layer2_outputs(4011)));
    outputs(11304) <= layer2_outputs(3455);
    outputs(11305) <= (layer2_outputs(11409)) xor (layer2_outputs(2281));
    outputs(11306) <= (layer2_outputs(1902)) xor (layer2_outputs(2177));
    outputs(11307) <= (layer2_outputs(10612)) xor (layer2_outputs(5546));
    outputs(11308) <= (layer2_outputs(3456)) xor (layer2_outputs(2349));
    outputs(11309) <= not((layer2_outputs(12603)) or (layer2_outputs(902)));
    outputs(11310) <= not((layer2_outputs(5064)) or (layer2_outputs(7817)));
    outputs(11311) <= not((layer2_outputs(6433)) or (layer2_outputs(11393)));
    outputs(11312) <= (layer2_outputs(1224)) xor (layer2_outputs(5294));
    outputs(11313) <= not((layer2_outputs(9517)) xor (layer2_outputs(252)));
    outputs(11314) <= not(layer2_outputs(6059));
    outputs(11315) <= layer2_outputs(5920);
    outputs(11316) <= layer2_outputs(11966);
    outputs(11317) <= not(layer2_outputs(1225)) or (layer2_outputs(9941));
    outputs(11318) <= layer2_outputs(2321);
    outputs(11319) <= not(layer2_outputs(7164));
    outputs(11320) <= (layer2_outputs(11663)) xor (layer2_outputs(10080));
    outputs(11321) <= not(layer2_outputs(906));
    outputs(11322) <= layer2_outputs(12631);
    outputs(11323) <= not(layer2_outputs(2037));
    outputs(11324) <= not((layer2_outputs(11898)) and (layer2_outputs(5370)));
    outputs(11325) <= layer2_outputs(1242);
    outputs(11326) <= (layer2_outputs(10562)) xor (layer2_outputs(1897));
    outputs(11327) <= (layer2_outputs(2041)) xor (layer2_outputs(7343));
    outputs(11328) <= not((layer2_outputs(2739)) xor (layer2_outputs(6363)));
    outputs(11329) <= not((layer2_outputs(10959)) and (layer2_outputs(7688)));
    outputs(11330) <= layer2_outputs(4916);
    outputs(11331) <= not((layer2_outputs(5542)) xor (layer2_outputs(6088)));
    outputs(11332) <= (layer2_outputs(4507)) xor (layer2_outputs(5306));
    outputs(11333) <= layer2_outputs(12031);
    outputs(11334) <= layer2_outputs(6893);
    outputs(11335) <= (layer2_outputs(3133)) and (layer2_outputs(1587));
    outputs(11336) <= (layer2_outputs(8452)) xor (layer2_outputs(3661));
    outputs(11337) <= (layer2_outputs(9505)) or (layer2_outputs(4509));
    outputs(11338) <= not((layer2_outputs(4575)) or (layer2_outputs(5612)));
    outputs(11339) <= layer2_outputs(12113);
    outputs(11340) <= layer2_outputs(970);
    outputs(11341) <= not((layer2_outputs(4226)) xor (layer2_outputs(12156)));
    outputs(11342) <= layer2_outputs(10732);
    outputs(11343) <= not((layer2_outputs(12785)) and (layer2_outputs(631)));
    outputs(11344) <= not((layer2_outputs(256)) xor (layer2_outputs(5700)));
    outputs(11345) <= layer2_outputs(9468);
    outputs(11346) <= not(layer2_outputs(167));
    outputs(11347) <= not(layer2_outputs(8741));
    outputs(11348) <= not((layer2_outputs(6054)) xor (layer2_outputs(10613)));
    outputs(11349) <= (layer2_outputs(6747)) and (layer2_outputs(8747));
    outputs(11350) <= (layer2_outputs(11481)) xor (layer2_outputs(6652));
    outputs(11351) <= layer2_outputs(7684);
    outputs(11352) <= layer2_outputs(11987);
    outputs(11353) <= not(layer2_outputs(2175));
    outputs(11354) <= (layer2_outputs(9715)) xor (layer2_outputs(5004));
    outputs(11355) <= layer2_outputs(10985);
    outputs(11356) <= not((layer2_outputs(12370)) xor (layer2_outputs(11994)));
    outputs(11357) <= layer2_outputs(8150);
    outputs(11358) <= layer2_outputs(7474);
    outputs(11359) <= not((layer2_outputs(9138)) and (layer2_outputs(8812)));
    outputs(11360) <= not((layer2_outputs(7156)) xor (layer2_outputs(4519)));
    outputs(11361) <= not(layer2_outputs(7434)) or (layer2_outputs(2832));
    outputs(11362) <= layer2_outputs(7010);
    outputs(11363) <= (layer2_outputs(4044)) xor (layer2_outputs(4285));
    outputs(11364) <= layer2_outputs(12430);
    outputs(11365) <= layer2_outputs(4857);
    outputs(11366) <= not(layer2_outputs(11268));
    outputs(11367) <= layer2_outputs(5627);
    outputs(11368) <= (layer2_outputs(7722)) xor (layer2_outputs(9182));
    outputs(11369) <= not(layer2_outputs(9783));
    outputs(11370) <= (layer2_outputs(10132)) xor (layer2_outputs(10130));
    outputs(11371) <= (layer2_outputs(1473)) or (layer2_outputs(7066));
    outputs(11372) <= not((layer2_outputs(6232)) and (layer2_outputs(2775)));
    outputs(11373) <= (layer2_outputs(9902)) xor (layer2_outputs(5698));
    outputs(11374) <= (layer2_outputs(2428)) and not (layer2_outputs(7128));
    outputs(11375) <= not(layer2_outputs(11646));
    outputs(11376) <= not((layer2_outputs(2330)) xor (layer2_outputs(10638)));
    outputs(11377) <= layer2_outputs(11115);
    outputs(11378) <= not(layer2_outputs(6175));
    outputs(11379) <= not(layer2_outputs(2759));
    outputs(11380) <= (layer2_outputs(2631)) xor (layer2_outputs(7044));
    outputs(11381) <= layer2_outputs(681);
    outputs(11382) <= not((layer2_outputs(9508)) xor (layer2_outputs(9285)));
    outputs(11383) <= layer2_outputs(3646);
    outputs(11384) <= not((layer2_outputs(12596)) xor (layer2_outputs(6255)));
    outputs(11385) <= not((layer2_outputs(11256)) xor (layer2_outputs(593)));
    outputs(11386) <= layer2_outputs(9598);
    outputs(11387) <= not((layer2_outputs(1844)) xor (layer2_outputs(12292)));
    outputs(11388) <= (layer2_outputs(6479)) xor (layer2_outputs(6272));
    outputs(11389) <= not(layer2_outputs(11649));
    outputs(11390) <= (layer2_outputs(12227)) or (layer2_outputs(6899));
    outputs(11391) <= not(layer2_outputs(10284));
    outputs(11392) <= not(layer2_outputs(8186));
    outputs(11393) <= not(layer2_outputs(4632));
    outputs(11394) <= not(layer2_outputs(8928)) or (layer2_outputs(11852));
    outputs(11395) <= layer2_outputs(6261);
    outputs(11396) <= layer2_outputs(5371);
    outputs(11397) <= not(layer2_outputs(11548));
    outputs(11398) <= (layer2_outputs(6221)) xor (layer2_outputs(8709));
    outputs(11399) <= not((layer2_outputs(8099)) and (layer2_outputs(12641)));
    outputs(11400) <= not(layer2_outputs(5239)) or (layer2_outputs(7472));
    outputs(11401) <= not(layer2_outputs(12115));
    outputs(11402) <= not(layer2_outputs(2070));
    outputs(11403) <= not(layer2_outputs(1468));
    outputs(11404) <= not(layer2_outputs(284));
    outputs(11405) <= layer2_outputs(1798);
    outputs(11406) <= (layer2_outputs(6301)) xor (layer2_outputs(11163));
    outputs(11407) <= (layer2_outputs(11089)) or (layer2_outputs(7190));
    outputs(11408) <= not((layer2_outputs(2636)) xor (layer2_outputs(11318)));
    outputs(11409) <= (layer2_outputs(9350)) or (layer2_outputs(5464));
    outputs(11410) <= layer2_outputs(9854);
    outputs(11411) <= not((layer2_outputs(5419)) xor (layer2_outputs(2499)));
    outputs(11412) <= (layer2_outputs(5825)) xor (layer2_outputs(5443));
    outputs(11413) <= not(layer2_outputs(7478)) or (layer2_outputs(2053));
    outputs(11414) <= (layer2_outputs(2015)) and (layer2_outputs(3345));
    outputs(11415) <= layer2_outputs(4043);
    outputs(11416) <= not(layer2_outputs(9096));
    outputs(11417) <= layer2_outputs(7349);
    outputs(11418) <= layer2_outputs(1254);
    outputs(11419) <= not(layer2_outputs(10790)) or (layer2_outputs(5841));
    outputs(11420) <= not((layer2_outputs(10025)) xor (layer2_outputs(11579)));
    outputs(11421) <= layer2_outputs(2330);
    outputs(11422) <= not(layer2_outputs(1854));
    outputs(11423) <= not((layer2_outputs(6114)) and (layer2_outputs(4037)));
    outputs(11424) <= layer2_outputs(10718);
    outputs(11425) <= not((layer2_outputs(6126)) xor (layer2_outputs(6689)));
    outputs(11426) <= not(layer2_outputs(9924)) or (layer2_outputs(9));
    outputs(11427) <= layer2_outputs(11327);
    outputs(11428) <= not((layer2_outputs(3991)) xor (layer2_outputs(6543)));
    outputs(11429) <= not((layer2_outputs(8799)) and (layer2_outputs(1732)));
    outputs(11430) <= not((layer2_outputs(6545)) xor (layer2_outputs(10900)));
    outputs(11431) <= not(layer2_outputs(7831)) or (layer2_outputs(6115));
    outputs(11432) <= not((layer2_outputs(10465)) xor (layer2_outputs(10492)));
    outputs(11433) <= layer2_outputs(7828);
    outputs(11434) <= not((layer2_outputs(1988)) xor (layer2_outputs(11534)));
    outputs(11435) <= not(layer2_outputs(2474));
    outputs(11436) <= (layer2_outputs(12358)) and (layer2_outputs(6730));
    outputs(11437) <= not(layer2_outputs(5179));
    outputs(11438) <= (layer2_outputs(11274)) xor (layer2_outputs(3090));
    outputs(11439) <= layer2_outputs(2076);
    outputs(11440) <= not(layer2_outputs(3081)) or (layer2_outputs(4726));
    outputs(11441) <= layer2_outputs(9923);
    outputs(11442) <= not(layer2_outputs(7617)) or (layer2_outputs(2828));
    outputs(11443) <= (layer2_outputs(7966)) xor (layer2_outputs(3470));
    outputs(11444) <= layer2_outputs(2808);
    outputs(11445) <= not(layer2_outputs(6129));
    outputs(11446) <= not((layer2_outputs(9679)) xor (layer2_outputs(4213)));
    outputs(11447) <= (layer2_outputs(2085)) or (layer2_outputs(11423));
    outputs(11448) <= not(layer2_outputs(2161));
    outputs(11449) <= layer2_outputs(6436);
    outputs(11450) <= (layer2_outputs(264)) xor (layer2_outputs(8923));
    outputs(11451) <= (layer2_outputs(7347)) and (layer2_outputs(6636));
    outputs(11452) <= not((layer2_outputs(1203)) xor (layer2_outputs(7889)));
    outputs(11453) <= not(layer2_outputs(10233));
    outputs(11454) <= not((layer2_outputs(128)) xor (layer2_outputs(8909)));
    outputs(11455) <= not((layer2_outputs(12493)) xor (layer2_outputs(2732)));
    outputs(11456) <= not(layer2_outputs(12094));
    outputs(11457) <= (layer2_outputs(3773)) xor (layer2_outputs(767));
    outputs(11458) <= not((layer2_outputs(9925)) xor (layer2_outputs(1037)));
    outputs(11459) <= not((layer2_outputs(1671)) and (layer2_outputs(9511)));
    outputs(11460) <= layer2_outputs(8323);
    outputs(11461) <= not(layer2_outputs(2394)) or (layer2_outputs(1471));
    outputs(11462) <= not((layer2_outputs(5118)) xor (layer2_outputs(10178)));
    outputs(11463) <= not(layer2_outputs(12367)) or (layer2_outputs(1859));
    outputs(11464) <= not(layer2_outputs(11849)) or (layer2_outputs(2873));
    outputs(11465) <= (layer2_outputs(4751)) xor (layer2_outputs(6678));
    outputs(11466) <= layer2_outputs(8856);
    outputs(11467) <= not((layer2_outputs(12718)) or (layer2_outputs(3498)));
    outputs(11468) <= not((layer2_outputs(7661)) xor (layer2_outputs(2249)));
    outputs(11469) <= (layer2_outputs(42)) xor (layer2_outputs(2820));
    outputs(11470) <= not(layer2_outputs(6412));
    outputs(11471) <= (layer2_outputs(11206)) xor (layer2_outputs(2431));
    outputs(11472) <= (layer2_outputs(5450)) or (layer2_outputs(11662));
    outputs(11473) <= (layer2_outputs(11532)) xor (layer2_outputs(12070));
    outputs(11474) <= not((layer2_outputs(11882)) xor (layer2_outputs(1393)));
    outputs(11475) <= (layer2_outputs(7843)) xor (layer2_outputs(3663));
    outputs(11476) <= (layer2_outputs(16)) xor (layer2_outputs(5453));
    outputs(11477) <= (layer2_outputs(1161)) or (layer2_outputs(9010));
    outputs(11478) <= (layer2_outputs(12343)) xor (layer2_outputs(8263));
    outputs(11479) <= layer2_outputs(6956);
    outputs(11480) <= (layer2_outputs(10306)) xor (layer2_outputs(2324));
    outputs(11481) <= (layer2_outputs(2418)) xor (layer2_outputs(8181));
    outputs(11482) <= not(layer2_outputs(8579));
    outputs(11483) <= layer2_outputs(7372);
    outputs(11484) <= not(layer2_outputs(4894));
    outputs(11485) <= layer2_outputs(3841);
    outputs(11486) <= layer2_outputs(5308);
    outputs(11487) <= layer2_outputs(170);
    outputs(11488) <= (layer2_outputs(9944)) and (layer2_outputs(9124));
    outputs(11489) <= not(layer2_outputs(2907));
    outputs(11490) <= not(layer2_outputs(10493));
    outputs(11491) <= not(layer2_outputs(9430));
    outputs(11492) <= (layer2_outputs(11671)) xor (layer2_outputs(10667));
    outputs(11493) <= not((layer2_outputs(6858)) xor (layer2_outputs(5175)));
    outputs(11494) <= not(layer2_outputs(9269));
    outputs(11495) <= layer2_outputs(2935);
    outputs(11496) <= (layer2_outputs(628)) xor (layer2_outputs(7070));
    outputs(11497) <= (layer2_outputs(12321)) xor (layer2_outputs(12538));
    outputs(11498) <= layer2_outputs(8449);
    outputs(11499) <= not(layer2_outputs(2803));
    outputs(11500) <= layer2_outputs(5015);
    outputs(11501) <= not(layer2_outputs(11741));
    outputs(11502) <= layer2_outputs(4834);
    outputs(11503) <= not(layer2_outputs(8902));
    outputs(11504) <= not(layer2_outputs(3095));
    outputs(11505) <= not((layer2_outputs(416)) xor (layer2_outputs(376)));
    outputs(11506) <= not(layer2_outputs(6186));
    outputs(11507) <= not(layer2_outputs(4522));
    outputs(11508) <= not(layer2_outputs(8791)) or (layer2_outputs(3176));
    outputs(11509) <= (layer2_outputs(2719)) xor (layer2_outputs(2915));
    outputs(11510) <= not(layer2_outputs(1078)) or (layer2_outputs(6577));
    outputs(11511) <= (layer2_outputs(1131)) and not (layer2_outputs(5146));
    outputs(11512) <= not(layer2_outputs(9534)) or (layer2_outputs(4081));
    outputs(11513) <= not(layer2_outputs(9927)) or (layer2_outputs(11125));
    outputs(11514) <= layer2_outputs(11590);
    outputs(11515) <= not(layer2_outputs(6932));
    outputs(11516) <= not(layer2_outputs(1715));
    outputs(11517) <= not((layer2_outputs(10691)) or (layer2_outputs(1767)));
    outputs(11518) <= layer2_outputs(1852);
    outputs(11519) <= (layer2_outputs(11541)) xor (layer2_outputs(2042));
    outputs(11520) <= layer2_outputs(6806);
    outputs(11521) <= layer2_outputs(12021);
    outputs(11522) <= not((layer2_outputs(5126)) xor (layer2_outputs(5861)));
    outputs(11523) <= (layer2_outputs(8478)) xor (layer2_outputs(6598));
    outputs(11524) <= (layer2_outputs(12462)) and not (layer2_outputs(6424));
    outputs(11525) <= (layer2_outputs(7384)) xor (layer2_outputs(2038));
    outputs(11526) <= layer2_outputs(10903);
    outputs(11527) <= not(layer2_outputs(12396));
    outputs(11528) <= (layer2_outputs(3590)) and (layer2_outputs(12198));
    outputs(11529) <= not(layer2_outputs(2035));
    outputs(11530) <= (layer2_outputs(4596)) or (layer2_outputs(11545));
    outputs(11531) <= not((layer2_outputs(9489)) xor (layer2_outputs(4178)));
    outputs(11532) <= not(layer2_outputs(6424));
    outputs(11533) <= layer2_outputs(5383);
    outputs(11534) <= (layer2_outputs(1869)) xor (layer2_outputs(12632));
    outputs(11535) <= not(layer2_outputs(5198));
    outputs(11536) <= not((layer2_outputs(642)) xor (layer2_outputs(12075)));
    outputs(11537) <= not((layer2_outputs(8258)) xor (layer2_outputs(4228)));
    outputs(11538) <= not(layer2_outputs(10151));
    outputs(11539) <= not(layer2_outputs(6109)) or (layer2_outputs(6600));
    outputs(11540) <= (layer2_outputs(3589)) and not (layer2_outputs(1401));
    outputs(11541) <= layer2_outputs(1900);
    outputs(11542) <= layer2_outputs(895);
    outputs(11543) <= layer2_outputs(936);
    outputs(11544) <= not((layer2_outputs(12485)) xor (layer2_outputs(4149)));
    outputs(11545) <= not(layer2_outputs(380));
    outputs(11546) <= layer2_outputs(5220);
    outputs(11547) <= (layer2_outputs(1374)) xor (layer2_outputs(8545));
    outputs(11548) <= not(layer2_outputs(190));
    outputs(11549) <= not((layer2_outputs(7331)) or (layer2_outputs(4270)));
    outputs(11550) <= not(layer2_outputs(11492));
    outputs(11551) <= not(layer2_outputs(8655));
    outputs(11552) <= layer2_outputs(10682);
    outputs(11553) <= not(layer2_outputs(12276));
    outputs(11554) <= not(layer2_outputs(3717));
    outputs(11555) <= layer2_outputs(7778);
    outputs(11556) <= not(layer2_outputs(10378));
    outputs(11557) <= (layer2_outputs(8418)) and not (layer2_outputs(2137));
    outputs(11558) <= not(layer2_outputs(3035));
    outputs(11559) <= not(layer2_outputs(6693));
    outputs(11560) <= layer2_outputs(12514);
    outputs(11561) <= not(layer2_outputs(10799));
    outputs(11562) <= not((layer2_outputs(3454)) xor (layer2_outputs(4021)));
    outputs(11563) <= not(layer2_outputs(10253));
    outputs(11564) <= layer2_outputs(3127);
    outputs(11565) <= not(layer2_outputs(12784));
    outputs(11566) <= (layer2_outputs(1345)) xor (layer2_outputs(9985));
    outputs(11567) <= not(layer2_outputs(4243));
    outputs(11568) <= not((layer2_outputs(5337)) xor (layer2_outputs(8987)));
    outputs(11569) <= layer2_outputs(4370);
    outputs(11570) <= layer2_outputs(387);
    outputs(11571) <= layer2_outputs(9468);
    outputs(11572) <= layer2_outputs(7485);
    outputs(11573) <= not((layer2_outputs(11457)) and (layer2_outputs(4140)));
    outputs(11574) <= layer2_outputs(4263);
    outputs(11575) <= (layer2_outputs(350)) and not (layer2_outputs(5879));
    outputs(11576) <= not(layer2_outputs(3630));
    outputs(11577) <= layer2_outputs(5622);
    outputs(11578) <= layer2_outputs(568);
    outputs(11579) <= layer2_outputs(3801);
    outputs(11580) <= not(layer2_outputs(3782));
    outputs(11581) <= (layer2_outputs(9248)) xor (layer2_outputs(12608));
    outputs(11582) <= not(layer2_outputs(12025)) or (layer2_outputs(10579));
    outputs(11583) <= layer2_outputs(3772);
    outputs(11584) <= (layer2_outputs(6243)) xor (layer2_outputs(324));
    outputs(11585) <= not(layer2_outputs(2737));
    outputs(11586) <= not(layer2_outputs(984));
    outputs(11587) <= not(layer2_outputs(11445));
    outputs(11588) <= not(layer2_outputs(4406));
    outputs(11589) <= not(layer2_outputs(3422));
    outputs(11590) <= not((layer2_outputs(5373)) and (layer2_outputs(11375)));
    outputs(11591) <= not(layer2_outputs(1057));
    outputs(11592) <= (layer2_outputs(6710)) xor (layer2_outputs(2955));
    outputs(11593) <= not((layer2_outputs(24)) xor (layer2_outputs(9081)));
    outputs(11594) <= not(layer2_outputs(12611));
    outputs(11595) <= (layer2_outputs(11794)) or (layer2_outputs(12277));
    outputs(11596) <= not(layer2_outputs(3200)) or (layer2_outputs(6136));
    outputs(11597) <= not(layer2_outputs(9869));
    outputs(11598) <= layer2_outputs(12254);
    outputs(11599) <= layer2_outputs(10414);
    outputs(11600) <= (layer2_outputs(202)) and (layer2_outputs(4182));
    outputs(11601) <= layer2_outputs(776);
    outputs(11602) <= not(layer2_outputs(7968));
    outputs(11603) <= layer2_outputs(8777);
    outputs(11604) <= layer2_outputs(7231);
    outputs(11605) <= not((layer2_outputs(4441)) and (layer2_outputs(3320)));
    outputs(11606) <= (layer2_outputs(8715)) xor (layer2_outputs(2877));
    outputs(11607) <= layer2_outputs(7965);
    outputs(11608) <= (layer2_outputs(447)) xor (layer2_outputs(5607));
    outputs(11609) <= not(layer2_outputs(11841)) or (layer2_outputs(7032));
    outputs(11610) <= not((layer2_outputs(2336)) or (layer2_outputs(11177)));
    outputs(11611) <= not(layer2_outputs(2078)) or (layer2_outputs(8617));
    outputs(11612) <= layer2_outputs(260);
    outputs(11613) <= layer2_outputs(2456);
    outputs(11614) <= not(layer2_outputs(2846));
    outputs(11615) <= layer2_outputs(3325);
    outputs(11616) <= not(layer2_outputs(972));
    outputs(11617) <= (layer2_outputs(2655)) and not (layer2_outputs(1753));
    outputs(11618) <= (layer2_outputs(12610)) xor (layer2_outputs(1136));
    outputs(11619) <= (layer2_outputs(4307)) xor (layer2_outputs(11417));
    outputs(11620) <= not(layer2_outputs(6903));
    outputs(11621) <= layer2_outputs(1812);
    outputs(11622) <= (layer2_outputs(9417)) and not (layer2_outputs(7443));
    outputs(11623) <= (layer2_outputs(4420)) and not (layer2_outputs(8778));
    outputs(11624) <= (layer2_outputs(5271)) xor (layer2_outputs(6927));
    outputs(11625) <= not((layer2_outputs(8696)) xor (layer2_outputs(5492)));
    outputs(11626) <= not((layer2_outputs(10456)) xor (layer2_outputs(9692)));
    outputs(11627) <= not((layer2_outputs(4061)) or (layer2_outputs(7417)));
    outputs(11628) <= not(layer2_outputs(6467)) or (layer2_outputs(3375));
    outputs(11629) <= (layer2_outputs(1011)) and (layer2_outputs(5872));
    outputs(11630) <= not(layer2_outputs(12181)) or (layer2_outputs(5620));
    outputs(11631) <= not(layer2_outputs(8550));
    outputs(11632) <= layer2_outputs(6814);
    outputs(11633) <= not((layer2_outputs(12633)) xor (layer2_outputs(5116)));
    outputs(11634) <= not(layer2_outputs(8892));
    outputs(11635) <= (layer2_outputs(3557)) and not (layer2_outputs(12664));
    outputs(11636) <= not((layer2_outputs(5139)) xor (layer2_outputs(7739)));
    outputs(11637) <= (layer2_outputs(1218)) xor (layer2_outputs(3379));
    outputs(11638) <= not((layer2_outputs(2346)) xor (layer2_outputs(4469)));
    outputs(11639) <= not(layer2_outputs(5566));
    outputs(11640) <= layer2_outputs(6429);
    outputs(11641) <= (layer2_outputs(12155)) xor (layer2_outputs(4196));
    outputs(11642) <= not((layer2_outputs(8205)) xor (layer2_outputs(971)));
    outputs(11643) <= not(layer2_outputs(9215));
    outputs(11644) <= not((layer2_outputs(6410)) xor (layer2_outputs(4286)));
    outputs(11645) <= not(layer2_outputs(754)) or (layer2_outputs(7223));
    outputs(11646) <= (layer2_outputs(11389)) and not (layer2_outputs(10879));
    outputs(11647) <= (layer2_outputs(3835)) and (layer2_outputs(8669));
    outputs(11648) <= layer2_outputs(9620);
    outputs(11649) <= layer2_outputs(1723);
    outputs(11650) <= not(layer2_outputs(2940));
    outputs(11651) <= layer2_outputs(2985);
    outputs(11652) <= not(layer2_outputs(8647));
    outputs(11653) <= not(layer2_outputs(2001));
    outputs(11654) <= not((layer2_outputs(915)) xor (layer2_outputs(2579)));
    outputs(11655) <= not((layer2_outputs(6138)) or (layer2_outputs(2475)));
    outputs(11656) <= not(layer2_outputs(9576));
    outputs(11657) <= not(layer2_outputs(11860)) or (layer2_outputs(11819));
    outputs(11658) <= (layer2_outputs(2080)) xor (layer2_outputs(11517));
    outputs(11659) <= not(layer2_outputs(4918));
    outputs(11660) <= not(layer2_outputs(11499));
    outputs(11661) <= layer2_outputs(10234);
    outputs(11662) <= layer2_outputs(4204);
    outputs(11663) <= (layer2_outputs(4206)) xor (layer2_outputs(7638));
    outputs(11664) <= layer2_outputs(5460);
    outputs(11665) <= not(layer2_outputs(4078)) or (layer2_outputs(5153));
    outputs(11666) <= not(layer2_outputs(7053));
    outputs(11667) <= not(layer2_outputs(12190));
    outputs(11668) <= not((layer2_outputs(11221)) xor (layer2_outputs(11077)));
    outputs(11669) <= not((layer2_outputs(4477)) xor (layer2_outputs(10998)));
    outputs(11670) <= layer2_outputs(7767);
    outputs(11671) <= not((layer2_outputs(1397)) xor (layer2_outputs(6171)));
    outputs(11672) <= not(layer2_outputs(1234));
    outputs(11673) <= layer2_outputs(10246);
    outputs(11674) <= layer2_outputs(3431);
    outputs(11675) <= not(layer2_outputs(4048));
    outputs(11676) <= layer2_outputs(5383);
    outputs(11677) <= (layer2_outputs(8834)) and (layer2_outputs(3409));
    outputs(11678) <= layer2_outputs(12081);
    outputs(11679) <= (layer2_outputs(3608)) xor (layer2_outputs(998));
    outputs(11680) <= not(layer2_outputs(9132));
    outputs(11681) <= not((layer2_outputs(8650)) xor (layer2_outputs(3764)));
    outputs(11682) <= layer2_outputs(4998);
    outputs(11683) <= not(layer2_outputs(11689));
    outputs(11684) <= (layer2_outputs(6160)) or (layer2_outputs(4718));
    outputs(11685) <= layer2_outputs(10724);
    outputs(11686) <= not((layer2_outputs(3386)) xor (layer2_outputs(148)));
    outputs(11687) <= not(layer2_outputs(5677));
    outputs(11688) <= not((layer2_outputs(4414)) and (layer2_outputs(2286)));
    outputs(11689) <= layer2_outputs(2173);
    outputs(11690) <= (layer2_outputs(2926)) or (layer2_outputs(7512));
    outputs(11691) <= layer2_outputs(9518);
    outputs(11692) <= not(layer2_outputs(73));
    outputs(11693) <= (layer2_outputs(7803)) and not (layer2_outputs(11766));
    outputs(11694) <= layer2_outputs(7540);
    outputs(11695) <= layer2_outputs(7936);
    outputs(11696) <= not((layer2_outputs(10868)) and (layer2_outputs(6152)));
    outputs(11697) <= not(layer2_outputs(4553));
    outputs(11698) <= layer2_outputs(1240);
    outputs(11699) <= not(layer2_outputs(3109));
    outputs(11700) <= (layer2_outputs(6200)) xor (layer2_outputs(8480));
    outputs(11701) <= not((layer2_outputs(2819)) xor (layer2_outputs(8277)));
    outputs(11702) <= not(layer2_outputs(10181));
    outputs(11703) <= layer2_outputs(12043);
    outputs(11704) <= layer2_outputs(3003);
    outputs(11705) <= not(layer2_outputs(5531));
    outputs(11706) <= not(layer2_outputs(9873));
    outputs(11707) <= not(layer2_outputs(1925));
    outputs(11708) <= (layer2_outputs(6720)) or (layer2_outputs(813));
    outputs(11709) <= (layer2_outputs(5180)) and (layer2_outputs(7767));
    outputs(11710) <= not(layer2_outputs(10254));
    outputs(11711) <= not(layer2_outputs(5961));
    outputs(11712) <= (layer2_outputs(1463)) xor (layer2_outputs(5904));
    outputs(11713) <= layer2_outputs(11783);
    outputs(11714) <= (layer2_outputs(10747)) and not (layer2_outputs(3338));
    outputs(11715) <= not((layer2_outputs(8574)) xor (layer2_outputs(8855)));
    outputs(11716) <= layer2_outputs(4775);
    outputs(11717) <= layer2_outputs(533);
    outputs(11718) <= not(layer2_outputs(8294));
    outputs(11719) <= layer2_outputs(7707);
    outputs(11720) <= layer2_outputs(12794);
    outputs(11721) <= not(layer2_outputs(473));
    outputs(11722) <= (layer2_outputs(9617)) and not (layer2_outputs(12154));
    outputs(11723) <= not(layer2_outputs(7711));
    outputs(11724) <= not(layer2_outputs(8415));
    outputs(11725) <= layer2_outputs(2961);
    outputs(11726) <= (layer2_outputs(3567)) xor (layer2_outputs(6079));
    outputs(11727) <= not(layer2_outputs(9252));
    outputs(11728) <= not((layer2_outputs(3584)) or (layer2_outputs(1548)));
    outputs(11729) <= (layer2_outputs(8654)) xor (layer2_outputs(2881));
    outputs(11730) <= not((layer2_outputs(4893)) or (layer2_outputs(10542)));
    outputs(11731) <= (layer2_outputs(8090)) xor (layer2_outputs(1826));
    outputs(11732) <= not(layer2_outputs(3423));
    outputs(11733) <= layer2_outputs(3995);
    outputs(11734) <= not((layer2_outputs(3813)) and (layer2_outputs(9149)));
    outputs(11735) <= not((layer2_outputs(11489)) and (layer2_outputs(8571)));
    outputs(11736) <= (layer2_outputs(10963)) xor (layer2_outputs(5332));
    outputs(11737) <= not(layer2_outputs(6155));
    outputs(11738) <= layer2_outputs(1170);
    outputs(11739) <= (layer2_outputs(6288)) and not (layer2_outputs(923));
    outputs(11740) <= not(layer2_outputs(11440));
    outputs(11741) <= (layer2_outputs(8328)) xor (layer2_outputs(6651));
    outputs(11742) <= not((layer2_outputs(9210)) and (layer2_outputs(6340)));
    outputs(11743) <= layer2_outputs(6045);
    outputs(11744) <= layer2_outputs(7576);
    outputs(11745) <= not(layer2_outputs(3946));
    outputs(11746) <= not(layer2_outputs(9932));
    outputs(11747) <= (layer2_outputs(5514)) xor (layer2_outputs(4328));
    outputs(11748) <= (layer2_outputs(9628)) xor (layer2_outputs(7459));
    outputs(11749) <= not((layer2_outputs(6841)) xor (layer2_outputs(2287)));
    outputs(11750) <= not(layer2_outputs(10671));
    outputs(11751) <= (layer2_outputs(7729)) and not (layer2_outputs(8504));
    outputs(11752) <= not(layer2_outputs(11430)) or (layer2_outputs(4571));
    outputs(11753) <= not(layer2_outputs(322));
    outputs(11754) <= not(layer2_outputs(55));
    outputs(11755) <= not(layer2_outputs(573));
    outputs(11756) <= not(layer2_outputs(6903));
    outputs(11757) <= layer2_outputs(7013);
    outputs(11758) <= (layer2_outputs(10668)) xor (layer2_outputs(9956));
    outputs(11759) <= layer2_outputs(6453);
    outputs(11760) <= (layer2_outputs(1899)) xor (layer2_outputs(1851));
    outputs(11761) <= not(layer2_outputs(6558));
    outputs(11762) <= layer2_outputs(6099);
    outputs(11763) <= not(layer2_outputs(10205));
    outputs(11764) <= not((layer2_outputs(8283)) xor (layer2_outputs(3310)));
    outputs(11765) <= layer2_outputs(179);
    outputs(11766) <= layer2_outputs(6690);
    outputs(11767) <= not(layer2_outputs(9079)) or (layer2_outputs(3641));
    outputs(11768) <= not((layer2_outputs(10194)) and (layer2_outputs(1351)));
    outputs(11769) <= not(layer2_outputs(1022));
    outputs(11770) <= not(layer2_outputs(5806)) or (layer2_outputs(10922));
    outputs(11771) <= layer2_outputs(676);
    outputs(11772) <= (layer2_outputs(7642)) xor (layer2_outputs(11611));
    outputs(11773) <= (layer2_outputs(7618)) xor (layer2_outputs(1582));
    outputs(11774) <= layer2_outputs(7187);
    outputs(11775) <= (layer2_outputs(4994)) and (layer2_outputs(3408));
    outputs(11776) <= not((layer2_outputs(9429)) xor (layer2_outputs(2297)));
    outputs(11777) <= (layer2_outputs(1795)) and (layer2_outputs(10414));
    outputs(11778) <= not(layer2_outputs(1766));
    outputs(11779) <= (layer2_outputs(1640)) xor (layer2_outputs(3281));
    outputs(11780) <= (layer2_outputs(10529)) xor (layer2_outputs(12536));
    outputs(11781) <= layer2_outputs(8610);
    outputs(11782) <= layer2_outputs(4272);
    outputs(11783) <= not((layer2_outputs(7676)) xor (layer2_outputs(1634)));
    outputs(11784) <= layer2_outputs(7360);
    outputs(11785) <= (layer2_outputs(3196)) xor (layer2_outputs(4640));
    outputs(11786) <= not(layer2_outputs(5488)) or (layer2_outputs(9994));
    outputs(11787) <= (layer2_outputs(862)) xor (layer2_outputs(5837));
    outputs(11788) <= not(layer2_outputs(10054)) or (layer2_outputs(7659));
    outputs(11789) <= not(layer2_outputs(492));
    outputs(11790) <= (layer2_outputs(11910)) and not (layer2_outputs(6427));
    outputs(11791) <= (layer2_outputs(8079)) xor (layer2_outputs(8975));
    outputs(11792) <= layer2_outputs(11730);
    outputs(11793) <= (layer2_outputs(6499)) xor (layer2_outputs(1374));
    outputs(11794) <= not(layer2_outputs(6826));
    outputs(11795) <= not(layer2_outputs(5283));
    outputs(11796) <= not(layer2_outputs(7348)) or (layer2_outputs(9267));
    outputs(11797) <= not(layer2_outputs(4462));
    outputs(11798) <= not(layer2_outputs(9000));
    outputs(11799) <= not(layer2_outputs(7851));
    outputs(11800) <= not((layer2_outputs(3796)) xor (layer2_outputs(11854)));
    outputs(11801) <= not(layer2_outputs(629));
    outputs(11802) <= layer2_outputs(3680);
    outputs(11803) <= layer2_outputs(846);
    outputs(11804) <= layer2_outputs(6736);
    outputs(11805) <= not((layer2_outputs(2644)) xor (layer2_outputs(2176)));
    outputs(11806) <= not(layer2_outputs(1378)) or (layer2_outputs(7656));
    outputs(11807) <= not(layer2_outputs(1578));
    outputs(11808) <= (layer2_outputs(2353)) and (layer2_outputs(2224));
    outputs(11809) <= not((layer2_outputs(3696)) xor (layer2_outputs(6295)));
    outputs(11810) <= not(layer2_outputs(3160));
    outputs(11811) <= layer2_outputs(11782);
    outputs(11812) <= not((layer2_outputs(1301)) xor (layer2_outputs(11573)));
    outputs(11813) <= (layer2_outputs(11739)) and (layer2_outputs(9131));
    outputs(11814) <= (layer2_outputs(11425)) and not (layer2_outputs(684));
    outputs(11815) <= layer2_outputs(7884);
    outputs(11816) <= layer2_outputs(2662);
    outputs(11817) <= layer2_outputs(11022);
    outputs(11818) <= not((layer2_outputs(6476)) or (layer2_outputs(4059)));
    outputs(11819) <= not(layer2_outputs(9699));
    outputs(11820) <= not(layer2_outputs(573));
    outputs(11821) <= not((layer2_outputs(6629)) xor (layer2_outputs(1375)));
    outputs(11822) <= not(layer2_outputs(9898));
    outputs(11823) <= (layer2_outputs(252)) xor (layer2_outputs(11768));
    outputs(11824) <= not((layer2_outputs(12265)) xor (layer2_outputs(2365)));
    outputs(11825) <= not((layer2_outputs(5966)) xor (layer2_outputs(3793)));
    outputs(11826) <= not(layer2_outputs(12371)) or (layer2_outputs(11));
    outputs(11827) <= not(layer2_outputs(3994));
    outputs(11828) <= layer2_outputs(10307);
    outputs(11829) <= layer2_outputs(12636);
    outputs(11830) <= layer2_outputs(6438);
    outputs(11831) <= not(layer2_outputs(4943));
    outputs(11832) <= layer2_outputs(9917);
    outputs(11833) <= not((layer2_outputs(989)) xor (layer2_outputs(10641)));
    outputs(11834) <= not(layer2_outputs(11135));
    outputs(11835) <= layer2_outputs(6077);
    outputs(11836) <= (layer2_outputs(7052)) xor (layer2_outputs(45));
    outputs(11837) <= not(layer2_outputs(3940)) or (layer2_outputs(3849));
    outputs(11838) <= layer2_outputs(621);
    outputs(11839) <= layer2_outputs(6618);
    outputs(11840) <= layer2_outputs(11564);
    outputs(11841) <= not(layer2_outputs(2086));
    outputs(11842) <= layer2_outputs(9173);
    outputs(11843) <= (layer2_outputs(5104)) and not (layer2_outputs(2848));
    outputs(11844) <= (layer2_outputs(2523)) xor (layer2_outputs(4938));
    outputs(11845) <= (layer2_outputs(8986)) and not (layer2_outputs(6419));
    outputs(11846) <= not(layer2_outputs(12695));
    outputs(11847) <= (layer2_outputs(10535)) and (layer2_outputs(6761));
    outputs(11848) <= not(layer2_outputs(1143));
    outputs(11849) <= not((layer2_outputs(9791)) xor (layer2_outputs(7391)));
    outputs(11850) <= layer2_outputs(2690);
    outputs(11851) <= not(layer2_outputs(8104));
    outputs(11852) <= layer2_outputs(925);
    outputs(11853) <= (layer2_outputs(6786)) xor (layer2_outputs(5898));
    outputs(11854) <= not(layer2_outputs(7546));
    outputs(11855) <= not((layer2_outputs(12665)) xor (layer2_outputs(7250)));
    outputs(11856) <= (layer2_outputs(3372)) xor (layer2_outputs(836));
    outputs(11857) <= not((layer2_outputs(1406)) xor (layer2_outputs(1047)));
    outputs(11858) <= layer2_outputs(5399);
    outputs(11859) <= not(layer2_outputs(5969));
    outputs(11860) <= (layer2_outputs(511)) and not (layer2_outputs(7328));
    outputs(11861) <= not((layer2_outputs(4624)) xor (layer2_outputs(12286)));
    outputs(11862) <= not(layer2_outputs(6123));
    outputs(11863) <= layer2_outputs(6563);
    outputs(11864) <= (layer2_outputs(4841)) and not (layer2_outputs(2756));
    outputs(11865) <= layer2_outputs(6056);
    outputs(11866) <= layer2_outputs(10461);
    outputs(11867) <= not(layer2_outputs(10192));
    outputs(11868) <= layer2_outputs(12206);
    outputs(11869) <= layer2_outputs(4095);
    outputs(11870) <= layer2_outputs(11887);
    outputs(11871) <= not((layer2_outputs(3397)) xor (layer2_outputs(7056)));
    outputs(11872) <= (layer2_outputs(8607)) xor (layer2_outputs(705));
    outputs(11873) <= layer2_outputs(7772);
    outputs(11874) <= layer2_outputs(4117);
    outputs(11875) <= not(layer2_outputs(1442));
    outputs(11876) <= not(layer2_outputs(12382));
    outputs(11877) <= not((layer2_outputs(8569)) xor (layer2_outputs(5367)));
    outputs(11878) <= layer2_outputs(5453);
    outputs(11879) <= not(layer2_outputs(5693));
    outputs(11880) <= not((layer2_outputs(5570)) and (layer2_outputs(4303)));
    outputs(11881) <= layer2_outputs(1725);
    outputs(11882) <= (layer2_outputs(11986)) xor (layer2_outputs(10118));
    outputs(11883) <= not(layer2_outputs(5139));
    outputs(11884) <= not((layer2_outputs(12406)) xor (layer2_outputs(1190)));
    outputs(11885) <= (layer2_outputs(9706)) and (layer2_outputs(8984));
    outputs(11886) <= not((layer2_outputs(3991)) xor (layer2_outputs(3734)));
    outputs(11887) <= not(layer2_outputs(12758));
    outputs(11888) <= not(layer2_outputs(4054));
    outputs(11889) <= not(layer2_outputs(6207));
    outputs(11890) <= layer2_outputs(10222);
    outputs(11891) <= not(layer2_outputs(10300));
    outputs(11892) <= (layer2_outputs(7344)) and not (layer2_outputs(5309));
    outputs(11893) <= layer2_outputs(12416);
    outputs(11894) <= not((layer2_outputs(1499)) and (layer2_outputs(8042)));
    outputs(11895) <= not((layer2_outputs(12524)) xor (layer2_outputs(8280)));
    outputs(11896) <= not(layer2_outputs(9800));
    outputs(11897) <= layer2_outputs(6658);
    outputs(11898) <= not(layer2_outputs(11180));
    outputs(11899) <= (layer2_outputs(11068)) xor (layer2_outputs(3036));
    outputs(11900) <= (layer2_outputs(9649)) and not (layer2_outputs(7364));
    outputs(11901) <= not(layer2_outputs(8211));
    outputs(11902) <= layer2_outputs(4066);
    outputs(11903) <= layer2_outputs(8926);
    outputs(11904) <= not((layer2_outputs(3936)) xor (layer2_outputs(10392)));
    outputs(11905) <= (layer2_outputs(10045)) xor (layer2_outputs(9151));
    outputs(11906) <= layer2_outputs(11734);
    outputs(11907) <= (layer2_outputs(3279)) and (layer2_outputs(3705));
    outputs(11908) <= (layer2_outputs(10923)) xor (layer2_outputs(11363));
    outputs(11909) <= not(layer2_outputs(3182));
    outputs(11910) <= layer2_outputs(7035);
    outputs(11911) <= not((layer2_outputs(1636)) xor (layer2_outputs(876)));
    outputs(11912) <= layer2_outputs(11494);
    outputs(11913) <= not(layer2_outputs(3452));
    outputs(11914) <= not(layer2_outputs(8445));
    outputs(11915) <= layer2_outputs(7092);
    outputs(11916) <= layer2_outputs(4714);
    outputs(11917) <= (layer2_outputs(905)) xor (layer2_outputs(12793));
    outputs(11918) <= not(layer2_outputs(2022));
    outputs(11919) <= (layer2_outputs(5569)) xor (layer2_outputs(10438));
    outputs(11920) <= layer2_outputs(5114);
    outputs(11921) <= not((layer2_outputs(9740)) xor (layer2_outputs(2895)));
    outputs(11922) <= not((layer2_outputs(1050)) and (layer2_outputs(7164)));
    outputs(11923) <= (layer2_outputs(11875)) or (layer2_outputs(8879));
    outputs(11924) <= not(layer2_outputs(7199));
    outputs(11925) <= layer2_outputs(6602);
    outputs(11926) <= (layer2_outputs(2453)) and (layer2_outputs(2750));
    outputs(11927) <= layer2_outputs(8946);
    outputs(11928) <= not(layer2_outputs(7240));
    outputs(11929) <= not(layer2_outputs(121));
    outputs(11930) <= not((layer2_outputs(273)) or (layer2_outputs(1190)));
    outputs(11931) <= not(layer2_outputs(5797));
    outputs(11932) <= not(layer2_outputs(8660)) or (layer2_outputs(8121));
    outputs(11933) <= layer2_outputs(7997);
    outputs(11934) <= not((layer2_outputs(7802)) or (layer2_outputs(3246)));
    outputs(11935) <= not(layer2_outputs(995));
    outputs(11936) <= not((layer2_outputs(4413)) xor (layer2_outputs(2979)));
    outputs(11937) <= (layer2_outputs(9030)) and not (layer2_outputs(1034));
    outputs(11938) <= layer2_outputs(4981);
    outputs(11939) <= not(layer2_outputs(10336));
    outputs(11940) <= layer2_outputs(3137);
    outputs(11941) <= (layer2_outputs(8954)) and not (layer2_outputs(1163));
    outputs(11942) <= not(layer2_outputs(3588));
    outputs(11943) <= (layer2_outputs(3273)) and not (layer2_outputs(2516));
    outputs(11944) <= not(layer2_outputs(7379));
    outputs(11945) <= layer2_outputs(9135);
    outputs(11946) <= (layer2_outputs(123)) or (layer2_outputs(9336));
    outputs(11947) <= not((layer2_outputs(9305)) xor (layer2_outputs(6489)));
    outputs(11948) <= not((layer2_outputs(10098)) xor (layer2_outputs(12031)));
    outputs(11949) <= not(layer2_outputs(10090));
    outputs(11950) <= not(layer2_outputs(1410)) or (layer2_outputs(6456));
    outputs(11951) <= not(layer2_outputs(4202));
    outputs(11952) <= not((layer2_outputs(2819)) and (layer2_outputs(10828)));
    outputs(11953) <= layer2_outputs(6539);
    outputs(11954) <= (layer2_outputs(10950)) and not (layer2_outputs(10902));
    outputs(11955) <= not(layer2_outputs(10026));
    outputs(11956) <= layer2_outputs(1995);
    outputs(11957) <= not(layer2_outputs(624)) or (layer2_outputs(2251));
    outputs(11958) <= not(layer2_outputs(7499)) or (layer2_outputs(2634));
    outputs(11959) <= (layer2_outputs(7314)) xor (layer2_outputs(3934));
    outputs(11960) <= (layer2_outputs(4738)) and (layer2_outputs(12267));
    outputs(11961) <= layer2_outputs(3570);
    outputs(11962) <= not(layer2_outputs(12095));
    outputs(11963) <= layer2_outputs(785);
    outputs(11964) <= layer2_outputs(11541);
    outputs(11965) <= not(layer2_outputs(10705));
    outputs(11966) <= not((layer2_outputs(7504)) xor (layer2_outputs(11614)));
    outputs(11967) <= not(layer2_outputs(3414)) or (layer2_outputs(8236));
    outputs(11968) <= not(layer2_outputs(5583));
    outputs(11969) <= not((layer2_outputs(4846)) xor (layer2_outputs(3818)));
    outputs(11970) <= (layer2_outputs(5267)) and not (layer2_outputs(11653));
    outputs(11971) <= not(layer2_outputs(10504));
    outputs(11972) <= not(layer2_outputs(65));
    outputs(11973) <= layer2_outputs(12189);
    outputs(11974) <= not(layer2_outputs(5493));
    outputs(11975) <= not((layer2_outputs(5834)) or (layer2_outputs(5404)));
    outputs(11976) <= not(layer2_outputs(6604)) or (layer2_outputs(11558));
    outputs(11977) <= not((layer2_outputs(7201)) xor (layer2_outputs(1113)));
    outputs(11978) <= not((layer2_outputs(660)) and (layer2_outputs(6198)));
    outputs(11979) <= not(layer2_outputs(1996));
    outputs(11980) <= (layer2_outputs(11604)) xor (layer2_outputs(2513));
    outputs(11981) <= layer2_outputs(6010);
    outputs(11982) <= not(layer2_outputs(7759)) or (layer2_outputs(2769));
    outputs(11983) <= layer2_outputs(5448);
    outputs(11984) <= (layer2_outputs(11048)) and (layer2_outputs(6336));
    outputs(11985) <= (layer2_outputs(12)) and not (layer2_outputs(8458));
    outputs(11986) <= layer2_outputs(2189);
    outputs(11987) <= not(layer2_outputs(1875));
    outputs(11988) <= layer2_outputs(884);
    outputs(11989) <= not((layer2_outputs(4226)) or (layer2_outputs(12008)));
    outputs(11990) <= (layer2_outputs(4562)) or (layer2_outputs(1714));
    outputs(11991) <= not(layer2_outputs(2975));
    outputs(11992) <= layer2_outputs(12374);
    outputs(11993) <= (layer2_outputs(9390)) xor (layer2_outputs(9856));
    outputs(11994) <= not(layer2_outputs(7008));
    outputs(11995) <= (layer2_outputs(11813)) xor (layer2_outputs(5169));
    outputs(11996) <= (layer2_outputs(4242)) xor (layer2_outputs(5046));
    outputs(11997) <= not(layer2_outputs(5145));
    outputs(11998) <= (layer2_outputs(12102)) xor (layer2_outputs(5687));
    outputs(11999) <= not(layer2_outputs(9839));
    outputs(12000) <= not(layer2_outputs(5656));
    outputs(12001) <= (layer2_outputs(1830)) xor (layer2_outputs(5123));
    outputs(12002) <= (layer2_outputs(6960)) xor (layer2_outputs(6991));
    outputs(12003) <= (layer2_outputs(8951)) and (layer2_outputs(659));
    outputs(12004) <= (layer2_outputs(3244)) or (layer2_outputs(3577));
    outputs(12005) <= layer2_outputs(5756);
    outputs(12006) <= not(layer2_outputs(8516));
    outputs(12007) <= (layer2_outputs(1075)) or (layer2_outputs(5827));
    outputs(12008) <= not(layer2_outputs(4065));
    outputs(12009) <= layer2_outputs(11421);
    outputs(12010) <= layer2_outputs(10672);
    outputs(12011) <= layer2_outputs(8493);
    outputs(12012) <= not(layer2_outputs(11500));
    outputs(12013) <= layer2_outputs(8591);
    outputs(12014) <= not(layer2_outputs(1691));
    outputs(12015) <= not((layer2_outputs(6622)) xor (layer2_outputs(3662)));
    outputs(12016) <= layer2_outputs(5539);
    outputs(12017) <= not(layer2_outputs(11693));
    outputs(12018) <= (layer2_outputs(11797)) xor (layer2_outputs(372));
    outputs(12019) <= not((layer2_outputs(64)) or (layer2_outputs(6657)));
    outputs(12020) <= not((layer2_outputs(8494)) xor (layer2_outputs(9960)));
    outputs(12021) <= not(layer2_outputs(6016));
    outputs(12022) <= (layer2_outputs(6377)) xor (layer2_outputs(627));
    outputs(12023) <= not(layer2_outputs(10241));
    outputs(12024) <= not(layer2_outputs(2114));
    outputs(12025) <= not(layer2_outputs(9903)) or (layer2_outputs(4508));
    outputs(12026) <= not(layer2_outputs(4345));
    outputs(12027) <= layer2_outputs(12202);
    outputs(12028) <= not(layer2_outputs(6712));
    outputs(12029) <= not((layer2_outputs(8133)) or (layer2_outputs(4384)));
    outputs(12030) <= not(layer2_outputs(7849));
    outputs(12031) <= not((layer2_outputs(2356)) or (layer2_outputs(12682)));
    outputs(12032) <= (layer2_outputs(1125)) xor (layer2_outputs(1618));
    outputs(12033) <= not(layer2_outputs(3907));
    outputs(12034) <= (layer2_outputs(3258)) xor (layer2_outputs(298));
    outputs(12035) <= not(layer2_outputs(4586));
    outputs(12036) <= not(layer2_outputs(940));
    outputs(12037) <= layer2_outputs(8426);
    outputs(12038) <= layer2_outputs(4888);
    outputs(12039) <= not((layer2_outputs(7143)) xor (layer2_outputs(3344)));
    outputs(12040) <= not((layer2_outputs(643)) xor (layer2_outputs(1796)));
    outputs(12041) <= not(layer2_outputs(7516));
    outputs(12042) <= layer2_outputs(9193);
    outputs(12043) <= not((layer2_outputs(5430)) xor (layer2_outputs(3762)));
    outputs(12044) <= not(layer2_outputs(8766));
    outputs(12045) <= layer2_outputs(8981);
    outputs(12046) <= layer2_outputs(878);
    outputs(12047) <= not(layer2_outputs(2439));
    outputs(12048) <= (layer2_outputs(6949)) xor (layer2_outputs(5783));
    outputs(12049) <= layer2_outputs(2360);
    outputs(12050) <= not((layer2_outputs(11138)) and (layer2_outputs(2551)));
    outputs(12051) <= (layer2_outputs(6270)) and (layer2_outputs(8692));
    outputs(12052) <= layer2_outputs(6620);
    outputs(12053) <= (layer2_outputs(9826)) xor (layer2_outputs(4019));
    outputs(12054) <= not(layer2_outputs(12302));
    outputs(12055) <= not(layer2_outputs(10297));
    outputs(12056) <= layer2_outputs(10347);
    outputs(12057) <= not((layer2_outputs(8645)) xor (layer2_outputs(888)));
    outputs(12058) <= not(layer2_outputs(2367));
    outputs(12059) <= (layer2_outputs(6337)) xor (layer2_outputs(8089));
    outputs(12060) <= not(layer2_outputs(3755));
    outputs(12061) <= layer2_outputs(6976);
    outputs(12062) <= not((layer2_outputs(7850)) and (layer2_outputs(2165)));
    outputs(12063) <= layer2_outputs(1312);
    outputs(12064) <= (layer2_outputs(2801)) or (layer2_outputs(3361));
    outputs(12065) <= layer2_outputs(2422);
    outputs(12066) <= layer2_outputs(12773);
    outputs(12067) <= (layer2_outputs(1940)) xor (layer2_outputs(9607));
    outputs(12068) <= layer2_outputs(5261);
    outputs(12069) <= layer2_outputs(8527);
    outputs(12070) <= (layer2_outputs(12244)) xor (layer2_outputs(4259));
    outputs(12071) <= not((layer2_outputs(736)) or (layer2_outputs(11087)));
    outputs(12072) <= not(layer2_outputs(11648));
    outputs(12073) <= not(layer2_outputs(7644));
    outputs(12074) <= layer2_outputs(452);
    outputs(12075) <= not(layer2_outputs(5272));
    outputs(12076) <= not((layer2_outputs(3513)) xor (layer2_outputs(3581)));
    outputs(12077) <= (layer2_outputs(1156)) and (layer2_outputs(2968));
    outputs(12078) <= layer2_outputs(9107);
    outputs(12079) <= (layer2_outputs(2997)) and (layer2_outputs(8462));
    outputs(12080) <= not(layer2_outputs(12025));
    outputs(12081) <= not(layer2_outputs(6820));
    outputs(12082) <= (layer2_outputs(4097)) xor (layer2_outputs(11818));
    outputs(12083) <= (layer2_outputs(9731)) and (layer2_outputs(4916));
    outputs(12084) <= not((layer2_outputs(12777)) xor (layer2_outputs(5292)));
    outputs(12085) <= not(layer2_outputs(11185));
    outputs(12086) <= (layer2_outputs(8121)) and not (layer2_outputs(6118));
    outputs(12087) <= not(layer2_outputs(5530));
    outputs(12088) <= layer2_outputs(936);
    outputs(12089) <= not(layer2_outputs(638)) or (layer2_outputs(1437));
    outputs(12090) <= not((layer2_outputs(2262)) and (layer2_outputs(8281)));
    outputs(12091) <= (layer2_outputs(5320)) xor (layer2_outputs(9526));
    outputs(12092) <= not(layer2_outputs(6743)) or (layer2_outputs(2461));
    outputs(12093) <= layer2_outputs(7318);
    outputs(12094) <= (layer2_outputs(2540)) and not (layer2_outputs(7483));
    outputs(12095) <= (layer2_outputs(5344)) xor (layer2_outputs(2743));
    outputs(12096) <= (layer2_outputs(8496)) xor (layer2_outputs(12546));
    outputs(12097) <= not(layer2_outputs(7216));
    outputs(12098) <= not((layer2_outputs(10055)) xor (layer2_outputs(8241)));
    outputs(12099) <= not((layer2_outputs(9014)) xor (layer2_outputs(755)));
    outputs(12100) <= not((layer2_outputs(10240)) xor (layer2_outputs(4675)));
    outputs(12101) <= not(layer2_outputs(1824));
    outputs(12102) <= (layer2_outputs(728)) and not (layer2_outputs(247));
    outputs(12103) <= not(layer2_outputs(3614));
    outputs(12104) <= layer2_outputs(8260);
    outputs(12105) <= layer2_outputs(5434);
    outputs(12106) <= layer2_outputs(9069);
    outputs(12107) <= layer2_outputs(4371);
    outputs(12108) <= (layer2_outputs(9425)) xor (layer2_outputs(8492));
    outputs(12109) <= not((layer2_outputs(6546)) xor (layer2_outputs(5934)));
    outputs(12110) <= layer2_outputs(12565);
    outputs(12111) <= not(layer2_outputs(5182)) or (layer2_outputs(2662));
    outputs(12112) <= layer2_outputs(5444);
    outputs(12113) <= not(layer2_outputs(6098));
    outputs(12114) <= (layer2_outputs(8834)) and not (layer2_outputs(11985));
    outputs(12115) <= (layer2_outputs(15)) xor (layer2_outputs(7396));
    outputs(12116) <= layer2_outputs(1177);
    outputs(12117) <= layer2_outputs(8343);
    outputs(12118) <= not(layer2_outputs(11095)) or (layer2_outputs(455));
    outputs(12119) <= layer2_outputs(8483);
    outputs(12120) <= not(layer2_outputs(12484));
    outputs(12121) <= layer2_outputs(2963);
    outputs(12122) <= (layer2_outputs(2009)) and (layer2_outputs(12186));
    outputs(12123) <= (layer2_outputs(4173)) xor (layer2_outputs(10285));
    outputs(12124) <= layer2_outputs(7351);
    outputs(12125) <= not(layer2_outputs(5046)) or (layer2_outputs(11015));
    outputs(12126) <= not(layer2_outputs(9548));
    outputs(12127) <= not((layer2_outputs(7220)) xor (layer2_outputs(3922)));
    outputs(12128) <= not((layer2_outputs(2734)) and (layer2_outputs(12356)));
    outputs(12129) <= (layer2_outputs(10764)) and (layer2_outputs(9013));
    outputs(12130) <= not(layer2_outputs(1308));
    outputs(12131) <= (layer2_outputs(12412)) xor (layer2_outputs(4786));
    outputs(12132) <= (layer2_outputs(2108)) xor (layer2_outputs(928));
    outputs(12133) <= layer2_outputs(6804);
    outputs(12134) <= not((layer2_outputs(7679)) and (layer2_outputs(6988)));
    outputs(12135) <= (layer2_outputs(82)) xor (layer2_outputs(7891));
    outputs(12136) <= not((layer2_outputs(5501)) or (layer2_outputs(6582)));
    outputs(12137) <= layer2_outputs(8735);
    outputs(12138) <= layer2_outputs(4602);
    outputs(12139) <= not(layer2_outputs(9571));
    outputs(12140) <= not(layer2_outputs(10974));
    outputs(12141) <= not(layer2_outputs(976));
    outputs(12142) <= (layer2_outputs(10078)) xor (layer2_outputs(7988));
    outputs(12143) <= layer2_outputs(11837);
    outputs(12144) <= (layer2_outputs(11210)) and not (layer2_outputs(12182));
    outputs(12145) <= (layer2_outputs(9660)) xor (layer2_outputs(8896));
    outputs(12146) <= layer2_outputs(680);
    outputs(12147) <= layer2_outputs(6751);
    outputs(12148) <= not(layer2_outputs(1145));
    outputs(12149) <= not((layer2_outputs(7939)) xor (layer2_outputs(4511)));
    outputs(12150) <= not((layer2_outputs(9052)) xor (layer2_outputs(11717)));
    outputs(12151) <= layer2_outputs(3153);
    outputs(12152) <= not(layer2_outputs(7942));
    outputs(12153) <= not(layer2_outputs(11500));
    outputs(12154) <= layer2_outputs(7502);
    outputs(12155) <= not(layer2_outputs(4115));
    outputs(12156) <= not(layer2_outputs(8233));
    outputs(12157) <= not(layer2_outputs(5084));
    outputs(12158) <= not(layer2_outputs(9356));
    outputs(12159) <= layer2_outputs(3277);
    outputs(12160) <= not((layer2_outputs(8832)) xor (layer2_outputs(10432)));
    outputs(12161) <= (layer2_outputs(3543)) xor (layer2_outputs(8366));
    outputs(12162) <= layer2_outputs(7230);
    outputs(12163) <= not(layer2_outputs(9584));
    outputs(12164) <= (layer2_outputs(11760)) and (layer2_outputs(3239));
    outputs(12165) <= not(layer2_outputs(2073));
    outputs(12166) <= not(layer2_outputs(6516));
    outputs(12167) <= (layer2_outputs(6399)) xor (layer2_outputs(123));
    outputs(12168) <= (layer2_outputs(5171)) xor (layer2_outputs(12115));
    outputs(12169) <= not(layer2_outputs(5801));
    outputs(12170) <= not((layer2_outputs(6402)) xor (layer2_outputs(475)));
    outputs(12171) <= (layer2_outputs(1092)) xor (layer2_outputs(7801));
    outputs(12172) <= layer2_outputs(10801);
    outputs(12173) <= not(layer2_outputs(4386));
    outputs(12174) <= layer2_outputs(2609);
    outputs(12175) <= (layer2_outputs(880)) and not (layer2_outputs(10510));
    outputs(12176) <= layer2_outputs(3059);
    outputs(12177) <= not((layer2_outputs(5829)) xor (layer2_outputs(5342)));
    outputs(12178) <= layer2_outputs(5959);
    outputs(12179) <= not(layer2_outputs(6541));
    outputs(12180) <= not(layer2_outputs(3529));
    outputs(12181) <= layer2_outputs(1073);
    outputs(12182) <= (layer2_outputs(6993)) and not (layer2_outputs(6799));
    outputs(12183) <= not(layer2_outputs(4660));
    outputs(12184) <= '1';
    outputs(12185) <= layer2_outputs(4775);
    outputs(12186) <= (layer2_outputs(11494)) and (layer2_outputs(3923));
    outputs(12187) <= layer2_outputs(1874);
    outputs(12188) <= layer2_outputs(5597);
    outputs(12189) <= not(layer2_outputs(294));
    outputs(12190) <= not((layer2_outputs(3952)) or (layer2_outputs(3219)));
    outputs(12191) <= layer2_outputs(3287);
    outputs(12192) <= not(layer2_outputs(9644));
    outputs(12193) <= not(layer2_outputs(4637));
    outputs(12194) <= (layer2_outputs(3972)) or (layer2_outputs(10099));
    outputs(12195) <= not((layer2_outputs(10895)) or (layer2_outputs(1130)));
    outputs(12196) <= not((layer2_outputs(1203)) xor (layer2_outputs(218)));
    outputs(12197) <= not((layer2_outputs(5347)) xor (layer2_outputs(10055)));
    outputs(12198) <= not((layer2_outputs(6856)) xor (layer2_outputs(5376)));
    outputs(12199) <= not((layer2_outputs(5009)) xor (layer2_outputs(8543)));
    outputs(12200) <= (layer2_outputs(7705)) xor (layer2_outputs(7572));
    outputs(12201) <= not((layer2_outputs(11846)) or (layer2_outputs(10615)));
    outputs(12202) <= not((layer2_outputs(7980)) and (layer2_outputs(11925)));
    outputs(12203) <= not(layer2_outputs(6817));
    outputs(12204) <= not(layer2_outputs(10711));
    outputs(12205) <= layer2_outputs(10371);
    outputs(12206) <= not((layer2_outputs(10268)) xor (layer2_outputs(6561)));
    outputs(12207) <= layer2_outputs(2270);
    outputs(12208) <= (layer2_outputs(7960)) and not (layer2_outputs(4499));
    outputs(12209) <= (layer2_outputs(1812)) xor (layer2_outputs(144));
    outputs(12210) <= not(layer2_outputs(10388));
    outputs(12211) <= not(layer2_outputs(9095));
    outputs(12212) <= (layer2_outputs(9568)) xor (layer2_outputs(12274));
    outputs(12213) <= layer2_outputs(7605);
    outputs(12214) <= not(layer2_outputs(12180));
    outputs(12215) <= not(layer2_outputs(5003)) or (layer2_outputs(535));
    outputs(12216) <= layer2_outputs(3919);
    outputs(12217) <= not(layer2_outputs(5451)) or (layer2_outputs(4101));
    outputs(12218) <= not((layer2_outputs(1683)) xor (layer2_outputs(7669)));
    outputs(12219) <= not((layer2_outputs(8803)) xor (layer2_outputs(10799)));
    outputs(12220) <= not(layer2_outputs(6420)) or (layer2_outputs(10285));
    outputs(12221) <= layer2_outputs(6312);
    outputs(12222) <= (layer2_outputs(3130)) and not (layer2_outputs(9110));
    outputs(12223) <= not(layer2_outputs(6896));
    outputs(12224) <= not(layer2_outputs(1463));
    outputs(12225) <= (layer2_outputs(8242)) and not (layer2_outputs(7099));
    outputs(12226) <= layer2_outputs(1289);
    outputs(12227) <= layer2_outputs(10264);
    outputs(12228) <= (layer2_outputs(4954)) and not (layer2_outputs(860));
    outputs(12229) <= not(layer2_outputs(2020));
    outputs(12230) <= layer2_outputs(12414);
    outputs(12231) <= (layer2_outputs(9431)) and (layer2_outputs(7814));
    outputs(12232) <= not(layer2_outputs(6604)) or (layer2_outputs(8096));
    outputs(12233) <= (layer2_outputs(3826)) and not (layer2_outputs(1196));
    outputs(12234) <= not(layer2_outputs(6667));
    outputs(12235) <= not(layer2_outputs(6351));
    outputs(12236) <= not((layer2_outputs(7023)) or (layer2_outputs(10173)));
    outputs(12237) <= (layer2_outputs(11567)) xor (layer2_outputs(2075));
    outputs(12238) <= not((layer2_outputs(6855)) xor (layer2_outputs(4476)));
    outputs(12239) <= not((layer2_outputs(9980)) and (layer2_outputs(3635)));
    outputs(12240) <= not(layer2_outputs(5573));
    outputs(12241) <= not(layer2_outputs(11583));
    outputs(12242) <= not(layer2_outputs(10935));
    outputs(12243) <= not(layer2_outputs(10168));
    outputs(12244) <= (layer2_outputs(11535)) xor (layer2_outputs(1226));
    outputs(12245) <= (layer2_outputs(10279)) and not (layer2_outputs(2146));
    outputs(12246) <= layer2_outputs(9645);
    outputs(12247) <= (layer2_outputs(9205)) and not (layer2_outputs(1162));
    outputs(12248) <= not(layer2_outputs(2913));
    outputs(12249) <= layer2_outputs(9717);
    outputs(12250) <= not(layer2_outputs(7914));
    outputs(12251) <= not(layer2_outputs(11307));
    outputs(12252) <= layer2_outputs(4773);
    outputs(12253) <= not(layer2_outputs(9862));
    outputs(12254) <= layer2_outputs(7029);
    outputs(12255) <= layer2_outputs(4265);
    outputs(12256) <= (layer2_outputs(975)) xor (layer2_outputs(5670));
    outputs(12257) <= (layer2_outputs(5335)) xor (layer2_outputs(4280));
    outputs(12258) <= layer2_outputs(4);
    outputs(12259) <= layer2_outputs(4587);
    outputs(12260) <= layer2_outputs(5614);
    outputs(12261) <= not(layer2_outputs(1038));
    outputs(12262) <= not(layer2_outputs(10913));
    outputs(12263) <= not(layer2_outputs(2401));
    outputs(12264) <= not(layer2_outputs(2960));
    outputs(12265) <= (layer2_outputs(4361)) xor (layer2_outputs(6713));
    outputs(12266) <= not(layer2_outputs(10967));
    outputs(12267) <= not(layer2_outputs(5285));
    outputs(12268) <= (layer2_outputs(12413)) and not (layer2_outputs(12419));
    outputs(12269) <= not(layer2_outputs(5762));
    outputs(12270) <= layer2_outputs(4790);
    outputs(12271) <= layer2_outputs(4923);
    outputs(12272) <= (layer2_outputs(9662)) xor (layer2_outputs(3123));
    outputs(12273) <= layer2_outputs(10137);
    outputs(12274) <= layer2_outputs(386);
    outputs(12275) <= layer2_outputs(979);
    outputs(12276) <= layer2_outputs(8476);
    outputs(12277) <= (layer2_outputs(4827)) xor (layer2_outputs(1728));
    outputs(12278) <= not(layer2_outputs(3502));
    outputs(12279) <= layer2_outputs(3408);
    outputs(12280) <= not(layer2_outputs(2250));
    outputs(12281) <= not((layer2_outputs(11332)) xor (layer2_outputs(11708)));
    outputs(12282) <= layer2_outputs(4799);
    outputs(12283) <= not(layer2_outputs(1890));
    outputs(12284) <= not((layer2_outputs(3330)) or (layer2_outputs(6869)));
    outputs(12285) <= (layer2_outputs(3013)) xor (layer2_outputs(11617));
    outputs(12286) <= not(layer2_outputs(10192));
    outputs(12287) <= layer2_outputs(3509);
    outputs(12288) <= not(layer2_outputs(9191));
    outputs(12289) <= (layer2_outputs(956)) xor (layer2_outputs(10551));
    outputs(12290) <= not((layer2_outputs(8651)) xor (layer2_outputs(1434)));
    outputs(12291) <= layer2_outputs(8243);
    outputs(12292) <= (layer2_outputs(5643)) xor (layer2_outputs(7698));
    outputs(12293) <= not((layer2_outputs(10197)) xor (layer2_outputs(7844)));
    outputs(12294) <= layer2_outputs(11415);
    outputs(12295) <= not(layer2_outputs(11017));
    outputs(12296) <= layer2_outputs(4141);
    outputs(12297) <= not(layer2_outputs(10468));
    outputs(12298) <= not(layer2_outputs(5743));
    outputs(12299) <= layer2_outputs(9289);
    outputs(12300) <= not((layer2_outputs(2079)) or (layer2_outputs(10141)));
    outputs(12301) <= layer2_outputs(403);
    outputs(12302) <= not(layer2_outputs(10864));
    outputs(12303) <= (layer2_outputs(7120)) xor (layer2_outputs(3004));
    outputs(12304) <= layer2_outputs(10186);
    outputs(12305) <= not(layer2_outputs(917));
    outputs(12306) <= (layer2_outputs(11265)) xor (layer2_outputs(7866));
    outputs(12307) <= (layer2_outputs(3920)) xor (layer2_outputs(11460));
    outputs(12308) <= (layer2_outputs(8223)) and not (layer2_outputs(9171));
    outputs(12309) <= not(layer2_outputs(3985));
    outputs(12310) <= (layer2_outputs(2766)) xor (layer2_outputs(9072));
    outputs(12311) <= layer2_outputs(5304);
    outputs(12312) <= (layer2_outputs(11791)) xor (layer2_outputs(12177));
    outputs(12313) <= not((layer2_outputs(1110)) xor (layer2_outputs(2977)));
    outputs(12314) <= not((layer2_outputs(2895)) xor (layer2_outputs(1453)));
    outputs(12315) <= (layer2_outputs(9604)) and not (layer2_outputs(6973));
    outputs(12316) <= not((layer2_outputs(3659)) xor (layer2_outputs(1084)));
    outputs(12317) <= (layer2_outputs(5593)) xor (layer2_outputs(3708));
    outputs(12318) <= layer2_outputs(7457);
    outputs(12319) <= not((layer2_outputs(8756)) or (layer2_outputs(10401)));
    outputs(12320) <= not((layer2_outputs(9804)) xor (layer2_outputs(1990)));
    outputs(12321) <= layer2_outputs(7959);
    outputs(12322) <= layer2_outputs(12519);
    outputs(12323) <= (layer2_outputs(8839)) xor (layer2_outputs(1063));
    outputs(12324) <= not(layer2_outputs(71));
    outputs(12325) <= not(layer2_outputs(6750));
    outputs(12326) <= not(layer2_outputs(12728)) or (layer2_outputs(7737));
    outputs(12327) <= not((layer2_outputs(2283)) xor (layer2_outputs(154)));
    outputs(12328) <= not(layer2_outputs(1755));
    outputs(12329) <= layer2_outputs(2655);
    outputs(12330) <= not(layer2_outputs(11193));
    outputs(12331) <= layer2_outputs(12788);
    outputs(12332) <= not((layer2_outputs(6578)) or (layer2_outputs(4741)));
    outputs(12333) <= not((layer2_outputs(5071)) xor (layer2_outputs(9343)));
    outputs(12334) <= not(layer2_outputs(8026));
    outputs(12335) <= not(layer2_outputs(3336)) or (layer2_outputs(6395));
    outputs(12336) <= (layer2_outputs(4320)) and (layer2_outputs(6377));
    outputs(12337) <= not(layer2_outputs(11143)) or (layer2_outputs(12479));
    outputs(12338) <= layer2_outputs(12756);
    outputs(12339) <= not((layer2_outputs(7573)) or (layer2_outputs(6151)));
    outputs(12340) <= layer2_outputs(6393);
    outputs(12341) <= (layer2_outputs(11245)) or (layer2_outputs(1261));
    outputs(12342) <= layer2_outputs(7664);
    outputs(12343) <= layer2_outputs(1144);
    outputs(12344) <= not(layer2_outputs(6036));
    outputs(12345) <= layer2_outputs(2856);
    outputs(12346) <= layer2_outputs(11424);
    outputs(12347) <= not(layer2_outputs(7375));
    outputs(12348) <= not((layer2_outputs(3183)) and (layer2_outputs(882)));
    outputs(12349) <= (layer2_outputs(8053)) and (layer2_outputs(2109));
    outputs(12350) <= (layer2_outputs(9316)) xor (layer2_outputs(2462));
    outputs(12351) <= (layer2_outputs(58)) xor (layer2_outputs(6158));
    outputs(12352) <= layer2_outputs(3127);
    outputs(12353) <= layer2_outputs(3480);
    outputs(12354) <= not(layer2_outputs(7715));
    outputs(12355) <= not((layer2_outputs(10252)) xor (layer2_outputs(6457)));
    outputs(12356) <= not((layer2_outputs(9596)) xor (layer2_outputs(9304)));
    outputs(12357) <= layer2_outputs(11780);
    outputs(12358) <= layer2_outputs(10921);
    outputs(12359) <= not(layer2_outputs(482));
    outputs(12360) <= not(layer2_outputs(12611));
    outputs(12361) <= layer2_outputs(4070);
    outputs(12362) <= layer2_outputs(3093);
    outputs(12363) <= not(layer2_outputs(1738));
    outputs(12364) <= not(layer2_outputs(10931));
    outputs(12365) <= layer2_outputs(139);
    outputs(12366) <= (layer2_outputs(11053)) xor (layer2_outputs(3115));
    outputs(12367) <= layer2_outputs(6628);
    outputs(12368) <= not(layer2_outputs(12158)) or (layer2_outputs(951));
    outputs(12369) <= layer2_outputs(4407);
    outputs(12370) <= not(layer2_outputs(262)) or (layer2_outputs(5300));
    outputs(12371) <= not((layer2_outputs(4702)) and (layer2_outputs(8538)));
    outputs(12372) <= layer2_outputs(5942);
    outputs(12373) <= layer2_outputs(10555);
    outputs(12374) <= (layer2_outputs(2781)) xor (layer2_outputs(56));
    outputs(12375) <= not((layer2_outputs(9417)) xor (layer2_outputs(6917)));
    outputs(12376) <= (layer2_outputs(5479)) xor (layer2_outputs(4229));
    outputs(12377) <= layer2_outputs(11814);
    outputs(12378) <= (layer2_outputs(9070)) xor (layer2_outputs(6268));
    outputs(12379) <= layer2_outputs(5100);
    outputs(12380) <= not((layer2_outputs(3410)) xor (layer2_outputs(12187)));
    outputs(12381) <= not((layer2_outputs(5318)) and (layer2_outputs(4314)));
    outputs(12382) <= (layer2_outputs(7472)) and not (layer2_outputs(10036));
    outputs(12383) <= layer2_outputs(4948);
    outputs(12384) <= not(layer2_outputs(9601));
    outputs(12385) <= not(layer2_outputs(6464));
    outputs(12386) <= layer2_outputs(7108);
    outputs(12387) <= (layer2_outputs(1239)) xor (layer2_outputs(1458));
    outputs(12388) <= not(layer2_outputs(328));
    outputs(12389) <= layer2_outputs(7725);
    outputs(12390) <= not((layer2_outputs(12344)) xor (layer2_outputs(4669)));
    outputs(12391) <= (layer2_outputs(11461)) or (layer2_outputs(1035));
    outputs(12392) <= not(layer2_outputs(7406));
    outputs(12393) <= not(layer2_outputs(7203)) or (layer2_outputs(5385));
    outputs(12394) <= (layer2_outputs(3039)) xor (layer2_outputs(12531));
    outputs(12395) <= layer2_outputs(12111);
    outputs(12396) <= not((layer2_outputs(8932)) xor (layer2_outputs(2797)));
    outputs(12397) <= not(layer2_outputs(7047));
    outputs(12398) <= layer2_outputs(7523);
    outputs(12399) <= not((layer2_outputs(12209)) xor (layer2_outputs(11304)));
    outputs(12400) <= not(layer2_outputs(1967));
    outputs(12401) <= not((layer2_outputs(1355)) xor (layer2_outputs(482)));
    outputs(12402) <= not(layer2_outputs(7357));
    outputs(12403) <= not((layer2_outputs(12782)) or (layer2_outputs(4115)));
    outputs(12404) <= not(layer2_outputs(10410));
    outputs(12405) <= not(layer2_outputs(6069));
    outputs(12406) <= layer2_outputs(9054);
    outputs(12407) <= not(layer2_outputs(3957));
    outputs(12408) <= not((layer2_outputs(1036)) xor (layer2_outputs(6184)));
    outputs(12409) <= (layer2_outputs(4277)) or (layer2_outputs(142));
    outputs(12410) <= not((layer2_outputs(11216)) xor (layer2_outputs(11616)));
    outputs(12411) <= not((layer2_outputs(11504)) xor (layer2_outputs(10558)));
    outputs(12412) <= layer2_outputs(6880);
    outputs(12413) <= not(layer2_outputs(27)) or (layer2_outputs(11699));
    outputs(12414) <= not((layer2_outputs(6226)) or (layer2_outputs(10538)));
    outputs(12415) <= not((layer2_outputs(6974)) xor (layer2_outputs(5581)));
    outputs(12416) <= not((layer2_outputs(6943)) xor (layer2_outputs(9360)));
    outputs(12417) <= layer2_outputs(9994);
    outputs(12418) <= not(layer2_outputs(6153));
    outputs(12419) <= not(layer2_outputs(9329));
    outputs(12420) <= (layer2_outputs(9565)) xor (layer2_outputs(563));
    outputs(12421) <= layer2_outputs(12373);
    outputs(12422) <= not(layer2_outputs(513));
    outputs(12423) <= layer2_outputs(5315);
    outputs(12424) <= not(layer2_outputs(8132));
    outputs(12425) <= not(layer2_outputs(4544));
    outputs(12426) <= not(layer2_outputs(8075));
    outputs(12427) <= not((layer2_outputs(514)) xor (layer2_outputs(5849)));
    outputs(12428) <= not(layer2_outputs(1977));
    outputs(12429) <= not(layer2_outputs(4304));
    outputs(12430) <= not(layer2_outputs(1067));
    outputs(12431) <= not(layer2_outputs(180)) or (layer2_outputs(4735));
    outputs(12432) <= (layer2_outputs(10685)) and (layer2_outputs(9949));
    outputs(12433) <= (layer2_outputs(7308)) and (layer2_outputs(7317));
    outputs(12434) <= not((layer2_outputs(3177)) or (layer2_outputs(10710)));
    outputs(12435) <= not((layer2_outputs(9247)) xor (layer2_outputs(255)));
    outputs(12436) <= not((layer2_outputs(3563)) and (layer2_outputs(2094)));
    outputs(12437) <= layer2_outputs(3326);
    outputs(12438) <= layer2_outputs(11875);
    outputs(12439) <= not(layer2_outputs(5549)) or (layer2_outputs(11058));
    outputs(12440) <= not(layer2_outputs(2059));
    outputs(12441) <= not(layer2_outputs(12509));
    outputs(12442) <= not(layer2_outputs(10096)) or (layer2_outputs(973));
    outputs(12443) <= (layer2_outputs(5439)) xor (layer2_outputs(8682));
    outputs(12444) <= not(layer2_outputs(4962));
    outputs(12445) <= not((layer2_outputs(10844)) xor (layer2_outputs(5591)));
    outputs(12446) <= layer2_outputs(7873);
    outputs(12447) <= layer2_outputs(7605);
    outputs(12448) <= not(layer2_outputs(9299));
    outputs(12449) <= not(layer2_outputs(2573));
    outputs(12450) <= layer2_outputs(1764);
    outputs(12451) <= (layer2_outputs(5962)) and not (layer2_outputs(2029));
    outputs(12452) <= layer2_outputs(7554);
    outputs(12453) <= not(layer2_outputs(11329));
    outputs(12454) <= layer2_outputs(2241);
    outputs(12455) <= layer2_outputs(5804);
    outputs(12456) <= layer2_outputs(12088);
    outputs(12457) <= layer2_outputs(1520);
    outputs(12458) <= not(layer2_outputs(5977));
    outputs(12459) <= (layer2_outputs(6347)) or (layer2_outputs(8196));
    outputs(12460) <= not((layer2_outputs(9075)) xor (layer2_outputs(7888)));
    outputs(12461) <= not(layer2_outputs(4724));
    outputs(12462) <= not(layer2_outputs(5049));
    outputs(12463) <= (layer2_outputs(8815)) and not (layer2_outputs(4715));
    outputs(12464) <= layer2_outputs(6627);
    outputs(12465) <= (layer2_outputs(6214)) and not (layer2_outputs(8883));
    outputs(12466) <= (layer2_outputs(3484)) xor (layer2_outputs(6196));
    outputs(12467) <= (layer2_outputs(10908)) xor (layer2_outputs(6684));
    outputs(12468) <= not(layer2_outputs(5625));
    outputs(12469) <= not(layer2_outputs(10933));
    outputs(12470) <= not(layer2_outputs(8676));
    outputs(12471) <= (layer2_outputs(5865)) or (layer2_outputs(1211));
    outputs(12472) <= not(layer2_outputs(3312));
    outputs(12473) <= layer2_outputs(3239);
    outputs(12474) <= not(layer2_outputs(6465));
    outputs(12475) <= not(layer2_outputs(12169));
    outputs(12476) <= not((layer2_outputs(525)) or (layer2_outputs(12524)));
    outputs(12477) <= not(layer2_outputs(9779));
    outputs(12478) <= (layer2_outputs(70)) xor (layer2_outputs(4179));
    outputs(12479) <= layer2_outputs(7374);
    outputs(12480) <= not((layer2_outputs(8669)) xor (layer2_outputs(2729)));
    outputs(12481) <= layer2_outputs(8723);
    outputs(12482) <= not(layer2_outputs(601)) or (layer2_outputs(11120));
    outputs(12483) <= layer2_outputs(6335);
    outputs(12484) <= (layer2_outputs(9388)) xor (layer2_outputs(2152));
    outputs(12485) <= (layer2_outputs(8113)) xor (layer2_outputs(12028));
    outputs(12486) <= layer2_outputs(538);
    outputs(12487) <= not(layer2_outputs(3479)) or (layer2_outputs(12392));
    outputs(12488) <= (layer2_outputs(8175)) xor (layer2_outputs(423));
    outputs(12489) <= not(layer2_outputs(12096)) or (layer2_outputs(7868));
    outputs(12490) <= not(layer2_outputs(1630));
    outputs(12491) <= layer2_outputs(3276);
    outputs(12492) <= layer2_outputs(10531);
    outputs(12493) <= not(layer2_outputs(4724)) or (layer2_outputs(11072));
    outputs(12494) <= not(layer2_outputs(3286));
    outputs(12495) <= (layer2_outputs(3551)) and not (layer2_outputs(10060));
    outputs(12496) <= layer2_outputs(4709);
    outputs(12497) <= (layer2_outputs(2340)) xor (layer2_outputs(5633));
    outputs(12498) <= (layer2_outputs(4640)) xor (layer2_outputs(7652));
    outputs(12499) <= (layer2_outputs(6962)) and not (layer2_outputs(3934));
    outputs(12500) <= not(layer2_outputs(2282));
    outputs(12501) <= not(layer2_outputs(3049));
    outputs(12502) <= layer2_outputs(3509);
    outputs(12503) <= (layer2_outputs(10893)) and not (layer2_outputs(4983));
    outputs(12504) <= not(layer2_outputs(7361));
    outputs(12505) <= not(layer2_outputs(11082));
    outputs(12506) <= (layer2_outputs(10787)) and (layer2_outputs(12016));
    outputs(12507) <= layer2_outputs(9938);
    outputs(12508) <= not(layer2_outputs(9987));
    outputs(12509) <= (layer2_outputs(8716)) and not (layer2_outputs(332));
    outputs(12510) <= not(layer2_outputs(1062));
    outputs(12511) <= layer2_outputs(4432);
    outputs(12512) <= not(layer2_outputs(2552));
    outputs(12513) <= layer2_outputs(9064);
    outputs(12514) <= not(layer2_outputs(9969));
    outputs(12515) <= (layer2_outputs(9831)) xor (layer2_outputs(2629));
    outputs(12516) <= layer2_outputs(10164);
    outputs(12517) <= not((layer2_outputs(1091)) xor (layer2_outputs(5642)));
    outputs(12518) <= not(layer2_outputs(7926)) or (layer2_outputs(9625));
    outputs(12519) <= not((layer2_outputs(12063)) and (layer2_outputs(3770)));
    outputs(12520) <= not(layer2_outputs(3699));
    outputs(12521) <= (layer2_outputs(6369)) and not (layer2_outputs(9752));
    outputs(12522) <= not(layer2_outputs(1992)) or (layer2_outputs(462));
    outputs(12523) <= not((layer2_outputs(6884)) xor (layer2_outputs(6724)));
    outputs(12524) <= (layer2_outputs(4516)) and (layer2_outputs(10210));
    outputs(12525) <= not((layer2_outputs(12328)) or (layer2_outputs(10001)));
    outputs(12526) <= (layer2_outputs(2845)) xor (layer2_outputs(6635));
    outputs(12527) <= not(layer2_outputs(1260));
    outputs(12528) <= layer2_outputs(1500);
    outputs(12529) <= not((layer2_outputs(11385)) xor (layer2_outputs(11406)));
    outputs(12530) <= (layer2_outputs(10615)) xor (layer2_outputs(4365));
    outputs(12531) <= layer2_outputs(6300);
    outputs(12532) <= layer2_outputs(1501);
    outputs(12533) <= (layer2_outputs(3144)) or (layer2_outputs(309));
    outputs(12534) <= (layer2_outputs(11057)) xor (layer2_outputs(9836));
    outputs(12535) <= layer2_outputs(1207);
    outputs(12536) <= not((layer2_outputs(299)) xor (layer2_outputs(6100)));
    outputs(12537) <= (layer2_outputs(179)) and (layer2_outputs(9346));
    outputs(12538) <= not(layer2_outputs(3469));
    outputs(12539) <= (layer2_outputs(2103)) or (layer2_outputs(777));
    outputs(12540) <= not(layer2_outputs(5397));
    outputs(12541) <= layer2_outputs(7131);
    outputs(12542) <= layer2_outputs(1721);
    outputs(12543) <= not((layer2_outputs(4581)) xor (layer2_outputs(5654)));
    outputs(12544) <= (layer2_outputs(10915)) and (layer2_outputs(5948));
    outputs(12545) <= (layer2_outputs(6169)) xor (layer2_outputs(12212));
    outputs(12546) <= layer2_outputs(5436);
    outputs(12547) <= not((layer2_outputs(11404)) xor (layer2_outputs(6219)));
    outputs(12548) <= (layer2_outputs(692)) and not (layer2_outputs(10142));
    outputs(12549) <= not((layer2_outputs(1029)) and (layer2_outputs(5278)));
    outputs(12550) <= not(layer2_outputs(10139));
    outputs(12551) <= not(layer2_outputs(7239));
    outputs(12552) <= layer2_outputs(3290);
    outputs(12553) <= not((layer2_outputs(3056)) and (layer2_outputs(4300)));
    outputs(12554) <= not(layer2_outputs(716));
    outputs(12555) <= not((layer2_outputs(7555)) xor (layer2_outputs(12205)));
    outputs(12556) <= not((layer2_outputs(620)) xor (layer2_outputs(9892)));
    outputs(12557) <= (layer2_outputs(3184)) xor (layer2_outputs(4630));
    outputs(12558) <= not((layer2_outputs(8248)) xor (layer2_outputs(8460)));
    outputs(12559) <= not(layer2_outputs(2608));
    outputs(12560) <= not((layer2_outputs(2859)) xor (layer2_outputs(4364)));
    outputs(12561) <= not((layer2_outputs(10145)) xor (layer2_outputs(11263)));
    outputs(12562) <= not((layer2_outputs(11636)) xor (layer2_outputs(2242)));
    outputs(12563) <= not(layer2_outputs(11382));
    outputs(12564) <= layer2_outputs(7834);
    outputs(12565) <= layer2_outputs(2406);
    outputs(12566) <= not((layer2_outputs(548)) or (layer2_outputs(5843)));
    outputs(12567) <= (layer2_outputs(2809)) and (layer2_outputs(10207));
    outputs(12568) <= not(layer2_outputs(7281));
    outputs(12569) <= (layer2_outputs(8239)) xor (layer2_outputs(1048));
    outputs(12570) <= layer2_outputs(7295);
    outputs(12571) <= layer2_outputs(7324);
    outputs(12572) <= not(layer2_outputs(11753));
    outputs(12573) <= (layer2_outputs(1157)) and not (layer2_outputs(10928));
    outputs(12574) <= not((layer2_outputs(1794)) and (layer2_outputs(404)));
    outputs(12575) <= not(layer2_outputs(1843));
    outputs(12576) <= not((layer2_outputs(4071)) xor (layer2_outputs(8762)));
    outputs(12577) <= not(layer2_outputs(10785));
    outputs(12578) <= not(layer2_outputs(408));
    outputs(12579) <= layer2_outputs(11021);
    outputs(12580) <= (layer2_outputs(7141)) xor (layer2_outputs(12640));
    outputs(12581) <= not(layer2_outputs(2681));
    outputs(12582) <= layer2_outputs(3057);
    outputs(12583) <= not((layer2_outputs(8608)) xor (layer2_outputs(6503)));
    outputs(12584) <= not((layer2_outputs(7461)) xor (layer2_outputs(2137)));
    outputs(12585) <= (layer2_outputs(349)) xor (layer2_outputs(1734));
    outputs(12586) <= (layer2_outputs(3626)) and (layer2_outputs(1721));
    outputs(12587) <= not(layer2_outputs(7117));
    outputs(12588) <= (layer2_outputs(7170)) and not (layer2_outputs(11512));
    outputs(12589) <= (layer2_outputs(7387)) or (layer2_outputs(6713));
    outputs(12590) <= not((layer2_outputs(9959)) xor (layer2_outputs(6426)));
    outputs(12591) <= layer2_outputs(7524);
    outputs(12592) <= (layer2_outputs(12553)) and not (layer2_outputs(9275));
    outputs(12593) <= not((layer2_outputs(5626)) and (layer2_outputs(4064)));
    outputs(12594) <= not((layer2_outputs(12632)) xor (layer2_outputs(3125)));
    outputs(12595) <= not(layer2_outputs(7396));
    outputs(12596) <= not(layer2_outputs(8157));
    outputs(12597) <= (layer2_outputs(650)) xor (layer2_outputs(6749));
    outputs(12598) <= not(layer2_outputs(9356));
    outputs(12599) <= (layer2_outputs(3531)) xor (layer2_outputs(10346));
    outputs(12600) <= layer2_outputs(8816);
    outputs(12601) <= (layer2_outputs(5648)) and not (layer2_outputs(3598));
    outputs(12602) <= not(layer2_outputs(2970));
    outputs(12603) <= not((layer2_outputs(5750)) or (layer2_outputs(4266)));
    outputs(12604) <= layer2_outputs(4555);
    outputs(12605) <= not(layer2_outputs(3672));
    outputs(12606) <= not(layer2_outputs(824));
    outputs(12607) <= not((layer2_outputs(602)) and (layer2_outputs(5075)));
    outputs(12608) <= (layer2_outputs(1865)) xor (layer2_outputs(7332));
    outputs(12609) <= (layer2_outputs(7885)) xor (layer2_outputs(780));
    outputs(12610) <= layer2_outputs(12241);
    outputs(12611) <= not((layer2_outputs(5623)) xor (layer2_outputs(11301)));
    outputs(12612) <= layer2_outputs(7848);
    outputs(12613) <= (layer2_outputs(8056)) and not (layer2_outputs(5403));
    outputs(12614) <= not(layer2_outputs(8509));
    outputs(12615) <= layer2_outputs(4096);
    outputs(12616) <= (layer2_outputs(1068)) and not (layer2_outputs(9414));
    outputs(12617) <= (layer2_outputs(8240)) xor (layer2_outputs(5252));
    outputs(12618) <= layer2_outputs(402);
    outputs(12619) <= layer2_outputs(10067);
    outputs(12620) <= not((layer2_outputs(8027)) or (layer2_outputs(11498)));
    outputs(12621) <= (layer2_outputs(12654)) xor (layer2_outputs(10999));
    outputs(12622) <= layer2_outputs(667);
    outputs(12623) <= not(layer2_outputs(4042));
    outputs(12624) <= not((layer2_outputs(9966)) xor (layer2_outputs(6518)));
    outputs(12625) <= not(layer2_outputs(401));
    outputs(12626) <= not(layer2_outputs(804));
    outputs(12627) <= not(layer2_outputs(11993));
    outputs(12628) <= layer2_outputs(2374);
    outputs(12629) <= layer2_outputs(6997);
    outputs(12630) <= (layer2_outputs(2178)) xor (layer2_outputs(9115));
    outputs(12631) <= layer2_outputs(11911);
    outputs(12632) <= not((layer2_outputs(1661)) xor (layer2_outputs(11230)));
    outputs(12633) <= (layer2_outputs(872)) and not (layer2_outputs(5683));
    outputs(12634) <= (layer2_outputs(8022)) xor (layer2_outputs(1407));
    outputs(12635) <= not((layer2_outputs(11981)) xor (layer2_outputs(12054)));
    outputs(12636) <= (layer2_outputs(9469)) and not (layer2_outputs(9133));
    outputs(12637) <= not(layer2_outputs(248)) or (layer2_outputs(8996));
    outputs(12638) <= (layer2_outputs(7258)) and (layer2_outputs(3417));
    outputs(12639) <= layer2_outputs(9380);
    outputs(12640) <= layer2_outputs(6962);
    outputs(12641) <= not(layer2_outputs(7781)) or (layer2_outputs(8053));
    outputs(12642) <= not((layer2_outputs(10658)) xor (layer2_outputs(3477)));
    outputs(12643) <= not((layer2_outputs(8648)) xor (layer2_outputs(6514)));
    outputs(12644) <= (layer2_outputs(366)) and not (layer2_outputs(12391));
    outputs(12645) <= not((layer2_outputs(2547)) or (layer2_outputs(3736)));
    outputs(12646) <= not(layer2_outputs(157));
    outputs(12647) <= not(layer2_outputs(2306));
    outputs(12648) <= layer2_outputs(8292);
    outputs(12649) <= (layer2_outputs(3006)) and not (layer2_outputs(12333));
    outputs(12650) <= not((layer2_outputs(12772)) xor (layer2_outputs(2427)));
    outputs(12651) <= not(layer2_outputs(12310));
    outputs(12652) <= not((layer2_outputs(11908)) xor (layer2_outputs(5537)));
    outputs(12653) <= not(layer2_outputs(2670));
    outputs(12654) <= layer2_outputs(10276);
    outputs(12655) <= not(layer2_outputs(8183));
    outputs(12656) <= (layer2_outputs(7513)) xor (layer2_outputs(4940));
    outputs(12657) <= layer2_outputs(1823);
    outputs(12658) <= (layer2_outputs(11810)) xor (layer2_outputs(11214));
    outputs(12659) <= (layer2_outputs(3014)) xor (layer2_outputs(5130));
    outputs(12660) <= not(layer2_outputs(250));
    outputs(12661) <= (layer2_outputs(5293)) xor (layer2_outputs(6524));
    outputs(12662) <= layer2_outputs(9036);
    outputs(12663) <= (layer2_outputs(8470)) or (layer2_outputs(8188));
    outputs(12664) <= not((layer2_outputs(5959)) xor (layer2_outputs(6100)));
    outputs(12665) <= not(layer2_outputs(10757));
    outputs(12666) <= layer2_outputs(6645);
    outputs(12667) <= (layer2_outputs(658)) xor (layer2_outputs(2728));
    outputs(12668) <= layer2_outputs(2985);
    outputs(12669) <= (layer2_outputs(6998)) and (layer2_outputs(11959));
    outputs(12670) <= not(layer2_outputs(28));
    outputs(12671) <= layer2_outputs(9157);
    outputs(12672) <= not(layer2_outputs(3501));
    outputs(12673) <= layer2_outputs(341);
    outputs(12674) <= not(layer2_outputs(12620));
    outputs(12675) <= (layer2_outputs(2417)) or (layer2_outputs(488));
    outputs(12676) <= not((layer2_outputs(11145)) xor (layer2_outputs(1148)));
    outputs(12677) <= (layer2_outputs(5547)) and (layer2_outputs(11853));
    outputs(12678) <= (layer2_outputs(6178)) and not (layer2_outputs(10600));
    outputs(12679) <= (layer2_outputs(11827)) or (layer2_outputs(7941));
    outputs(12680) <= (layer2_outputs(5211)) and not (layer2_outputs(5237));
    outputs(12681) <= (layer2_outputs(10633)) xor (layer2_outputs(10982));
    outputs(12682) <= not(layer2_outputs(5210));
    outputs(12683) <= layer2_outputs(8070);
    outputs(12684) <= layer2_outputs(11036);
    outputs(12685) <= layer2_outputs(1170);
    outputs(12686) <= (layer2_outputs(6119)) and not (layer2_outputs(11720));
    outputs(12687) <= not(layer2_outputs(7254));
    outputs(12688) <= (layer2_outputs(1174)) xor (layer2_outputs(10093));
    outputs(12689) <= not((layer2_outputs(5640)) xor (layer2_outputs(12478)));
    outputs(12690) <= not(layer2_outputs(253));
    outputs(12691) <= not(layer2_outputs(4946));
    outputs(12692) <= layer2_outputs(1898);
    outputs(12693) <= not((layer2_outputs(3687)) xor (layer2_outputs(409)));
    outputs(12694) <= not(layer2_outputs(11061));
    outputs(12695) <= not((layer2_outputs(1582)) xor (layer2_outputs(9162)));
    outputs(12696) <= (layer2_outputs(5375)) or (layer2_outputs(6917));
    outputs(12697) <= not(layer2_outputs(9494)) or (layer2_outputs(268));
    outputs(12698) <= (layer2_outputs(3607)) and not (layer2_outputs(8374));
    outputs(12699) <= (layer2_outputs(5318)) xor (layer2_outputs(1589));
    outputs(12700) <= not((layer2_outputs(152)) xor (layer2_outputs(6348)));
    outputs(12701) <= not((layer2_outputs(372)) xor (layer2_outputs(7986)));
    outputs(12702) <= (layer2_outputs(7782)) and (layer2_outputs(2751));
    outputs(12703) <= not((layer2_outputs(722)) xor (layer2_outputs(6800)));
    outputs(12704) <= not(layer2_outputs(10945));
    outputs(12705) <= not((layer2_outputs(1074)) xor (layer2_outputs(8305)));
    outputs(12706) <= layer2_outputs(11271);
    outputs(12707) <= layer2_outputs(8885);
    outputs(12708) <= layer2_outputs(8293);
    outputs(12709) <= (layer2_outputs(1552)) and (layer2_outputs(4520));
    outputs(12710) <= not((layer2_outputs(1928)) xor (layer2_outputs(2084)));
    outputs(12711) <= layer2_outputs(1437);
    outputs(12712) <= layer2_outputs(11051);
    outputs(12713) <= not(layer2_outputs(5186));
    outputs(12714) <= not((layer2_outputs(9630)) xor (layer2_outputs(3188)));
    outputs(12715) <= not(layer2_outputs(3064));
    outputs(12716) <= not((layer2_outputs(11855)) xor (layer2_outputs(9804)));
    outputs(12717) <= (layer2_outputs(1271)) and (layer2_outputs(5680));
    outputs(12718) <= layer2_outputs(5942);
    outputs(12719) <= layer2_outputs(1177);
    outputs(12720) <= layer2_outputs(10366);
    outputs(12721) <= (layer2_outputs(9002)) xor (layer2_outputs(2807));
    outputs(12722) <= (layer2_outputs(10979)) xor (layer2_outputs(11248));
    outputs(12723) <= not(layer2_outputs(7104));
    outputs(12724) <= not((layer2_outputs(7339)) xor (layer2_outputs(6378)));
    outputs(12725) <= (layer2_outputs(11940)) and not (layer2_outputs(2429));
    outputs(12726) <= layer2_outputs(8564);
    outputs(12727) <= layer2_outputs(11936);
    outputs(12728) <= (layer2_outputs(9821)) xor (layer2_outputs(9683));
    outputs(12729) <= not(layer2_outputs(4003));
    outputs(12730) <= (layer2_outputs(11309)) xor (layer2_outputs(5604));
    outputs(12731) <= (layer2_outputs(1591)) or (layer2_outputs(10159));
    outputs(12732) <= layer2_outputs(5434);
    outputs(12733) <= not(layer2_outputs(526));
    outputs(12734) <= not(layer2_outputs(9026)) or (layer2_outputs(1970));
    outputs(12735) <= not(layer2_outputs(8506));
    outputs(12736) <= (layer2_outputs(12418)) or (layer2_outputs(9821));
    outputs(12737) <= (layer2_outputs(2107)) or (layer2_outputs(8376));
    outputs(12738) <= (layer2_outputs(4182)) and (layer2_outputs(1408));
    outputs(12739) <= not((layer2_outputs(864)) xor (layer2_outputs(8747)));
    outputs(12740) <= layer2_outputs(4688);
    outputs(12741) <= not((layer2_outputs(2465)) xor (layer2_outputs(3272)));
    outputs(12742) <= (layer2_outputs(3202)) xor (layer2_outputs(3015));
    outputs(12743) <= layer2_outputs(5047);
    outputs(12744) <= not(layer2_outputs(10381));
    outputs(12745) <= (layer2_outputs(11232)) xor (layer2_outputs(11253));
    outputs(12746) <= layer2_outputs(10350);
    outputs(12747) <= not(layer2_outputs(4454));
    outputs(12748) <= layer2_outputs(10177);
    outputs(12749) <= layer2_outputs(10486);
    outputs(12750) <= layer2_outputs(11748);
    outputs(12751) <= layer2_outputs(529);
    outputs(12752) <= not(layer2_outputs(6508)) or (layer2_outputs(1832));
    outputs(12753) <= not(layer2_outputs(3585));
    outputs(12754) <= layer2_outputs(6755);
    outputs(12755) <= (layer2_outputs(106)) xor (layer2_outputs(7280));
    outputs(12756) <= layer2_outputs(8998);
    outputs(12757) <= not(layer2_outputs(6009));
    outputs(12758) <= not(layer2_outputs(8675));
    outputs(12759) <= not((layer2_outputs(12556)) and (layer2_outputs(6665)));
    outputs(12760) <= not((layer2_outputs(10189)) xor (layer2_outputs(6253)));
    outputs(12761) <= not(layer2_outputs(1505));
    outputs(12762) <= (layer2_outputs(11700)) and not (layer2_outputs(7826));
    outputs(12763) <= layer2_outputs(1295);
    outputs(12764) <= not(layer2_outputs(10036));
    outputs(12765) <= not((layer2_outputs(7543)) xor (layer2_outputs(3012)));
    outputs(12766) <= not(layer2_outputs(10601)) or (layer2_outputs(7718));
    outputs(12767) <= not(layer2_outputs(8848));
    outputs(12768) <= not(layer2_outputs(6401));
    outputs(12769) <= layer2_outputs(8570);
    outputs(12770) <= not(layer2_outputs(7111));
    outputs(12771) <= not(layer2_outputs(78));
    outputs(12772) <= not(layer2_outputs(7161));
    outputs(12773) <= not(layer2_outputs(1136)) or (layer2_outputs(2395));
    outputs(12774) <= layer2_outputs(9053);
    outputs(12775) <= not(layer2_outputs(765));
    outputs(12776) <= not((layer2_outputs(3462)) xor (layer2_outputs(6319)));
    outputs(12777) <= not((layer2_outputs(1031)) xor (layer2_outputs(5863)));
    outputs(12778) <= (layer2_outputs(11173)) and not (layer2_outputs(9325));
    outputs(12779) <= layer2_outputs(2847);
    outputs(12780) <= not(layer2_outputs(2918));
    outputs(12781) <= not((layer2_outputs(6666)) and (layer2_outputs(8356)));
    outputs(12782) <= (layer2_outputs(5951)) xor (layer2_outputs(3941));
    outputs(12783) <= not(layer2_outputs(11811));
    outputs(12784) <= layer2_outputs(8869);
    outputs(12785) <= not(layer2_outputs(8124));
    outputs(12786) <= (layer2_outputs(12380)) xor (layer2_outputs(10074));
    outputs(12787) <= not(layer2_outputs(8102));
    outputs(12788) <= (layer2_outputs(360)) and not (layer2_outputs(90));
    outputs(12789) <= (layer2_outputs(4435)) xor (layer2_outputs(11019));
    outputs(12790) <= layer2_outputs(2598);
    outputs(12791) <= (layer2_outputs(5860)) and (layer2_outputs(6752));
    outputs(12792) <= not((layer2_outputs(9664)) xor (layer2_outputs(45)));
    outputs(12793) <= layer2_outputs(3027);
    outputs(12794) <= not(layer2_outputs(3452));
    outputs(12795) <= layer2_outputs(10427);
    outputs(12796) <= not(layer2_outputs(11737));
    outputs(12797) <= (layer2_outputs(12561)) and not (layer2_outputs(4439));
    outputs(12798) <= layer2_outputs(6690);
    outputs(12799) <= (layer2_outputs(3714)) xor (layer2_outputs(7591));

end Behavioral;
