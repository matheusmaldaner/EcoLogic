library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs: in std_logic_vector(1023 downto 0);
        outputs: out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs: std_logic_vector(7679 downto 0);

begin
    layer0_outputs(0) <= b;
    layer0_outputs(1) <= not b;
    layer0_outputs(2) <= not a;
    layer0_outputs(3) <= not (a or b);
    layer0_outputs(4) <= not (a or b);
    layer0_outputs(5) <= a xor b;
    layer0_outputs(6) <= a xor b;
    layer0_outputs(7) <= not (a or b);
    layer0_outputs(8) <= not b;
    layer0_outputs(9) <= a or b;
    layer0_outputs(10) <= a or b;
    layer0_outputs(11) <= not b;
    layer0_outputs(12) <= a xor b;
    layer0_outputs(13) <= b;
    layer0_outputs(14) <= 1'b1;
    layer0_outputs(15) <= not (a xor b);
    layer0_outputs(16) <= not (a or b);
    layer0_outputs(17) <= a or b;
    layer0_outputs(18) <= a or b;
    layer0_outputs(19) <= not a;
    layer0_outputs(20) <= not b or a;
    layer0_outputs(21) <= not b or a;
    layer0_outputs(22) <= b;
    layer0_outputs(23) <= not b;
    layer0_outputs(24) <= a xor b;
    layer0_outputs(25) <= a or b;
    layer0_outputs(26) <= not (a or b);
    layer0_outputs(27) <= not b or a;
    layer0_outputs(28) <= not (a or b);
    layer0_outputs(29) <= not b;
    layer0_outputs(30) <= not (a or b);
    layer0_outputs(31) <= b;
    layer0_outputs(32) <= b;
    layer0_outputs(33) <= not a or b;
    layer0_outputs(34) <= not (a or b);
    layer0_outputs(35) <= not (a or b);
    layer0_outputs(36) <= not (a or b);
    layer0_outputs(37) <= not (a or b);
    layer0_outputs(38) <= not (a or b);
    layer0_outputs(39) <= a xor b;
    layer0_outputs(40) <= not (a or b);
    layer0_outputs(41) <= a and not b;
    layer0_outputs(42) <= a xor b;
    layer0_outputs(43) <= b;
    layer0_outputs(44) <= not (a xor b);
    layer0_outputs(45) <= not (a xor b);
    layer0_outputs(46) <= not (a and b);
    layer0_outputs(47) <= not a or b;
    layer0_outputs(48) <= not (a or b);
    layer0_outputs(49) <= b and not a;
    layer0_outputs(50) <= not (a xor b);
    layer0_outputs(51) <= not a;
    layer0_outputs(52) <= not a;
    layer0_outputs(53) <= not a;
    layer0_outputs(54) <= b and not a;
    layer0_outputs(55) <= a and not b;
    layer0_outputs(56) <= not (a or b);
    layer0_outputs(57) <= a xor b;
    layer0_outputs(58) <= b and not a;
    layer0_outputs(59) <= a xor b;
    layer0_outputs(60) <= not a or b;
    layer0_outputs(61) <= a xor b;
    layer0_outputs(62) <= b and not a;
    layer0_outputs(63) <= not b or a;
    layer0_outputs(64) <= a and b;
    layer0_outputs(65) <= not b or a;
    layer0_outputs(66) <= a;
    layer0_outputs(67) <= not (a xor b);
    layer0_outputs(68) <= b and not a;
    layer0_outputs(69) <= not b or a;
    layer0_outputs(70) <= a;
    layer0_outputs(71) <= a;
    layer0_outputs(72) <= not a or b;
    layer0_outputs(73) <= a and not b;
    layer0_outputs(74) <= a and not b;
    layer0_outputs(75) <= not b or a;
    layer0_outputs(76) <= a or b;
    layer0_outputs(77) <= a;
    layer0_outputs(78) <= not (a and b);
    layer0_outputs(79) <= b and not a;
    layer0_outputs(80) <= a and not b;
    layer0_outputs(81) <= b;
    layer0_outputs(82) <= a or b;
    layer0_outputs(83) <= not b or a;
    layer0_outputs(84) <= not (a xor b);
    layer0_outputs(85) <= not b or a;
    layer0_outputs(86) <= a or b;
    layer0_outputs(87) <= not a;
    layer0_outputs(88) <= not (a xor b);
    layer0_outputs(89) <= a xor b;
    layer0_outputs(90) <= a or b;
    layer0_outputs(91) <= a or b;
    layer0_outputs(92) <= not b or a;
    layer0_outputs(93) <= not (a or b);
    layer0_outputs(94) <= a or b;
    layer0_outputs(95) <= a xor b;
    layer0_outputs(96) <= 1'b0;
    layer0_outputs(97) <= not b;
    layer0_outputs(98) <= b and not a;
    layer0_outputs(99) <= a and not b;
    layer0_outputs(100) <= not b;
    layer0_outputs(101) <= b;
    layer0_outputs(102) <= a;
    layer0_outputs(103) <= not a;
    layer0_outputs(104) <= a or b;
    layer0_outputs(105) <= a xor b;
    layer0_outputs(106) <= not (a or b);
    layer0_outputs(107) <= b and not a;
    layer0_outputs(108) <= b;
    layer0_outputs(109) <= a or b;
    layer0_outputs(110) <= a or b;
    layer0_outputs(111) <= a and not b;
    layer0_outputs(112) <= b and not a;
    layer0_outputs(113) <= not (a and b);
    layer0_outputs(114) <= a or b;
    layer0_outputs(115) <= not a or b;
    layer0_outputs(116) <= not a;
    layer0_outputs(117) <= a xor b;
    layer0_outputs(118) <= not (a or b);
    layer0_outputs(119) <= a;
    layer0_outputs(120) <= a xor b;
    layer0_outputs(121) <= a or b;
    layer0_outputs(122) <= not (a or b);
    layer0_outputs(123) <= not (a or b);
    layer0_outputs(124) <= a;
    layer0_outputs(125) <= 1'b0;
    layer0_outputs(126) <= b;
    layer0_outputs(127) <= a xor b;
    layer0_outputs(128) <= not (a xor b);
    layer0_outputs(129) <= a or b;
    layer0_outputs(130) <= not (a or b);
    layer0_outputs(131) <= not b or a;
    layer0_outputs(132) <= a and not b;
    layer0_outputs(133) <= not a;
    layer0_outputs(134) <= a or b;
    layer0_outputs(135) <= a;
    layer0_outputs(136) <= a or b;
    layer0_outputs(137) <= a or b;
    layer0_outputs(138) <= not (a or b);
    layer0_outputs(139) <= a;
    layer0_outputs(140) <= not (a or b);
    layer0_outputs(141) <= not b;
    layer0_outputs(142) <= not a;
    layer0_outputs(143) <= not a;
    layer0_outputs(144) <= a or b;
    layer0_outputs(145) <= a and not b;
    layer0_outputs(146) <= a;
    layer0_outputs(147) <= a and not b;
    layer0_outputs(148) <= b and not a;
    layer0_outputs(149) <= a;
    layer0_outputs(150) <= a xor b;
    layer0_outputs(151) <= not (a or b);
    layer0_outputs(152) <= not a;
    layer0_outputs(153) <= not (a xor b);
    layer0_outputs(154) <= not (a or b);
    layer0_outputs(155) <= not (a or b);
    layer0_outputs(156) <= a;
    layer0_outputs(157) <= 1'b0;
    layer0_outputs(158) <= not b or a;
    layer0_outputs(159) <= a or b;
    layer0_outputs(160) <= not (a xor b);
    layer0_outputs(161) <= not b or a;
    layer0_outputs(162) <= not b or a;
    layer0_outputs(163) <= a or b;
    layer0_outputs(164) <= b and not a;
    layer0_outputs(165) <= a xor b;
    layer0_outputs(166) <= not b or a;
    layer0_outputs(167) <= not a or b;
    layer0_outputs(168) <= not (a and b);
    layer0_outputs(169) <= b;
    layer0_outputs(170) <= a xor b;
    layer0_outputs(171) <= not a or b;
    layer0_outputs(172) <= not a;
    layer0_outputs(173) <= not (a or b);
    layer0_outputs(174) <= a xor b;
    layer0_outputs(175) <= a and b;
    layer0_outputs(176) <= b and not a;
    layer0_outputs(177) <= not (a and b);
    layer0_outputs(178) <= a;
    layer0_outputs(179) <= not (a xor b);
    layer0_outputs(180) <= a or b;
    layer0_outputs(181) <= b;
    layer0_outputs(182) <= not a;
    layer0_outputs(183) <= a and not b;
    layer0_outputs(184) <= not (a xor b);
    layer0_outputs(185) <= a or b;
    layer0_outputs(186) <= not (a xor b);
    layer0_outputs(187) <= not (a or b);
    layer0_outputs(188) <= a or b;
    layer0_outputs(189) <= not b;
    layer0_outputs(190) <= not (a or b);
    layer0_outputs(191) <= a and b;
    layer0_outputs(192) <= not a or b;
    layer0_outputs(193) <= not (a and b);
    layer0_outputs(194) <= not (a xor b);
    layer0_outputs(195) <= a xor b;
    layer0_outputs(196) <= not a or b;
    layer0_outputs(197) <= a or b;
    layer0_outputs(198) <= a or b;
    layer0_outputs(199) <= not b or a;
    layer0_outputs(200) <= a or b;
    layer0_outputs(201) <= not b;
    layer0_outputs(202) <= a;
    layer0_outputs(203) <= a and not b;
    layer0_outputs(204) <= b;
    layer0_outputs(205) <= 1'b0;
    layer0_outputs(206) <= not b;
    layer0_outputs(207) <= b and not a;
    layer0_outputs(208) <= a or b;
    layer0_outputs(209) <= a;
    layer0_outputs(210) <= not (a and b);
    layer0_outputs(211) <= a and not b;
    layer0_outputs(212) <= a;
    layer0_outputs(213) <= a or b;
    layer0_outputs(214) <= not a;
    layer0_outputs(215) <= not b or a;
    layer0_outputs(216) <= not b or a;
    layer0_outputs(217) <= not a or b;
    layer0_outputs(218) <= b and not a;
    layer0_outputs(219) <= not a;
    layer0_outputs(220) <= b;
    layer0_outputs(221) <= a and not b;
    layer0_outputs(222) <= not (a xor b);
    layer0_outputs(223) <= a xor b;
    layer0_outputs(224) <= a or b;
    layer0_outputs(225) <= b and not a;
    layer0_outputs(226) <= a and not b;
    layer0_outputs(227) <= not a or b;
    layer0_outputs(228) <= b and not a;
    layer0_outputs(229) <= not b;
    layer0_outputs(230) <= b and not a;
    layer0_outputs(231) <= not (a or b);
    layer0_outputs(232) <= a;
    layer0_outputs(233) <= a;
    layer0_outputs(234) <= not b;
    layer0_outputs(235) <= a and not b;
    layer0_outputs(236) <= b and not a;
    layer0_outputs(237) <= a or b;
    layer0_outputs(238) <= not a or b;
    layer0_outputs(239) <= not b;
    layer0_outputs(240) <= not (a or b);
    layer0_outputs(241) <= not b;
    layer0_outputs(242) <= not (a xor b);
    layer0_outputs(243) <= a or b;
    layer0_outputs(244) <= not (a or b);
    layer0_outputs(245) <= not b;
    layer0_outputs(246) <= b;
    layer0_outputs(247) <= 1'b1;
    layer0_outputs(248) <= not b;
    layer0_outputs(249) <= not b or a;
    layer0_outputs(250) <= a xor b;
    layer0_outputs(251) <= a or b;
    layer0_outputs(252) <= not (a xor b);
    layer0_outputs(253) <= not (a or b);
    layer0_outputs(254) <= not a;
    layer0_outputs(255) <= not (a or b);
    layer0_outputs(256) <= a or b;
    layer0_outputs(257) <= not a or b;
    layer0_outputs(258) <= 1'b0;
    layer0_outputs(259) <= a and not b;
    layer0_outputs(260) <= a and not b;
    layer0_outputs(261) <= a and not b;
    layer0_outputs(262) <= not (a or b);
    layer0_outputs(263) <= not (a or b);
    layer0_outputs(264) <= not b or a;
    layer0_outputs(265) <= not (a xor b);
    layer0_outputs(266) <= a or b;
    layer0_outputs(267) <= a and b;
    layer0_outputs(268) <= not (a xor b);
    layer0_outputs(269) <= a or b;
    layer0_outputs(270) <= b and not a;
    layer0_outputs(271) <= a and not b;
    layer0_outputs(272) <= not (a or b);
    layer0_outputs(273) <= a or b;
    layer0_outputs(274) <= not (a xor b);
    layer0_outputs(275) <= a or b;
    layer0_outputs(276) <= a or b;
    layer0_outputs(277) <= b;
    layer0_outputs(278) <= not b;
    layer0_outputs(279) <= not (a and b);
    layer0_outputs(280) <= a or b;
    layer0_outputs(281) <= not (a or b);
    layer0_outputs(282) <= not (a xor b);
    layer0_outputs(283) <= a xor b;
    layer0_outputs(284) <= not a;
    layer0_outputs(285) <= a;
    layer0_outputs(286) <= b and not a;
    layer0_outputs(287) <= a xor b;
    layer0_outputs(288) <= a or b;
    layer0_outputs(289) <= b and not a;
    layer0_outputs(290) <= b;
    layer0_outputs(291) <= not a;
    layer0_outputs(292) <= a;
    layer0_outputs(293) <= a xor b;
    layer0_outputs(294) <= not (a xor b);
    layer0_outputs(295) <= not b or a;
    layer0_outputs(296) <= not (a or b);
    layer0_outputs(297) <= not b or a;
    layer0_outputs(298) <= 1'b1;
    layer0_outputs(299) <= not (a or b);
    layer0_outputs(300) <= not a;
    layer0_outputs(301) <= not b or a;
    layer0_outputs(302) <= a and not b;
    layer0_outputs(303) <= b and not a;
    layer0_outputs(304) <= a and not b;
    layer0_outputs(305) <= 1'b0;
    layer0_outputs(306) <= not (a or b);
    layer0_outputs(307) <= a or b;
    layer0_outputs(308) <= not a or b;
    layer0_outputs(309) <= b and not a;
    layer0_outputs(310) <= not (a xor b);
    layer0_outputs(311) <= not (a xor b);
    layer0_outputs(312) <= a;
    layer0_outputs(313) <= not a or b;
    layer0_outputs(314) <= not b;
    layer0_outputs(315) <= not (a xor b);
    layer0_outputs(316) <= not (a xor b);
    layer0_outputs(317) <= not (a or b);
    layer0_outputs(318) <= not (a or b);
    layer0_outputs(319) <= not a or b;
    layer0_outputs(320) <= a xor b;
    layer0_outputs(321) <= not (a xor b);
    layer0_outputs(322) <= not a;
    layer0_outputs(323) <= not b or a;
    layer0_outputs(324) <= b and not a;
    layer0_outputs(325) <= a xor b;
    layer0_outputs(326) <= a xor b;
    layer0_outputs(327) <= a xor b;
    layer0_outputs(328) <= a xor b;
    layer0_outputs(329) <= a and not b;
    layer0_outputs(330) <= b and not a;
    layer0_outputs(331) <= not (a or b);
    layer0_outputs(332) <= not (a or b);
    layer0_outputs(333) <= a and not b;
    layer0_outputs(334) <= a xor b;
    layer0_outputs(335) <= b;
    layer0_outputs(336) <= b;
    layer0_outputs(337) <= not b or a;
    layer0_outputs(338) <= a or b;
    layer0_outputs(339) <= b and not a;
    layer0_outputs(340) <= a and b;
    layer0_outputs(341) <= not a or b;
    layer0_outputs(342) <= not (a or b);
    layer0_outputs(343) <= not b;
    layer0_outputs(344) <= a xor b;
    layer0_outputs(345) <= a;
    layer0_outputs(346) <= not a;
    layer0_outputs(347) <= a xor b;
    layer0_outputs(348) <= 1'b1;
    layer0_outputs(349) <= not (a xor b);
    layer0_outputs(350) <= not (a or b);
    layer0_outputs(351) <= not b;
    layer0_outputs(352) <= not (a or b);
    layer0_outputs(353) <= a xor b;
    layer0_outputs(354) <= 1'b0;
    layer0_outputs(355) <= not (a and b);
    layer0_outputs(356) <= not b or a;
    layer0_outputs(357) <= not (a xor b);
    layer0_outputs(358) <= b;
    layer0_outputs(359) <= a;
    layer0_outputs(360) <= a;
    layer0_outputs(361) <= not b;
    layer0_outputs(362) <= not b;
    layer0_outputs(363) <= a xor b;
    layer0_outputs(364) <= not b;
    layer0_outputs(365) <= a xor b;
    layer0_outputs(366) <= a;
    layer0_outputs(367) <= not (a xor b);
    layer0_outputs(368) <= b and not a;
    layer0_outputs(369) <= b and not a;
    layer0_outputs(370) <= not (a xor b);
    layer0_outputs(371) <= a;
    layer0_outputs(372) <= a or b;
    layer0_outputs(373) <= not a;
    layer0_outputs(374) <= a;
    layer0_outputs(375) <= a or b;
    layer0_outputs(376) <= b and not a;
    layer0_outputs(377) <= not (a xor b);
    layer0_outputs(378) <= not b;
    layer0_outputs(379) <= not (a xor b);
    layer0_outputs(380) <= a;
    layer0_outputs(381) <= a;
    layer0_outputs(382) <= not b or a;
    layer0_outputs(383) <= not (a xor b);
    layer0_outputs(384) <= a;
    layer0_outputs(385) <= a and b;
    layer0_outputs(386) <= b;
    layer0_outputs(387) <= not b;
    layer0_outputs(388) <= a or b;
    layer0_outputs(389) <= not a;
    layer0_outputs(390) <= not b;
    layer0_outputs(391) <= a;
    layer0_outputs(392) <= a xor b;
    layer0_outputs(393) <= not b or a;
    layer0_outputs(394) <= not b;
    layer0_outputs(395) <= a and not b;
    layer0_outputs(396) <= not a or b;
    layer0_outputs(397) <= not (a or b);
    layer0_outputs(398) <= b;
    layer0_outputs(399) <= not a;
    layer0_outputs(400) <= a xor b;
    layer0_outputs(401) <= not (a xor b);
    layer0_outputs(402) <= a and b;
    layer0_outputs(403) <= not b;
    layer0_outputs(404) <= not b;
    layer0_outputs(405) <= b;
    layer0_outputs(406) <= not (a xor b);
    layer0_outputs(407) <= not b;
    layer0_outputs(408) <= not b;
    layer0_outputs(409) <= not b or a;
    layer0_outputs(410) <= not b or a;
    layer0_outputs(411) <= not a;
    layer0_outputs(412) <= b and not a;
    layer0_outputs(413) <= not a or b;
    layer0_outputs(414) <= a and b;
    layer0_outputs(415) <= a or b;
    layer0_outputs(416) <= not a;
    layer0_outputs(417) <= not (a or b);
    layer0_outputs(418) <= a or b;
    layer0_outputs(419) <= not (a or b);
    layer0_outputs(420) <= a and not b;
    layer0_outputs(421) <= not b;
    layer0_outputs(422) <= a;
    layer0_outputs(423) <= b and not a;
    layer0_outputs(424) <= a and b;
    layer0_outputs(425) <= b and not a;
    layer0_outputs(426) <= b;
    layer0_outputs(427) <= not (a xor b);
    layer0_outputs(428) <= not b;
    layer0_outputs(429) <= a or b;
    layer0_outputs(430) <= not b or a;
    layer0_outputs(431) <= b;
    layer0_outputs(432) <= a or b;
    layer0_outputs(433) <= not (a xor b);
    layer0_outputs(434) <= not (a or b);
    layer0_outputs(435) <= a or b;
    layer0_outputs(436) <= b and not a;
    layer0_outputs(437) <= not a or b;
    layer0_outputs(438) <= not (a or b);
    layer0_outputs(439) <= a and not b;
    layer0_outputs(440) <= a or b;
    layer0_outputs(441) <= a and not b;
    layer0_outputs(442) <= not b;
    layer0_outputs(443) <= a;
    layer0_outputs(444) <= b and not a;
    layer0_outputs(445) <= a xor b;
    layer0_outputs(446) <= a;
    layer0_outputs(447) <= a and not b;
    layer0_outputs(448) <= not a;
    layer0_outputs(449) <= not a or b;
    layer0_outputs(450) <= not a or b;
    layer0_outputs(451) <= not a;
    layer0_outputs(452) <= a or b;
    layer0_outputs(453) <= a xor b;
    layer0_outputs(454) <= not (a or b);
    layer0_outputs(455) <= a xor b;
    layer0_outputs(456) <= not b or a;
    layer0_outputs(457) <= not (a or b);
    layer0_outputs(458) <= not (a or b);
    layer0_outputs(459) <= a xor b;
    layer0_outputs(460) <= b and not a;
    layer0_outputs(461) <= not a or b;
    layer0_outputs(462) <= b;
    layer0_outputs(463) <= a and b;
    layer0_outputs(464) <= not b;
    layer0_outputs(465) <= a xor b;
    layer0_outputs(466) <= not (a or b);
    layer0_outputs(467) <= a and b;
    layer0_outputs(468) <= a or b;
    layer0_outputs(469) <= not b;
    layer0_outputs(470) <= 1'b1;
    layer0_outputs(471) <= 1'b0;
    layer0_outputs(472) <= not b or a;
    layer0_outputs(473) <= not (a or b);
    layer0_outputs(474) <= a;
    layer0_outputs(475) <= 1'b0;
    layer0_outputs(476) <= a and not b;
    layer0_outputs(477) <= a or b;
    layer0_outputs(478) <= b and not a;
    layer0_outputs(479) <= a and not b;
    layer0_outputs(480) <= not (a or b);
    layer0_outputs(481) <= not a;
    layer0_outputs(482) <= a and b;
    layer0_outputs(483) <= a or b;
    layer0_outputs(484) <= 1'b0;
    layer0_outputs(485) <= not (a xor b);
    layer0_outputs(486) <= a or b;
    layer0_outputs(487) <= not b or a;
    layer0_outputs(488) <= a or b;
    layer0_outputs(489) <= a or b;
    layer0_outputs(490) <= not (a or b);
    layer0_outputs(491) <= a and not b;
    layer0_outputs(492) <= not b or a;
    layer0_outputs(493) <= not a or b;
    layer0_outputs(494) <= not (a or b);
    layer0_outputs(495) <= b;
    layer0_outputs(496) <= not b or a;
    layer0_outputs(497) <= not (a or b);
    layer0_outputs(498) <= not b;
    layer0_outputs(499) <= not (a xor b);
    layer0_outputs(500) <= not a;
    layer0_outputs(501) <= b and not a;
    layer0_outputs(502) <= not (a xor b);
    layer0_outputs(503) <= not a or b;
    layer0_outputs(504) <= not (a xor b);
    layer0_outputs(505) <= not (a and b);
    layer0_outputs(506) <= not (a or b);
    layer0_outputs(507) <= a or b;
    layer0_outputs(508) <= a;
    layer0_outputs(509) <= b;
    layer0_outputs(510) <= not b;
    layer0_outputs(511) <= not (a xor b);
    layer0_outputs(512) <= not (a xor b);
    layer0_outputs(513) <= 1'b1;
    layer0_outputs(514) <= not a or b;
    layer0_outputs(515) <= not (a or b);
    layer0_outputs(516) <= a;
    layer0_outputs(517) <= a or b;
    layer0_outputs(518) <= a and not b;
    layer0_outputs(519) <= not a;
    layer0_outputs(520) <= not (a xor b);
    layer0_outputs(521) <= a or b;
    layer0_outputs(522) <= not (a xor b);
    layer0_outputs(523) <= a and b;
    layer0_outputs(524) <= not b;
    layer0_outputs(525) <= a xor b;
    layer0_outputs(526) <= not b;
    layer0_outputs(527) <= not (a and b);
    layer0_outputs(528) <= a;
    layer0_outputs(529) <= not (a or b);
    layer0_outputs(530) <= a and not b;
    layer0_outputs(531) <= not (a xor b);
    layer0_outputs(532) <= a;
    layer0_outputs(533) <= not b or a;
    layer0_outputs(534) <= b and not a;
    layer0_outputs(535) <= not a or b;
    layer0_outputs(536) <= b;
    layer0_outputs(537) <= b;
    layer0_outputs(538) <= not b or a;
    layer0_outputs(539) <= 1'b1;
    layer0_outputs(540) <= a and b;
    layer0_outputs(541) <= not (a xor b);
    layer0_outputs(542) <= a or b;
    layer0_outputs(543) <= a xor b;
    layer0_outputs(544) <= not b or a;
    layer0_outputs(545) <= a;
    layer0_outputs(546) <= not (a or b);
    layer0_outputs(547) <= not (a xor b);
    layer0_outputs(548) <= a and not b;
    layer0_outputs(549) <= a and not b;
    layer0_outputs(550) <= b;
    layer0_outputs(551) <= a and b;
    layer0_outputs(552) <= not a or b;
    layer0_outputs(553) <= a or b;
    layer0_outputs(554) <= a or b;
    layer0_outputs(555) <= a xor b;
    layer0_outputs(556) <= not a;
    layer0_outputs(557) <= a;
    layer0_outputs(558) <= b;
    layer0_outputs(559) <= not a;
    layer0_outputs(560) <= not (a and b);
    layer0_outputs(561) <= not (a or b);
    layer0_outputs(562) <= a xor b;
    layer0_outputs(563) <= a or b;
    layer0_outputs(564) <= not a or b;
    layer0_outputs(565) <= b;
    layer0_outputs(566) <= not a or b;
    layer0_outputs(567) <= not (a or b);
    layer0_outputs(568) <= a xor b;
    layer0_outputs(569) <= b and not a;
    layer0_outputs(570) <= not a or b;
    layer0_outputs(571) <= a;
    layer0_outputs(572) <= a or b;
    layer0_outputs(573) <= a or b;
    layer0_outputs(574) <= a or b;
    layer0_outputs(575) <= not b or a;
    layer0_outputs(576) <= not (a and b);
    layer0_outputs(577) <= not a;
    layer0_outputs(578) <= a xor b;
    layer0_outputs(579) <= a;
    layer0_outputs(580) <= a or b;
    layer0_outputs(581) <= a and not b;
    layer0_outputs(582) <= not a;
    layer0_outputs(583) <= a or b;
    layer0_outputs(584) <= not b;
    layer0_outputs(585) <= a;
    layer0_outputs(586) <= a and not b;
    layer0_outputs(587) <= b and not a;
    layer0_outputs(588) <= not (a xor b);
    layer0_outputs(589) <= not (a or b);
    layer0_outputs(590) <= not (a or b);
    layer0_outputs(591) <= 1'b1;
    layer0_outputs(592) <= a or b;
    layer0_outputs(593) <= not a;
    layer0_outputs(594) <= not a;
    layer0_outputs(595) <= not (a or b);
    layer0_outputs(596) <= a;
    layer0_outputs(597) <= not (a or b);
    layer0_outputs(598) <= not (a and b);
    layer0_outputs(599) <= a or b;
    layer0_outputs(600) <= not (a xor b);
    layer0_outputs(601) <= not (a or b);
    layer0_outputs(602) <= not (a xor b);
    layer0_outputs(603) <= a or b;
    layer0_outputs(604) <= a;
    layer0_outputs(605) <= b;
    layer0_outputs(606) <= a or b;
    layer0_outputs(607) <= b;
    layer0_outputs(608) <= b;
    layer0_outputs(609) <= not b or a;
    layer0_outputs(610) <= 1'b0;
    layer0_outputs(611) <= not (a or b);
    layer0_outputs(612) <= a or b;
    layer0_outputs(613) <= b;
    layer0_outputs(614) <= a or b;
    layer0_outputs(615) <= 1'b1;
    layer0_outputs(616) <= b;
    layer0_outputs(617) <= not b;
    layer0_outputs(618) <= not (a xor b);
    layer0_outputs(619) <= a xor b;
    layer0_outputs(620) <= not (a or b);
    layer0_outputs(621) <= not (a xor b);
    layer0_outputs(622) <= not b or a;
    layer0_outputs(623) <= not (a or b);
    layer0_outputs(624) <= b;
    layer0_outputs(625) <= not (a or b);
    layer0_outputs(626) <= a and not b;
    layer0_outputs(627) <= not b or a;
    layer0_outputs(628) <= not (a xor b);
    layer0_outputs(629) <= not (a xor b);
    layer0_outputs(630) <= a or b;
    layer0_outputs(631) <= a or b;
    layer0_outputs(632) <= a or b;
    layer0_outputs(633) <= not (a or b);
    layer0_outputs(634) <= a xor b;
    layer0_outputs(635) <= not b;
    layer0_outputs(636) <= a and not b;
    layer0_outputs(637) <= not (a or b);
    layer0_outputs(638) <= a or b;
    layer0_outputs(639) <= a and not b;
    layer0_outputs(640) <= a;
    layer0_outputs(641) <= not (a or b);
    layer0_outputs(642) <= not (a or b);
    layer0_outputs(643) <= a and not b;
    layer0_outputs(644) <= b and not a;
    layer0_outputs(645) <= a xor b;
    layer0_outputs(646) <= not b or a;
    layer0_outputs(647) <= not a;
    layer0_outputs(648) <= a;
    layer0_outputs(649) <= not (a or b);
    layer0_outputs(650) <= not (a or b);
    layer0_outputs(651) <= a and not b;
    layer0_outputs(652) <= 1'b1;
    layer0_outputs(653) <= a or b;
    layer0_outputs(654) <= not (a or b);
    layer0_outputs(655) <= a or b;
    layer0_outputs(656) <= b and not a;
    layer0_outputs(657) <= a;
    layer0_outputs(658) <= not a;
    layer0_outputs(659) <= a or b;
    layer0_outputs(660) <= a or b;
    layer0_outputs(661) <= not (a or b);
    layer0_outputs(662) <= not (a or b);
    layer0_outputs(663) <= a or b;
    layer0_outputs(664) <= a;
    layer0_outputs(665) <= not (a xor b);
    layer0_outputs(666) <= not a or b;
    layer0_outputs(667) <= a xor b;
    layer0_outputs(668) <= not a or b;
    layer0_outputs(669) <= not a or b;
    layer0_outputs(670) <= not a or b;
    layer0_outputs(671) <= a or b;
    layer0_outputs(672) <= a;
    layer0_outputs(673) <= a or b;
    layer0_outputs(674) <= a or b;
    layer0_outputs(675) <= not (a or b);
    layer0_outputs(676) <= a or b;
    layer0_outputs(677) <= a or b;
    layer0_outputs(678) <= a xor b;
    layer0_outputs(679) <= not a;
    layer0_outputs(680) <= not (a and b);
    layer0_outputs(681) <= a and not b;
    layer0_outputs(682) <= not a or b;
    layer0_outputs(683) <= a or b;
    layer0_outputs(684) <= not (a or b);
    layer0_outputs(685) <= not b or a;
    layer0_outputs(686) <= b and not a;
    layer0_outputs(687) <= not (a xor b);
    layer0_outputs(688) <= a and not b;
    layer0_outputs(689) <= a xor b;
    layer0_outputs(690) <= a;
    layer0_outputs(691) <= b and not a;
    layer0_outputs(692) <= a xor b;
    layer0_outputs(693) <= not a or b;
    layer0_outputs(694) <= not b;
    layer0_outputs(695) <= a and not b;
    layer0_outputs(696) <= a xor b;
    layer0_outputs(697) <= b and not a;
    layer0_outputs(698) <= a or b;
    layer0_outputs(699) <= a and not b;
    layer0_outputs(700) <= not (a xor b);
    layer0_outputs(701) <= not b or a;
    layer0_outputs(702) <= not b or a;
    layer0_outputs(703) <= b;
    layer0_outputs(704) <= not (a or b);
    layer0_outputs(705) <= a and not b;
    layer0_outputs(706) <= a and not b;
    layer0_outputs(707) <= not b;
    layer0_outputs(708) <= not a;
    layer0_outputs(709) <= not (a or b);
    layer0_outputs(710) <= a xor b;
    layer0_outputs(711) <= not (a or b);
    layer0_outputs(712) <= not a;
    layer0_outputs(713) <= not a or b;
    layer0_outputs(714) <= not (a and b);
    layer0_outputs(715) <= a and not b;
    layer0_outputs(716) <= a or b;
    layer0_outputs(717) <= not (a xor b);
    layer0_outputs(718) <= not (a or b);
    layer0_outputs(719) <= b;
    layer0_outputs(720) <= a;
    layer0_outputs(721) <= 1'b1;
    layer0_outputs(722) <= b;
    layer0_outputs(723) <= not b;
    layer0_outputs(724) <= not b or a;
    layer0_outputs(725) <= a or b;
    layer0_outputs(726) <= not a or b;
    layer0_outputs(727) <= a and not b;
    layer0_outputs(728) <= not a or b;
    layer0_outputs(729) <= not (a or b);
    layer0_outputs(730) <= not b or a;
    layer0_outputs(731) <= a xor b;
    layer0_outputs(732) <= a and not b;
    layer0_outputs(733) <= a or b;
    layer0_outputs(734) <= a or b;
    layer0_outputs(735) <= a or b;
    layer0_outputs(736) <= b;
    layer0_outputs(737) <= not (a xor b);
    layer0_outputs(738) <= a and not b;
    layer0_outputs(739) <= not (a or b);
    layer0_outputs(740) <= not (a xor b);
    layer0_outputs(741) <= a or b;
    layer0_outputs(742) <= not b or a;
    layer0_outputs(743) <= b;
    layer0_outputs(744) <= not b;
    layer0_outputs(745) <= a or b;
    layer0_outputs(746) <= not b or a;
    layer0_outputs(747) <= a;
    layer0_outputs(748) <= not b or a;
    layer0_outputs(749) <= not b;
    layer0_outputs(750) <= b and not a;
    layer0_outputs(751) <= not b or a;
    layer0_outputs(752) <= not b or a;
    layer0_outputs(753) <= a or b;
    layer0_outputs(754) <= not b;
    layer0_outputs(755) <= a and not b;
    layer0_outputs(756) <= a or b;
    layer0_outputs(757) <= not a or b;
    layer0_outputs(758) <= not (a xor b);
    layer0_outputs(759) <= 1'b1;
    layer0_outputs(760) <= not (a xor b);
    layer0_outputs(761) <= not a or b;
    layer0_outputs(762) <= a;
    layer0_outputs(763) <= a xor b;
    layer0_outputs(764) <= b and not a;
    layer0_outputs(765) <= a or b;
    layer0_outputs(766) <= a xor b;
    layer0_outputs(767) <= a xor b;
    layer0_outputs(768) <= a xor b;
    layer0_outputs(769) <= a and not b;
    layer0_outputs(770) <= not (a or b);
    layer0_outputs(771) <= a or b;
    layer0_outputs(772) <= not b;
    layer0_outputs(773) <= not a or b;
    layer0_outputs(774) <= b;
    layer0_outputs(775) <= a xor b;
    layer0_outputs(776) <= not (a xor b);
    layer0_outputs(777) <= not (a or b);
    layer0_outputs(778) <= not a;
    layer0_outputs(779) <= 1'b0;
    layer0_outputs(780) <= not b;
    layer0_outputs(781) <= a and not b;
    layer0_outputs(782) <= not b or a;
    layer0_outputs(783) <= not a or b;
    layer0_outputs(784) <= not (a xor b);
    layer0_outputs(785) <= a;
    layer0_outputs(786) <= not (a xor b);
    layer0_outputs(787) <= not (a or b);
    layer0_outputs(788) <= a xor b;
    layer0_outputs(789) <= b;
    layer0_outputs(790) <= 1'b0;
    layer0_outputs(791) <= a xor b;
    layer0_outputs(792) <= not (a or b);
    layer0_outputs(793) <= b;
    layer0_outputs(794) <= b;
    layer0_outputs(795) <= a xor b;
    layer0_outputs(796) <= not (a or b);
    layer0_outputs(797) <= not b or a;
    layer0_outputs(798) <= b;
    layer0_outputs(799) <= not (a or b);
    layer0_outputs(800) <= not a or b;
    layer0_outputs(801) <= b and not a;
    layer0_outputs(802) <= not b;
    layer0_outputs(803) <= a and not b;
    layer0_outputs(804) <= not (a or b);
    layer0_outputs(805) <= not (a or b);
    layer0_outputs(806) <= not (a or b);
    layer0_outputs(807) <= b;
    layer0_outputs(808) <= not a;
    layer0_outputs(809) <= not (a or b);
    layer0_outputs(810) <= a or b;
    layer0_outputs(811) <= not (a xor b);
    layer0_outputs(812) <= a and not b;
    layer0_outputs(813) <= a xor b;
    layer0_outputs(814) <= a and b;
    layer0_outputs(815) <= a and not b;
    layer0_outputs(816) <= not a or b;
    layer0_outputs(817) <= a or b;
    layer0_outputs(818) <= not (a or b);
    layer0_outputs(819) <= a xor b;
    layer0_outputs(820) <= not a;
    layer0_outputs(821) <= not b;
    layer0_outputs(822) <= not (a or b);
    layer0_outputs(823) <= not (a or b);
    layer0_outputs(824) <= not (a or b);
    layer0_outputs(825) <= not (a or b);
    layer0_outputs(826) <= not a or b;
    layer0_outputs(827) <= 1'b1;
    layer0_outputs(828) <= not (a or b);
    layer0_outputs(829) <= a xor b;
    layer0_outputs(830) <= not (a xor b);
    layer0_outputs(831) <= b;
    layer0_outputs(832) <= not (a or b);
    layer0_outputs(833) <= not b or a;
    layer0_outputs(834) <= not a;
    layer0_outputs(835) <= a or b;
    layer0_outputs(836) <= a xor b;
    layer0_outputs(837) <= a or b;
    layer0_outputs(838) <= a and not b;
    layer0_outputs(839) <= a xor b;
    layer0_outputs(840) <= a or b;
    layer0_outputs(841) <= 1'b1;
    layer0_outputs(842) <= a;
    layer0_outputs(843) <= not a or b;
    layer0_outputs(844) <= b;
    layer0_outputs(845) <= a xor b;
    layer0_outputs(846) <= a and not b;
    layer0_outputs(847) <= a;
    layer0_outputs(848) <= a or b;
    layer0_outputs(849) <= a xor b;
    layer0_outputs(850) <= not (a or b);
    layer0_outputs(851) <= not (a xor b);
    layer0_outputs(852) <= not b or a;
    layer0_outputs(853) <= a and not b;
    layer0_outputs(854) <= a;
    layer0_outputs(855) <= a;
    layer0_outputs(856) <= a or b;
    layer0_outputs(857) <= b;
    layer0_outputs(858) <= a and not b;
    layer0_outputs(859) <= a or b;
    layer0_outputs(860) <= not (a or b);
    layer0_outputs(861) <= not (a and b);
    layer0_outputs(862) <= a xor b;
    layer0_outputs(863) <= a and b;
    layer0_outputs(864) <= not b or a;
    layer0_outputs(865) <= b and not a;
    layer0_outputs(866) <= a;
    layer0_outputs(867) <= not (a xor b);
    layer0_outputs(868) <= a xor b;
    layer0_outputs(869) <= 1'b1;
    layer0_outputs(870) <= not (a xor b);
    layer0_outputs(871) <= a or b;
    layer0_outputs(872) <= b;
    layer0_outputs(873) <= a xor b;
    layer0_outputs(874) <= b and not a;
    layer0_outputs(875) <= a or b;
    layer0_outputs(876) <= not (a or b);
    layer0_outputs(877) <= not (a and b);
    layer0_outputs(878) <= 1'b1;
    layer0_outputs(879) <= a and b;
    layer0_outputs(880) <= not (a or b);
    layer0_outputs(881) <= a xor b;
    layer0_outputs(882) <= b and not a;
    layer0_outputs(883) <= b and not a;
    layer0_outputs(884) <= not (a or b);
    layer0_outputs(885) <= a or b;
    layer0_outputs(886) <= a;
    layer0_outputs(887) <= b;
    layer0_outputs(888) <= a xor b;
    layer0_outputs(889) <= a xor b;
    layer0_outputs(890) <= not b or a;
    layer0_outputs(891) <= b;
    layer0_outputs(892) <= not (a or b);
    layer0_outputs(893) <= a or b;
    layer0_outputs(894) <= not (a xor b);
    layer0_outputs(895) <= not (a or b);
    layer0_outputs(896) <= not a or b;
    layer0_outputs(897) <= not (a or b);
    layer0_outputs(898) <= a;
    layer0_outputs(899) <= a or b;
    layer0_outputs(900) <= a and not b;
    layer0_outputs(901) <= not b;
    layer0_outputs(902) <= b;
    layer0_outputs(903) <= not (a or b);
    layer0_outputs(904) <= not (a or b);
    layer0_outputs(905) <= not (a or b);
    layer0_outputs(906) <= not a or b;
    layer0_outputs(907) <= b;
    layer0_outputs(908) <= not a;
    layer0_outputs(909) <= not b;
    layer0_outputs(910) <= not a;
    layer0_outputs(911) <= 1'b0;
    layer0_outputs(912) <= not a or b;
    layer0_outputs(913) <= a or b;
    layer0_outputs(914) <= not a;
    layer0_outputs(915) <= not a or b;
    layer0_outputs(916) <= not b;
    layer0_outputs(917) <= a xor b;
    layer0_outputs(918) <= not b or a;
    layer0_outputs(919) <= not (a and b);
    layer0_outputs(920) <= not b or a;
    layer0_outputs(921) <= a or b;
    layer0_outputs(922) <= a or b;
    layer0_outputs(923) <= not a or b;
    layer0_outputs(924) <= a;
    layer0_outputs(925) <= not a or b;
    layer0_outputs(926) <= not (a or b);
    layer0_outputs(927) <= 1'b0;
    layer0_outputs(928) <= a;
    layer0_outputs(929) <= a or b;
    layer0_outputs(930) <= not (a or b);
    layer0_outputs(931) <= b and not a;
    layer0_outputs(932) <= not b or a;
    layer0_outputs(933) <= a and b;
    layer0_outputs(934) <= a and b;
    layer0_outputs(935) <= a and b;
    layer0_outputs(936) <= not b or a;
    layer0_outputs(937) <= not b;
    layer0_outputs(938) <= not (a xor b);
    layer0_outputs(939) <= not (a or b);
    layer0_outputs(940) <= b;
    layer0_outputs(941) <= a or b;
    layer0_outputs(942) <= a or b;
    layer0_outputs(943) <= not (a or b);
    layer0_outputs(944) <= 1'b0;
    layer0_outputs(945) <= not (a or b);
    layer0_outputs(946) <= not (a or b);
    layer0_outputs(947) <= a xor b;
    layer0_outputs(948) <= not (a or b);
    layer0_outputs(949) <= not b;
    layer0_outputs(950) <= a xor b;
    layer0_outputs(951) <= not b;
    layer0_outputs(952) <= not (a or b);
    layer0_outputs(953) <= a or b;
    layer0_outputs(954) <= a;
    layer0_outputs(955) <= a;
    layer0_outputs(956) <= not (a or b);
    layer0_outputs(957) <= a xor b;
    layer0_outputs(958) <= b and not a;
    layer0_outputs(959) <= not (a or b);
    layer0_outputs(960) <= a and not b;
    layer0_outputs(961) <= a or b;
    layer0_outputs(962) <= a;
    layer0_outputs(963) <= not b;
    layer0_outputs(964) <= not (a xor b);
    layer0_outputs(965) <= not (a or b);
    layer0_outputs(966) <= not a;
    layer0_outputs(967) <= b;
    layer0_outputs(968) <= not a or b;
    layer0_outputs(969) <= a xor b;
    layer0_outputs(970) <= b;
    layer0_outputs(971) <= not a or b;
    layer0_outputs(972) <= a or b;
    layer0_outputs(973) <= a xor b;
    layer0_outputs(974) <= not (a or b);
    layer0_outputs(975) <= not b or a;
    layer0_outputs(976) <= not (a xor b);
    layer0_outputs(977) <= a;
    layer0_outputs(978) <= b;
    layer0_outputs(979) <= b;
    layer0_outputs(980) <= a and not b;
    layer0_outputs(981) <= a xor b;
    layer0_outputs(982) <= a or b;
    layer0_outputs(983) <= a or b;
    layer0_outputs(984) <= not a or b;
    layer0_outputs(985) <= b;
    layer0_outputs(986) <= b;
    layer0_outputs(987) <= a or b;
    layer0_outputs(988) <= a or b;
    layer0_outputs(989) <= a or b;
    layer0_outputs(990) <= a;
    layer0_outputs(991) <= b and not a;
    layer0_outputs(992) <= not b or a;
    layer0_outputs(993) <= not a or b;
    layer0_outputs(994) <= not (a xor b);
    layer0_outputs(995) <= a or b;
    layer0_outputs(996) <= not (a or b);
    layer0_outputs(997) <= b;
    layer0_outputs(998) <= a;
    layer0_outputs(999) <= a or b;
    layer0_outputs(1000) <= a or b;
    layer0_outputs(1001) <= not a or b;
    layer0_outputs(1002) <= not (a or b);
    layer0_outputs(1003) <= not (a or b);
    layer0_outputs(1004) <= not (a or b);
    layer0_outputs(1005) <= not b;
    layer0_outputs(1006) <= a or b;
    layer0_outputs(1007) <= a;
    layer0_outputs(1008) <= not a or b;
    layer0_outputs(1009) <= a or b;
    layer0_outputs(1010) <= not (a xor b);
    layer0_outputs(1011) <= not (a or b);
    layer0_outputs(1012) <= b;
    layer0_outputs(1013) <= not a;
    layer0_outputs(1014) <= not b or a;
    layer0_outputs(1015) <= a xor b;
    layer0_outputs(1016) <= not (a xor b);
    layer0_outputs(1017) <= 1'b1;
    layer0_outputs(1018) <= not (a xor b);
    layer0_outputs(1019) <= not (a and b);
    layer0_outputs(1020) <= b;
    layer0_outputs(1021) <= not a;
    layer0_outputs(1022) <= not b;
    layer0_outputs(1023) <= b;
    layer0_outputs(1024) <= a and not b;
    layer0_outputs(1025) <= a;
    layer0_outputs(1026) <= a and not b;
    layer0_outputs(1027) <= not (a or b);
    layer0_outputs(1028) <= a and not b;
    layer0_outputs(1029) <= a xor b;
    layer0_outputs(1030) <= b;
    layer0_outputs(1031) <= a;
    layer0_outputs(1032) <= not b;
    layer0_outputs(1033) <= not a;
    layer0_outputs(1034) <= b and not a;
    layer0_outputs(1035) <= not (a or b);
    layer0_outputs(1036) <= not (a or b);
    layer0_outputs(1037) <= not (a xor b);
    layer0_outputs(1038) <= not (a xor b);
    layer0_outputs(1039) <= 1'b0;
    layer0_outputs(1040) <= a xor b;
    layer0_outputs(1041) <= not (a or b);
    layer0_outputs(1042) <= not a or b;
    layer0_outputs(1043) <= b;
    layer0_outputs(1044) <= a and not b;
    layer0_outputs(1045) <= not b;
    layer0_outputs(1046) <= a and b;
    layer0_outputs(1047) <= not (a or b);
    layer0_outputs(1048) <= not (a and b);
    layer0_outputs(1049) <= a and not b;
    layer0_outputs(1050) <= a or b;
    layer0_outputs(1051) <= not (a xor b);
    layer0_outputs(1052) <= a or b;
    layer0_outputs(1053) <= a and not b;
    layer0_outputs(1054) <= not b;
    layer0_outputs(1055) <= a;
    layer0_outputs(1056) <= b and not a;
    layer0_outputs(1057) <= not a or b;
    layer0_outputs(1058) <= not b or a;
    layer0_outputs(1059) <= a or b;
    layer0_outputs(1060) <= 1'b0;
    layer0_outputs(1061) <= not b;
    layer0_outputs(1062) <= b;
    layer0_outputs(1063) <= b and not a;
    layer0_outputs(1064) <= not (a xor b);
    layer0_outputs(1065) <= not a;
    layer0_outputs(1066) <= a or b;
    layer0_outputs(1067) <= a or b;
    layer0_outputs(1068) <= b and not a;
    layer0_outputs(1069) <= a xor b;
    layer0_outputs(1070) <= a xor b;
    layer0_outputs(1071) <= a or b;
    layer0_outputs(1072) <= a or b;
    layer0_outputs(1073) <= a or b;
    layer0_outputs(1074) <= a xor b;
    layer0_outputs(1075) <= not (a or b);
    layer0_outputs(1076) <= not (a or b);
    layer0_outputs(1077) <= a or b;
    layer0_outputs(1078) <= a or b;
    layer0_outputs(1079) <= a or b;
    layer0_outputs(1080) <= not a;
    layer0_outputs(1081) <= a or b;
    layer0_outputs(1082) <= a or b;
    layer0_outputs(1083) <= 1'b0;
    layer0_outputs(1084) <= b and not a;
    layer0_outputs(1085) <= not a or b;
    layer0_outputs(1086) <= not (a xor b);
    layer0_outputs(1087) <= a;
    layer0_outputs(1088) <= a xor b;
    layer0_outputs(1089) <= not b;
    layer0_outputs(1090) <= a and not b;
    layer0_outputs(1091) <= not (a xor b);
    layer0_outputs(1092) <= a xor b;
    layer0_outputs(1093) <= a xor b;
    layer0_outputs(1094) <= not b or a;
    layer0_outputs(1095) <= a;
    layer0_outputs(1096) <= not b;
    layer0_outputs(1097) <= not (a xor b);
    layer0_outputs(1098) <= not (a xor b);
    layer0_outputs(1099) <= not (a or b);
    layer0_outputs(1100) <= not (a or b);
    layer0_outputs(1101) <= a xor b;
    layer0_outputs(1102) <= 1'b1;
    layer0_outputs(1103) <= a and not b;
    layer0_outputs(1104) <= a or b;
    layer0_outputs(1105) <= b;
    layer0_outputs(1106) <= not b;
    layer0_outputs(1107) <= b and not a;
    layer0_outputs(1108) <= not (a xor b);
    layer0_outputs(1109) <= not (a or b);
    layer0_outputs(1110) <= not b;
    layer0_outputs(1111) <= a xor b;
    layer0_outputs(1112) <= a;
    layer0_outputs(1113) <= a or b;
    layer0_outputs(1114) <= not (a xor b);
    layer0_outputs(1115) <= a or b;
    layer0_outputs(1116) <= not a;
    layer0_outputs(1117) <= b;
    layer0_outputs(1118) <= a and not b;
    layer0_outputs(1119) <= b and not a;
    layer0_outputs(1120) <= not (a or b);
    layer0_outputs(1121) <= not b or a;
    layer0_outputs(1122) <= a and not b;
    layer0_outputs(1123) <= not a;
    layer0_outputs(1124) <= not (a xor b);
    layer0_outputs(1125) <= not (a or b);
    layer0_outputs(1126) <= not (a xor b);
    layer0_outputs(1127) <= b and not a;
    layer0_outputs(1128) <= not b;
    layer0_outputs(1129) <= not b;
    layer0_outputs(1130) <= a or b;
    layer0_outputs(1131) <= a and not b;
    layer0_outputs(1132) <= not (a or b);
    layer0_outputs(1133) <= not (a xor b);
    layer0_outputs(1134) <= a and not b;
    layer0_outputs(1135) <= b and not a;
    layer0_outputs(1136) <= a xor b;
    layer0_outputs(1137) <= 1'b1;
    layer0_outputs(1138) <= not (a or b);
    layer0_outputs(1139) <= b and not a;
    layer0_outputs(1140) <= not (a or b);
    layer0_outputs(1141) <= not a or b;
    layer0_outputs(1142) <= a;
    layer0_outputs(1143) <= not a;
    layer0_outputs(1144) <= not (a or b);
    layer0_outputs(1145) <= not b or a;
    layer0_outputs(1146) <= not a or b;
    layer0_outputs(1147) <= a and not b;
    layer0_outputs(1148) <= a xor b;
    layer0_outputs(1149) <= not a or b;
    layer0_outputs(1150) <= a or b;
    layer0_outputs(1151) <= not a or b;
    layer0_outputs(1152) <= a or b;
    layer0_outputs(1153) <= b and not a;
    layer0_outputs(1154) <= b and not a;
    layer0_outputs(1155) <= a;
    layer0_outputs(1156) <= a;
    layer0_outputs(1157) <= b and not a;
    layer0_outputs(1158) <= not b or a;
    layer0_outputs(1159) <= not b;
    layer0_outputs(1160) <= not b;
    layer0_outputs(1161) <= not (a or b);
    layer0_outputs(1162) <= a or b;
    layer0_outputs(1163) <= not a;
    layer0_outputs(1164) <= not b or a;
    layer0_outputs(1165) <= b and not a;
    layer0_outputs(1166) <= a or b;
    layer0_outputs(1167) <= not b;
    layer0_outputs(1168) <= not a;
    layer0_outputs(1169) <= a or b;
    layer0_outputs(1170) <= b;
    layer0_outputs(1171) <= 1'b0;
    layer0_outputs(1172) <= not (a or b);
    layer0_outputs(1173) <= not (a xor b);
    layer0_outputs(1174) <= not b or a;
    layer0_outputs(1175) <= not (a xor b);
    layer0_outputs(1176) <= a and not b;
    layer0_outputs(1177) <= not a or b;
    layer0_outputs(1178) <= 1'b1;
    layer0_outputs(1179) <= not (a or b);
    layer0_outputs(1180) <= a or b;
    layer0_outputs(1181) <= a xor b;
    layer0_outputs(1182) <= not (a or b);
    layer0_outputs(1183) <= a or b;
    layer0_outputs(1184) <= a;
    layer0_outputs(1185) <= not (a xor b);
    layer0_outputs(1186) <= not (a or b);
    layer0_outputs(1187) <= not b;
    layer0_outputs(1188) <= not (a or b);
    layer0_outputs(1189) <= not (a xor b);
    layer0_outputs(1190) <= not (a or b);
    layer0_outputs(1191) <= not (a or b);
    layer0_outputs(1192) <= a or b;
    layer0_outputs(1193) <= 1'b1;
    layer0_outputs(1194) <= not a;
    layer0_outputs(1195) <= a and not b;
    layer0_outputs(1196) <= a;
    layer0_outputs(1197) <= b;
    layer0_outputs(1198) <= 1'b0;
    layer0_outputs(1199) <= a xor b;
    layer0_outputs(1200) <= not a;
    layer0_outputs(1201) <= not (a xor b);
    layer0_outputs(1202) <= b;
    layer0_outputs(1203) <= a and not b;
    layer0_outputs(1204) <= not a;
    layer0_outputs(1205) <= a xor b;
    layer0_outputs(1206) <= a xor b;
    layer0_outputs(1207) <= b;
    layer0_outputs(1208) <= not (a or b);
    layer0_outputs(1209) <= not (a and b);
    layer0_outputs(1210) <= not b or a;
    layer0_outputs(1211) <= a;
    layer0_outputs(1212) <= not b or a;
    layer0_outputs(1213) <= b;
    layer0_outputs(1214) <= not b;
    layer0_outputs(1215) <= not b or a;
    layer0_outputs(1216) <= a or b;
    layer0_outputs(1217) <= a or b;
    layer0_outputs(1218) <= not a;
    layer0_outputs(1219) <= a or b;
    layer0_outputs(1220) <= a and not b;
    layer0_outputs(1221) <= a and not b;
    layer0_outputs(1222) <= a or b;
    layer0_outputs(1223) <= not (a xor b);
    layer0_outputs(1224) <= not a;
    layer0_outputs(1225) <= not (a or b);
    layer0_outputs(1226) <= a or b;
    layer0_outputs(1227) <= b and not a;
    layer0_outputs(1228) <= not (a or b);
    layer0_outputs(1229) <= a or b;
    layer0_outputs(1230) <= not b;
    layer0_outputs(1231) <= a or b;
    layer0_outputs(1232) <= not (a xor b);
    layer0_outputs(1233) <= not (a or b);
    layer0_outputs(1234) <= not (a xor b);
    layer0_outputs(1235) <= a xor b;
    layer0_outputs(1236) <= b and not a;
    layer0_outputs(1237) <= not b or a;
    layer0_outputs(1238) <= not (a xor b);
    layer0_outputs(1239) <= a xor b;
    layer0_outputs(1240) <= a xor b;
    layer0_outputs(1241) <= not (a or b);
    layer0_outputs(1242) <= a xor b;
    layer0_outputs(1243) <= not b;
    layer0_outputs(1244) <= not (a or b);
    layer0_outputs(1245) <= a or b;
    layer0_outputs(1246) <= not (a or b);
    layer0_outputs(1247) <= not a;
    layer0_outputs(1248) <= not (a or b);
    layer0_outputs(1249) <= b;
    layer0_outputs(1250) <= not b;
    layer0_outputs(1251) <= b;
    layer0_outputs(1252) <= not a;
    layer0_outputs(1253) <= not b or a;
    layer0_outputs(1254) <= b;
    layer0_outputs(1255) <= b and not a;
    layer0_outputs(1256) <= a or b;
    layer0_outputs(1257) <= not a or b;
    layer0_outputs(1258) <= not (a or b);
    layer0_outputs(1259) <= a or b;
    layer0_outputs(1260) <= a xor b;
    layer0_outputs(1261) <= not a;
    layer0_outputs(1262) <= a or b;
    layer0_outputs(1263) <= b;
    layer0_outputs(1264) <= not (a xor b);
    layer0_outputs(1265) <= a or b;
    layer0_outputs(1266) <= a or b;
    layer0_outputs(1267) <= a xor b;
    layer0_outputs(1268) <= not (a or b);
    layer0_outputs(1269) <= not b;
    layer0_outputs(1270) <= not b or a;
    layer0_outputs(1271) <= b and not a;
    layer0_outputs(1272) <= not (a or b);
    layer0_outputs(1273) <= a or b;
    layer0_outputs(1274) <= a and not b;
    layer0_outputs(1275) <= a xor b;
    layer0_outputs(1276) <= not (a or b);
    layer0_outputs(1277) <= a;
    layer0_outputs(1278) <= not b;
    layer0_outputs(1279) <= not b or a;
    layer0_outputs(1280) <= a xor b;
    layer0_outputs(1281) <= b and not a;
    layer0_outputs(1282) <= a or b;
    layer0_outputs(1283) <= not b or a;
    layer0_outputs(1284) <= a or b;
    layer0_outputs(1285) <= a xor b;
    layer0_outputs(1286) <= a or b;
    layer0_outputs(1287) <= 1'b1;
    layer0_outputs(1288) <= a;
    layer0_outputs(1289) <= a and b;
    layer0_outputs(1290) <= not (a or b);
    layer0_outputs(1291) <= not b or a;
    layer0_outputs(1292) <= not a;
    layer0_outputs(1293) <= a and not b;
    layer0_outputs(1294) <= a and not b;
    layer0_outputs(1295) <= not a;
    layer0_outputs(1296) <= 1'b0;
    layer0_outputs(1297) <= a and not b;
    layer0_outputs(1298) <= a or b;
    layer0_outputs(1299) <= not (a or b);
    layer0_outputs(1300) <= not a or b;
    layer0_outputs(1301) <= not (a or b);
    layer0_outputs(1302) <= b and not a;
    layer0_outputs(1303) <= not a;
    layer0_outputs(1304) <= not (a xor b);
    layer0_outputs(1305) <= 1'b1;
    layer0_outputs(1306) <= not a or b;
    layer0_outputs(1307) <= a or b;
    layer0_outputs(1308) <= not b or a;
    layer0_outputs(1309) <= a or b;
    layer0_outputs(1310) <= not a or b;
    layer0_outputs(1311) <= not (a and b);
    layer0_outputs(1312) <= not a;
    layer0_outputs(1313) <= b and not a;
    layer0_outputs(1314) <= not a;
    layer0_outputs(1315) <= not a or b;
    layer0_outputs(1316) <= b and not a;
    layer0_outputs(1317) <= a or b;
    layer0_outputs(1318) <= b and not a;
    layer0_outputs(1319) <= not (a xor b);
    layer0_outputs(1320) <= not (a or b);
    layer0_outputs(1321) <= a or b;
    layer0_outputs(1322) <= not (a xor b);
    layer0_outputs(1323) <= not (a and b);
    layer0_outputs(1324) <= not (a or b);
    layer0_outputs(1325) <= not a or b;
    layer0_outputs(1326) <= b and not a;
    layer0_outputs(1327) <= a;
    layer0_outputs(1328) <= not a;
    layer0_outputs(1329) <= b and not a;
    layer0_outputs(1330) <= not (a or b);
    layer0_outputs(1331) <= a or b;
    layer0_outputs(1332) <= b and not a;
    layer0_outputs(1333) <= not a;
    layer0_outputs(1334) <= a xor b;
    layer0_outputs(1335) <= not (a xor b);
    layer0_outputs(1336) <= not (a or b);
    layer0_outputs(1337) <= b;
    layer0_outputs(1338) <= a;
    layer0_outputs(1339) <= a or b;
    layer0_outputs(1340) <= not (a xor b);
    layer0_outputs(1341) <= not (a or b);
    layer0_outputs(1342) <= not (a xor b);
    layer0_outputs(1343) <= a;
    layer0_outputs(1344) <= a or b;
    layer0_outputs(1345) <= a or b;
    layer0_outputs(1346) <= not (a or b);
    layer0_outputs(1347) <= not b;
    layer0_outputs(1348) <= not a or b;
    layer0_outputs(1349) <= not (a or b);
    layer0_outputs(1350) <= not a;
    layer0_outputs(1351) <= a;
    layer0_outputs(1352) <= not a or b;
    layer0_outputs(1353) <= not a;
    layer0_outputs(1354) <= a or b;
    layer0_outputs(1355) <= 1'b1;
    layer0_outputs(1356) <= b and not a;
    layer0_outputs(1357) <= not b or a;
    layer0_outputs(1358) <= not (a xor b);
    layer0_outputs(1359) <= a and not b;
    layer0_outputs(1360) <= a;
    layer0_outputs(1361) <= not (a and b);
    layer0_outputs(1362) <= not (a or b);
    layer0_outputs(1363) <= not a;
    layer0_outputs(1364) <= a or b;
    layer0_outputs(1365) <= a xor b;
    layer0_outputs(1366) <= 1'b1;
    layer0_outputs(1367) <= not a or b;
    layer0_outputs(1368) <= a xor b;
    layer0_outputs(1369) <= not b or a;
    layer0_outputs(1370) <= b and not a;
    layer0_outputs(1371) <= not (a or b);
    layer0_outputs(1372) <= not a;
    layer0_outputs(1373) <= not (a or b);
    layer0_outputs(1374) <= a and not b;
    layer0_outputs(1375) <= not (a and b);
    layer0_outputs(1376) <= not b or a;
    layer0_outputs(1377) <= a xor b;
    layer0_outputs(1378) <= not (a or b);
    layer0_outputs(1379) <= not a or b;
    layer0_outputs(1380) <= a and not b;
    layer0_outputs(1381) <= a or b;
    layer0_outputs(1382) <= not a;
    layer0_outputs(1383) <= b;
    layer0_outputs(1384) <= not a or b;
    layer0_outputs(1385) <= a and b;
    layer0_outputs(1386) <= b and not a;
    layer0_outputs(1387) <= a or b;
    layer0_outputs(1388) <= a or b;
    layer0_outputs(1389) <= b and not a;
    layer0_outputs(1390) <= b and not a;
    layer0_outputs(1391) <= not b;
    layer0_outputs(1392) <= not (a or b);
    layer0_outputs(1393) <= not a;
    layer0_outputs(1394) <= a xor b;
    layer0_outputs(1395) <= not (a xor b);
    layer0_outputs(1396) <= a or b;
    layer0_outputs(1397) <= a or b;
    layer0_outputs(1398) <= a;
    layer0_outputs(1399) <= not a or b;
    layer0_outputs(1400) <= a or b;
    layer0_outputs(1401) <= a;
    layer0_outputs(1402) <= a;
    layer0_outputs(1403) <= not (a or b);
    layer0_outputs(1404) <= a xor b;
    layer0_outputs(1405) <= not (a or b);
    layer0_outputs(1406) <= not a;
    layer0_outputs(1407) <= a xor b;
    layer0_outputs(1408) <= not (a or b);
    layer0_outputs(1409) <= not (a or b);
    layer0_outputs(1410) <= not (a or b);
    layer0_outputs(1411) <= not b;
    layer0_outputs(1412) <= a;
    layer0_outputs(1413) <= a xor b;
    layer0_outputs(1414) <= a xor b;
    layer0_outputs(1415) <= not (a or b);
    layer0_outputs(1416) <= a;
    layer0_outputs(1417) <= not b or a;
    layer0_outputs(1418) <= a or b;
    layer0_outputs(1419) <= b and not a;
    layer0_outputs(1420) <= not a;
    layer0_outputs(1421) <= not (a or b);
    layer0_outputs(1422) <= not (a or b);
    layer0_outputs(1423) <= b;
    layer0_outputs(1424) <= not (a xor b);
    layer0_outputs(1425) <= a or b;
    layer0_outputs(1426) <= a or b;
    layer0_outputs(1427) <= a and not b;
    layer0_outputs(1428) <= not b or a;
    layer0_outputs(1429) <= a or b;
    layer0_outputs(1430) <= a xor b;
    layer0_outputs(1431) <= not a;
    layer0_outputs(1432) <= not b;
    layer0_outputs(1433) <= not (a or b);
    layer0_outputs(1434) <= not b;
    layer0_outputs(1435) <= a or b;
    layer0_outputs(1436) <= 1'b1;
    layer0_outputs(1437) <= b;
    layer0_outputs(1438) <= not a;
    layer0_outputs(1439) <= a or b;
    layer0_outputs(1440) <= not a or b;
    layer0_outputs(1441) <= b and not a;
    layer0_outputs(1442) <= not a or b;
    layer0_outputs(1443) <= not (a xor b);
    layer0_outputs(1444) <= a or b;
    layer0_outputs(1445) <= not b or a;
    layer0_outputs(1446) <= not (a or b);
    layer0_outputs(1447) <= a and not b;
    layer0_outputs(1448) <= a and not b;
    layer0_outputs(1449) <= not b or a;
    layer0_outputs(1450) <= a;
    layer0_outputs(1451) <= not a or b;
    layer0_outputs(1452) <= b;
    layer0_outputs(1453) <= not (a xor b);
    layer0_outputs(1454) <= b;
    layer0_outputs(1455) <= not (a or b);
    layer0_outputs(1456) <= not (a or b);
    layer0_outputs(1457) <= a xor b;
    layer0_outputs(1458) <= b;
    layer0_outputs(1459) <= not (a or b);
    layer0_outputs(1460) <= a xor b;
    layer0_outputs(1461) <= a and b;
    layer0_outputs(1462) <= a and not b;
    layer0_outputs(1463) <= not a;
    layer0_outputs(1464) <= not b;
    layer0_outputs(1465) <= a xor b;
    layer0_outputs(1466) <= b;
    layer0_outputs(1467) <= not (a xor b);
    layer0_outputs(1468) <= not (a or b);
    layer0_outputs(1469) <= not (a or b);
    layer0_outputs(1470) <= a;
    layer0_outputs(1471) <= not (a and b);
    layer0_outputs(1472) <= not a;
    layer0_outputs(1473) <= b and not a;
    layer0_outputs(1474) <= not (a or b);
    layer0_outputs(1475) <= not a;
    layer0_outputs(1476) <= a or b;
    layer0_outputs(1477) <= a;
    layer0_outputs(1478) <= not (a or b);
    layer0_outputs(1479) <= 1'b1;
    layer0_outputs(1480) <= b and not a;
    layer0_outputs(1481) <= a or b;
    layer0_outputs(1482) <= not (a and b);
    layer0_outputs(1483) <= a and not b;
    layer0_outputs(1484) <= b;
    layer0_outputs(1485) <= not a or b;
    layer0_outputs(1486) <= a xor b;
    layer0_outputs(1487) <= a xor b;
    layer0_outputs(1488) <= a xor b;
    layer0_outputs(1489) <= a or b;
    layer0_outputs(1490) <= a xor b;
    layer0_outputs(1491) <= b and not a;
    layer0_outputs(1492) <= not b or a;
    layer0_outputs(1493) <= not a;
    layer0_outputs(1494) <= not (a or b);
    layer0_outputs(1495) <= not a;
    layer0_outputs(1496) <= a or b;
    layer0_outputs(1497) <= not b;
    layer0_outputs(1498) <= not (a or b);
    layer0_outputs(1499) <= a xor b;
    layer0_outputs(1500) <= not a or b;
    layer0_outputs(1501) <= not b or a;
    layer0_outputs(1502) <= not a or b;
    layer0_outputs(1503) <= not a;
    layer0_outputs(1504) <= b and not a;
    layer0_outputs(1505) <= a;
    layer0_outputs(1506) <= a or b;
    layer0_outputs(1507) <= not b or a;
    layer0_outputs(1508) <= not a or b;
    layer0_outputs(1509) <= a;
    layer0_outputs(1510) <= not (a and b);
    layer0_outputs(1511) <= 1'b0;
    layer0_outputs(1512) <= a and not b;
    layer0_outputs(1513) <= a or b;
    layer0_outputs(1514) <= not (a or b);
    layer0_outputs(1515) <= a xor b;
    layer0_outputs(1516) <= a xor b;
    layer0_outputs(1517) <= a or b;
    layer0_outputs(1518) <= b and not a;
    layer0_outputs(1519) <= not a or b;
    layer0_outputs(1520) <= a xor b;
    layer0_outputs(1521) <= not (a or b);
    layer0_outputs(1522) <= b and not a;
    layer0_outputs(1523) <= b;
    layer0_outputs(1524) <= 1'b1;
    layer0_outputs(1525) <= a;
    layer0_outputs(1526) <= not b or a;
    layer0_outputs(1527) <= a or b;
    layer0_outputs(1528) <= a or b;
    layer0_outputs(1529) <= not (a xor b);
    layer0_outputs(1530) <= not b;
    layer0_outputs(1531) <= b;
    layer0_outputs(1532) <= not a;
    layer0_outputs(1533) <= not a;
    layer0_outputs(1534) <= a xor b;
    layer0_outputs(1535) <= not b;
    layer0_outputs(1536) <= a xor b;
    layer0_outputs(1537) <= not (a xor b);
    layer0_outputs(1538) <= a or b;
    layer0_outputs(1539) <= not a;
    layer0_outputs(1540) <= not b or a;
    layer0_outputs(1541) <= a and not b;
    layer0_outputs(1542) <= not (a xor b);
    layer0_outputs(1543) <= not (a xor b);
    layer0_outputs(1544) <= not b;
    layer0_outputs(1545) <= not b or a;
    layer0_outputs(1546) <= not (a xor b);
    layer0_outputs(1547) <= not (a or b);
    layer0_outputs(1548) <= a xor b;
    layer0_outputs(1549) <= not b or a;
    layer0_outputs(1550) <= a;
    layer0_outputs(1551) <= a and not b;
    layer0_outputs(1552) <= not b or a;
    layer0_outputs(1553) <= a or b;
    layer0_outputs(1554) <= a or b;
    layer0_outputs(1555) <= a or b;
    layer0_outputs(1556) <= a;
    layer0_outputs(1557) <= b;
    layer0_outputs(1558) <= not a or b;
    layer0_outputs(1559) <= a and not b;
    layer0_outputs(1560) <= not (a or b);
    layer0_outputs(1561) <= not (a or b);
    layer0_outputs(1562) <= not b or a;
    layer0_outputs(1563) <= not (a or b);
    layer0_outputs(1564) <= not (a or b);
    layer0_outputs(1565) <= not b;
    layer0_outputs(1566) <= a and b;
    layer0_outputs(1567) <= a xor b;
    layer0_outputs(1568) <= a or b;
    layer0_outputs(1569) <= not a or b;
    layer0_outputs(1570) <= a xor b;
    layer0_outputs(1571) <= a;
    layer0_outputs(1572) <= a or b;
    layer0_outputs(1573) <= a or b;
    layer0_outputs(1574) <= a;
    layer0_outputs(1575) <= not a or b;
    layer0_outputs(1576) <= not (a xor b);
    layer0_outputs(1577) <= not b;
    layer0_outputs(1578) <= b and not a;
    layer0_outputs(1579) <= a or b;
    layer0_outputs(1580) <= a;
    layer0_outputs(1581) <= not b or a;
    layer0_outputs(1582) <= b and not a;
    layer0_outputs(1583) <= b and not a;
    layer0_outputs(1584) <= b and not a;
    layer0_outputs(1585) <= a or b;
    layer0_outputs(1586) <= not (a or b);
    layer0_outputs(1587) <= 1'b1;
    layer0_outputs(1588) <= a or b;
    layer0_outputs(1589) <= not b or a;
    layer0_outputs(1590) <= not (a xor b);
    layer0_outputs(1591) <= a or b;
    layer0_outputs(1592) <= not b or a;
    layer0_outputs(1593) <= a and not b;
    layer0_outputs(1594) <= not (a or b);
    layer0_outputs(1595) <= a or b;
    layer0_outputs(1596) <= a and b;
    layer0_outputs(1597) <= b;
    layer0_outputs(1598) <= not b or a;
    layer0_outputs(1599) <= not (a or b);
    layer0_outputs(1600) <= a and not b;
    layer0_outputs(1601) <= a xor b;
    layer0_outputs(1602) <= not b;
    layer0_outputs(1603) <= not (a xor b);
    layer0_outputs(1604) <= a or b;
    layer0_outputs(1605) <= not b;
    layer0_outputs(1606) <= not b or a;
    layer0_outputs(1607) <= not b;
    layer0_outputs(1608) <= a or b;
    layer0_outputs(1609) <= not (a xor b);
    layer0_outputs(1610) <= not (a and b);
    layer0_outputs(1611) <= not a;
    layer0_outputs(1612) <= not (a xor b);
    layer0_outputs(1613) <= a;
    layer0_outputs(1614) <= not (a or b);
    layer0_outputs(1615) <= a xor b;
    layer0_outputs(1616) <= b;
    layer0_outputs(1617) <= b;
    layer0_outputs(1618) <= a and b;
    layer0_outputs(1619) <= not (a xor b);
    layer0_outputs(1620) <= not a or b;
    layer0_outputs(1621) <= a;
    layer0_outputs(1622) <= b;
    layer0_outputs(1623) <= a;
    layer0_outputs(1624) <= a or b;
    layer0_outputs(1625) <= 1'b1;
    layer0_outputs(1626) <= not a;
    layer0_outputs(1627) <= not (a xor b);
    layer0_outputs(1628) <= b and not a;
    layer0_outputs(1629) <= a and not b;
    layer0_outputs(1630) <= b and not a;
    layer0_outputs(1631) <= not b or a;
    layer0_outputs(1632) <= a or b;
    layer0_outputs(1633) <= a xor b;
    layer0_outputs(1634) <= not b;
    layer0_outputs(1635) <= not (a or b);
    layer0_outputs(1636) <= not (a xor b);
    layer0_outputs(1637) <= not a or b;
    layer0_outputs(1638) <= a;
    layer0_outputs(1639) <= a or b;
    layer0_outputs(1640) <= not (a xor b);
    layer0_outputs(1641) <= not (a and b);
    layer0_outputs(1642) <= not a;
    layer0_outputs(1643) <= not (a or b);
    layer0_outputs(1644) <= not b;
    layer0_outputs(1645) <= not a or b;
    layer0_outputs(1646) <= not (a or b);
    layer0_outputs(1647) <= not a or b;
    layer0_outputs(1648) <= b and not a;
    layer0_outputs(1649) <= not (a or b);
    layer0_outputs(1650) <= a or b;
    layer0_outputs(1651) <= not a or b;
    layer0_outputs(1652) <= b and not a;
    layer0_outputs(1653) <= not a;
    layer0_outputs(1654) <= a xor b;
    layer0_outputs(1655) <= not b;
    layer0_outputs(1656) <= not (a or b);
    layer0_outputs(1657) <= not (a xor b);
    layer0_outputs(1658) <= a and b;
    layer0_outputs(1659) <= a or b;
    layer0_outputs(1660) <= a and not b;
    layer0_outputs(1661) <= not (a or b);
    layer0_outputs(1662) <= a or b;
    layer0_outputs(1663) <= not b or a;
    layer0_outputs(1664) <= a xor b;
    layer0_outputs(1665) <= a;
    layer0_outputs(1666) <= b and not a;
    layer0_outputs(1667) <= a and not b;
    layer0_outputs(1668) <= b;
    layer0_outputs(1669) <= b and not a;
    layer0_outputs(1670) <= a;
    layer0_outputs(1671) <= not b;
    layer0_outputs(1672) <= not (a or b);
    layer0_outputs(1673) <= a xor b;
    layer0_outputs(1674) <= not b or a;
    layer0_outputs(1675) <= not a or b;
    layer0_outputs(1676) <= b and not a;
    layer0_outputs(1677) <= a and not b;
    layer0_outputs(1678) <= not (a or b);
    layer0_outputs(1679) <= a;
    layer0_outputs(1680) <= a and not b;
    layer0_outputs(1681) <= b and not a;
    layer0_outputs(1682) <= not b;
    layer0_outputs(1683) <= b;
    layer0_outputs(1684) <= a xor b;
    layer0_outputs(1685) <= not (a xor b);
    layer0_outputs(1686) <= a and not b;
    layer0_outputs(1687) <= not a or b;
    layer0_outputs(1688) <= not b or a;
    layer0_outputs(1689) <= a;
    layer0_outputs(1690) <= not b;
    layer0_outputs(1691) <= not b or a;
    layer0_outputs(1692) <= not b;
    layer0_outputs(1693) <= a or b;
    layer0_outputs(1694) <= b;
    layer0_outputs(1695) <= a or b;
    layer0_outputs(1696) <= not a or b;
    layer0_outputs(1697) <= not (a xor b);
    layer0_outputs(1698) <= not b or a;
    layer0_outputs(1699) <= not (a or b);
    layer0_outputs(1700) <= a and b;
    layer0_outputs(1701) <= a and not b;
    layer0_outputs(1702) <= not a or b;
    layer0_outputs(1703) <= b;
    layer0_outputs(1704) <= a or b;
    layer0_outputs(1705) <= not (a or b);
    layer0_outputs(1706) <= a xor b;
    layer0_outputs(1707) <= not b;
    layer0_outputs(1708) <= a and b;
    layer0_outputs(1709) <= not b;
    layer0_outputs(1710) <= a or b;
    layer0_outputs(1711) <= a and not b;
    layer0_outputs(1712) <= not (a xor b);
    layer0_outputs(1713) <= a or b;
    layer0_outputs(1714) <= not (a or b);
    layer0_outputs(1715) <= not b or a;
    layer0_outputs(1716) <= not (a xor b);
    layer0_outputs(1717) <= 1'b1;
    layer0_outputs(1718) <= not (a or b);
    layer0_outputs(1719) <= a;
    layer0_outputs(1720) <= not b or a;
    layer0_outputs(1721) <= not (a xor b);
    layer0_outputs(1722) <= not (a or b);
    layer0_outputs(1723) <= not b;
    layer0_outputs(1724) <= a;
    layer0_outputs(1725) <= not (a or b);
    layer0_outputs(1726) <= not a;
    layer0_outputs(1727) <= a or b;
    layer0_outputs(1728) <= not (a or b);
    layer0_outputs(1729) <= not a or b;
    layer0_outputs(1730) <= not (a xor b);
    layer0_outputs(1731) <= not a;
    layer0_outputs(1732) <= not b;
    layer0_outputs(1733) <= a or b;
    layer0_outputs(1734) <= not (a xor b);
    layer0_outputs(1735) <= b and not a;
    layer0_outputs(1736) <= b;
    layer0_outputs(1737) <= a or b;
    layer0_outputs(1738) <= b and not a;
    layer0_outputs(1739) <= a or b;
    layer0_outputs(1740) <= b and not a;
    layer0_outputs(1741) <= not (a xor b);
    layer0_outputs(1742) <= not b;
    layer0_outputs(1743) <= not (a or b);
    layer0_outputs(1744) <= 1'b0;
    layer0_outputs(1745) <= not a;
    layer0_outputs(1746) <= a or b;
    layer0_outputs(1747) <= not (a xor b);
    layer0_outputs(1748) <= a or b;
    layer0_outputs(1749) <= b;
    layer0_outputs(1750) <= not (a or b);
    layer0_outputs(1751) <= not b;
    layer0_outputs(1752) <= not (a or b);
    layer0_outputs(1753) <= a and not b;
    layer0_outputs(1754) <= a xor b;
    layer0_outputs(1755) <= not a;
    layer0_outputs(1756) <= a and not b;
    layer0_outputs(1757) <= not b;
    layer0_outputs(1758) <= 1'b0;
    layer0_outputs(1759) <= not (a xor b);
    layer0_outputs(1760) <= not a;
    layer0_outputs(1761) <= a;
    layer0_outputs(1762) <= 1'b1;
    layer0_outputs(1763) <= b and not a;
    layer0_outputs(1764) <= not b or a;
    layer0_outputs(1765) <= not (a or b);
    layer0_outputs(1766) <= a or b;
    layer0_outputs(1767) <= not b or a;
    layer0_outputs(1768) <= b and not a;
    layer0_outputs(1769) <= not (a or b);
    layer0_outputs(1770) <= a or b;
    layer0_outputs(1771) <= not (a or b);
    layer0_outputs(1772) <= a;
    layer0_outputs(1773) <= not (a or b);
    layer0_outputs(1774) <= not a;
    layer0_outputs(1775) <= a or b;
    layer0_outputs(1776) <= not (a or b);
    layer0_outputs(1777) <= not (a or b);
    layer0_outputs(1778) <= not a or b;
    layer0_outputs(1779) <= a or b;
    layer0_outputs(1780) <= not a or b;
    layer0_outputs(1781) <= b and not a;
    layer0_outputs(1782) <= a;
    layer0_outputs(1783) <= not (a xor b);
    layer0_outputs(1784) <= not b or a;
    layer0_outputs(1785) <= a and not b;
    layer0_outputs(1786) <= a and not b;
    layer0_outputs(1787) <= not (a xor b);
    layer0_outputs(1788) <= not (a xor b);
    layer0_outputs(1789) <= not b or a;
    layer0_outputs(1790) <= b and not a;
    layer0_outputs(1791) <= a;
    layer0_outputs(1792) <= a or b;
    layer0_outputs(1793) <= not b;
    layer0_outputs(1794) <= a or b;
    layer0_outputs(1795) <= a or b;
    layer0_outputs(1796) <= not b or a;
    layer0_outputs(1797) <= b and not a;
    layer0_outputs(1798) <= not b;
    layer0_outputs(1799) <= a and not b;
    layer0_outputs(1800) <= a;
    layer0_outputs(1801) <= 1'b1;
    layer0_outputs(1802) <= not a or b;
    layer0_outputs(1803) <= not a;
    layer0_outputs(1804) <= not a or b;
    layer0_outputs(1805) <= not (a or b);
    layer0_outputs(1806) <= not (a xor b);
    layer0_outputs(1807) <= not (a or b);
    layer0_outputs(1808) <= not (a xor b);
    layer0_outputs(1809) <= not (a or b);
    layer0_outputs(1810) <= a or b;
    layer0_outputs(1811) <= a;
    layer0_outputs(1812) <= a and not b;
    layer0_outputs(1813) <= a xor b;
    layer0_outputs(1814) <= b and not a;
    layer0_outputs(1815) <= a and not b;
    layer0_outputs(1816) <= a xor b;
    layer0_outputs(1817) <= not b or a;
    layer0_outputs(1818) <= not b or a;
    layer0_outputs(1819) <= not a or b;
    layer0_outputs(1820) <= not (a xor b);
    layer0_outputs(1821) <= not (a or b);
    layer0_outputs(1822) <= a or b;
    layer0_outputs(1823) <= a or b;
    layer0_outputs(1824) <= b and not a;
    layer0_outputs(1825) <= not b or a;
    layer0_outputs(1826) <= not (a or b);
    layer0_outputs(1827) <= not (a xor b);
    layer0_outputs(1828) <= not (a or b);
    layer0_outputs(1829) <= not a;
    layer0_outputs(1830) <= not (a xor b);
    layer0_outputs(1831) <= not (a or b);
    layer0_outputs(1832) <= b;
    layer0_outputs(1833) <= not b or a;
    layer0_outputs(1834) <= not (a or b);
    layer0_outputs(1835) <= a;
    layer0_outputs(1836) <= a or b;
    layer0_outputs(1837) <= not a or b;
    layer0_outputs(1838) <= not a;
    layer0_outputs(1839) <= not a or b;
    layer0_outputs(1840) <= a or b;
    layer0_outputs(1841) <= not b or a;
    layer0_outputs(1842) <= a and not b;
    layer0_outputs(1843) <= b;
    layer0_outputs(1844) <= not (a xor b);
    layer0_outputs(1845) <= b and not a;
    layer0_outputs(1846) <= a;
    layer0_outputs(1847) <= a;
    layer0_outputs(1848) <= b and not a;
    layer0_outputs(1849) <= not b;
    layer0_outputs(1850) <= b;
    layer0_outputs(1851) <= b;
    layer0_outputs(1852) <= b and not a;
    layer0_outputs(1853) <= not (a xor b);
    layer0_outputs(1854) <= 1'b0;
    layer0_outputs(1855) <= a or b;
    layer0_outputs(1856) <= a and not b;
    layer0_outputs(1857) <= a;
    layer0_outputs(1858) <= not a;
    layer0_outputs(1859) <= not (a or b);
    layer0_outputs(1860) <= a and not b;
    layer0_outputs(1861) <= not a or b;
    layer0_outputs(1862) <= a or b;
    layer0_outputs(1863) <= not (a or b);
    layer0_outputs(1864) <= not a or b;
    layer0_outputs(1865) <= a;
    layer0_outputs(1866) <= not (a xor b);
    layer0_outputs(1867) <= not a;
    layer0_outputs(1868) <= a and not b;
    layer0_outputs(1869) <= not (a xor b);
    layer0_outputs(1870) <= not (a or b);
    layer0_outputs(1871) <= not b;
    layer0_outputs(1872) <= a xor b;
    layer0_outputs(1873) <= a and not b;
    layer0_outputs(1874) <= not b;
    layer0_outputs(1875) <= not b or a;
    layer0_outputs(1876) <= not (a or b);
    layer0_outputs(1877) <= not b or a;
    layer0_outputs(1878) <= a xor b;
    layer0_outputs(1879) <= 1'b1;
    layer0_outputs(1880) <= a xor b;
    layer0_outputs(1881) <= a xor b;
    layer0_outputs(1882) <= a xor b;
    layer0_outputs(1883) <= not a;
    layer0_outputs(1884) <= b and not a;
    layer0_outputs(1885) <= not (a xor b);
    layer0_outputs(1886) <= not b;
    layer0_outputs(1887) <= not (a or b);
    layer0_outputs(1888) <= a;
    layer0_outputs(1889) <= not b or a;
    layer0_outputs(1890) <= not a or b;
    layer0_outputs(1891) <= a or b;
    layer0_outputs(1892) <= 1'b1;
    layer0_outputs(1893) <= a xor b;
    layer0_outputs(1894) <= not a or b;
    layer0_outputs(1895) <= b;
    layer0_outputs(1896) <= not b;
    layer0_outputs(1897) <= not (a or b);
    layer0_outputs(1898) <= 1'b0;
    layer0_outputs(1899) <= a or b;
    layer0_outputs(1900) <= not b;
    layer0_outputs(1901) <= not a;
    layer0_outputs(1902) <= not (a or b);
    layer0_outputs(1903) <= not b;
    layer0_outputs(1904) <= not b or a;
    layer0_outputs(1905) <= not (a or b);
    layer0_outputs(1906) <= a or b;
    layer0_outputs(1907) <= 1'b0;
    layer0_outputs(1908) <= not a;
    layer0_outputs(1909) <= a;
    layer0_outputs(1910) <= not b;
    layer0_outputs(1911) <= not (a xor b);
    layer0_outputs(1912) <= not b or a;
    layer0_outputs(1913) <= not a or b;
    layer0_outputs(1914) <= not (a or b);
    layer0_outputs(1915) <= a and not b;
    layer0_outputs(1916) <= b;
    layer0_outputs(1917) <= a xor b;
    layer0_outputs(1918) <= a;
    layer0_outputs(1919) <= not (a xor b);
    layer0_outputs(1920) <= not (a xor b);
    layer0_outputs(1921) <= a;
    layer0_outputs(1922) <= not (a xor b);
    layer0_outputs(1923) <= not (a and b);
    layer0_outputs(1924) <= a or b;
    layer0_outputs(1925) <= not a or b;
    layer0_outputs(1926) <= a or b;
    layer0_outputs(1927) <= not (a or b);
    layer0_outputs(1928) <= not (a xor b);
    layer0_outputs(1929) <= not b or a;
    layer0_outputs(1930) <= not b or a;
    layer0_outputs(1931) <= not b;
    layer0_outputs(1932) <= not b or a;
    layer0_outputs(1933) <= not b or a;
    layer0_outputs(1934) <= not b or a;
    layer0_outputs(1935) <= a;
    layer0_outputs(1936) <= not b or a;
    layer0_outputs(1937) <= b;
    layer0_outputs(1938) <= not (a or b);
    layer0_outputs(1939) <= not (a or b);
    layer0_outputs(1940) <= a and not b;
    layer0_outputs(1941) <= not (a xor b);
    layer0_outputs(1942) <= a xor b;
    layer0_outputs(1943) <= not (a or b);
    layer0_outputs(1944) <= not a or b;
    layer0_outputs(1945) <= a xor b;
    layer0_outputs(1946) <= not a or b;
    layer0_outputs(1947) <= not (a or b);
    layer0_outputs(1948) <= not a or b;
    layer0_outputs(1949) <= a xor b;
    layer0_outputs(1950) <= not a or b;
    layer0_outputs(1951) <= not (a xor b);
    layer0_outputs(1952) <= not b;
    layer0_outputs(1953) <= 1'b0;
    layer0_outputs(1954) <= a;
    layer0_outputs(1955) <= not a or b;
    layer0_outputs(1956) <= not (a and b);
    layer0_outputs(1957) <= a or b;
    layer0_outputs(1958) <= not a or b;
    layer0_outputs(1959) <= not (a or b);
    layer0_outputs(1960) <= a or b;
    layer0_outputs(1961) <= b and not a;
    layer0_outputs(1962) <= a and b;
    layer0_outputs(1963) <= a xor b;
    layer0_outputs(1964) <= a and not b;
    layer0_outputs(1965) <= a and b;
    layer0_outputs(1966) <= a xor b;
    layer0_outputs(1967) <= 1'b0;
    layer0_outputs(1968) <= a or b;
    layer0_outputs(1969) <= not (a xor b);
    layer0_outputs(1970) <= not b;
    layer0_outputs(1971) <= not a or b;
    layer0_outputs(1972) <= not b or a;
    layer0_outputs(1973) <= not b or a;
    layer0_outputs(1974) <= a xor b;
    layer0_outputs(1975) <= not (a or b);
    layer0_outputs(1976) <= a xor b;
    layer0_outputs(1977) <= a or b;
    layer0_outputs(1978) <= b and not a;
    layer0_outputs(1979) <= a and not b;
    layer0_outputs(1980) <= not a;
    layer0_outputs(1981) <= b and not a;
    layer0_outputs(1982) <= not a or b;
    layer0_outputs(1983) <= not b;
    layer0_outputs(1984) <= not (a or b);
    layer0_outputs(1985) <= b and not a;
    layer0_outputs(1986) <= not a;
    layer0_outputs(1987) <= a and not b;
    layer0_outputs(1988) <= a or b;
    layer0_outputs(1989) <= b and not a;
    layer0_outputs(1990) <= not a;
    layer0_outputs(1991) <= b and not a;
    layer0_outputs(1992) <= a;
    layer0_outputs(1993) <= not b or a;
    layer0_outputs(1994) <= not (a xor b);
    layer0_outputs(1995) <= a or b;
    layer0_outputs(1996) <= a xor b;
    layer0_outputs(1997) <= not (a or b);
    layer0_outputs(1998) <= b;
    layer0_outputs(1999) <= a;
    layer0_outputs(2000) <= not (a and b);
    layer0_outputs(2001) <= not (a or b);
    layer0_outputs(2002) <= not (a or b);
    layer0_outputs(2003) <= b and not a;
    layer0_outputs(2004) <= a or b;
    layer0_outputs(2005) <= not (a and b);
    layer0_outputs(2006) <= not b;
    layer0_outputs(2007) <= not b or a;
    layer0_outputs(2008) <= a xor b;
    layer0_outputs(2009) <= not a or b;
    layer0_outputs(2010) <= a xor b;
    layer0_outputs(2011) <= not a or b;
    layer0_outputs(2012) <= a xor b;
    layer0_outputs(2013) <= b and not a;
    layer0_outputs(2014) <= not a or b;
    layer0_outputs(2015) <= a xor b;
    layer0_outputs(2016) <= not a or b;
    layer0_outputs(2017) <= a or b;
    layer0_outputs(2018) <= not b or a;
    layer0_outputs(2019) <= a and not b;
    layer0_outputs(2020) <= a and b;
    layer0_outputs(2021) <= a;
    layer0_outputs(2022) <= not (a or b);
    layer0_outputs(2023) <= not (a or b);
    layer0_outputs(2024) <= a xor b;
    layer0_outputs(2025) <= b and not a;
    layer0_outputs(2026) <= a or b;
    layer0_outputs(2027) <= not b or a;
    layer0_outputs(2028) <= not b or a;
    layer0_outputs(2029) <= not (a or b);
    layer0_outputs(2030) <= not a or b;
    layer0_outputs(2031) <= a and not b;
    layer0_outputs(2032) <= not (a or b);
    layer0_outputs(2033) <= a xor b;
    layer0_outputs(2034) <= 1'b0;
    layer0_outputs(2035) <= b;
    layer0_outputs(2036) <= b;
    layer0_outputs(2037) <= not (a or b);
    layer0_outputs(2038) <= not (a or b);
    layer0_outputs(2039) <= not b;
    layer0_outputs(2040) <= not (a or b);
    layer0_outputs(2041) <= a or b;
    layer0_outputs(2042) <= a xor b;
    layer0_outputs(2043) <= a or b;
    layer0_outputs(2044) <= a;
    layer0_outputs(2045) <= a or b;
    layer0_outputs(2046) <= a xor b;
    layer0_outputs(2047) <= a or b;
    layer0_outputs(2048) <= not b;
    layer0_outputs(2049) <= not a;
    layer0_outputs(2050) <= not (a and b);
    layer0_outputs(2051) <= not a or b;
    layer0_outputs(2052) <= a;
    layer0_outputs(2053) <= b;
    layer0_outputs(2054) <= a or b;
    layer0_outputs(2055) <= a and not b;
    layer0_outputs(2056) <= not b;
    layer0_outputs(2057) <= a and b;
    layer0_outputs(2058) <= b;
    layer0_outputs(2059) <= b;
    layer0_outputs(2060) <= not (a or b);
    layer0_outputs(2061) <= not (a xor b);
    layer0_outputs(2062) <= not (a and b);
    layer0_outputs(2063) <= a or b;
    layer0_outputs(2064) <= b and not a;
    layer0_outputs(2065) <= a and not b;
    layer0_outputs(2066) <= not a or b;
    layer0_outputs(2067) <= not a;
    layer0_outputs(2068) <= a or b;
    layer0_outputs(2069) <= a and b;
    layer0_outputs(2070) <= a xor b;
    layer0_outputs(2071) <= b;
    layer0_outputs(2072) <= not (a or b);
    layer0_outputs(2073) <= not (a xor b);
    layer0_outputs(2074) <= a or b;
    layer0_outputs(2075) <= not (a xor b);
    layer0_outputs(2076) <= not b;
    layer0_outputs(2077) <= not (a or b);
    layer0_outputs(2078) <= a or b;
    layer0_outputs(2079) <= a xor b;
    layer0_outputs(2080) <= not b;
    layer0_outputs(2081) <= not (a xor b);
    layer0_outputs(2082) <= not (a or b);
    layer0_outputs(2083) <= not (a xor b);
    layer0_outputs(2084) <= b;
    layer0_outputs(2085) <= a and not b;
    layer0_outputs(2086) <= not a;
    layer0_outputs(2087) <= not a or b;
    layer0_outputs(2088) <= a xor b;
    layer0_outputs(2089) <= a;
    layer0_outputs(2090) <= a;
    layer0_outputs(2091) <= not (a or b);
    layer0_outputs(2092) <= a and not b;
    layer0_outputs(2093) <= not a or b;
    layer0_outputs(2094) <= a xor b;
    layer0_outputs(2095) <= b;
    layer0_outputs(2096) <= b and not a;
    layer0_outputs(2097) <= a xor b;
    layer0_outputs(2098) <= a xor b;
    layer0_outputs(2099) <= a or b;
    layer0_outputs(2100) <= not b;
    layer0_outputs(2101) <= not b or a;
    layer0_outputs(2102) <= a or b;
    layer0_outputs(2103) <= not a or b;
    layer0_outputs(2104) <= a or b;
    layer0_outputs(2105) <= a or b;
    layer0_outputs(2106) <= a xor b;
    layer0_outputs(2107) <= not a;
    layer0_outputs(2108) <= b and not a;
    layer0_outputs(2109) <= a;
    layer0_outputs(2110) <= b and not a;
    layer0_outputs(2111) <= b;
    layer0_outputs(2112) <= not b or a;
    layer0_outputs(2113) <= not b;
    layer0_outputs(2114) <= not (a xor b);
    layer0_outputs(2115) <= a;
    layer0_outputs(2116) <= b;
    layer0_outputs(2117) <= not b;
    layer0_outputs(2118) <= not a;
    layer0_outputs(2119) <= not (a xor b);
    layer0_outputs(2120) <= b and not a;
    layer0_outputs(2121) <= not b or a;
    layer0_outputs(2122) <= b and not a;
    layer0_outputs(2123) <= not (a or b);
    layer0_outputs(2124) <= 1'b1;
    layer0_outputs(2125) <= a or b;
    layer0_outputs(2126) <= a and not b;
    layer0_outputs(2127) <= b;
    layer0_outputs(2128) <= b and not a;
    layer0_outputs(2129) <= a xor b;
    layer0_outputs(2130) <= not b;
    layer0_outputs(2131) <= not a or b;
    layer0_outputs(2132) <= not a or b;
    layer0_outputs(2133) <= not b;
    layer0_outputs(2134) <= b;
    layer0_outputs(2135) <= a or b;
    layer0_outputs(2136) <= a and b;
    layer0_outputs(2137) <= a xor b;
    layer0_outputs(2138) <= a or b;
    layer0_outputs(2139) <= a and not b;
    layer0_outputs(2140) <= not (a or b);
    layer0_outputs(2141) <= a xor b;
    layer0_outputs(2142) <= a;
    layer0_outputs(2143) <= not (a and b);
    layer0_outputs(2144) <= not b;
    layer0_outputs(2145) <= a and not b;
    layer0_outputs(2146) <= a xor b;
    layer0_outputs(2147) <= not (a or b);
    layer0_outputs(2148) <= not b;
    layer0_outputs(2149) <= not b or a;
    layer0_outputs(2150) <= not a or b;
    layer0_outputs(2151) <= a or b;
    layer0_outputs(2152) <= not (a or b);
    layer0_outputs(2153) <= not b;
    layer0_outputs(2154) <= not (a or b);
    layer0_outputs(2155) <= not a or b;
    layer0_outputs(2156) <= b and not a;
    layer0_outputs(2157) <= not b;
    layer0_outputs(2158) <= not b;
    layer0_outputs(2159) <= a xor b;
    layer0_outputs(2160) <= not b;
    layer0_outputs(2161) <= 1'b1;
    layer0_outputs(2162) <= not (a xor b);
    layer0_outputs(2163) <= not (a xor b);
    layer0_outputs(2164) <= a and not b;
    layer0_outputs(2165) <= not a;
    layer0_outputs(2166) <= not a or b;
    layer0_outputs(2167) <= a xor b;
    layer0_outputs(2168) <= a;
    layer0_outputs(2169) <= b and not a;
    layer0_outputs(2170) <= not (a or b);
    layer0_outputs(2171) <= not (a or b);
    layer0_outputs(2172) <= not (a or b);
    layer0_outputs(2173) <= a;
    layer0_outputs(2174) <= a xor b;
    layer0_outputs(2175) <= a or b;
    layer0_outputs(2176) <= a or b;
    layer0_outputs(2177) <= b;
    layer0_outputs(2178) <= not b;
    layer0_outputs(2179) <= b;
    layer0_outputs(2180) <= 1'b1;
    layer0_outputs(2181) <= not (a or b);
    layer0_outputs(2182) <= a or b;
    layer0_outputs(2183) <= b;
    layer0_outputs(2184) <= not b or a;
    layer0_outputs(2185) <= not (a or b);
    layer0_outputs(2186) <= b and not a;
    layer0_outputs(2187) <= a or b;
    layer0_outputs(2188) <= a and not b;
    layer0_outputs(2189) <= a xor b;
    layer0_outputs(2190) <= not (a xor b);
    layer0_outputs(2191) <= not (a or b);
    layer0_outputs(2192) <= not (a xor b);
    layer0_outputs(2193) <= not b or a;
    layer0_outputs(2194) <= a xor b;
    layer0_outputs(2195) <= not b or a;
    layer0_outputs(2196) <= b and not a;
    layer0_outputs(2197) <= not (a or b);
    layer0_outputs(2198) <= not b or a;
    layer0_outputs(2199) <= not (a xor b);
    layer0_outputs(2200) <= a or b;
    layer0_outputs(2201) <= b and not a;
    layer0_outputs(2202) <= a or b;
    layer0_outputs(2203) <= not a or b;
    layer0_outputs(2204) <= a or b;
    layer0_outputs(2205) <= a or b;
    layer0_outputs(2206) <= not (a or b);
    layer0_outputs(2207) <= not b;
    layer0_outputs(2208) <= b and not a;
    layer0_outputs(2209) <= 1'b1;
    layer0_outputs(2210) <= not a or b;
    layer0_outputs(2211) <= a xor b;
    layer0_outputs(2212) <= a and not b;
    layer0_outputs(2213) <= b;
    layer0_outputs(2214) <= a xor b;
    layer0_outputs(2215) <= a xor b;
    layer0_outputs(2216) <= a xor b;
    layer0_outputs(2217) <= a or b;
    layer0_outputs(2218) <= b and not a;
    layer0_outputs(2219) <= a or b;
    layer0_outputs(2220) <= b and not a;
    layer0_outputs(2221) <= not (a or b);
    layer0_outputs(2222) <= a;
    layer0_outputs(2223) <= a;
    layer0_outputs(2224) <= a or b;
    layer0_outputs(2225) <= a xor b;
    layer0_outputs(2226) <= not (a or b);
    layer0_outputs(2227) <= a;
    layer0_outputs(2228) <= not (a or b);
    layer0_outputs(2229) <= a xor b;
    layer0_outputs(2230) <= a and not b;
    layer0_outputs(2231) <= a;
    layer0_outputs(2232) <= not (a xor b);
    layer0_outputs(2233) <= not a or b;
    layer0_outputs(2234) <= not b or a;
    layer0_outputs(2235) <= not a or b;
    layer0_outputs(2236) <= not (a or b);
    layer0_outputs(2237) <= not a or b;
    layer0_outputs(2238) <= not a or b;
    layer0_outputs(2239) <= a;
    layer0_outputs(2240) <= not (a or b);
    layer0_outputs(2241) <= b;
    layer0_outputs(2242) <= not b or a;
    layer0_outputs(2243) <= b and not a;
    layer0_outputs(2244) <= a or b;
    layer0_outputs(2245) <= not b;
    layer0_outputs(2246) <= a or b;
    layer0_outputs(2247) <= b and not a;
    layer0_outputs(2248) <= a or b;
    layer0_outputs(2249) <= a or b;
    layer0_outputs(2250) <= a or b;
    layer0_outputs(2251) <= not (a or b);
    layer0_outputs(2252) <= a or b;
    layer0_outputs(2253) <= not (a or b);
    layer0_outputs(2254) <= not (a xor b);
    layer0_outputs(2255) <= not (a or b);
    layer0_outputs(2256) <= not a or b;
    layer0_outputs(2257) <= not a;
    layer0_outputs(2258) <= not b or a;
    layer0_outputs(2259) <= not (a xor b);
    layer0_outputs(2260) <= 1'b0;
    layer0_outputs(2261) <= not a;
    layer0_outputs(2262) <= a xor b;
    layer0_outputs(2263) <= a and not b;
    layer0_outputs(2264) <= not (a or b);
    layer0_outputs(2265) <= a or b;
    layer0_outputs(2266) <= not (a xor b);
    layer0_outputs(2267) <= b and not a;
    layer0_outputs(2268) <= not (a or b);
    layer0_outputs(2269) <= a or b;
    layer0_outputs(2270) <= not a;
    layer0_outputs(2271) <= not a;
    layer0_outputs(2272) <= a;
    layer0_outputs(2273) <= not b or a;
    layer0_outputs(2274) <= not (a or b);
    layer0_outputs(2275) <= a or b;
    layer0_outputs(2276) <= not (a or b);
    layer0_outputs(2277) <= a xor b;
    layer0_outputs(2278) <= a or b;
    layer0_outputs(2279) <= not a or b;
    layer0_outputs(2280) <= not b or a;
    layer0_outputs(2281) <= a or b;
    layer0_outputs(2282) <= a or b;
    layer0_outputs(2283) <= a and not b;
    layer0_outputs(2284) <= a;
    layer0_outputs(2285) <= a or b;
    layer0_outputs(2286) <= not a or b;
    layer0_outputs(2287) <= b and not a;
    layer0_outputs(2288) <= not (a or b);
    layer0_outputs(2289) <= not b or a;
    layer0_outputs(2290) <= not (a xor b);
    layer0_outputs(2291) <= not (a xor b);
    layer0_outputs(2292) <= not (a or b);
    layer0_outputs(2293) <= a and not b;
    layer0_outputs(2294) <= a and not b;
    layer0_outputs(2295) <= not (a or b);
    layer0_outputs(2296) <= not (a and b);
    layer0_outputs(2297) <= not a;
    layer0_outputs(2298) <= a xor b;
    layer0_outputs(2299) <= a xor b;
    layer0_outputs(2300) <= a xor b;
    layer0_outputs(2301) <= b;
    layer0_outputs(2302) <= b;
    layer0_outputs(2303) <= a;
    layer0_outputs(2304) <= a;
    layer0_outputs(2305) <= a and not b;
    layer0_outputs(2306) <= not (a or b);
    layer0_outputs(2307) <= not a or b;
    layer0_outputs(2308) <= not a;
    layer0_outputs(2309) <= b and not a;
    layer0_outputs(2310) <= a or b;
    layer0_outputs(2311) <= a;
    layer0_outputs(2312) <= not (a and b);
    layer0_outputs(2313) <= b;
    layer0_outputs(2314) <= not (a xor b);
    layer0_outputs(2315) <= not (a xor b);
    layer0_outputs(2316) <= a xor b;
    layer0_outputs(2317) <= a or b;
    layer0_outputs(2318) <= b;
    layer0_outputs(2319) <= not (a xor b);
    layer0_outputs(2320) <= a;
    layer0_outputs(2321) <= not b or a;
    layer0_outputs(2322) <= b;
    layer0_outputs(2323) <= a and b;
    layer0_outputs(2324) <= a;
    layer0_outputs(2325) <= a or b;
    layer0_outputs(2326) <= not (a or b);
    layer0_outputs(2327) <= not (a and b);
    layer0_outputs(2328) <= b;
    layer0_outputs(2329) <= not a or b;
    layer0_outputs(2330) <= b;
    layer0_outputs(2331) <= not (a xor b);
    layer0_outputs(2332) <= b;
    layer0_outputs(2333) <= 1'b1;
    layer0_outputs(2334) <= not (a xor b);
    layer0_outputs(2335) <= a and b;
    layer0_outputs(2336) <= not (a or b);
    layer0_outputs(2337) <= a;
    layer0_outputs(2338) <= a and not b;
    layer0_outputs(2339) <= not (a or b);
    layer0_outputs(2340) <= not b;
    layer0_outputs(2341) <= a;
    layer0_outputs(2342) <= a;
    layer0_outputs(2343) <= not a or b;
    layer0_outputs(2344) <= not (a or b);
    layer0_outputs(2345) <= not (a or b);
    layer0_outputs(2346) <= not (a or b);
    layer0_outputs(2347) <= not b or a;
    layer0_outputs(2348) <= not a or b;
    layer0_outputs(2349) <= a or b;
    layer0_outputs(2350) <= not b;
    layer0_outputs(2351) <= 1'b1;
    layer0_outputs(2352) <= not a;
    layer0_outputs(2353) <= a;
    layer0_outputs(2354) <= not (a xor b);
    layer0_outputs(2355) <= not (a xor b);
    layer0_outputs(2356) <= not a;
    layer0_outputs(2357) <= not (a xor b);
    layer0_outputs(2358) <= not a;
    layer0_outputs(2359) <= 1'b0;
    layer0_outputs(2360) <= a or b;
    layer0_outputs(2361) <= not a or b;
    layer0_outputs(2362) <= a or b;
    layer0_outputs(2363) <= not b or a;
    layer0_outputs(2364) <= a or b;
    layer0_outputs(2365) <= a xor b;
    layer0_outputs(2366) <= not b or a;
    layer0_outputs(2367) <= not b;
    layer0_outputs(2368) <= not (a and b);
    layer0_outputs(2369) <= not (a or b);
    layer0_outputs(2370) <= not a or b;
    layer0_outputs(2371) <= a and not b;
    layer0_outputs(2372) <= not (a or b);
    layer0_outputs(2373) <= not a;
    layer0_outputs(2374) <= not (a or b);
    layer0_outputs(2375) <= b and not a;
    layer0_outputs(2376) <= a and b;
    layer0_outputs(2377) <= not (a or b);
    layer0_outputs(2378) <= a and b;
    layer0_outputs(2379) <= 1'b0;
    layer0_outputs(2380) <= not (a or b);
    layer0_outputs(2381) <= a or b;
    layer0_outputs(2382) <= a or b;
    layer0_outputs(2383) <= not (a xor b);
    layer0_outputs(2384) <= not (a xor b);
    layer0_outputs(2385) <= not (a xor b);
    layer0_outputs(2386) <= not (a or b);
    layer0_outputs(2387) <= a and not b;
    layer0_outputs(2388) <= not b;
    layer0_outputs(2389) <= b and not a;
    layer0_outputs(2390) <= b and not a;
    layer0_outputs(2391) <= a and not b;
    layer0_outputs(2392) <= a or b;
    layer0_outputs(2393) <= not (a or b);
    layer0_outputs(2394) <= a and b;
    layer0_outputs(2395) <= not (a xor b);
    layer0_outputs(2396) <= not a;
    layer0_outputs(2397) <= a and not b;
    layer0_outputs(2398) <= not b;
    layer0_outputs(2399) <= not a or b;
    layer0_outputs(2400) <= not (a xor b);
    layer0_outputs(2401) <= not a;
    layer0_outputs(2402) <= a or b;
    layer0_outputs(2403) <= a or b;
    layer0_outputs(2404) <= not b or a;
    layer0_outputs(2405) <= 1'b0;
    layer0_outputs(2406) <= a xor b;
    layer0_outputs(2407) <= not b or a;
    layer0_outputs(2408) <= 1'b0;
    layer0_outputs(2409) <= a xor b;
    layer0_outputs(2410) <= not a;
    layer0_outputs(2411) <= not (a xor b);
    layer0_outputs(2412) <= b;
    layer0_outputs(2413) <= a xor b;
    layer0_outputs(2414) <= a or b;
    layer0_outputs(2415) <= not b or a;
    layer0_outputs(2416) <= 1'b0;
    layer0_outputs(2417) <= not (a or b);
    layer0_outputs(2418) <= not b;
    layer0_outputs(2419) <= not (a or b);
    layer0_outputs(2420) <= not (a xor b);
    layer0_outputs(2421) <= a xor b;
    layer0_outputs(2422) <= not (a or b);
    layer0_outputs(2423) <= b;
    layer0_outputs(2424) <= b;
    layer0_outputs(2425) <= not b or a;
    layer0_outputs(2426) <= a or b;
    layer0_outputs(2427) <= b;
    layer0_outputs(2428) <= not (a xor b);
    layer0_outputs(2429) <= not a;
    layer0_outputs(2430) <= not (a or b);
    layer0_outputs(2431) <= not (a or b);
    layer0_outputs(2432) <= not (a xor b);
    layer0_outputs(2433) <= not (a xor b);
    layer0_outputs(2434) <= a and b;
    layer0_outputs(2435) <= not (a or b);
    layer0_outputs(2436) <= a or b;
    layer0_outputs(2437) <= b and not a;
    layer0_outputs(2438) <= a or b;
    layer0_outputs(2439) <= a and b;
    layer0_outputs(2440) <= not (a or b);
    layer0_outputs(2441) <= not (a or b);
    layer0_outputs(2442) <= b and not a;
    layer0_outputs(2443) <= not a or b;
    layer0_outputs(2444) <= b and not a;
    layer0_outputs(2445) <= not (a or b);
    layer0_outputs(2446) <= a;
    layer0_outputs(2447) <= a and b;
    layer0_outputs(2448) <= a or b;
    layer0_outputs(2449) <= a xor b;
    layer0_outputs(2450) <= b;
    layer0_outputs(2451) <= a or b;
    layer0_outputs(2452) <= not (a and b);
    layer0_outputs(2453) <= a or b;
    layer0_outputs(2454) <= a;
    layer0_outputs(2455) <= not (a or b);
    layer0_outputs(2456) <= not b or a;
    layer0_outputs(2457) <= not (a or b);
    layer0_outputs(2458) <= not b or a;
    layer0_outputs(2459) <= not b or a;
    layer0_outputs(2460) <= 1'b0;
    layer0_outputs(2461) <= not (a or b);
    layer0_outputs(2462) <= a;
    layer0_outputs(2463) <= not (a or b);
    layer0_outputs(2464) <= not a or b;
    layer0_outputs(2465) <= 1'b1;
    layer0_outputs(2466) <= not (a or b);
    layer0_outputs(2467) <= a or b;
    layer0_outputs(2468) <= not a;
    layer0_outputs(2469) <= not a or b;
    layer0_outputs(2470) <= a xor b;
    layer0_outputs(2471) <= a and b;
    layer0_outputs(2472) <= b;
    layer0_outputs(2473) <= a and not b;
    layer0_outputs(2474) <= a xor b;
    layer0_outputs(2475) <= not (a or b);
    layer0_outputs(2476) <= not (a xor b);
    layer0_outputs(2477) <= a or b;
    layer0_outputs(2478) <= 1'b1;
    layer0_outputs(2479) <= b;
    layer0_outputs(2480) <= not b;
    layer0_outputs(2481) <= not (a or b);
    layer0_outputs(2482) <= a xor b;
    layer0_outputs(2483) <= not a or b;
    layer0_outputs(2484) <= not b;
    layer0_outputs(2485) <= not b;
    layer0_outputs(2486) <= 1'b1;
    layer0_outputs(2487) <= a and b;
    layer0_outputs(2488) <= b and not a;
    layer0_outputs(2489) <= not b;
    layer0_outputs(2490) <= a and b;
    layer0_outputs(2491) <= not (a xor b);
    layer0_outputs(2492) <= not (a and b);
    layer0_outputs(2493) <= not b;
    layer0_outputs(2494) <= not (a or b);
    layer0_outputs(2495) <= a xor b;
    layer0_outputs(2496) <= a;
    layer0_outputs(2497) <= b and not a;
    layer0_outputs(2498) <= not a or b;
    layer0_outputs(2499) <= not (a or b);
    layer0_outputs(2500) <= not (a or b);
    layer0_outputs(2501) <= not b;
    layer0_outputs(2502) <= not (a xor b);
    layer0_outputs(2503) <= not (a or b);
    layer0_outputs(2504) <= a xor b;
    layer0_outputs(2505) <= not (a or b);
    layer0_outputs(2506) <= 1'b0;
    layer0_outputs(2507) <= a or b;
    layer0_outputs(2508) <= not a or b;
    layer0_outputs(2509) <= not b;
    layer0_outputs(2510) <= b and not a;
    layer0_outputs(2511) <= a and not b;
    layer0_outputs(2512) <= b;
    layer0_outputs(2513) <= b;
    layer0_outputs(2514) <= a and not b;
    layer0_outputs(2515) <= not (a xor b);
    layer0_outputs(2516) <= not a;
    layer0_outputs(2517) <= not a;
    layer0_outputs(2518) <= not a or b;
    layer0_outputs(2519) <= a;
    layer0_outputs(2520) <= b and not a;
    layer0_outputs(2521) <= a or b;
    layer0_outputs(2522) <= not (a xor b);
    layer0_outputs(2523) <= 1'b0;
    layer0_outputs(2524) <= a xor b;
    layer0_outputs(2525) <= a and not b;
    layer0_outputs(2526) <= a;
    layer0_outputs(2527) <= not (a and b);
    layer0_outputs(2528) <= b;
    layer0_outputs(2529) <= not (a xor b);
    layer0_outputs(2530) <= a or b;
    layer0_outputs(2531) <= not (a xor b);
    layer0_outputs(2532) <= 1'b1;
    layer0_outputs(2533) <= not a or b;
    layer0_outputs(2534) <= b and not a;
    layer0_outputs(2535) <= a;
    layer0_outputs(2536) <= not b or a;
    layer0_outputs(2537) <= not a or b;
    layer0_outputs(2538) <= not (a or b);
    layer0_outputs(2539) <= b and not a;
    layer0_outputs(2540) <= a xor b;
    layer0_outputs(2541) <= not (a or b);
    layer0_outputs(2542) <= not a;
    layer0_outputs(2543) <= a xor b;
    layer0_outputs(2544) <= not b;
    layer0_outputs(2545) <= not b;
    layer0_outputs(2546) <= not a or b;
    layer0_outputs(2547) <= not (a or b);
    layer0_outputs(2548) <= a and not b;
    layer0_outputs(2549) <= a xor b;
    layer0_outputs(2550) <= not b or a;
    layer0_outputs(2551) <= not (a or b);
    layer0_outputs(2552) <= not a or b;
    layer0_outputs(2553) <= a and not b;
    layer0_outputs(2554) <= b;
    layer0_outputs(2555) <= a xor b;
    layer0_outputs(2556) <= a xor b;
    layer0_outputs(2557) <= not b;
    layer0_outputs(2558) <= not b;
    layer0_outputs(2559) <= not (a or b);
    layer0_outputs(2560) <= 1'b0;
    layer0_outputs(2561) <= a or b;
    layer0_outputs(2562) <= not (a xor b);
    layer0_outputs(2563) <= not b or a;
    layer0_outputs(2564) <= not a or b;
    layer0_outputs(2565) <= not (a or b);
    layer0_outputs(2566) <= not (a xor b);
    layer0_outputs(2567) <= not (a or b);
    layer0_outputs(2568) <= b;
    layer0_outputs(2569) <= a xor b;
    layer0_outputs(2570) <= not (a xor b);
    layer0_outputs(2571) <= 1'b1;
    layer0_outputs(2572) <= 1'b1;
    layer0_outputs(2573) <= not a;
    layer0_outputs(2574) <= a or b;
    layer0_outputs(2575) <= not (a or b);
    layer0_outputs(2576) <= not b or a;
    layer0_outputs(2577) <= b;
    layer0_outputs(2578) <= a or b;
    layer0_outputs(2579) <= not (a or b);
    layer0_outputs(2580) <= not b or a;
    layer0_outputs(2581) <= a or b;
    layer0_outputs(2582) <= a xor b;
    layer0_outputs(2583) <= a or b;
    layer0_outputs(2584) <= a xor b;
    layer0_outputs(2585) <= a;
    layer0_outputs(2586) <= a xor b;
    layer0_outputs(2587) <= b and not a;
    layer0_outputs(2588) <= 1'b0;
    layer0_outputs(2589) <= a or b;
    layer0_outputs(2590) <= not (a xor b);
    layer0_outputs(2591) <= a or b;
    layer0_outputs(2592) <= a xor b;
    layer0_outputs(2593) <= not (a xor b);
    layer0_outputs(2594) <= b;
    layer0_outputs(2595) <= not (a or b);
    layer0_outputs(2596) <= 1'b0;
    layer0_outputs(2597) <= not a or b;
    layer0_outputs(2598) <= b and not a;
    layer0_outputs(2599) <= a and not b;
    layer0_outputs(2600) <= not (a or b);
    layer0_outputs(2601) <= a and not b;
    layer0_outputs(2602) <= not (a xor b);
    layer0_outputs(2603) <= not (a or b);
    layer0_outputs(2604) <= a and not b;
    layer0_outputs(2605) <= a;
    layer0_outputs(2606) <= not a or b;
    layer0_outputs(2607) <= b;
    layer0_outputs(2608) <= not a or b;
    layer0_outputs(2609) <= not (a xor b);
    layer0_outputs(2610) <= a and b;
    layer0_outputs(2611) <= not (a xor b);
    layer0_outputs(2612) <= not (a or b);
    layer0_outputs(2613) <= 1'b1;
    layer0_outputs(2614) <= not a or b;
    layer0_outputs(2615) <= a;
    layer0_outputs(2616) <= not a;
    layer0_outputs(2617) <= not (a and b);
    layer0_outputs(2618) <= b;
    layer0_outputs(2619) <= not (a xor b);
    layer0_outputs(2620) <= b;
    layer0_outputs(2621) <= 1'b1;
    layer0_outputs(2622) <= not (a or b);
    layer0_outputs(2623) <= not (a or b);
    layer0_outputs(2624) <= not a or b;
    layer0_outputs(2625) <= a or b;
    layer0_outputs(2626) <= a and not b;
    layer0_outputs(2627) <= not (a or b);
    layer0_outputs(2628) <= b;
    layer0_outputs(2629) <= a xor b;
    layer0_outputs(2630) <= not (a or b);
    layer0_outputs(2631) <= b and not a;
    layer0_outputs(2632) <= a or b;
    layer0_outputs(2633) <= b;
    layer0_outputs(2634) <= a xor b;
    layer0_outputs(2635) <= not b;
    layer0_outputs(2636) <= not a;
    layer0_outputs(2637) <= a or b;
    layer0_outputs(2638) <= not b;
    layer0_outputs(2639) <= not b;
    layer0_outputs(2640) <= not b;
    layer0_outputs(2641) <= not a or b;
    layer0_outputs(2642) <= a or b;
    layer0_outputs(2643) <= not b;
    layer0_outputs(2644) <= not a;
    layer0_outputs(2645) <= not (a or b);
    layer0_outputs(2646) <= b and not a;
    layer0_outputs(2647) <= not (a or b);
    layer0_outputs(2648) <= not (a xor b);
    layer0_outputs(2649) <= a or b;
    layer0_outputs(2650) <= 1'b0;
    layer0_outputs(2651) <= a xor b;
    layer0_outputs(2652) <= 1'b1;
    layer0_outputs(2653) <= not (a or b);
    layer0_outputs(2654) <= 1'b1;
    layer0_outputs(2655) <= not b;
    layer0_outputs(2656) <= not a or b;
    layer0_outputs(2657) <= not b;
    layer0_outputs(2658) <= not a;
    layer0_outputs(2659) <= a or b;
    layer0_outputs(2660) <= a xor b;
    layer0_outputs(2661) <= b;
    layer0_outputs(2662) <= not b;
    layer0_outputs(2663) <= a or b;
    layer0_outputs(2664) <= not (a xor b);
    layer0_outputs(2665) <= not b;
    layer0_outputs(2666) <= not b or a;
    layer0_outputs(2667) <= not (a xor b);
    layer0_outputs(2668) <= not (a xor b);
    layer0_outputs(2669) <= a xor b;
    layer0_outputs(2670) <= a or b;
    layer0_outputs(2671) <= not (a xor b);
    layer0_outputs(2672) <= 1'b0;
    layer0_outputs(2673) <= not a or b;
    layer0_outputs(2674) <= a xor b;
    layer0_outputs(2675) <= a;
    layer0_outputs(2676) <= a xor b;
    layer0_outputs(2677) <= a;
    layer0_outputs(2678) <= not (a xor b);
    layer0_outputs(2679) <= not a or b;
    layer0_outputs(2680) <= a xor b;
    layer0_outputs(2681) <= a;
    layer0_outputs(2682) <= not a;
    layer0_outputs(2683) <= b;
    layer0_outputs(2684) <= a or b;
    layer0_outputs(2685) <= not b or a;
    layer0_outputs(2686) <= a;
    layer0_outputs(2687) <= a and b;
    layer0_outputs(2688) <= a and b;
    layer0_outputs(2689) <= b;
    layer0_outputs(2690) <= not b;
    layer0_outputs(2691) <= not b;
    layer0_outputs(2692) <= a or b;
    layer0_outputs(2693) <= not (a xor b);
    layer0_outputs(2694) <= a xor b;
    layer0_outputs(2695) <= a or b;
    layer0_outputs(2696) <= not a;
    layer0_outputs(2697) <= not a or b;
    layer0_outputs(2698) <= b;
    layer0_outputs(2699) <= not (a or b);
    layer0_outputs(2700) <= b;
    layer0_outputs(2701) <= not (a or b);
    layer0_outputs(2702) <= not (a and b);
    layer0_outputs(2703) <= not (a xor b);
    layer0_outputs(2704) <= a and not b;
    layer0_outputs(2705) <= a xor b;
    layer0_outputs(2706) <= a and not b;
    layer0_outputs(2707) <= a;
    layer0_outputs(2708) <= a or b;
    layer0_outputs(2709) <= not (a xor b);
    layer0_outputs(2710) <= a xor b;
    layer0_outputs(2711) <= a;
    layer0_outputs(2712) <= b;
    layer0_outputs(2713) <= not (a and b);
    layer0_outputs(2714) <= not b;
    layer0_outputs(2715) <= not (a xor b);
    layer0_outputs(2716) <= a and b;
    layer0_outputs(2717) <= not a or b;
    layer0_outputs(2718) <= a xor b;
    layer0_outputs(2719) <= not b or a;
    layer0_outputs(2720) <= not (a xor b);
    layer0_outputs(2721) <= not a;
    layer0_outputs(2722) <= b;
    layer0_outputs(2723) <= not b or a;
    layer0_outputs(2724) <= a xor b;
    layer0_outputs(2725) <= not a or b;
    layer0_outputs(2726) <= a xor b;
    layer0_outputs(2727) <= a and not b;
    layer0_outputs(2728) <= not a;
    layer0_outputs(2729) <= 1'b0;
    layer0_outputs(2730) <= a;
    layer0_outputs(2731) <= a;
    layer0_outputs(2732) <= b;
    layer0_outputs(2733) <= a;
    layer0_outputs(2734) <= a or b;
    layer0_outputs(2735) <= not a or b;
    layer0_outputs(2736) <= 1'b0;
    layer0_outputs(2737) <= b;
    layer0_outputs(2738) <= not (a xor b);
    layer0_outputs(2739) <= not (a or b);
    layer0_outputs(2740) <= a and not b;
    layer0_outputs(2741) <= not b;
    layer0_outputs(2742) <= a or b;
    layer0_outputs(2743) <= b;
    layer0_outputs(2744) <= b;
    layer0_outputs(2745) <= a or b;
    layer0_outputs(2746) <= not (a or b);
    layer0_outputs(2747) <= not (a xor b);
    layer0_outputs(2748) <= a and not b;
    layer0_outputs(2749) <= a and not b;
    layer0_outputs(2750) <= not (a xor b);
    layer0_outputs(2751) <= not (a xor b);
    layer0_outputs(2752) <= not (a or b);
    layer0_outputs(2753) <= a xor b;
    layer0_outputs(2754) <= not a;
    layer0_outputs(2755) <= a or b;
    layer0_outputs(2756) <= not a;
    layer0_outputs(2757) <= not a;
    layer0_outputs(2758) <= not (a or b);
    layer0_outputs(2759) <= not (a xor b);
    layer0_outputs(2760) <= a and not b;
    layer0_outputs(2761) <= a;
    layer0_outputs(2762) <= b;
    layer0_outputs(2763) <= not b;
    layer0_outputs(2764) <= not (a or b);
    layer0_outputs(2765) <= b and not a;
    layer0_outputs(2766) <= not a;
    layer0_outputs(2767) <= not a;
    layer0_outputs(2768) <= not (a xor b);
    layer0_outputs(2769) <= not (a and b);
    layer0_outputs(2770) <= a or b;
    layer0_outputs(2771) <= b and not a;
    layer0_outputs(2772) <= not (a and b);
    layer0_outputs(2773) <= a xor b;
    layer0_outputs(2774) <= a or b;
    layer0_outputs(2775) <= not a;
    layer0_outputs(2776) <= a and not b;
    layer0_outputs(2777) <= a and not b;
    layer0_outputs(2778) <= not a;
    layer0_outputs(2779) <= not (a or b);
    layer0_outputs(2780) <= a;
    layer0_outputs(2781) <= not b;
    layer0_outputs(2782) <= a or b;
    layer0_outputs(2783) <= a;
    layer0_outputs(2784) <= a xor b;
    layer0_outputs(2785) <= not (a or b);
    layer0_outputs(2786) <= a and not b;
    layer0_outputs(2787) <= b;
    layer0_outputs(2788) <= not (a or b);
    layer0_outputs(2789) <= b;
    layer0_outputs(2790) <= a or b;
    layer0_outputs(2791) <= not a;
    layer0_outputs(2792) <= a or b;
    layer0_outputs(2793) <= a xor b;
    layer0_outputs(2794) <= not (a xor b);
    layer0_outputs(2795) <= not (a xor b);
    layer0_outputs(2796) <= b and not a;
    layer0_outputs(2797) <= a or b;
    layer0_outputs(2798) <= 1'b1;
    layer0_outputs(2799) <= not a;
    layer0_outputs(2800) <= a and not b;
    layer0_outputs(2801) <= not (a xor b);
    layer0_outputs(2802) <= a and b;
    layer0_outputs(2803) <= not b;
    layer0_outputs(2804) <= a xor b;
    layer0_outputs(2805) <= not (a xor b);
    layer0_outputs(2806) <= a xor b;
    layer0_outputs(2807) <= a or b;
    layer0_outputs(2808) <= not a or b;
    layer0_outputs(2809) <= a xor b;
    layer0_outputs(2810) <= a and not b;
    layer0_outputs(2811) <= not (a xor b);
    layer0_outputs(2812) <= not (a and b);
    layer0_outputs(2813) <= a and not b;
    layer0_outputs(2814) <= a or b;
    layer0_outputs(2815) <= not a;
    layer0_outputs(2816) <= not b;
    layer0_outputs(2817) <= a and not b;
    layer0_outputs(2818) <= not a;
    layer0_outputs(2819) <= not (a or b);
    layer0_outputs(2820) <= not a;
    layer0_outputs(2821) <= not (a or b);
    layer0_outputs(2822) <= a or b;
    layer0_outputs(2823) <= not b;
    layer0_outputs(2824) <= not a or b;
    layer0_outputs(2825) <= not a or b;
    layer0_outputs(2826) <= not b or a;
    layer0_outputs(2827) <= a and not b;
    layer0_outputs(2828) <= b;
    layer0_outputs(2829) <= not (a or b);
    layer0_outputs(2830) <= 1'b1;
    layer0_outputs(2831) <= not b;
    layer0_outputs(2832) <= not a;
    layer0_outputs(2833) <= 1'b0;
    layer0_outputs(2834) <= not (a xor b);
    layer0_outputs(2835) <= a;
    layer0_outputs(2836) <= a and not b;
    layer0_outputs(2837) <= not a or b;
    layer0_outputs(2838) <= a xor b;
    layer0_outputs(2839) <= b;
    layer0_outputs(2840) <= b;
    layer0_outputs(2841) <= not (a or b);
    layer0_outputs(2842) <= not (a or b);
    layer0_outputs(2843) <= b;
    layer0_outputs(2844) <= a and not b;
    layer0_outputs(2845) <= a xor b;
    layer0_outputs(2846) <= a xor b;
    layer0_outputs(2847) <= a xor b;
    layer0_outputs(2848) <= not a or b;
    layer0_outputs(2849) <= a or b;
    layer0_outputs(2850) <= a or b;
    layer0_outputs(2851) <= not (a xor b);
    layer0_outputs(2852) <= not (a or b);
    layer0_outputs(2853) <= b and not a;
    layer0_outputs(2854) <= not (a xor b);
    layer0_outputs(2855) <= not a or b;
    layer0_outputs(2856) <= a xor b;
    layer0_outputs(2857) <= not (a or b);
    layer0_outputs(2858) <= a and not b;
    layer0_outputs(2859) <= not (a or b);
    layer0_outputs(2860) <= not (a xor b);
    layer0_outputs(2861) <= a and not b;
    layer0_outputs(2862) <= not (a xor b);
    layer0_outputs(2863) <= a or b;
    layer0_outputs(2864) <= not (a or b);
    layer0_outputs(2865) <= not (a and b);
    layer0_outputs(2866) <= not (a or b);
    layer0_outputs(2867) <= not (a xor b);
    layer0_outputs(2868) <= a or b;
    layer0_outputs(2869) <= not a or b;
    layer0_outputs(2870) <= a and not b;
    layer0_outputs(2871) <= not b;
    layer0_outputs(2872) <= 1'b1;
    layer0_outputs(2873) <= not (a or b);
    layer0_outputs(2874) <= not (a xor b);
    layer0_outputs(2875) <= not b or a;
    layer0_outputs(2876) <= a and b;
    layer0_outputs(2877) <= not b;
    layer0_outputs(2878) <= b;
    layer0_outputs(2879) <= a;
    layer0_outputs(2880) <= a xor b;
    layer0_outputs(2881) <= a or b;
    layer0_outputs(2882) <= not b or a;
    layer0_outputs(2883) <= a and not b;
    layer0_outputs(2884) <= a;
    layer0_outputs(2885) <= a and not b;
    layer0_outputs(2886) <= not (a or b);
    layer0_outputs(2887) <= 1'b1;
    layer0_outputs(2888) <= a;
    layer0_outputs(2889) <= a or b;
    layer0_outputs(2890) <= b;
    layer0_outputs(2891) <= b and not a;
    layer0_outputs(2892) <= a or b;
    layer0_outputs(2893) <= 1'b0;
    layer0_outputs(2894) <= a or b;
    layer0_outputs(2895) <= a xor b;
    layer0_outputs(2896) <= a or b;
    layer0_outputs(2897) <= not b;
    layer0_outputs(2898) <= not a or b;
    layer0_outputs(2899) <= not b or a;
    layer0_outputs(2900) <= a and b;
    layer0_outputs(2901) <= not a or b;
    layer0_outputs(2902) <= a or b;
    layer0_outputs(2903) <= 1'b1;
    layer0_outputs(2904) <= a;
    layer0_outputs(2905) <= not b or a;
    layer0_outputs(2906) <= 1'b0;
    layer0_outputs(2907) <= a and not b;
    layer0_outputs(2908) <= b and not a;
    layer0_outputs(2909) <= a and b;
    layer0_outputs(2910) <= not (a or b);
    layer0_outputs(2911) <= not a or b;
    layer0_outputs(2912) <= not (a xor b);
    layer0_outputs(2913) <= a xor b;
    layer0_outputs(2914) <= b;
    layer0_outputs(2915) <= a and not b;
    layer0_outputs(2916) <= a or b;
    layer0_outputs(2917) <= a xor b;
    layer0_outputs(2918) <= b;
    layer0_outputs(2919) <= not (a or b);
    layer0_outputs(2920) <= b and not a;
    layer0_outputs(2921) <= not (a xor b);
    layer0_outputs(2922) <= a xor b;
    layer0_outputs(2923) <= a and not b;
    layer0_outputs(2924) <= not (a xor b);
    layer0_outputs(2925) <= not b or a;
    layer0_outputs(2926) <= not b;
    layer0_outputs(2927) <= b and not a;
    layer0_outputs(2928) <= a or b;
    layer0_outputs(2929) <= not (a or b);
    layer0_outputs(2930) <= not (a and b);
    layer0_outputs(2931) <= not b or a;
    layer0_outputs(2932) <= not b;
    layer0_outputs(2933) <= b;
    layer0_outputs(2934) <= 1'b1;
    layer0_outputs(2935) <= not b or a;
    layer0_outputs(2936) <= not b;
    layer0_outputs(2937) <= a or b;
    layer0_outputs(2938) <= not a;
    layer0_outputs(2939) <= a or b;
    layer0_outputs(2940) <= a;
    layer0_outputs(2941) <= not b or a;
    layer0_outputs(2942) <= a and not b;
    layer0_outputs(2943) <= b;
    layer0_outputs(2944) <= not b or a;
    layer0_outputs(2945) <= not a;
    layer0_outputs(2946) <= not a or b;
    layer0_outputs(2947) <= not a or b;
    layer0_outputs(2948) <= not (a or b);
    layer0_outputs(2949) <= a;
    layer0_outputs(2950) <= not b;
    layer0_outputs(2951) <= not (a and b);
    layer0_outputs(2952) <= a or b;
    layer0_outputs(2953) <= a or b;
    layer0_outputs(2954) <= a and not b;
    layer0_outputs(2955) <= not b or a;
    layer0_outputs(2956) <= b and not a;
    layer0_outputs(2957) <= a and not b;
    layer0_outputs(2958) <= not a;
    layer0_outputs(2959) <= b and not a;
    layer0_outputs(2960) <= a and not b;
    layer0_outputs(2961) <= a xor b;
    layer0_outputs(2962) <= not (a or b);
    layer0_outputs(2963) <= not a;
    layer0_outputs(2964) <= 1'b1;
    layer0_outputs(2965) <= not (a xor b);
    layer0_outputs(2966) <= a or b;
    layer0_outputs(2967) <= not (a or b);
    layer0_outputs(2968) <= a xor b;
    layer0_outputs(2969) <= not (a or b);
    layer0_outputs(2970) <= not (a or b);
    layer0_outputs(2971) <= not (a or b);
    layer0_outputs(2972) <= not b or a;
    layer0_outputs(2973) <= not (a xor b);
    layer0_outputs(2974) <= a xor b;
    layer0_outputs(2975) <= not (a or b);
    layer0_outputs(2976) <= not (a or b);
    layer0_outputs(2977) <= a xor b;
    layer0_outputs(2978) <= a or b;
    layer0_outputs(2979) <= not b;
    layer0_outputs(2980) <= b;
    layer0_outputs(2981) <= not (a or b);
    layer0_outputs(2982) <= not b;
    layer0_outputs(2983) <= not (a xor b);
    layer0_outputs(2984) <= a or b;
    layer0_outputs(2985) <= a;
    layer0_outputs(2986) <= b;
    layer0_outputs(2987) <= not a or b;
    layer0_outputs(2988) <= not (a or b);
    layer0_outputs(2989) <= a or b;
    layer0_outputs(2990) <= not (a or b);
    layer0_outputs(2991) <= not (a or b);
    layer0_outputs(2992) <= not (a or b);
    layer0_outputs(2993) <= a or b;
    layer0_outputs(2994) <= a or b;
    layer0_outputs(2995) <= not b or a;
    layer0_outputs(2996) <= a or b;
    layer0_outputs(2997) <= not (a or b);
    layer0_outputs(2998) <= not a or b;
    layer0_outputs(2999) <= not b;
    layer0_outputs(3000) <= 1'b0;
    layer0_outputs(3001) <= not b;
    layer0_outputs(3002) <= a and b;
    layer0_outputs(3003) <= b and not a;
    layer0_outputs(3004) <= a and b;
    layer0_outputs(3005) <= not b;
    layer0_outputs(3006) <= a and b;
    layer0_outputs(3007) <= a xor b;
    layer0_outputs(3008) <= a xor b;
    layer0_outputs(3009) <= not (a or b);
    layer0_outputs(3010) <= not (a xor b);
    layer0_outputs(3011) <= a and b;
    layer0_outputs(3012) <= a;
    layer0_outputs(3013) <= not b;
    layer0_outputs(3014) <= not (a xor b);
    layer0_outputs(3015) <= a;
    layer0_outputs(3016) <= not b;
    layer0_outputs(3017) <= b and not a;
    layer0_outputs(3018) <= not (a or b);
    layer0_outputs(3019) <= a;
    layer0_outputs(3020) <= a or b;
    layer0_outputs(3021) <= b;
    layer0_outputs(3022) <= not (a xor b);
    layer0_outputs(3023) <= not (a xor b);
    layer0_outputs(3024) <= 1'b1;
    layer0_outputs(3025) <= a and not b;
    layer0_outputs(3026) <= not (a xor b);
    layer0_outputs(3027) <= b;
    layer0_outputs(3028) <= not b or a;
    layer0_outputs(3029) <= a xor b;
    layer0_outputs(3030) <= not (a xor b);
    layer0_outputs(3031) <= b and not a;
    layer0_outputs(3032) <= a or b;
    layer0_outputs(3033) <= not (a xor b);
    layer0_outputs(3034) <= b and not a;
    layer0_outputs(3035) <= a;
    layer0_outputs(3036) <= b;
    layer0_outputs(3037) <= not (a xor b);
    layer0_outputs(3038) <= a or b;
    layer0_outputs(3039) <= a xor b;
    layer0_outputs(3040) <= b and not a;
    layer0_outputs(3041) <= not a;
    layer0_outputs(3042) <= b;
    layer0_outputs(3043) <= not (a or b);
    layer0_outputs(3044) <= not (a or b);
    layer0_outputs(3045) <= not b or a;
    layer0_outputs(3046) <= a or b;
    layer0_outputs(3047) <= not b;
    layer0_outputs(3048) <= not a;
    layer0_outputs(3049) <= a;
    layer0_outputs(3050) <= 1'b1;
    layer0_outputs(3051) <= a and b;
    layer0_outputs(3052) <= a or b;
    layer0_outputs(3053) <= a;
    layer0_outputs(3054) <= not (a xor b);
    layer0_outputs(3055) <= not (a xor b);
    layer0_outputs(3056) <= not (a or b);
    layer0_outputs(3057) <= a or b;
    layer0_outputs(3058) <= a or b;
    layer0_outputs(3059) <= not b;
    layer0_outputs(3060) <= a xor b;
    layer0_outputs(3061) <= b;
    layer0_outputs(3062) <= a;
    layer0_outputs(3063) <= not (a or b);
    layer0_outputs(3064) <= a or b;
    layer0_outputs(3065) <= a or b;
    layer0_outputs(3066) <= a;
    layer0_outputs(3067) <= a and not b;
    layer0_outputs(3068) <= not (a xor b);
    layer0_outputs(3069) <= b and not a;
    layer0_outputs(3070) <= not a or b;
    layer0_outputs(3071) <= a;
    layer0_outputs(3072) <= not b or a;
    layer0_outputs(3073) <= not a;
    layer0_outputs(3074) <= not b;
    layer0_outputs(3075) <= not a or b;
    layer0_outputs(3076) <= a xor b;
    layer0_outputs(3077) <= not (a or b);
    layer0_outputs(3078) <= not (a xor b);
    layer0_outputs(3079) <= not (a or b);
    layer0_outputs(3080) <= b and not a;
    layer0_outputs(3081) <= not a or b;
    layer0_outputs(3082) <= not (a or b);
    layer0_outputs(3083) <= not b or a;
    layer0_outputs(3084) <= not a or b;
    layer0_outputs(3085) <= b and not a;
    layer0_outputs(3086) <= a xor b;
    layer0_outputs(3087) <= not (a xor b);
    layer0_outputs(3088) <= not a;
    layer0_outputs(3089) <= a;
    layer0_outputs(3090) <= a xor b;
    layer0_outputs(3091) <= a or b;
    layer0_outputs(3092) <= not a or b;
    layer0_outputs(3093) <= a or b;
    layer0_outputs(3094) <= a xor b;
    layer0_outputs(3095) <= a or b;
    layer0_outputs(3096) <= not (a xor b);
    layer0_outputs(3097) <= not b or a;
    layer0_outputs(3098) <= not (a or b);
    layer0_outputs(3099) <= not (a or b);
    layer0_outputs(3100) <= not (a or b);
    layer0_outputs(3101) <= b;
    layer0_outputs(3102) <= a or b;
    layer0_outputs(3103) <= not (a or b);
    layer0_outputs(3104) <= a xor b;
    layer0_outputs(3105) <= not (a xor b);
    layer0_outputs(3106) <= a xor b;
    layer0_outputs(3107) <= a;
    layer0_outputs(3108) <= not (a and b);
    layer0_outputs(3109) <= not a or b;
    layer0_outputs(3110) <= not b;
    layer0_outputs(3111) <= not b;
    layer0_outputs(3112) <= a and not b;
    layer0_outputs(3113) <= not a or b;
    layer0_outputs(3114) <= a xor b;
    layer0_outputs(3115) <= b;
    layer0_outputs(3116) <= b;
    layer0_outputs(3117) <= not (a or b);
    layer0_outputs(3118) <= not a or b;
    layer0_outputs(3119) <= not a;
    layer0_outputs(3120) <= not b or a;
    layer0_outputs(3121) <= a and not b;
    layer0_outputs(3122) <= a or b;
    layer0_outputs(3123) <= not (a xor b);
    layer0_outputs(3124) <= not b or a;
    layer0_outputs(3125) <= a or b;
    layer0_outputs(3126) <= a;
    layer0_outputs(3127) <= not b or a;
    layer0_outputs(3128) <= a;
    layer0_outputs(3129) <= not b or a;
    layer0_outputs(3130) <= a and b;
    layer0_outputs(3131) <= not (a or b);
    layer0_outputs(3132) <= a;
    layer0_outputs(3133) <= not b;
    layer0_outputs(3134) <= 1'b1;
    layer0_outputs(3135) <= b and not a;
    layer0_outputs(3136) <= a xor b;
    layer0_outputs(3137) <= a;
    layer0_outputs(3138) <= not a or b;
    layer0_outputs(3139) <= b and not a;
    layer0_outputs(3140) <= a or b;
    layer0_outputs(3141) <= not (a xor b);
    layer0_outputs(3142) <= b;
    layer0_outputs(3143) <= not a;
    layer0_outputs(3144) <= not b;
    layer0_outputs(3145) <= b;
    layer0_outputs(3146) <= 1'b1;
    layer0_outputs(3147) <= a xor b;
    layer0_outputs(3148) <= not b or a;
    layer0_outputs(3149) <= not (a xor b);
    layer0_outputs(3150) <= a or b;
    layer0_outputs(3151) <= a xor b;
    layer0_outputs(3152) <= not (a or b);
    layer0_outputs(3153) <= not b or a;
    layer0_outputs(3154) <= a xor b;
    layer0_outputs(3155) <= a and b;
    layer0_outputs(3156) <= not (a xor b);
    layer0_outputs(3157) <= not a or b;
    layer0_outputs(3158) <= a xor b;
    layer0_outputs(3159) <= b;
    layer0_outputs(3160) <= a or b;
    layer0_outputs(3161) <= b and not a;
    layer0_outputs(3162) <= b;
    layer0_outputs(3163) <= a;
    layer0_outputs(3164) <= not a;
    layer0_outputs(3165) <= not a;
    layer0_outputs(3166) <= a xor b;
    layer0_outputs(3167) <= not (a or b);
    layer0_outputs(3168) <= not a;
    layer0_outputs(3169) <= not a;
    layer0_outputs(3170) <= not (a xor b);
    layer0_outputs(3171) <= not a;
    layer0_outputs(3172) <= a or b;
    layer0_outputs(3173) <= not (a xor b);
    layer0_outputs(3174) <= not a or b;
    layer0_outputs(3175) <= a or b;
    layer0_outputs(3176) <= b;
    layer0_outputs(3177) <= a xor b;
    layer0_outputs(3178) <= not a or b;
    layer0_outputs(3179) <= not a or b;
    layer0_outputs(3180) <= b;
    layer0_outputs(3181) <= not a or b;
    layer0_outputs(3182) <= b and not a;
    layer0_outputs(3183) <= not b;
    layer0_outputs(3184) <= not (a or b);
    layer0_outputs(3185) <= b;
    layer0_outputs(3186) <= b;
    layer0_outputs(3187) <= not b;
    layer0_outputs(3188) <= a or b;
    layer0_outputs(3189) <= not (a or b);
    layer0_outputs(3190) <= a xor b;
    layer0_outputs(3191) <= a xor b;
    layer0_outputs(3192) <= not (a xor b);
    layer0_outputs(3193) <= a or b;
    layer0_outputs(3194) <= not (a or b);
    layer0_outputs(3195) <= a xor b;
    layer0_outputs(3196) <= a;
    layer0_outputs(3197) <= not b or a;
    layer0_outputs(3198) <= b;
    layer0_outputs(3199) <= not b;
    layer0_outputs(3200) <= a and b;
    layer0_outputs(3201) <= 1'b0;
    layer0_outputs(3202) <= a and not b;
    layer0_outputs(3203) <= not b;
    layer0_outputs(3204) <= a;
    layer0_outputs(3205) <= not a;
    layer0_outputs(3206) <= not a;
    layer0_outputs(3207) <= a or b;
    layer0_outputs(3208) <= not b;
    layer0_outputs(3209) <= not (a or b);
    layer0_outputs(3210) <= a xor b;
    layer0_outputs(3211) <= a xor b;
    layer0_outputs(3212) <= not b or a;
    layer0_outputs(3213) <= a or b;
    layer0_outputs(3214) <= a;
    layer0_outputs(3215) <= not a;
    layer0_outputs(3216) <= a;
    layer0_outputs(3217) <= not (a xor b);
    layer0_outputs(3218) <= a or b;
    layer0_outputs(3219) <= not (a xor b);
    layer0_outputs(3220) <= a or b;
    layer0_outputs(3221) <= a;
    layer0_outputs(3222) <= b;
    layer0_outputs(3223) <= a xor b;
    layer0_outputs(3224) <= a or b;
    layer0_outputs(3225) <= not b or a;
    layer0_outputs(3226) <= a and not b;
    layer0_outputs(3227) <= not b or a;
    layer0_outputs(3228) <= a or b;
    layer0_outputs(3229) <= not b;
    layer0_outputs(3230) <= b and not a;
    layer0_outputs(3231) <= b and not a;
    layer0_outputs(3232) <= a or b;
    layer0_outputs(3233) <= a xor b;
    layer0_outputs(3234) <= not b;
    layer0_outputs(3235) <= not (a xor b);
    layer0_outputs(3236) <= not a;
    layer0_outputs(3237) <= b and not a;
    layer0_outputs(3238) <= a or b;
    layer0_outputs(3239) <= a or b;
    layer0_outputs(3240) <= not (a xor b);
    layer0_outputs(3241) <= not a or b;
    layer0_outputs(3242) <= not a or b;
    layer0_outputs(3243) <= not (a xor b);
    layer0_outputs(3244) <= b;
    layer0_outputs(3245) <= a;
    layer0_outputs(3246) <= a or b;
    layer0_outputs(3247) <= b;
    layer0_outputs(3248) <= not (a or b);
    layer0_outputs(3249) <= a xor b;
    layer0_outputs(3250) <= a;
    layer0_outputs(3251) <= not (a xor b);
    layer0_outputs(3252) <= not (a or b);
    layer0_outputs(3253) <= b;
    layer0_outputs(3254) <= a and not b;
    layer0_outputs(3255) <= a or b;
    layer0_outputs(3256) <= not (a or b);
    layer0_outputs(3257) <= a or b;
    layer0_outputs(3258) <= not (a or b);
    layer0_outputs(3259) <= not (a or b);
    layer0_outputs(3260) <= a and b;
    layer0_outputs(3261) <= a;
    layer0_outputs(3262) <= not a or b;
    layer0_outputs(3263) <= a and not b;
    layer0_outputs(3264) <= a and not b;
    layer0_outputs(3265) <= not b;
    layer0_outputs(3266) <= not (a or b);
    layer0_outputs(3267) <= not b or a;
    layer0_outputs(3268) <= a or b;
    layer0_outputs(3269) <= not (a xor b);
    layer0_outputs(3270) <= a or b;
    layer0_outputs(3271) <= not b or a;
    layer0_outputs(3272) <= a xor b;
    layer0_outputs(3273) <= a or b;
    layer0_outputs(3274) <= a;
    layer0_outputs(3275) <= not (a or b);
    layer0_outputs(3276) <= a or b;
    layer0_outputs(3277) <= a or b;
    layer0_outputs(3278) <= not (a or b);
    layer0_outputs(3279) <= a xor b;
    layer0_outputs(3280) <= a or b;
    layer0_outputs(3281) <= not (a xor b);
    layer0_outputs(3282) <= a or b;
    layer0_outputs(3283) <= not b or a;
    layer0_outputs(3284) <= not b or a;
    layer0_outputs(3285) <= b and not a;
    layer0_outputs(3286) <= a or b;
    layer0_outputs(3287) <= b;
    layer0_outputs(3288) <= a or b;
    layer0_outputs(3289) <= a xor b;
    layer0_outputs(3290) <= a and not b;
    layer0_outputs(3291) <= not (a or b);
    layer0_outputs(3292) <= a or b;
    layer0_outputs(3293) <= not a;
    layer0_outputs(3294) <= not a or b;
    layer0_outputs(3295) <= not (a xor b);
    layer0_outputs(3296) <= a and b;
    layer0_outputs(3297) <= b;
    layer0_outputs(3298) <= a or b;
    layer0_outputs(3299) <= not (a or b);
    layer0_outputs(3300) <= not (a xor b);
    layer0_outputs(3301) <= not (a xor b);
    layer0_outputs(3302) <= not (a and b);
    layer0_outputs(3303) <= a and not b;
    layer0_outputs(3304) <= a xor b;
    layer0_outputs(3305) <= not (a or b);
    layer0_outputs(3306) <= not a or b;
    layer0_outputs(3307) <= not (a xor b);
    layer0_outputs(3308) <= b and not a;
    layer0_outputs(3309) <= not b;
    layer0_outputs(3310) <= a xor b;
    layer0_outputs(3311) <= not (a or b);
    layer0_outputs(3312) <= a or b;
    layer0_outputs(3313) <= b and not a;
    layer0_outputs(3314) <= not (a or b);
    layer0_outputs(3315) <= not a;
    layer0_outputs(3316) <= a xor b;
    layer0_outputs(3317) <= not (a or b);
    layer0_outputs(3318) <= not a or b;
    layer0_outputs(3319) <= b and not a;
    layer0_outputs(3320) <= not (a or b);
    layer0_outputs(3321) <= b;
    layer0_outputs(3322) <= a xor b;
    layer0_outputs(3323) <= not (a xor b);
    layer0_outputs(3324) <= b and not a;
    layer0_outputs(3325) <= not a or b;
    layer0_outputs(3326) <= not (a or b);
    layer0_outputs(3327) <= b;
    layer0_outputs(3328) <= b and not a;
    layer0_outputs(3329) <= b and not a;
    layer0_outputs(3330) <= not (a xor b);
    layer0_outputs(3331) <= not b;
    layer0_outputs(3332) <= b and not a;
    layer0_outputs(3333) <= not b;
    layer0_outputs(3334) <= not a or b;
    layer0_outputs(3335) <= not (a or b);
    layer0_outputs(3336) <= a xor b;
    layer0_outputs(3337) <= not a;
    layer0_outputs(3338) <= not b or a;
    layer0_outputs(3339) <= not a;
    layer0_outputs(3340) <= a and not b;
    layer0_outputs(3341) <= not (a or b);
    layer0_outputs(3342) <= a xor b;
    layer0_outputs(3343) <= not b;
    layer0_outputs(3344) <= not a or b;
    layer0_outputs(3345) <= not b or a;
    layer0_outputs(3346) <= a xor b;
    layer0_outputs(3347) <= not a or b;
    layer0_outputs(3348) <= 1'b0;
    layer0_outputs(3349) <= not (a or b);
    layer0_outputs(3350) <= not a or b;
    layer0_outputs(3351) <= not b;
    layer0_outputs(3352) <= 1'b0;
    layer0_outputs(3353) <= b;
    layer0_outputs(3354) <= not (a and b);
    layer0_outputs(3355) <= b;
    layer0_outputs(3356) <= a and not b;
    layer0_outputs(3357) <= not a or b;
    layer0_outputs(3358) <= not a or b;
    layer0_outputs(3359) <= not b;
    layer0_outputs(3360) <= not (a and b);
    layer0_outputs(3361) <= a xor b;
    layer0_outputs(3362) <= a or b;
    layer0_outputs(3363) <= a xor b;
    layer0_outputs(3364) <= not (a xor b);
    layer0_outputs(3365) <= a and not b;
    layer0_outputs(3366) <= a or b;
    layer0_outputs(3367) <= not a or b;
    layer0_outputs(3368) <= a xor b;
    layer0_outputs(3369) <= b;
    layer0_outputs(3370) <= not (a xor b);
    layer0_outputs(3371) <= not (a xor b);
    layer0_outputs(3372) <= not (a or b);
    layer0_outputs(3373) <= not b;
    layer0_outputs(3374) <= a or b;
    layer0_outputs(3375) <= a or b;
    layer0_outputs(3376) <= a and not b;
    layer0_outputs(3377) <= b and not a;
    layer0_outputs(3378) <= b;
    layer0_outputs(3379) <= not a or b;
    layer0_outputs(3380) <= a;
    layer0_outputs(3381) <= not (a or b);
    layer0_outputs(3382) <= not (a and b);
    layer0_outputs(3383) <= b;
    layer0_outputs(3384) <= not b;
    layer0_outputs(3385) <= not b;
    layer0_outputs(3386) <= a;
    layer0_outputs(3387) <= not b or a;
    layer0_outputs(3388) <= not a or b;
    layer0_outputs(3389) <= a;
    layer0_outputs(3390) <= not (a or b);
    layer0_outputs(3391) <= b;
    layer0_outputs(3392) <= 1'b1;
    layer0_outputs(3393) <= a xor b;
    layer0_outputs(3394) <= a and not b;
    layer0_outputs(3395) <= a;
    layer0_outputs(3396) <= a xor b;
    layer0_outputs(3397) <= a or b;
    layer0_outputs(3398) <= not a or b;
    layer0_outputs(3399) <= not a or b;
    layer0_outputs(3400) <= not b or a;
    layer0_outputs(3401) <= not (a xor b);
    layer0_outputs(3402) <= a and not b;
    layer0_outputs(3403) <= a or b;
    layer0_outputs(3404) <= a or b;
    layer0_outputs(3405) <= b and not a;
    layer0_outputs(3406) <= b;
    layer0_outputs(3407) <= 1'b1;
    layer0_outputs(3408) <= a;
    layer0_outputs(3409) <= a and not b;
    layer0_outputs(3410) <= a and not b;
    layer0_outputs(3411) <= not (a or b);
    layer0_outputs(3412) <= a or b;
    layer0_outputs(3413) <= a xor b;
    layer0_outputs(3414) <= b and not a;
    layer0_outputs(3415) <= not (a or b);
    layer0_outputs(3416) <= b and not a;
    layer0_outputs(3417) <= a or b;
    layer0_outputs(3418) <= not (a or b);
    layer0_outputs(3419) <= a and not b;
    layer0_outputs(3420) <= b and not a;
    layer0_outputs(3421) <= a or b;
    layer0_outputs(3422) <= not (a or b);
    layer0_outputs(3423) <= not a or b;
    layer0_outputs(3424) <= not b;
    layer0_outputs(3425) <= not (a or b);
    layer0_outputs(3426) <= a or b;
    layer0_outputs(3427) <= not b;
    layer0_outputs(3428) <= not b or a;
    layer0_outputs(3429) <= not (a or b);
    layer0_outputs(3430) <= a;
    layer0_outputs(3431) <= not b or a;
    layer0_outputs(3432) <= a and b;
    layer0_outputs(3433) <= not a or b;
    layer0_outputs(3434) <= a xor b;
    layer0_outputs(3435) <= not (a and b);
    layer0_outputs(3436) <= a or b;
    layer0_outputs(3437) <= not (a xor b);
    layer0_outputs(3438) <= b and not a;
    layer0_outputs(3439) <= not b or a;
    layer0_outputs(3440) <= a or b;
    layer0_outputs(3441) <= not (a and b);
    layer0_outputs(3442) <= a or b;
    layer0_outputs(3443) <= not (a or b);
    layer0_outputs(3444) <= b and not a;
    layer0_outputs(3445) <= a or b;
    layer0_outputs(3446) <= not b or a;
    layer0_outputs(3447) <= a or b;
    layer0_outputs(3448) <= a xor b;
    layer0_outputs(3449) <= not a or b;
    layer0_outputs(3450) <= not (a xor b);
    layer0_outputs(3451) <= not b;
    layer0_outputs(3452) <= a;
    layer0_outputs(3453) <= not b;
    layer0_outputs(3454) <= not a;
    layer0_outputs(3455) <= a or b;
    layer0_outputs(3456) <= a or b;
    layer0_outputs(3457) <= b;
    layer0_outputs(3458) <= not b or a;
    layer0_outputs(3459) <= not a;
    layer0_outputs(3460) <= a xor b;
    layer0_outputs(3461) <= not b or a;
    layer0_outputs(3462) <= a or b;
    layer0_outputs(3463) <= not (a or b);
    layer0_outputs(3464) <= a xor b;
    layer0_outputs(3465) <= b;
    layer0_outputs(3466) <= a and not b;
    layer0_outputs(3467) <= not (a and b);
    layer0_outputs(3468) <= b and not a;
    layer0_outputs(3469) <= a or b;
    layer0_outputs(3470) <= not (a xor b);
    layer0_outputs(3471) <= b and not a;
    layer0_outputs(3472) <= not a;
    layer0_outputs(3473) <= a;
    layer0_outputs(3474) <= b;
    layer0_outputs(3475) <= not (a or b);
    layer0_outputs(3476) <= not (a xor b);
    layer0_outputs(3477) <= not a;
    layer0_outputs(3478) <= not (a xor b);
    layer0_outputs(3479) <= not (a xor b);
    layer0_outputs(3480) <= a or b;
    layer0_outputs(3481) <= b and not a;
    layer0_outputs(3482) <= 1'b1;
    layer0_outputs(3483) <= b and not a;
    layer0_outputs(3484) <= a or b;
    layer0_outputs(3485) <= not (a or b);
    layer0_outputs(3486) <= a or b;
    layer0_outputs(3487) <= 1'b0;
    layer0_outputs(3488) <= b and not a;
    layer0_outputs(3489) <= b and not a;
    layer0_outputs(3490) <= b and not a;
    layer0_outputs(3491) <= a xor b;
    layer0_outputs(3492) <= not b;
    layer0_outputs(3493) <= not (a or b);
    layer0_outputs(3494) <= not (a or b);
    layer0_outputs(3495) <= not a;
    layer0_outputs(3496) <= not a;
    layer0_outputs(3497) <= not a or b;
    layer0_outputs(3498) <= not a;
    layer0_outputs(3499) <= not b or a;
    layer0_outputs(3500) <= not a;
    layer0_outputs(3501) <= a or b;
    layer0_outputs(3502) <= not (a xor b);
    layer0_outputs(3503) <= a or b;
    layer0_outputs(3504) <= a and not b;
    layer0_outputs(3505) <= b;
    layer0_outputs(3506) <= a;
    layer0_outputs(3507) <= a xor b;
    layer0_outputs(3508) <= not (a or b);
    layer0_outputs(3509) <= not (a or b);
    layer0_outputs(3510) <= b and not a;
    layer0_outputs(3511) <= not (a or b);
    layer0_outputs(3512) <= a or b;
    layer0_outputs(3513) <= not (a or b);
    layer0_outputs(3514) <= not (a xor b);
    layer0_outputs(3515) <= a xor b;
    layer0_outputs(3516) <= not (a or b);
    layer0_outputs(3517) <= b;
    layer0_outputs(3518) <= not (a or b);
    layer0_outputs(3519) <= not (a or b);
    layer0_outputs(3520) <= not a;
    layer0_outputs(3521) <= a or b;
    layer0_outputs(3522) <= not a;
    layer0_outputs(3523) <= a xor b;
    layer0_outputs(3524) <= not (a xor b);
    layer0_outputs(3525) <= a and not b;
    layer0_outputs(3526) <= not b or a;
    layer0_outputs(3527) <= b;
    layer0_outputs(3528) <= a xor b;
    layer0_outputs(3529) <= not b or a;
    layer0_outputs(3530) <= a xor b;
    layer0_outputs(3531) <= not (a or b);
    layer0_outputs(3532) <= a;
    layer0_outputs(3533) <= a or b;
    layer0_outputs(3534) <= a or b;
    layer0_outputs(3535) <= not a;
    layer0_outputs(3536) <= not (a xor b);
    layer0_outputs(3537) <= a xor b;
    layer0_outputs(3538) <= b and not a;
    layer0_outputs(3539) <= a and not b;
    layer0_outputs(3540) <= not b;
    layer0_outputs(3541) <= a and b;
    layer0_outputs(3542) <= a xor b;
    layer0_outputs(3543) <= not b or a;
    layer0_outputs(3544) <= a or b;
    layer0_outputs(3545) <= not b or a;
    layer0_outputs(3546) <= not (a or b);
    layer0_outputs(3547) <= not (a and b);
    layer0_outputs(3548) <= not (a or b);
    layer0_outputs(3549) <= not (a or b);
    layer0_outputs(3550) <= not (a and b);
    layer0_outputs(3551) <= b and not a;
    layer0_outputs(3552) <= 1'b1;
    layer0_outputs(3553) <= a xor b;
    layer0_outputs(3554) <= not a;
    layer0_outputs(3555) <= a;
    layer0_outputs(3556) <= not b or a;
    layer0_outputs(3557) <= not a;
    layer0_outputs(3558) <= a xor b;
    layer0_outputs(3559) <= not b or a;
    layer0_outputs(3560) <= a or b;
    layer0_outputs(3561) <= not a;
    layer0_outputs(3562) <= a and not b;
    layer0_outputs(3563) <= not b or a;
    layer0_outputs(3564) <= a xor b;
    layer0_outputs(3565) <= b and not a;
    layer0_outputs(3566) <= a;
    layer0_outputs(3567) <= not (a or b);
    layer0_outputs(3568) <= not b;
    layer0_outputs(3569) <= a;
    layer0_outputs(3570) <= a or b;
    layer0_outputs(3571) <= a or b;
    layer0_outputs(3572) <= b and not a;
    layer0_outputs(3573) <= not a;
    layer0_outputs(3574) <= a or b;
    layer0_outputs(3575) <= not a or b;
    layer0_outputs(3576) <= a xor b;
    layer0_outputs(3577) <= a xor b;
    layer0_outputs(3578) <= a and not b;
    layer0_outputs(3579) <= b and not a;
    layer0_outputs(3580) <= a and not b;
    layer0_outputs(3581) <= not (a or b);
    layer0_outputs(3582) <= not a or b;
    layer0_outputs(3583) <= a xor b;
    layer0_outputs(3584) <= a or b;
    layer0_outputs(3585) <= not a;
    layer0_outputs(3586) <= not (a xor b);
    layer0_outputs(3587) <= b and not a;
    layer0_outputs(3588) <= a or b;
    layer0_outputs(3589) <= not a;
    layer0_outputs(3590) <= a and b;
    layer0_outputs(3591) <= b and not a;
    layer0_outputs(3592) <= not a or b;
    layer0_outputs(3593) <= not (a or b);
    layer0_outputs(3594) <= a xor b;
    layer0_outputs(3595) <= a or b;
    layer0_outputs(3596) <= a and b;
    layer0_outputs(3597) <= b;
    layer0_outputs(3598) <= not b;
    layer0_outputs(3599) <= not a or b;
    layer0_outputs(3600) <= not (a xor b);
    layer0_outputs(3601) <= not (a or b);
    layer0_outputs(3602) <= a and b;
    layer0_outputs(3603) <= not a or b;
    layer0_outputs(3604) <= b;
    layer0_outputs(3605) <= a xor b;
    layer0_outputs(3606) <= not a or b;
    layer0_outputs(3607) <= a or b;
    layer0_outputs(3608) <= not (a or b);
    layer0_outputs(3609) <= not b or a;
    layer0_outputs(3610) <= not a or b;
    layer0_outputs(3611) <= not b;
    layer0_outputs(3612) <= not b;
    layer0_outputs(3613) <= a and b;
    layer0_outputs(3614) <= not (a or b);
    layer0_outputs(3615) <= a or b;
    layer0_outputs(3616) <= a;
    layer0_outputs(3617) <= a xor b;
    layer0_outputs(3618) <= a xor b;
    layer0_outputs(3619) <= a or b;
    layer0_outputs(3620) <= not (a xor b);
    layer0_outputs(3621) <= not (a or b);
    layer0_outputs(3622) <= not (a and b);
    layer0_outputs(3623) <= b;
    layer0_outputs(3624) <= b and not a;
    layer0_outputs(3625) <= not b or a;
    layer0_outputs(3626) <= not a or b;
    layer0_outputs(3627) <= a;
    layer0_outputs(3628) <= a and not b;
    layer0_outputs(3629) <= a;
    layer0_outputs(3630) <= a and not b;
    layer0_outputs(3631) <= a xor b;
    layer0_outputs(3632) <= a or b;
    layer0_outputs(3633) <= not (a or b);
    layer0_outputs(3634) <= 1'b0;
    layer0_outputs(3635) <= not (a or b);
    layer0_outputs(3636) <= b and not a;
    layer0_outputs(3637) <= a or b;
    layer0_outputs(3638) <= b and not a;
    layer0_outputs(3639) <= b;
    layer0_outputs(3640) <= a and not b;
    layer0_outputs(3641) <= not a or b;
    layer0_outputs(3642) <= not b;
    layer0_outputs(3643) <= a or b;
    layer0_outputs(3644) <= not (a or b);
    layer0_outputs(3645) <= not a or b;
    layer0_outputs(3646) <= a or b;
    layer0_outputs(3647) <= a or b;
    layer0_outputs(3648) <= not (a or b);
    layer0_outputs(3649) <= not (a xor b);
    layer0_outputs(3650) <= a xor b;
    layer0_outputs(3651) <= a and b;
    layer0_outputs(3652) <= b;
    layer0_outputs(3653) <= b;
    layer0_outputs(3654) <= not a or b;
    layer0_outputs(3655) <= a or b;
    layer0_outputs(3656) <= not a;
    layer0_outputs(3657) <= a or b;
    layer0_outputs(3658) <= not (a xor b);
    layer0_outputs(3659) <= not (a and b);
    layer0_outputs(3660) <= not b;
    layer0_outputs(3661) <= a and not b;
    layer0_outputs(3662) <= not (a or b);
    layer0_outputs(3663) <= not (a xor b);
    layer0_outputs(3664) <= not b or a;
    layer0_outputs(3665) <= not b;
    layer0_outputs(3666) <= b;
    layer0_outputs(3667) <= a or b;
    layer0_outputs(3668) <= not (a or b);
    layer0_outputs(3669) <= not (a xor b);
    layer0_outputs(3670) <= b and not a;
    layer0_outputs(3671) <= a and not b;
    layer0_outputs(3672) <= a or b;
    layer0_outputs(3673) <= b and not a;
    layer0_outputs(3674) <= not (a or b);
    layer0_outputs(3675) <= a and b;
    layer0_outputs(3676) <= a xor b;
    layer0_outputs(3677) <= b and not a;
    layer0_outputs(3678) <= a or b;
    layer0_outputs(3679) <= not a or b;
    layer0_outputs(3680) <= not (a or b);
    layer0_outputs(3681) <= a xor b;
    layer0_outputs(3682) <= a or b;
    layer0_outputs(3683) <= not a;
    layer0_outputs(3684) <= a and not b;
    layer0_outputs(3685) <= a;
    layer0_outputs(3686) <= b;
    layer0_outputs(3687) <= not b;
    layer0_outputs(3688) <= a or b;
    layer0_outputs(3689) <= b and not a;
    layer0_outputs(3690) <= b;
    layer0_outputs(3691) <= not (a or b);
    layer0_outputs(3692) <= not b or a;
    layer0_outputs(3693) <= not a or b;
    layer0_outputs(3694) <= 1'b0;
    layer0_outputs(3695) <= b and not a;
    layer0_outputs(3696) <= a and not b;
    layer0_outputs(3697) <= b and not a;
    layer0_outputs(3698) <= a or b;
    layer0_outputs(3699) <= a and not b;
    layer0_outputs(3700) <= not b;
    layer0_outputs(3701) <= not a or b;
    layer0_outputs(3702) <= a and b;
    layer0_outputs(3703) <= not (a or b);
    layer0_outputs(3704) <= not a;
    layer0_outputs(3705) <= a;
    layer0_outputs(3706) <= a or b;
    layer0_outputs(3707) <= not (a xor b);
    layer0_outputs(3708) <= not a;
    layer0_outputs(3709) <= a xor b;
    layer0_outputs(3710) <= a or b;
    layer0_outputs(3711) <= not (a xor b);
    layer0_outputs(3712) <= not (a or b);
    layer0_outputs(3713) <= a xor b;
    layer0_outputs(3714) <= not (a or b);
    layer0_outputs(3715) <= a or b;
    layer0_outputs(3716) <= a xor b;
    layer0_outputs(3717) <= not (a and b);
    layer0_outputs(3718) <= not (a xor b);
    layer0_outputs(3719) <= a xor b;
    layer0_outputs(3720) <= a xor b;
    layer0_outputs(3721) <= not (a xor b);
    layer0_outputs(3722) <= not a or b;
    layer0_outputs(3723) <= a and not b;
    layer0_outputs(3724) <= a or b;
    layer0_outputs(3725) <= not (a xor b);
    layer0_outputs(3726) <= not (a or b);
    layer0_outputs(3727) <= a xor b;
    layer0_outputs(3728) <= a xor b;
    layer0_outputs(3729) <= not (a or b);
    layer0_outputs(3730) <= b;
    layer0_outputs(3731) <= not (a or b);
    layer0_outputs(3732) <= not a or b;
    layer0_outputs(3733) <= a and not b;
    layer0_outputs(3734) <= b and not a;
    layer0_outputs(3735) <= a;
    layer0_outputs(3736) <= a xor b;
    layer0_outputs(3737) <= a and b;
    layer0_outputs(3738) <= a or b;
    layer0_outputs(3739) <= a or b;
    layer0_outputs(3740) <= not b or a;
    layer0_outputs(3741) <= not (a or b);
    layer0_outputs(3742) <= a and b;
    layer0_outputs(3743) <= not (a xor b);
    layer0_outputs(3744) <= a or b;
    layer0_outputs(3745) <= b;
    layer0_outputs(3746) <= not (a or b);
    layer0_outputs(3747) <= b and not a;
    layer0_outputs(3748) <= a or b;
    layer0_outputs(3749) <= not (a or b);
    layer0_outputs(3750) <= not (a xor b);
    layer0_outputs(3751) <= a or b;
    layer0_outputs(3752) <= a xor b;
    layer0_outputs(3753) <= 1'b1;
    layer0_outputs(3754) <= b;
    layer0_outputs(3755) <= not (a xor b);
    layer0_outputs(3756) <= not b;
    layer0_outputs(3757) <= a or b;
    layer0_outputs(3758) <= a and not b;
    layer0_outputs(3759) <= a xor b;
    layer0_outputs(3760) <= a xor b;
    layer0_outputs(3761) <= not (a or b);
    layer0_outputs(3762) <= 1'b0;
    layer0_outputs(3763) <= not b or a;
    layer0_outputs(3764) <= not b;
    layer0_outputs(3765) <= a;
    layer0_outputs(3766) <= not b;
    layer0_outputs(3767) <= a or b;
    layer0_outputs(3768) <= a or b;
    layer0_outputs(3769) <= not (a or b);
    layer0_outputs(3770) <= a;
    layer0_outputs(3771) <= not (a or b);
    layer0_outputs(3772) <= not b;
    layer0_outputs(3773) <= 1'b1;
    layer0_outputs(3774) <= not (a xor b);
    layer0_outputs(3775) <= a or b;
    layer0_outputs(3776) <= not b;
    layer0_outputs(3777) <= a;
    layer0_outputs(3778) <= not (a or b);
    layer0_outputs(3779) <= b and not a;
    layer0_outputs(3780) <= a or b;
    layer0_outputs(3781) <= a;
    layer0_outputs(3782) <= a or b;
    layer0_outputs(3783) <= not (a or b);
    layer0_outputs(3784) <= not (a xor b);
    layer0_outputs(3785) <= not b;
    layer0_outputs(3786) <= a or b;
    layer0_outputs(3787) <= b and not a;
    layer0_outputs(3788) <= a and not b;
    layer0_outputs(3789) <= not a or b;
    layer0_outputs(3790) <= not (a xor b);
    layer0_outputs(3791) <= a;
    layer0_outputs(3792) <= not a;
    layer0_outputs(3793) <= b;
    layer0_outputs(3794) <= not b;
    layer0_outputs(3795) <= not (a xor b);
    layer0_outputs(3796) <= a and not b;
    layer0_outputs(3797) <= not a;
    layer0_outputs(3798) <= not (a xor b);
    layer0_outputs(3799) <= not (a or b);
    layer0_outputs(3800) <= a or b;
    layer0_outputs(3801) <= a or b;
    layer0_outputs(3802) <= not (a xor b);
    layer0_outputs(3803) <= not a or b;
    layer0_outputs(3804) <= not a;
    layer0_outputs(3805) <= a xor b;
    layer0_outputs(3806) <= not a;
    layer0_outputs(3807) <= a xor b;
    layer0_outputs(3808) <= not a or b;
    layer0_outputs(3809) <= a or b;
    layer0_outputs(3810) <= a xor b;
    layer0_outputs(3811) <= not a;
    layer0_outputs(3812) <= a and not b;
    layer0_outputs(3813) <= not (a or b);
    layer0_outputs(3814) <= not b or a;
    layer0_outputs(3815) <= a xor b;
    layer0_outputs(3816) <= not b or a;
    layer0_outputs(3817) <= not (a or b);
    layer0_outputs(3818) <= not b;
    layer0_outputs(3819) <= not a;
    layer0_outputs(3820) <= a or b;
    layer0_outputs(3821) <= not a;
    layer0_outputs(3822) <= not b or a;
    layer0_outputs(3823) <= not (a xor b);
    layer0_outputs(3824) <= not (a or b);
    layer0_outputs(3825) <= not (a or b);
    layer0_outputs(3826) <= not a;
    layer0_outputs(3827) <= not (a or b);
    layer0_outputs(3828) <= not b;
    layer0_outputs(3829) <= a or b;
    layer0_outputs(3830) <= a;
    layer0_outputs(3831) <= not (a or b);
    layer0_outputs(3832) <= a and b;
    layer0_outputs(3833) <= a and not b;
    layer0_outputs(3834) <= not (a or b);
    layer0_outputs(3835) <= a or b;
    layer0_outputs(3836) <= a and b;
    layer0_outputs(3837) <= not a;
    layer0_outputs(3838) <= not (a xor b);
    layer0_outputs(3839) <= not (a or b);
    layer0_outputs(3840) <= not (a xor b);
    layer0_outputs(3841) <= 1'b0;
    layer0_outputs(3842) <= a;
    layer0_outputs(3843) <= a xor b;
    layer0_outputs(3844) <= not (a and b);
    layer0_outputs(3845) <= not (a xor b);
    layer0_outputs(3846) <= not (a or b);
    layer0_outputs(3847) <= a or b;
    layer0_outputs(3848) <= a and not b;
    layer0_outputs(3849) <= not b;
    layer0_outputs(3850) <= not a;
    layer0_outputs(3851) <= not a or b;
    layer0_outputs(3852) <= not (a or b);
    layer0_outputs(3853) <= not (a or b);
    layer0_outputs(3854) <= not (a or b);
    layer0_outputs(3855) <= not (a xor b);
    layer0_outputs(3856) <= not (a xor b);
    layer0_outputs(3857) <= not b or a;
    layer0_outputs(3858) <= a or b;
    layer0_outputs(3859) <= not b or a;
    layer0_outputs(3860) <= a;
    layer0_outputs(3861) <= not b;
    layer0_outputs(3862) <= a or b;
    layer0_outputs(3863) <= not b;
    layer0_outputs(3864) <= a xor b;
    layer0_outputs(3865) <= not (a or b);
    layer0_outputs(3866) <= a or b;
    layer0_outputs(3867) <= a or b;
    layer0_outputs(3868) <= not b;
    layer0_outputs(3869) <= a or b;
    layer0_outputs(3870) <= a xor b;
    layer0_outputs(3871) <= not b or a;
    layer0_outputs(3872) <= not (a and b);
    layer0_outputs(3873) <= not a;
    layer0_outputs(3874) <= not (a or b);
    layer0_outputs(3875) <= a or b;
    layer0_outputs(3876) <= not (a or b);
    layer0_outputs(3877) <= a xor b;
    layer0_outputs(3878) <= not (a or b);
    layer0_outputs(3879) <= 1'b0;
    layer0_outputs(3880) <= b;
    layer0_outputs(3881) <= a and not b;
    layer0_outputs(3882) <= not (a or b);
    layer0_outputs(3883) <= b and not a;
    layer0_outputs(3884) <= not a;
    layer0_outputs(3885) <= a or b;
    layer0_outputs(3886) <= not a;
    layer0_outputs(3887) <= b and not a;
    layer0_outputs(3888) <= not (a xor b);
    layer0_outputs(3889) <= not (a xor b);
    layer0_outputs(3890) <= a and not b;
    layer0_outputs(3891) <= not (a xor b);
    layer0_outputs(3892) <= not a or b;
    layer0_outputs(3893) <= a and b;
    layer0_outputs(3894) <= not (a or b);
    layer0_outputs(3895) <= not b or a;
    layer0_outputs(3896) <= b and not a;
    layer0_outputs(3897) <= a or b;
    layer0_outputs(3898) <= a and b;
    layer0_outputs(3899) <= a;
    layer0_outputs(3900) <= a xor b;
    layer0_outputs(3901) <= not b;
    layer0_outputs(3902) <= a xor b;
    layer0_outputs(3903) <= not (a and b);
    layer0_outputs(3904) <= b and not a;
    layer0_outputs(3905) <= not (a or b);
    layer0_outputs(3906) <= not (a or b);
    layer0_outputs(3907) <= a and not b;
    layer0_outputs(3908) <= a or b;
    layer0_outputs(3909) <= not b;
    layer0_outputs(3910) <= not a;
    layer0_outputs(3911) <= 1'b0;
    layer0_outputs(3912) <= b and not a;
    layer0_outputs(3913) <= b and not a;
    layer0_outputs(3914) <= not (a and b);
    layer0_outputs(3915) <= a;
    layer0_outputs(3916) <= not a or b;
    layer0_outputs(3917) <= not (a xor b);
    layer0_outputs(3918) <= a or b;
    layer0_outputs(3919) <= a or b;
    layer0_outputs(3920) <= not (a or b);
    layer0_outputs(3921) <= 1'b0;
    layer0_outputs(3922) <= b;
    layer0_outputs(3923) <= b;
    layer0_outputs(3924) <= not (a or b);
    layer0_outputs(3925) <= not a;
    layer0_outputs(3926) <= not (a xor b);
    layer0_outputs(3927) <= not (a or b);
    layer0_outputs(3928) <= a xor b;
    layer0_outputs(3929) <= a or b;
    layer0_outputs(3930) <= not (a or b);
    layer0_outputs(3931) <= a and not b;
    layer0_outputs(3932) <= a or b;
    layer0_outputs(3933) <= not (a or b);
    layer0_outputs(3934) <= b and not a;
    layer0_outputs(3935) <= not a;
    layer0_outputs(3936) <= not (a or b);
    layer0_outputs(3937) <= a xor b;
    layer0_outputs(3938) <= not (a xor b);
    layer0_outputs(3939) <= not (a and b);
    layer0_outputs(3940) <= not b or a;
    layer0_outputs(3941) <= not (a or b);
    layer0_outputs(3942) <= b and not a;
    layer0_outputs(3943) <= not a;
    layer0_outputs(3944) <= not (a xor b);
    layer0_outputs(3945) <= a and b;
    layer0_outputs(3946) <= not a or b;
    layer0_outputs(3947) <= not b;
    layer0_outputs(3948) <= not (a or b);
    layer0_outputs(3949) <= not (a and b);
    layer0_outputs(3950) <= a xor b;
    layer0_outputs(3951) <= a and not b;
    layer0_outputs(3952) <= a;
    layer0_outputs(3953) <= a xor b;
    layer0_outputs(3954) <= a;
    layer0_outputs(3955) <= not (a xor b);
    layer0_outputs(3956) <= not (a or b);
    layer0_outputs(3957) <= not (a or b);
    layer0_outputs(3958) <= not a or b;
    layer0_outputs(3959) <= not (a or b);
    layer0_outputs(3960) <= a or b;
    layer0_outputs(3961) <= not (a or b);
    layer0_outputs(3962) <= a or b;
    layer0_outputs(3963) <= not (a or b);
    layer0_outputs(3964) <= a or b;
    layer0_outputs(3965) <= b and not a;
    layer0_outputs(3966) <= not a or b;
    layer0_outputs(3967) <= a or b;
    layer0_outputs(3968) <= not b;
    layer0_outputs(3969) <= not (a or b);
    layer0_outputs(3970) <= a;
    layer0_outputs(3971) <= not (a or b);
    layer0_outputs(3972) <= not (a or b);
    layer0_outputs(3973) <= not a or b;
    layer0_outputs(3974) <= b;
    layer0_outputs(3975) <= a or b;
    layer0_outputs(3976) <= not b or a;
    layer0_outputs(3977) <= not a or b;
    layer0_outputs(3978) <= not b or a;
    layer0_outputs(3979) <= a and b;
    layer0_outputs(3980) <= a and b;
    layer0_outputs(3981) <= not b;
    layer0_outputs(3982) <= not (a or b);
    layer0_outputs(3983) <= not a;
    layer0_outputs(3984) <= a;
    layer0_outputs(3985) <= not (a xor b);
    layer0_outputs(3986) <= not a or b;
    layer0_outputs(3987) <= a xor b;
    layer0_outputs(3988) <= b;
    layer0_outputs(3989) <= not a;
    layer0_outputs(3990) <= a and b;
    layer0_outputs(3991) <= not a or b;
    layer0_outputs(3992) <= not (a xor b);
    layer0_outputs(3993) <= a and not b;
    layer0_outputs(3994) <= a or b;
    layer0_outputs(3995) <= b and not a;
    layer0_outputs(3996) <= not (a xor b);
    layer0_outputs(3997) <= not (a or b);
    layer0_outputs(3998) <= a and b;
    layer0_outputs(3999) <= a or b;
    layer0_outputs(4000) <= b and not a;
    layer0_outputs(4001) <= b;
    layer0_outputs(4002) <= not (a or b);
    layer0_outputs(4003) <= a xor b;
    layer0_outputs(4004) <= b;
    layer0_outputs(4005) <= a or b;
    layer0_outputs(4006) <= a or b;
    layer0_outputs(4007) <= not (a or b);
    layer0_outputs(4008) <= not (a xor b);
    layer0_outputs(4009) <= not b or a;
    layer0_outputs(4010) <= not (a or b);
    layer0_outputs(4011) <= b and not a;
    layer0_outputs(4012) <= a and not b;
    layer0_outputs(4013) <= a or b;
    layer0_outputs(4014) <= a xor b;
    layer0_outputs(4015) <= b;
    layer0_outputs(4016) <= not (a or b);
    layer0_outputs(4017) <= not a or b;
    layer0_outputs(4018) <= a or b;
    layer0_outputs(4019) <= not (a xor b);
    layer0_outputs(4020) <= a;
    layer0_outputs(4021) <= a and b;
    layer0_outputs(4022) <= not b;
    layer0_outputs(4023) <= a;
    layer0_outputs(4024) <= not a;
    layer0_outputs(4025) <= b and not a;
    layer0_outputs(4026) <= not (a or b);
    layer0_outputs(4027) <= a and not b;
    layer0_outputs(4028) <= not (a xor b);
    layer0_outputs(4029) <= not (a xor b);
    layer0_outputs(4030) <= a and not b;
    layer0_outputs(4031) <= a;
    layer0_outputs(4032) <= b and not a;
    layer0_outputs(4033) <= a xor b;
    layer0_outputs(4034) <= b;
    layer0_outputs(4035) <= a and not b;
    layer0_outputs(4036) <= not (a xor b);
    layer0_outputs(4037) <= b and not a;
    layer0_outputs(4038) <= a xor b;
    layer0_outputs(4039) <= b;
    layer0_outputs(4040) <= b;
    layer0_outputs(4041) <= b;
    layer0_outputs(4042) <= a and b;
    layer0_outputs(4043) <= a and not b;
    layer0_outputs(4044) <= not (a or b);
    layer0_outputs(4045) <= a xor b;
    layer0_outputs(4046) <= not b;
    layer0_outputs(4047) <= a and not b;
    layer0_outputs(4048) <= not (a or b);
    layer0_outputs(4049) <= not a or b;
    layer0_outputs(4050) <= a and not b;
    layer0_outputs(4051) <= not (a or b);
    layer0_outputs(4052) <= not (a xor b);
    layer0_outputs(4053) <= a and not b;
    layer0_outputs(4054) <= not b;
    layer0_outputs(4055) <= a and b;
    layer0_outputs(4056) <= a;
    layer0_outputs(4057) <= not (a xor b);
    layer0_outputs(4058) <= b and not a;
    layer0_outputs(4059) <= not b;
    layer0_outputs(4060) <= not b or a;
    layer0_outputs(4061) <= not (a or b);
    layer0_outputs(4062) <= a or b;
    layer0_outputs(4063) <= not a or b;
    layer0_outputs(4064) <= not b or a;
    layer0_outputs(4065) <= a and not b;
    layer0_outputs(4066) <= a and b;
    layer0_outputs(4067) <= not b;
    layer0_outputs(4068) <= a xor b;
    layer0_outputs(4069) <= a xor b;
    layer0_outputs(4070) <= a xor b;
    layer0_outputs(4071) <= a xor b;
    layer0_outputs(4072) <= not b or a;
    layer0_outputs(4073) <= a or b;
    layer0_outputs(4074) <= a xor b;
    layer0_outputs(4075) <= not b;
    layer0_outputs(4076) <= not (a or b);
    layer0_outputs(4077) <= not b;
    layer0_outputs(4078) <= a and b;
    layer0_outputs(4079) <= b and not a;
    layer0_outputs(4080) <= not (a or b);
    layer0_outputs(4081) <= not b;
    layer0_outputs(4082) <= a xor b;
    layer0_outputs(4083) <= a xor b;
    layer0_outputs(4084) <= not a or b;
    layer0_outputs(4085) <= a or b;
    layer0_outputs(4086) <= not (a xor b);
    layer0_outputs(4087) <= not (a or b);
    layer0_outputs(4088) <= not (a or b);
    layer0_outputs(4089) <= not b or a;
    layer0_outputs(4090) <= not a;
    layer0_outputs(4091) <= 1'b0;
    layer0_outputs(4092) <= not b or a;
    layer0_outputs(4093) <= a and b;
    layer0_outputs(4094) <= a xor b;
    layer0_outputs(4095) <= a or b;
    layer0_outputs(4096) <= not (a xor b);
    layer0_outputs(4097) <= a;
    layer0_outputs(4098) <= not a;
    layer0_outputs(4099) <= not (a xor b);
    layer0_outputs(4100) <= b;
    layer0_outputs(4101) <= 1'b0;
    layer0_outputs(4102) <= not (a xor b);
    layer0_outputs(4103) <= a and not b;
    layer0_outputs(4104) <= not b;
    layer0_outputs(4105) <= a or b;
    layer0_outputs(4106) <= not b or a;
    layer0_outputs(4107) <= a or b;
    layer0_outputs(4108) <= not a or b;
    layer0_outputs(4109) <= a xor b;
    layer0_outputs(4110) <= b;
    layer0_outputs(4111) <= not (a or b);
    layer0_outputs(4112) <= a or b;
    layer0_outputs(4113) <= not (a xor b);
    layer0_outputs(4114) <= a xor b;
    layer0_outputs(4115) <= a and not b;
    layer0_outputs(4116) <= a xor b;
    layer0_outputs(4117) <= a or b;
    layer0_outputs(4118) <= not b;
    layer0_outputs(4119) <= a or b;
    layer0_outputs(4120) <= a and b;
    layer0_outputs(4121) <= not b or a;
    layer0_outputs(4122) <= not a or b;
    layer0_outputs(4123) <= a or b;
    layer0_outputs(4124) <= not b;
    layer0_outputs(4125) <= not b;
    layer0_outputs(4126) <= not (a or b);
    layer0_outputs(4127) <= a and not b;
    layer0_outputs(4128) <= a xor b;
    layer0_outputs(4129) <= not (a or b);
    layer0_outputs(4130) <= not a;
    layer0_outputs(4131) <= not (a xor b);
    layer0_outputs(4132) <= not b;
    layer0_outputs(4133) <= not b;
    layer0_outputs(4134) <= a or b;
    layer0_outputs(4135) <= a and not b;
    layer0_outputs(4136) <= a and b;
    layer0_outputs(4137) <= a;
    layer0_outputs(4138) <= not b;
    layer0_outputs(4139) <= a xor b;
    layer0_outputs(4140) <= not b or a;
    layer0_outputs(4141) <= not b;
    layer0_outputs(4142) <= not (a xor b);
    layer0_outputs(4143) <= not (a or b);
    layer0_outputs(4144) <= not (a or b);
    layer0_outputs(4145) <= a xor b;
    layer0_outputs(4146) <= b;
    layer0_outputs(4147) <= a xor b;
    layer0_outputs(4148) <= not a;
    layer0_outputs(4149) <= a xor b;
    layer0_outputs(4150) <= not (a xor b);
    layer0_outputs(4151) <= not (a or b);
    layer0_outputs(4152) <= a or b;
    layer0_outputs(4153) <= a and b;
    layer0_outputs(4154) <= not (a or b);
    layer0_outputs(4155) <= b and not a;
    layer0_outputs(4156) <= a or b;
    layer0_outputs(4157) <= not a or b;
    layer0_outputs(4158) <= not (a xor b);
    layer0_outputs(4159) <= a xor b;
    layer0_outputs(4160) <= not (a or b);
    layer0_outputs(4161) <= a and not b;
    layer0_outputs(4162) <= 1'b1;
    layer0_outputs(4163) <= not a;
    layer0_outputs(4164) <= not a;
    layer0_outputs(4165) <= a xor b;
    layer0_outputs(4166) <= not (a or b);
    layer0_outputs(4167) <= a and b;
    layer0_outputs(4168) <= a xor b;
    layer0_outputs(4169) <= a and not b;
    layer0_outputs(4170) <= a or b;
    layer0_outputs(4171) <= a and b;
    layer0_outputs(4172) <= a;
    layer0_outputs(4173) <= a;
    layer0_outputs(4174) <= not (a or b);
    layer0_outputs(4175) <= a or b;
    layer0_outputs(4176) <= a and b;
    layer0_outputs(4177) <= not (a or b);
    layer0_outputs(4178) <= not (a or b);
    layer0_outputs(4179) <= not a;
    layer0_outputs(4180) <= not (a or b);
    layer0_outputs(4181) <= a or b;
    layer0_outputs(4182) <= not (a or b);
    layer0_outputs(4183) <= not b;
    layer0_outputs(4184) <= a xor b;
    layer0_outputs(4185) <= a and not b;
    layer0_outputs(4186) <= a or b;
    layer0_outputs(4187) <= not (a xor b);
    layer0_outputs(4188) <= 1'b1;
    layer0_outputs(4189) <= a or b;
    layer0_outputs(4190) <= not (a or b);
    layer0_outputs(4191) <= a xor b;
    layer0_outputs(4192) <= a xor b;
    layer0_outputs(4193) <= not b or a;
    layer0_outputs(4194) <= not (a or b);
    layer0_outputs(4195) <= a;
    layer0_outputs(4196) <= a or b;
    layer0_outputs(4197) <= not a;
    layer0_outputs(4198) <= b and not a;
    layer0_outputs(4199) <= a and not b;
    layer0_outputs(4200) <= b;
    layer0_outputs(4201) <= not b or a;
    layer0_outputs(4202) <= not (a and b);
    layer0_outputs(4203) <= not a;
    layer0_outputs(4204) <= not a;
    layer0_outputs(4205) <= not b or a;
    layer0_outputs(4206) <= a xor b;
    layer0_outputs(4207) <= not b or a;
    layer0_outputs(4208) <= b;
    layer0_outputs(4209) <= a xor b;
    layer0_outputs(4210) <= 1'b1;
    layer0_outputs(4211) <= not (a xor b);
    layer0_outputs(4212) <= not (a or b);
    layer0_outputs(4213) <= a or b;
    layer0_outputs(4214) <= a or b;
    layer0_outputs(4215) <= a and b;
    layer0_outputs(4216) <= not a or b;
    layer0_outputs(4217) <= b;
    layer0_outputs(4218) <= not (a xor b);
    layer0_outputs(4219) <= not (a or b);
    layer0_outputs(4220) <= a and not b;
    layer0_outputs(4221) <= b and not a;
    layer0_outputs(4222) <= not (a or b);
    layer0_outputs(4223) <= b and not a;
    layer0_outputs(4224) <= not a or b;
    layer0_outputs(4225) <= b;
    layer0_outputs(4226) <= not (a or b);
    layer0_outputs(4227) <= a or b;
    layer0_outputs(4228) <= not b;
    layer0_outputs(4229) <= 1'b1;
    layer0_outputs(4230) <= not (a or b);
    layer0_outputs(4231) <= b;
    layer0_outputs(4232) <= b;
    layer0_outputs(4233) <= not a;
    layer0_outputs(4234) <= a and not b;
    layer0_outputs(4235) <= not a;
    layer0_outputs(4236) <= not b;
    layer0_outputs(4237) <= a and not b;
    layer0_outputs(4238) <= not (a or b);
    layer0_outputs(4239) <= not (a or b);
    layer0_outputs(4240) <= not (a xor b);
    layer0_outputs(4241) <= 1'b0;
    layer0_outputs(4242) <= a or b;
    layer0_outputs(4243) <= a xor b;
    layer0_outputs(4244) <= not (a xor b);
    layer0_outputs(4245) <= not a or b;
    layer0_outputs(4246) <= not a;
    layer0_outputs(4247) <= 1'b1;
    layer0_outputs(4248) <= not b or a;
    layer0_outputs(4249) <= not a or b;
    layer0_outputs(4250) <= a;
    layer0_outputs(4251) <= a and b;
    layer0_outputs(4252) <= not a;
    layer0_outputs(4253) <= a xor b;
    layer0_outputs(4254) <= not (a or b);
    layer0_outputs(4255) <= a;
    layer0_outputs(4256) <= 1'b1;
    layer0_outputs(4257) <= b;
    layer0_outputs(4258) <= b and not a;
    layer0_outputs(4259) <= not (a or b);
    layer0_outputs(4260) <= not (a or b);
    layer0_outputs(4261) <= b;
    layer0_outputs(4262) <= not (a xor b);
    layer0_outputs(4263) <= not a;
    layer0_outputs(4264) <= not b;
    layer0_outputs(4265) <= not a or b;
    layer0_outputs(4266) <= not b or a;
    layer0_outputs(4267) <= a xor b;
    layer0_outputs(4268) <= a or b;
    layer0_outputs(4269) <= a xor b;
    layer0_outputs(4270) <= a or b;
    layer0_outputs(4271) <= 1'b1;
    layer0_outputs(4272) <= a or b;
    layer0_outputs(4273) <= a or b;
    layer0_outputs(4274) <= b and not a;
    layer0_outputs(4275) <= not (a xor b);
    layer0_outputs(4276) <= a and not b;
    layer0_outputs(4277) <= a;
    layer0_outputs(4278) <= 1'b1;
    layer0_outputs(4279) <= a or b;
    layer0_outputs(4280) <= a or b;
    layer0_outputs(4281) <= not (a or b);
    layer0_outputs(4282) <= not b;
    layer0_outputs(4283) <= a xor b;
    layer0_outputs(4284) <= a and not b;
    layer0_outputs(4285) <= not b;
    layer0_outputs(4286) <= b;
    layer0_outputs(4287) <= not (a or b);
    layer0_outputs(4288) <= not a;
    layer0_outputs(4289) <= not b;
    layer0_outputs(4290) <= not b or a;
    layer0_outputs(4291) <= not b;
    layer0_outputs(4292) <= a or b;
    layer0_outputs(4293) <= a or b;
    layer0_outputs(4294) <= not (a or b);
    layer0_outputs(4295) <= 1'b1;
    layer0_outputs(4296) <= not (a or b);
    layer0_outputs(4297) <= 1'b1;
    layer0_outputs(4298) <= a or b;
    layer0_outputs(4299) <= not (a xor b);
    layer0_outputs(4300) <= b and not a;
    layer0_outputs(4301) <= a and not b;
    layer0_outputs(4302) <= b and not a;
    layer0_outputs(4303) <= not a;
    layer0_outputs(4304) <= not (a or b);
    layer0_outputs(4305) <= not b;
    layer0_outputs(4306) <= 1'b0;
    layer0_outputs(4307) <= not (a or b);
    layer0_outputs(4308) <= not a or b;
    layer0_outputs(4309) <= a;
    layer0_outputs(4310) <= not a or b;
    layer0_outputs(4311) <= not b;
    layer0_outputs(4312) <= not b;
    layer0_outputs(4313) <= a xor b;
    layer0_outputs(4314) <= not b or a;
    layer0_outputs(4315) <= not b;
    layer0_outputs(4316) <= 1'b0;
    layer0_outputs(4317) <= not (a or b);
    layer0_outputs(4318) <= not a;
    layer0_outputs(4319) <= b;
    layer0_outputs(4320) <= a or b;
    layer0_outputs(4321) <= a and not b;
    layer0_outputs(4322) <= a and b;
    layer0_outputs(4323) <= not (a or b);
    layer0_outputs(4324) <= a or b;
    layer0_outputs(4325) <= not b;
    layer0_outputs(4326) <= a and b;
    layer0_outputs(4327) <= a or b;
    layer0_outputs(4328) <= not (a or b);
    layer0_outputs(4329) <= not a or b;
    layer0_outputs(4330) <= b;
    layer0_outputs(4331) <= a or b;
    layer0_outputs(4332) <= not b or a;
    layer0_outputs(4333) <= a and not b;
    layer0_outputs(4334) <= not (a xor b);
    layer0_outputs(4335) <= a or b;
    layer0_outputs(4336) <= b and not a;
    layer0_outputs(4337) <= not a;
    layer0_outputs(4338) <= a or b;
    layer0_outputs(4339) <= not (a or b);
    layer0_outputs(4340) <= not a;
    layer0_outputs(4341) <= a xor b;
    layer0_outputs(4342) <= b;
    layer0_outputs(4343) <= b;
    layer0_outputs(4344) <= not a;
    layer0_outputs(4345) <= not a or b;
    layer0_outputs(4346) <= not (a or b);
    layer0_outputs(4347) <= b;
    layer0_outputs(4348) <= 1'b0;
    layer0_outputs(4349) <= b;
    layer0_outputs(4350) <= a or b;
    layer0_outputs(4351) <= not b or a;
    layer0_outputs(4352) <= not (a xor b);
    layer0_outputs(4353) <= not (a or b);
    layer0_outputs(4354) <= not b;
    layer0_outputs(4355) <= b;
    layer0_outputs(4356) <= a or b;
    layer0_outputs(4357) <= a or b;
    layer0_outputs(4358) <= not (a xor b);
    layer0_outputs(4359) <= not a or b;
    layer0_outputs(4360) <= not (a and b);
    layer0_outputs(4361) <= not b or a;
    layer0_outputs(4362) <= a or b;
    layer0_outputs(4363) <= not (a or b);
    layer0_outputs(4364) <= b and not a;
    layer0_outputs(4365) <= b;
    layer0_outputs(4366) <= b;
    layer0_outputs(4367) <= 1'b1;
    layer0_outputs(4368) <= a or b;
    layer0_outputs(4369) <= not b or a;
    layer0_outputs(4370) <= a and not b;
    layer0_outputs(4371) <= a xor b;
    layer0_outputs(4372) <= a;
    layer0_outputs(4373) <= not (a or b);
    layer0_outputs(4374) <= a xor b;
    layer0_outputs(4375) <= a or b;
    layer0_outputs(4376) <= not (a xor b);
    layer0_outputs(4377) <= not a;
    layer0_outputs(4378) <= a;
    layer0_outputs(4379) <= not b or a;
    layer0_outputs(4380) <= not a or b;
    layer0_outputs(4381) <= b and not a;
    layer0_outputs(4382) <= a;
    layer0_outputs(4383) <= not b;
    layer0_outputs(4384) <= a and not b;
    layer0_outputs(4385) <= a and b;
    layer0_outputs(4386) <= not b;
    layer0_outputs(4387) <= not a;
    layer0_outputs(4388) <= a and not b;
    layer0_outputs(4389) <= b and not a;
    layer0_outputs(4390) <= a and not b;
    layer0_outputs(4391) <= not (a or b);
    layer0_outputs(4392) <= a or b;
    layer0_outputs(4393) <= not (a or b);
    layer0_outputs(4394) <= not (a or b);
    layer0_outputs(4395) <= not b or a;
    layer0_outputs(4396) <= 1'b1;
    layer0_outputs(4397) <= a or b;
    layer0_outputs(4398) <= not (a or b);
    layer0_outputs(4399) <= a or b;
    layer0_outputs(4400) <= not b;
    layer0_outputs(4401) <= a and not b;
    layer0_outputs(4402) <= a or b;
    layer0_outputs(4403) <= a or b;
    layer0_outputs(4404) <= a or b;
    layer0_outputs(4405) <= a or b;
    layer0_outputs(4406) <= a;
    layer0_outputs(4407) <= not b or a;
    layer0_outputs(4408) <= not (a xor b);
    layer0_outputs(4409) <= not a;
    layer0_outputs(4410) <= b and not a;
    layer0_outputs(4411) <= not a;
    layer0_outputs(4412) <= not (a or b);
    layer0_outputs(4413) <= not (a and b);
    layer0_outputs(4414) <= not a or b;
    layer0_outputs(4415) <= a or b;
    layer0_outputs(4416) <= not a or b;
    layer0_outputs(4417) <= not (a or b);
    layer0_outputs(4418) <= not a or b;
    layer0_outputs(4419) <= a xor b;
    layer0_outputs(4420) <= b and not a;
    layer0_outputs(4421) <= a xor b;
    layer0_outputs(4422) <= a or b;
    layer0_outputs(4423) <= not (a or b);
    layer0_outputs(4424) <= a;
    layer0_outputs(4425) <= not (a or b);
    layer0_outputs(4426) <= b and not a;
    layer0_outputs(4427) <= a xor b;
    layer0_outputs(4428) <= not (a or b);
    layer0_outputs(4429) <= a;
    layer0_outputs(4430) <= not a;
    layer0_outputs(4431) <= not (a or b);
    layer0_outputs(4432) <= not (a or b);
    layer0_outputs(4433) <= not b;
    layer0_outputs(4434) <= a or b;
    layer0_outputs(4435) <= not b or a;
    layer0_outputs(4436) <= a or b;
    layer0_outputs(4437) <= a;
    layer0_outputs(4438) <= not b or a;
    layer0_outputs(4439) <= not (a xor b);
    layer0_outputs(4440) <= not b or a;
    layer0_outputs(4441) <= not (a or b);
    layer0_outputs(4442) <= a;
    layer0_outputs(4443) <= not a;
    layer0_outputs(4444) <= not (a or b);
    layer0_outputs(4445) <= a and b;
    layer0_outputs(4446) <= not a;
    layer0_outputs(4447) <= b;
    layer0_outputs(4448) <= not (a or b);
    layer0_outputs(4449) <= b;
    layer0_outputs(4450) <= b;
    layer0_outputs(4451) <= not b;
    layer0_outputs(4452) <= a xor b;
    layer0_outputs(4453) <= a and not b;
    layer0_outputs(4454) <= a;
    layer0_outputs(4455) <= not a or b;
    layer0_outputs(4456) <= a or b;
    layer0_outputs(4457) <= not b;
    layer0_outputs(4458) <= a or b;
    layer0_outputs(4459) <= a xor b;
    layer0_outputs(4460) <= not (a xor b);
    layer0_outputs(4461) <= a xor b;
    layer0_outputs(4462) <= not a or b;
    layer0_outputs(4463) <= not a or b;
    layer0_outputs(4464) <= not (a and b);
    layer0_outputs(4465) <= a and not b;
    layer0_outputs(4466) <= a;
    layer0_outputs(4467) <= b;
    layer0_outputs(4468) <= a and b;
    layer0_outputs(4469) <= a or b;
    layer0_outputs(4470) <= not (a or b);
    layer0_outputs(4471) <= a and b;
    layer0_outputs(4472) <= a or b;
    layer0_outputs(4473) <= not b or a;
    layer0_outputs(4474) <= not b or a;
    layer0_outputs(4475) <= not (a or b);
    layer0_outputs(4476) <= a and b;
    layer0_outputs(4477) <= 1'b0;
    layer0_outputs(4478) <= not (a xor b);
    layer0_outputs(4479) <= not (a or b);
    layer0_outputs(4480) <= b;
    layer0_outputs(4481) <= 1'b0;
    layer0_outputs(4482) <= not b;
    layer0_outputs(4483) <= not (a xor b);
    layer0_outputs(4484) <= not (a or b);
    layer0_outputs(4485) <= b and not a;
    layer0_outputs(4486) <= b and not a;
    layer0_outputs(4487) <= not a or b;
    layer0_outputs(4488) <= 1'b1;
    layer0_outputs(4489) <= not b or a;
    layer0_outputs(4490) <= 1'b0;
    layer0_outputs(4491) <= not b or a;
    layer0_outputs(4492) <= not (a xor b);
    layer0_outputs(4493) <= a or b;
    layer0_outputs(4494) <= not (a or b);
    layer0_outputs(4495) <= a or b;
    layer0_outputs(4496) <= b;
    layer0_outputs(4497) <= not a or b;
    layer0_outputs(4498) <= not b or a;
    layer0_outputs(4499) <= not (a or b);
    layer0_outputs(4500) <= not (a or b);
    layer0_outputs(4501) <= a xor b;
    layer0_outputs(4502) <= not (a or b);
    layer0_outputs(4503) <= not (a xor b);
    layer0_outputs(4504) <= not a or b;
    layer0_outputs(4505) <= b and not a;
    layer0_outputs(4506) <= a xor b;
    layer0_outputs(4507) <= not b or a;
    layer0_outputs(4508) <= not (a or b);
    layer0_outputs(4509) <= not a;
    layer0_outputs(4510) <= b;
    layer0_outputs(4511) <= b and not a;
    layer0_outputs(4512) <= not (a xor b);
    layer0_outputs(4513) <= not a;
    layer0_outputs(4514) <= not (a xor b);
    layer0_outputs(4515) <= not (a xor b);
    layer0_outputs(4516) <= b;
    layer0_outputs(4517) <= not (a or b);
    layer0_outputs(4518) <= a or b;
    layer0_outputs(4519) <= not b or a;
    layer0_outputs(4520) <= not a;
    layer0_outputs(4521) <= a;
    layer0_outputs(4522) <= not a or b;
    layer0_outputs(4523) <= not (a xor b);
    layer0_outputs(4524) <= a or b;
    layer0_outputs(4525) <= not (a xor b);
    layer0_outputs(4526) <= not b;
    layer0_outputs(4527) <= 1'b0;
    layer0_outputs(4528) <= b and not a;
    layer0_outputs(4529) <= not (a or b);
    layer0_outputs(4530) <= b;
    layer0_outputs(4531) <= not b;
    layer0_outputs(4532) <= a or b;
    layer0_outputs(4533) <= b and not a;
    layer0_outputs(4534) <= a xor b;
    layer0_outputs(4535) <= not (a xor b);
    layer0_outputs(4536) <= a or b;
    layer0_outputs(4537) <= not b;
    layer0_outputs(4538) <= not b;
    layer0_outputs(4539) <= b;
    layer0_outputs(4540) <= a xor b;
    layer0_outputs(4541) <= b;
    layer0_outputs(4542) <= 1'b1;
    layer0_outputs(4543) <= a xor b;
    layer0_outputs(4544) <= b and not a;
    layer0_outputs(4545) <= a or b;
    layer0_outputs(4546) <= not b or a;
    layer0_outputs(4547) <= a and b;
    layer0_outputs(4548) <= not b or a;
    layer0_outputs(4549) <= a or b;
    layer0_outputs(4550) <= not (a xor b);
    layer0_outputs(4551) <= b;
    layer0_outputs(4552) <= a xor b;
    layer0_outputs(4553) <= not (a xor b);
    layer0_outputs(4554) <= not a;
    layer0_outputs(4555) <= a or b;
    layer0_outputs(4556) <= not b or a;
    layer0_outputs(4557) <= b and not a;
    layer0_outputs(4558) <= not b or a;
    layer0_outputs(4559) <= not (a xor b);
    layer0_outputs(4560) <= a and not b;
    layer0_outputs(4561) <= not (a xor b);
    layer0_outputs(4562) <= a and not b;
    layer0_outputs(4563) <= a and not b;
    layer0_outputs(4564) <= not (a xor b);
    layer0_outputs(4565) <= a xor b;
    layer0_outputs(4566) <= not (a or b);
    layer0_outputs(4567) <= not b or a;
    layer0_outputs(4568) <= not (a or b);
    layer0_outputs(4569) <= not a;
    layer0_outputs(4570) <= not b;
    layer0_outputs(4571) <= 1'b0;
    layer0_outputs(4572) <= a xor b;
    layer0_outputs(4573) <= b and not a;
    layer0_outputs(4574) <= not (a or b);
    layer0_outputs(4575) <= not (a or b);
    layer0_outputs(4576) <= not (a xor b);
    layer0_outputs(4577) <= not b;
    layer0_outputs(4578) <= not (a or b);
    layer0_outputs(4579) <= not (a xor b);
    layer0_outputs(4580) <= a;
    layer0_outputs(4581) <= not (a and b);
    layer0_outputs(4582) <= not b or a;
    layer0_outputs(4583) <= not (a or b);
    layer0_outputs(4584) <= a or b;
    layer0_outputs(4585) <= not b;
    layer0_outputs(4586) <= a xor b;
    layer0_outputs(4587) <= a or b;
    layer0_outputs(4588) <= not (a or b);
    layer0_outputs(4589) <= a xor b;
    layer0_outputs(4590) <= a xor b;
    layer0_outputs(4591) <= b and not a;
    layer0_outputs(4592) <= not (a xor b);
    layer0_outputs(4593) <= not b;
    layer0_outputs(4594) <= not (a xor b);
    layer0_outputs(4595) <= not b or a;
    layer0_outputs(4596) <= not a;
    layer0_outputs(4597) <= not b or a;
    layer0_outputs(4598) <= b and not a;
    layer0_outputs(4599) <= b;
    layer0_outputs(4600) <= not b or a;
    layer0_outputs(4601) <= not a or b;
    layer0_outputs(4602) <= not b;
    layer0_outputs(4603) <= b;
    layer0_outputs(4604) <= not (a or b);
    layer0_outputs(4605) <= b and not a;
    layer0_outputs(4606) <= b and not a;
    layer0_outputs(4607) <= 1'b1;
    layer0_outputs(4608) <= a or b;
    layer0_outputs(4609) <= a and not b;
    layer0_outputs(4610) <= not b or a;
    layer0_outputs(4611) <= 1'b1;
    layer0_outputs(4612) <= a or b;
    layer0_outputs(4613) <= b and not a;
    layer0_outputs(4614) <= not (a xor b);
    layer0_outputs(4615) <= a;
    layer0_outputs(4616) <= a or b;
    layer0_outputs(4617) <= not (a or b);
    layer0_outputs(4618) <= not b;
    layer0_outputs(4619) <= b;
    layer0_outputs(4620) <= not a or b;
    layer0_outputs(4621) <= not b;
    layer0_outputs(4622) <= not a or b;
    layer0_outputs(4623) <= not (a or b);
    layer0_outputs(4624) <= a or b;
    layer0_outputs(4625) <= not (a xor b);
    layer0_outputs(4626) <= not (a xor b);
    layer0_outputs(4627) <= not (a or b);
    layer0_outputs(4628) <= not a;
    layer0_outputs(4629) <= not b;
    layer0_outputs(4630) <= not (a xor b);
    layer0_outputs(4631) <= b;
    layer0_outputs(4632) <= not (a xor b);
    layer0_outputs(4633) <= not b or a;
    layer0_outputs(4634) <= not (a or b);
    layer0_outputs(4635) <= not a or b;
    layer0_outputs(4636) <= not b or a;
    layer0_outputs(4637) <= not (a xor b);
    layer0_outputs(4638) <= a or b;
    layer0_outputs(4639) <= a or b;
    layer0_outputs(4640) <= b;
    layer0_outputs(4641) <= not (a xor b);
    layer0_outputs(4642) <= 1'b1;
    layer0_outputs(4643) <= not (a or b);
    layer0_outputs(4644) <= not (a xor b);
    layer0_outputs(4645) <= not (a xor b);
    layer0_outputs(4646) <= not b or a;
    layer0_outputs(4647) <= a xor b;
    layer0_outputs(4648) <= not (a or b);
    layer0_outputs(4649) <= not (a xor b);
    layer0_outputs(4650) <= not (a or b);
    layer0_outputs(4651) <= b;
    layer0_outputs(4652) <= not a;
    layer0_outputs(4653) <= not a or b;
    layer0_outputs(4654) <= not a or b;
    layer0_outputs(4655) <= a or b;
    layer0_outputs(4656) <= not (a or b);
    layer0_outputs(4657) <= a or b;
    layer0_outputs(4658) <= not (a or b);
    layer0_outputs(4659) <= a and not b;
    layer0_outputs(4660) <= a or b;
    layer0_outputs(4661) <= b;
    layer0_outputs(4662) <= not a or b;
    layer0_outputs(4663) <= a;
    layer0_outputs(4664) <= a or b;
    layer0_outputs(4665) <= a or b;
    layer0_outputs(4666) <= b;
    layer0_outputs(4667) <= 1'b1;
    layer0_outputs(4668) <= 1'b0;
    layer0_outputs(4669) <= a or b;
    layer0_outputs(4670) <= not a;
    layer0_outputs(4671) <= 1'b0;
    layer0_outputs(4672) <= a or b;
    layer0_outputs(4673) <= not b;
    layer0_outputs(4674) <= a or b;
    layer0_outputs(4675) <= not (a xor b);
    layer0_outputs(4676) <= not a;
    layer0_outputs(4677) <= a or b;
    layer0_outputs(4678) <= not a;
    layer0_outputs(4679) <= a or b;
    layer0_outputs(4680) <= b;
    layer0_outputs(4681) <= not (a xor b);
    layer0_outputs(4682) <= not b;
    layer0_outputs(4683) <= not a or b;
    layer0_outputs(4684) <= a xor b;
    layer0_outputs(4685) <= not (a or b);
    layer0_outputs(4686) <= b;
    layer0_outputs(4687) <= not (a xor b);
    layer0_outputs(4688) <= b;
    layer0_outputs(4689) <= a or b;
    layer0_outputs(4690) <= not (a or b);
    layer0_outputs(4691) <= not (a xor b);
    layer0_outputs(4692) <= a xor b;
    layer0_outputs(4693) <= b;
    layer0_outputs(4694) <= a or b;
    layer0_outputs(4695) <= not a;
    layer0_outputs(4696) <= not (a or b);
    layer0_outputs(4697) <= not a;
    layer0_outputs(4698) <= not (a or b);
    layer0_outputs(4699) <= a or b;
    layer0_outputs(4700) <= b and not a;
    layer0_outputs(4701) <= not a;
    layer0_outputs(4702) <= not (a and b);
    layer0_outputs(4703) <= not (a or b);
    layer0_outputs(4704) <= not (a or b);
    layer0_outputs(4705) <= not (a xor b);
    layer0_outputs(4706) <= a;
    layer0_outputs(4707) <= b and not a;
    layer0_outputs(4708) <= a;
    layer0_outputs(4709) <= 1'b1;
    layer0_outputs(4710) <= not a or b;
    layer0_outputs(4711) <= a or b;
    layer0_outputs(4712) <= a or b;
    layer0_outputs(4713) <= not b;
    layer0_outputs(4714) <= not a or b;
    layer0_outputs(4715) <= not (a or b);
    layer0_outputs(4716) <= a xor b;
    layer0_outputs(4717) <= 1'b0;
    layer0_outputs(4718) <= a and not b;
    layer0_outputs(4719) <= not (a or b);
    layer0_outputs(4720) <= a;
    layer0_outputs(4721) <= not (a and b);
    layer0_outputs(4722) <= b;
    layer0_outputs(4723) <= a or b;
    layer0_outputs(4724) <= a or b;
    layer0_outputs(4725) <= a xor b;
    layer0_outputs(4726) <= b and not a;
    layer0_outputs(4727) <= not (a xor b);
    layer0_outputs(4728) <= a or b;
    layer0_outputs(4729) <= a and b;
    layer0_outputs(4730) <= not a;
    layer0_outputs(4731) <= not a or b;
    layer0_outputs(4732) <= not (a or b);
    layer0_outputs(4733) <= a xor b;
    layer0_outputs(4734) <= a or b;
    layer0_outputs(4735) <= a xor b;
    layer0_outputs(4736) <= not (a or b);
    layer0_outputs(4737) <= b;
    layer0_outputs(4738) <= 1'b0;
    layer0_outputs(4739) <= not b or a;
    layer0_outputs(4740) <= not (a xor b);
    layer0_outputs(4741) <= not a or b;
    layer0_outputs(4742) <= not b or a;
    layer0_outputs(4743) <= b;
    layer0_outputs(4744) <= a xor b;
    layer0_outputs(4745) <= not (a xor b);
    layer0_outputs(4746) <= not a;
    layer0_outputs(4747) <= not a or b;
    layer0_outputs(4748) <= b and not a;
    layer0_outputs(4749) <= b and not a;
    layer0_outputs(4750) <= a xor b;
    layer0_outputs(4751) <= not (a or b);
    layer0_outputs(4752) <= not a;
    layer0_outputs(4753) <= b;
    layer0_outputs(4754) <= a and b;
    layer0_outputs(4755) <= 1'b1;
    layer0_outputs(4756) <= not (a or b);
    layer0_outputs(4757) <= not a or b;
    layer0_outputs(4758) <= not a;
    layer0_outputs(4759) <= a or b;
    layer0_outputs(4760) <= not b;
    layer0_outputs(4761) <= 1'b0;
    layer0_outputs(4762) <= b and not a;
    layer0_outputs(4763) <= a or b;
    layer0_outputs(4764) <= not (a and b);
    layer0_outputs(4765) <= not (a or b);
    layer0_outputs(4766) <= b;
    layer0_outputs(4767) <= not a or b;
    layer0_outputs(4768) <= b;
    layer0_outputs(4769) <= a;
    layer0_outputs(4770) <= a or b;
    layer0_outputs(4771) <= b;
    layer0_outputs(4772) <= not (a xor b);
    layer0_outputs(4773) <= a or b;
    layer0_outputs(4774) <= a or b;
    layer0_outputs(4775) <= 1'b1;
    layer0_outputs(4776) <= a xor b;
    layer0_outputs(4777) <= a xor b;
    layer0_outputs(4778) <= not a;
    layer0_outputs(4779) <= not a;
    layer0_outputs(4780) <= a or b;
    layer0_outputs(4781) <= not a or b;
    layer0_outputs(4782) <= a xor b;
    layer0_outputs(4783) <= a xor b;
    layer0_outputs(4784) <= not a;
    layer0_outputs(4785) <= not b;
    layer0_outputs(4786) <= a and b;
    layer0_outputs(4787) <= a;
    layer0_outputs(4788) <= not (a or b);
    layer0_outputs(4789) <= a or b;
    layer0_outputs(4790) <= a xor b;
    layer0_outputs(4791) <= not (a xor b);
    layer0_outputs(4792) <= a;
    layer0_outputs(4793) <= a or b;
    layer0_outputs(4794) <= a;
    layer0_outputs(4795) <= not b or a;
    layer0_outputs(4796) <= not (a or b);
    layer0_outputs(4797) <= a and b;
    layer0_outputs(4798) <= b and not a;
    layer0_outputs(4799) <= b;
    layer0_outputs(4800) <= a and not b;
    layer0_outputs(4801) <= not (a xor b);
    layer0_outputs(4802) <= not a or b;
    layer0_outputs(4803) <= a or b;
    layer0_outputs(4804) <= not a or b;
    layer0_outputs(4805) <= not (a xor b);
    layer0_outputs(4806) <= not (a or b);
    layer0_outputs(4807) <= not (a xor b);
    layer0_outputs(4808) <= a xor b;
    layer0_outputs(4809) <= a or b;
    layer0_outputs(4810) <= not (a and b);
    layer0_outputs(4811) <= a xor b;
    layer0_outputs(4812) <= a or b;
    layer0_outputs(4813) <= a or b;
    layer0_outputs(4814) <= a or b;
    layer0_outputs(4815) <= a xor b;
    layer0_outputs(4816) <= a xor b;
    layer0_outputs(4817) <= not (a xor b);
    layer0_outputs(4818) <= not (a xor b);
    layer0_outputs(4819) <= not a;
    layer0_outputs(4820) <= a or b;
    layer0_outputs(4821) <= not (a or b);
    layer0_outputs(4822) <= 1'b0;
    layer0_outputs(4823) <= a xor b;
    layer0_outputs(4824) <= not (a or b);
    layer0_outputs(4825) <= a and not b;
    layer0_outputs(4826) <= not (a or b);
    layer0_outputs(4827) <= not a;
    layer0_outputs(4828) <= a xor b;
    layer0_outputs(4829) <= not b or a;
    layer0_outputs(4830) <= not a;
    layer0_outputs(4831) <= not a or b;
    layer0_outputs(4832) <= not a;
    layer0_outputs(4833) <= a;
    layer0_outputs(4834) <= not (a or b);
    layer0_outputs(4835) <= not (a or b);
    layer0_outputs(4836) <= not b;
    layer0_outputs(4837) <= not (a xor b);
    layer0_outputs(4838) <= not b or a;
    layer0_outputs(4839) <= b and not a;
    layer0_outputs(4840) <= not a;
    layer0_outputs(4841) <= b;
    layer0_outputs(4842) <= a xor b;
    layer0_outputs(4843) <= a xor b;
    layer0_outputs(4844) <= a xor b;
    layer0_outputs(4845) <= not b;
    layer0_outputs(4846) <= not (a xor b);
    layer0_outputs(4847) <= a or b;
    layer0_outputs(4848) <= b and not a;
    layer0_outputs(4849) <= a and b;
    layer0_outputs(4850) <= not (a or b);
    layer0_outputs(4851) <= a;
    layer0_outputs(4852) <= not (a or b);
    layer0_outputs(4853) <= a and not b;
    layer0_outputs(4854) <= not a or b;
    layer0_outputs(4855) <= not (a xor b);
    layer0_outputs(4856) <= a;
    layer0_outputs(4857) <= a or b;
    layer0_outputs(4858) <= not a;
    layer0_outputs(4859) <= not (a or b);
    layer0_outputs(4860) <= a;
    layer0_outputs(4861) <= not (a xor b);
    layer0_outputs(4862) <= not b;
    layer0_outputs(4863) <= not b;
    layer0_outputs(4864) <= a xor b;
    layer0_outputs(4865) <= not (a or b);
    layer0_outputs(4866) <= not (a or b);
    layer0_outputs(4867) <= not b;
    layer0_outputs(4868) <= not (a or b);
    layer0_outputs(4869) <= 1'b0;
    layer0_outputs(4870) <= a or b;
    layer0_outputs(4871) <= 1'b1;
    layer0_outputs(4872) <= b and not a;
    layer0_outputs(4873) <= not (a or b);
    layer0_outputs(4874) <= not (a xor b);
    layer0_outputs(4875) <= b and not a;
    layer0_outputs(4876) <= a or b;
    layer0_outputs(4877) <= 1'b0;
    layer0_outputs(4878) <= not b;
    layer0_outputs(4879) <= a or b;
    layer0_outputs(4880) <= a or b;
    layer0_outputs(4881) <= not (a or b);
    layer0_outputs(4882) <= not b;
    layer0_outputs(4883) <= a xor b;
    layer0_outputs(4884) <= not a;
    layer0_outputs(4885) <= a or b;
    layer0_outputs(4886) <= a;
    layer0_outputs(4887) <= b;
    layer0_outputs(4888) <= not b;
    layer0_outputs(4889) <= not (a or b);
    layer0_outputs(4890) <= a;
    layer0_outputs(4891) <= a or b;
    layer0_outputs(4892) <= not a or b;
    layer0_outputs(4893) <= b and not a;
    layer0_outputs(4894) <= not (a xor b);
    layer0_outputs(4895) <= not b or a;
    layer0_outputs(4896) <= a and not b;
    layer0_outputs(4897) <= a or b;
    layer0_outputs(4898) <= 1'b0;
    layer0_outputs(4899) <= not b;
    layer0_outputs(4900) <= not (a xor b);
    layer0_outputs(4901) <= b and not a;
    layer0_outputs(4902) <= not a;
    layer0_outputs(4903) <= not (a or b);
    layer0_outputs(4904) <= not b;
    layer0_outputs(4905) <= not (a or b);
    layer0_outputs(4906) <= a;
    layer0_outputs(4907) <= a;
    layer0_outputs(4908) <= not b;
    layer0_outputs(4909) <= not (a xor b);
    layer0_outputs(4910) <= a and not b;
    layer0_outputs(4911) <= not b;
    layer0_outputs(4912) <= a;
    layer0_outputs(4913) <= not a or b;
    layer0_outputs(4914) <= 1'b1;
    layer0_outputs(4915) <= not a;
    layer0_outputs(4916) <= 1'b0;
    layer0_outputs(4917) <= not b;
    layer0_outputs(4918) <= b;
    layer0_outputs(4919) <= not a;
    layer0_outputs(4920) <= a;
    layer0_outputs(4921) <= not b or a;
    layer0_outputs(4922) <= b;
    layer0_outputs(4923) <= not b;
    layer0_outputs(4924) <= not (a or b);
    layer0_outputs(4925) <= not b or a;
    layer0_outputs(4926) <= b and not a;
    layer0_outputs(4927) <= b and not a;
    layer0_outputs(4928) <= a xor b;
    layer0_outputs(4929) <= not b;
    layer0_outputs(4930) <= not a or b;
    layer0_outputs(4931) <= b;
    layer0_outputs(4932) <= not (a xor b);
    layer0_outputs(4933) <= b and not a;
    layer0_outputs(4934) <= a or b;
    layer0_outputs(4935) <= b and not a;
    layer0_outputs(4936) <= not a;
    layer0_outputs(4937) <= not (a or b);
    layer0_outputs(4938) <= a or b;
    layer0_outputs(4939) <= a or b;
    layer0_outputs(4940) <= a;
    layer0_outputs(4941) <= a or b;
    layer0_outputs(4942) <= a;
    layer0_outputs(4943) <= b;
    layer0_outputs(4944) <= a or b;
    layer0_outputs(4945) <= not a;
    layer0_outputs(4946) <= a;
    layer0_outputs(4947) <= a and not b;
    layer0_outputs(4948) <= b and not a;
    layer0_outputs(4949) <= a;
    layer0_outputs(4950) <= not (a xor b);
    layer0_outputs(4951) <= b and not a;
    layer0_outputs(4952) <= not b;
    layer0_outputs(4953) <= not (a or b);
    layer0_outputs(4954) <= a xor b;
    layer0_outputs(4955) <= not (a or b);
    layer0_outputs(4956) <= b and not a;
    layer0_outputs(4957) <= a or b;
    layer0_outputs(4958) <= b and not a;
    layer0_outputs(4959) <= 1'b1;
    layer0_outputs(4960) <= not (a xor b);
    layer0_outputs(4961) <= not b;
    layer0_outputs(4962) <= not (a or b);
    layer0_outputs(4963) <= a and not b;
    layer0_outputs(4964) <= b and not a;
    layer0_outputs(4965) <= a xor b;
    layer0_outputs(4966) <= a and not b;
    layer0_outputs(4967) <= a;
    layer0_outputs(4968) <= a or b;
    layer0_outputs(4969) <= b;
    layer0_outputs(4970) <= not (a xor b);
    layer0_outputs(4971) <= a or b;
    layer0_outputs(4972) <= not (a xor b);
    layer0_outputs(4973) <= a and not b;
    layer0_outputs(4974) <= a or b;
    layer0_outputs(4975) <= not (a or b);
    layer0_outputs(4976) <= b and not a;
    layer0_outputs(4977) <= not b or a;
    layer0_outputs(4978) <= not (a or b);
    layer0_outputs(4979) <= a or b;
    layer0_outputs(4980) <= a or b;
    layer0_outputs(4981) <= not (a xor b);
    layer0_outputs(4982) <= a and not b;
    layer0_outputs(4983) <= not (a or b);
    layer0_outputs(4984) <= not (a and b);
    layer0_outputs(4985) <= a or b;
    layer0_outputs(4986) <= a or b;
    layer0_outputs(4987) <= not a;
    layer0_outputs(4988) <= a or b;
    layer0_outputs(4989) <= a;
    layer0_outputs(4990) <= b;
    layer0_outputs(4991) <= not b or a;
    layer0_outputs(4992) <= not b;
    layer0_outputs(4993) <= a and not b;
    layer0_outputs(4994) <= a xor b;
    layer0_outputs(4995) <= a or b;
    layer0_outputs(4996) <= not (a or b);
    layer0_outputs(4997) <= not (a or b);
    layer0_outputs(4998) <= a or b;
    layer0_outputs(4999) <= not (a and b);
    layer0_outputs(5000) <= not (a or b);
    layer0_outputs(5001) <= not b or a;
    layer0_outputs(5002) <= not a;
    layer0_outputs(5003) <= 1'b1;
    layer0_outputs(5004) <= not (a xor b);
    layer0_outputs(5005) <= not b or a;
    layer0_outputs(5006) <= b and not a;
    layer0_outputs(5007) <= a or b;
    layer0_outputs(5008) <= a xor b;
    layer0_outputs(5009) <= a or b;
    layer0_outputs(5010) <= not b;
    layer0_outputs(5011) <= a or b;
    layer0_outputs(5012) <= b and not a;
    layer0_outputs(5013) <= a;
    layer0_outputs(5014) <= a xor b;
    layer0_outputs(5015) <= not (a or b);
    layer0_outputs(5016) <= a or b;
    layer0_outputs(5017) <= not a or b;
    layer0_outputs(5018) <= not (a or b);
    layer0_outputs(5019) <= not (a or b);
    layer0_outputs(5020) <= a xor b;
    layer0_outputs(5021) <= not (a or b);
    layer0_outputs(5022) <= a or b;
    layer0_outputs(5023) <= a xor b;
    layer0_outputs(5024) <= not a or b;
    layer0_outputs(5025) <= not b;
    layer0_outputs(5026) <= a and not b;
    layer0_outputs(5027) <= b and not a;
    layer0_outputs(5028) <= a or b;
    layer0_outputs(5029) <= not a or b;
    layer0_outputs(5030) <= not (a xor b);
    layer0_outputs(5031) <= not (a or b);
    layer0_outputs(5032) <= b and not a;
    layer0_outputs(5033) <= b;
    layer0_outputs(5034) <= a and not b;
    layer0_outputs(5035) <= a;
    layer0_outputs(5036) <= 1'b1;
    layer0_outputs(5037) <= not a;
    layer0_outputs(5038) <= a or b;
    layer0_outputs(5039) <= b and not a;
    layer0_outputs(5040) <= b;
    layer0_outputs(5041) <= a and not b;
    layer0_outputs(5042) <= not b or a;
    layer0_outputs(5043) <= not b or a;
    layer0_outputs(5044) <= not (a and b);
    layer0_outputs(5045) <= not b;
    layer0_outputs(5046) <= not b;
    layer0_outputs(5047) <= not a;
    layer0_outputs(5048) <= a;
    layer0_outputs(5049) <= not b;
    layer0_outputs(5050) <= not a or b;
    layer0_outputs(5051) <= not (a xor b);
    layer0_outputs(5052) <= b;
    layer0_outputs(5053) <= not b or a;
    layer0_outputs(5054) <= not b;
    layer0_outputs(5055) <= not a or b;
    layer0_outputs(5056) <= not (a or b);
    layer0_outputs(5057) <= a or b;
    layer0_outputs(5058) <= a or b;
    layer0_outputs(5059) <= a or b;
    layer0_outputs(5060) <= b;
    layer0_outputs(5061) <= not (a xor b);
    layer0_outputs(5062) <= not a;
    layer0_outputs(5063) <= not (a xor b);
    layer0_outputs(5064) <= a xor b;
    layer0_outputs(5065) <= not (a xor b);
    layer0_outputs(5066) <= not a;
    layer0_outputs(5067) <= a and not b;
    layer0_outputs(5068) <= b;
    layer0_outputs(5069) <= a and b;
    layer0_outputs(5070) <= b and not a;
    layer0_outputs(5071) <= not b or a;
    layer0_outputs(5072) <= b;
    layer0_outputs(5073) <= a or b;
    layer0_outputs(5074) <= a xor b;
    layer0_outputs(5075) <= b;
    layer0_outputs(5076) <= not b;
    layer0_outputs(5077) <= not (a or b);
    layer0_outputs(5078) <= not (a xor b);
    layer0_outputs(5079) <= not b;
    layer0_outputs(5080) <= a xor b;
    layer0_outputs(5081) <= not a or b;
    layer0_outputs(5082) <= a xor b;
    layer0_outputs(5083) <= not a;
    layer0_outputs(5084) <= a or b;
    layer0_outputs(5085) <= a xor b;
    layer0_outputs(5086) <= not (a or b);
    layer0_outputs(5087) <= b;
    layer0_outputs(5088) <= not b;
    layer0_outputs(5089) <= a or b;
    layer0_outputs(5090) <= not (a xor b);
    layer0_outputs(5091) <= 1'b0;
    layer0_outputs(5092) <= not (a and b);
    layer0_outputs(5093) <= b and not a;
    layer0_outputs(5094) <= a;
    layer0_outputs(5095) <= not (a xor b);
    layer0_outputs(5096) <= a xor b;
    layer0_outputs(5097) <= b;
    layer0_outputs(5098) <= not (a or b);
    layer0_outputs(5099) <= a and not b;
    layer0_outputs(5100) <= b and not a;
    layer0_outputs(5101) <= a;
    layer0_outputs(5102) <= a or b;
    layer0_outputs(5103) <= 1'b0;
    layer0_outputs(5104) <= not b;
    layer0_outputs(5105) <= not (a or b);
    layer0_outputs(5106) <= a or b;
    layer0_outputs(5107) <= not a or b;
    layer0_outputs(5108) <= not b;
    layer0_outputs(5109) <= b and not a;
    layer0_outputs(5110) <= not (a or b);
    layer0_outputs(5111) <= not b;
    layer0_outputs(5112) <= a or b;
    layer0_outputs(5113) <= not (a or b);
    layer0_outputs(5114) <= a;
    layer0_outputs(5115) <= a and not b;
    layer0_outputs(5116) <= 1'b0;
    layer0_outputs(5117) <= b;
    layer0_outputs(5118) <= not a or b;
    layer0_outputs(5119) <= not (a xor b);
    layer0_outputs(5120) <= a xor b;
    layer0_outputs(5121) <= a;
    layer0_outputs(5122) <= a xor b;
    layer0_outputs(5123) <= not (a and b);
    layer0_outputs(5124) <= b and not a;
    layer0_outputs(5125) <= b and not a;
    layer0_outputs(5126) <= not (a or b);
    layer0_outputs(5127) <= b;
    layer0_outputs(5128) <= a and not b;
    layer0_outputs(5129) <= not (a or b);
    layer0_outputs(5130) <= not (a or b);
    layer0_outputs(5131) <= not (a or b);
    layer0_outputs(5132) <= not b or a;
    layer0_outputs(5133) <= not b or a;
    layer0_outputs(5134) <= b and not a;
    layer0_outputs(5135) <= not (a or b);
    layer0_outputs(5136) <= b;
    layer0_outputs(5137) <= a xor b;
    layer0_outputs(5138) <= not (a or b);
    layer0_outputs(5139) <= a xor b;
    layer0_outputs(5140) <= not a or b;
    layer0_outputs(5141) <= a or b;
    layer0_outputs(5142) <= a xor b;
    layer0_outputs(5143) <= not b;
    layer0_outputs(5144) <= a and not b;
    layer0_outputs(5145) <= a;
    layer0_outputs(5146) <= b and not a;
    layer0_outputs(5147) <= a xor b;
    layer0_outputs(5148) <= not (a or b);
    layer0_outputs(5149) <= not b;
    layer0_outputs(5150) <= a or b;
    layer0_outputs(5151) <= not (a or b);
    layer0_outputs(5152) <= a xor b;
    layer0_outputs(5153) <= not a;
    layer0_outputs(5154) <= b and not a;
    layer0_outputs(5155) <= not (a or b);
    layer0_outputs(5156) <= not (a or b);
    layer0_outputs(5157) <= b and not a;
    layer0_outputs(5158) <= a or b;
    layer0_outputs(5159) <= a or b;
    layer0_outputs(5160) <= not a;
    layer0_outputs(5161) <= a or b;
    layer0_outputs(5162) <= b;
    layer0_outputs(5163) <= not b;
    layer0_outputs(5164) <= not (a or b);
    layer0_outputs(5165) <= a or b;
    layer0_outputs(5166) <= not b;
    layer0_outputs(5167) <= not (a xor b);
    layer0_outputs(5168) <= a;
    layer0_outputs(5169) <= a or b;
    layer0_outputs(5170) <= b;
    layer0_outputs(5171) <= b;
    layer0_outputs(5172) <= a and b;
    layer0_outputs(5173) <= b;
    layer0_outputs(5174) <= a;
    layer0_outputs(5175) <= a and not b;
    layer0_outputs(5176) <= b;
    layer0_outputs(5177) <= a or b;
    layer0_outputs(5178) <= a or b;
    layer0_outputs(5179) <= a and not b;
    layer0_outputs(5180) <= not b or a;
    layer0_outputs(5181) <= a xor b;
    layer0_outputs(5182) <= not (a or b);
    layer0_outputs(5183) <= not (a or b);
    layer0_outputs(5184) <= b and not a;
    layer0_outputs(5185) <= a and b;
    layer0_outputs(5186) <= not (a xor b);
    layer0_outputs(5187) <= a and not b;
    layer0_outputs(5188) <= 1'b1;
    layer0_outputs(5189) <= b and not a;
    layer0_outputs(5190) <= 1'b1;
    layer0_outputs(5191) <= b and not a;
    layer0_outputs(5192) <= a and not b;
    layer0_outputs(5193) <= 1'b0;
    layer0_outputs(5194) <= b;
    layer0_outputs(5195) <= not b or a;
    layer0_outputs(5196) <= not a or b;
    layer0_outputs(5197) <= not (a or b);
    layer0_outputs(5198) <= a xor b;
    layer0_outputs(5199) <= not (a and b);
    layer0_outputs(5200) <= 1'b1;
    layer0_outputs(5201) <= b and not a;
    layer0_outputs(5202) <= not (a xor b);
    layer0_outputs(5203) <= not (a and b);
    layer0_outputs(5204) <= a and not b;
    layer0_outputs(5205) <= not a or b;
    layer0_outputs(5206) <= not (a or b);
    layer0_outputs(5207) <= a or b;
    layer0_outputs(5208) <= not (a and b);
    layer0_outputs(5209) <= not a;
    layer0_outputs(5210) <= b;
    layer0_outputs(5211) <= not (a xor b);
    layer0_outputs(5212) <= a;
    layer0_outputs(5213) <= not (a xor b);
    layer0_outputs(5214) <= not a or b;
    layer0_outputs(5215) <= b;
    layer0_outputs(5216) <= a xor b;
    layer0_outputs(5217) <= not (a or b);
    layer0_outputs(5218) <= not (a xor b);
    layer0_outputs(5219) <= not (a or b);
    layer0_outputs(5220) <= a xor b;
    layer0_outputs(5221) <= a or b;
    layer0_outputs(5222) <= b and not a;
    layer0_outputs(5223) <= not b;
    layer0_outputs(5224) <= not (a or b);
    layer0_outputs(5225) <= b;
    layer0_outputs(5226) <= a or b;
    layer0_outputs(5227) <= not b or a;
    layer0_outputs(5228) <= a or b;
    layer0_outputs(5229) <= a xor b;
    layer0_outputs(5230) <= not a or b;
    layer0_outputs(5231) <= a xor b;
    layer0_outputs(5232) <= b and not a;
    layer0_outputs(5233) <= a xor b;
    layer0_outputs(5234) <= a;
    layer0_outputs(5235) <= a or b;
    layer0_outputs(5236) <= b and not a;
    layer0_outputs(5237) <= a xor b;
    layer0_outputs(5238) <= not (a or b);
    layer0_outputs(5239) <= b and not a;
    layer0_outputs(5240) <= not (a or b);
    layer0_outputs(5241) <= b;
    layer0_outputs(5242) <= not a or b;
    layer0_outputs(5243) <= not b or a;
    layer0_outputs(5244) <= a or b;
    layer0_outputs(5245) <= not a;
    layer0_outputs(5246) <= a;
    layer0_outputs(5247) <= not (a or b);
    layer0_outputs(5248) <= not (a or b);
    layer0_outputs(5249) <= not a or b;
    layer0_outputs(5250) <= a or b;
    layer0_outputs(5251) <= a or b;
    layer0_outputs(5252) <= a or b;
    layer0_outputs(5253) <= a xor b;
    layer0_outputs(5254) <= b and not a;
    layer0_outputs(5255) <= not (a or b);
    layer0_outputs(5256) <= not a;
    layer0_outputs(5257) <= a xor b;
    layer0_outputs(5258) <= not (a or b);
    layer0_outputs(5259) <= not b or a;
    layer0_outputs(5260) <= not (a or b);
    layer0_outputs(5261) <= a;
    layer0_outputs(5262) <= 1'b0;
    layer0_outputs(5263) <= a or b;
    layer0_outputs(5264) <= 1'b1;
    layer0_outputs(5265) <= not (a xor b);
    layer0_outputs(5266) <= not b;
    layer0_outputs(5267) <= not b or a;
    layer0_outputs(5268) <= a or b;
    layer0_outputs(5269) <= a or b;
    layer0_outputs(5270) <= not (a xor b);
    layer0_outputs(5271) <= not a;
    layer0_outputs(5272) <= b;
    layer0_outputs(5273) <= b;
    layer0_outputs(5274) <= not (a xor b);
    layer0_outputs(5275) <= a xor b;
    layer0_outputs(5276) <= 1'b1;
    layer0_outputs(5277) <= b and not a;
    layer0_outputs(5278) <= not b or a;
    layer0_outputs(5279) <= not (a or b);
    layer0_outputs(5280) <= not b or a;
    layer0_outputs(5281) <= not b;
    layer0_outputs(5282) <= a or b;
    layer0_outputs(5283) <= not (a xor b);
    layer0_outputs(5284) <= not (a xor b);
    layer0_outputs(5285) <= not (a xor b);
    layer0_outputs(5286) <= not a;
    layer0_outputs(5287) <= 1'b0;
    layer0_outputs(5288) <= not b or a;
    layer0_outputs(5289) <= a xor b;
    layer0_outputs(5290) <= not a;
    layer0_outputs(5291) <= b;
    layer0_outputs(5292) <= not b;
    layer0_outputs(5293) <= b;
    layer0_outputs(5294) <= a and not b;
    layer0_outputs(5295) <= a;
    layer0_outputs(5296) <= not b;
    layer0_outputs(5297) <= a xor b;
    layer0_outputs(5298) <= not a;
    layer0_outputs(5299) <= not a or b;
    layer0_outputs(5300) <= a;
    layer0_outputs(5301) <= not (a or b);
    layer0_outputs(5302) <= not b or a;
    layer0_outputs(5303) <= b and not a;
    layer0_outputs(5304) <= a;
    layer0_outputs(5305) <= not b;
    layer0_outputs(5306) <= a or b;
    layer0_outputs(5307) <= not (a or b);
    layer0_outputs(5308) <= not a or b;
    layer0_outputs(5309) <= not a;
    layer0_outputs(5310) <= not (a xor b);
    layer0_outputs(5311) <= not (a xor b);
    layer0_outputs(5312) <= not (a or b);
    layer0_outputs(5313) <= a xor b;
    layer0_outputs(5314) <= b;
    layer0_outputs(5315) <= not a;
    layer0_outputs(5316) <= b;
    layer0_outputs(5317) <= b;
    layer0_outputs(5318) <= b;
    layer0_outputs(5319) <= a xor b;
    layer0_outputs(5320) <= not a;
    layer0_outputs(5321) <= a or b;
    layer0_outputs(5322) <= not (a or b);
    layer0_outputs(5323) <= not a;
    layer0_outputs(5324) <= not a;
    layer0_outputs(5325) <= not (a or b);
    layer0_outputs(5326) <= not a;
    layer0_outputs(5327) <= not a or b;
    layer0_outputs(5328) <= a and not b;
    layer0_outputs(5329) <= not (a or b);
    layer0_outputs(5330) <= b;
    layer0_outputs(5331) <= not (a or b);
    layer0_outputs(5332) <= not b or a;
    layer0_outputs(5333) <= not (a and b);
    layer0_outputs(5334) <= a;
    layer0_outputs(5335) <= a xor b;
    layer0_outputs(5336) <= not b or a;
    layer0_outputs(5337) <= not a or b;
    layer0_outputs(5338) <= b and not a;
    layer0_outputs(5339) <= a and not b;
    layer0_outputs(5340) <= a or b;
    layer0_outputs(5341) <= a xor b;
    layer0_outputs(5342) <= a;
    layer0_outputs(5343) <= a;
    layer0_outputs(5344) <= not (a or b);
    layer0_outputs(5345) <= 1'b1;
    layer0_outputs(5346) <= not b;
    layer0_outputs(5347) <= a xor b;
    layer0_outputs(5348) <= not (a or b);
    layer0_outputs(5349) <= not (a xor b);
    layer0_outputs(5350) <= not a or b;
    layer0_outputs(5351) <= b;
    layer0_outputs(5352) <= a or b;
    layer0_outputs(5353) <= not (a or b);
    layer0_outputs(5354) <= not b or a;
    layer0_outputs(5355) <= a;
    layer0_outputs(5356) <= not (a or b);
    layer0_outputs(5357) <= not b or a;
    layer0_outputs(5358) <= not (a xor b);
    layer0_outputs(5359) <= a or b;
    layer0_outputs(5360) <= not (a or b);
    layer0_outputs(5361) <= a or b;
    layer0_outputs(5362) <= b;
    layer0_outputs(5363) <= a;
    layer0_outputs(5364) <= a;
    layer0_outputs(5365) <= not (a xor b);
    layer0_outputs(5366) <= a or b;
    layer0_outputs(5367) <= not (a xor b);
    layer0_outputs(5368) <= not (a or b);
    layer0_outputs(5369) <= not b;
    layer0_outputs(5370) <= not a or b;
    layer0_outputs(5371) <= 1'b0;
    layer0_outputs(5372) <= not (a xor b);
    layer0_outputs(5373) <= 1'b1;
    layer0_outputs(5374) <= not (a or b);
    layer0_outputs(5375) <= not (a and b);
    layer0_outputs(5376) <= b;
    layer0_outputs(5377) <= a and not b;
    layer0_outputs(5378) <= a xor b;
    layer0_outputs(5379) <= a or b;
    layer0_outputs(5380) <= a xor b;
    layer0_outputs(5381) <= not (a or b);
    layer0_outputs(5382) <= not (a or b);
    layer0_outputs(5383) <= b;
    layer0_outputs(5384) <= a or b;
    layer0_outputs(5385) <= not a or b;
    layer0_outputs(5386) <= a or b;
    layer0_outputs(5387) <= not a or b;
    layer0_outputs(5388) <= not b or a;
    layer0_outputs(5389) <= not (a xor b);
    layer0_outputs(5390) <= not a;
    layer0_outputs(5391) <= not b;
    layer0_outputs(5392) <= not (a and b);
    layer0_outputs(5393) <= a;
    layer0_outputs(5394) <= not (a or b);
    layer0_outputs(5395) <= 1'b0;
    layer0_outputs(5396) <= a xor b;
    layer0_outputs(5397) <= a;
    layer0_outputs(5398) <= b;
    layer0_outputs(5399) <= not b or a;
    layer0_outputs(5400) <= b;
    layer0_outputs(5401) <= a and not b;
    layer0_outputs(5402) <= 1'b0;
    layer0_outputs(5403) <= not b;
    layer0_outputs(5404) <= not (a or b);
    layer0_outputs(5405) <= a or b;
    layer0_outputs(5406) <= a or b;
    layer0_outputs(5407) <= not a;
    layer0_outputs(5408) <= not (a or b);
    layer0_outputs(5409) <= not (a and b);
    layer0_outputs(5410) <= a or b;
    layer0_outputs(5411) <= b;
    layer0_outputs(5412) <= b;
    layer0_outputs(5413) <= a xor b;
    layer0_outputs(5414) <= not b;
    layer0_outputs(5415) <= not b;
    layer0_outputs(5416) <= not b or a;
    layer0_outputs(5417) <= not (a and b);
    layer0_outputs(5418) <= not a;
    layer0_outputs(5419) <= a xor b;
    layer0_outputs(5420) <= not a or b;
    layer0_outputs(5421) <= a or b;
    layer0_outputs(5422) <= not b;
    layer0_outputs(5423) <= not b or a;
    layer0_outputs(5424) <= not (a or b);
    layer0_outputs(5425) <= a and not b;
    layer0_outputs(5426) <= a or b;
    layer0_outputs(5427) <= not (a xor b);
    layer0_outputs(5428) <= not b or a;
    layer0_outputs(5429) <= not (a or b);
    layer0_outputs(5430) <= not b or a;
    layer0_outputs(5431) <= not a;
    layer0_outputs(5432) <= a and not b;
    layer0_outputs(5433) <= a xor b;
    layer0_outputs(5434) <= not (a or b);
    layer0_outputs(5435) <= not (a or b);
    layer0_outputs(5436) <= not (a or b);
    layer0_outputs(5437) <= a and b;
    layer0_outputs(5438) <= b and not a;
    layer0_outputs(5439) <= not a or b;
    layer0_outputs(5440) <= a;
    layer0_outputs(5441) <= not (a or b);
    layer0_outputs(5442) <= a or b;
    layer0_outputs(5443) <= b;
    layer0_outputs(5444) <= b;
    layer0_outputs(5445) <= a or b;
    layer0_outputs(5446) <= not (a or b);
    layer0_outputs(5447) <= a and not b;
    layer0_outputs(5448) <= a xor b;
    layer0_outputs(5449) <= a xor b;
    layer0_outputs(5450) <= b;
    layer0_outputs(5451) <= not b;
    layer0_outputs(5452) <= b and not a;
    layer0_outputs(5453) <= b;
    layer0_outputs(5454) <= not (a or b);
    layer0_outputs(5455) <= a xor b;
    layer0_outputs(5456) <= not (a or b);
    layer0_outputs(5457) <= a;
    layer0_outputs(5458) <= a or b;
    layer0_outputs(5459) <= b;
    layer0_outputs(5460) <= not a or b;
    layer0_outputs(5461) <= a;
    layer0_outputs(5462) <= not (a or b);
    layer0_outputs(5463) <= not (a or b);
    layer0_outputs(5464) <= not a or b;
    layer0_outputs(5465) <= not (a xor b);
    layer0_outputs(5466) <= not a or b;
    layer0_outputs(5467) <= not (a or b);
    layer0_outputs(5468) <= a or b;
    layer0_outputs(5469) <= not a;
    layer0_outputs(5470) <= not b;
    layer0_outputs(5471) <= not a;
    layer0_outputs(5472) <= a xor b;
    layer0_outputs(5473) <= not (a xor b);
    layer0_outputs(5474) <= a xor b;
    layer0_outputs(5475) <= b;
    layer0_outputs(5476) <= not a or b;
    layer0_outputs(5477) <= a or b;
    layer0_outputs(5478) <= not a;
    layer0_outputs(5479) <= not b;
    layer0_outputs(5480) <= not (a or b);
    layer0_outputs(5481) <= not (a xor b);
    layer0_outputs(5482) <= a xor b;
    layer0_outputs(5483) <= a or b;
    layer0_outputs(5484) <= a and b;
    layer0_outputs(5485) <= b and not a;
    layer0_outputs(5486) <= a xor b;
    layer0_outputs(5487) <= a and not b;
    layer0_outputs(5488) <= a;
    layer0_outputs(5489) <= not b;
    layer0_outputs(5490) <= a;
    layer0_outputs(5491) <= a and b;
    layer0_outputs(5492) <= a or b;
    layer0_outputs(5493) <= not a or b;
    layer0_outputs(5494) <= b;
    layer0_outputs(5495) <= a or b;
    layer0_outputs(5496) <= a and not b;
    layer0_outputs(5497) <= a or b;
    layer0_outputs(5498) <= not (a xor b);
    layer0_outputs(5499) <= a and not b;
    layer0_outputs(5500) <= not (a or b);
    layer0_outputs(5501) <= 1'b0;
    layer0_outputs(5502) <= not a;
    layer0_outputs(5503) <= a;
    layer0_outputs(5504) <= b and not a;
    layer0_outputs(5505) <= not (a and b);
    layer0_outputs(5506) <= not a or b;
    layer0_outputs(5507) <= a xor b;
    layer0_outputs(5508) <= not a;
    layer0_outputs(5509) <= 1'b1;
    layer0_outputs(5510) <= not a;
    layer0_outputs(5511) <= a or b;
    layer0_outputs(5512) <= not a;
    layer0_outputs(5513) <= not (a or b);
    layer0_outputs(5514) <= not (a or b);
    layer0_outputs(5515) <= not (a or b);
    layer0_outputs(5516) <= not b or a;
    layer0_outputs(5517) <= not b;
    layer0_outputs(5518) <= not (a or b);
    layer0_outputs(5519) <= not (a xor b);
    layer0_outputs(5520) <= 1'b0;
    layer0_outputs(5521) <= not b;
    layer0_outputs(5522) <= not a;
    layer0_outputs(5523) <= a;
    layer0_outputs(5524) <= not (a and b);
    layer0_outputs(5525) <= a or b;
    layer0_outputs(5526) <= a or b;
    layer0_outputs(5527) <= b and not a;
    layer0_outputs(5528) <= a or b;
    layer0_outputs(5529) <= a and b;
    layer0_outputs(5530) <= a xor b;
    layer0_outputs(5531) <= a and not b;
    layer0_outputs(5532) <= not b;
    layer0_outputs(5533) <= b;
    layer0_outputs(5534) <= b;
    layer0_outputs(5535) <= a or b;
    layer0_outputs(5536) <= a or b;
    layer0_outputs(5537) <= not (a xor b);
    layer0_outputs(5538) <= not a or b;
    layer0_outputs(5539) <= 1'b0;
    layer0_outputs(5540) <= a;
    layer0_outputs(5541) <= a xor b;
    layer0_outputs(5542) <= b and not a;
    layer0_outputs(5543) <= b;
    layer0_outputs(5544) <= a or b;
    layer0_outputs(5545) <= a or b;
    layer0_outputs(5546) <= b;
    layer0_outputs(5547) <= b and not a;
    layer0_outputs(5548) <= not (a or b);
    layer0_outputs(5549) <= a and not b;
    layer0_outputs(5550) <= a xor b;
    layer0_outputs(5551) <= a xor b;
    layer0_outputs(5552) <= not (a xor b);
    layer0_outputs(5553) <= not (a or b);
    layer0_outputs(5554) <= a and not b;
    layer0_outputs(5555) <= 1'b0;
    layer0_outputs(5556) <= not (a or b);
    layer0_outputs(5557) <= not a;
    layer0_outputs(5558) <= b and not a;
    layer0_outputs(5559) <= a xor b;
    layer0_outputs(5560) <= not (a or b);
    layer0_outputs(5561) <= not (a or b);
    layer0_outputs(5562) <= not (a or b);
    layer0_outputs(5563) <= a and not b;
    layer0_outputs(5564) <= b and not a;
    layer0_outputs(5565) <= a and b;
    layer0_outputs(5566) <= b;
    layer0_outputs(5567) <= not a;
    layer0_outputs(5568) <= not (a xor b);
    layer0_outputs(5569) <= not b or a;
    layer0_outputs(5570) <= 1'b1;
    layer0_outputs(5571) <= b;
    layer0_outputs(5572) <= a;
    layer0_outputs(5573) <= a and not b;
    layer0_outputs(5574) <= not (a or b);
    layer0_outputs(5575) <= a or b;
    layer0_outputs(5576) <= a or b;
    layer0_outputs(5577) <= not (a xor b);
    layer0_outputs(5578) <= not (a or b);
    layer0_outputs(5579) <= 1'b1;
    layer0_outputs(5580) <= b and not a;
    layer0_outputs(5581) <= not a or b;
    layer0_outputs(5582) <= not (a or b);
    layer0_outputs(5583) <= a;
    layer0_outputs(5584) <= not a or b;
    layer0_outputs(5585) <= a xor b;
    layer0_outputs(5586) <= not (a or b);
    layer0_outputs(5587) <= a and not b;
    layer0_outputs(5588) <= a xor b;
    layer0_outputs(5589) <= not a;
    layer0_outputs(5590) <= a xor b;
    layer0_outputs(5591) <= a xor b;
    layer0_outputs(5592) <= b;
    layer0_outputs(5593) <= a or b;
    layer0_outputs(5594) <= not (a xor b);
    layer0_outputs(5595) <= not (a xor b);
    layer0_outputs(5596) <= not b or a;
    layer0_outputs(5597) <= not (a xor b);
    layer0_outputs(5598) <= a or b;
    layer0_outputs(5599) <= not (a xor b);
    layer0_outputs(5600) <= a and not b;
    layer0_outputs(5601) <= not (a or b);
    layer0_outputs(5602) <= not b or a;
    layer0_outputs(5603) <= not b;
    layer0_outputs(5604) <= not (a or b);
    layer0_outputs(5605) <= not a or b;
    layer0_outputs(5606) <= 1'b1;
    layer0_outputs(5607) <= not b;
    layer0_outputs(5608) <= not a;
    layer0_outputs(5609) <= not b;
    layer0_outputs(5610) <= a or b;
    layer0_outputs(5611) <= not b;
    layer0_outputs(5612) <= 1'b1;
    layer0_outputs(5613) <= not b;
    layer0_outputs(5614) <= a or b;
    layer0_outputs(5615) <= b and not a;
    layer0_outputs(5616) <= not (a xor b);
    layer0_outputs(5617) <= a xor b;
    layer0_outputs(5618) <= 1'b0;
    layer0_outputs(5619) <= a;
    layer0_outputs(5620) <= 1'b1;
    layer0_outputs(5621) <= a or b;
    layer0_outputs(5622) <= a;
    layer0_outputs(5623) <= a or b;
    layer0_outputs(5624) <= not (a or b);
    layer0_outputs(5625) <= not (a or b);
    layer0_outputs(5626) <= not b;
    layer0_outputs(5627) <= not (a or b);
    layer0_outputs(5628) <= a;
    layer0_outputs(5629) <= a;
    layer0_outputs(5630) <= not a;
    layer0_outputs(5631) <= a and not b;
    layer0_outputs(5632) <= not (a xor b);
    layer0_outputs(5633) <= a and not b;
    layer0_outputs(5634) <= not b;
    layer0_outputs(5635) <= b;
    layer0_outputs(5636) <= b;
    layer0_outputs(5637) <= not a;
    layer0_outputs(5638) <= a xor b;
    layer0_outputs(5639) <= a xor b;
    layer0_outputs(5640) <= not b;
    layer0_outputs(5641) <= not a;
    layer0_outputs(5642) <= not (a or b);
    layer0_outputs(5643) <= a xor b;
    layer0_outputs(5644) <= a xor b;
    layer0_outputs(5645) <= a or b;
    layer0_outputs(5646) <= b and not a;
    layer0_outputs(5647) <= b;
    layer0_outputs(5648) <= b and not a;
    layer0_outputs(5649) <= 1'b1;
    layer0_outputs(5650) <= not (a or b);
    layer0_outputs(5651) <= a;
    layer0_outputs(5652) <= a or b;
    layer0_outputs(5653) <= not (a xor b);
    layer0_outputs(5654) <= not (a xor b);
    layer0_outputs(5655) <= not b;
    layer0_outputs(5656) <= a or b;
    layer0_outputs(5657) <= 1'b0;
    layer0_outputs(5658) <= a and not b;
    layer0_outputs(5659) <= a or b;
    layer0_outputs(5660) <= not (a or b);
    layer0_outputs(5661) <= a xor b;
    layer0_outputs(5662) <= a or b;
    layer0_outputs(5663) <= not (a or b);
    layer0_outputs(5664) <= not b;
    layer0_outputs(5665) <= a or b;
    layer0_outputs(5666) <= not a;
    layer0_outputs(5667) <= not (a xor b);
    layer0_outputs(5668) <= a or b;
    layer0_outputs(5669) <= not b;
    layer0_outputs(5670) <= a;
    layer0_outputs(5671) <= not (a or b);
    layer0_outputs(5672) <= not a or b;
    layer0_outputs(5673) <= b and not a;
    layer0_outputs(5674) <= not b;
    layer0_outputs(5675) <= a;
    layer0_outputs(5676) <= a or b;
    layer0_outputs(5677) <= a xor b;
    layer0_outputs(5678) <= not a or b;
    layer0_outputs(5679) <= a xor b;
    layer0_outputs(5680) <= not (a or b);
    layer0_outputs(5681) <= a or b;
    layer0_outputs(5682) <= a xor b;
    layer0_outputs(5683) <= not (a or b);
    layer0_outputs(5684) <= not a;
    layer0_outputs(5685) <= a xor b;
    layer0_outputs(5686) <= b;
    layer0_outputs(5687) <= a or b;
    layer0_outputs(5688) <= not (a or b);
    layer0_outputs(5689) <= not (a xor b);
    layer0_outputs(5690) <= not (a or b);
    layer0_outputs(5691) <= not a;
    layer0_outputs(5692) <= a and not b;
    layer0_outputs(5693) <= b and not a;
    layer0_outputs(5694) <= b;
    layer0_outputs(5695) <= not a or b;
    layer0_outputs(5696) <= a;
    layer0_outputs(5697) <= not b or a;
    layer0_outputs(5698) <= not a or b;
    layer0_outputs(5699) <= a and not b;
    layer0_outputs(5700) <= a or b;
    layer0_outputs(5701) <= not a or b;
    layer0_outputs(5702) <= a and not b;
    layer0_outputs(5703) <= not b;
    layer0_outputs(5704) <= b and not a;
    layer0_outputs(5705) <= 1'b0;
    layer0_outputs(5706) <= not b;
    layer0_outputs(5707) <= b;
    layer0_outputs(5708) <= not (a or b);
    layer0_outputs(5709) <= b;
    layer0_outputs(5710) <= a xor b;
    layer0_outputs(5711) <= 1'b1;
    layer0_outputs(5712) <= not (a and b);
    layer0_outputs(5713) <= a and b;
    layer0_outputs(5714) <= a xor b;
    layer0_outputs(5715) <= a;
    layer0_outputs(5716) <= a or b;
    layer0_outputs(5717) <= a;
    layer0_outputs(5718) <= a xor b;
    layer0_outputs(5719) <= not b;
    layer0_outputs(5720) <= b and not a;
    layer0_outputs(5721) <= 1'b1;
    layer0_outputs(5722) <= not b;
    layer0_outputs(5723) <= not b;
    layer0_outputs(5724) <= a and b;
    layer0_outputs(5725) <= a or b;
    layer0_outputs(5726) <= a or b;
    layer0_outputs(5727) <= a or b;
    layer0_outputs(5728) <= not b;
    layer0_outputs(5729) <= a xor b;
    layer0_outputs(5730) <= not (a or b);
    layer0_outputs(5731) <= not a;
    layer0_outputs(5732) <= not (a or b);
    layer0_outputs(5733) <= not b or a;
    layer0_outputs(5734) <= b and not a;
    layer0_outputs(5735) <= a or b;
    layer0_outputs(5736) <= a and b;
    layer0_outputs(5737) <= not b or a;
    layer0_outputs(5738) <= b;
    layer0_outputs(5739) <= not b or a;
    layer0_outputs(5740) <= b;
    layer0_outputs(5741) <= not a;
    layer0_outputs(5742) <= a and not b;
    layer0_outputs(5743) <= not b or a;
    layer0_outputs(5744) <= a;
    layer0_outputs(5745) <= b;
    layer0_outputs(5746) <= not a;
    layer0_outputs(5747) <= not (a xor b);
    layer0_outputs(5748) <= a or b;
    layer0_outputs(5749) <= a xor b;
    layer0_outputs(5750) <= a and not b;
    layer0_outputs(5751) <= a;
    layer0_outputs(5752) <= not a;
    layer0_outputs(5753) <= a and not b;
    layer0_outputs(5754) <= not (a or b);
    layer0_outputs(5755) <= a xor b;
    layer0_outputs(5756) <= not a;
    layer0_outputs(5757) <= a and b;
    layer0_outputs(5758) <= not b or a;
    layer0_outputs(5759) <= b;
    layer0_outputs(5760) <= not a or b;
    layer0_outputs(5761) <= a and not b;
    layer0_outputs(5762) <= a xor b;
    layer0_outputs(5763) <= not a or b;
    layer0_outputs(5764) <= b;
    layer0_outputs(5765) <= a and not b;
    layer0_outputs(5766) <= a or b;
    layer0_outputs(5767) <= not a;
    layer0_outputs(5768) <= not a or b;
    layer0_outputs(5769) <= not b or a;
    layer0_outputs(5770) <= not a;
    layer0_outputs(5771) <= not (a xor b);
    layer0_outputs(5772) <= a or b;
    layer0_outputs(5773) <= not (a or b);
    layer0_outputs(5774) <= 1'b1;
    layer0_outputs(5775) <= a or b;
    layer0_outputs(5776) <= not (a or b);
    layer0_outputs(5777) <= a and not b;
    layer0_outputs(5778) <= a xor b;
    layer0_outputs(5779) <= a xor b;
    layer0_outputs(5780) <= a xor b;
    layer0_outputs(5781) <= a or b;
    layer0_outputs(5782) <= a and not b;
    layer0_outputs(5783) <= a;
    layer0_outputs(5784) <= b and not a;
    layer0_outputs(5785) <= not (a or b);
    layer0_outputs(5786) <= not a;
    layer0_outputs(5787) <= not (a or b);
    layer0_outputs(5788) <= a;
    layer0_outputs(5789) <= not (a or b);
    layer0_outputs(5790) <= not a or b;
    layer0_outputs(5791) <= a and not b;
    layer0_outputs(5792) <= not a;
    layer0_outputs(5793) <= b and not a;
    layer0_outputs(5794) <= not a;
    layer0_outputs(5795) <= not (a or b);
    layer0_outputs(5796) <= a and not b;
    layer0_outputs(5797) <= not (a or b);
    layer0_outputs(5798) <= not a or b;
    layer0_outputs(5799) <= not (a xor b);
    layer0_outputs(5800) <= a;
    layer0_outputs(5801) <= not a or b;
    layer0_outputs(5802) <= a or b;
    layer0_outputs(5803) <= a;
    layer0_outputs(5804) <= a or b;
    layer0_outputs(5805) <= not (a or b);
    layer0_outputs(5806) <= a and not b;
    layer0_outputs(5807) <= a and not b;
    layer0_outputs(5808) <= not (a or b);
    layer0_outputs(5809) <= not (a or b);
    layer0_outputs(5810) <= a or b;
    layer0_outputs(5811) <= a;
    layer0_outputs(5812) <= a and b;
    layer0_outputs(5813) <= not (a or b);
    layer0_outputs(5814) <= not b;
    layer0_outputs(5815) <= a or b;
    layer0_outputs(5816) <= a or b;
    layer0_outputs(5817) <= a or b;
    layer0_outputs(5818) <= not b;
    layer0_outputs(5819) <= not (a or b);
    layer0_outputs(5820) <= a or b;
    layer0_outputs(5821) <= b and not a;
    layer0_outputs(5822) <= a or b;
    layer0_outputs(5823) <= not b or a;
    layer0_outputs(5824) <= not b;
    layer0_outputs(5825) <= b and not a;
    layer0_outputs(5826) <= a xor b;
    layer0_outputs(5827) <= a xor b;
    layer0_outputs(5828) <= not (a or b);
    layer0_outputs(5829) <= a;
    layer0_outputs(5830) <= not (a xor b);
    layer0_outputs(5831) <= a xor b;
    layer0_outputs(5832) <= not (a xor b);
    layer0_outputs(5833) <= b;
    layer0_outputs(5834) <= a xor b;
    layer0_outputs(5835) <= not b;
    layer0_outputs(5836) <= not (a xor b);
    layer0_outputs(5837) <= b and not a;
    layer0_outputs(5838) <= not (a or b);
    layer0_outputs(5839) <= b;
    layer0_outputs(5840) <= a or b;
    layer0_outputs(5841) <= not (a or b);
    layer0_outputs(5842) <= not b or a;
    layer0_outputs(5843) <= not b;
    layer0_outputs(5844) <= a;
    layer0_outputs(5845) <= b;
    layer0_outputs(5846) <= a xor b;
    layer0_outputs(5847) <= not (a xor b);
    layer0_outputs(5848) <= b and not a;
    layer0_outputs(5849) <= 1'b1;
    layer0_outputs(5850) <= a and not b;
    layer0_outputs(5851) <= not (a and b);
    layer0_outputs(5852) <= a;
    layer0_outputs(5853) <= not (a or b);
    layer0_outputs(5854) <= not (a and b);
    layer0_outputs(5855) <= 1'b1;
    layer0_outputs(5856) <= b;
    layer0_outputs(5857) <= not (a xor b);
    layer0_outputs(5858) <= not (a xor b);
    layer0_outputs(5859) <= not b;
    layer0_outputs(5860) <= not a;
    layer0_outputs(5861) <= not a;
    layer0_outputs(5862) <= not b or a;
    layer0_outputs(5863) <= 1'b1;
    layer0_outputs(5864) <= not (a and b);
    layer0_outputs(5865) <= not (a or b);
    layer0_outputs(5866) <= not b or a;
    layer0_outputs(5867) <= b and not a;
    layer0_outputs(5868) <= a or b;
    layer0_outputs(5869) <= a;
    layer0_outputs(5870) <= b;
    layer0_outputs(5871) <= not a or b;
    layer0_outputs(5872) <= not (a xor b);
    layer0_outputs(5873) <= not (a xor b);
    layer0_outputs(5874) <= not b;
    layer0_outputs(5875) <= not a or b;
    layer0_outputs(5876) <= a or b;
    layer0_outputs(5877) <= not (a or b);
    layer0_outputs(5878) <= b;
    layer0_outputs(5879) <= not a;
    layer0_outputs(5880) <= a or b;
    layer0_outputs(5881) <= a xor b;
    layer0_outputs(5882) <= not a;
    layer0_outputs(5883) <= a or b;
    layer0_outputs(5884) <= not (a or b);
    layer0_outputs(5885) <= a or b;
    layer0_outputs(5886) <= not b;
    layer0_outputs(5887) <= a;
    layer0_outputs(5888) <= not (a xor b);
    layer0_outputs(5889) <= b;
    layer0_outputs(5890) <= a xor b;
    layer0_outputs(5891) <= not b or a;
    layer0_outputs(5892) <= not b;
    layer0_outputs(5893) <= a or b;
    layer0_outputs(5894) <= not a or b;
    layer0_outputs(5895) <= b;
    layer0_outputs(5896) <= 1'b1;
    layer0_outputs(5897) <= not a;
    layer0_outputs(5898) <= 1'b1;
    layer0_outputs(5899) <= not b or a;
    layer0_outputs(5900) <= 1'b0;
    layer0_outputs(5901) <= a;
    layer0_outputs(5902) <= a and not b;
    layer0_outputs(5903) <= not (a and b);
    layer0_outputs(5904) <= not b or a;
    layer0_outputs(5905) <= a;
    layer0_outputs(5906) <= b and not a;
    layer0_outputs(5907) <= a xor b;
    layer0_outputs(5908) <= not b or a;
    layer0_outputs(5909) <= a;
    layer0_outputs(5910) <= not (a xor b);
    layer0_outputs(5911) <= not (a xor b);
    layer0_outputs(5912) <= a or b;
    layer0_outputs(5913) <= not (a or b);
    layer0_outputs(5914) <= 1'b1;
    layer0_outputs(5915) <= not (a and b);
    layer0_outputs(5916) <= a xor b;
    layer0_outputs(5917) <= not (a xor b);
    layer0_outputs(5918) <= not (a xor b);
    layer0_outputs(5919) <= b;
    layer0_outputs(5920) <= not b;
    layer0_outputs(5921) <= a xor b;
    layer0_outputs(5922) <= b;
    layer0_outputs(5923) <= a and not b;
    layer0_outputs(5924) <= b and not a;
    layer0_outputs(5925) <= a xor b;
    layer0_outputs(5926) <= a;
    layer0_outputs(5927) <= a and not b;
    layer0_outputs(5928) <= not b or a;
    layer0_outputs(5929) <= not b or a;
    layer0_outputs(5930) <= a;
    layer0_outputs(5931) <= b;
    layer0_outputs(5932) <= a xor b;
    layer0_outputs(5933) <= not (a or b);
    layer0_outputs(5934) <= not a or b;
    layer0_outputs(5935) <= not (a or b);
    layer0_outputs(5936) <= not (a xor b);
    layer0_outputs(5937) <= not (a xor b);
    layer0_outputs(5938) <= a xor b;
    layer0_outputs(5939) <= not (a xor b);
    layer0_outputs(5940) <= not (a or b);
    layer0_outputs(5941) <= a xor b;
    layer0_outputs(5942) <= a xor b;
    layer0_outputs(5943) <= a xor b;
    layer0_outputs(5944) <= not a;
    layer0_outputs(5945) <= a and not b;
    layer0_outputs(5946) <= not b or a;
    layer0_outputs(5947) <= not (a or b);
    layer0_outputs(5948) <= not (a xor b);
    layer0_outputs(5949) <= not (a xor b);
    layer0_outputs(5950) <= not (a or b);
    layer0_outputs(5951) <= a;
    layer0_outputs(5952) <= not (a xor b);
    layer0_outputs(5953) <= 1'b0;
    layer0_outputs(5954) <= a;
    layer0_outputs(5955) <= 1'b0;
    layer0_outputs(5956) <= a or b;
    layer0_outputs(5957) <= a or b;
    layer0_outputs(5958) <= b;
    layer0_outputs(5959) <= a and not b;
    layer0_outputs(5960) <= not b;
    layer0_outputs(5961) <= not b;
    layer0_outputs(5962) <= not (a or b);
    layer0_outputs(5963) <= not (a or b);
    layer0_outputs(5964) <= not (a or b);
    layer0_outputs(5965) <= a or b;
    layer0_outputs(5966) <= not a or b;
    layer0_outputs(5967) <= not a or b;
    layer0_outputs(5968) <= not (a xor b);
    layer0_outputs(5969) <= a xor b;
    layer0_outputs(5970) <= not (a xor b);
    layer0_outputs(5971) <= b and not a;
    layer0_outputs(5972) <= not a or b;
    layer0_outputs(5973) <= not (a or b);
    layer0_outputs(5974) <= not b;
    layer0_outputs(5975) <= not (a xor b);
    layer0_outputs(5976) <= a or b;
    layer0_outputs(5977) <= not (a or b);
    layer0_outputs(5978) <= a;
    layer0_outputs(5979) <= not (a or b);
    layer0_outputs(5980) <= not (a or b);
    layer0_outputs(5981) <= a or b;
    layer0_outputs(5982) <= a;
    layer0_outputs(5983) <= a or b;
    layer0_outputs(5984) <= not (a or b);
    layer0_outputs(5985) <= not a;
    layer0_outputs(5986) <= not (a xor b);
    layer0_outputs(5987) <= not (a or b);
    layer0_outputs(5988) <= not (a and b);
    layer0_outputs(5989) <= a or b;
    layer0_outputs(5990) <= not (a or b);
    layer0_outputs(5991) <= a and b;
    layer0_outputs(5992) <= b and not a;
    layer0_outputs(5993) <= not (a or b);
    layer0_outputs(5994) <= a xor b;
    layer0_outputs(5995) <= b;
    layer0_outputs(5996) <= 1'b1;
    layer0_outputs(5997) <= not b or a;
    layer0_outputs(5998) <= not b or a;
    layer0_outputs(5999) <= a xor b;
    layer0_outputs(6000) <= not (a or b);
    layer0_outputs(6001) <= 1'b0;
    layer0_outputs(6002) <= a or b;
    layer0_outputs(6003) <= b and not a;
    layer0_outputs(6004) <= b and not a;
    layer0_outputs(6005) <= a or b;
    layer0_outputs(6006) <= a;
    layer0_outputs(6007) <= not b or a;
    layer0_outputs(6008) <= not b;
    layer0_outputs(6009) <= 1'b0;
    layer0_outputs(6010) <= b and not a;
    layer0_outputs(6011) <= not a;
    layer0_outputs(6012) <= not (a or b);
    layer0_outputs(6013) <= not a or b;
    layer0_outputs(6014) <= not a or b;
    layer0_outputs(6015) <= a and not b;
    layer0_outputs(6016) <= not (a and b);
    layer0_outputs(6017) <= 1'b1;
    layer0_outputs(6018) <= not b;
    layer0_outputs(6019) <= not a or b;
    layer0_outputs(6020) <= a;
    layer0_outputs(6021) <= not a;
    layer0_outputs(6022) <= not (a or b);
    layer0_outputs(6023) <= not b or a;
    layer0_outputs(6024) <= a and not b;
    layer0_outputs(6025) <= b;
    layer0_outputs(6026) <= b and not a;
    layer0_outputs(6027) <= not b or a;
    layer0_outputs(6028) <= not (a or b);
    layer0_outputs(6029) <= b and not a;
    layer0_outputs(6030) <= not a or b;
    layer0_outputs(6031) <= a or b;
    layer0_outputs(6032) <= not b or a;
    layer0_outputs(6033) <= not (a xor b);
    layer0_outputs(6034) <= not (a and b);
    layer0_outputs(6035) <= b;
    layer0_outputs(6036) <= not b or a;
    layer0_outputs(6037) <= not a or b;
    layer0_outputs(6038) <= b and not a;
    layer0_outputs(6039) <= a xor b;
    layer0_outputs(6040) <= b and not a;
    layer0_outputs(6041) <= not b or a;
    layer0_outputs(6042) <= a and not b;
    layer0_outputs(6043) <= a xor b;
    layer0_outputs(6044) <= not (a or b);
    layer0_outputs(6045) <= not b;
    layer0_outputs(6046) <= a or b;
    layer0_outputs(6047) <= a;
    layer0_outputs(6048) <= b;
    layer0_outputs(6049) <= a;
    layer0_outputs(6050) <= not (a or b);
    layer0_outputs(6051) <= not b;
    layer0_outputs(6052) <= b and not a;
    layer0_outputs(6053) <= a or b;
    layer0_outputs(6054) <= not b;
    layer0_outputs(6055) <= a or b;
    layer0_outputs(6056) <= b and not a;
    layer0_outputs(6057) <= a and not b;
    layer0_outputs(6058) <= a or b;
    layer0_outputs(6059) <= a or b;
    layer0_outputs(6060) <= a or b;
    layer0_outputs(6061) <= not (a xor b);
    layer0_outputs(6062) <= a or b;
    layer0_outputs(6063) <= 1'b0;
    layer0_outputs(6064) <= a xor b;
    layer0_outputs(6065) <= a or b;
    layer0_outputs(6066) <= b and not a;
    layer0_outputs(6067) <= b;
    layer0_outputs(6068) <= not b or a;
    layer0_outputs(6069) <= a or b;
    layer0_outputs(6070) <= not a;
    layer0_outputs(6071) <= not (a or b);
    layer0_outputs(6072) <= b;
    layer0_outputs(6073) <= not b or a;
    layer0_outputs(6074) <= not b or a;
    layer0_outputs(6075) <= a xor b;
    layer0_outputs(6076) <= b and not a;
    layer0_outputs(6077) <= not a or b;
    layer0_outputs(6078) <= a;
    layer0_outputs(6079) <= a or b;
    layer0_outputs(6080) <= not a or b;
    layer0_outputs(6081) <= not (a xor b);
    layer0_outputs(6082) <= not (a xor b);
    layer0_outputs(6083) <= b and not a;
    layer0_outputs(6084) <= a or b;
    layer0_outputs(6085) <= a;
    layer0_outputs(6086) <= not b;
    layer0_outputs(6087) <= not (a xor b);
    layer0_outputs(6088) <= not (a or b);
    layer0_outputs(6089) <= a xor b;
    layer0_outputs(6090) <= a or b;
    layer0_outputs(6091) <= a xor b;
    layer0_outputs(6092) <= b and not a;
    layer0_outputs(6093) <= b;
    layer0_outputs(6094) <= not b;
    layer0_outputs(6095) <= a and not b;
    layer0_outputs(6096) <= a;
    layer0_outputs(6097) <= b and not a;
    layer0_outputs(6098) <= a;
    layer0_outputs(6099) <= a or b;
    layer0_outputs(6100) <= a;
    layer0_outputs(6101) <= not (a xor b);
    layer0_outputs(6102) <= not a;
    layer0_outputs(6103) <= not a;
    layer0_outputs(6104) <= a and not b;
    layer0_outputs(6105) <= b and not a;
    layer0_outputs(6106) <= a and b;
    layer0_outputs(6107) <= a or b;
    layer0_outputs(6108) <= 1'b1;
    layer0_outputs(6109) <= not b or a;
    layer0_outputs(6110) <= b and not a;
    layer0_outputs(6111) <= not a or b;
    layer0_outputs(6112) <= b;
    layer0_outputs(6113) <= b and not a;
    layer0_outputs(6114) <= a;
    layer0_outputs(6115) <= a or b;
    layer0_outputs(6116) <= a or b;
    layer0_outputs(6117) <= not a or b;
    layer0_outputs(6118) <= not (a or b);
    layer0_outputs(6119) <= not a;
    layer0_outputs(6120) <= a xor b;
    layer0_outputs(6121) <= a or b;
    layer0_outputs(6122) <= not (a or b);
    layer0_outputs(6123) <= not (a xor b);
    layer0_outputs(6124) <= not b;
    layer0_outputs(6125) <= not (a or b);
    layer0_outputs(6126) <= not b or a;
    layer0_outputs(6127) <= not b;
    layer0_outputs(6128) <= not (a or b);
    layer0_outputs(6129) <= not (a or b);
    layer0_outputs(6130) <= 1'b0;
    layer0_outputs(6131) <= a or b;
    layer0_outputs(6132) <= a and b;
    layer0_outputs(6133) <= a or b;
    layer0_outputs(6134) <= not (a xor b);
    layer0_outputs(6135) <= a and b;
    layer0_outputs(6136) <= a or b;
    layer0_outputs(6137) <= 1'b1;
    layer0_outputs(6138) <= a or b;
    layer0_outputs(6139) <= b;
    layer0_outputs(6140) <= not a;
    layer0_outputs(6141) <= not b;
    layer0_outputs(6142) <= not b or a;
    layer0_outputs(6143) <= a xor b;
    layer0_outputs(6144) <= 1'b0;
    layer0_outputs(6145) <= not a or b;
    layer0_outputs(6146) <= a or b;
    layer0_outputs(6147) <= a xor b;
    layer0_outputs(6148) <= not a;
    layer0_outputs(6149) <= b and not a;
    layer0_outputs(6150) <= a;
    layer0_outputs(6151) <= a xor b;
    layer0_outputs(6152) <= not a;
    layer0_outputs(6153) <= 1'b1;
    layer0_outputs(6154) <= b and not a;
    layer0_outputs(6155) <= not (a or b);
    layer0_outputs(6156) <= b;
    layer0_outputs(6157) <= not b or a;
    layer0_outputs(6158) <= not (a or b);
    layer0_outputs(6159) <= not b;
    layer0_outputs(6160) <= b and not a;
    layer0_outputs(6161) <= not (a or b);
    layer0_outputs(6162) <= not (a or b);
    layer0_outputs(6163) <= not a;
    layer0_outputs(6164) <= not a;
    layer0_outputs(6165) <= not a or b;
    layer0_outputs(6166) <= not a;
    layer0_outputs(6167) <= not (a or b);
    layer0_outputs(6168) <= 1'b0;
    layer0_outputs(6169) <= a xor b;
    layer0_outputs(6170) <= a or b;
    layer0_outputs(6171) <= b and not a;
    layer0_outputs(6172) <= not (a xor b);
    layer0_outputs(6173) <= not a;
    layer0_outputs(6174) <= a and b;
    layer0_outputs(6175) <= b;
    layer0_outputs(6176) <= not (a or b);
    layer0_outputs(6177) <= not (a or b);
    layer0_outputs(6178) <= not b or a;
    layer0_outputs(6179) <= a or b;
    layer0_outputs(6180) <= a or b;
    layer0_outputs(6181) <= a or b;
    layer0_outputs(6182) <= a or b;
    layer0_outputs(6183) <= not a;
    layer0_outputs(6184) <= b and not a;
    layer0_outputs(6185) <= not a or b;
    layer0_outputs(6186) <= a or b;
    layer0_outputs(6187) <= b and not a;
    layer0_outputs(6188) <= not b;
    layer0_outputs(6189) <= not a;
    layer0_outputs(6190) <= a xor b;
    layer0_outputs(6191) <= not (a or b);
    layer0_outputs(6192) <= not b;
    layer0_outputs(6193) <= a;
    layer0_outputs(6194) <= not a or b;
    layer0_outputs(6195) <= not b;
    layer0_outputs(6196) <= a or b;
    layer0_outputs(6197) <= not b;
    layer0_outputs(6198) <= not b;
    layer0_outputs(6199) <= not (a xor b);
    layer0_outputs(6200) <= not a or b;
    layer0_outputs(6201) <= not (a or b);
    layer0_outputs(6202) <= a;
    layer0_outputs(6203) <= a or b;
    layer0_outputs(6204) <= a and not b;
    layer0_outputs(6205) <= a and not b;
    layer0_outputs(6206) <= a or b;
    layer0_outputs(6207) <= a xor b;
    layer0_outputs(6208) <= not a or b;
    layer0_outputs(6209) <= b and not a;
    layer0_outputs(6210) <= not (a xor b);
    layer0_outputs(6211) <= 1'b0;
    layer0_outputs(6212) <= a or b;
    layer0_outputs(6213) <= 1'b0;
    layer0_outputs(6214) <= not b;
    layer0_outputs(6215) <= a or b;
    layer0_outputs(6216) <= not b or a;
    layer0_outputs(6217) <= b and not a;
    layer0_outputs(6218) <= not (a xor b);
    layer0_outputs(6219) <= not (a or b);
    layer0_outputs(6220) <= a xor b;
    layer0_outputs(6221) <= a and not b;
    layer0_outputs(6222) <= not a;
    layer0_outputs(6223) <= a and b;
    layer0_outputs(6224) <= not (a xor b);
    layer0_outputs(6225) <= not b;
    layer0_outputs(6226) <= a xor b;
    layer0_outputs(6227) <= not (a xor b);
    layer0_outputs(6228) <= not (a or b);
    layer0_outputs(6229) <= not (a or b);
    layer0_outputs(6230) <= b and not a;
    layer0_outputs(6231) <= a and b;
    layer0_outputs(6232) <= 1'b1;
    layer0_outputs(6233) <= a and not b;
    layer0_outputs(6234) <= not b;
    layer0_outputs(6235) <= not a or b;
    layer0_outputs(6236) <= not (a xor b);
    layer0_outputs(6237) <= 1'b1;
    layer0_outputs(6238) <= a;
    layer0_outputs(6239) <= not b or a;
    layer0_outputs(6240) <= a xor b;
    layer0_outputs(6241) <= a;
    layer0_outputs(6242) <= 1'b0;
    layer0_outputs(6243) <= not (a or b);
    layer0_outputs(6244) <= b and not a;
    layer0_outputs(6245) <= not a or b;
    layer0_outputs(6246) <= a and not b;
    layer0_outputs(6247) <= not a;
    layer0_outputs(6248) <= a and b;
    layer0_outputs(6249) <= a or b;
    layer0_outputs(6250) <= a or b;
    layer0_outputs(6251) <= a xor b;
    layer0_outputs(6252) <= not a;
    layer0_outputs(6253) <= not (a xor b);
    layer0_outputs(6254) <= not b;
    layer0_outputs(6255) <= not (a xor b);
    layer0_outputs(6256) <= a;
    layer0_outputs(6257) <= not b;
    layer0_outputs(6258) <= not (a or b);
    layer0_outputs(6259) <= a or b;
    layer0_outputs(6260) <= b and not a;
    layer0_outputs(6261) <= a and not b;
    layer0_outputs(6262) <= a;
    layer0_outputs(6263) <= not b or a;
    layer0_outputs(6264) <= not b or a;
    layer0_outputs(6265) <= not a;
    layer0_outputs(6266) <= not b or a;
    layer0_outputs(6267) <= a;
    layer0_outputs(6268) <= not b;
    layer0_outputs(6269) <= b;
    layer0_outputs(6270) <= not a;
    layer0_outputs(6271) <= not b or a;
    layer0_outputs(6272) <= not a or b;
    layer0_outputs(6273) <= not a or b;
    layer0_outputs(6274) <= a xor b;
    layer0_outputs(6275) <= not (a or b);
    layer0_outputs(6276) <= not b;
    layer0_outputs(6277) <= not a;
    layer0_outputs(6278) <= not (a xor b);
    layer0_outputs(6279) <= b;
    layer0_outputs(6280) <= not (a or b);
    layer0_outputs(6281) <= 1'b0;
    layer0_outputs(6282) <= not a;
    layer0_outputs(6283) <= not b or a;
    layer0_outputs(6284) <= not b;
    layer0_outputs(6285) <= b and not a;
    layer0_outputs(6286) <= a xor b;
    layer0_outputs(6287) <= a xor b;
    layer0_outputs(6288) <= a or b;
    layer0_outputs(6289) <= b;
    layer0_outputs(6290) <= b;
    layer0_outputs(6291) <= b and not a;
    layer0_outputs(6292) <= a xor b;
    layer0_outputs(6293) <= not a or b;
    layer0_outputs(6294) <= not a or b;
    layer0_outputs(6295) <= not b;
    layer0_outputs(6296) <= a or b;
    layer0_outputs(6297) <= a and not b;
    layer0_outputs(6298) <= a and not b;
    layer0_outputs(6299) <= a xor b;
    layer0_outputs(6300) <= a or b;
    layer0_outputs(6301) <= b and not a;
    layer0_outputs(6302) <= a or b;
    layer0_outputs(6303) <= b and not a;
    layer0_outputs(6304) <= b;
    layer0_outputs(6305) <= a or b;
    layer0_outputs(6306) <= not b or a;
    layer0_outputs(6307) <= a xor b;
    layer0_outputs(6308) <= not (a xor b);
    layer0_outputs(6309) <= not a or b;
    layer0_outputs(6310) <= 1'b1;
    layer0_outputs(6311) <= a or b;
    layer0_outputs(6312) <= a or b;
    layer0_outputs(6313) <= not b or a;
    layer0_outputs(6314) <= b;
    layer0_outputs(6315) <= not a;
    layer0_outputs(6316) <= not (a xor b);
    layer0_outputs(6317) <= a xor b;
    layer0_outputs(6318) <= a xor b;
    layer0_outputs(6319) <= a and not b;
    layer0_outputs(6320) <= a or b;
    layer0_outputs(6321) <= a or b;
    layer0_outputs(6322) <= not (a or b);
    layer0_outputs(6323) <= not (a xor b);
    layer0_outputs(6324) <= not (a or b);
    layer0_outputs(6325) <= not (a or b);
    layer0_outputs(6326) <= not (a and b);
    layer0_outputs(6327) <= a or b;
    layer0_outputs(6328) <= not (a or b);
    layer0_outputs(6329) <= not a;
    layer0_outputs(6330) <= a xor b;
    layer0_outputs(6331) <= a;
    layer0_outputs(6332) <= a or b;
    layer0_outputs(6333) <= not b;
    layer0_outputs(6334) <= 1'b0;
    layer0_outputs(6335) <= a xor b;
    layer0_outputs(6336) <= 1'b1;
    layer0_outputs(6337) <= not a or b;
    layer0_outputs(6338) <= not b;
    layer0_outputs(6339) <= a and b;
    layer0_outputs(6340) <= not (a xor b);
    layer0_outputs(6341) <= a or b;
    layer0_outputs(6342) <= not (a and b);
    layer0_outputs(6343) <= a and not b;
    layer0_outputs(6344) <= a and not b;
    layer0_outputs(6345) <= b and not a;
    layer0_outputs(6346) <= not b;
    layer0_outputs(6347) <= not (a or b);
    layer0_outputs(6348) <= a and b;
    layer0_outputs(6349) <= a xor b;
    layer0_outputs(6350) <= not b;
    layer0_outputs(6351) <= a;
    layer0_outputs(6352) <= not b or a;
    layer0_outputs(6353) <= a xor b;
    layer0_outputs(6354) <= not (a or b);
    layer0_outputs(6355) <= not (a or b);
    layer0_outputs(6356) <= a or b;
    layer0_outputs(6357) <= a and b;
    layer0_outputs(6358) <= not (a or b);
    layer0_outputs(6359) <= b;
    layer0_outputs(6360) <= not (a or b);
    layer0_outputs(6361) <= a xor b;
    layer0_outputs(6362) <= not a or b;
    layer0_outputs(6363) <= a or b;
    layer0_outputs(6364) <= not b or a;
    layer0_outputs(6365) <= 1'b0;
    layer0_outputs(6366) <= a xor b;
    layer0_outputs(6367) <= not (a or b);
    layer0_outputs(6368) <= not a or b;
    layer0_outputs(6369) <= not (a or b);
    layer0_outputs(6370) <= b;
    layer0_outputs(6371) <= a;
    layer0_outputs(6372) <= not a or b;
    layer0_outputs(6373) <= a;
    layer0_outputs(6374) <= not a or b;
    layer0_outputs(6375) <= b and not a;
    layer0_outputs(6376) <= b and not a;
    layer0_outputs(6377) <= a and not b;
    layer0_outputs(6378) <= a or b;
    layer0_outputs(6379) <= b;
    layer0_outputs(6380) <= not b;
    layer0_outputs(6381) <= a xor b;
    layer0_outputs(6382) <= a and not b;
    layer0_outputs(6383) <= a or b;
    layer0_outputs(6384) <= a xor b;
    layer0_outputs(6385) <= a and not b;
    layer0_outputs(6386) <= b;
    layer0_outputs(6387) <= b;
    layer0_outputs(6388) <= a and not b;
    layer0_outputs(6389) <= not (a xor b);
    layer0_outputs(6390) <= not a;
    layer0_outputs(6391) <= not a or b;
    layer0_outputs(6392) <= not (a or b);
    layer0_outputs(6393) <= a;
    layer0_outputs(6394) <= not (a or b);
    layer0_outputs(6395) <= not b or a;
    layer0_outputs(6396) <= not a or b;
    layer0_outputs(6397) <= a or b;
    layer0_outputs(6398) <= not a or b;
    layer0_outputs(6399) <= not (a or b);
    layer0_outputs(6400) <= not a;
    layer0_outputs(6401) <= not b;
    layer0_outputs(6402) <= not b;
    layer0_outputs(6403) <= a;
    layer0_outputs(6404) <= b and not a;
    layer0_outputs(6405) <= a and not b;
    layer0_outputs(6406) <= a;
    layer0_outputs(6407) <= not b or a;
    layer0_outputs(6408) <= not (a and b);
    layer0_outputs(6409) <= not (a or b);
    layer0_outputs(6410) <= not a;
    layer0_outputs(6411) <= not a or b;
    layer0_outputs(6412) <= a or b;
    layer0_outputs(6413) <= a or b;
    layer0_outputs(6414) <= not (a xor b);
    layer0_outputs(6415) <= b;
    layer0_outputs(6416) <= a xor b;
    layer0_outputs(6417) <= b;
    layer0_outputs(6418) <= not a or b;
    layer0_outputs(6419) <= not b or a;
    layer0_outputs(6420) <= not b;
    layer0_outputs(6421) <= a;
    layer0_outputs(6422) <= a and not b;
    layer0_outputs(6423) <= a and not b;
    layer0_outputs(6424) <= 1'b1;
    layer0_outputs(6425) <= a and not b;
    layer0_outputs(6426) <= not b;
    layer0_outputs(6427) <= not a;
    layer0_outputs(6428) <= a;
    layer0_outputs(6429) <= not b or a;
    layer0_outputs(6430) <= a or b;
    layer0_outputs(6431) <= a;
    layer0_outputs(6432) <= a xor b;
    layer0_outputs(6433) <= not (a or b);
    layer0_outputs(6434) <= a or b;
    layer0_outputs(6435) <= not (a or b);
    layer0_outputs(6436) <= not a;
    layer0_outputs(6437) <= not (a xor b);
    layer0_outputs(6438) <= not b or a;
    layer0_outputs(6439) <= a or b;
    layer0_outputs(6440) <= not a or b;
    layer0_outputs(6441) <= 1'b0;
    layer0_outputs(6442) <= a or b;
    layer0_outputs(6443) <= 1'b1;
    layer0_outputs(6444) <= not (a xor b);
    layer0_outputs(6445) <= 1'b1;
    layer0_outputs(6446) <= not (a or b);
    layer0_outputs(6447) <= not (a or b);
    layer0_outputs(6448) <= a or b;
    layer0_outputs(6449) <= not (a or b);
    layer0_outputs(6450) <= not (a and b);
    layer0_outputs(6451) <= not (a xor b);
    layer0_outputs(6452) <= not (a or b);
    layer0_outputs(6453) <= not (a and b);
    layer0_outputs(6454) <= b;
    layer0_outputs(6455) <= a xor b;
    layer0_outputs(6456) <= not b or a;
    layer0_outputs(6457) <= not a or b;
    layer0_outputs(6458) <= a xor b;
    layer0_outputs(6459) <= not a or b;
    layer0_outputs(6460) <= a or b;
    layer0_outputs(6461) <= 1'b0;
    layer0_outputs(6462) <= a xor b;
    layer0_outputs(6463) <= not (a or b);
    layer0_outputs(6464) <= a or b;
    layer0_outputs(6465) <= not a;
    layer0_outputs(6466) <= not a or b;
    layer0_outputs(6467) <= a;
    layer0_outputs(6468) <= a;
    layer0_outputs(6469) <= b;
    layer0_outputs(6470) <= a xor b;
    layer0_outputs(6471) <= not a;
    layer0_outputs(6472) <= not (a or b);
    layer0_outputs(6473) <= a or b;
    layer0_outputs(6474) <= not (a xor b);
    layer0_outputs(6475) <= a;
    layer0_outputs(6476) <= not (a or b);
    layer0_outputs(6477) <= b and not a;
    layer0_outputs(6478) <= a xor b;
    layer0_outputs(6479) <= not (a or b);
    layer0_outputs(6480) <= not (a xor b);
    layer0_outputs(6481) <= not (a or b);
    layer0_outputs(6482) <= not (a xor b);
    layer0_outputs(6483) <= a or b;
    layer0_outputs(6484) <= a and not b;
    layer0_outputs(6485) <= not b;
    layer0_outputs(6486) <= not (a xor b);
    layer0_outputs(6487) <= a and not b;
    layer0_outputs(6488) <= not b or a;
    layer0_outputs(6489) <= a xor b;
    layer0_outputs(6490) <= a xor b;
    layer0_outputs(6491) <= not (a or b);
    layer0_outputs(6492) <= b and not a;
    layer0_outputs(6493) <= not (a or b);
    layer0_outputs(6494) <= not (a or b);
    layer0_outputs(6495) <= a or b;
    layer0_outputs(6496) <= a;
    layer0_outputs(6497) <= not a or b;
    layer0_outputs(6498) <= 1'b1;
    layer0_outputs(6499) <= a or b;
    layer0_outputs(6500) <= a and not b;
    layer0_outputs(6501) <= a and not b;
    layer0_outputs(6502) <= not a;
    layer0_outputs(6503) <= a and b;
    layer0_outputs(6504) <= a;
    layer0_outputs(6505) <= not (a xor b);
    layer0_outputs(6506) <= not (a xor b);
    layer0_outputs(6507) <= a and b;
    layer0_outputs(6508) <= a;
    layer0_outputs(6509) <= not b or a;
    layer0_outputs(6510) <= a xor b;
    layer0_outputs(6511) <= a;
    layer0_outputs(6512) <= b and not a;
    layer0_outputs(6513) <= not (a or b);
    layer0_outputs(6514) <= a or b;
    layer0_outputs(6515) <= a and not b;
    layer0_outputs(6516) <= not b or a;
    layer0_outputs(6517) <= b;
    layer0_outputs(6518) <= not a;
    layer0_outputs(6519) <= not (a or b);
    layer0_outputs(6520) <= a or b;
    layer0_outputs(6521) <= not (a or b);
    layer0_outputs(6522) <= a xor b;
    layer0_outputs(6523) <= a or b;
    layer0_outputs(6524) <= not a or b;
    layer0_outputs(6525) <= a;
    layer0_outputs(6526) <= not a or b;
    layer0_outputs(6527) <= not b;
    layer0_outputs(6528) <= not a;
    layer0_outputs(6529) <= b;
    layer0_outputs(6530) <= not (a xor b);
    layer0_outputs(6531) <= not b;
    layer0_outputs(6532) <= not b;
    layer0_outputs(6533) <= a xor b;
    layer0_outputs(6534) <= b;
    layer0_outputs(6535) <= a or b;
    layer0_outputs(6536) <= a xor b;
    layer0_outputs(6537) <= not b;
    layer0_outputs(6538) <= 1'b0;
    layer0_outputs(6539) <= a xor b;
    layer0_outputs(6540) <= a or b;
    layer0_outputs(6541) <= 1'b1;
    layer0_outputs(6542) <= a xor b;
    layer0_outputs(6543) <= b and not a;
    layer0_outputs(6544) <= not (a and b);
    layer0_outputs(6545) <= not b;
    layer0_outputs(6546) <= not (a xor b);
    layer0_outputs(6547) <= not (a or b);
    layer0_outputs(6548) <= b;
    layer0_outputs(6549) <= not a;
    layer0_outputs(6550) <= not b or a;
    layer0_outputs(6551) <= not b or a;
    layer0_outputs(6552) <= a;
    layer0_outputs(6553) <= a or b;
    layer0_outputs(6554) <= a or b;
    layer0_outputs(6555) <= a or b;
    layer0_outputs(6556) <= a and not b;
    layer0_outputs(6557) <= a;
    layer0_outputs(6558) <= not (a xor b);
    layer0_outputs(6559) <= not a;
    layer0_outputs(6560) <= not (a xor b);
    layer0_outputs(6561) <= not (a or b);
    layer0_outputs(6562) <= b;
    layer0_outputs(6563) <= a or b;
    layer0_outputs(6564) <= not a;
    layer0_outputs(6565) <= a or b;
    layer0_outputs(6566) <= b;
    layer0_outputs(6567) <= not (a xor b);
    layer0_outputs(6568) <= a xor b;
    layer0_outputs(6569) <= a or b;
    layer0_outputs(6570) <= 1'b0;
    layer0_outputs(6571) <= not (a xor b);
    layer0_outputs(6572) <= not a or b;
    layer0_outputs(6573) <= a and not b;
    layer0_outputs(6574) <= 1'b1;
    layer0_outputs(6575) <= not (a xor b);
    layer0_outputs(6576) <= b;
    layer0_outputs(6577) <= a and b;
    layer0_outputs(6578) <= a xor b;
    layer0_outputs(6579) <= not a or b;
    layer0_outputs(6580) <= a or b;
    layer0_outputs(6581) <= not (a or b);
    layer0_outputs(6582) <= b and not a;
    layer0_outputs(6583) <= not a;
    layer0_outputs(6584) <= b and not a;
    layer0_outputs(6585) <= a or b;
    layer0_outputs(6586) <= not a or b;
    layer0_outputs(6587) <= a xor b;
    layer0_outputs(6588) <= not a or b;
    layer0_outputs(6589) <= not (a xor b);
    layer0_outputs(6590) <= not (a xor b);
    layer0_outputs(6591) <= b;
    layer0_outputs(6592) <= a xor b;
    layer0_outputs(6593) <= not (a or b);
    layer0_outputs(6594) <= not (a xor b);
    layer0_outputs(6595) <= a or b;
    layer0_outputs(6596) <= b;
    layer0_outputs(6597) <= not (a or b);
    layer0_outputs(6598) <= not (a xor b);
    layer0_outputs(6599) <= 1'b1;
    layer0_outputs(6600) <= a;
    layer0_outputs(6601) <= a xor b;
    layer0_outputs(6602) <= not b;
    layer0_outputs(6603) <= a or b;
    layer0_outputs(6604) <= not b;
    layer0_outputs(6605) <= b;
    layer0_outputs(6606) <= a and b;
    layer0_outputs(6607) <= a or b;
    layer0_outputs(6608) <= a and b;
    layer0_outputs(6609) <= not a or b;
    layer0_outputs(6610) <= not (a and b);
    layer0_outputs(6611) <= b;
    layer0_outputs(6612) <= not a;
    layer0_outputs(6613) <= a;
    layer0_outputs(6614) <= a xor b;
    layer0_outputs(6615) <= a;
    layer0_outputs(6616) <= not b;
    layer0_outputs(6617) <= a or b;
    layer0_outputs(6618) <= a xor b;
    layer0_outputs(6619) <= not (a xor b);
    layer0_outputs(6620) <= not a or b;
    layer0_outputs(6621) <= a or b;
    layer0_outputs(6622) <= a or b;
    layer0_outputs(6623) <= a and b;
    layer0_outputs(6624) <= b;
    layer0_outputs(6625) <= a or b;
    layer0_outputs(6626) <= b and not a;
    layer0_outputs(6627) <= not b or a;
    layer0_outputs(6628) <= not (a or b);
    layer0_outputs(6629) <= a or b;
    layer0_outputs(6630) <= a and not b;
    layer0_outputs(6631) <= b;
    layer0_outputs(6632) <= 1'b1;
    layer0_outputs(6633) <= a and not b;
    layer0_outputs(6634) <= not (a xor b);
    layer0_outputs(6635) <= not (a xor b);
    layer0_outputs(6636) <= a or b;
    layer0_outputs(6637) <= not (a xor b);
    layer0_outputs(6638) <= a;
    layer0_outputs(6639) <= not (a or b);
    layer0_outputs(6640) <= not b or a;
    layer0_outputs(6641) <= b;
    layer0_outputs(6642) <= a;
    layer0_outputs(6643) <= a;
    layer0_outputs(6644) <= not (a or b);
    layer0_outputs(6645) <= not b;
    layer0_outputs(6646) <= not a or b;
    layer0_outputs(6647) <= a or b;
    layer0_outputs(6648) <= a xor b;
    layer0_outputs(6649) <= 1'b1;
    layer0_outputs(6650) <= a or b;
    layer0_outputs(6651) <= a;
    layer0_outputs(6652) <= a xor b;
    layer0_outputs(6653) <= b;
    layer0_outputs(6654) <= not (a or b);
    layer0_outputs(6655) <= not (a or b);
    layer0_outputs(6656) <= not (a or b);
    layer0_outputs(6657) <= not b;
    layer0_outputs(6658) <= b;
    layer0_outputs(6659) <= not a or b;
    layer0_outputs(6660) <= a or b;
    layer0_outputs(6661) <= not (a xor b);
    layer0_outputs(6662) <= not a or b;
    layer0_outputs(6663) <= not a;
    layer0_outputs(6664) <= not (a xor b);
    layer0_outputs(6665) <= not a or b;
    layer0_outputs(6666) <= not (a xor b);
    layer0_outputs(6667) <= b;
    layer0_outputs(6668) <= not b or a;
    layer0_outputs(6669) <= a;
    layer0_outputs(6670) <= not b or a;
    layer0_outputs(6671) <= a or b;
    layer0_outputs(6672) <= not (a xor b);
    layer0_outputs(6673) <= a or b;
    layer0_outputs(6674) <= a and b;
    layer0_outputs(6675) <= a xor b;
    layer0_outputs(6676) <= not a;
    layer0_outputs(6677) <= b;
    layer0_outputs(6678) <= not b or a;
    layer0_outputs(6679) <= a or b;
    layer0_outputs(6680) <= not (a or b);
    layer0_outputs(6681) <= b and not a;
    layer0_outputs(6682) <= not a or b;
    layer0_outputs(6683) <= a xor b;
    layer0_outputs(6684) <= a or b;
    layer0_outputs(6685) <= a;
    layer0_outputs(6686) <= a or b;
    layer0_outputs(6687) <= a and not b;
    layer0_outputs(6688) <= not (a or b);
    layer0_outputs(6689) <= a or b;
    layer0_outputs(6690) <= not b;
    layer0_outputs(6691) <= not (a xor b);
    layer0_outputs(6692) <= not (a or b);
    layer0_outputs(6693) <= a and not b;
    layer0_outputs(6694) <= b;
    layer0_outputs(6695) <= not a or b;
    layer0_outputs(6696) <= not a or b;
    layer0_outputs(6697) <= a or b;
    layer0_outputs(6698) <= not a or b;
    layer0_outputs(6699) <= a and not b;
    layer0_outputs(6700) <= a and b;
    layer0_outputs(6701) <= a;
    layer0_outputs(6702) <= not (a or b);
    layer0_outputs(6703) <= not b or a;
    layer0_outputs(6704) <= not a;
    layer0_outputs(6705) <= b and not a;
    layer0_outputs(6706) <= a xor b;
    layer0_outputs(6707) <= a and not b;
    layer0_outputs(6708) <= a and not b;
    layer0_outputs(6709) <= a;
    layer0_outputs(6710) <= not a or b;
    layer0_outputs(6711) <= not (a or b);
    layer0_outputs(6712) <= 1'b0;
    layer0_outputs(6713) <= a or b;
    layer0_outputs(6714) <= not a;
    layer0_outputs(6715) <= 1'b0;
    layer0_outputs(6716) <= a and not b;
    layer0_outputs(6717) <= a and not b;
    layer0_outputs(6718) <= b and not a;
    layer0_outputs(6719) <= not b or a;
    layer0_outputs(6720) <= a and not b;
    layer0_outputs(6721) <= a or b;
    layer0_outputs(6722) <= not a;
    layer0_outputs(6723) <= not (a or b);
    layer0_outputs(6724) <= b;
    layer0_outputs(6725) <= not a or b;
    layer0_outputs(6726) <= a;
    layer0_outputs(6727) <= not a or b;
    layer0_outputs(6728) <= not b or a;
    layer0_outputs(6729) <= not b;
    layer0_outputs(6730) <= not (a or b);
    layer0_outputs(6731) <= not b or a;
    layer0_outputs(6732) <= a or b;
    layer0_outputs(6733) <= not (a xor b);
    layer0_outputs(6734) <= not (a or b);
    layer0_outputs(6735) <= b and not a;
    layer0_outputs(6736) <= b and not a;
    layer0_outputs(6737) <= not a;
    layer0_outputs(6738) <= a;
    layer0_outputs(6739) <= not (a or b);
    layer0_outputs(6740) <= a xor b;
    layer0_outputs(6741) <= a;
    layer0_outputs(6742) <= not (a or b);
    layer0_outputs(6743) <= not b or a;
    layer0_outputs(6744) <= not (a xor b);
    layer0_outputs(6745) <= a or b;
    layer0_outputs(6746) <= a xor b;
    layer0_outputs(6747) <= not a;
    layer0_outputs(6748) <= b;
    layer0_outputs(6749) <= a xor b;
    layer0_outputs(6750) <= not a;
    layer0_outputs(6751) <= not a or b;
    layer0_outputs(6752) <= not (a or b);
    layer0_outputs(6753) <= not b;
    layer0_outputs(6754) <= a xor b;
    layer0_outputs(6755) <= a or b;
    layer0_outputs(6756) <= not b;
    layer0_outputs(6757) <= not b;
    layer0_outputs(6758) <= a and not b;
    layer0_outputs(6759) <= not (a or b);
    layer0_outputs(6760) <= not (a xor b);
    layer0_outputs(6761) <= a xor b;
    layer0_outputs(6762) <= not (a xor b);
    layer0_outputs(6763) <= not a or b;
    layer0_outputs(6764) <= not b;
    layer0_outputs(6765) <= not (a xor b);
    layer0_outputs(6766) <= not b;
    layer0_outputs(6767) <= not (a or b);
    layer0_outputs(6768) <= a or b;
    layer0_outputs(6769) <= not a or b;
    layer0_outputs(6770) <= not a;
    layer0_outputs(6771) <= not a or b;
    layer0_outputs(6772) <= a and not b;
    layer0_outputs(6773) <= not b or a;
    layer0_outputs(6774) <= a or b;
    layer0_outputs(6775) <= b;
    layer0_outputs(6776) <= a or b;
    layer0_outputs(6777) <= a;
    layer0_outputs(6778) <= not b;
    layer0_outputs(6779) <= b and not a;
    layer0_outputs(6780) <= not (a or b);
    layer0_outputs(6781) <= a xor b;
    layer0_outputs(6782) <= not (a or b);
    layer0_outputs(6783) <= not (a or b);
    layer0_outputs(6784) <= not (a or b);
    layer0_outputs(6785) <= b;
    layer0_outputs(6786) <= a xor b;
    layer0_outputs(6787) <= not a or b;
    layer0_outputs(6788) <= not b;
    layer0_outputs(6789) <= not b or a;
    layer0_outputs(6790) <= a or b;
    layer0_outputs(6791) <= a xor b;
    layer0_outputs(6792) <= a;
    layer0_outputs(6793) <= not b;
    layer0_outputs(6794) <= not (a xor b);
    layer0_outputs(6795) <= b and not a;
    layer0_outputs(6796) <= b and not a;
    layer0_outputs(6797) <= not a or b;
    layer0_outputs(6798) <= a and b;
    layer0_outputs(6799) <= b and not a;
    layer0_outputs(6800) <= a or b;
    layer0_outputs(6801) <= a;
    layer0_outputs(6802) <= a and not b;
    layer0_outputs(6803) <= not (a xor b);
    layer0_outputs(6804) <= not b;
    layer0_outputs(6805) <= a or b;
    layer0_outputs(6806) <= not (a or b);
    layer0_outputs(6807) <= not (a or b);
    layer0_outputs(6808) <= not (a xor b);
    layer0_outputs(6809) <= not a or b;
    layer0_outputs(6810) <= not (a xor b);
    layer0_outputs(6811) <= not a or b;
    layer0_outputs(6812) <= a xor b;
    layer0_outputs(6813) <= not (a xor b);
    layer0_outputs(6814) <= not b or a;
    layer0_outputs(6815) <= not (a xor b);
    layer0_outputs(6816) <= a xor b;
    layer0_outputs(6817) <= a and not b;
    layer0_outputs(6818) <= a or b;
    layer0_outputs(6819) <= b;
    layer0_outputs(6820) <= not (a or b);
    layer0_outputs(6821) <= a or b;
    layer0_outputs(6822) <= not a;
    layer0_outputs(6823) <= not a or b;
    layer0_outputs(6824) <= not (a or b);
    layer0_outputs(6825) <= not b or a;
    layer0_outputs(6826) <= not b;
    layer0_outputs(6827) <= a and b;
    layer0_outputs(6828) <= a xor b;
    layer0_outputs(6829) <= not a or b;
    layer0_outputs(6830) <= a or b;
    layer0_outputs(6831) <= not (a or b);
    layer0_outputs(6832) <= a or b;
    layer0_outputs(6833) <= a;
    layer0_outputs(6834) <= b and not a;
    layer0_outputs(6835) <= not b or a;
    layer0_outputs(6836) <= not (a or b);
    layer0_outputs(6837) <= a or b;
    layer0_outputs(6838) <= not b or a;
    layer0_outputs(6839) <= not a or b;
    layer0_outputs(6840) <= a xor b;
    layer0_outputs(6841) <= not (a xor b);
    layer0_outputs(6842) <= not (a or b);
    layer0_outputs(6843) <= a and not b;
    layer0_outputs(6844) <= not (a xor b);
    layer0_outputs(6845) <= not (a or b);
    layer0_outputs(6846) <= a or b;
    layer0_outputs(6847) <= not (a xor b);
    layer0_outputs(6848) <= not (a or b);
    layer0_outputs(6849) <= a and not b;
    layer0_outputs(6850) <= not a;
    layer0_outputs(6851) <= a;
    layer0_outputs(6852) <= not b or a;
    layer0_outputs(6853) <= not a or b;
    layer0_outputs(6854) <= not (a or b);
    layer0_outputs(6855) <= a or b;
    layer0_outputs(6856) <= not b or a;
    layer0_outputs(6857) <= not (a or b);
    layer0_outputs(6858) <= 1'b1;
    layer0_outputs(6859) <= not b or a;
    layer0_outputs(6860) <= a and not b;
    layer0_outputs(6861) <= not (a or b);
    layer0_outputs(6862) <= a or b;
    layer0_outputs(6863) <= not (a or b);
    layer0_outputs(6864) <= a and not b;
    layer0_outputs(6865) <= not (a and b);
    layer0_outputs(6866) <= not (a xor b);
    layer0_outputs(6867) <= not b;
    layer0_outputs(6868) <= b;
    layer0_outputs(6869) <= a and not b;
    layer0_outputs(6870) <= not (a xor b);
    layer0_outputs(6871) <= a or b;
    layer0_outputs(6872) <= a and not b;
    layer0_outputs(6873) <= not b;
    layer0_outputs(6874) <= not b or a;
    layer0_outputs(6875) <= not (a and b);
    layer0_outputs(6876) <= not b or a;
    layer0_outputs(6877) <= not (a or b);
    layer0_outputs(6878) <= not a;
    layer0_outputs(6879) <= a and not b;
    layer0_outputs(6880) <= not (a or b);
    layer0_outputs(6881) <= a and not b;
    layer0_outputs(6882) <= not (a xor b);
    layer0_outputs(6883) <= a or b;
    layer0_outputs(6884) <= not (a or b);
    layer0_outputs(6885) <= b and not a;
    layer0_outputs(6886) <= not b or a;
    layer0_outputs(6887) <= not b or a;
    layer0_outputs(6888) <= a and not b;
    layer0_outputs(6889) <= not b;
    layer0_outputs(6890) <= a;
    layer0_outputs(6891) <= not a or b;
    layer0_outputs(6892) <= a or b;
    layer0_outputs(6893) <= a xor b;
    layer0_outputs(6894) <= b;
    layer0_outputs(6895) <= not b or a;
    layer0_outputs(6896) <= not b or a;
    layer0_outputs(6897) <= not a;
    layer0_outputs(6898) <= not b;
    layer0_outputs(6899) <= not (a xor b);
    layer0_outputs(6900) <= not (a or b);
    layer0_outputs(6901) <= b;
    layer0_outputs(6902) <= not (a xor b);
    layer0_outputs(6903) <= a;
    layer0_outputs(6904) <= a and not b;
    layer0_outputs(6905) <= a xor b;
    layer0_outputs(6906) <= a or b;
    layer0_outputs(6907) <= not a;
    layer0_outputs(6908) <= a or b;
    layer0_outputs(6909) <= b;
    layer0_outputs(6910) <= a;
    layer0_outputs(6911) <= a and not b;
    layer0_outputs(6912) <= not a or b;
    layer0_outputs(6913) <= a;
    layer0_outputs(6914) <= not a or b;
    layer0_outputs(6915) <= not b or a;
    layer0_outputs(6916) <= a xor b;
    layer0_outputs(6917) <= b;
    layer0_outputs(6918) <= not a;
    layer0_outputs(6919) <= not a;
    layer0_outputs(6920) <= a or b;
    layer0_outputs(6921) <= not a or b;
    layer0_outputs(6922) <= a or b;
    layer0_outputs(6923) <= a or b;
    layer0_outputs(6924) <= not a;
    layer0_outputs(6925) <= a;
    layer0_outputs(6926) <= not (a or b);
    layer0_outputs(6927) <= not b;
    layer0_outputs(6928) <= not a or b;
    layer0_outputs(6929) <= not (a xor b);
    layer0_outputs(6930) <= not b;
    layer0_outputs(6931) <= not (a or b);
    layer0_outputs(6932) <= not a or b;
    layer0_outputs(6933) <= a xor b;
    layer0_outputs(6934) <= not a;
    layer0_outputs(6935) <= a or b;
    layer0_outputs(6936) <= not (a or b);
    layer0_outputs(6937) <= b;
    layer0_outputs(6938) <= b;
    layer0_outputs(6939) <= b;
    layer0_outputs(6940) <= not (a or b);
    layer0_outputs(6941) <= a xor b;
    layer0_outputs(6942) <= not a or b;
    layer0_outputs(6943) <= not b or a;
    layer0_outputs(6944) <= not (a or b);
    layer0_outputs(6945) <= 1'b1;
    layer0_outputs(6946) <= a xor b;
    layer0_outputs(6947) <= not (a or b);
    layer0_outputs(6948) <= not (a or b);
    layer0_outputs(6949) <= b and not a;
    layer0_outputs(6950) <= a xor b;
    layer0_outputs(6951) <= 1'b1;
    layer0_outputs(6952) <= not a;
    layer0_outputs(6953) <= b;
    layer0_outputs(6954) <= a;
    layer0_outputs(6955) <= b;
    layer0_outputs(6956) <= 1'b0;
    layer0_outputs(6957) <= not (a or b);
    layer0_outputs(6958) <= not b or a;
    layer0_outputs(6959) <= b;
    layer0_outputs(6960) <= not b or a;
    layer0_outputs(6961) <= a;
    layer0_outputs(6962) <= a;
    layer0_outputs(6963) <= not (a or b);
    layer0_outputs(6964) <= a or b;
    layer0_outputs(6965) <= b and not a;
    layer0_outputs(6966) <= a and not b;
    layer0_outputs(6967) <= a or b;
    layer0_outputs(6968) <= a and b;
    layer0_outputs(6969) <= a;
    layer0_outputs(6970) <= not (a or b);
    layer0_outputs(6971) <= not (a or b);
    layer0_outputs(6972) <= not (a xor b);
    layer0_outputs(6973) <= a or b;
    layer0_outputs(6974) <= a or b;
    layer0_outputs(6975) <= b;
    layer0_outputs(6976) <= a;
    layer0_outputs(6977) <= a xor b;
    layer0_outputs(6978) <= not (a or b);
    layer0_outputs(6979) <= not b;
    layer0_outputs(6980) <= not (a xor b);
    layer0_outputs(6981) <= not (a or b);
    layer0_outputs(6982) <= not b;
    layer0_outputs(6983) <= not (a or b);
    layer0_outputs(6984) <= not (a or b);
    layer0_outputs(6985) <= 1'b0;
    layer0_outputs(6986) <= b;
    layer0_outputs(6987) <= not b or a;
    layer0_outputs(6988) <= not (a xor b);
    layer0_outputs(6989) <= not b;
    layer0_outputs(6990) <= b;
    layer0_outputs(6991) <= not (a or b);
    layer0_outputs(6992) <= a or b;
    layer0_outputs(6993) <= not (a and b);
    layer0_outputs(6994) <= a and not b;
    layer0_outputs(6995) <= a and not b;
    layer0_outputs(6996) <= a or b;
    layer0_outputs(6997) <= not a;
    layer0_outputs(6998) <= a and b;
    layer0_outputs(6999) <= a or b;
    layer0_outputs(7000) <= b;
    layer0_outputs(7001) <= b;
    layer0_outputs(7002) <= a xor b;
    layer0_outputs(7003) <= a or b;
    layer0_outputs(7004) <= a xor b;
    layer0_outputs(7005) <= not a or b;
    layer0_outputs(7006) <= not (a xor b);
    layer0_outputs(7007) <= a or b;
    layer0_outputs(7008) <= a and not b;
    layer0_outputs(7009) <= not (a or b);
    layer0_outputs(7010) <= not (a or b);
    layer0_outputs(7011) <= 1'b0;
    layer0_outputs(7012) <= b and not a;
    layer0_outputs(7013) <= b;
    layer0_outputs(7014) <= not (a or b);
    layer0_outputs(7015) <= a;
    layer0_outputs(7016) <= b and not a;
    layer0_outputs(7017) <= b and not a;
    layer0_outputs(7018) <= not b or a;
    layer0_outputs(7019) <= not (a xor b);
    layer0_outputs(7020) <= not (a or b);
    layer0_outputs(7021) <= a or b;
    layer0_outputs(7022) <= a xor b;
    layer0_outputs(7023) <= b and not a;
    layer0_outputs(7024) <= not (a xor b);
    layer0_outputs(7025) <= not (a xor b);
    layer0_outputs(7026) <= not (a xor b);
    layer0_outputs(7027) <= a xor b;
    layer0_outputs(7028) <= not a or b;
    layer0_outputs(7029) <= not a;
    layer0_outputs(7030) <= a xor b;
    layer0_outputs(7031) <= a and not b;
    layer0_outputs(7032) <= a and not b;
    layer0_outputs(7033) <= b and not a;
    layer0_outputs(7034) <= a or b;
    layer0_outputs(7035) <= not (a or b);
    layer0_outputs(7036) <= not (a xor b);
    layer0_outputs(7037) <= a xor b;
    layer0_outputs(7038) <= not b;
    layer0_outputs(7039) <= b;
    layer0_outputs(7040) <= a;
    layer0_outputs(7041) <= not a or b;
    layer0_outputs(7042) <= a;
    layer0_outputs(7043) <= not (a or b);
    layer0_outputs(7044) <= b and not a;
    layer0_outputs(7045) <= a;
    layer0_outputs(7046) <= not b;
    layer0_outputs(7047) <= b;
    layer0_outputs(7048) <= not (a or b);
    layer0_outputs(7049) <= not (a or b);
    layer0_outputs(7050) <= not b;
    layer0_outputs(7051) <= not (a or b);
    layer0_outputs(7052) <= not (a or b);
    layer0_outputs(7053) <= not b;
    layer0_outputs(7054) <= b;
    layer0_outputs(7055) <= a or b;
    layer0_outputs(7056) <= not a or b;
    layer0_outputs(7057) <= not b or a;
    layer0_outputs(7058) <= a or b;
    layer0_outputs(7059) <= not (a or b);
    layer0_outputs(7060) <= a xor b;
    layer0_outputs(7061) <= b and not a;
    layer0_outputs(7062) <= a xor b;
    layer0_outputs(7063) <= 1'b1;
    layer0_outputs(7064) <= a and not b;
    layer0_outputs(7065) <= not (a or b);
    layer0_outputs(7066) <= a;
    layer0_outputs(7067) <= not a or b;
    layer0_outputs(7068) <= not a;
    layer0_outputs(7069) <= a xor b;
    layer0_outputs(7070) <= not (a or b);
    layer0_outputs(7071) <= b and not a;
    layer0_outputs(7072) <= a xor b;
    layer0_outputs(7073) <= not (a or b);
    layer0_outputs(7074) <= not a;
    layer0_outputs(7075) <= b and not a;
    layer0_outputs(7076) <= not b or a;
    layer0_outputs(7077) <= a or b;
    layer0_outputs(7078) <= a and b;
    layer0_outputs(7079) <= a;
    layer0_outputs(7080) <= b;
    layer0_outputs(7081) <= not (a xor b);
    layer0_outputs(7082) <= not (a or b);
    layer0_outputs(7083) <= not (a or b);
    layer0_outputs(7084) <= not (a or b);
    layer0_outputs(7085) <= not a;
    layer0_outputs(7086) <= not b;
    layer0_outputs(7087) <= a;
    layer0_outputs(7088) <= a xor b;
    layer0_outputs(7089) <= not (a or b);
    layer0_outputs(7090) <= a;
    layer0_outputs(7091) <= a or b;
    layer0_outputs(7092) <= not b;
    layer0_outputs(7093) <= not b;
    layer0_outputs(7094) <= a;
    layer0_outputs(7095) <= a and not b;
    layer0_outputs(7096) <= not a;
    layer0_outputs(7097) <= a and not b;
    layer0_outputs(7098) <= a and not b;
    layer0_outputs(7099) <= not (a and b);
    layer0_outputs(7100) <= not b or a;
    layer0_outputs(7101) <= b and not a;
    layer0_outputs(7102) <= a;
    layer0_outputs(7103) <= a and not b;
    layer0_outputs(7104) <= a or b;
    layer0_outputs(7105) <= not (a xor b);
    layer0_outputs(7106) <= b;
    layer0_outputs(7107) <= a or b;
    layer0_outputs(7108) <= not (a and b);
    layer0_outputs(7109) <= not a;
    layer0_outputs(7110) <= a or b;
    layer0_outputs(7111) <= not (a or b);
    layer0_outputs(7112) <= not (a xor b);
    layer0_outputs(7113) <= not b;
    layer0_outputs(7114) <= not (a xor b);
    layer0_outputs(7115) <= not (a xor b);
    layer0_outputs(7116) <= not a;
    layer0_outputs(7117) <= not b or a;
    layer0_outputs(7118) <= not (a and b);
    layer0_outputs(7119) <= a;
    layer0_outputs(7120) <= not (a or b);
    layer0_outputs(7121) <= b and not a;
    layer0_outputs(7122) <= b;
    layer0_outputs(7123) <= not b or a;
    layer0_outputs(7124) <= not (a or b);
    layer0_outputs(7125) <= a or b;
    layer0_outputs(7126) <= not a or b;
    layer0_outputs(7127) <= not (a xor b);
    layer0_outputs(7128) <= a or b;
    layer0_outputs(7129) <= not (a xor b);
    layer0_outputs(7130) <= b;
    layer0_outputs(7131) <= not (a and b);
    layer0_outputs(7132) <= b;
    layer0_outputs(7133) <= not a;
    layer0_outputs(7134) <= not (a or b);
    layer0_outputs(7135) <= a xor b;
    layer0_outputs(7136) <= not (a xor b);
    layer0_outputs(7137) <= not b or a;
    layer0_outputs(7138) <= not (a or b);
    layer0_outputs(7139) <= not a;
    layer0_outputs(7140) <= not (a xor b);
    layer0_outputs(7141) <= a;
    layer0_outputs(7142) <= a or b;
    layer0_outputs(7143) <= not a;
    layer0_outputs(7144) <= a and not b;
    layer0_outputs(7145) <= b and not a;
    layer0_outputs(7146) <= not a or b;
    layer0_outputs(7147) <= b and not a;
    layer0_outputs(7148) <= not (a or b);
    layer0_outputs(7149) <= not a;
    layer0_outputs(7150) <= not a or b;
    layer0_outputs(7151) <= not (a xor b);
    layer0_outputs(7152) <= not a or b;
    layer0_outputs(7153) <= not (a or b);
    layer0_outputs(7154) <= not (a or b);
    layer0_outputs(7155) <= a and not b;
    layer0_outputs(7156) <= b and not a;
    layer0_outputs(7157) <= not (a or b);
    layer0_outputs(7158) <= a xor b;
    layer0_outputs(7159) <= a;
    layer0_outputs(7160) <= a xor b;
    layer0_outputs(7161) <= not b;
    layer0_outputs(7162) <= b and not a;
    layer0_outputs(7163) <= not b;
    layer0_outputs(7164) <= a or b;
    layer0_outputs(7165) <= not a or b;
    layer0_outputs(7166) <= not (a or b);
    layer0_outputs(7167) <= not (a or b);
    layer0_outputs(7168) <= not (a or b);
    layer0_outputs(7169) <= not (a xor b);
    layer0_outputs(7170) <= a or b;
    layer0_outputs(7171) <= not b or a;
    layer0_outputs(7172) <= not a or b;
    layer0_outputs(7173) <= b and not a;
    layer0_outputs(7174) <= not b or a;
    layer0_outputs(7175) <= not b;
    layer0_outputs(7176) <= not (a xor b);
    layer0_outputs(7177) <= not a;
    layer0_outputs(7178) <= 1'b0;
    layer0_outputs(7179) <= not b or a;
    layer0_outputs(7180) <= a and not b;
    layer0_outputs(7181) <= not (a xor b);
    layer0_outputs(7182) <= not a;
    layer0_outputs(7183) <= not a or b;
    layer0_outputs(7184) <= not b or a;
    layer0_outputs(7185) <= not a or b;
    layer0_outputs(7186) <= a or b;
    layer0_outputs(7187) <= a and not b;
    layer0_outputs(7188) <= a xor b;
    layer0_outputs(7189) <= not (a or b);
    layer0_outputs(7190) <= a or b;
    layer0_outputs(7191) <= not (a or b);
    layer0_outputs(7192) <= not (a xor b);
    layer0_outputs(7193) <= a or b;
    layer0_outputs(7194) <= a and not b;
    layer0_outputs(7195) <= a and not b;
    layer0_outputs(7196) <= not b;
    layer0_outputs(7197) <= a or b;
    layer0_outputs(7198) <= b and not a;
    layer0_outputs(7199) <= not (a or b);
    layer0_outputs(7200) <= a or b;
    layer0_outputs(7201) <= a or b;
    layer0_outputs(7202) <= a and not b;
    layer0_outputs(7203) <= not (a xor b);
    layer0_outputs(7204) <= not (a xor b);
    layer0_outputs(7205) <= a or b;
    layer0_outputs(7206) <= 1'b1;
    layer0_outputs(7207) <= a or b;
    layer0_outputs(7208) <= b and not a;
    layer0_outputs(7209) <= not b;
    layer0_outputs(7210) <= not b or a;
    layer0_outputs(7211) <= not (a and b);
    layer0_outputs(7212) <= a;
    layer0_outputs(7213) <= not a or b;
    layer0_outputs(7214) <= b and not a;
    layer0_outputs(7215) <= not a;
    layer0_outputs(7216) <= not (a xor b);
    layer0_outputs(7217) <= a or b;
    layer0_outputs(7218) <= not b or a;
    layer0_outputs(7219) <= not (a xor b);
    layer0_outputs(7220) <= b and not a;
    layer0_outputs(7221) <= not b;
    layer0_outputs(7222) <= a xor b;
    layer0_outputs(7223) <= not (a or b);
    layer0_outputs(7224) <= not b or a;
    layer0_outputs(7225) <= a and not b;
    layer0_outputs(7226) <= not b;
    layer0_outputs(7227) <= not (a xor b);
    layer0_outputs(7228) <= not (a xor b);
    layer0_outputs(7229) <= not (a xor b);
    layer0_outputs(7230) <= a;
    layer0_outputs(7231) <= a;
    layer0_outputs(7232) <= not (a xor b);
    layer0_outputs(7233) <= b;
    layer0_outputs(7234) <= not (a or b);
    layer0_outputs(7235) <= not a;
    layer0_outputs(7236) <= not b;
    layer0_outputs(7237) <= not a;
    layer0_outputs(7238) <= not (a xor b);
    layer0_outputs(7239) <= a or b;
    layer0_outputs(7240) <= not a;
    layer0_outputs(7241) <= not (a or b);
    layer0_outputs(7242) <= b and not a;
    layer0_outputs(7243) <= a or b;
    layer0_outputs(7244) <= not b or a;
    layer0_outputs(7245) <= not b or a;
    layer0_outputs(7246) <= b and not a;
    layer0_outputs(7247) <= not a or b;
    layer0_outputs(7248) <= 1'b0;
    layer0_outputs(7249) <= not (a or b);
    layer0_outputs(7250) <= not a or b;
    layer0_outputs(7251) <= b;
    layer0_outputs(7252) <= not b or a;
    layer0_outputs(7253) <= a or b;
    layer0_outputs(7254) <= not a or b;
    layer0_outputs(7255) <= not a or b;
    layer0_outputs(7256) <= not b or a;
    layer0_outputs(7257) <= not (a and b);
    layer0_outputs(7258) <= a xor b;
    layer0_outputs(7259) <= a or b;
    layer0_outputs(7260) <= a and b;
    layer0_outputs(7261) <= a;
    layer0_outputs(7262) <= 1'b0;
    layer0_outputs(7263) <= not a or b;
    layer0_outputs(7264) <= a;
    layer0_outputs(7265) <= not b or a;
    layer0_outputs(7266) <= a xor b;
    layer0_outputs(7267) <= not a or b;
    layer0_outputs(7268) <= not (a xor b);
    layer0_outputs(7269) <= not (a xor b);
    layer0_outputs(7270) <= a or b;
    layer0_outputs(7271) <= not b;
    layer0_outputs(7272) <= not (a or b);
    layer0_outputs(7273) <= b and not a;
    layer0_outputs(7274) <= not a;
    layer0_outputs(7275) <= not (a xor b);
    layer0_outputs(7276) <= 1'b1;
    layer0_outputs(7277) <= a xor b;
    layer0_outputs(7278) <= not (a or b);
    layer0_outputs(7279) <= not (a or b);
    layer0_outputs(7280) <= a or b;
    layer0_outputs(7281) <= not (a xor b);
    layer0_outputs(7282) <= not a or b;
    layer0_outputs(7283) <= not (a xor b);
    layer0_outputs(7284) <= b;
    layer0_outputs(7285) <= b and not a;
    layer0_outputs(7286) <= not (a or b);
    layer0_outputs(7287) <= not (a xor b);
    layer0_outputs(7288) <= not b;
    layer0_outputs(7289) <= a;
    layer0_outputs(7290) <= not a or b;
    layer0_outputs(7291) <= b;
    layer0_outputs(7292) <= 1'b1;
    layer0_outputs(7293) <= a or b;
    layer0_outputs(7294) <= not (a or b);
    layer0_outputs(7295) <= a or b;
    layer0_outputs(7296) <= not (a or b);
    layer0_outputs(7297) <= not b or a;
    layer0_outputs(7298) <= b and not a;
    layer0_outputs(7299) <= not a;
    layer0_outputs(7300) <= not (a or b);
    layer0_outputs(7301) <= not a or b;
    layer0_outputs(7302) <= not a;
    layer0_outputs(7303) <= b and not a;
    layer0_outputs(7304) <= not (a xor b);
    layer0_outputs(7305) <= a xor b;
    layer0_outputs(7306) <= not b;
    layer0_outputs(7307) <= not (a or b);
    layer0_outputs(7308) <= b;
    layer0_outputs(7309) <= a xor b;
    layer0_outputs(7310) <= b;
    layer0_outputs(7311) <= not b or a;
    layer0_outputs(7312) <= b and not a;
    layer0_outputs(7313) <= not (a or b);
    layer0_outputs(7314) <= b and not a;
    layer0_outputs(7315) <= a and b;
    layer0_outputs(7316) <= a or b;
    layer0_outputs(7317) <= not b;
    layer0_outputs(7318) <= a and b;
    layer0_outputs(7319) <= not b;
    layer0_outputs(7320) <= not (a or b);
    layer0_outputs(7321) <= a and not b;
    layer0_outputs(7322) <= not (a or b);
    layer0_outputs(7323) <= not a;
    layer0_outputs(7324) <= a or b;
    layer0_outputs(7325) <= not a or b;
    layer0_outputs(7326) <= b and not a;
    layer0_outputs(7327) <= not (a or b);
    layer0_outputs(7328) <= 1'b0;
    layer0_outputs(7329) <= a and b;
    layer0_outputs(7330) <= b;
    layer0_outputs(7331) <= a and not b;
    layer0_outputs(7332) <= not a;
    layer0_outputs(7333) <= not (a xor b);
    layer0_outputs(7334) <= a or b;
    layer0_outputs(7335) <= not a;
    layer0_outputs(7336) <= a or b;
    layer0_outputs(7337) <= not (a or b);
    layer0_outputs(7338) <= b;
    layer0_outputs(7339) <= not (a and b);
    layer0_outputs(7340) <= b and not a;
    layer0_outputs(7341) <= a or b;
    layer0_outputs(7342) <= a or b;
    layer0_outputs(7343) <= a or b;
    layer0_outputs(7344) <= a xor b;
    layer0_outputs(7345) <= a;
    layer0_outputs(7346) <= a or b;
    layer0_outputs(7347) <= not (a xor b);
    layer0_outputs(7348) <= not (a xor b);
    layer0_outputs(7349) <= a and not b;
    layer0_outputs(7350) <= a or b;
    layer0_outputs(7351) <= a and b;
    layer0_outputs(7352) <= 1'b1;
    layer0_outputs(7353) <= a and b;
    layer0_outputs(7354) <= b and not a;
    layer0_outputs(7355) <= not b;
    layer0_outputs(7356) <= b and not a;
    layer0_outputs(7357) <= b and not a;
    layer0_outputs(7358) <= not (a or b);
    layer0_outputs(7359) <= not a;
    layer0_outputs(7360) <= a and not b;
    layer0_outputs(7361) <= b;
    layer0_outputs(7362) <= a;
    layer0_outputs(7363) <= a or b;
    layer0_outputs(7364) <= not (a or b);
    layer0_outputs(7365) <= not a;
    layer0_outputs(7366) <= a and not b;
    layer0_outputs(7367) <= not a;
    layer0_outputs(7368) <= a xor b;
    layer0_outputs(7369) <= a and not b;
    layer0_outputs(7370) <= b;
    layer0_outputs(7371) <= a xor b;
    layer0_outputs(7372) <= a or b;
    layer0_outputs(7373) <= not (a xor b);
    layer0_outputs(7374) <= not a;
    layer0_outputs(7375) <= a xor b;
    layer0_outputs(7376) <= not a or b;
    layer0_outputs(7377) <= not (a xor b);
    layer0_outputs(7378) <= a or b;
    layer0_outputs(7379) <= not a or b;
    layer0_outputs(7380) <= not b or a;
    layer0_outputs(7381) <= a and b;
    layer0_outputs(7382) <= 1'b0;
    layer0_outputs(7383) <= not (a xor b);
    layer0_outputs(7384) <= not b or a;
    layer0_outputs(7385) <= b and not a;
    layer0_outputs(7386) <= not b or a;
    layer0_outputs(7387) <= a or b;
    layer0_outputs(7388) <= a or b;
    layer0_outputs(7389) <= a xor b;
    layer0_outputs(7390) <= not a or b;
    layer0_outputs(7391) <= b;
    layer0_outputs(7392) <= not a;
    layer0_outputs(7393) <= a;
    layer0_outputs(7394) <= not b or a;
    layer0_outputs(7395) <= not (a or b);
    layer0_outputs(7396) <= not (a or b);
    layer0_outputs(7397) <= a xor b;
    layer0_outputs(7398) <= not b or a;
    layer0_outputs(7399) <= not (a or b);
    layer0_outputs(7400) <= not (a or b);
    layer0_outputs(7401) <= not a or b;
    layer0_outputs(7402) <= a xor b;
    layer0_outputs(7403) <= a;
    layer0_outputs(7404) <= not (a xor b);
    layer0_outputs(7405) <= a xor b;
    layer0_outputs(7406) <= not a or b;
    layer0_outputs(7407) <= not (a or b);
    layer0_outputs(7408) <= not (a xor b);
    layer0_outputs(7409) <= not (a xor b);
    layer0_outputs(7410) <= a;
    layer0_outputs(7411) <= a xor b;
    layer0_outputs(7412) <= a xor b;
    layer0_outputs(7413) <= not b or a;
    layer0_outputs(7414) <= a or b;
    layer0_outputs(7415) <= not b or a;
    layer0_outputs(7416) <= not b or a;
    layer0_outputs(7417) <= not (a xor b);
    layer0_outputs(7418) <= a;
    layer0_outputs(7419) <= b;
    layer0_outputs(7420) <= a xor b;
    layer0_outputs(7421) <= not b;
    layer0_outputs(7422) <= not a or b;
    layer0_outputs(7423) <= not (a xor b);
    layer0_outputs(7424) <= not b;
    layer0_outputs(7425) <= a or b;
    layer0_outputs(7426) <= a xor b;
    layer0_outputs(7427) <= a xor b;
    layer0_outputs(7428) <= a and b;
    layer0_outputs(7429) <= a;
    layer0_outputs(7430) <= not (a or b);
    layer0_outputs(7431) <= not (a and b);
    layer0_outputs(7432) <= a and b;
    layer0_outputs(7433) <= not a or b;
    layer0_outputs(7434) <= not (a or b);
    layer0_outputs(7435) <= a and not b;
    layer0_outputs(7436) <= a xor b;
    layer0_outputs(7437) <= b;
    layer0_outputs(7438) <= a xor b;
    layer0_outputs(7439) <= not a or b;
    layer0_outputs(7440) <= a xor b;
    layer0_outputs(7441) <= not (a or b);
    layer0_outputs(7442) <= not (a xor b);
    layer0_outputs(7443) <= a xor b;
    layer0_outputs(7444) <= a or b;
    layer0_outputs(7445) <= a or b;
    layer0_outputs(7446) <= not (a xor b);
    layer0_outputs(7447) <= a or b;
    layer0_outputs(7448) <= b and not a;
    layer0_outputs(7449) <= a xor b;
    layer0_outputs(7450) <= not b;
    layer0_outputs(7451) <= a xor b;
    layer0_outputs(7452) <= a or b;
    layer0_outputs(7453) <= a or b;
    layer0_outputs(7454) <= not b;
    layer0_outputs(7455) <= not (a xor b);
    layer0_outputs(7456) <= not (a or b);
    layer0_outputs(7457) <= b and not a;
    layer0_outputs(7458) <= b and not a;
    layer0_outputs(7459) <= not (a xor b);
    layer0_outputs(7460) <= not b;
    layer0_outputs(7461) <= a;
    layer0_outputs(7462) <= not b;
    layer0_outputs(7463) <= not (a or b);
    layer0_outputs(7464) <= not (a or b);
    layer0_outputs(7465) <= not a;
    layer0_outputs(7466) <= a xor b;
    layer0_outputs(7467) <= b and not a;
    layer0_outputs(7468) <= not (a xor b);
    layer0_outputs(7469) <= a;
    layer0_outputs(7470) <= a;
    layer0_outputs(7471) <= a;
    layer0_outputs(7472) <= a xor b;
    layer0_outputs(7473) <= a or b;
    layer0_outputs(7474) <= a and not b;
    layer0_outputs(7475) <= not b;
    layer0_outputs(7476) <= not b;
    layer0_outputs(7477) <= a and b;
    layer0_outputs(7478) <= not (a or b);
    layer0_outputs(7479) <= b and not a;
    layer0_outputs(7480) <= a or b;
    layer0_outputs(7481) <= not (a xor b);
    layer0_outputs(7482) <= not a or b;
    layer0_outputs(7483) <= not b;
    layer0_outputs(7484) <= a and not b;
    layer0_outputs(7485) <= a or b;
    layer0_outputs(7486) <= a and not b;
    layer0_outputs(7487) <= not b;
    layer0_outputs(7488) <= not (a or b);
    layer0_outputs(7489) <= a xor b;
    layer0_outputs(7490) <= not b or a;
    layer0_outputs(7491) <= not (a or b);
    layer0_outputs(7492) <= a;
    layer0_outputs(7493) <= a xor b;
    layer0_outputs(7494) <= b;
    layer0_outputs(7495) <= not (a xor b);
    layer0_outputs(7496) <= not (a or b);
    layer0_outputs(7497) <= a xor b;
    layer0_outputs(7498) <= not a or b;
    layer0_outputs(7499) <= a or b;
    layer0_outputs(7500) <= a or b;
    layer0_outputs(7501) <= b and not a;
    layer0_outputs(7502) <= not (a or b);
    layer0_outputs(7503) <= a or b;
    layer0_outputs(7504) <= not (a or b);
    layer0_outputs(7505) <= not (a or b);
    layer0_outputs(7506) <= not a or b;
    layer0_outputs(7507) <= not b;
    layer0_outputs(7508) <= not a;
    layer0_outputs(7509) <= not (a or b);
    layer0_outputs(7510) <= a xor b;
    layer0_outputs(7511) <= not (a xor b);
    layer0_outputs(7512) <= a;
    layer0_outputs(7513) <= not b;
    layer0_outputs(7514) <= not b or a;
    layer0_outputs(7515) <= a or b;
    layer0_outputs(7516) <= not a or b;
    layer0_outputs(7517) <= not (a or b);
    layer0_outputs(7518) <= a or b;
    layer0_outputs(7519) <= a and not b;
    layer0_outputs(7520) <= a or b;
    layer0_outputs(7521) <= not b;
    layer0_outputs(7522) <= a xor b;
    layer0_outputs(7523) <= not (a or b);
    layer0_outputs(7524) <= not (a xor b);
    layer0_outputs(7525) <= a xor b;
    layer0_outputs(7526) <= not a or b;
    layer0_outputs(7527) <= a or b;
    layer0_outputs(7528) <= a xor b;
    layer0_outputs(7529) <= not a or b;
    layer0_outputs(7530) <= b and not a;
    layer0_outputs(7531) <= not (a xor b);
    layer0_outputs(7532) <= not a;
    layer0_outputs(7533) <= not a or b;
    layer0_outputs(7534) <= a or b;
    layer0_outputs(7535) <= not a or b;
    layer0_outputs(7536) <= not (a xor b);
    layer0_outputs(7537) <= not b or a;
    layer0_outputs(7538) <= not (a or b);
    layer0_outputs(7539) <= a xor b;
    layer0_outputs(7540) <= not a or b;
    layer0_outputs(7541) <= a or b;
    layer0_outputs(7542) <= not (a or b);
    layer0_outputs(7543) <= not b or a;
    layer0_outputs(7544) <= a xor b;
    layer0_outputs(7545) <= b;
    layer0_outputs(7546) <= not b or a;
    layer0_outputs(7547) <= b;
    layer0_outputs(7548) <= b and not a;
    layer0_outputs(7549) <= not a;
    layer0_outputs(7550) <= not a;
    layer0_outputs(7551) <= a xor b;
    layer0_outputs(7552) <= a or b;
    layer0_outputs(7553) <= not b or a;
    layer0_outputs(7554) <= a or b;
    layer0_outputs(7555) <= not (a or b);
    layer0_outputs(7556) <= a or b;
    layer0_outputs(7557) <= a or b;
    layer0_outputs(7558) <= a;
    layer0_outputs(7559) <= a xor b;
    layer0_outputs(7560) <= not (a or b);
    layer0_outputs(7561) <= not a or b;
    layer0_outputs(7562) <= 1'b1;
    layer0_outputs(7563) <= not (a or b);
    layer0_outputs(7564) <= not (a or b);
    layer0_outputs(7565) <= a xor b;
    layer0_outputs(7566) <= a xor b;
    layer0_outputs(7567) <= a;
    layer0_outputs(7568) <= a and b;
    layer0_outputs(7569) <= not b or a;
    layer0_outputs(7570) <= not (a or b);
    layer0_outputs(7571) <= not (a and b);
    layer0_outputs(7572) <= not (a or b);
    layer0_outputs(7573) <= not (a xor b);
    layer0_outputs(7574) <= b;
    layer0_outputs(7575) <= not a;
    layer0_outputs(7576) <= not a;
    layer0_outputs(7577) <= a;
    layer0_outputs(7578) <= not a or b;
    layer0_outputs(7579) <= b;
    layer0_outputs(7580) <= 1'b0;
    layer0_outputs(7581) <= b;
    layer0_outputs(7582) <= a and not b;
    layer0_outputs(7583) <= a and not b;
    layer0_outputs(7584) <= not (a xor b);
    layer0_outputs(7585) <= not (a or b);
    layer0_outputs(7586) <= 1'b1;
    layer0_outputs(7587) <= a or b;
    layer0_outputs(7588) <= a or b;
    layer0_outputs(7589) <= a xor b;
    layer0_outputs(7590) <= not a;
    layer0_outputs(7591) <= not a;
    layer0_outputs(7592) <= a or b;
    layer0_outputs(7593) <= not (a xor b);
    layer0_outputs(7594) <= not (a or b);
    layer0_outputs(7595) <= b and not a;
    layer0_outputs(7596) <= a xor b;
    layer0_outputs(7597) <= b and not a;
    layer0_outputs(7598) <= a or b;
    layer0_outputs(7599) <= not (a or b);
    layer0_outputs(7600) <= not a;
    layer0_outputs(7601) <= a and b;
    layer0_outputs(7602) <= a or b;
    layer0_outputs(7603) <= 1'b0;
    layer0_outputs(7604) <= not a;
    layer0_outputs(7605) <= a or b;
    layer0_outputs(7606) <= not (a xor b);
    layer0_outputs(7607) <= a or b;
    layer0_outputs(7608) <= a or b;
    layer0_outputs(7609) <= a or b;
    layer0_outputs(7610) <= not a;
    layer0_outputs(7611) <= b;
    layer0_outputs(7612) <= b;
    layer0_outputs(7613) <= b and not a;
    layer0_outputs(7614) <= not a;
    layer0_outputs(7615) <= not a;
    layer0_outputs(7616) <= not a or b;
    layer0_outputs(7617) <= a and not b;
    layer0_outputs(7618) <= not b or a;
    layer0_outputs(7619) <= not a;
    layer0_outputs(7620) <= b;
    layer0_outputs(7621) <= a xor b;
    layer0_outputs(7622) <= a or b;
    layer0_outputs(7623) <= a or b;
    layer0_outputs(7624) <= a and not b;
    layer0_outputs(7625) <= not (a or b);
    layer0_outputs(7626) <= a or b;
    layer0_outputs(7627) <= not (a or b);
    layer0_outputs(7628) <= b;
    layer0_outputs(7629) <= not b;
    layer0_outputs(7630) <= a or b;
    layer0_outputs(7631) <= not a or b;
    layer0_outputs(7632) <= not (a or b);
    layer0_outputs(7633) <= a xor b;
    layer0_outputs(7634) <= b;
    layer0_outputs(7635) <= not (a or b);
    layer0_outputs(7636) <= not b or a;
    layer0_outputs(7637) <= not a or b;
    layer0_outputs(7638) <= a and not b;
    layer0_outputs(7639) <= not (a or b);
    layer0_outputs(7640) <= not (a or b);
    layer0_outputs(7641) <= a or b;
    layer0_outputs(7642) <= b and not a;
    layer0_outputs(7643) <= not a;
    layer0_outputs(7644) <= a and not b;
    layer0_outputs(7645) <= a or b;
    layer0_outputs(7646) <= not b or a;
    layer0_outputs(7647) <= a or b;
    layer0_outputs(7648) <= a and not b;
    layer0_outputs(7649) <= b and not a;
    layer0_outputs(7650) <= b;
    layer0_outputs(7651) <= not b or a;
    layer0_outputs(7652) <= not (a or b);
    layer0_outputs(7653) <= a and not b;
    layer0_outputs(7654) <= not (a xor b);
    layer0_outputs(7655) <= not b or a;
    layer0_outputs(7656) <= not (a xor b);
    layer0_outputs(7657) <= a;
    layer0_outputs(7658) <= not (a or b);
    layer0_outputs(7659) <= a xor b;
    layer0_outputs(7660) <= not (a xor b);
    layer0_outputs(7661) <= a;
    layer0_outputs(7662) <= a or b;
    layer0_outputs(7663) <= not a;
    layer0_outputs(7664) <= not a or b;
    layer0_outputs(7665) <= not b or a;
    layer0_outputs(7666) <= a or b;
    layer0_outputs(7667) <= a xor b;
    layer0_outputs(7668) <= not a or b;
    layer0_outputs(7669) <= not (a xor b);
    layer0_outputs(7670) <= not a or b;
    layer0_outputs(7671) <= a or b;
    layer0_outputs(7672) <= not a;
    layer0_outputs(7673) <= a;
    layer0_outputs(7674) <= not a or b;
    layer0_outputs(7675) <= not (a and b);
    layer0_outputs(7676) <= a and not b;
    layer0_outputs(7677) <= not (a or b);
    layer0_outputs(7678) <= a or b;
    layer0_outputs(7679) <= 1'b0;
    outputs(0) <= a and b;
    outputs(1) <= a xor b;
    outputs(2) <= b;
    outputs(3) <= not (a xor b);
    outputs(4) <= not a;
    outputs(5) <= not (a xor b);
    outputs(6) <= not b;
    outputs(7) <= not a;
    outputs(8) <= not (a xor b);
    outputs(9) <= not (a xor b);
    outputs(10) <= b and not a;
    outputs(11) <= not (a and b);
    outputs(12) <= b and not a;
    outputs(13) <= not (a and b);
    outputs(14) <= a;
    outputs(15) <= not b;
    outputs(16) <= not a;
    outputs(17) <= a and not b;
    outputs(18) <= a xor b;
    outputs(19) <= a and not b;
    outputs(20) <= a or b;
    outputs(21) <= a;
    outputs(22) <= not a;
    outputs(23) <= a xor b;
    outputs(24) <= a xor b;
    outputs(25) <= b;
    outputs(26) <= not b;
    outputs(27) <= not b;
    outputs(28) <= a xor b;
    outputs(29) <= b;
    outputs(30) <= a xor b;
    outputs(31) <= not b;
    outputs(32) <= b and not a;
    outputs(33) <= b;
    outputs(34) <= not b;
    outputs(35) <= not (a xor b);
    outputs(36) <= a xor b;
    outputs(37) <= not a;
    outputs(38) <= not (a or b);
    outputs(39) <= a and b;
    outputs(40) <= b;
    outputs(41) <= not b;
    outputs(42) <= not (a xor b);
    outputs(43) <= b;
    outputs(44) <= a xor b;
    outputs(45) <= not a;
    outputs(46) <= a xor b;
    outputs(47) <= not (a and b);
    outputs(48) <= b;
    outputs(49) <= not a or b;
    outputs(50) <= a xor b;
    outputs(51) <= not a;
    outputs(52) <= not (a or b);
    outputs(53) <= not a or b;
    outputs(54) <= a;
    outputs(55) <= not b;
    outputs(56) <= a;
    outputs(57) <= a;
    outputs(58) <= not a;
    outputs(59) <= a;
    outputs(60) <= b and not a;
    outputs(61) <= a;
    outputs(62) <= not (a or b);
    outputs(63) <= not b;
    outputs(64) <= a;
    outputs(65) <= b;
    outputs(66) <= not a or b;
    outputs(67) <= a xor b;
    outputs(68) <= a and not b;
    outputs(69) <= a and not b;
    outputs(70) <= a xor b;
    outputs(71) <= not (a or b);
    outputs(72) <= b;
    outputs(73) <= a and not b;
    outputs(74) <= not (a xor b);
    outputs(75) <= not (a and b);
    outputs(76) <= not a;
    outputs(77) <= not (a or b);
    outputs(78) <= a and b;
    outputs(79) <= a and b;
    outputs(80) <= not (a or b);
    outputs(81) <= not a;
    outputs(82) <= b;
    outputs(83) <= a and b;
    outputs(84) <= not a;
    outputs(85) <= a xor b;
    outputs(86) <= not a;
    outputs(87) <= not a;
    outputs(88) <= not b;
    outputs(89) <= not b;
    outputs(90) <= b and not a;
    outputs(91) <= not a;
    outputs(92) <= a and b;
    outputs(93) <= a or b;
    outputs(94) <= not a;
    outputs(95) <= a;
    outputs(96) <= a and not b;
    outputs(97) <= not b;
    outputs(98) <= a;
    outputs(99) <= not (a xor b);
    outputs(100) <= a;
    outputs(101) <= a and b;
    outputs(102) <= a or b;
    outputs(103) <= a or b;
    outputs(104) <= a xor b;
    outputs(105) <= a xor b;
    outputs(106) <= not a;
    outputs(107) <= a and not b;
    outputs(108) <= a and not b;
    outputs(109) <= not (a and b);
    outputs(110) <= not b;
    outputs(111) <= not b or a;
    outputs(112) <= b;
    outputs(113) <= b;
    outputs(114) <= a and not b;
    outputs(115) <= not a;
    outputs(116) <= not (a xor b);
    outputs(117) <= b and not a;
    outputs(118) <= not b or a;
    outputs(119) <= a;
    outputs(120) <= not a or b;
    outputs(121) <= not (a xor b);
    outputs(122) <= a or b;
    outputs(123) <= not b;
    outputs(124) <= b;
    outputs(125) <= not a;
    outputs(126) <= not (a xor b);
    outputs(127) <= a xor b;
    outputs(128) <= a xor b;
    outputs(129) <= a;
    outputs(130) <= b;
    outputs(131) <= a;
    outputs(132) <= a;
    outputs(133) <= a and not b;
    outputs(134) <= not a;
    outputs(135) <= not (a xor b);
    outputs(136) <= a;
    outputs(137) <= not b or a;
    outputs(138) <= not b;
    outputs(139) <= not (a xor b);
    outputs(140) <= not b;
    outputs(141) <= a xor b;
    outputs(142) <= a and b;
    outputs(143) <= not b;
    outputs(144) <= not (a and b);
    outputs(145) <= not (a or b);
    outputs(146) <= a or b;
    outputs(147) <= not b or a;
    outputs(148) <= not (a or b);
    outputs(149) <= b;
    outputs(150) <= not (a or b);
    outputs(151) <= b;
    outputs(152) <= not (a xor b);
    outputs(153) <= a;
    outputs(154) <= a;
    outputs(155) <= b;
    outputs(156) <= a;
    outputs(157) <= a xor b;
    outputs(158) <= a and not b;
    outputs(159) <= a xor b;
    outputs(160) <= not b or a;
    outputs(161) <= not (a or b);
    outputs(162) <= not b;
    outputs(163) <= not (a or b);
    outputs(164) <= b;
    outputs(165) <= not a;
    outputs(166) <= a and not b;
    outputs(167) <= b;
    outputs(168) <= a xor b;
    outputs(169) <= a;
    outputs(170) <= a;
    outputs(171) <= not b;
    outputs(172) <= not b or a;
    outputs(173) <= a or b;
    outputs(174) <= b;
    outputs(175) <= not a;
    outputs(176) <= a;
    outputs(177) <= a;
    outputs(178) <= not a or b;
    outputs(179) <= not (a xor b);
    outputs(180) <= a;
    outputs(181) <= not a;
    outputs(182) <= b;
    outputs(183) <= a xor b;
    outputs(184) <= b and not a;
    outputs(185) <= a;
    outputs(186) <= not b or a;
    outputs(187) <= a or b;
    outputs(188) <= b and not a;
    outputs(189) <= not (a xor b);
    outputs(190) <= a xor b;
    outputs(191) <= not (a and b);
    outputs(192) <= a and not b;
    outputs(193) <= b;
    outputs(194) <= not b;
    outputs(195) <= b and not a;
    outputs(196) <= a;
    outputs(197) <= a xor b;
    outputs(198) <= b and not a;
    outputs(199) <= a xor b;
    outputs(200) <= b;
    outputs(201) <= a;
    outputs(202) <= a and not b;
    outputs(203) <= not a;
    outputs(204) <= not (a xor b);
    outputs(205) <= a and not b;
    outputs(206) <= a;
    outputs(207) <= not b;
    outputs(208) <= a xor b;
    outputs(209) <= not a;
    outputs(210) <= b;
    outputs(211) <= not b;
    outputs(212) <= a and b;
    outputs(213) <= not a;
    outputs(214) <= not a;
    outputs(215) <= a and not b;
    outputs(216) <= not (a xor b);
    outputs(217) <= a and not b;
    outputs(218) <= a;
    outputs(219) <= a xor b;
    outputs(220) <= b;
    outputs(221) <= a;
    outputs(222) <= a xor b;
    outputs(223) <= not b or a;
    outputs(224) <= not (a and b);
    outputs(225) <= not (a xor b);
    outputs(226) <= not a or b;
    outputs(227) <= not (a xor b);
    outputs(228) <= a and not b;
    outputs(229) <= a and not b;
    outputs(230) <= a xor b;
    outputs(231) <= not a;
    outputs(232) <= not b;
    outputs(233) <= a xor b;
    outputs(234) <= not b;
    outputs(235) <= a xor b;
    outputs(236) <= b and not a;
    outputs(237) <= a and b;
    outputs(238) <= a;
    outputs(239) <= a xor b;
    outputs(240) <= not b;
    outputs(241) <= a and b;
    outputs(242) <= b;
    outputs(243) <= not (a xor b);
    outputs(244) <= not a;
    outputs(245) <= a and b;
    outputs(246) <= a and b;
    outputs(247) <= a and not b;
    outputs(248) <= not b;
    outputs(249) <= a;
    outputs(250) <= not a;
    outputs(251) <= b;
    outputs(252) <= a;
    outputs(253) <= not b;
    outputs(254) <= a and not b;
    outputs(255) <= not (a xor b);
    outputs(256) <= a;
    outputs(257) <= not (a xor b);
    outputs(258) <= not (a xor b);
    outputs(259) <= b;
    outputs(260) <= b;
    outputs(261) <= not b or a;
    outputs(262) <= a xor b;
    outputs(263) <= a xor b;
    outputs(264) <= a xor b;
    outputs(265) <= a;
    outputs(266) <= a;
    outputs(267) <= a;
    outputs(268) <= not a;
    outputs(269) <= not b;
    outputs(270) <= not (a xor b);
    outputs(271) <= b;
    outputs(272) <= a xor b;
    outputs(273) <= not (a and b);
    outputs(274) <= not (a and b);
    outputs(275) <= a xor b;
    outputs(276) <= not (a and b);
    outputs(277) <= b;
    outputs(278) <= a;
    outputs(279) <= not b;
    outputs(280) <= a and not b;
    outputs(281) <= a and not b;
    outputs(282) <= a xor b;
    outputs(283) <= not a or b;
    outputs(284) <= a xor b;
    outputs(285) <= not a;
    outputs(286) <= a and not b;
    outputs(287) <= b;
    outputs(288) <= not a or b;
    outputs(289) <= not b;
    outputs(290) <= not b;
    outputs(291) <= a;
    outputs(292) <= not (a xor b);
    outputs(293) <= a;
    outputs(294) <= b and not a;
    outputs(295) <= a;
    outputs(296) <= b;
    outputs(297) <= not (a xor b);
    outputs(298) <= a;
    outputs(299) <= b;
    outputs(300) <= b;
    outputs(301) <= a and not b;
    outputs(302) <= b and not a;
    outputs(303) <= a;
    outputs(304) <= b and not a;
    outputs(305) <= b and not a;
    outputs(306) <= a;
    outputs(307) <= b and not a;
    outputs(308) <= not b;
    outputs(309) <= a xor b;
    outputs(310) <= not (a xor b);
    outputs(311) <= a;
    outputs(312) <= a xor b;
    outputs(313) <= not (a xor b);
    outputs(314) <= not b;
    outputs(315) <= not a;
    outputs(316) <= b;
    outputs(317) <= b;
    outputs(318) <= a;
    outputs(319) <= not a or b;
    outputs(320) <= a and not b;
    outputs(321) <= not (a or b);
    outputs(322) <= a and not b;
    outputs(323) <= a or b;
    outputs(324) <= a and not b;
    outputs(325) <= b;
    outputs(326) <= not b;
    outputs(327) <= not b;
    outputs(328) <= not a;
    outputs(329) <= b;
    outputs(330) <= not (a xor b);
    outputs(331) <= b;
    outputs(332) <= not a;
    outputs(333) <= a and b;
    outputs(334) <= not b;
    outputs(335) <= a;
    outputs(336) <= not (a xor b);
    outputs(337) <= not (a xor b);
    outputs(338) <= not (a or b);
    outputs(339) <= not b;
    outputs(340) <= not a;
    outputs(341) <= not (a xor b);
    outputs(342) <= not b;
    outputs(343) <= a;
    outputs(344) <= a xor b;
    outputs(345) <= not (a and b);
    outputs(346) <= not (a xor b);
    outputs(347) <= not (a xor b);
    outputs(348) <= not (a xor b);
    outputs(349) <= a and not b;
    outputs(350) <= b and not a;
    outputs(351) <= a;
    outputs(352) <= a and not b;
    outputs(353) <= not (a xor b);
    outputs(354) <= not a;
    outputs(355) <= not (a xor b);
    outputs(356) <= not a;
    outputs(357) <= not (a or b);
    outputs(358) <= a;
    outputs(359) <= not a;
    outputs(360) <= a and b;
    outputs(361) <= b;
    outputs(362) <= not a;
    outputs(363) <= not (a or b);
    outputs(364) <= b and not a;
    outputs(365) <= b and not a;
    outputs(366) <= a and not b;
    outputs(367) <= b;
    outputs(368) <= not b;
    outputs(369) <= b;
    outputs(370) <= not a;
    outputs(371) <= not (a or b);
    outputs(372) <= a and b;
    outputs(373) <= a and not b;
    outputs(374) <= not b;
    outputs(375) <= a and b;
    outputs(376) <= b;
    outputs(377) <= not a;
    outputs(378) <= a xor b;
    outputs(379) <= a xor b;
    outputs(380) <= a xor b;
    outputs(381) <= a;
    outputs(382) <= a or b;
    outputs(383) <= not a;
    outputs(384) <= a xor b;
    outputs(385) <= a or b;
    outputs(386) <= not b or a;
    outputs(387) <= not (a xor b);
    outputs(388) <= b and not a;
    outputs(389) <= not a;
    outputs(390) <= a and b;
    outputs(391) <= a and b;
    outputs(392) <= not b;
    outputs(393) <= not b or a;
    outputs(394) <= not a or b;
    outputs(395) <= not a;
    outputs(396) <= not a or b;
    outputs(397) <= not (a and b);
    outputs(398) <= not (a or b);
    outputs(399) <= a and b;
    outputs(400) <= a and b;
    outputs(401) <= not b;
    outputs(402) <= not (a xor b);
    outputs(403) <= b and not a;
    outputs(404) <= not b;
    outputs(405) <= a xor b;
    outputs(406) <= not b;
    outputs(407) <= b;
    outputs(408) <= not (a xor b);
    outputs(409) <= a xor b;
    outputs(410) <= b and not a;
    outputs(411) <= a and b;
    outputs(412) <= not b;
    outputs(413) <= a;
    outputs(414) <= not (a xor b);
    outputs(415) <= a;
    outputs(416) <= a;
    outputs(417) <= b and not a;
    outputs(418) <= a xor b;
    outputs(419) <= a and b;
    outputs(420) <= a and not b;
    outputs(421) <= not (a and b);
    outputs(422) <= a xor b;
    outputs(423) <= b;
    outputs(424) <= a and not b;
    outputs(425) <= b and not a;
    outputs(426) <= b and not a;
    outputs(427) <= not b;
    outputs(428) <= b;
    outputs(429) <= not b;
    outputs(430) <= not a;
    outputs(431) <= not (a xor b);
    outputs(432) <= not b or a;
    outputs(433) <= not b;
    outputs(434) <= b and not a;
    outputs(435) <= a and not b;
    outputs(436) <= not (a xor b);
    outputs(437) <= not b;
    outputs(438) <= not (a xor b);
    outputs(439) <= a xor b;
    outputs(440) <= not b or a;
    outputs(441) <= not (a xor b);
    outputs(442) <= b;
    outputs(443) <= a xor b;
    outputs(444) <= a;
    outputs(445) <= not (a xor b);
    outputs(446) <= not (a or b);
    outputs(447) <= not b;
    outputs(448) <= not b;
    outputs(449) <= a;
    outputs(450) <= a and b;
    outputs(451) <= not a;
    outputs(452) <= not b;
    outputs(453) <= b;
    outputs(454) <= not b;
    outputs(455) <= not b;
    outputs(456) <= not a;
    outputs(457) <= b;
    outputs(458) <= not (a or b);
    outputs(459) <= not b or a;
    outputs(460) <= not b;
    outputs(461) <= b and not a;
    outputs(462) <= b;
    outputs(463) <= not (a xor b);
    outputs(464) <= b and not a;
    outputs(465) <= not b;
    outputs(466) <= not a;
    outputs(467) <= a;
    outputs(468) <= not b;
    outputs(469) <= not (a xor b);
    outputs(470) <= not (a and b);
    outputs(471) <= not a;
    outputs(472) <= not a;
    outputs(473) <= not a;
    outputs(474) <= b;
    outputs(475) <= a;
    outputs(476) <= a and not b;
    outputs(477) <= a;
    outputs(478) <= b;
    outputs(479) <= not (a xor b);
    outputs(480) <= not (a or b);
    outputs(481) <= not a;
    outputs(482) <= not (a xor b);
    outputs(483) <= not (a xor b);
    outputs(484) <= b and not a;
    outputs(485) <= b;
    outputs(486) <= a;
    outputs(487) <= a and not b;
    outputs(488) <= b and not a;
    outputs(489) <= not b;
    outputs(490) <= b;
    outputs(491) <= not (a or b);
    outputs(492) <= a;
    outputs(493) <= a xor b;
    outputs(494) <= not a;
    outputs(495) <= not a;
    outputs(496) <= a xor b;
    outputs(497) <= not (a and b);
    outputs(498) <= not a;
    outputs(499) <= not b;
    outputs(500) <= a xor b;
    outputs(501) <= not b or a;
    outputs(502) <= b;
    outputs(503) <= a xor b;
    outputs(504) <= not a;
    outputs(505) <= not (a xor b);
    outputs(506) <= a;
    outputs(507) <= a and not b;
    outputs(508) <= not b;
    outputs(509) <= not a;
    outputs(510) <= a and not b;
    outputs(511) <= not b;
    outputs(512) <= not a;
    outputs(513) <= b and not a;
    outputs(514) <= a or b;
    outputs(515) <= not a or b;
    outputs(516) <= not a;
    outputs(517) <= a or b;
    outputs(518) <= not (a or b);
    outputs(519) <= a and not b;
    outputs(520) <= not (a xor b);
    outputs(521) <= b;
    outputs(522) <= not b;
    outputs(523) <= not (a xor b);
    outputs(524) <= a and not b;
    outputs(525) <= b;
    outputs(526) <= b;
    outputs(527) <= a and not b;
    outputs(528) <= not (a or b);
    outputs(529) <= a xor b;
    outputs(530) <= not a;
    outputs(531) <= not b;
    outputs(532) <= not b;
    outputs(533) <= a xor b;
    outputs(534) <= not (a or b);
    outputs(535) <= a xor b;
    outputs(536) <= a xor b;
    outputs(537) <= a;
    outputs(538) <= not (a or b);
    outputs(539) <= not a or b;
    outputs(540) <= a and not b;
    outputs(541) <= not b;
    outputs(542) <= not b;
    outputs(543) <= a;
    outputs(544) <= not b;
    outputs(545) <= a or b;
    outputs(546) <= not b;
    outputs(547) <= not b;
    outputs(548) <= not b;
    outputs(549) <= a and b;
    outputs(550) <= not a;
    outputs(551) <= not a;
    outputs(552) <= a;
    outputs(553) <= not a;
    outputs(554) <= not b;
    outputs(555) <= not b;
    outputs(556) <= a xor b;
    outputs(557) <= b;
    outputs(558) <= b;
    outputs(559) <= b and not a;
    outputs(560) <= a xor b;
    outputs(561) <= b and not a;
    outputs(562) <= not b;
    outputs(563) <= not (a xor b);
    outputs(564) <= not (a xor b);
    outputs(565) <= a;
    outputs(566) <= not a;
    outputs(567) <= b;
    outputs(568) <= not b;
    outputs(569) <= a;
    outputs(570) <= not (a or b);
    outputs(571) <= not a;
    outputs(572) <= not (a xor b);
    outputs(573) <= a;
    outputs(574) <= not a;
    outputs(575) <= not b;
    outputs(576) <= a xor b;
    outputs(577) <= not b;
    outputs(578) <= not b;
    outputs(579) <= not b or a;
    outputs(580) <= a and not b;
    outputs(581) <= a xor b;
    outputs(582) <= a;
    outputs(583) <= a and not b;
    outputs(584) <= a xor b;
    outputs(585) <= a;
    outputs(586) <= a xor b;
    outputs(587) <= a and not b;
    outputs(588) <= a xor b;
    outputs(589) <= not (a and b);
    outputs(590) <= b;
    outputs(591) <= a;
    outputs(592) <= b;
    outputs(593) <= a;
    outputs(594) <= not a;
    outputs(595) <= not (a and b);
    outputs(596) <= b and not a;
    outputs(597) <= a xor b;
    outputs(598) <= not b;
    outputs(599) <= not a;
    outputs(600) <= not a;
    outputs(601) <= not a;
    outputs(602) <= a and b;
    outputs(603) <= 1'b0;
    outputs(604) <= b;
    outputs(605) <= a xor b;
    outputs(606) <= a or b;
    outputs(607) <= not b;
    outputs(608) <= not (a or b);
    outputs(609) <= not (a or b);
    outputs(610) <= not b;
    outputs(611) <= a and b;
    outputs(612) <= not b or a;
    outputs(613) <= a;
    outputs(614) <= a and not b;
    outputs(615) <= not (a xor b);
    outputs(616) <= not (a xor b);
    outputs(617) <= a and not b;
    outputs(618) <= not b or a;
    outputs(619) <= not b;
    outputs(620) <= a and not b;
    outputs(621) <= b and not a;
    outputs(622) <= not (a xor b);
    outputs(623) <= not (a or b);
    outputs(624) <= a and b;
    outputs(625) <= not (a xor b);
    outputs(626) <= not b;
    outputs(627) <= a xor b;
    outputs(628) <= b and not a;
    outputs(629) <= a;
    outputs(630) <= not b;
    outputs(631) <= not (a xor b);
    outputs(632) <= a xor b;
    outputs(633) <= b;
    outputs(634) <= a and not b;
    outputs(635) <= a;
    outputs(636) <= not (a xor b);
    outputs(637) <= a or b;
    outputs(638) <= a and b;
    outputs(639) <= a;
    outputs(640) <= not b or a;
    outputs(641) <= a;
    outputs(642) <= a;
    outputs(643) <= a xor b;
    outputs(644) <= a xor b;
    outputs(645) <= b;
    outputs(646) <= b and not a;
    outputs(647) <= a and not b;
    outputs(648) <= a xor b;
    outputs(649) <= not b;
    outputs(650) <= not a;
    outputs(651) <= a and b;
    outputs(652) <= not a or b;
    outputs(653) <= b and not a;
    outputs(654) <= not b;
    outputs(655) <= b;
    outputs(656) <= b and not a;
    outputs(657) <= a;
    outputs(658) <= not (a xor b);
    outputs(659) <= not a or b;
    outputs(660) <= a;
    outputs(661) <= not (a xor b);
    outputs(662) <= a xor b;
    outputs(663) <= a and not b;
    outputs(664) <= a and not b;
    outputs(665) <= not b;
    outputs(666) <= not (a xor b);
    outputs(667) <= a xor b;
    outputs(668) <= not (a and b);
    outputs(669) <= not (a xor b);
    outputs(670) <= b and not a;
    outputs(671) <= a;
    outputs(672) <= a or b;
    outputs(673) <= not a;
    outputs(674) <= not b;
    outputs(675) <= not (a or b);
    outputs(676) <= not a;
    outputs(677) <= not b or a;
    outputs(678) <= a and b;
    outputs(679) <= b;
    outputs(680) <= not (a xor b);
    outputs(681) <= not (a xor b);
    outputs(682) <= a;
    outputs(683) <= b;
    outputs(684) <= a or b;
    outputs(685) <= not a or b;
    outputs(686) <= a xor b;
    outputs(687) <= b;
    outputs(688) <= a and b;
    outputs(689) <= not b;
    outputs(690) <= not a;
    outputs(691) <= b;
    outputs(692) <= not (a xor b);
    outputs(693) <= a xor b;
    outputs(694) <= not a;
    outputs(695) <= b;
    outputs(696) <= a xor b;
    outputs(697) <= a and b;
    outputs(698) <= not a;
    outputs(699) <= a xor b;
    outputs(700) <= b and not a;
    outputs(701) <= a xor b;
    outputs(702) <= not a;
    outputs(703) <= not (a xor b);
    outputs(704) <= a;
    outputs(705) <= not a;
    outputs(706) <= not b;
    outputs(707) <= not a;
    outputs(708) <= not a or b;
    outputs(709) <= not (a xor b);
    outputs(710) <= a xor b;
    outputs(711) <= b and not a;
    outputs(712) <= a and b;
    outputs(713) <= not a;
    outputs(714) <= b;
    outputs(715) <= a and not b;
    outputs(716) <= not b or a;
    outputs(717) <= not (a xor b);
    outputs(718) <= b;
    outputs(719) <= not a or b;
    outputs(720) <= not (a and b);
    outputs(721) <= not b;
    outputs(722) <= a;
    outputs(723) <= b;
    outputs(724) <= b;
    outputs(725) <= not b;
    outputs(726) <= not (a and b);
    outputs(727) <= b;
    outputs(728) <= not (a xor b);
    outputs(729) <= a;
    outputs(730) <= not b;
    outputs(731) <= not (a xor b);
    outputs(732) <= a;
    outputs(733) <= b;
    outputs(734) <= b;
    outputs(735) <= a xor b;
    outputs(736) <= b;
    outputs(737) <= not a or b;
    outputs(738) <= not a;
    outputs(739) <= not (a xor b);
    outputs(740) <= not a;
    outputs(741) <= not b or a;
    outputs(742) <= not b or a;
    outputs(743) <= not (a xor b);
    outputs(744) <= a xor b;
    outputs(745) <= b;
    outputs(746) <= not (a or b);
    outputs(747) <= b;
    outputs(748) <= not (a xor b);
    outputs(749) <= not a;
    outputs(750) <= b and not a;
    outputs(751) <= not a;
    outputs(752) <= not (a or b);
    outputs(753) <= a;
    outputs(754) <= b;
    outputs(755) <= a;
    outputs(756) <= not b;
    outputs(757) <= not (a or b);
    outputs(758) <= not (a or b);
    outputs(759) <= not a;
    outputs(760) <= a xor b;
    outputs(761) <= b and not a;
    outputs(762) <= not (a xor b);
    outputs(763) <= a and b;
    outputs(764) <= not (a xor b);
    outputs(765) <= not (a or b);
    outputs(766) <= a;
    outputs(767) <= a and b;
    outputs(768) <= a and b;
    outputs(769) <= a xor b;
    outputs(770) <= a;
    outputs(771) <= a and b;
    outputs(772) <= not a;
    outputs(773) <= b;
    outputs(774) <= not (a or b);
    outputs(775) <= not b or a;
    outputs(776) <= b;
    outputs(777) <= a and not b;
    outputs(778) <= not a;
    outputs(779) <= a;
    outputs(780) <= not (a or b);
    outputs(781) <= b;
    outputs(782) <= b and not a;
    outputs(783) <= b and not a;
    outputs(784) <= not (a xor b);
    outputs(785) <= b;
    outputs(786) <= a and b;
    outputs(787) <= a and not b;
    outputs(788) <= not (a or b);
    outputs(789) <= not (a or b);
    outputs(790) <= a and b;
    outputs(791) <= a xor b;
    outputs(792) <= b and not a;
    outputs(793) <= b and not a;
    outputs(794) <= a xor b;
    outputs(795) <= not b;
    outputs(796) <= not (a or b);
    outputs(797) <= not (a or b);
    outputs(798) <= b and not a;
    outputs(799) <= a xor b;
    outputs(800) <= a and not b;
    outputs(801) <= not (a or b);
    outputs(802) <= a xor b;
    outputs(803) <= b;
    outputs(804) <= b and not a;
    outputs(805) <= a and b;
    outputs(806) <= b and not a;
    outputs(807) <= a and not b;
    outputs(808) <= b and not a;
    outputs(809) <= not a;
    outputs(810) <= b and not a;
    outputs(811) <= b;
    outputs(812) <= a and b;
    outputs(813) <= a xor b;
    outputs(814) <= b and not a;
    outputs(815) <= a and not b;
    outputs(816) <= not a;
    outputs(817) <= a and not b;
    outputs(818) <= a and b;
    outputs(819) <= a and not b;
    outputs(820) <= not (a xor b);
    outputs(821) <= not (a or b);
    outputs(822) <= a xor b;
    outputs(823) <= a and b;
    outputs(824) <= a and b;
    outputs(825) <= a and not b;
    outputs(826) <= not (a or b);
    outputs(827) <= not (a or b);
    outputs(828) <= not (a or b);
    outputs(829) <= b and not a;
    outputs(830) <= a and not b;
    outputs(831) <= not (a xor b);
    outputs(832) <= not a;
    outputs(833) <= a and not b;
    outputs(834) <= a;
    outputs(835) <= not a;
    outputs(836) <= a and b;
    outputs(837) <= a and b;
    outputs(838) <= not b;
    outputs(839) <= not (a or b);
    outputs(840) <= not (a or b);
    outputs(841) <= a and b;
    outputs(842) <= a and not b;
    outputs(843) <= not (a xor b);
    outputs(844) <= b;
    outputs(845) <= b and not a;
    outputs(846) <= not (a or b);
    outputs(847) <= b;
    outputs(848) <= 1'b0;
    outputs(849) <= not a;
    outputs(850) <= a;
    outputs(851) <= not (a or b);
    outputs(852) <= not b;
    outputs(853) <= b and not a;
    outputs(854) <= a and not b;
    outputs(855) <= b and not a;
    outputs(856) <= 1'b0;
    outputs(857) <= not a;
    outputs(858) <= b and not a;
    outputs(859) <= not (a or b);
    outputs(860) <= not a;
    outputs(861) <= a and not b;
    outputs(862) <= a and b;
    outputs(863) <= a and not b;
    outputs(864) <= not b;
    outputs(865) <= a;
    outputs(866) <= not (a or b);
    outputs(867) <= a and not b;
    outputs(868) <= not (a or b);
    outputs(869) <= 1'b0;
    outputs(870) <= a and not b;
    outputs(871) <= a and b;
    outputs(872) <= not (a xor b);
    outputs(873) <= b and not a;
    outputs(874) <= a and b;
    outputs(875) <= not b;
    outputs(876) <= a;
    outputs(877) <= not (a or b);
    outputs(878) <= b and not a;
    outputs(879) <= a and b;
    outputs(880) <= a and b;
    outputs(881) <= a xor b;
    outputs(882) <= a and not b;
    outputs(883) <= b and not a;
    outputs(884) <= a xor b;
    outputs(885) <= not (a xor b);
    outputs(886) <= not (a xor b);
    outputs(887) <= not b;
    outputs(888) <= b and not a;
    outputs(889) <= not (a xor b);
    outputs(890) <= b and not a;
    outputs(891) <= b and not a;
    outputs(892) <= not a;
    outputs(893) <= b and not a;
    outputs(894) <= a and b;
    outputs(895) <= a and b;
    outputs(896) <= not a;
    outputs(897) <= a and not b;
    outputs(898) <= b;
    outputs(899) <= a;
    outputs(900) <= not (a or b);
    outputs(901) <= a xor b;
    outputs(902) <= a and b;
    outputs(903) <= b;
    outputs(904) <= not (a or b);
    outputs(905) <= a and b;
    outputs(906) <= b and not a;
    outputs(907) <= not b;
    outputs(908) <= b and not a;
    outputs(909) <= not b;
    outputs(910) <= a and not b;
    outputs(911) <= a and not b;
    outputs(912) <= not b or a;
    outputs(913) <= a xor b;
    outputs(914) <= b and not a;
    outputs(915) <= not b;
    outputs(916) <= b and not a;
    outputs(917) <= b;
    outputs(918) <= not (a or b);
    outputs(919) <= b;
    outputs(920) <= not b;
    outputs(921) <= a and b;
    outputs(922) <= not (a or b);
    outputs(923) <= a and not b;
    outputs(924) <= b;
    outputs(925) <= b and not a;
    outputs(926) <= b and not a;
    outputs(927) <= not a;
    outputs(928) <= not (a xor b);
    outputs(929) <= b and not a;
    outputs(930) <= not a;
    outputs(931) <= b and not a;
    outputs(932) <= b and not a;
    outputs(933) <= not (a or b);
    outputs(934) <= not (a or b);
    outputs(935) <= a and not b;
    outputs(936) <= not b;
    outputs(937) <= a and b;
    outputs(938) <= a xor b;
    outputs(939) <= a;
    outputs(940) <= a xor b;
    outputs(941) <= b and not a;
    outputs(942) <= not (a or b);
    outputs(943) <= b and not a;
    outputs(944) <= not (a or b);
    outputs(945) <= b and not a;
    outputs(946) <= a xor b;
    outputs(947) <= not (a or b);
    outputs(948) <= a and b;
    outputs(949) <= not b;
    outputs(950) <= not a;
    outputs(951) <= not (a xor b);
    outputs(952) <= a and b;
    outputs(953) <= a and not b;
    outputs(954) <= a and not b;
    outputs(955) <= not b;
    outputs(956) <= b and not a;
    outputs(957) <= a and not b;
    outputs(958) <= b and not a;
    outputs(959) <= b and not a;
    outputs(960) <= b and not a;
    outputs(961) <= a and b;
    outputs(962) <= a and b;
    outputs(963) <= not a;
    outputs(964) <= a and b;
    outputs(965) <= a and not b;
    outputs(966) <= a and b;
    outputs(967) <= b and not a;
    outputs(968) <= b and not a;
    outputs(969) <= a;
    outputs(970) <= a and not b;
    outputs(971) <= a and not b;
    outputs(972) <= not (a xor b);
    outputs(973) <= not (a xor b);
    outputs(974) <= not a;
    outputs(975) <= not (a or b);
    outputs(976) <= a and b;
    outputs(977) <= b;
    outputs(978) <= b;
    outputs(979) <= not (a or b);
    outputs(980) <= a xor b;
    outputs(981) <= not (a xor b);
    outputs(982) <= b and not a;
    outputs(983) <= not (a xor b);
    outputs(984) <= a;
    outputs(985) <= a and b;
    outputs(986) <= not b;
    outputs(987) <= a and not b;
    outputs(988) <= not (a or b);
    outputs(989) <= not (a or b);
    outputs(990) <= not b;
    outputs(991) <= a and b;
    outputs(992) <= a and b;
    outputs(993) <= not (a xor b);
    outputs(994) <= a;
    outputs(995) <= b and not a;
    outputs(996) <= a xor b;
    outputs(997) <= a and b;
    outputs(998) <= b and not a;
    outputs(999) <= not (a or b);
    outputs(1000) <= b;
    outputs(1001) <= a;
    outputs(1002) <= not a;
    outputs(1003) <= not (a or b);
    outputs(1004) <= a and b;
    outputs(1005) <= not (a or b);
    outputs(1006) <= 1'b0;
    outputs(1007) <= 1'b0;
    outputs(1008) <= a and not b;
    outputs(1009) <= a and not b;
    outputs(1010) <= a and not b;
    outputs(1011) <= b and not a;
    outputs(1012) <= not (a xor b);
    outputs(1013) <= a;
    outputs(1014) <= not (a xor b);
    outputs(1015) <= not (a or b);
    outputs(1016) <= a xor b;
    outputs(1017) <= not (a xor b);
    outputs(1018) <= not (a or b);
    outputs(1019) <= not (a xor b);
    outputs(1020) <= not a;
    outputs(1021) <= not b;
    outputs(1022) <= a and not b;
    outputs(1023) <= a and not b;
    outputs(1024) <= a and not b;
    outputs(1025) <= not (a or b);
    outputs(1026) <= b;
    outputs(1027) <= a and b;
    outputs(1028) <= not a or b;
    outputs(1029) <= a;
    outputs(1030) <= not a;
    outputs(1031) <= not b;
    outputs(1032) <= not a;
    outputs(1033) <= a and not b;
    outputs(1034) <= 1'b0;
    outputs(1035) <= a and not b;
    outputs(1036) <= not b;
    outputs(1037) <= not (a or b);
    outputs(1038) <= a and b;
    outputs(1039) <= b and not a;
    outputs(1040) <= not b;
    outputs(1041) <= a and b;
    outputs(1042) <= a and not b;
    outputs(1043) <= not (a or b);
    outputs(1044) <= not (a xor b);
    outputs(1045) <= not (a or b);
    outputs(1046) <= a and not b;
    outputs(1047) <= not (a xor b);
    outputs(1048) <= b and not a;
    outputs(1049) <= a and not b;
    outputs(1050) <= not (a xor b);
    outputs(1051) <= a and not b;
    outputs(1052) <= a xor b;
    outputs(1053) <= a and not b;
    outputs(1054) <= not (a xor b);
    outputs(1055) <= not (a xor b);
    outputs(1056) <= not (a xor b);
    outputs(1057) <= a and not b;
    outputs(1058) <= a xor b;
    outputs(1059) <= a and not b;
    outputs(1060) <= a and b;
    outputs(1061) <= not a;
    outputs(1062) <= a and not b;
    outputs(1063) <= a;
    outputs(1064) <= a and not b;
    outputs(1065) <= a;
    outputs(1066) <= a and not b;
    outputs(1067) <= a and b;
    outputs(1068) <= a;
    outputs(1069) <= a and b;
    outputs(1070) <= not (a or b);
    outputs(1071) <= a;
    outputs(1072) <= not (a and b);
    outputs(1073) <= not a;
    outputs(1074) <= not a;
    outputs(1075) <= a and b;
    outputs(1076) <= a and b;
    outputs(1077) <= not (a or b);
    outputs(1078) <= not (a or b);
    outputs(1079) <= b and not a;
    outputs(1080) <= a and not b;
    outputs(1081) <= a and b;
    outputs(1082) <= a and not b;
    outputs(1083) <= b and not a;
    outputs(1084) <= a xor b;
    outputs(1085) <= a xor b;
    outputs(1086) <= not (a or b);
    outputs(1087) <= a and not b;
    outputs(1088) <= not a;
    outputs(1089) <= not (a or b);
    outputs(1090) <= not (a xor b);
    outputs(1091) <= a;
    outputs(1092) <= a xor b;
    outputs(1093) <= a and not b;
    outputs(1094) <= not (a xor b);
    outputs(1095) <= b and not a;
    outputs(1096) <= b and not a;
    outputs(1097) <= not (a or b);
    outputs(1098) <= not (a xor b);
    outputs(1099) <= a and not b;
    outputs(1100) <= a xor b;
    outputs(1101) <= a and not b;
    outputs(1102) <= not b;
    outputs(1103) <= a and b;
    outputs(1104) <= b and not a;
    outputs(1105) <= a xor b;
    outputs(1106) <= a and not b;
    outputs(1107) <= a and b;
    outputs(1108) <= not (a or b);
    outputs(1109) <= a and not b;
    outputs(1110) <= not (a or b);
    outputs(1111) <= b and not a;
    outputs(1112) <= not (a or b);
    outputs(1113) <= b;
    outputs(1114) <= b;
    outputs(1115) <= b and not a;
    outputs(1116) <= b and not a;
    outputs(1117) <= a;
    outputs(1118) <= b;
    outputs(1119) <= b and not a;
    outputs(1120) <= b;
    outputs(1121) <= not (a or b);
    outputs(1122) <= a and not b;
    outputs(1123) <= not (a xor b);
    outputs(1124) <= a and not b;
    outputs(1125) <= a and b;
    outputs(1126) <= a and not b;
    outputs(1127) <= a;
    outputs(1128) <= 1'b0;
    outputs(1129) <= a and not b;
    outputs(1130) <= b and not a;
    outputs(1131) <= a and b;
    outputs(1132) <= not b;
    outputs(1133) <= not b;
    outputs(1134) <= b and not a;
    outputs(1135) <= not (a or b);
    outputs(1136) <= a and not b;
    outputs(1137) <= not a;
    outputs(1138) <= a;
    outputs(1139) <= a and b;
    outputs(1140) <= a;
    outputs(1141) <= a and b;
    outputs(1142) <= a and not b;
    outputs(1143) <= not b;
    outputs(1144) <= 1'b0;
    outputs(1145) <= not (a or b);
    outputs(1146) <= not (a or b);
    outputs(1147) <= not (a or b);
    outputs(1148) <= a xor b;
    outputs(1149) <= a and not b;
    outputs(1150) <= a xor b;
    outputs(1151) <= not (a or b);
    outputs(1152) <= 1'b0;
    outputs(1153) <= not (a xor b);
    outputs(1154) <= b and not a;
    outputs(1155) <= not (a or b);
    outputs(1156) <= not a;
    outputs(1157) <= not (a or b);
    outputs(1158) <= a and not b;
    outputs(1159) <= b and not a;
    outputs(1160) <= not (a or b);
    outputs(1161) <= a;
    outputs(1162) <= a;
    outputs(1163) <= a and not b;
    outputs(1164) <= b;
    outputs(1165) <= not (a xor b);
    outputs(1166) <= a and not b;
    outputs(1167) <= 1'b0;
    outputs(1168) <= a and not b;
    outputs(1169) <= a and not b;
    outputs(1170) <= a and b;
    outputs(1171) <= a xor b;
    outputs(1172) <= b;
    outputs(1173) <= not (a or b);
    outputs(1174) <= a and not b;
    outputs(1175) <= not a;
    outputs(1176) <= b and not a;
    outputs(1177) <= a and not b;
    outputs(1178) <= not a;
    outputs(1179) <= b and not a;
    outputs(1180) <= not a;
    outputs(1181) <= not (a or b);
    outputs(1182) <= a xor b;
    outputs(1183) <= a and b;
    outputs(1184) <= 1'b0;
    outputs(1185) <= a xor b;
    outputs(1186) <= not (a or b);
    outputs(1187) <= b and not a;
    outputs(1188) <= b and not a;
    outputs(1189) <= a and b;
    outputs(1190) <= a;
    outputs(1191) <= a xor b;
    outputs(1192) <= a xor b;
    outputs(1193) <= a and b;
    outputs(1194) <= a and b;
    outputs(1195) <= not a;
    outputs(1196) <= not b or a;
    outputs(1197) <= not (a or b);
    outputs(1198) <= a and b;
    outputs(1199) <= not (a or b);
    outputs(1200) <= not a;
    outputs(1201) <= not b;
    outputs(1202) <= a and not b;
    outputs(1203) <= a and not b;
    outputs(1204) <= a and not b;
    outputs(1205) <= b and not a;
    outputs(1206) <= 1'b0;
    outputs(1207) <= a;
    outputs(1208) <= a and not b;
    outputs(1209) <= not b;
    outputs(1210) <= 1'b0;
    outputs(1211) <= a;
    outputs(1212) <= not (a xor b);
    outputs(1213) <= a;
    outputs(1214) <= a;
    outputs(1215) <= a and not b;
    outputs(1216) <= not (a or b);
    outputs(1217) <= not (a xor b);
    outputs(1218) <= not (a xor b);
    outputs(1219) <= not (a or b);
    outputs(1220) <= a and not b;
    outputs(1221) <= not b;
    outputs(1222) <= not (a xor b);
    outputs(1223) <= not (a xor b);
    outputs(1224) <= a and b;
    outputs(1225) <= not a or b;
    outputs(1226) <= b;
    outputs(1227) <= a and b;
    outputs(1228) <= a;
    outputs(1229) <= a;
    outputs(1230) <= a and not b;
    outputs(1231) <= a xor b;
    outputs(1232) <= a and b;
    outputs(1233) <= a xor b;
    outputs(1234) <= a xor b;
    outputs(1235) <= b and not a;
    outputs(1236) <= b and not a;
    outputs(1237) <= b and not a;
    outputs(1238) <= a and b;
    outputs(1239) <= not b;
    outputs(1240) <= not a;
    outputs(1241) <= a;
    outputs(1242) <= not b;
    outputs(1243) <= a xor b;
    outputs(1244) <= a and b;
    outputs(1245) <= b and not a;
    outputs(1246) <= not b;
    outputs(1247) <= b;
    outputs(1248) <= a and not b;
    outputs(1249) <= not (a xor b);
    outputs(1250) <= b;
    outputs(1251) <= b and not a;
    outputs(1252) <= b and not a;
    outputs(1253) <= a and not b;
    outputs(1254) <= a xor b;
    outputs(1255) <= a and not b;
    outputs(1256) <= not (a or b);
    outputs(1257) <= not a or b;
    outputs(1258) <= not b;
    outputs(1259) <= b and not a;
    outputs(1260) <= a and not b;
    outputs(1261) <= a and b;
    outputs(1262) <= not (a or b);
    outputs(1263) <= not (a xor b);
    outputs(1264) <= not (a or b);
    outputs(1265) <= not (a xor b);
    outputs(1266) <= a and b;
    outputs(1267) <= not b;
    outputs(1268) <= 1'b0;
    outputs(1269) <= not (a or b);
    outputs(1270) <= a and b;
    outputs(1271) <= b and not a;
    outputs(1272) <= not (a or b);
    outputs(1273) <= not (a or b);
    outputs(1274) <= not b;
    outputs(1275) <= b and not a;
    outputs(1276) <= not a;
    outputs(1277) <= a;
    outputs(1278) <= b and not a;
    outputs(1279) <= not (a xor b);
    outputs(1280) <= not (a xor b);
    outputs(1281) <= b and not a;
    outputs(1282) <= a and b;
    outputs(1283) <= not (a xor b);
    outputs(1284) <= not (a or b);
    outputs(1285) <= a and not b;
    outputs(1286) <= not (a or b);
    outputs(1287) <= b and not a;
    outputs(1288) <= a and not b;
    outputs(1289) <= a;
    outputs(1290) <= a and b;
    outputs(1291) <= a and not b;
    outputs(1292) <= a and b;
    outputs(1293) <= a xor b;
    outputs(1294) <= a and not b;
    outputs(1295) <= not (a or b);
    outputs(1296) <= b and not a;
    outputs(1297) <= a and b;
    outputs(1298) <= a xor b;
    outputs(1299) <= a and b;
    outputs(1300) <= b and not a;
    outputs(1301) <= a and not b;
    outputs(1302) <= b and not a;
    outputs(1303) <= b and not a;
    outputs(1304) <= a xor b;
    outputs(1305) <= b;
    outputs(1306) <= not (a or b);
    outputs(1307) <= a xor b;
    outputs(1308) <= a and not b;
    outputs(1309) <= not b;
    outputs(1310) <= a and not b;
    outputs(1311) <= b and not a;
    outputs(1312) <= a and b;
    outputs(1313) <= a;
    outputs(1314) <= b and not a;
    outputs(1315) <= not b;
    outputs(1316) <= a and not b;
    outputs(1317) <= not (a or b);
    outputs(1318) <= b;
    outputs(1319) <= 1'b0;
    outputs(1320) <= b and not a;
    outputs(1321) <= not a;
    outputs(1322) <= 1'b0;
    outputs(1323) <= a and b;
    outputs(1324) <= not (a or b);
    outputs(1325) <= a and not b;
    outputs(1326) <= not b;
    outputs(1327) <= b and not a;
    outputs(1328) <= not (a or b);
    outputs(1329) <= a and not b;
    outputs(1330) <= not (a or b);
    outputs(1331) <= not (a xor b);
    outputs(1332) <= not (a xor b);
    outputs(1333) <= a and b;
    outputs(1334) <= a and not b;
    outputs(1335) <= a and not b;
    outputs(1336) <= b and not a;
    outputs(1337) <= not (a or b);
    outputs(1338) <= not (a xor b);
    outputs(1339) <= b and not a;
    outputs(1340) <= not (a or b);
    outputs(1341) <= a and not b;
    outputs(1342) <= b;
    outputs(1343) <= a and not b;
    outputs(1344) <= not (a xor b);
    outputs(1345) <= not a;
    outputs(1346) <= a;
    outputs(1347) <= a and b;
    outputs(1348) <= a and b;
    outputs(1349) <= not (a xor b);
    outputs(1350) <= not (a or b);
    outputs(1351) <= a and not b;
    outputs(1352) <= 1'b0;
    outputs(1353) <= b and not a;
    outputs(1354) <= a;
    outputs(1355) <= b and not a;
    outputs(1356) <= b and not a;
    outputs(1357) <= a and b;
    outputs(1358) <= a xor b;
    outputs(1359) <= a;
    outputs(1360) <= not a;
    outputs(1361) <= a xor b;
    outputs(1362) <= b and not a;
    outputs(1363) <= b and not a;
    outputs(1364) <= not (a xor b);
    outputs(1365) <= not a;
    outputs(1366) <= not (a xor b);
    outputs(1367) <= a and b;
    outputs(1368) <= b;
    outputs(1369) <= a and b;
    outputs(1370) <= a xor b;
    outputs(1371) <= a and b;
    outputs(1372) <= a xor b;
    outputs(1373) <= b and not a;
    outputs(1374) <= not b;
    outputs(1375) <= a and b;
    outputs(1376) <= not (a xor b);
    outputs(1377) <= not (a xor b);
    outputs(1378) <= b and not a;
    outputs(1379) <= b and not a;
    outputs(1380) <= not (a xor b);
    outputs(1381) <= a and not b;
    outputs(1382) <= a and b;
    outputs(1383) <= not (a or b);
    outputs(1384) <= a and not b;
    outputs(1385) <= a;
    outputs(1386) <= not (a or b);
    outputs(1387) <= b and not a;
    outputs(1388) <= a and b;
    outputs(1389) <= not (a or b);
    outputs(1390) <= not (a or b);
    outputs(1391) <= a xor b;
    outputs(1392) <= a and not b;
    outputs(1393) <= a and not b;
    outputs(1394) <= not (a or b);
    outputs(1395) <= b;
    outputs(1396) <= a;
    outputs(1397) <= not (a or b);
    outputs(1398) <= a;
    outputs(1399) <= a;
    outputs(1400) <= a and not b;
    outputs(1401) <= not (a xor b);
    outputs(1402) <= a and not b;
    outputs(1403) <= a and b;
    outputs(1404) <= b and not a;
    outputs(1405) <= a and not b;
    outputs(1406) <= not (a or b);
    outputs(1407) <= a and b;
    outputs(1408) <= b and not a;
    outputs(1409) <= not (a xor b);
    outputs(1410) <= a and b;
    outputs(1411) <= not a;
    outputs(1412) <= not (a or b);
    outputs(1413) <= not b;
    outputs(1414) <= a and b;
    outputs(1415) <= a and not b;
    outputs(1416) <= not (a or b);
    outputs(1417) <= not a;
    outputs(1418) <= b and not a;
    outputs(1419) <= a and b;
    outputs(1420) <= a and b;
    outputs(1421) <= a;
    outputs(1422) <= a and b;
    outputs(1423) <= a and b;
    outputs(1424) <= b and not a;
    outputs(1425) <= b and not a;
    outputs(1426) <= a and b;
    outputs(1427) <= a and b;
    outputs(1428) <= a xor b;
    outputs(1429) <= 1'b0;
    outputs(1430) <= b and not a;
    outputs(1431) <= a and not b;
    outputs(1432) <= a and not b;
    outputs(1433) <= a;
    outputs(1434) <= 1'b0;
    outputs(1435) <= a and b;
    outputs(1436) <= b and not a;
    outputs(1437) <= a and b;
    outputs(1438) <= b;
    outputs(1439) <= b and not a;
    outputs(1440) <= not (a or b);
    outputs(1441) <= a and not b;
    outputs(1442) <= a and not b;
    outputs(1443) <= a and b;
    outputs(1444) <= not (a or b);
    outputs(1445) <= a xor b;
    outputs(1446) <= a and b;
    outputs(1447) <= a and b;
    outputs(1448) <= a and not b;
    outputs(1449) <= b and not a;
    outputs(1450) <= not (a xor b);
    outputs(1451) <= not (a xor b);
    outputs(1452) <= b;
    outputs(1453) <= a and not b;
    outputs(1454) <= a xor b;
    outputs(1455) <= not a;
    outputs(1456) <= 1'b0;
    outputs(1457) <= a and b;
    outputs(1458) <= b;
    outputs(1459) <= a;
    outputs(1460) <= 1'b0;
    outputs(1461) <= a and b;
    outputs(1462) <= a and not b;
    outputs(1463) <= a and b;
    outputs(1464) <= a and not b;
    outputs(1465) <= b and not a;
    outputs(1466) <= a and b;
    outputs(1467) <= b and not a;
    outputs(1468) <= not b;
    outputs(1469) <= not (a xor b);
    outputs(1470) <= not a;
    outputs(1471) <= b and not a;
    outputs(1472) <= b and not a;
    outputs(1473) <= a or b;
    outputs(1474) <= not (a xor b);
    outputs(1475) <= b and not a;
    outputs(1476) <= 1'b0;
    outputs(1477) <= not (a or b);
    outputs(1478) <= not b;
    outputs(1479) <= not a;
    outputs(1480) <= not (a or b);
    outputs(1481) <= a and not b;
    outputs(1482) <= a xor b;
    outputs(1483) <= a and b;
    outputs(1484) <= a and not b;
    outputs(1485) <= b and not a;
    outputs(1486) <= not (a or b);
    outputs(1487) <= a and not b;
    outputs(1488) <= a and b;
    outputs(1489) <= not (a or b);
    outputs(1490) <= not b;
    outputs(1491) <= not (a or b);
    outputs(1492) <= not (a or b);
    outputs(1493) <= a and not b;
    outputs(1494) <= b and not a;
    outputs(1495) <= a and b;
    outputs(1496) <= b and not a;
    outputs(1497) <= not (a xor b);
    outputs(1498) <= a and b;
    outputs(1499) <= b;
    outputs(1500) <= a and b;
    outputs(1501) <= b and not a;
    outputs(1502) <= a and not b;
    outputs(1503) <= not a;
    outputs(1504) <= a and b;
    outputs(1505) <= a and not b;
    outputs(1506) <= a and b;
    outputs(1507) <= b;
    outputs(1508) <= a and b;
    outputs(1509) <= not (a xor b);
    outputs(1510) <= a and b;
    outputs(1511) <= not (a or b);
    outputs(1512) <= a and not b;
    outputs(1513) <= a and b;
    outputs(1514) <= b and not a;
    outputs(1515) <= not a;
    outputs(1516) <= a;
    outputs(1517) <= b;
    outputs(1518) <= not a;
    outputs(1519) <= not a;
    outputs(1520) <= a and not b;
    outputs(1521) <= a and not b;
    outputs(1522) <= not (a xor b);
    outputs(1523) <= not b;
    outputs(1524) <= a and not b;
    outputs(1525) <= not (a or b);
    outputs(1526) <= not (a or b);
    outputs(1527) <= a and not b;
    outputs(1528) <= b and not a;
    outputs(1529) <= b and not a;
    outputs(1530) <= b;
    outputs(1531) <= b;
    outputs(1532) <= a;
    outputs(1533) <= not a;
    outputs(1534) <= not (a or b);
    outputs(1535) <= a and not b;
    outputs(1536) <= not (a or b);
    outputs(1537) <= 1'b1;
    outputs(1538) <= a;
    outputs(1539) <= a xor b;
    outputs(1540) <= not b;
    outputs(1541) <= not b or a;
    outputs(1542) <= not a or b;
    outputs(1543) <= not a;
    outputs(1544) <= not (a or b);
    outputs(1545) <= b and not a;
    outputs(1546) <= b;
    outputs(1547) <= not b or a;
    outputs(1548) <= not (a xor b);
    outputs(1549) <= not a or b;
    outputs(1550) <= b;
    outputs(1551) <= not (a xor b);
    outputs(1552) <= b;
    outputs(1553) <= not b;
    outputs(1554) <= a and not b;
    outputs(1555) <= b;
    outputs(1556) <= not (a or b);
    outputs(1557) <= a xor b;
    outputs(1558) <= not (a or b);
    outputs(1559) <= b and not a;
    outputs(1560) <= a;
    outputs(1561) <= not b or a;
    outputs(1562) <= not b or a;
    outputs(1563) <= not (a and b);
    outputs(1564) <= not (a or b);
    outputs(1565) <= not a or b;
    outputs(1566) <= not a;
    outputs(1567) <= b and not a;
    outputs(1568) <= not b;
    outputs(1569) <= not b or a;
    outputs(1570) <= a and not b;
    outputs(1571) <= b;
    outputs(1572) <= not b;
    outputs(1573) <= b;
    outputs(1574) <= a;
    outputs(1575) <= a and b;
    outputs(1576) <= a xor b;
    outputs(1577) <= b;
    outputs(1578) <= not b;
    outputs(1579) <= a or b;
    outputs(1580) <= not a or b;
    outputs(1581) <= a xor b;
    outputs(1582) <= not a;
    outputs(1583) <= a xor b;
    outputs(1584) <= b;
    outputs(1585) <= a;
    outputs(1586) <= b;
    outputs(1587) <= not (a and b);
    outputs(1588) <= not (a and b);
    outputs(1589) <= b;
    outputs(1590) <= not a;
    outputs(1591) <= not (a or b);
    outputs(1592) <= a;
    outputs(1593) <= not b;
    outputs(1594) <= not (a and b);
    outputs(1595) <= a and not b;
    outputs(1596) <= not (a xor b);
    outputs(1597) <= a or b;
    outputs(1598) <= not b;
    outputs(1599) <= b;
    outputs(1600) <= a;
    outputs(1601) <= a or b;
    outputs(1602) <= not b;
    outputs(1603) <= not b or a;
    outputs(1604) <= not a or b;
    outputs(1605) <= not (a xor b);
    outputs(1606) <= b and not a;
    outputs(1607) <= a xor b;
    outputs(1608) <= not (a xor b);
    outputs(1609) <= a;
    outputs(1610) <= a;
    outputs(1611) <= a xor b;
    outputs(1612) <= b and not a;
    outputs(1613) <= not a or b;
    outputs(1614) <= not b or a;
    outputs(1615) <= not a;
    outputs(1616) <= a;
    outputs(1617) <= not (a xor b);
    outputs(1618) <= a xor b;
    outputs(1619) <= a;
    outputs(1620) <= a xor b;
    outputs(1621) <= not a or b;
    outputs(1622) <= not (a or b);
    outputs(1623) <= not a;
    outputs(1624) <= a xor b;
    outputs(1625) <= a xor b;
    outputs(1626) <= not (a xor b);
    outputs(1627) <= b;
    outputs(1628) <= not (a or b);
    outputs(1629) <= a and b;
    outputs(1630) <= a;
    outputs(1631) <= b and not a;
    outputs(1632) <= a;
    outputs(1633) <= a and not b;
    outputs(1634) <= a or b;
    outputs(1635) <= not (a and b);
    outputs(1636) <= not b;
    outputs(1637) <= not (a xor b);
    outputs(1638) <= not (a xor b);
    outputs(1639) <= not (a and b);
    outputs(1640) <= a xor b;
    outputs(1641) <= b and not a;
    outputs(1642) <= a and b;
    outputs(1643) <= not (a and b);
    outputs(1644) <= a;
    outputs(1645) <= b;
    outputs(1646) <= not (a or b);
    outputs(1647) <= a and b;
    outputs(1648) <= a xor b;
    outputs(1649) <= b;
    outputs(1650) <= a or b;
    outputs(1651) <= a xor b;
    outputs(1652) <= a and b;
    outputs(1653) <= not (a and b);
    outputs(1654) <= a and not b;
    outputs(1655) <= not a;
    outputs(1656) <= a xor b;
    outputs(1657) <= not (a and b);
    outputs(1658) <= not b;
    outputs(1659) <= a and not b;
    outputs(1660) <= a xor b;
    outputs(1661) <= not (a xor b);
    outputs(1662) <= not a;
    outputs(1663) <= a xor b;
    outputs(1664) <= not a;
    outputs(1665) <= not (a xor b);
    outputs(1666) <= not b or a;
    outputs(1667) <= not a;
    outputs(1668) <= not (a xor b);
    outputs(1669) <= b;
    outputs(1670) <= not a;
    outputs(1671) <= not (a xor b);
    outputs(1672) <= not a;
    outputs(1673) <= not b;
    outputs(1674) <= a xor b;
    outputs(1675) <= a and not b;
    outputs(1676) <= not b;
    outputs(1677) <= not a or b;
    outputs(1678) <= a;
    outputs(1679) <= b;
    outputs(1680) <= not a;
    outputs(1681) <= a xor b;
    outputs(1682) <= a;
    outputs(1683) <= b;
    outputs(1684) <= a;
    outputs(1685) <= not (a and b);
    outputs(1686) <= not (a xor b);
    outputs(1687) <= a xor b;
    outputs(1688) <= not (a xor b);
    outputs(1689) <= not a;
    outputs(1690) <= not a;
    outputs(1691) <= not (a or b);
    outputs(1692) <= not (a or b);
    outputs(1693) <= a and b;
    outputs(1694) <= not a or b;
    outputs(1695) <= not (a and b);
    outputs(1696) <= b;
    outputs(1697) <= not a;
    outputs(1698) <= not b;
    outputs(1699) <= not a;
    outputs(1700) <= not a;
    outputs(1701) <= a xor b;
    outputs(1702) <= a;
    outputs(1703) <= a xor b;
    outputs(1704) <= a or b;
    outputs(1705) <= a;
    outputs(1706) <= b;
    outputs(1707) <= not b;
    outputs(1708) <= not (a xor b);
    outputs(1709) <= not a;
    outputs(1710) <= b;
    outputs(1711) <= not a or b;
    outputs(1712) <= a;
    outputs(1713) <= not a;
    outputs(1714) <= b;
    outputs(1715) <= not a or b;
    outputs(1716) <= a;
    outputs(1717) <= a;
    outputs(1718) <= not b or a;
    outputs(1719) <= b;
    outputs(1720) <= a and b;
    outputs(1721) <= a or b;
    outputs(1722) <= not (a xor b);
    outputs(1723) <= a;
    outputs(1724) <= a or b;
    outputs(1725) <= a;
    outputs(1726) <= not a;
    outputs(1727) <= a and not b;
    outputs(1728) <= a or b;
    outputs(1729) <= a and b;
    outputs(1730) <= not b or a;
    outputs(1731) <= a and b;
    outputs(1732) <= not (a xor b);
    outputs(1733) <= not b;
    outputs(1734) <= not b;
    outputs(1735) <= not b or a;
    outputs(1736) <= a;
    outputs(1737) <= not a;
    outputs(1738) <= a;
    outputs(1739) <= not a or b;
    outputs(1740) <= not b;
    outputs(1741) <= a;
    outputs(1742) <= not (a xor b);
    outputs(1743) <= a;
    outputs(1744) <= not b;
    outputs(1745) <= a xor b;
    outputs(1746) <= not b or a;
    outputs(1747) <= a and b;
    outputs(1748) <= not a or b;
    outputs(1749) <= not (a or b);
    outputs(1750) <= not (a xor b);
    outputs(1751) <= a;
    outputs(1752) <= b and not a;
    outputs(1753) <= not (a and b);
    outputs(1754) <= not a or b;
    outputs(1755) <= not a or b;
    outputs(1756) <= not a or b;
    outputs(1757) <= not (a xor b);
    outputs(1758) <= b;
    outputs(1759) <= not (a and b);
    outputs(1760) <= not (a xor b);
    outputs(1761) <= a and not b;
    outputs(1762) <= not (a xor b);
    outputs(1763) <= not b or a;
    outputs(1764) <= a or b;
    outputs(1765) <= not b;
    outputs(1766) <= b;
    outputs(1767) <= a xor b;
    outputs(1768) <= not b or a;
    outputs(1769) <= not b;
    outputs(1770) <= not b or a;
    outputs(1771) <= not a or b;
    outputs(1772) <= not b;
    outputs(1773) <= a or b;
    outputs(1774) <= not (a xor b);
    outputs(1775) <= not a;
    outputs(1776) <= a and not b;
    outputs(1777) <= a and not b;
    outputs(1778) <= a;
    outputs(1779) <= not b or a;
    outputs(1780) <= a or b;
    outputs(1781) <= not b or a;
    outputs(1782) <= a or b;
    outputs(1783) <= a and b;
    outputs(1784) <= b;
    outputs(1785) <= not b;
    outputs(1786) <= a and not b;
    outputs(1787) <= a xor b;
    outputs(1788) <= a;
    outputs(1789) <= b;
    outputs(1790) <= not b;
    outputs(1791) <= a and not b;
    outputs(1792) <= b;
    outputs(1793) <= not (a or b);
    outputs(1794) <= a;
    outputs(1795) <= b;
    outputs(1796) <= a and not b;
    outputs(1797) <= not a or b;
    outputs(1798) <= not a or b;
    outputs(1799) <= b;
    outputs(1800) <= not b;
    outputs(1801) <= b;
    outputs(1802) <= not a;
    outputs(1803) <= not a;
    outputs(1804) <= a and b;
    outputs(1805) <= not a;
    outputs(1806) <= not (a xor b);
    outputs(1807) <= not a;
    outputs(1808) <= not a;
    outputs(1809) <= not (a or b);
    outputs(1810) <= b and not a;
    outputs(1811) <= b;
    outputs(1812) <= not b or a;
    outputs(1813) <= a xor b;
    outputs(1814) <= a and not b;
    outputs(1815) <= not b;
    outputs(1816) <= a and b;
    outputs(1817) <= b;
    outputs(1818) <= a xor b;
    outputs(1819) <= a;
    outputs(1820) <= a and b;
    outputs(1821) <= not a;
    outputs(1822) <= not a;
    outputs(1823) <= not a;
    outputs(1824) <= not a;
    outputs(1825) <= not (a xor b);
    outputs(1826) <= a or b;
    outputs(1827) <= a xor b;
    outputs(1828) <= not b;
    outputs(1829) <= a xor b;
    outputs(1830) <= b and not a;
    outputs(1831) <= a;
    outputs(1832) <= not a;
    outputs(1833) <= not (a or b);
    outputs(1834) <= not b or a;
    outputs(1835) <= not (a xor b);
    outputs(1836) <= b;
    outputs(1837) <= b;
    outputs(1838) <= not (a xor b);
    outputs(1839) <= not b;
    outputs(1840) <= not (a and b);
    outputs(1841) <= not (a or b);
    outputs(1842) <= a;
    outputs(1843) <= b;
    outputs(1844) <= not (a or b);
    outputs(1845) <= b;
    outputs(1846) <= a;
    outputs(1847) <= not (a or b);
    outputs(1848) <= not a;
    outputs(1849) <= not (a and b);
    outputs(1850) <= not (a or b);
    outputs(1851) <= a xor b;
    outputs(1852) <= not b;
    outputs(1853) <= not (a or b);
    outputs(1854) <= b;
    outputs(1855) <= b;
    outputs(1856) <= not a;
    outputs(1857) <= not (a or b);
    outputs(1858) <= a;
    outputs(1859) <= a;
    outputs(1860) <= a;
    outputs(1861) <= not a;
    outputs(1862) <= not a;
    outputs(1863) <= not (a and b);
    outputs(1864) <= not b;
    outputs(1865) <= a or b;
    outputs(1866) <= a xor b;
    outputs(1867) <= a and not b;
    outputs(1868) <= not (a or b);
    outputs(1869) <= a and b;
    outputs(1870) <= a;
    outputs(1871) <= not a or b;
    outputs(1872) <= a;
    outputs(1873) <= b;
    outputs(1874) <= not (a xor b);
    outputs(1875) <= a and not b;
    outputs(1876) <= not b;
    outputs(1877) <= a or b;
    outputs(1878) <= a xor b;
    outputs(1879) <= a;
    outputs(1880) <= not b or a;
    outputs(1881) <= not (a xor b);
    outputs(1882) <= b;
    outputs(1883) <= not b;
    outputs(1884) <= a or b;
    outputs(1885) <= not (a and b);
    outputs(1886) <= not (a and b);
    outputs(1887) <= b and not a;
    outputs(1888) <= not (a and b);
    outputs(1889) <= not (a xor b);
    outputs(1890) <= a xor b;
    outputs(1891) <= not a;
    outputs(1892) <= b and not a;
    outputs(1893) <= not (a xor b);
    outputs(1894) <= a xor b;
    outputs(1895) <= not (a and b);
    outputs(1896) <= not a;
    outputs(1897) <= not (a and b);
    outputs(1898) <= a xor b;
    outputs(1899) <= not (a xor b);
    outputs(1900) <= a and not b;
    outputs(1901) <= a or b;
    outputs(1902) <= a or b;
    outputs(1903) <= b;
    outputs(1904) <= not a or b;
    outputs(1905) <= b;
    outputs(1906) <= not (a xor b);
    outputs(1907) <= a and not b;
    outputs(1908) <= not b or a;
    outputs(1909) <= not (a and b);
    outputs(1910) <= not b;
    outputs(1911) <= not a;
    outputs(1912) <= a;
    outputs(1913) <= not a;
    outputs(1914) <= b and not a;
    outputs(1915) <= not a;
    outputs(1916) <= a xor b;
    outputs(1917) <= b and not a;
    outputs(1918) <= not (a and b);
    outputs(1919) <= not (a or b);
    outputs(1920) <= b;
    outputs(1921) <= not a or b;
    outputs(1922) <= a or b;
    outputs(1923) <= b and not a;
    outputs(1924) <= not b or a;
    outputs(1925) <= not a;
    outputs(1926) <= b;
    outputs(1927) <= not a or b;
    outputs(1928) <= a or b;
    outputs(1929) <= a or b;
    outputs(1930) <= a and not b;
    outputs(1931) <= a xor b;
    outputs(1932) <= b;
    outputs(1933) <= a;
    outputs(1934) <= not b;
    outputs(1935) <= not (a or b);
    outputs(1936) <= b and not a;
    outputs(1937) <= not a;
    outputs(1938) <= a and not b;
    outputs(1939) <= not b;
    outputs(1940) <= not a;
    outputs(1941) <= a and b;
    outputs(1942) <= not b;
    outputs(1943) <= not a or b;
    outputs(1944) <= not b;
    outputs(1945) <= a or b;
    outputs(1946) <= a xor b;
    outputs(1947) <= not (a xor b);
    outputs(1948) <= not a;
    outputs(1949) <= not (a xor b);
    outputs(1950) <= a or b;
    outputs(1951) <= not (a or b);
    outputs(1952) <= not a;
    outputs(1953) <= a and b;
    outputs(1954) <= not (a and b);
    outputs(1955) <= b and not a;
    outputs(1956) <= a;
    outputs(1957) <= not (a or b);
    outputs(1958) <= b and not a;
    outputs(1959) <= not b;
    outputs(1960) <= not (a and b);
    outputs(1961) <= not b or a;
    outputs(1962) <= a or b;
    outputs(1963) <= a and b;
    outputs(1964) <= not (a xor b);
    outputs(1965) <= b;
    outputs(1966) <= not (a xor b);
    outputs(1967) <= not (a or b);
    outputs(1968) <= a;
    outputs(1969) <= a;
    outputs(1970) <= a;
    outputs(1971) <= not (a or b);
    outputs(1972) <= a or b;
    outputs(1973) <= a and b;
    outputs(1974) <= a or b;
    outputs(1975) <= a;
    outputs(1976) <= b and not a;
    outputs(1977) <= a or b;
    outputs(1978) <= not b;
    outputs(1979) <= b;
    outputs(1980) <= not (a and b);
    outputs(1981) <= b and not a;
    outputs(1982) <= not b;
    outputs(1983) <= not a or b;
    outputs(1984) <= a xor b;
    outputs(1985) <= not b or a;
    outputs(1986) <= a or b;
    outputs(1987) <= a;
    outputs(1988) <= not b or a;
    outputs(1989) <= b;
    outputs(1990) <= a or b;
    outputs(1991) <= a;
    outputs(1992) <= not (a xor b);
    outputs(1993) <= a xor b;
    outputs(1994) <= not (a xor b);
    outputs(1995) <= not a;
    outputs(1996) <= not (a and b);
    outputs(1997) <= a or b;
    outputs(1998) <= not (a xor b);
    outputs(1999) <= not a;
    outputs(2000) <= a and b;
    outputs(2001) <= not b;
    outputs(2002) <= not (a xor b);
    outputs(2003) <= a or b;
    outputs(2004) <= a;
    outputs(2005) <= b and not a;
    outputs(2006) <= a and b;
    outputs(2007) <= not (a and b);
    outputs(2008) <= a;
    outputs(2009) <= not a;
    outputs(2010) <= a xor b;
    outputs(2011) <= not (a xor b);
    outputs(2012) <= b and not a;
    outputs(2013) <= not a;
    outputs(2014) <= not (a xor b);
    outputs(2015) <= not b;
    outputs(2016) <= not b;
    outputs(2017) <= not a;
    outputs(2018) <= not (a or b);
    outputs(2019) <= not (a xor b);
    outputs(2020) <= not (a or b);
    outputs(2021) <= not a;
    outputs(2022) <= a and not b;
    outputs(2023) <= a xor b;
    outputs(2024) <= a and not b;
    outputs(2025) <= not b or a;
    outputs(2026) <= b;
    outputs(2027) <= not (a xor b);
    outputs(2028) <= a xor b;
    outputs(2029) <= b and not a;
    outputs(2030) <= b;
    outputs(2031) <= not b;
    outputs(2032) <= a;
    outputs(2033) <= a and not b;
    outputs(2034) <= not a;
    outputs(2035) <= a;
    outputs(2036) <= a and not b;
    outputs(2037) <= b;
    outputs(2038) <= a xor b;
    outputs(2039) <= not a or b;
    outputs(2040) <= b and not a;
    outputs(2041) <= not a;
    outputs(2042) <= b and not a;
    outputs(2043) <= not b;
    outputs(2044) <= a and not b;
    outputs(2045) <= a xor b;
    outputs(2046) <= not b or a;
    outputs(2047) <= a and not b;
    outputs(2048) <= a;
    outputs(2049) <= not a;
    outputs(2050) <= not (a and b);
    outputs(2051) <= a;
    outputs(2052) <= not b;
    outputs(2053) <= not b;
    outputs(2054) <= not b;
    outputs(2055) <= not a;
    outputs(2056) <= not a;
    outputs(2057) <= not b;
    outputs(2058) <= not (a and b);
    outputs(2059) <= b;
    outputs(2060) <= a;
    outputs(2061) <= b and not a;
    outputs(2062) <= a xor b;
    outputs(2063) <= not (a xor b);
    outputs(2064) <= not (a and b);
    outputs(2065) <= not a or b;
    outputs(2066) <= not (a or b);
    outputs(2067) <= not a or b;
    outputs(2068) <= a and b;
    outputs(2069) <= not (a xor b);
    outputs(2070) <= a xor b;
    outputs(2071) <= b and not a;
    outputs(2072) <= a;
    outputs(2073) <= not b;
    outputs(2074) <= b and not a;
    outputs(2075) <= a or b;
    outputs(2076) <= b and not a;
    outputs(2077) <= not (a xor b);
    outputs(2078) <= not a or b;
    outputs(2079) <= b and not a;
    outputs(2080) <= not b or a;
    outputs(2081) <= a;
    outputs(2082) <= a and not b;
    outputs(2083) <= a and not b;
    outputs(2084) <= b and not a;
    outputs(2085) <= not b;
    outputs(2086) <= not a or b;
    outputs(2087) <= a or b;
    outputs(2088) <= not (a or b);
    outputs(2089) <= a;
    outputs(2090) <= a and not b;
    outputs(2091) <= not (a and b);
    outputs(2092) <= not b;
    outputs(2093) <= b;
    outputs(2094) <= not (a and b);
    outputs(2095) <= a and not b;
    outputs(2096) <= not (a xor b);
    outputs(2097) <= a or b;
    outputs(2098) <= b;
    outputs(2099) <= not a or b;
    outputs(2100) <= not b;
    outputs(2101) <= not b or a;
    outputs(2102) <= a;
    outputs(2103) <= b and not a;
    outputs(2104) <= a xor b;
    outputs(2105) <= b;
    outputs(2106) <= not b or a;
    outputs(2107) <= not b or a;
    outputs(2108) <= not b;
    outputs(2109) <= b;
    outputs(2110) <= a xor b;
    outputs(2111) <= a or b;
    outputs(2112) <= b and not a;
    outputs(2113) <= not a;
    outputs(2114) <= not (a and b);
    outputs(2115) <= b and not a;
    outputs(2116) <= not b;
    outputs(2117) <= not (a or b);
    outputs(2118) <= a and b;
    outputs(2119) <= a xor b;
    outputs(2120) <= b and not a;
    outputs(2121) <= not (a xor b);
    outputs(2122) <= not a or b;
    outputs(2123) <= not a;
    outputs(2124) <= not (a and b);
    outputs(2125) <= not b;
    outputs(2126) <= not (a and b);
    outputs(2127) <= not (a xor b);
    outputs(2128) <= not b or a;
    outputs(2129) <= not (a and b);
    outputs(2130) <= a xor b;
    outputs(2131) <= a and b;
    outputs(2132) <= b;
    outputs(2133) <= not b;
    outputs(2134) <= not b;
    outputs(2135) <= a or b;
    outputs(2136) <= not (a xor b);
    outputs(2137) <= a;
    outputs(2138) <= a xor b;
    outputs(2139) <= not a;
    outputs(2140) <= not (a xor b);
    outputs(2141) <= not a or b;
    outputs(2142) <= a;
    outputs(2143) <= not (a xor b);
    outputs(2144) <= not (a xor b);
    outputs(2145) <= not (a xor b);
    outputs(2146) <= not a;
    outputs(2147) <= a and not b;
    outputs(2148) <= a and b;
    outputs(2149) <= b;
    outputs(2150) <= not b;
    outputs(2151) <= a or b;
    outputs(2152) <= a or b;
    outputs(2153) <= a or b;
    outputs(2154) <= a xor b;
    outputs(2155) <= a or b;
    outputs(2156) <= not (a xor b);
    outputs(2157) <= a xor b;
    outputs(2158) <= not b or a;
    outputs(2159) <= a and b;
    outputs(2160) <= not (a xor b);
    outputs(2161) <= not b;
    outputs(2162) <= a xor b;
    outputs(2163) <= a xor b;
    outputs(2164) <= b;
    outputs(2165) <= not (a and b);
    outputs(2166) <= not a;
    outputs(2167) <= not b;
    outputs(2168) <= not (a and b);
    outputs(2169) <= b;
    outputs(2170) <= not (a xor b);
    outputs(2171) <= not (a and b);
    outputs(2172) <= b;
    outputs(2173) <= not (a xor b);
    outputs(2174) <= a and b;
    outputs(2175) <= a and not b;
    outputs(2176) <= not a;
    outputs(2177) <= a;
    outputs(2178) <= a;
    outputs(2179) <= not a or b;
    outputs(2180) <= not (a xor b);
    outputs(2181) <= not (a or b);
    outputs(2182) <= a or b;
    outputs(2183) <= a;
    outputs(2184) <= not b;
    outputs(2185) <= not a;
    outputs(2186) <= a or b;
    outputs(2187) <= not a or b;
    outputs(2188) <= not a;
    outputs(2189) <= not b;
    outputs(2190) <= a and not b;
    outputs(2191) <= b;
    outputs(2192) <= not b or a;
    outputs(2193) <= not a;
    outputs(2194) <= not (a xor b);
    outputs(2195) <= a or b;
    outputs(2196) <= not (a xor b);
    outputs(2197) <= a or b;
    outputs(2198) <= b and not a;
    outputs(2199) <= b;
    outputs(2200) <= a and not b;
    outputs(2201) <= not a;
    outputs(2202) <= not a;
    outputs(2203) <= not (a xor b);
    outputs(2204) <= not (a xor b);
    outputs(2205) <= a xor b;
    outputs(2206) <= not (a xor b);
    outputs(2207) <= b;
    outputs(2208) <= a;
    outputs(2209) <= not (a xor b);
    outputs(2210) <= not a or b;
    outputs(2211) <= not a or b;
    outputs(2212) <= not b;
    outputs(2213) <= not (a xor b);
    outputs(2214) <= not a;
    outputs(2215) <= a xor b;
    outputs(2216) <= not a;
    outputs(2217) <= not (a or b);
    outputs(2218) <= a xor b;
    outputs(2219) <= not a;
    outputs(2220) <= a;
    outputs(2221) <= a or b;
    outputs(2222) <= not a;
    outputs(2223) <= not b;
    outputs(2224) <= not a or b;
    outputs(2225) <= b;
    outputs(2226) <= not (a xor b);
    outputs(2227) <= not b or a;
    outputs(2228) <= a;
    outputs(2229) <= not b;
    outputs(2230) <= not a;
    outputs(2231) <= b and not a;
    outputs(2232) <= a xor b;
    outputs(2233) <= not b;
    outputs(2234) <= a and not b;
    outputs(2235) <= a xor b;
    outputs(2236) <= not a;
    outputs(2237) <= a;
    outputs(2238) <= not (a xor b);
    outputs(2239) <= not a;
    outputs(2240) <= not a;
    outputs(2241) <= a and b;
    outputs(2242) <= not b;
    outputs(2243) <= not a;
    outputs(2244) <= a xor b;
    outputs(2245) <= a and not b;
    outputs(2246) <= not (a and b);
    outputs(2247) <= not a;
    outputs(2248) <= not a or b;
    outputs(2249) <= a xor b;
    outputs(2250) <= b;
    outputs(2251) <= a;
    outputs(2252) <= a xor b;
    outputs(2253) <= not a or b;
    outputs(2254) <= not a;
    outputs(2255) <= a;
    outputs(2256) <= a and not b;
    outputs(2257) <= not b;
    outputs(2258) <= a;
    outputs(2259) <= a xor b;
    outputs(2260) <= not (a xor b);
    outputs(2261) <= not (a xor b);
    outputs(2262) <= b;
    outputs(2263) <= not a or b;
    outputs(2264) <= not a;
    outputs(2265) <= a;
    outputs(2266) <= b and not a;
    outputs(2267) <= not b;
    outputs(2268) <= a xor b;
    outputs(2269) <= a or b;
    outputs(2270) <= not a or b;
    outputs(2271) <= not b;
    outputs(2272) <= not (a xor b);
    outputs(2273) <= not a;
    outputs(2274) <= a or b;
    outputs(2275) <= not (a and b);
    outputs(2276) <= not (a or b);
    outputs(2277) <= a xor b;
    outputs(2278) <= a xor b;
    outputs(2279) <= not b;
    outputs(2280) <= a and b;
    outputs(2281) <= not (a xor b);
    outputs(2282) <= a and not b;
    outputs(2283) <= not b;
    outputs(2284) <= not b or a;
    outputs(2285) <= a and not b;
    outputs(2286) <= not (a or b);
    outputs(2287) <= b and not a;
    outputs(2288) <= not b or a;
    outputs(2289) <= not (a or b);
    outputs(2290) <= a xor b;
    outputs(2291) <= not (a and b);
    outputs(2292) <= b;
    outputs(2293) <= not (a xor b);
    outputs(2294) <= not (a xor b);
    outputs(2295) <= a xor b;
    outputs(2296) <= not a;
    outputs(2297) <= a or b;
    outputs(2298) <= not b;
    outputs(2299) <= a;
    outputs(2300) <= not (a or b);
    outputs(2301) <= b;
    outputs(2302) <= not b;
    outputs(2303) <= a or b;
    outputs(2304) <= not a;
    outputs(2305) <= b and not a;
    outputs(2306) <= not a;
    outputs(2307) <= b;
    outputs(2308) <= a and not b;
    outputs(2309) <= not b or a;
    outputs(2310) <= not b;
    outputs(2311) <= a;
    outputs(2312) <= a and b;
    outputs(2313) <= not a;
    outputs(2314) <= a or b;
    outputs(2315) <= a;
    outputs(2316) <= not b or a;
    outputs(2317) <= not b or a;
    outputs(2318) <= not (a xor b);
    outputs(2319) <= b and not a;
    outputs(2320) <= a and b;
    outputs(2321) <= not (a xor b);
    outputs(2322) <= not a or b;
    outputs(2323) <= b and not a;
    outputs(2324) <= not (a xor b);
    outputs(2325) <= a and not b;
    outputs(2326) <= a or b;
    outputs(2327) <= not (a xor b);
    outputs(2328) <= a or b;
    outputs(2329) <= not (a or b);
    outputs(2330) <= not b;
    outputs(2331) <= not a or b;
    outputs(2332) <= b and not a;
    outputs(2333) <= not b or a;
    outputs(2334) <= not b;
    outputs(2335) <= not a;
    outputs(2336) <= a and not b;
    outputs(2337) <= not (a xor b);
    outputs(2338) <= b and not a;
    outputs(2339) <= b and not a;
    outputs(2340) <= not b;
    outputs(2341) <= b;
    outputs(2342) <= a and not b;
    outputs(2343) <= b and not a;
    outputs(2344) <= not a or b;
    outputs(2345) <= a and not b;
    outputs(2346) <= not a or b;
    outputs(2347) <= not (a and b);
    outputs(2348) <= a xor b;
    outputs(2349) <= not b or a;
    outputs(2350) <= a xor b;
    outputs(2351) <= not (a xor b);
    outputs(2352) <= a and not b;
    outputs(2353) <= b and not a;
    outputs(2354) <= a and not b;
    outputs(2355) <= a;
    outputs(2356) <= a;
    outputs(2357) <= b;
    outputs(2358) <= a and b;
    outputs(2359) <= a;
    outputs(2360) <= not b;
    outputs(2361) <= not b;
    outputs(2362) <= not a or b;
    outputs(2363) <= not (a xor b);
    outputs(2364) <= not (a and b);
    outputs(2365) <= b and not a;
    outputs(2366) <= a xor b;
    outputs(2367) <= not (a and b);
    outputs(2368) <= b;
    outputs(2369) <= a and not b;
    outputs(2370) <= not (a xor b);
    outputs(2371) <= not (a and b);
    outputs(2372) <= not b;
    outputs(2373) <= a and b;
    outputs(2374) <= b;
    outputs(2375) <= not a;
    outputs(2376) <= b;
    outputs(2377) <= a and not b;
    outputs(2378) <= not b or a;
    outputs(2379) <= b;
    outputs(2380) <= b;
    outputs(2381) <= not a;
    outputs(2382) <= a and b;
    outputs(2383) <= not (a or b);
    outputs(2384) <= a and b;
    outputs(2385) <= not a;
    outputs(2386) <= a or b;
    outputs(2387) <= a or b;
    outputs(2388) <= a xor b;
    outputs(2389) <= not b;
    outputs(2390) <= b;
    outputs(2391) <= not b or a;
    outputs(2392) <= a xor b;
    outputs(2393) <= not b;
    outputs(2394) <= not b;
    outputs(2395) <= not (a xor b);
    outputs(2396) <= a xor b;
    outputs(2397) <= a and not b;
    outputs(2398) <= not b;
    outputs(2399) <= b and not a;
    outputs(2400) <= a xor b;
    outputs(2401) <= not b;
    outputs(2402) <= a;
    outputs(2403) <= not a;
    outputs(2404) <= not b or a;
    outputs(2405) <= not a;
    outputs(2406) <= not a or b;
    outputs(2407) <= not a or b;
    outputs(2408) <= not (a and b);
    outputs(2409) <= b;
    outputs(2410) <= not b;
    outputs(2411) <= a xor b;
    outputs(2412) <= a and not b;
    outputs(2413) <= a xor b;
    outputs(2414) <= not a;
    outputs(2415) <= b;
    outputs(2416) <= a xor b;
    outputs(2417) <= not a;
    outputs(2418) <= a;
    outputs(2419) <= not b or a;
    outputs(2420) <= not b;
    outputs(2421) <= not a;
    outputs(2422) <= a and b;
    outputs(2423) <= b and not a;
    outputs(2424) <= not b or a;
    outputs(2425) <= a and b;
    outputs(2426) <= not (a and b);
    outputs(2427) <= not (a and b);
    outputs(2428) <= not (a xor b);
    outputs(2429) <= not a;
    outputs(2430) <= b and not a;
    outputs(2431) <= not b;
    outputs(2432) <= a xor b;
    outputs(2433) <= not (a xor b);
    outputs(2434) <= not (a xor b);
    outputs(2435) <= not (a xor b);
    outputs(2436) <= a xor b;
    outputs(2437) <= not a;
    outputs(2438) <= not a;
    outputs(2439) <= a;
    outputs(2440) <= a xor b;
    outputs(2441) <= a xor b;
    outputs(2442) <= not a;
    outputs(2443) <= a;
    outputs(2444) <= not (a xor b);
    outputs(2445) <= not a or b;
    outputs(2446) <= not b or a;
    outputs(2447) <= a and not b;
    outputs(2448) <= not a;
    outputs(2449) <= b;
    outputs(2450) <= a or b;
    outputs(2451) <= a xor b;
    outputs(2452) <= not (a and b);
    outputs(2453) <= b and not a;
    outputs(2454) <= not (a or b);
    outputs(2455) <= not b;
    outputs(2456) <= a xor b;
    outputs(2457) <= not a;
    outputs(2458) <= not a or b;
    outputs(2459) <= not (a and b);
    outputs(2460) <= a or b;
    outputs(2461) <= not (a and b);
    outputs(2462) <= a and b;
    outputs(2463) <= a and b;
    outputs(2464) <= a xor b;
    outputs(2465) <= not b;
    outputs(2466) <= not b;
    outputs(2467) <= not b;
    outputs(2468) <= a;
    outputs(2469) <= not (a xor b);
    outputs(2470) <= not b;
    outputs(2471) <= not a;
    outputs(2472) <= not (a or b);
    outputs(2473) <= b;
    outputs(2474) <= not b;
    outputs(2475) <= not (a or b);
    outputs(2476) <= a xor b;
    outputs(2477) <= not (a xor b);
    outputs(2478) <= not a or b;
    outputs(2479) <= a or b;
    outputs(2480) <= a or b;
    outputs(2481) <= a;
    outputs(2482) <= a;
    outputs(2483) <= not (a xor b);
    outputs(2484) <= a;
    outputs(2485) <= b and not a;
    outputs(2486) <= not (a or b);
    outputs(2487) <= not a;
    outputs(2488) <= not (a and b);
    outputs(2489) <= a xor b;
    outputs(2490) <= a xor b;
    outputs(2491) <= a;
    outputs(2492) <= a;
    outputs(2493) <= not (a and b);
    outputs(2494) <= b;
    outputs(2495) <= not (a xor b);
    outputs(2496) <= not (a xor b);
    outputs(2497) <= a xor b;
    outputs(2498) <= a or b;
    outputs(2499) <= b and not a;
    outputs(2500) <= not a;
    outputs(2501) <= a xor b;
    outputs(2502) <= not b;
    outputs(2503) <= not a;
    outputs(2504) <= not (a or b);
    outputs(2505) <= not (a or b);
    outputs(2506) <= not a;
    outputs(2507) <= not (a xor b);
    outputs(2508) <= b and not a;
    outputs(2509) <= not (a or b);
    outputs(2510) <= not (a xor b);
    outputs(2511) <= b;
    outputs(2512) <= not b or a;
    outputs(2513) <= not (a xor b);
    outputs(2514) <= not b;
    outputs(2515) <= a and not b;
    outputs(2516) <= not a;
    outputs(2517) <= a xor b;
    outputs(2518) <= not b;
    outputs(2519) <= a or b;
    outputs(2520) <= not (a xor b);
    outputs(2521) <= a and b;
    outputs(2522) <= a or b;
    outputs(2523) <= a;
    outputs(2524) <= not a or b;
    outputs(2525) <= b;
    outputs(2526) <= not a or b;
    outputs(2527) <= not a;
    outputs(2528) <= not b;
    outputs(2529) <= b and not a;
    outputs(2530) <= not b;
    outputs(2531) <= not b;
    outputs(2532) <= a;
    outputs(2533) <= not a or b;
    outputs(2534) <= not (a xor b);
    outputs(2535) <= not a or b;
    outputs(2536) <= a and not b;
    outputs(2537) <= b and not a;
    outputs(2538) <= not a;
    outputs(2539) <= b and not a;
    outputs(2540) <= not a;
    outputs(2541) <= a or b;
    outputs(2542) <= not (a and b);
    outputs(2543) <= not a;
    outputs(2544) <= a and not b;
    outputs(2545) <= not (a xor b);
    outputs(2546) <= a;
    outputs(2547) <= not (a xor b);
    outputs(2548) <= not b or a;
    outputs(2549) <= a xor b;
    outputs(2550) <= b and not a;
    outputs(2551) <= not a or b;
    outputs(2552) <= not (a xor b);
    outputs(2553) <= not (a and b);
    outputs(2554) <= not a;
    outputs(2555) <= a;
    outputs(2556) <= not (a xor b);
    outputs(2557) <= not (a xor b);
    outputs(2558) <= not (a and b);
    outputs(2559) <= not (a xor b);
    outputs(2560) <= not (a or b);
    outputs(2561) <= a xor b;
    outputs(2562) <= a and b;
    outputs(2563) <= not b;
    outputs(2564) <= not b;
    outputs(2565) <= not (a or b);
    outputs(2566) <= a;
    outputs(2567) <= not (a xor b);
    outputs(2568) <= not a;
    outputs(2569) <= not (a and b);
    outputs(2570) <= b;
    outputs(2571) <= a;
    outputs(2572) <= a and b;
    outputs(2573) <= not b;
    outputs(2574) <= not a or b;
    outputs(2575) <= a and not b;
    outputs(2576) <= not (a and b);
    outputs(2577) <= not (a xor b);
    outputs(2578) <= b and not a;
    outputs(2579) <= a;
    outputs(2580) <= not b;
    outputs(2581) <= a and not b;
    outputs(2582) <= a;
    outputs(2583) <= not (a and b);
    outputs(2584) <= a;
    outputs(2585) <= a;
    outputs(2586) <= not a;
    outputs(2587) <= not a;
    outputs(2588) <= not b;
    outputs(2589) <= not (a or b);
    outputs(2590) <= not b;
    outputs(2591) <= a xor b;
    outputs(2592) <= b;
    outputs(2593) <= not a or b;
    outputs(2594) <= a xor b;
    outputs(2595) <= not (a xor b);
    outputs(2596) <= b and not a;
    outputs(2597) <= b;
    outputs(2598) <= not a;
    outputs(2599) <= a or b;
    outputs(2600) <= b;
    outputs(2601) <= a and not b;
    outputs(2602) <= not (a xor b);
    outputs(2603) <= not a;
    outputs(2604) <= not a;
    outputs(2605) <= not (a xor b);
    outputs(2606) <= not a;
    outputs(2607) <= not b;
    outputs(2608) <= not a;
    outputs(2609) <= b;
    outputs(2610) <= a xor b;
    outputs(2611) <= not (a and b);
    outputs(2612) <= a;
    outputs(2613) <= not (a and b);
    outputs(2614) <= b;
    outputs(2615) <= a xor b;
    outputs(2616) <= a or b;
    outputs(2617) <= not (a or b);
    outputs(2618) <= not b or a;
    outputs(2619) <= a xor b;
    outputs(2620) <= not (a or b);
    outputs(2621) <= not a;
    outputs(2622) <= a xor b;
    outputs(2623) <= b and not a;
    outputs(2624) <= not b;
    outputs(2625) <= not a or b;
    outputs(2626) <= a xor b;
    outputs(2627) <= not a;
    outputs(2628) <= b;
    outputs(2629) <= not b or a;
    outputs(2630) <= not (a or b);
    outputs(2631) <= not (a xor b);
    outputs(2632) <= a xor b;
    outputs(2633) <= a xor b;
    outputs(2634) <= a or b;
    outputs(2635) <= not (a and b);
    outputs(2636) <= not b;
    outputs(2637) <= not (a and b);
    outputs(2638) <= b;
    outputs(2639) <= a;
    outputs(2640) <= not a or b;
    outputs(2641) <= not (a and b);
    outputs(2642) <= a xor b;
    outputs(2643) <= not (a and b);
    outputs(2644) <= not a or b;
    outputs(2645) <= not a or b;
    outputs(2646) <= not (a xor b);
    outputs(2647) <= a xor b;
    outputs(2648) <= not (a xor b);
    outputs(2649) <= b and not a;
    outputs(2650) <= a and not b;
    outputs(2651) <= not (a xor b);
    outputs(2652) <= not (a or b);
    outputs(2653) <= not (a and b);
    outputs(2654) <= a;
    outputs(2655) <= a xor b;
    outputs(2656) <= not a or b;
    outputs(2657) <= a and b;
    outputs(2658) <= a xor b;
    outputs(2659) <= not (a and b);
    outputs(2660) <= not b or a;
    outputs(2661) <= a xor b;
    outputs(2662) <= not a;
    outputs(2663) <= not a or b;
    outputs(2664) <= a and b;
    outputs(2665) <= b;
    outputs(2666) <= not a;
    outputs(2667) <= a;
    outputs(2668) <= a xor b;
    outputs(2669) <= b;
    outputs(2670) <= not b or a;
    outputs(2671) <= not (a or b);
    outputs(2672) <= not a;
    outputs(2673) <= not a;
    outputs(2674) <= b and not a;
    outputs(2675) <= a and not b;
    outputs(2676) <= not (a and b);
    outputs(2677) <= not (a or b);
    outputs(2678) <= not (a or b);
    outputs(2679) <= not a or b;
    outputs(2680) <= a xor b;
    outputs(2681) <= not (a or b);
    outputs(2682) <= a;
    outputs(2683) <= a;
    outputs(2684) <= a;
    outputs(2685) <= not b;
    outputs(2686) <= a and not b;
    outputs(2687) <= a;
    outputs(2688) <= a xor b;
    outputs(2689) <= not b or a;
    outputs(2690) <= not a;
    outputs(2691) <= a or b;
    outputs(2692) <= b;
    outputs(2693) <= a xor b;
    outputs(2694) <= not a or b;
    outputs(2695) <= not a or b;
    outputs(2696) <= not (a xor b);
    outputs(2697) <= not b or a;
    outputs(2698) <= b;
    outputs(2699) <= b and not a;
    outputs(2700) <= not (a or b);
    outputs(2701) <= a xor b;
    outputs(2702) <= not (a or b);
    outputs(2703) <= b;
    outputs(2704) <= not b;
    outputs(2705) <= a xor b;
    outputs(2706) <= a xor b;
    outputs(2707) <= a or b;
    outputs(2708) <= not (a xor b);
    outputs(2709) <= a and not b;
    outputs(2710) <= b;
    outputs(2711) <= not (a or b);
    outputs(2712) <= a xor b;
    outputs(2713) <= a xor b;
    outputs(2714) <= a and not b;
    outputs(2715) <= a;
    outputs(2716) <= not (a xor b);
    outputs(2717) <= not (a xor b);
    outputs(2718) <= not a;
    outputs(2719) <= a xor b;
    outputs(2720) <= not (a xor b);
    outputs(2721) <= a or b;
    outputs(2722) <= a xor b;
    outputs(2723) <= a and not b;
    outputs(2724) <= a and not b;
    outputs(2725) <= a or b;
    outputs(2726) <= a xor b;
    outputs(2727) <= a xor b;
    outputs(2728) <= not b;
    outputs(2729) <= not a;
    outputs(2730) <= b and not a;
    outputs(2731) <= not (a xor b);
    outputs(2732) <= b and not a;
    outputs(2733) <= not (a or b);
    outputs(2734) <= not b or a;
    outputs(2735) <= a;
    outputs(2736) <= a and not b;
    outputs(2737) <= not a or b;
    outputs(2738) <= a;
    outputs(2739) <= not b;
    outputs(2740) <= not a;
    outputs(2741) <= not (a xor b);
    outputs(2742) <= not a or b;
    outputs(2743) <= not (a or b);
    outputs(2744) <= not b;
    outputs(2745) <= not (a or b);
    outputs(2746) <= not a;
    outputs(2747) <= not a;
    outputs(2748) <= b;
    outputs(2749) <= not b or a;
    outputs(2750) <= a;
    outputs(2751) <= not b;
    outputs(2752) <= not a or b;
    outputs(2753) <= not a;
    outputs(2754) <= not a;
    outputs(2755) <= not (a xor b);
    outputs(2756) <= not a or b;
    outputs(2757) <= a and b;
    outputs(2758) <= not a;
    outputs(2759) <= a;
    outputs(2760) <= a xor b;
    outputs(2761) <= not (a and b);
    outputs(2762) <= not a;
    outputs(2763) <= not a or b;
    outputs(2764) <= not b;
    outputs(2765) <= a;
    outputs(2766) <= not a or b;
    outputs(2767) <= not b or a;
    outputs(2768) <= a xor b;
    outputs(2769) <= a and b;
    outputs(2770) <= a xor b;
    outputs(2771) <= a;
    outputs(2772) <= not (a and b);
    outputs(2773) <= not (a or b);
    outputs(2774) <= not a or b;
    outputs(2775) <= a xor b;
    outputs(2776) <= not (a and b);
    outputs(2777) <= not (a or b);
    outputs(2778) <= not a or b;
    outputs(2779) <= not b or a;
    outputs(2780) <= a and b;
    outputs(2781) <= not (a or b);
    outputs(2782) <= a xor b;
    outputs(2783) <= a xor b;
    outputs(2784) <= not b or a;
    outputs(2785) <= b and not a;
    outputs(2786) <= a;
    outputs(2787) <= a;
    outputs(2788) <= a xor b;
    outputs(2789) <= a or b;
    outputs(2790) <= not b;
    outputs(2791) <= b and not a;
    outputs(2792) <= b and not a;
    outputs(2793) <= b;
    outputs(2794) <= b;
    outputs(2795) <= not (a or b);
    outputs(2796) <= a xor b;
    outputs(2797) <= not b;
    outputs(2798) <= not a or b;
    outputs(2799) <= a and not b;
    outputs(2800) <= not (a or b);
    outputs(2801) <= a;
    outputs(2802) <= not a;
    outputs(2803) <= b;
    outputs(2804) <= a xor b;
    outputs(2805) <= not (a xor b);
    outputs(2806) <= not b;
    outputs(2807) <= a xor b;
    outputs(2808) <= a and b;
    outputs(2809) <= not a or b;
    outputs(2810) <= a and not b;
    outputs(2811) <= not a;
    outputs(2812) <= not (a xor b);
    outputs(2813) <= b and not a;
    outputs(2814) <= a and b;
    outputs(2815) <= a xor b;
    outputs(2816) <= not a;
    outputs(2817) <= a and not b;
    outputs(2818) <= not (a or b);
    outputs(2819) <= not b;
    outputs(2820) <= not (a and b);
    outputs(2821) <= a and not b;
    outputs(2822) <= a;
    outputs(2823) <= a or b;
    outputs(2824) <= not (a xor b);
    outputs(2825) <= not b or a;
    outputs(2826) <= a and not b;
    outputs(2827) <= not (a xor b);
    outputs(2828) <= a xor b;
    outputs(2829) <= b;
    outputs(2830) <= a;
    outputs(2831) <= not b or a;
    outputs(2832) <= not a or b;
    outputs(2833) <= a xor b;
    outputs(2834) <= not a or b;
    outputs(2835) <= not a or b;
    outputs(2836) <= a xor b;
    outputs(2837) <= not b or a;
    outputs(2838) <= b;
    outputs(2839) <= a;
    outputs(2840) <= a and not b;
    outputs(2841) <= not b or a;
    outputs(2842) <= b and not a;
    outputs(2843) <= not (a or b);
    outputs(2844) <= not a;
    outputs(2845) <= b and not a;
    outputs(2846) <= not b;
    outputs(2847) <= not a or b;
    outputs(2848) <= not (a xor b);
    outputs(2849) <= not a;
    outputs(2850) <= a and not b;
    outputs(2851) <= not a or b;
    outputs(2852) <= not a;
    outputs(2853) <= not a;
    outputs(2854) <= not (a or b);
    outputs(2855) <= a and b;
    outputs(2856) <= b;
    outputs(2857) <= not a;
    outputs(2858) <= not (a and b);
    outputs(2859) <= not (a or b);
    outputs(2860) <= a xor b;
    outputs(2861) <= not (a and b);
    outputs(2862) <= not (a or b);
    outputs(2863) <= a and not b;
    outputs(2864) <= not (a xor b);
    outputs(2865) <= not b or a;
    outputs(2866) <= not (a and b);
    outputs(2867) <= a and not b;
    outputs(2868) <= b;
    outputs(2869) <= a;
    outputs(2870) <= not (a or b);
    outputs(2871) <= not a or b;
    outputs(2872) <= not (a xor b);
    outputs(2873) <= b;
    outputs(2874) <= not (a and b);
    outputs(2875) <= b and not a;
    outputs(2876) <= b;
    outputs(2877) <= not b or a;
    outputs(2878) <= a;
    outputs(2879) <= a xor b;
    outputs(2880) <= b and not a;
    outputs(2881) <= a xor b;
    outputs(2882) <= not a or b;
    outputs(2883) <= not b or a;
    outputs(2884) <= not (a xor b);
    outputs(2885) <= b and not a;
    outputs(2886) <= not (a and b);
    outputs(2887) <= a or b;
    outputs(2888) <= not (a xor b);
    outputs(2889) <= a and not b;
    outputs(2890) <= a and not b;
    outputs(2891) <= a xor b;
    outputs(2892) <= a xor b;
    outputs(2893) <= not b;
    outputs(2894) <= b;
    outputs(2895) <= not b;
    outputs(2896) <= not (a and b);
    outputs(2897) <= not b or a;
    outputs(2898) <= not a;
    outputs(2899) <= a or b;
    outputs(2900) <= b;
    outputs(2901) <= not (a and b);
    outputs(2902) <= b and not a;
    outputs(2903) <= not b or a;
    outputs(2904) <= not (a or b);
    outputs(2905) <= not a;
    outputs(2906) <= not b;
    outputs(2907) <= not a;
    outputs(2908) <= not a;
    outputs(2909) <= b and not a;
    outputs(2910) <= a xor b;
    outputs(2911) <= a and b;
    outputs(2912) <= not (a xor b);
    outputs(2913) <= not b;
    outputs(2914) <= a xor b;
    outputs(2915) <= not a or b;
    outputs(2916) <= not b;
    outputs(2917) <= a;
    outputs(2918) <= b and not a;
    outputs(2919) <= not (a and b);
    outputs(2920) <= not (a xor b);
    outputs(2921) <= b and not a;
    outputs(2922) <= b and not a;
    outputs(2923) <= b;
    outputs(2924) <= a xor b;
    outputs(2925) <= a and b;
    outputs(2926) <= a and not b;
    outputs(2927) <= a;
    outputs(2928) <= not a;
    outputs(2929) <= not b;
    outputs(2930) <= a or b;
    outputs(2931) <= not (a xor b);
    outputs(2932) <= not a or b;
    outputs(2933) <= a xor b;
    outputs(2934) <= a xor b;
    outputs(2935) <= not b;
    outputs(2936) <= b and not a;
    outputs(2937) <= not a;
    outputs(2938) <= not a or b;
    outputs(2939) <= not b;
    outputs(2940) <= not (a xor b);
    outputs(2941) <= a and b;
    outputs(2942) <= b;
    outputs(2943) <= not (a xor b);
    outputs(2944) <= not b or a;
    outputs(2945) <= not b;
    outputs(2946) <= not (a or b);
    outputs(2947) <= a and not b;
    outputs(2948) <= a;
    outputs(2949) <= a;
    outputs(2950) <= a and b;
    outputs(2951) <= a or b;
    outputs(2952) <= not b or a;
    outputs(2953) <= a or b;
    outputs(2954) <= a and b;
    outputs(2955) <= a and not b;
    outputs(2956) <= not b or a;
    outputs(2957) <= not a or b;
    outputs(2958) <= not (a xor b);
    outputs(2959) <= not (a xor b);
    outputs(2960) <= not b;
    outputs(2961) <= a and not b;
    outputs(2962) <= b and not a;
    outputs(2963) <= not (a xor b);
    outputs(2964) <= not (a xor b);
    outputs(2965) <= not a;
    outputs(2966) <= not b;
    outputs(2967) <= b;
    outputs(2968) <= not (a xor b);
    outputs(2969) <= a or b;
    outputs(2970) <= a xor b;
    outputs(2971) <= a;
    outputs(2972) <= a;
    outputs(2973) <= a;
    outputs(2974) <= not a;
    outputs(2975) <= a and not b;
    outputs(2976) <= not a or b;
    outputs(2977) <= a or b;
    outputs(2978) <= a xor b;
    outputs(2979) <= not b;
    outputs(2980) <= b;
    outputs(2981) <= b;
    outputs(2982) <= not (a xor b);
    outputs(2983) <= a or b;
    outputs(2984) <= not a;
    outputs(2985) <= a or b;
    outputs(2986) <= a xor b;
    outputs(2987) <= a xor b;
    outputs(2988) <= b and not a;
    outputs(2989) <= not (a and b);
    outputs(2990) <= b;
    outputs(2991) <= a;
    outputs(2992) <= not b;
    outputs(2993) <= a xor b;
    outputs(2994) <= b;
    outputs(2995) <= not (a or b);
    outputs(2996) <= a xor b;
    outputs(2997) <= b;
    outputs(2998) <= a or b;
    outputs(2999) <= not b;
    outputs(3000) <= a or b;
    outputs(3001) <= not b;
    outputs(3002) <= not (a xor b);
    outputs(3003) <= a xor b;
    outputs(3004) <= not a;
    outputs(3005) <= not (a xor b);
    outputs(3006) <= not (a xor b);
    outputs(3007) <= b and not a;
    outputs(3008) <= not a;
    outputs(3009) <= a xor b;
    outputs(3010) <= a;
    outputs(3011) <= not a;
    outputs(3012) <= not b;
    outputs(3013) <= b and not a;
    outputs(3014) <= not (a and b);
    outputs(3015) <= a or b;
    outputs(3016) <= a or b;
    outputs(3017) <= not (a xor b);
    outputs(3018) <= a;
    outputs(3019) <= not (a and b);
    outputs(3020) <= not a;
    outputs(3021) <= not (a or b);
    outputs(3022) <= a xor b;
    outputs(3023) <= not a;
    outputs(3024) <= a xor b;
    outputs(3025) <= not (a and b);
    outputs(3026) <= a and not b;
    outputs(3027) <= not a or b;
    outputs(3028) <= b and not a;
    outputs(3029) <= not a;
    outputs(3030) <= not b or a;
    outputs(3031) <= a and not b;
    outputs(3032) <= a and b;
    outputs(3033) <= a or b;
    outputs(3034) <= a or b;
    outputs(3035) <= a and not b;
    outputs(3036) <= a;
    outputs(3037) <= a xor b;
    outputs(3038) <= a xor b;
    outputs(3039) <= a;
    outputs(3040) <= b;
    outputs(3041) <= a;
    outputs(3042) <= a or b;
    outputs(3043) <= not a;
    outputs(3044) <= not (a xor b);
    outputs(3045) <= not (a xor b);
    outputs(3046) <= a and not b;
    outputs(3047) <= not b;
    outputs(3048) <= b and not a;
    outputs(3049) <= not (a xor b);
    outputs(3050) <= a or b;
    outputs(3051) <= a;
    outputs(3052) <= a;
    outputs(3053) <= a;
    outputs(3054) <= not b;
    outputs(3055) <= not a;
    outputs(3056) <= not (a xor b);
    outputs(3057) <= not a or b;
    outputs(3058) <= not a;
    outputs(3059) <= not (a or b);
    outputs(3060) <= a;
    outputs(3061) <= not a or b;
    outputs(3062) <= not (a and b);
    outputs(3063) <= not b;
    outputs(3064) <= not a;
    outputs(3065) <= not b;
    outputs(3066) <= not a;
    outputs(3067) <= not (a xor b);
    outputs(3068) <= not b;
    outputs(3069) <= b;
    outputs(3070) <= not (a xor b);
    outputs(3071) <= a xor b;
    outputs(3072) <= a and b;
    outputs(3073) <= not (a or b);
    outputs(3074) <= a and not b;
    outputs(3075) <= b;
    outputs(3076) <= b;
    outputs(3077) <= a;
    outputs(3078) <= not (a or b);
    outputs(3079) <= not (a or b);
    outputs(3080) <= a;
    outputs(3081) <= a xor b;
    outputs(3082) <= not (a and b);
    outputs(3083) <= not b;
    outputs(3084) <= b and not a;
    outputs(3085) <= a xor b;
    outputs(3086) <= not b;
    outputs(3087) <= not a;
    outputs(3088) <= b and not a;
    outputs(3089) <= not b;
    outputs(3090) <= not (a xor b);
    outputs(3091) <= not (a xor b);
    outputs(3092) <= not (a or b);
    outputs(3093) <= a;
    outputs(3094) <= a;
    outputs(3095) <= b and not a;
    outputs(3096) <= 1'b0;
    outputs(3097) <= not (a xor b);
    outputs(3098) <= b and not a;
    outputs(3099) <= b;
    outputs(3100) <= b;
    outputs(3101) <= a;
    outputs(3102) <= a;
    outputs(3103) <= b and not a;
    outputs(3104) <= not (a xor b);
    outputs(3105) <= b;
    outputs(3106) <= b and not a;
    outputs(3107) <= not (a and b);
    outputs(3108) <= a;
    outputs(3109) <= a xor b;
    outputs(3110) <= a and b;
    outputs(3111) <= not (a or b);
    outputs(3112) <= a and b;
    outputs(3113) <= not (a xor b);
    outputs(3114) <= not a;
    outputs(3115) <= a or b;
    outputs(3116) <= a xor b;
    outputs(3117) <= not a;
    outputs(3118) <= b and not a;
    outputs(3119) <= a or b;
    outputs(3120) <= not (a xor b);
    outputs(3121) <= a and not b;
    outputs(3122) <= not (a and b);
    outputs(3123) <= not b;
    outputs(3124) <= not (a or b);
    outputs(3125) <= not (a xor b);
    outputs(3126) <= b and not a;
    outputs(3127) <= a and b;
    outputs(3128) <= not a;
    outputs(3129) <= not (a or b);
    outputs(3130) <= b and not a;
    outputs(3131) <= not (a xor b);
    outputs(3132) <= not a or b;
    outputs(3133) <= not (a xor b);
    outputs(3134) <= a xor b;
    outputs(3135) <= not b or a;
    outputs(3136) <= not b;
    outputs(3137) <= not (a xor b);
    outputs(3138) <= a and b;
    outputs(3139) <= a xor b;
    outputs(3140) <= b;
    outputs(3141) <= not b or a;
    outputs(3142) <= a xor b;
    outputs(3143) <= not (a xor b);
    outputs(3144) <= not a;
    outputs(3145) <= not a;
    outputs(3146) <= b;
    outputs(3147) <= not a;
    outputs(3148) <= not (a xor b);
    outputs(3149) <= b and not a;
    outputs(3150) <= a xor b;
    outputs(3151) <= a and b;
    outputs(3152) <= a;
    outputs(3153) <= a xor b;
    outputs(3154) <= not a;
    outputs(3155) <= not b;
    outputs(3156) <= a and not b;
    outputs(3157) <= a xor b;
    outputs(3158) <= not (a or b);
    outputs(3159) <= a and not b;
    outputs(3160) <= not (a xor b);
    outputs(3161) <= not a;
    outputs(3162) <= not a;
    outputs(3163) <= b and not a;
    outputs(3164) <= not a;
    outputs(3165) <= a xor b;
    outputs(3166) <= not (a xor b);
    outputs(3167) <= not (a xor b);
    outputs(3168) <= not (a and b);
    outputs(3169) <= not (a or b);
    outputs(3170) <= a;
    outputs(3171) <= a and b;
    outputs(3172) <= a and not b;
    outputs(3173) <= a and b;
    outputs(3174) <= a xor b;
    outputs(3175) <= not b;
    outputs(3176) <= a and not b;
    outputs(3177) <= a;
    outputs(3178) <= not b;
    outputs(3179) <= not (a or b);
    outputs(3180) <= a and not b;
    outputs(3181) <= a;
    outputs(3182) <= a and not b;
    outputs(3183) <= a;
    outputs(3184) <= a and not b;
    outputs(3185) <= not (a and b);
    outputs(3186) <= a xor b;
    outputs(3187) <= a;
    outputs(3188) <= a;
    outputs(3189) <= not (a xor b);
    outputs(3190) <= not a;
    outputs(3191) <= not b;
    outputs(3192) <= not a;
    outputs(3193) <= not (a xor b);
    outputs(3194) <= a or b;
    outputs(3195) <= a and not b;
    outputs(3196) <= a and not b;
    outputs(3197) <= a;
    outputs(3198) <= b;
    outputs(3199) <= not (a xor b);
    outputs(3200) <= not b;
    outputs(3201) <= not b;
    outputs(3202) <= b and not a;
    outputs(3203) <= not (a xor b);
    outputs(3204) <= not (a or b);
    outputs(3205) <= a and not b;
    outputs(3206) <= a and b;
    outputs(3207) <= not b or a;
    outputs(3208) <= 1'b0;
    outputs(3209) <= a and not b;
    outputs(3210) <= b and not a;
    outputs(3211) <= a xor b;
    outputs(3212) <= not (a xor b);
    outputs(3213) <= a;
    outputs(3214) <= b;
    outputs(3215) <= a;
    outputs(3216) <= b and not a;
    outputs(3217) <= b and not a;
    outputs(3218) <= a and b;
    outputs(3219) <= b;
    outputs(3220) <= b;
    outputs(3221) <= b;
    outputs(3222) <= a or b;
    outputs(3223) <= not b;
    outputs(3224) <= not a;
    outputs(3225) <= a and b;
    outputs(3226) <= b and not a;
    outputs(3227) <= not (a or b);
    outputs(3228) <= not (a xor b);
    outputs(3229) <= not (a or b);
    outputs(3230) <= a;
    outputs(3231) <= not (a or b);
    outputs(3232) <= not (a xor b);
    outputs(3233) <= not b;
    outputs(3234) <= not b;
    outputs(3235) <= not a;
    outputs(3236) <= not a;
    outputs(3237) <= a;
    outputs(3238) <= b;
    outputs(3239) <= not b or a;
    outputs(3240) <= not (a or b);
    outputs(3241) <= a xor b;
    outputs(3242) <= not (a xor b);
    outputs(3243) <= a and not b;
    outputs(3244) <= a xor b;
    outputs(3245) <= a and b;
    outputs(3246) <= a and b;
    outputs(3247) <= not a;
    outputs(3248) <= not (a xor b);
    outputs(3249) <= a and not b;
    outputs(3250) <= a and not b;
    outputs(3251) <= not b or a;
    outputs(3252) <= not b;
    outputs(3253) <= not (a or b);
    outputs(3254) <= not (a or b);
    outputs(3255) <= a xor b;
    outputs(3256) <= a;
    outputs(3257) <= not (a or b);
    outputs(3258) <= b and not a;
    outputs(3259) <= a and not b;
    outputs(3260) <= b and not a;
    outputs(3261) <= a and not b;
    outputs(3262) <= b and not a;
    outputs(3263) <= b and not a;
    outputs(3264) <= a xor b;
    outputs(3265) <= a or b;
    outputs(3266) <= a and b;
    outputs(3267) <= not (a xor b);
    outputs(3268) <= a xor b;
    outputs(3269) <= not (a or b);
    outputs(3270) <= 1'b0;
    outputs(3271) <= not (a xor b);
    outputs(3272) <= a and b;
    outputs(3273) <= a and b;
    outputs(3274) <= a xor b;
    outputs(3275) <= b;
    outputs(3276) <= not (a xor b);
    outputs(3277) <= b and not a;
    outputs(3278) <= b and not a;
    outputs(3279) <= b;
    outputs(3280) <= a and b;
    outputs(3281) <= b and not a;
    outputs(3282) <= not (a or b);
    outputs(3283) <= b and not a;
    outputs(3284) <= not (a or b);
    outputs(3285) <= b;
    outputs(3286) <= not (a or b);
    outputs(3287) <= b;
    outputs(3288) <= a;
    outputs(3289) <= a xor b;
    outputs(3290) <= not a;
    outputs(3291) <= a and b;
    outputs(3292) <= not (a xor b);
    outputs(3293) <= a and b;
    outputs(3294) <= a and b;
    outputs(3295) <= a xor b;
    outputs(3296) <= a;
    outputs(3297) <= b;
    outputs(3298) <= not (a or b);
    outputs(3299) <= a;
    outputs(3300) <= b and not a;
    outputs(3301) <= a xor b;
    outputs(3302) <= not b or a;
    outputs(3303) <= not (a or b);
    outputs(3304) <= not a;
    outputs(3305) <= not (a or b);
    outputs(3306) <= a;
    outputs(3307) <= not (a or b);
    outputs(3308) <= not (a xor b);
    outputs(3309) <= a and not b;
    outputs(3310) <= not (a or b);
    outputs(3311) <= a;
    outputs(3312) <= 1'b0;
    outputs(3313) <= not b;
    outputs(3314) <= b;
    outputs(3315) <= a and b;
    outputs(3316) <= a;
    outputs(3317) <= a and not b;
    outputs(3318) <= not (a or b);
    outputs(3319) <= not b;
    outputs(3320) <= a and b;
    outputs(3321) <= not a;
    outputs(3322) <= not b;
    outputs(3323) <= not (a xor b);
    outputs(3324) <= a and b;
    outputs(3325) <= not a;
    outputs(3326) <= not (a or b);
    outputs(3327) <= a and b;
    outputs(3328) <= not (a xor b);
    outputs(3329) <= a xor b;
    outputs(3330) <= not (a or b);
    outputs(3331) <= not (a or b);
    outputs(3332) <= a;
    outputs(3333) <= not (a or b);
    outputs(3334) <= not (a or b);
    outputs(3335) <= not a;
    outputs(3336) <= a and b;
    outputs(3337) <= a and not b;
    outputs(3338) <= not (a or b);
    outputs(3339) <= not a;
    outputs(3340) <= a and not b;
    outputs(3341) <= not (a xor b);
    outputs(3342) <= not (a xor b);
    outputs(3343) <= not b or a;
    outputs(3344) <= not b;
    outputs(3345) <= not b;
    outputs(3346) <= not (a xor b);
    outputs(3347) <= not a;
    outputs(3348) <= b;
    outputs(3349) <= a;
    outputs(3350) <= not (a or b);
    outputs(3351) <= a;
    outputs(3352) <= not (a xor b);
    outputs(3353) <= a and b;
    outputs(3354) <= a and not b;
    outputs(3355) <= not a or b;
    outputs(3356) <= a and not b;
    outputs(3357) <= a;
    outputs(3358) <= not b;
    outputs(3359) <= a;
    outputs(3360) <= not (a xor b);
    outputs(3361) <= a or b;
    outputs(3362) <= not (a xor b);
    outputs(3363) <= a and b;
    outputs(3364) <= not b;
    outputs(3365) <= a and not b;
    outputs(3366) <= b;
    outputs(3367) <= b and not a;
    outputs(3368) <= a and b;
    outputs(3369) <= a or b;
    outputs(3370) <= b and not a;
    outputs(3371) <= not b;
    outputs(3372) <= a xor b;
    outputs(3373) <= a;
    outputs(3374) <= not (a xor b);
    outputs(3375) <= not b;
    outputs(3376) <= not (a or b);
    outputs(3377) <= a and b;
    outputs(3378) <= not a;
    outputs(3379) <= not (a xor b);
    outputs(3380) <= a xor b;
    outputs(3381) <= a and not b;
    outputs(3382) <= b and not a;
    outputs(3383) <= not b;
    outputs(3384) <= not (a and b);
    outputs(3385) <= not b;
    outputs(3386) <= b;
    outputs(3387) <= b and not a;
    outputs(3388) <= a;
    outputs(3389) <= a and b;
    outputs(3390) <= not b;
    outputs(3391) <= not b;
    outputs(3392) <= not a;
    outputs(3393) <= not (a or b);
    outputs(3394) <= a and b;
    outputs(3395) <= not (a and b);
    outputs(3396) <= not (a and b);
    outputs(3397) <= a and b;
    outputs(3398) <= not b;
    outputs(3399) <= a xor b;
    outputs(3400) <= b and not a;
    outputs(3401) <= not (a xor b);
    outputs(3402) <= not b or a;
    outputs(3403) <= not (a or b);
    outputs(3404) <= b;
    outputs(3405) <= b;
    outputs(3406) <= not a;
    outputs(3407) <= not (a or b);
    outputs(3408) <= a and b;
    outputs(3409) <= a and b;
    outputs(3410) <= not (a or b);
    outputs(3411) <= a;
    outputs(3412) <= a;
    outputs(3413) <= a and b;
    outputs(3414) <= b;
    outputs(3415) <= a xor b;
    outputs(3416) <= not (a xor b);
    outputs(3417) <= b;
    outputs(3418) <= not (a or b);
    outputs(3419) <= not b;
    outputs(3420) <= not (a or b);
    outputs(3421) <= b;
    outputs(3422) <= a and b;
    outputs(3423) <= not (a xor b);
    outputs(3424) <= a xor b;
    outputs(3425) <= a;
    outputs(3426) <= a and not b;
    outputs(3427) <= not b;
    outputs(3428) <= not (a xor b);
    outputs(3429) <= not (a or b);
    outputs(3430) <= not (a xor b);
    outputs(3431) <= not (a xor b);
    outputs(3432) <= b and not a;
    outputs(3433) <= a and not b;
    outputs(3434) <= b and not a;
    outputs(3435) <= a xor b;
    outputs(3436) <= a or b;
    outputs(3437) <= a;
    outputs(3438) <= not b;
    outputs(3439) <= not a;
    outputs(3440) <= b;
    outputs(3441) <= a xor b;
    outputs(3442) <= b and not a;
    outputs(3443) <= b;
    outputs(3444) <= b;
    outputs(3445) <= a and not b;
    outputs(3446) <= a and b;
    outputs(3447) <= b and not a;
    outputs(3448) <= not (a xor b);
    outputs(3449) <= not (a or b);
    outputs(3450) <= a;
    outputs(3451) <= not (a or b);
    outputs(3452) <= a and b;
    outputs(3453) <= not (a xor b);
    outputs(3454) <= b;
    outputs(3455) <= a xor b;
    outputs(3456) <= not a or b;
    outputs(3457) <= not b or a;
    outputs(3458) <= a xor b;
    outputs(3459) <= a and not b;
    outputs(3460) <= b and not a;
    outputs(3461) <= not a;
    outputs(3462) <= b;
    outputs(3463) <= b and not a;
    outputs(3464) <= not (a or b);
    outputs(3465) <= b;
    outputs(3466) <= not (a and b);
    outputs(3467) <= a xor b;
    outputs(3468) <= b and not a;
    outputs(3469) <= a xor b;
    outputs(3470) <= a xor b;
    outputs(3471) <= a;
    outputs(3472) <= a and not b;
    outputs(3473) <= not (a or b);
    outputs(3474) <= not b;
    outputs(3475) <= not a;
    outputs(3476) <= not (a xor b);
    outputs(3477) <= not a;
    outputs(3478) <= not (a or b);
    outputs(3479) <= not (a xor b);
    outputs(3480) <= not b;
    outputs(3481) <= b and not a;
    outputs(3482) <= a and not b;
    outputs(3483) <= not b;
    outputs(3484) <= b;
    outputs(3485) <= a and not b;
    outputs(3486) <= not (a or b);
    outputs(3487) <= b and not a;
    outputs(3488) <= not b;
    outputs(3489) <= not (a or b);
    outputs(3490) <= not b;
    outputs(3491) <= not a;
    outputs(3492) <= not b;
    outputs(3493) <= not (a or b);
    outputs(3494) <= a;
    outputs(3495) <= not (a xor b);
    outputs(3496) <= b;
    outputs(3497) <= not a;
    outputs(3498) <= not (a or b);
    outputs(3499) <= not (a or b);
    outputs(3500) <= a;
    outputs(3501) <= a;
    outputs(3502) <= a and not b;
    outputs(3503) <= not b;
    outputs(3504) <= not (a and b);
    outputs(3505) <= not b;
    outputs(3506) <= b and not a;
    outputs(3507) <= b and not a;
    outputs(3508) <= a and b;
    outputs(3509) <= not (a or b);
    outputs(3510) <= not (a xor b);
    outputs(3511) <= not (a xor b);
    outputs(3512) <= b;
    outputs(3513) <= a and b;
    outputs(3514) <= a;
    outputs(3515) <= not (a or b);
    outputs(3516) <= b and not a;
    outputs(3517) <= not a;
    outputs(3518) <= not b or a;
    outputs(3519) <= a and b;
    outputs(3520) <= b;
    outputs(3521) <= not b;
    outputs(3522) <= not (a xor b);
    outputs(3523) <= not (a and b);
    outputs(3524) <= a;
    outputs(3525) <= a and not b;
    outputs(3526) <= b and not a;
    outputs(3527) <= not a;
    outputs(3528) <= a;
    outputs(3529) <= a;
    outputs(3530) <= b and not a;
    outputs(3531) <= b and not a;
    outputs(3532) <= not (a or b);
    outputs(3533) <= a xor b;
    outputs(3534) <= not (a xor b);
    outputs(3535) <= a and not b;
    outputs(3536) <= a xor b;
    outputs(3537) <= not b;
    outputs(3538) <= not (a or b);
    outputs(3539) <= a and not b;
    outputs(3540) <= not (a or b);
    outputs(3541) <= not a;
    outputs(3542) <= a xor b;
    outputs(3543) <= b and not a;
    outputs(3544) <= not (a or b);
    outputs(3545) <= not b;
    outputs(3546) <= not (a or b);
    outputs(3547) <= not (a xor b);
    outputs(3548) <= a xor b;
    outputs(3549) <= not b or a;
    outputs(3550) <= a and b;
    outputs(3551) <= not a;
    outputs(3552) <= a;
    outputs(3553) <= b and not a;
    outputs(3554) <= a;
    outputs(3555) <= not (a or b);
    outputs(3556) <= b and not a;
    outputs(3557) <= b;
    outputs(3558) <= a and not b;
    outputs(3559) <= a;
    outputs(3560) <= b and not a;
    outputs(3561) <= a and not b;
    outputs(3562) <= a xor b;
    outputs(3563) <= not (a or b);
    outputs(3564) <= not a;
    outputs(3565) <= a;
    outputs(3566) <= not (a or b);
    outputs(3567) <= not (a xor b);
    outputs(3568) <= b and not a;
    outputs(3569) <= a;
    outputs(3570) <= not (a xor b);
    outputs(3571) <= not (a or b);
    outputs(3572) <= b;
    outputs(3573) <= a;
    outputs(3574) <= a xor b;
    outputs(3575) <= b and not a;
    outputs(3576) <= not (a xor b);
    outputs(3577) <= a and b;
    outputs(3578) <= b;
    outputs(3579) <= a and not b;
    outputs(3580) <= not b or a;
    outputs(3581) <= b;
    outputs(3582) <= a and b;
    outputs(3583) <= not (a and b);
    outputs(3584) <= not (a xor b);
    outputs(3585) <= a and b;
    outputs(3586) <= not b;
    outputs(3587) <= b;
    outputs(3588) <= a;
    outputs(3589) <= a xor b;
    outputs(3590) <= a xor b;
    outputs(3591) <= a xor b;
    outputs(3592) <= not b;
    outputs(3593) <= a and not b;
    outputs(3594) <= not a;
    outputs(3595) <= not a;
    outputs(3596) <= a and b;
    outputs(3597) <= a or b;
    outputs(3598) <= not (a xor b);
    outputs(3599) <= not a;
    outputs(3600) <= not b;
    outputs(3601) <= a or b;
    outputs(3602) <= a;
    outputs(3603) <= not (a and b);
    outputs(3604) <= not a;
    outputs(3605) <= not (a xor b);
    outputs(3606) <= not b;
    outputs(3607) <= not b;
    outputs(3608) <= not b;
    outputs(3609) <= not a;
    outputs(3610) <= not a;
    outputs(3611) <= a and b;
    outputs(3612) <= not a;
    outputs(3613) <= not (a or b);
    outputs(3614) <= not (a or b);
    outputs(3615) <= not a;
    outputs(3616) <= a or b;
    outputs(3617) <= a and b;
    outputs(3618) <= not a;
    outputs(3619) <= not a;
    outputs(3620) <= not (a xor b);
    outputs(3621) <= not a;
    outputs(3622) <= not a;
    outputs(3623) <= not (a and b);
    outputs(3624) <= a and b;
    outputs(3625) <= not b;
    outputs(3626) <= b and not a;
    outputs(3627) <= b;
    outputs(3628) <= b;
    outputs(3629) <= a;
    outputs(3630) <= not a;
    outputs(3631) <= not b or a;
    outputs(3632) <= a and not b;
    outputs(3633) <= not b;
    outputs(3634) <= b and not a;
    outputs(3635) <= a and not b;
    outputs(3636) <= a;
    outputs(3637) <= not (a or b);
    outputs(3638) <= a and b;
    outputs(3639) <= a or b;
    outputs(3640) <= not (a and b);
    outputs(3641) <= not b;
    outputs(3642) <= not (a xor b);
    outputs(3643) <= a xor b;
    outputs(3644) <= a;
    outputs(3645) <= not b;
    outputs(3646) <= a and b;
    outputs(3647) <= not (a xor b);
    outputs(3648) <= b and not a;
    outputs(3649) <= a xor b;
    outputs(3650) <= not b;
    outputs(3651) <= a and b;
    outputs(3652) <= a;
    outputs(3653) <= not (a or b);
    outputs(3654) <= not (a or b);
    outputs(3655) <= not (a or b);
    outputs(3656) <= not b;
    outputs(3657) <= a xor b;
    outputs(3658) <= not (a or b);
    outputs(3659) <= b and not a;
    outputs(3660) <= b and not a;
    outputs(3661) <= a xor b;
    outputs(3662) <= not (a or b);
    outputs(3663) <= a;
    outputs(3664) <= a and b;
    outputs(3665) <= not a;
    outputs(3666) <= not b;
    outputs(3667) <= b and not a;
    outputs(3668) <= not (a xor b);
    outputs(3669) <= not a;
    outputs(3670) <= not (a xor b);
    outputs(3671) <= not b;
    outputs(3672) <= a and b;
    outputs(3673) <= not b;
    outputs(3674) <= not (a xor b);
    outputs(3675) <= not a;
    outputs(3676) <= b and not a;
    outputs(3677) <= not b;
    outputs(3678) <= a or b;
    outputs(3679) <= not a;
    outputs(3680) <= a and not b;
    outputs(3681) <= not (a or b);
    outputs(3682) <= not b or a;
    outputs(3683) <= not b;
    outputs(3684) <= a and b;
    outputs(3685) <= a;
    outputs(3686) <= not a;
    outputs(3687) <= a xor b;
    outputs(3688) <= not (a xor b);
    outputs(3689) <= a and b;
    outputs(3690) <= a xor b;
    outputs(3691) <= a and b;
    outputs(3692) <= not (a xor b);
    outputs(3693) <= a and not b;
    outputs(3694) <= not (a xor b);
    outputs(3695) <= not a;
    outputs(3696) <= not (a or b);
    outputs(3697) <= a xor b;
    outputs(3698) <= not b;
    outputs(3699) <= not (a or b);
    outputs(3700) <= a;
    outputs(3701) <= a;
    outputs(3702) <= a and b;
    outputs(3703) <= a and not b;
    outputs(3704) <= b and not a;
    outputs(3705) <= not (a xor b);
    outputs(3706) <= not (a xor b);
    outputs(3707) <= b and not a;
    outputs(3708) <= not (a or b);
    outputs(3709) <= a xor b;
    outputs(3710) <= a and not b;
    outputs(3711) <= not (a xor b);
    outputs(3712) <= not (a or b);
    outputs(3713) <= not a;
    outputs(3714) <= not (a xor b);
    outputs(3715) <= a and b;
    outputs(3716) <= a xor b;
    outputs(3717) <= not (a or b);
    outputs(3718) <= not a;
    outputs(3719) <= not a;
    outputs(3720) <= a xor b;
    outputs(3721) <= a xor b;
    outputs(3722) <= b and not a;
    outputs(3723) <= a and not b;
    outputs(3724) <= a;
    outputs(3725) <= a;
    outputs(3726) <= not a;
    outputs(3727) <= not a;
    outputs(3728) <= a xor b;
    outputs(3729) <= a xor b;
    outputs(3730) <= a and b;
    outputs(3731) <= not (a or b);
    outputs(3732) <= not (a xor b);
    outputs(3733) <= b;
    outputs(3734) <= not (a or b);
    outputs(3735) <= b and not a;
    outputs(3736) <= b;
    outputs(3737) <= not b;
    outputs(3738) <= not (a or b);
    outputs(3739) <= a and not b;
    outputs(3740) <= b;
    outputs(3741) <= not (a xor b);
    outputs(3742) <= b;
    outputs(3743) <= b and not a;
    outputs(3744) <= b;
    outputs(3745) <= not a;
    outputs(3746) <= a;
    outputs(3747) <= not (a xor b);
    outputs(3748) <= not (a or b);
    outputs(3749) <= a xor b;
    outputs(3750) <= not (a or b);
    outputs(3751) <= a and b;
    outputs(3752) <= not a;
    outputs(3753) <= not a;
    outputs(3754) <= a;
    outputs(3755) <= b and not a;
    outputs(3756) <= not b;
    outputs(3757) <= a and not b;
    outputs(3758) <= a and b;
    outputs(3759) <= not (a and b);
    outputs(3760) <= a and not b;
    outputs(3761) <= a and not b;
    outputs(3762) <= not (a xor b);
    outputs(3763) <= not b or a;
    outputs(3764) <= a;
    outputs(3765) <= a and b;
    outputs(3766) <= a;
    outputs(3767) <= b and not a;
    outputs(3768) <= a;
    outputs(3769) <= a and b;
    outputs(3770) <= not b;
    outputs(3771) <= not b;
    outputs(3772) <= b;
    outputs(3773) <= a xor b;
    outputs(3774) <= a xor b;
    outputs(3775) <= not (a or b);
    outputs(3776) <= not b;
    outputs(3777) <= b and not a;
    outputs(3778) <= not a;
    outputs(3779) <= not a or b;
    outputs(3780) <= a xor b;
    outputs(3781) <= not a;
    outputs(3782) <= a and not b;
    outputs(3783) <= a;
    outputs(3784) <= b;
    outputs(3785) <= a and b;
    outputs(3786) <= a;
    outputs(3787) <= not (a xor b);
    outputs(3788) <= not a;
    outputs(3789) <= a;
    outputs(3790) <= a xor b;
    outputs(3791) <= a;
    outputs(3792) <= not (a or b);
    outputs(3793) <= not (a xor b);
    outputs(3794) <= not (a or b);
    outputs(3795) <= not b;
    outputs(3796) <= b;
    outputs(3797) <= b and not a;
    outputs(3798) <= not (a or b);
    outputs(3799) <= a and not b;
    outputs(3800) <= b;
    outputs(3801) <= a and b;
    outputs(3802) <= a and not b;
    outputs(3803) <= not (a xor b);
    outputs(3804) <= not (a or b);
    outputs(3805) <= a and not b;
    outputs(3806) <= a;
    outputs(3807) <= a or b;
    outputs(3808) <= b;
    outputs(3809) <= a xor b;
    outputs(3810) <= not (a or b);
    outputs(3811) <= not a;
    outputs(3812) <= not (a and b);
    outputs(3813) <= not a;
    outputs(3814) <= not b;
    outputs(3815) <= a and not b;
    outputs(3816) <= not b or a;
    outputs(3817) <= a;
    outputs(3818) <= not a or b;
    outputs(3819) <= not a;
    outputs(3820) <= not (a xor b);
    outputs(3821) <= a xor b;
    outputs(3822) <= a and b;
    outputs(3823) <= a;
    outputs(3824) <= not a;
    outputs(3825) <= not (a or b);
    outputs(3826) <= not b;
    outputs(3827) <= b;
    outputs(3828) <= a and b;
    outputs(3829) <= not a;
    outputs(3830) <= not a or b;
    outputs(3831) <= a xor b;
    outputs(3832) <= b;
    outputs(3833) <= not (a or b);
    outputs(3834) <= a;
    outputs(3835) <= not (a or b);
    outputs(3836) <= a;
    outputs(3837) <= not b or a;
    outputs(3838) <= a and not b;
    outputs(3839) <= b;
    outputs(3840) <= b and not a;
    outputs(3841) <= b;
    outputs(3842) <= not a or b;
    outputs(3843) <= a xor b;
    outputs(3844) <= b and not a;
    outputs(3845) <= a xor b;
    outputs(3846) <= a;
    outputs(3847) <= not (a and b);
    outputs(3848) <= a xor b;
    outputs(3849) <= a and not b;
    outputs(3850) <= not b;
    outputs(3851) <= a and not b;
    outputs(3852) <= b and not a;
    outputs(3853) <= a and b;
    outputs(3854) <= a or b;
    outputs(3855) <= not b;
    outputs(3856) <= a;
    outputs(3857) <= not (a xor b);
    outputs(3858) <= b and not a;
    outputs(3859) <= not b;
    outputs(3860) <= b;
    outputs(3861) <= not (a or b);
    outputs(3862) <= not a;
    outputs(3863) <= not b or a;
    outputs(3864) <= not b;
    outputs(3865) <= not b;
    outputs(3866) <= not a;
    outputs(3867) <= not b;
    outputs(3868) <= not a;
    outputs(3869) <= not (a xor b);
    outputs(3870) <= not (a xor b);
    outputs(3871) <= not (a xor b);
    outputs(3872) <= a xor b;
    outputs(3873) <= not a;
    outputs(3874) <= a and b;
    outputs(3875) <= not (a and b);
    outputs(3876) <= not a;
    outputs(3877) <= a xor b;
    outputs(3878) <= not a or b;
    outputs(3879) <= not (a or b);
    outputs(3880) <= not (a xor b);
    outputs(3881) <= a xor b;
    outputs(3882) <= not a;
    outputs(3883) <= a;
    outputs(3884) <= a or b;
    outputs(3885) <= a xor b;
    outputs(3886) <= a;
    outputs(3887) <= not a or b;
    outputs(3888) <= not (a xor b);
    outputs(3889) <= not a;
    outputs(3890) <= a xor b;
    outputs(3891) <= a xor b;
    outputs(3892) <= not a;
    outputs(3893) <= a or b;
    outputs(3894) <= a xor b;
    outputs(3895) <= a or b;
    outputs(3896) <= not a;
    outputs(3897) <= not b;
    outputs(3898) <= not b;
    outputs(3899) <= b;
    outputs(3900) <= a xor b;
    outputs(3901) <= not (a xor b);
    outputs(3902) <= a xor b;
    outputs(3903) <= a xor b;
    outputs(3904) <= b;
    outputs(3905) <= not a;
    outputs(3906) <= b;
    outputs(3907) <= b;
    outputs(3908) <= not b;
    outputs(3909) <= b and not a;
    outputs(3910) <= a;
    outputs(3911) <= a xor b;
    outputs(3912) <= not a;
    outputs(3913) <= not b;
    outputs(3914) <= a and b;
    outputs(3915) <= not b or a;
    outputs(3916) <= not (a xor b);
    outputs(3917) <= not b or a;
    outputs(3918) <= not a;
    outputs(3919) <= not a or b;
    outputs(3920) <= b and not a;
    outputs(3921) <= b;
    outputs(3922) <= a or b;
    outputs(3923) <= a and b;
    outputs(3924) <= not a or b;
    outputs(3925) <= not a;
    outputs(3926) <= not (a xor b);
    outputs(3927) <= a;
    outputs(3928) <= not (a xor b);
    outputs(3929) <= a;
    outputs(3930) <= a and b;
    outputs(3931) <= not (a xor b);
    outputs(3932) <= not b;
    outputs(3933) <= not (a or b);
    outputs(3934) <= not (a and b);
    outputs(3935) <= a and not b;
    outputs(3936) <= not (a and b);
    outputs(3937) <= b and not a;
    outputs(3938) <= a;
    outputs(3939) <= not a;
    outputs(3940) <= not b;
    outputs(3941) <= a;
    outputs(3942) <= not (a or b);
    outputs(3943) <= not (a xor b);
    outputs(3944) <= b;
    outputs(3945) <= not (a or b);
    outputs(3946) <= a xor b;
    outputs(3947) <= a xor b;
    outputs(3948) <= not (a and b);
    outputs(3949) <= a xor b;
    outputs(3950) <= not a or b;
    outputs(3951) <= not a;
    outputs(3952) <= a;
    outputs(3953) <= b;
    outputs(3954) <= not (a xor b);
    outputs(3955) <= a xor b;
    outputs(3956) <= not a;
    outputs(3957) <= not (a or b);
    outputs(3958) <= not b;
    outputs(3959) <= not a;
    outputs(3960) <= a and b;
    outputs(3961) <= a xor b;
    outputs(3962) <= not (a or b);
    outputs(3963) <= not (a xor b);
    outputs(3964) <= not (a xor b);
    outputs(3965) <= not b;
    outputs(3966) <= a xor b;
    outputs(3967) <= b;
    outputs(3968) <= not a;
    outputs(3969) <= a xor b;
    outputs(3970) <= a xor b;
    outputs(3971) <= a xor b;
    outputs(3972) <= a xor b;
    outputs(3973) <= not b;
    outputs(3974) <= not b;
    outputs(3975) <= a xor b;
    outputs(3976) <= not b or a;
    outputs(3977) <= a and not b;
    outputs(3978) <= not (a xor b);
    outputs(3979) <= b;
    outputs(3980) <= a;
    outputs(3981) <= a xor b;
    outputs(3982) <= a;
    outputs(3983) <= b;
    outputs(3984) <= not a;
    outputs(3985) <= a and b;
    outputs(3986) <= not b;
    outputs(3987) <= a and not b;
    outputs(3988) <= not (a xor b);
    outputs(3989) <= a and not b;
    outputs(3990) <= not b or a;
    outputs(3991) <= b and not a;
    outputs(3992) <= not (a xor b);
    outputs(3993) <= a;
    outputs(3994) <= not b or a;
    outputs(3995) <= not a;
    outputs(3996) <= not a;
    outputs(3997) <= b;
    outputs(3998) <= not a or b;
    outputs(3999) <= a and b;
    outputs(4000) <= b and not a;
    outputs(4001) <= a xor b;
    outputs(4002) <= a xor b;
    outputs(4003) <= not (a or b);
    outputs(4004) <= a xor b;
    outputs(4005) <= not b;
    outputs(4006) <= not (a or b);
    outputs(4007) <= b;
    outputs(4008) <= not a;
    outputs(4009) <= not b;
    outputs(4010) <= a xor b;
    outputs(4011) <= not (a xor b);
    outputs(4012) <= a xor b;
    outputs(4013) <= b;
    outputs(4014) <= a xor b;
    outputs(4015) <= a xor b;
    outputs(4016) <= a and b;
    outputs(4017) <= not b;
    outputs(4018) <= a xor b;
    outputs(4019) <= b;
    outputs(4020) <= a;
    outputs(4021) <= a and not b;
    outputs(4022) <= b;
    outputs(4023) <= a or b;
    outputs(4024) <= b and not a;
    outputs(4025) <= not b;
    outputs(4026) <= a;
    outputs(4027) <= not a or b;
    outputs(4028) <= not a;
    outputs(4029) <= a;
    outputs(4030) <= b and not a;
    outputs(4031) <= not (a xor b);
    outputs(4032) <= a;
    outputs(4033) <= 1'b1;
    outputs(4034) <= a xor b;
    outputs(4035) <= not (a xor b);
    outputs(4036) <= a and not b;
    outputs(4037) <= b and not a;
    outputs(4038) <= not a;
    outputs(4039) <= not (a and b);
    outputs(4040) <= a or b;
    outputs(4041) <= not b or a;
    outputs(4042) <= a and not b;
    outputs(4043) <= not b or a;
    outputs(4044) <= not b or a;
    outputs(4045) <= a and not b;
    outputs(4046) <= a xor b;
    outputs(4047) <= b;
    outputs(4048) <= not a;
    outputs(4049) <= not a;
    outputs(4050) <= not b;
    outputs(4051) <= not b or a;
    outputs(4052) <= not b;
    outputs(4053) <= b;
    outputs(4054) <= a;
    outputs(4055) <= not a;
    outputs(4056) <= a;
    outputs(4057) <= not (a xor b);
    outputs(4058) <= not b or a;
    outputs(4059) <= not b or a;
    outputs(4060) <= not (a xor b);
    outputs(4061) <= b;
    outputs(4062) <= not b;
    outputs(4063) <= a or b;
    outputs(4064) <= not b;
    outputs(4065) <= a and b;
    outputs(4066) <= not b;
    outputs(4067) <= a xor b;
    outputs(4068) <= not b;
    outputs(4069) <= b;
    outputs(4070) <= b;
    outputs(4071) <= a xor b;
    outputs(4072) <= a;
    outputs(4073) <= not a or b;
    outputs(4074) <= not b;
    outputs(4075) <= not (a xor b);
    outputs(4076) <= a;
    outputs(4077) <= b and not a;
    outputs(4078) <= a xor b;
    outputs(4079) <= a xor b;
    outputs(4080) <= a;
    outputs(4081) <= not (a and b);
    outputs(4082) <= not a or b;
    outputs(4083) <= not (a and b);
    outputs(4084) <= not (a and b);
    outputs(4085) <= not a or b;
    outputs(4086) <= not (a and b);
    outputs(4087) <= not (a xor b);
    outputs(4088) <= not b;
    outputs(4089) <= a xor b;
    outputs(4090) <= b;
    outputs(4091) <= b;
    outputs(4092) <= b;
    outputs(4093) <= not (a and b);
    outputs(4094) <= b;
    outputs(4095) <= a xor b;
    outputs(4096) <= not (a xor b);
    outputs(4097) <= a and not b;
    outputs(4098) <= a and b;
    outputs(4099) <= not b;
    outputs(4100) <= a xor b;
    outputs(4101) <= not (a xor b);
    outputs(4102) <= not a;
    outputs(4103) <= a or b;
    outputs(4104) <= not (a and b);
    outputs(4105) <= a and not b;
    outputs(4106) <= a and b;
    outputs(4107) <= b;
    outputs(4108) <= b;
    outputs(4109) <= not a;
    outputs(4110) <= a xor b;
    outputs(4111) <= not b;
    outputs(4112) <= a and b;
    outputs(4113) <= a and b;
    outputs(4114) <= not (a xor b);
    outputs(4115) <= not a;
    outputs(4116) <= not (a xor b);
    outputs(4117) <= not b;
    outputs(4118) <= b;
    outputs(4119) <= a and b;
    outputs(4120) <= a xor b;
    outputs(4121) <= a xor b;
    outputs(4122) <= a xor b;
    outputs(4123) <= not b;
    outputs(4124) <= b;
    outputs(4125) <= a or b;
    outputs(4126) <= not (a or b);
    outputs(4127) <= a;
    outputs(4128) <= not a;
    outputs(4129) <= not (a or b);
    outputs(4130) <= a xor b;
    outputs(4131) <= b and not a;
    outputs(4132) <= b;
    outputs(4133) <= not (a xor b);
    outputs(4134) <= not b;
    outputs(4135) <= not (a xor b);
    outputs(4136) <= not b or a;
    outputs(4137) <= a;
    outputs(4138) <= not a;
    outputs(4139) <= a;
    outputs(4140) <= not b;
    outputs(4141) <= a or b;
    outputs(4142) <= not b or a;
    outputs(4143) <= not (a xor b);
    outputs(4144) <= not (a and b);
    outputs(4145) <= not (a xor b);
    outputs(4146) <= b;
    outputs(4147) <= b;
    outputs(4148) <= not (a xor b);
    outputs(4149) <= not (a xor b);
    outputs(4150) <= a;
    outputs(4151) <= not b;
    outputs(4152) <= not a;
    outputs(4153) <= not (a or b);
    outputs(4154) <= a and not b;
    outputs(4155) <= not a or b;
    outputs(4156) <= b and not a;
    outputs(4157) <= b;
    outputs(4158) <= a xor b;
    outputs(4159) <= not b;
    outputs(4160) <= b;
    outputs(4161) <= not (a and b);
    outputs(4162) <= a xor b;
    outputs(4163) <= not a;
    outputs(4164) <= b;
    outputs(4165) <= a xor b;
    outputs(4166) <= a and not b;
    outputs(4167) <= a xor b;
    outputs(4168) <= not a or b;
    outputs(4169) <= a;
    outputs(4170) <= a xor b;
    outputs(4171) <= not (a xor b);
    outputs(4172) <= a xor b;
    outputs(4173) <= not a or b;
    outputs(4174) <= b and not a;
    outputs(4175) <= b;
    outputs(4176) <= not (a or b);
    outputs(4177) <= a xor b;
    outputs(4178) <= not a;
    outputs(4179) <= not b or a;
    outputs(4180) <= a;
    outputs(4181) <= not b or a;
    outputs(4182) <= b;
    outputs(4183) <= not a;
    outputs(4184) <= not a or b;
    outputs(4185) <= a;
    outputs(4186) <= not b;
    outputs(4187) <= a xor b;
    outputs(4188) <= a;
    outputs(4189) <= a;
    outputs(4190) <= not a;
    outputs(4191) <= a xor b;
    outputs(4192) <= a xor b;
    outputs(4193) <= a;
    outputs(4194) <= not (a xor b);
    outputs(4195) <= not (a xor b);
    outputs(4196) <= a;
    outputs(4197) <= a xor b;
    outputs(4198) <= a xor b;
    outputs(4199) <= not (a xor b);
    outputs(4200) <= not (a and b);
    outputs(4201) <= not a;
    outputs(4202) <= not a;
    outputs(4203) <= a and not b;
    outputs(4204) <= a xor b;
    outputs(4205) <= not (a xor b);
    outputs(4206) <= b and not a;
    outputs(4207) <= not a;
    outputs(4208) <= not (a and b);
    outputs(4209) <= a xor b;
    outputs(4210) <= a and not b;
    outputs(4211) <= b;
    outputs(4212) <= a;
    outputs(4213) <= not (a or b);
    outputs(4214) <= not a;
    outputs(4215) <= a and b;
    outputs(4216) <= not a;
    outputs(4217) <= a and not b;
    outputs(4218) <= not (a xor b);
    outputs(4219) <= not (a and b);
    outputs(4220) <= b;
    outputs(4221) <= not (a xor b);
    outputs(4222) <= b;
    outputs(4223) <= not (a xor b);
    outputs(4224) <= not b;
    outputs(4225) <= not b or a;
    outputs(4226) <= a xor b;
    outputs(4227) <= a;
    outputs(4228) <= a and b;
    outputs(4229) <= not b;
    outputs(4230) <= not b;
    outputs(4231) <= not a or b;
    outputs(4232) <= a and not b;
    outputs(4233) <= not (a xor b);
    outputs(4234) <= a and b;
    outputs(4235) <= b;
    outputs(4236) <= a xor b;
    outputs(4237) <= a xor b;
    outputs(4238) <= not b;
    outputs(4239) <= a and b;
    outputs(4240) <= not a or b;
    outputs(4241) <= not a;
    outputs(4242) <= a and not b;
    outputs(4243) <= not b;
    outputs(4244) <= a;
    outputs(4245) <= not b;
    outputs(4246) <= a;
    outputs(4247) <= not (a xor b);
    outputs(4248) <= not a;
    outputs(4249) <= not (a xor b);
    outputs(4250) <= a or b;
    outputs(4251) <= a xor b;
    outputs(4252) <= b and not a;
    outputs(4253) <= a;
    outputs(4254) <= not (a and b);
    outputs(4255) <= not (a and b);
    outputs(4256) <= b and not a;
    outputs(4257) <= not b or a;
    outputs(4258) <= a and b;
    outputs(4259) <= not a;
    outputs(4260) <= not b;
    outputs(4261) <= not b;
    outputs(4262) <= a and b;
    outputs(4263) <= a xor b;
    outputs(4264) <= not (a xor b);
    outputs(4265) <= not (a xor b);
    outputs(4266) <= a or b;
    outputs(4267) <= not b;
    outputs(4268) <= not b;
    outputs(4269) <= not b or a;
    outputs(4270) <= not a;
    outputs(4271) <= b;
    outputs(4272) <= a or b;
    outputs(4273) <= a or b;
    outputs(4274) <= a;
    outputs(4275) <= not (a xor b);
    outputs(4276) <= a or b;
    outputs(4277) <= not b or a;
    outputs(4278) <= not a or b;
    outputs(4279) <= a or b;
    outputs(4280) <= a;
    outputs(4281) <= not a or b;
    outputs(4282) <= b;
    outputs(4283) <= a or b;
    outputs(4284) <= not (a or b);
    outputs(4285) <= not (a xor b);
    outputs(4286) <= a and not b;
    outputs(4287) <= b;
    outputs(4288) <= not b;
    outputs(4289) <= a and not b;
    outputs(4290) <= a and b;
    outputs(4291) <= a;
    outputs(4292) <= not (a and b);
    outputs(4293) <= not a;
    outputs(4294) <= not (a or b);
    outputs(4295) <= b;
    outputs(4296) <= not (a xor b);
    outputs(4297) <= a xor b;
    outputs(4298) <= not a or b;
    outputs(4299) <= a and not b;
    outputs(4300) <= a or b;
    outputs(4301) <= a and b;
    outputs(4302) <= not b;
    outputs(4303) <= not b;
    outputs(4304) <= a xor b;
    outputs(4305) <= a;
    outputs(4306) <= not (a or b);
    outputs(4307) <= not a;
    outputs(4308) <= a;
    outputs(4309) <= a;
    outputs(4310) <= a or b;
    outputs(4311) <= not (a xor b);
    outputs(4312) <= not b;
    outputs(4313) <= a xor b;
    outputs(4314) <= not b or a;
    outputs(4315) <= a or b;
    outputs(4316) <= a xor b;
    outputs(4317) <= a and b;
    outputs(4318) <= a or b;
    outputs(4319) <= not a;
    outputs(4320) <= not b or a;
    outputs(4321) <= a and not b;
    outputs(4322) <= a or b;
    outputs(4323) <= a or b;
    outputs(4324) <= not (a and b);
    outputs(4325) <= a xor b;
    outputs(4326) <= b;
    outputs(4327) <= not (a and b);
    outputs(4328) <= b;
    outputs(4329) <= a and not b;
    outputs(4330) <= a xor b;
    outputs(4331) <= b;
    outputs(4332) <= not a;
    outputs(4333) <= a xor b;
    outputs(4334) <= not b;
    outputs(4335) <= a and b;
    outputs(4336) <= not (a xor b);
    outputs(4337) <= not (a and b);
    outputs(4338) <= not (a and b);
    outputs(4339) <= a xor b;
    outputs(4340) <= a xor b;
    outputs(4341) <= a xor b;
    outputs(4342) <= b and not a;
    outputs(4343) <= not (a or b);
    outputs(4344) <= not (a and b);
    outputs(4345) <= not b or a;
    outputs(4346) <= a and b;
    outputs(4347) <= not (a xor b);
    outputs(4348) <= not a;
    outputs(4349) <= b;
    outputs(4350) <= not (a or b);
    outputs(4351) <= a xor b;
    outputs(4352) <= not a or b;
    outputs(4353) <= a and b;
    outputs(4354) <= b;
    outputs(4355) <= not (a xor b);
    outputs(4356) <= a;
    outputs(4357) <= a xor b;
    outputs(4358) <= not (a xor b);
    outputs(4359) <= b;
    outputs(4360) <= a xor b;
    outputs(4361) <= a;
    outputs(4362) <= a xor b;
    outputs(4363) <= not (a xor b);
    outputs(4364) <= a or b;
    outputs(4365) <= not a or b;
    outputs(4366) <= not (a and b);
    outputs(4367) <= a;
    outputs(4368) <= a;
    outputs(4369) <= not b;
    outputs(4370) <= not (a or b);
    outputs(4371) <= a xor b;
    outputs(4372) <= not (a and b);
    outputs(4373) <= not b;
    outputs(4374) <= not (a xor b);
    outputs(4375) <= not b;
    outputs(4376) <= b and not a;
    outputs(4377) <= a;
    outputs(4378) <= a and b;
    outputs(4379) <= not a or b;
    outputs(4380) <= a xor b;
    outputs(4381) <= a;
    outputs(4382) <= a and b;
    outputs(4383) <= a;
    outputs(4384) <= a and b;
    outputs(4385) <= a and b;
    outputs(4386) <= not a;
    outputs(4387) <= not a or b;
    outputs(4388) <= not a or b;
    outputs(4389) <= b;
    outputs(4390) <= b;
    outputs(4391) <= a;
    outputs(4392) <= a xor b;
    outputs(4393) <= not (a xor b);
    outputs(4394) <= not (a xor b);
    outputs(4395) <= not (a or b);
    outputs(4396) <= not a or b;
    outputs(4397) <= not b;
    outputs(4398) <= a xor b;
    outputs(4399) <= a xor b;
    outputs(4400) <= b;
    outputs(4401) <= not (a xor b);
    outputs(4402) <= not b or a;
    outputs(4403) <= a xor b;
    outputs(4404) <= a and not b;
    outputs(4405) <= b;
    outputs(4406) <= not (a xor b);
    outputs(4407) <= a xor b;
    outputs(4408) <= not (a xor b);
    outputs(4409) <= a or b;
    outputs(4410) <= not (a xor b);
    outputs(4411) <= a and b;
    outputs(4412) <= not a or b;
    outputs(4413) <= a;
    outputs(4414) <= not (a xor b);
    outputs(4415) <= a xor b;
    outputs(4416) <= a xor b;
    outputs(4417) <= a;
    outputs(4418) <= not b;
    outputs(4419) <= not (a and b);
    outputs(4420) <= not b or a;
    outputs(4421) <= not (a or b);
    outputs(4422) <= a and not b;
    outputs(4423) <= a;
    outputs(4424) <= not a;
    outputs(4425) <= not (a xor b);
    outputs(4426) <= b and not a;
    outputs(4427) <= not a;
    outputs(4428) <= not (a xor b);
    outputs(4429) <= b;
    outputs(4430) <= a and not b;
    outputs(4431) <= not a;
    outputs(4432) <= a or b;
    outputs(4433) <= a and b;
    outputs(4434) <= not a;
    outputs(4435) <= b;
    outputs(4436) <= b and not a;
    outputs(4437) <= not (a or b);
    outputs(4438) <= a;
    outputs(4439) <= a xor b;
    outputs(4440) <= a and b;
    outputs(4441) <= not a or b;
    outputs(4442) <= not a;
    outputs(4443) <= a or b;
    outputs(4444) <= not (a xor b);
    outputs(4445) <= not b;
    outputs(4446) <= not a;
    outputs(4447) <= a or b;
    outputs(4448) <= not (a xor b);
    outputs(4449) <= a and not b;
    outputs(4450) <= a and not b;
    outputs(4451) <= not (a xor b);
    outputs(4452) <= a;
    outputs(4453) <= b and not a;
    outputs(4454) <= not b;
    outputs(4455) <= a and b;
    outputs(4456) <= b and not a;
    outputs(4457) <= b;
    outputs(4458) <= not (a xor b);
    outputs(4459) <= a xor b;
    outputs(4460) <= not b or a;
    outputs(4461) <= a or b;
    outputs(4462) <= a;
    outputs(4463) <= not a;
    outputs(4464) <= not a or b;
    outputs(4465) <= b and not a;
    outputs(4466) <= not (a and b);
    outputs(4467) <= b;
    outputs(4468) <= a xor b;
    outputs(4469) <= b;
    outputs(4470) <= not (a xor b);
    outputs(4471) <= not a;
    outputs(4472) <= not (a xor b);
    outputs(4473) <= b;
    outputs(4474) <= not (a xor b);
    outputs(4475) <= not b;
    outputs(4476) <= not a or b;
    outputs(4477) <= b;
    outputs(4478) <= a;
    outputs(4479) <= not (a xor b);
    outputs(4480) <= b and not a;
    outputs(4481) <= not (a xor b);
    outputs(4482) <= b and not a;
    outputs(4483) <= not b or a;
    outputs(4484) <= a xor b;
    outputs(4485) <= a and not b;
    outputs(4486) <= not b;
    outputs(4487) <= not (a or b);
    outputs(4488) <= b;
    outputs(4489) <= a xor b;
    outputs(4490) <= not a;
    outputs(4491) <= a and b;
    outputs(4492) <= not (a or b);
    outputs(4493) <= not (a and b);
    outputs(4494) <= not (a and b);
    outputs(4495) <= a;
    outputs(4496) <= a xor b;
    outputs(4497) <= not a or b;
    outputs(4498) <= b;
    outputs(4499) <= b;
    outputs(4500) <= not (a xor b);
    outputs(4501) <= not (a xor b);
    outputs(4502) <= not b;
    outputs(4503) <= a and b;
    outputs(4504) <= not a;
    outputs(4505) <= not (a xor b);
    outputs(4506) <= not (a or b);
    outputs(4507) <= not a or b;
    outputs(4508) <= a;
    outputs(4509) <= not a;
    outputs(4510) <= a;
    outputs(4511) <= a and b;
    outputs(4512) <= not (a xor b);
    outputs(4513) <= a and b;
    outputs(4514) <= a and b;
    outputs(4515) <= not (a xor b);
    outputs(4516) <= not (a xor b);
    outputs(4517) <= a and b;
    outputs(4518) <= a and b;
    outputs(4519) <= a xor b;
    outputs(4520) <= not b;
    outputs(4521) <= a and not b;
    outputs(4522) <= a and b;
    outputs(4523) <= a and b;
    outputs(4524) <= not (a xor b);
    outputs(4525) <= a;
    outputs(4526) <= a or b;
    outputs(4527) <= a;
    outputs(4528) <= b;
    outputs(4529) <= not b or a;
    outputs(4530) <= a xor b;
    outputs(4531) <= b;
    outputs(4532) <= b;
    outputs(4533) <= not a or b;
    outputs(4534) <= a and not b;
    outputs(4535) <= not b;
    outputs(4536) <= not (a or b);
    outputs(4537) <= a;
    outputs(4538) <= a;
    outputs(4539) <= not b;
    outputs(4540) <= not (a and b);
    outputs(4541) <= not b or a;
    outputs(4542) <= not (a or b);
    outputs(4543) <= not a or b;
    outputs(4544) <= a xor b;
    outputs(4545) <= b;
    outputs(4546) <= not b;
    outputs(4547) <= a and b;
    outputs(4548) <= a;
    outputs(4549) <= not (a or b);
    outputs(4550) <= a or b;
    outputs(4551) <= not b or a;
    outputs(4552) <= a and b;
    outputs(4553) <= b;
    outputs(4554) <= a;
    outputs(4555) <= a;
    outputs(4556) <= b and not a;
    outputs(4557) <= a or b;
    outputs(4558) <= a or b;
    outputs(4559) <= not (a or b);
    outputs(4560) <= a and b;
    outputs(4561) <= a or b;
    outputs(4562) <= not a or b;
    outputs(4563) <= not b;
    outputs(4564) <= a;
    outputs(4565) <= b and not a;
    outputs(4566) <= a xor b;
    outputs(4567) <= a;
    outputs(4568) <= not a;
    outputs(4569) <= b;
    outputs(4570) <= not (a xor b);
    outputs(4571) <= not a;
    outputs(4572) <= b and not a;
    outputs(4573) <= not b;
    outputs(4574) <= a xor b;
    outputs(4575) <= not a;
    outputs(4576) <= a xor b;
    outputs(4577) <= not b or a;
    outputs(4578) <= a xor b;
    outputs(4579) <= a;
    outputs(4580) <= a;
    outputs(4581) <= a xor b;
    outputs(4582) <= not (a xor b);
    outputs(4583) <= a or b;
    outputs(4584) <= b and not a;
    outputs(4585) <= b;
    outputs(4586) <= b;
    outputs(4587) <= b and not a;
    outputs(4588) <= a and b;
    outputs(4589) <= not b;
    outputs(4590) <= b and not a;
    outputs(4591) <= not a;
    outputs(4592) <= not a or b;
    outputs(4593) <= not (a xor b);
    outputs(4594) <= not (a xor b);
    outputs(4595) <= a and not b;
    outputs(4596) <= a and not b;
    outputs(4597) <= not b;
    outputs(4598) <= a;
    outputs(4599) <= not (a xor b);
    outputs(4600) <= not b;
    outputs(4601) <= not a;
    outputs(4602) <= b and not a;
    outputs(4603) <= b;
    outputs(4604) <= a and not b;
    outputs(4605) <= b and not a;
    outputs(4606) <= not a or b;
    outputs(4607) <= a and b;
    outputs(4608) <= a and not b;
    outputs(4609) <= not b;
    outputs(4610) <= b and not a;
    outputs(4611) <= not (a xor b);
    outputs(4612) <= not (a xor b);
    outputs(4613) <= not (a or b);
    outputs(4614) <= not (a or b);
    outputs(4615) <= not (a or b);
    outputs(4616) <= a and not b;
    outputs(4617) <= not (a or b);
    outputs(4618) <= not (a or b);
    outputs(4619) <= not (a xor b);
    outputs(4620) <= not b;
    outputs(4621) <= a xor b;
    outputs(4622) <= not b;
    outputs(4623) <= not (a and b);
    outputs(4624) <= b and not a;
    outputs(4625) <= a or b;
    outputs(4626) <= a;
    outputs(4627) <= a and not b;
    outputs(4628) <= b and not a;
    outputs(4629) <= not b;
    outputs(4630) <= a xor b;
    outputs(4631) <= not (a or b);
    outputs(4632) <= a xor b;
    outputs(4633) <= not a;
    outputs(4634) <= not (a xor b);
    outputs(4635) <= b and not a;
    outputs(4636) <= not (a xor b);
    outputs(4637) <= not (a and b);
    outputs(4638) <= not (a and b);
    outputs(4639) <= b;
    outputs(4640) <= not (a xor b);
    outputs(4641) <= a and b;
    outputs(4642) <= a;
    outputs(4643) <= a;
    outputs(4644) <= a;
    outputs(4645) <= not b;
    outputs(4646) <= not a;
    outputs(4647) <= not (a and b);
    outputs(4648) <= b and not a;
    outputs(4649) <= not a;
    outputs(4650) <= not a;
    outputs(4651) <= not (a xor b);
    outputs(4652) <= a and b;
    outputs(4653) <= not b;
    outputs(4654) <= not (a xor b);
    outputs(4655) <= not (a or b);
    outputs(4656) <= not (a or b);
    outputs(4657) <= not a;
    outputs(4658) <= a and b;
    outputs(4659) <= b and not a;
    outputs(4660) <= a xor b;
    outputs(4661) <= not b;
    outputs(4662) <= b and not a;
    outputs(4663) <= a and b;
    outputs(4664) <= a and not b;
    outputs(4665) <= a or b;
    outputs(4666) <= a and not b;
    outputs(4667) <= a xor b;
    outputs(4668) <= b;
    outputs(4669) <= not (a or b);
    outputs(4670) <= b;
    outputs(4671) <= b;
    outputs(4672) <= a xor b;
    outputs(4673) <= not b or a;
    outputs(4674) <= a and b;
    outputs(4675) <= a;
    outputs(4676) <= a and b;
    outputs(4677) <= a;
    outputs(4678) <= a or b;
    outputs(4679) <= not b;
    outputs(4680) <= not (a and b);
    outputs(4681) <= a xor b;
    outputs(4682) <= b;
    outputs(4683) <= not (a or b);
    outputs(4684) <= a or b;
    outputs(4685) <= not a;
    outputs(4686) <= not (a or b);
    outputs(4687) <= a xor b;
    outputs(4688) <= not a or b;
    outputs(4689) <= a xor b;
    outputs(4690) <= a;
    outputs(4691) <= not b;
    outputs(4692) <= not (a or b);
    outputs(4693) <= not (a and b);
    outputs(4694) <= not b;
    outputs(4695) <= not b;
    outputs(4696) <= not b;
    outputs(4697) <= not a;
    outputs(4698) <= b and not a;
    outputs(4699) <= not a;
    outputs(4700) <= not (a xor b);
    outputs(4701) <= not a;
    outputs(4702) <= not b;
    outputs(4703) <= not a;
    outputs(4704) <= a or b;
    outputs(4705) <= a xor b;
    outputs(4706) <= a and not b;
    outputs(4707) <= a xor b;
    outputs(4708) <= not b;
    outputs(4709) <= a;
    outputs(4710) <= a and not b;
    outputs(4711) <= not a;
    outputs(4712) <= a and not b;
    outputs(4713) <= not b;
    outputs(4714) <= a;
    outputs(4715) <= a or b;
    outputs(4716) <= b and not a;
    outputs(4717) <= b and not a;
    outputs(4718) <= not b or a;
    outputs(4719) <= not (a or b);
    outputs(4720) <= b and not a;
    outputs(4721) <= b;
    outputs(4722) <= not a or b;
    outputs(4723) <= a;
    outputs(4724) <= not (a or b);
    outputs(4725) <= a;
    outputs(4726) <= a xor b;
    outputs(4727) <= not (a or b);
    outputs(4728) <= a and not b;
    outputs(4729) <= b;
    outputs(4730) <= not a or b;
    outputs(4731) <= a xor b;
    outputs(4732) <= a and not b;
    outputs(4733) <= not (a xor b);
    outputs(4734) <= not a;
    outputs(4735) <= not a;
    outputs(4736) <= a or b;
    outputs(4737) <= a and not b;
    outputs(4738) <= not a;
    outputs(4739) <= not a;
    outputs(4740) <= b and not a;
    outputs(4741) <= not (a or b);
    outputs(4742) <= not (a xor b);
    outputs(4743) <= a xor b;
    outputs(4744) <= a or b;
    outputs(4745) <= a and not b;
    outputs(4746) <= not b or a;
    outputs(4747) <= not a;
    outputs(4748) <= not (a xor b);
    outputs(4749) <= a and b;
    outputs(4750) <= not (a xor b);
    outputs(4751) <= not (a xor b);
    outputs(4752) <= b;
    outputs(4753) <= not a;
    outputs(4754) <= not b;
    outputs(4755) <= b;
    outputs(4756) <= not a;
    outputs(4757) <= a;
    outputs(4758) <= b;
    outputs(4759) <= b and not a;
    outputs(4760) <= a and b;
    outputs(4761) <= not a;
    outputs(4762) <= a or b;
    outputs(4763) <= a xor b;
    outputs(4764) <= b and not a;
    outputs(4765) <= b;
    outputs(4766) <= not a;
    outputs(4767) <= not b;
    outputs(4768) <= a and not b;
    outputs(4769) <= b;
    outputs(4770) <= not a or b;
    outputs(4771) <= not a or b;
    outputs(4772) <= not b;
    outputs(4773) <= a xor b;
    outputs(4774) <= a xor b;
    outputs(4775) <= not (a xor b);
    outputs(4776) <= b and not a;
    outputs(4777) <= not (a xor b);
    outputs(4778) <= not b;
    outputs(4779) <= not b or a;
    outputs(4780) <= not (a xor b);
    outputs(4781) <= not (a xor b);
    outputs(4782) <= not (a or b);
    outputs(4783) <= not a;
    outputs(4784) <= not (a xor b);
    outputs(4785) <= b;
    outputs(4786) <= b;
    outputs(4787) <= a and not b;
    outputs(4788) <= a and not b;
    outputs(4789) <= a and b;
    outputs(4790) <= not b;
    outputs(4791) <= a;
    outputs(4792) <= not (a xor b);
    outputs(4793) <= not (a xor b);
    outputs(4794) <= not a;
    outputs(4795) <= a;
    outputs(4796) <= a and not b;
    outputs(4797) <= a and b;
    outputs(4798) <= a and b;
    outputs(4799) <= not (a xor b);
    outputs(4800) <= not b;
    outputs(4801) <= b;
    outputs(4802) <= not (a xor b);
    outputs(4803) <= not (a or b);
    outputs(4804) <= not (a xor b);
    outputs(4805) <= b;
    outputs(4806) <= not b;
    outputs(4807) <= not b;
    outputs(4808) <= not (a xor b);
    outputs(4809) <= a;
    outputs(4810) <= b;
    outputs(4811) <= a and not b;
    outputs(4812) <= b and not a;
    outputs(4813) <= not b or a;
    outputs(4814) <= not a;
    outputs(4815) <= not b;
    outputs(4816) <= not a;
    outputs(4817) <= a and b;
    outputs(4818) <= not a or b;
    outputs(4819) <= a;
    outputs(4820) <= a xor b;
    outputs(4821) <= not a;
    outputs(4822) <= not a;
    outputs(4823) <= not (a and b);
    outputs(4824) <= not (a and b);
    outputs(4825) <= not (a or b);
    outputs(4826) <= a and not b;
    outputs(4827) <= a and b;
    outputs(4828) <= not a;
    outputs(4829) <= a;
    outputs(4830) <= a or b;
    outputs(4831) <= not a;
    outputs(4832) <= b and not a;
    outputs(4833) <= b and not a;
    outputs(4834) <= not b;
    outputs(4835) <= a or b;
    outputs(4836) <= a and b;
    outputs(4837) <= not b;
    outputs(4838) <= a xor b;
    outputs(4839) <= a and b;
    outputs(4840) <= a and not b;
    outputs(4841) <= not (a and b);
    outputs(4842) <= not b or a;
    outputs(4843) <= not (a and b);
    outputs(4844) <= not (a or b);
    outputs(4845) <= not (a or b);
    outputs(4846) <= not (a and b);
    outputs(4847) <= not b;
    outputs(4848) <= not (a xor b);
    outputs(4849) <= a and b;
    outputs(4850) <= not (a xor b);
    outputs(4851) <= a and not b;
    outputs(4852) <= not (a or b);
    outputs(4853) <= a and b;
    outputs(4854) <= not (a or b);
    outputs(4855) <= not a;
    outputs(4856) <= not (a xor b);
    outputs(4857) <= not a;
    outputs(4858) <= a xor b;
    outputs(4859) <= not b;
    outputs(4860) <= not (a and b);
    outputs(4861) <= b;
    outputs(4862) <= b;
    outputs(4863) <= not (a xor b);
    outputs(4864) <= b;
    outputs(4865) <= b and not a;
    outputs(4866) <= not b;
    outputs(4867) <= not (a or b);
    outputs(4868) <= not (a and b);
    outputs(4869) <= a and b;
    outputs(4870) <= not (a and b);
    outputs(4871) <= not (a or b);
    outputs(4872) <= not (a or b);
    outputs(4873) <= a;
    outputs(4874) <= not (a or b);
    outputs(4875) <= a and not b;
    outputs(4876) <= not (a xor b);
    outputs(4877) <= a and not b;
    outputs(4878) <= not (a and b);
    outputs(4879) <= a and not b;
    outputs(4880) <= b and not a;
    outputs(4881) <= not (a xor b);
    outputs(4882) <= a xor b;
    outputs(4883) <= not (a xor b);
    outputs(4884) <= not (a xor b);
    outputs(4885) <= not b;
    outputs(4886) <= a;
    outputs(4887) <= b;
    outputs(4888) <= not (a xor b);
    outputs(4889) <= not b or a;
    outputs(4890) <= b;
    outputs(4891) <= b and not a;
    outputs(4892) <= b;
    outputs(4893) <= a and not b;
    outputs(4894) <= a or b;
    outputs(4895) <= b and not a;
    outputs(4896) <= not a;
    outputs(4897) <= a and b;
    outputs(4898) <= a xor b;
    outputs(4899) <= b;
    outputs(4900) <= a xor b;
    outputs(4901) <= a xor b;
    outputs(4902) <= not b;
    outputs(4903) <= a xor b;
    outputs(4904) <= not b;
    outputs(4905) <= not a;
    outputs(4906) <= not (a or b);
    outputs(4907) <= a xor b;
    outputs(4908) <= b;
    outputs(4909) <= b;
    outputs(4910) <= a;
    outputs(4911) <= not a;
    outputs(4912) <= not b;
    outputs(4913) <= b;
    outputs(4914) <= not a;
    outputs(4915) <= not b;
    outputs(4916) <= not a;
    outputs(4917) <= not (a xor b);
    outputs(4918) <= not (a or b);
    outputs(4919) <= b;
    outputs(4920) <= not b;
    outputs(4921) <= a;
    outputs(4922) <= a;
    outputs(4923) <= a or b;
    outputs(4924) <= not b;
    outputs(4925) <= b and not a;
    outputs(4926) <= b;
    outputs(4927) <= not a;
    outputs(4928) <= b;
    outputs(4929) <= b and not a;
    outputs(4930) <= a;
    outputs(4931) <= b and not a;
    outputs(4932) <= a;
    outputs(4933) <= a;
    outputs(4934) <= a and not b;
    outputs(4935) <= not (a xor b);
    outputs(4936) <= a;
    outputs(4937) <= a;
    outputs(4938) <= not (a xor b);
    outputs(4939) <= not (a and b);
    outputs(4940) <= a xor b;
    outputs(4941) <= not b;
    outputs(4942) <= not a or b;
    outputs(4943) <= a and not b;
    outputs(4944) <= a and not b;
    outputs(4945) <= not a;
    outputs(4946) <= not (a or b);
    outputs(4947) <= a or b;
    outputs(4948) <= a;
    outputs(4949) <= a and not b;
    outputs(4950) <= b;
    outputs(4951) <= a;
    outputs(4952) <= not (a xor b);
    outputs(4953) <= not a;
    outputs(4954) <= not (a xor b);
    outputs(4955) <= b;
    outputs(4956) <= not b;
    outputs(4957) <= not a;
    outputs(4958) <= b;
    outputs(4959) <= a xor b;
    outputs(4960) <= not (a and b);
    outputs(4961) <= a or b;
    outputs(4962) <= b;
    outputs(4963) <= b;
    outputs(4964) <= not a or b;
    outputs(4965) <= not b;
    outputs(4966) <= a and b;
    outputs(4967) <= b;
    outputs(4968) <= not (a xor b);
    outputs(4969) <= not (a xor b);
    outputs(4970) <= a and b;
    outputs(4971) <= a and not b;
    outputs(4972) <= b and not a;
    outputs(4973) <= not (a xor b);
    outputs(4974) <= not b;
    outputs(4975) <= not a;
    outputs(4976) <= not b or a;
    outputs(4977) <= a and b;
    outputs(4978) <= a and not b;
    outputs(4979) <= not a;
    outputs(4980) <= a or b;
    outputs(4981) <= not b;
    outputs(4982) <= b and not a;
    outputs(4983) <= b;
    outputs(4984) <= not (a or b);
    outputs(4985) <= a and b;
    outputs(4986) <= not (a xor b);
    outputs(4987) <= a;
    outputs(4988) <= a or b;
    outputs(4989) <= not b;
    outputs(4990) <= not (a or b);
    outputs(4991) <= not (a xor b);
    outputs(4992) <= not (a xor b);
    outputs(4993) <= not a;
    outputs(4994) <= not (a or b);
    outputs(4995) <= b and not a;
    outputs(4996) <= a xor b;
    outputs(4997) <= not b;
    outputs(4998) <= not (a xor b);
    outputs(4999) <= a xor b;
    outputs(5000) <= not (a or b);
    outputs(5001) <= b;
    outputs(5002) <= a and not b;
    outputs(5003) <= a;
    outputs(5004) <= a;
    outputs(5005) <= not a;
    outputs(5006) <= a and b;
    outputs(5007) <= a and b;
    outputs(5008) <= not (a xor b);
    outputs(5009) <= not (a or b);
    outputs(5010) <= a xor b;
    outputs(5011) <= not (a xor b);
    outputs(5012) <= a and not b;
    outputs(5013) <= not a or b;
    outputs(5014) <= not (a and b);
    outputs(5015) <= a;
    outputs(5016) <= not (a xor b);
    outputs(5017) <= b;
    outputs(5018) <= a and not b;
    outputs(5019) <= not b;
    outputs(5020) <= not b;
    outputs(5021) <= a and b;
    outputs(5022) <= a or b;
    outputs(5023) <= a and not b;
    outputs(5024) <= not (a xor b);
    outputs(5025) <= not (a xor b);
    outputs(5026) <= not (a or b);
    outputs(5027) <= not b;
    outputs(5028) <= not b or a;
    outputs(5029) <= b and not a;
    outputs(5030) <= a xor b;
    outputs(5031) <= a and not b;
    outputs(5032) <= b;
    outputs(5033) <= a and b;
    outputs(5034) <= a;
    outputs(5035) <= a or b;
    outputs(5036) <= a and not b;
    outputs(5037) <= a and b;
    outputs(5038) <= a and not b;
    outputs(5039) <= not a;
    outputs(5040) <= a xor b;
    outputs(5041) <= a;
    outputs(5042) <= not a;
    outputs(5043) <= not a or b;
    outputs(5044) <= not a;
    outputs(5045) <= not a;
    outputs(5046) <= b and not a;
    outputs(5047) <= a or b;
    outputs(5048) <= a or b;
    outputs(5049) <= b;
    outputs(5050) <= not (a and b);
    outputs(5051) <= a xor b;
    outputs(5052) <= not a or b;
    outputs(5053) <= a and b;
    outputs(5054) <= not (a xor b);
    outputs(5055) <= b and not a;
    outputs(5056) <= not (a or b);
    outputs(5057) <= a;
    outputs(5058) <= not a;
    outputs(5059) <= a xor b;
    outputs(5060) <= not a;
    outputs(5061) <= not a;
    outputs(5062) <= a or b;
    outputs(5063) <= a and b;
    outputs(5064) <= a and not b;
    outputs(5065) <= a;
    outputs(5066) <= 1'b0;
    outputs(5067) <= a and not b;
    outputs(5068) <= a xor b;
    outputs(5069) <= b;
    outputs(5070) <= a xor b;
    outputs(5071) <= a and not b;
    outputs(5072) <= not a;
    outputs(5073) <= a or b;
    outputs(5074) <= not (a xor b);
    outputs(5075) <= not (a xor b);
    outputs(5076) <= not a;
    outputs(5077) <= a xor b;
    outputs(5078) <= not (a xor b);
    outputs(5079) <= not (a xor b);
    outputs(5080) <= not a;
    outputs(5081) <= a xor b;
    outputs(5082) <= b and not a;
    outputs(5083) <= not a;
    outputs(5084) <= b and not a;
    outputs(5085) <= not (a xor b);
    outputs(5086) <= a xor b;
    outputs(5087) <= not a;
    outputs(5088) <= a and not b;
    outputs(5089) <= not (a and b);
    outputs(5090) <= a and b;
    outputs(5091) <= not (a xor b);
    outputs(5092) <= not (a xor b);
    outputs(5093) <= a and b;
    outputs(5094) <= a and not b;
    outputs(5095) <= a and not b;
    outputs(5096) <= b and not a;
    outputs(5097) <= not a or b;
    outputs(5098) <= b;
    outputs(5099) <= a xor b;
    outputs(5100) <= a xor b;
    outputs(5101) <= not b;
    outputs(5102) <= a xor b;
    outputs(5103) <= not (a and b);
    outputs(5104) <= not a;
    outputs(5105) <= a xor b;
    outputs(5106) <= not b;
    outputs(5107) <= not (a or b);
    outputs(5108) <= not (a or b);
    outputs(5109) <= a;
    outputs(5110) <= not b;
    outputs(5111) <= not b;
    outputs(5112) <= not a or b;
    outputs(5113) <= not b;
    outputs(5114) <= a and not b;
    outputs(5115) <= not a or b;
    outputs(5116) <= b and not a;
    outputs(5117) <= not (a xor b);
    outputs(5118) <= not a or b;
    outputs(5119) <= b;
    outputs(5120) <= not (a xor b);
    outputs(5121) <= a and b;
    outputs(5122) <= not (a xor b);
    outputs(5123) <= a or b;
    outputs(5124) <= not b;
    outputs(5125) <= not (a or b);
    outputs(5126) <= not b or a;
    outputs(5127) <= b and not a;
    outputs(5128) <= not b or a;
    outputs(5129) <= a and b;
    outputs(5130) <= a;
    outputs(5131) <= a and not b;
    outputs(5132) <= not (a xor b);
    outputs(5133) <= a xor b;
    outputs(5134) <= a and not b;
    outputs(5135) <= a and not b;
    outputs(5136) <= not (a or b);
    outputs(5137) <= a and b;
    outputs(5138) <= b;
    outputs(5139) <= not b or a;
    outputs(5140) <= not b;
    outputs(5141) <= a xor b;
    outputs(5142) <= not a;
    outputs(5143) <= not b;
    outputs(5144) <= a;
    outputs(5145) <= not (a and b);
    outputs(5146) <= a and not b;
    outputs(5147) <= not (a or b);
    outputs(5148) <= a;
    outputs(5149) <= not b;
    outputs(5150) <= not (a or b);
    outputs(5151) <= a or b;
    outputs(5152) <= not a;
    outputs(5153) <= not a;
    outputs(5154) <= not b;
    outputs(5155) <= a xor b;
    outputs(5156) <= a and not b;
    outputs(5157) <= b and not a;
    outputs(5158) <= not b;
    outputs(5159) <= not (a xor b);
    outputs(5160) <= not (a xor b);
    outputs(5161) <= a and b;
    outputs(5162) <= b;
    outputs(5163) <= not (a xor b);
    outputs(5164) <= not (a or b);
    outputs(5165) <= not (a and b);
    outputs(5166) <= a;
    outputs(5167) <= 1'b0;
    outputs(5168) <= a xor b;
    outputs(5169) <= a xor b;
    outputs(5170) <= not b;
    outputs(5171) <= not b;
    outputs(5172) <= a xor b;
    outputs(5173) <= not a;
    outputs(5174) <= b and not a;
    outputs(5175) <= not (a xor b);
    outputs(5176) <= not b or a;
    outputs(5177) <= a or b;
    outputs(5178) <= a xor b;
    outputs(5179) <= b;
    outputs(5180) <= a xor b;
    outputs(5181) <= b;
    outputs(5182) <= a and not b;
    outputs(5183) <= a and not b;
    outputs(5184) <= not b;
    outputs(5185) <= not (a or b);
    outputs(5186) <= b and not a;
    outputs(5187) <= a;
    outputs(5188) <= b and not a;
    outputs(5189) <= a;
    outputs(5190) <= not (a xor b);
    outputs(5191) <= a xor b;
    outputs(5192) <= not b;
    outputs(5193) <= not a;
    outputs(5194) <= a;
    outputs(5195) <= b;
    outputs(5196) <= not (a xor b);
    outputs(5197) <= a xor b;
    outputs(5198) <= b and not a;
    outputs(5199) <= a xor b;
    outputs(5200) <= not (a xor b);
    outputs(5201) <= not a;
    outputs(5202) <= not b;
    outputs(5203) <= a and not b;
    outputs(5204) <= b;
    outputs(5205) <= a;
    outputs(5206) <= a xor b;
    outputs(5207) <= not (a xor b);
    outputs(5208) <= not (a and b);
    outputs(5209) <= not b;
    outputs(5210) <= not (a and b);
    outputs(5211) <= b and not a;
    outputs(5212) <= not (a or b);
    outputs(5213) <= b;
    outputs(5214) <= not a;
    outputs(5215) <= not b;
    outputs(5216) <= a;
    outputs(5217) <= not (a xor b);
    outputs(5218) <= a and b;
    outputs(5219) <= a;
    outputs(5220) <= a xor b;
    outputs(5221) <= not (a and b);
    outputs(5222) <= b;
    outputs(5223) <= a and not b;
    outputs(5224) <= a xor b;
    outputs(5225) <= not a;
    outputs(5226) <= not (a and b);
    outputs(5227) <= not (a and b);
    outputs(5228) <= not b or a;
    outputs(5229) <= b;
    outputs(5230) <= not (a xor b);
    outputs(5231) <= not (a xor b);
    outputs(5232) <= not b;
    outputs(5233) <= b and not a;
    outputs(5234) <= a and b;
    outputs(5235) <= not a;
    outputs(5236) <= b;
    outputs(5237) <= a;
    outputs(5238) <= not (a xor b);
    outputs(5239) <= not a;
    outputs(5240) <= b and not a;
    outputs(5241) <= a or b;
    outputs(5242) <= not (a or b);
    outputs(5243) <= b;
    outputs(5244) <= b;
    outputs(5245) <= not b or a;
    outputs(5246) <= not (a or b);
    outputs(5247) <= not (a xor b);
    outputs(5248) <= not (a or b);
    outputs(5249) <= a xor b;
    outputs(5250) <= a and b;
    outputs(5251) <= not (a or b);
    outputs(5252) <= not (a or b);
    outputs(5253) <= not b;
    outputs(5254) <= b;
    outputs(5255) <= not (a xor b);
    outputs(5256) <= not (a or b);
    outputs(5257) <= not (a xor b);
    outputs(5258) <= a and b;
    outputs(5259) <= b;
    outputs(5260) <= not (a xor b);
    outputs(5261) <= b and not a;
    outputs(5262) <= a xor b;
    outputs(5263) <= b;
    outputs(5264) <= not a;
    outputs(5265) <= a xor b;
    outputs(5266) <= not (a xor b);
    outputs(5267) <= not b;
    outputs(5268) <= not b or a;
    outputs(5269) <= b;
    outputs(5270) <= b;
    outputs(5271) <= a xor b;
    outputs(5272) <= not b or a;
    outputs(5273) <= b;
    outputs(5274) <= b and not a;
    outputs(5275) <= not (a or b);
    outputs(5276) <= b;
    outputs(5277) <= a xor b;
    outputs(5278) <= not b;
    outputs(5279) <= a;
    outputs(5280) <= b;
    outputs(5281) <= not a;
    outputs(5282) <= not (a xor b);
    outputs(5283) <= not b or a;
    outputs(5284) <= a;
    outputs(5285) <= not (a and b);
    outputs(5286) <= not (a or b);
    outputs(5287) <= a xor b;
    outputs(5288) <= not (a or b);
    outputs(5289) <= a or b;
    outputs(5290) <= not (a or b);
    outputs(5291) <= a xor b;
    outputs(5292) <= not (a and b);
    outputs(5293) <= not b;
    outputs(5294) <= not (a xor b);
    outputs(5295) <= not a;
    outputs(5296) <= not (a xor b);
    outputs(5297) <= not (a xor b);
    outputs(5298) <= a;
    outputs(5299) <= not (a xor b);
    outputs(5300) <= not (a and b);
    outputs(5301) <= not b;
    outputs(5302) <= a and b;
    outputs(5303) <= not a;
    outputs(5304) <= not a;
    outputs(5305) <= not (a and b);
    outputs(5306) <= b;
    outputs(5307) <= a or b;
    outputs(5308) <= not a;
    outputs(5309) <= not b or a;
    outputs(5310) <= b and not a;
    outputs(5311) <= not (a or b);
    outputs(5312) <= not a;
    outputs(5313) <= not (a xor b);
    outputs(5314) <= a;
    outputs(5315) <= not b;
    outputs(5316) <= not (a or b);
    outputs(5317) <= a xor b;
    outputs(5318) <= not a;
    outputs(5319) <= not b;
    outputs(5320) <= not b or a;
    outputs(5321) <= a and not b;
    outputs(5322) <= a and b;
    outputs(5323) <= b and not a;
    outputs(5324) <= b and not a;
    outputs(5325) <= not b;
    outputs(5326) <= b;
    outputs(5327) <= a or b;
    outputs(5328) <= not (a or b);
    outputs(5329) <= a and not b;
    outputs(5330) <= not b;
    outputs(5331) <= b;
    outputs(5332) <= not (a xor b);
    outputs(5333) <= not a or b;
    outputs(5334) <= b;
    outputs(5335) <= not a or b;
    outputs(5336) <= b and not a;
    outputs(5337) <= a xor b;
    outputs(5338) <= a and not b;
    outputs(5339) <= not b;
    outputs(5340) <= not (a and b);
    outputs(5341) <= not b;
    outputs(5342) <= a and b;
    outputs(5343) <= a or b;
    outputs(5344) <= a and b;
    outputs(5345) <= not b or a;
    outputs(5346) <= a and b;
    outputs(5347) <= not b;
    outputs(5348) <= b;
    outputs(5349) <= not (a or b);
    outputs(5350) <= a;
    outputs(5351) <= not b;
    outputs(5352) <= not b;
    outputs(5353) <= a and not b;
    outputs(5354) <= not b;
    outputs(5355) <= not (a and b);
    outputs(5356) <= not a or b;
    outputs(5357) <= not a or b;
    outputs(5358) <= a xor b;
    outputs(5359) <= a xor b;
    outputs(5360) <= a and b;
    outputs(5361) <= not b or a;
    outputs(5362) <= not b;
    outputs(5363) <= a;
    outputs(5364) <= a;
    outputs(5365) <= a;
    outputs(5366) <= a xor b;
    outputs(5367) <= a;
    outputs(5368) <= not b;
    outputs(5369) <= not (a or b);
    outputs(5370) <= not a;
    outputs(5371) <= b;
    outputs(5372) <= not (a xor b);
    outputs(5373) <= a and not b;
    outputs(5374) <= b;
    outputs(5375) <= not a;
    outputs(5376) <= b and not a;
    outputs(5377) <= a and b;
    outputs(5378) <= not a;
    outputs(5379) <= a;
    outputs(5380) <= not b;
    outputs(5381) <= not b;
    outputs(5382) <= a and not b;
    outputs(5383) <= not a;
    outputs(5384) <= not a or b;
    outputs(5385) <= not (a and b);
    outputs(5386) <= a;
    outputs(5387) <= a and not b;
    outputs(5388) <= a;
    outputs(5389) <= a and not b;
    outputs(5390) <= b;
    outputs(5391) <= b;
    outputs(5392) <= a xor b;
    outputs(5393) <= a and b;
    outputs(5394) <= b;
    outputs(5395) <= a and b;
    outputs(5396) <= not (a and b);
    outputs(5397) <= a and not b;
    outputs(5398) <= a;
    outputs(5399) <= b;
    outputs(5400) <= b;
    outputs(5401) <= not b or a;
    outputs(5402) <= not (a or b);
    outputs(5403) <= a and b;
    outputs(5404) <= not (a xor b);
    outputs(5405) <= not (a or b);
    outputs(5406) <= not a;
    outputs(5407) <= a or b;
    outputs(5408) <= a and b;
    outputs(5409) <= not (a xor b);
    outputs(5410) <= a xor b;
    outputs(5411) <= not b;
    outputs(5412) <= not b;
    outputs(5413) <= not b or a;
    outputs(5414) <= a and b;
    outputs(5415) <= not a;
    outputs(5416) <= not b;
    outputs(5417) <= not (a or b);
    outputs(5418) <= not (a or b);
    outputs(5419) <= not b or a;
    outputs(5420) <= not a;
    outputs(5421) <= b;
    outputs(5422) <= not (a xor b);
    outputs(5423) <= a and b;
    outputs(5424) <= b;
    outputs(5425) <= not a or b;
    outputs(5426) <= b and not a;
    outputs(5427) <= a and b;
    outputs(5428) <= not b;
    outputs(5429) <= not b;
    outputs(5430) <= not (a and b);
    outputs(5431) <= b;
    outputs(5432) <= not (a and b);
    outputs(5433) <= not a;
    outputs(5434) <= not (a and b);
    outputs(5435) <= a and not b;
    outputs(5436) <= not (a or b);
    outputs(5437) <= a and b;
    outputs(5438) <= a;
    outputs(5439) <= b and not a;
    outputs(5440) <= not b;
    outputs(5441) <= a xor b;
    outputs(5442) <= not b;
    outputs(5443) <= a;
    outputs(5444) <= a xor b;
    outputs(5445) <= b;
    outputs(5446) <= b;
    outputs(5447) <= a or b;
    outputs(5448) <= not (a or b);
    outputs(5449) <= a xor b;
    outputs(5450) <= b;
    outputs(5451) <= b and not a;
    outputs(5452) <= not (a xor b);
    outputs(5453) <= a and b;
    outputs(5454) <= not b;
    outputs(5455) <= not a;
    outputs(5456) <= not a;
    outputs(5457) <= a;
    outputs(5458) <= not b or a;
    outputs(5459) <= a xor b;
    outputs(5460) <= not (a xor b);
    outputs(5461) <= b and not a;
    outputs(5462) <= b;
    outputs(5463) <= b;
    outputs(5464) <= a and b;
    outputs(5465) <= not b or a;
    outputs(5466) <= a or b;
    outputs(5467) <= a or b;
    outputs(5468) <= not b;
    outputs(5469) <= a and b;
    outputs(5470) <= a and b;
    outputs(5471) <= not b;
    outputs(5472) <= b and not a;
    outputs(5473) <= not a;
    outputs(5474) <= not a;
    outputs(5475) <= a;
    outputs(5476) <= not (a or b);
    outputs(5477) <= a xor b;
    outputs(5478) <= a and b;
    outputs(5479) <= not b;
    outputs(5480) <= not a;
    outputs(5481) <= a and not b;
    outputs(5482) <= b and not a;
    outputs(5483) <= not a;
    outputs(5484) <= not (a or b);
    outputs(5485) <= a and b;
    outputs(5486) <= not b or a;
    outputs(5487) <= not (a or b);
    outputs(5488) <= not b;
    outputs(5489) <= not (a or b);
    outputs(5490) <= not (a xor b);
    outputs(5491) <= not a;
    outputs(5492) <= not a or b;
    outputs(5493) <= a xor b;
    outputs(5494) <= not b or a;
    outputs(5495) <= a;
    outputs(5496) <= a and not b;
    outputs(5497) <= a and not b;
    outputs(5498) <= not b;
    outputs(5499) <= not a;
    outputs(5500) <= a xor b;
    outputs(5501) <= not (a and b);
    outputs(5502) <= a and b;
    outputs(5503) <= b;
    outputs(5504) <= a;
    outputs(5505) <= not b;
    outputs(5506) <= a;
    outputs(5507) <= a;
    outputs(5508) <= a and b;
    outputs(5509) <= not (a xor b);
    outputs(5510) <= a and not b;
    outputs(5511) <= not (a xor b);
    outputs(5512) <= a and b;
    outputs(5513) <= b;
    outputs(5514) <= b and not a;
    outputs(5515) <= a and not b;
    outputs(5516) <= not b or a;
    outputs(5517) <= not b;
    outputs(5518) <= not (a xor b);
    outputs(5519) <= not a;
    outputs(5520) <= b and not a;
    outputs(5521) <= not (a and b);
    outputs(5522) <= a and b;
    outputs(5523) <= not (a or b);
    outputs(5524) <= not b;
    outputs(5525) <= a;
    outputs(5526) <= a and not b;
    outputs(5527) <= not (a or b);
    outputs(5528) <= not b or a;
    outputs(5529) <= b and not a;
    outputs(5530) <= a and not b;
    outputs(5531) <= a;
    outputs(5532) <= a and not b;
    outputs(5533) <= not b or a;
    outputs(5534) <= b;
    outputs(5535) <= a xor b;
    outputs(5536) <= a and not b;
    outputs(5537) <= b and not a;
    outputs(5538) <= a xor b;
    outputs(5539) <= a;
    outputs(5540) <= not a;
    outputs(5541) <= b;
    outputs(5542) <= a;
    outputs(5543) <= a and not b;
    outputs(5544) <= not b;
    outputs(5545) <= b;
    outputs(5546) <= a and b;
    outputs(5547) <= a and not b;
    outputs(5548) <= a;
    outputs(5549) <= not b;
    outputs(5550) <= not b;
    outputs(5551) <= not (a xor b);
    outputs(5552) <= not (a xor b);
    outputs(5553) <= not (a xor b);
    outputs(5554) <= a and b;
    outputs(5555) <= not (a xor b);
    outputs(5556) <= a xor b;
    outputs(5557) <= not a;
    outputs(5558) <= a and not b;
    outputs(5559) <= not b;
    outputs(5560) <= b;
    outputs(5561) <= not (a or b);
    outputs(5562) <= a or b;
    outputs(5563) <= not a or b;
    outputs(5564) <= not (a and b);
    outputs(5565) <= not b;
    outputs(5566) <= b;
    outputs(5567) <= not (a xor b);
    outputs(5568) <= b;
    outputs(5569) <= b and not a;
    outputs(5570) <= not (a or b);
    outputs(5571) <= a xor b;
    outputs(5572) <= a;
    outputs(5573) <= a;
    outputs(5574) <= a;
    outputs(5575) <= not b;
    outputs(5576) <= a;
    outputs(5577) <= not (a and b);
    outputs(5578) <= not b;
    outputs(5579) <= a and b;
    outputs(5580) <= b;
    outputs(5581) <= not a;
    outputs(5582) <= a xor b;
    outputs(5583) <= not a;
    outputs(5584) <= not (a and b);
    outputs(5585) <= a and b;
    outputs(5586) <= a;
    outputs(5587) <= not (a xor b);
    outputs(5588) <= a and b;
    outputs(5589) <= not (a and b);
    outputs(5590) <= b and not a;
    outputs(5591) <= not a;
    outputs(5592) <= not (a or b);
    outputs(5593) <= a;
    outputs(5594) <= a or b;
    outputs(5595) <= not (a or b);
    outputs(5596) <= a and not b;
    outputs(5597) <= not (a or b);
    outputs(5598) <= a and b;
    outputs(5599) <= not (a xor b);
    outputs(5600) <= not a;
    outputs(5601) <= a and not b;
    outputs(5602) <= not a or b;
    outputs(5603) <= a and not b;
    outputs(5604) <= a and not b;
    outputs(5605) <= a and b;
    outputs(5606) <= b and not a;
    outputs(5607) <= a and b;
    outputs(5608) <= b and not a;
    outputs(5609) <= a xor b;
    outputs(5610) <= b;
    outputs(5611) <= a;
    outputs(5612) <= a and b;
    outputs(5613) <= not (a or b);
    outputs(5614) <= a and not b;
    outputs(5615) <= a xor b;
    outputs(5616) <= not (a xor b);
    outputs(5617) <= not b;
    outputs(5618) <= a or b;
    outputs(5619) <= not b;
    outputs(5620) <= not b;
    outputs(5621) <= not (a or b);
    outputs(5622) <= not a or b;
    outputs(5623) <= b and not a;
    outputs(5624) <= not (a xor b);
    outputs(5625) <= b;
    outputs(5626) <= b;
    outputs(5627) <= not (a or b);
    outputs(5628) <= a and b;
    outputs(5629) <= not a;
    outputs(5630) <= a and not b;
    outputs(5631) <= not (a and b);
    outputs(5632) <= b;
    outputs(5633) <= b;
    outputs(5634) <= b;
    outputs(5635) <= not (a and b);
    outputs(5636) <= b and not a;
    outputs(5637) <= a;
    outputs(5638) <= a;
    outputs(5639) <= a xor b;
    outputs(5640) <= a;
    outputs(5641) <= a xor b;
    outputs(5642) <= b;
    outputs(5643) <= not a;
    outputs(5644) <= not b;
    outputs(5645) <= not a;
    outputs(5646) <= b and not a;
    outputs(5647) <= a xor b;
    outputs(5648) <= a or b;
    outputs(5649) <= not a;
    outputs(5650) <= b and not a;
    outputs(5651) <= not b;
    outputs(5652) <= not (a or b);
    outputs(5653) <= not (a xor b);
    outputs(5654) <= b and not a;
    outputs(5655) <= a and not b;
    outputs(5656) <= b and not a;
    outputs(5657) <= not b;
    outputs(5658) <= a;
    outputs(5659) <= not a;
    outputs(5660) <= a;
    outputs(5661) <= not b;
    outputs(5662) <= a and not b;
    outputs(5663) <= a xor b;
    outputs(5664) <= a xor b;
    outputs(5665) <= b;
    outputs(5666) <= not a;
    outputs(5667) <= not (a xor b);
    outputs(5668) <= not a;
    outputs(5669) <= not a;
    outputs(5670) <= a;
    outputs(5671) <= not (a xor b);
    outputs(5672) <= b and not a;
    outputs(5673) <= b and not a;
    outputs(5674) <= not a;
    outputs(5675) <= not b;
    outputs(5676) <= a or b;
    outputs(5677) <= not b;
    outputs(5678) <= not a;
    outputs(5679) <= b and not a;
    outputs(5680) <= a xor b;
    outputs(5681) <= not b;
    outputs(5682) <= a;
    outputs(5683) <= b;
    outputs(5684) <= a xor b;
    outputs(5685) <= b and not a;
    outputs(5686) <= a;
    outputs(5687) <= not (a xor b);
    outputs(5688) <= a xor b;
    outputs(5689) <= not (a xor b);
    outputs(5690) <= a;
    outputs(5691) <= b;
    outputs(5692) <= not (a xor b);
    outputs(5693) <= not a or b;
    outputs(5694) <= a xor b;
    outputs(5695) <= not a;
    outputs(5696) <= a and not b;
    outputs(5697) <= b;
    outputs(5698) <= a;
    outputs(5699) <= not b;
    outputs(5700) <= not (a xor b);
    outputs(5701) <= b and not a;
    outputs(5702) <= not (a or b);
    outputs(5703) <= a xor b;
    outputs(5704) <= a xor b;
    outputs(5705) <= a xor b;
    outputs(5706) <= not (a xor b);
    outputs(5707) <= a xor b;
    outputs(5708) <= a xor b;
    outputs(5709) <= not a;
    outputs(5710) <= a xor b;
    outputs(5711) <= a and b;
    outputs(5712) <= a and not b;
    outputs(5713) <= a;
    outputs(5714) <= a xor b;
    outputs(5715) <= not b or a;
    outputs(5716) <= a xor b;
    outputs(5717) <= a xor b;
    outputs(5718) <= not b;
    outputs(5719) <= not b;
    outputs(5720) <= b and not a;
    outputs(5721) <= a;
    outputs(5722) <= b;
    outputs(5723) <= b;
    outputs(5724) <= not (a and b);
    outputs(5725) <= not (a and b);
    outputs(5726) <= a and not b;
    outputs(5727) <= a xor b;
    outputs(5728) <= a and b;
    outputs(5729) <= a xor b;
    outputs(5730) <= not a or b;
    outputs(5731) <= not a;
    outputs(5732) <= a and b;
    outputs(5733) <= not (a xor b);
    outputs(5734) <= b and not a;
    outputs(5735) <= b and not a;
    outputs(5736) <= a and not b;
    outputs(5737) <= not b;
    outputs(5738) <= a and b;
    outputs(5739) <= not (a xor b);
    outputs(5740) <= not (a xor b);
    outputs(5741) <= a and not b;
    outputs(5742) <= not a or b;
    outputs(5743) <= not (a xor b);
    outputs(5744) <= a and b;
    outputs(5745) <= not (a xor b);
    outputs(5746) <= not a;
    outputs(5747) <= not a;
    outputs(5748) <= not (a and b);
    outputs(5749) <= a and not b;
    outputs(5750) <= b;
    outputs(5751) <= a xor b;
    outputs(5752) <= a and b;
    outputs(5753) <= not (a xor b);
    outputs(5754) <= a or b;
    outputs(5755) <= not b;
    outputs(5756) <= not b;
    outputs(5757) <= a;
    outputs(5758) <= a and b;
    outputs(5759) <= not b;
    outputs(5760) <= b;
    outputs(5761) <= b and not a;
    outputs(5762) <= not b;
    outputs(5763) <= a xor b;
    outputs(5764) <= not a;
    outputs(5765) <= b;
    outputs(5766) <= a xor b;
    outputs(5767) <= not (a xor b);
    outputs(5768) <= not (a xor b);
    outputs(5769) <= not a;
    outputs(5770) <= not (a xor b);
    outputs(5771) <= not (a xor b);
    outputs(5772) <= not (a xor b);
    outputs(5773) <= a xor b;
    outputs(5774) <= b;
    outputs(5775) <= a;
    outputs(5776) <= not b;
    outputs(5777) <= not a or b;
    outputs(5778) <= a;
    outputs(5779) <= not (a xor b);
    outputs(5780) <= a and not b;
    outputs(5781) <= a xor b;
    outputs(5782) <= b and not a;
    outputs(5783) <= not (a or b);
    outputs(5784) <= a or b;
    outputs(5785) <= a and not b;
    outputs(5786) <= not a;
    outputs(5787) <= a and b;
    outputs(5788) <= a;
    outputs(5789) <= b and not a;
    outputs(5790) <= 1'b1;
    outputs(5791) <= not b;
    outputs(5792) <= b;
    outputs(5793) <= a and b;
    outputs(5794) <= a or b;
    outputs(5795) <= b and not a;
    outputs(5796) <= not (a and b);
    outputs(5797) <= b and not a;
    outputs(5798) <= a and not b;
    outputs(5799) <= not a;
    outputs(5800) <= a xor b;
    outputs(5801) <= not b;
    outputs(5802) <= not (a and b);
    outputs(5803) <= a;
    outputs(5804) <= b;
    outputs(5805) <= a and not b;
    outputs(5806) <= not (a xor b);
    outputs(5807) <= a xor b;
    outputs(5808) <= a;
    outputs(5809) <= b and not a;
    outputs(5810) <= b;
    outputs(5811) <= not (a xor b);
    outputs(5812) <= not a;
    outputs(5813) <= b;
    outputs(5814) <= not b;
    outputs(5815) <= b and not a;
    outputs(5816) <= not a or b;
    outputs(5817) <= a;
    outputs(5818) <= a;
    outputs(5819) <= a;
    outputs(5820) <= not (a or b);
    outputs(5821) <= a or b;
    outputs(5822) <= a xor b;
    outputs(5823) <= a;
    outputs(5824) <= a xor b;
    outputs(5825) <= b;
    outputs(5826) <= a and b;
    outputs(5827) <= not a;
    outputs(5828) <= a;
    outputs(5829) <= not a or b;
    outputs(5830) <= a xor b;
    outputs(5831) <= a and not b;
    outputs(5832) <= b;
    outputs(5833) <= b;
    outputs(5834) <= not b;
    outputs(5835) <= b;
    outputs(5836) <= not (a xor b);
    outputs(5837) <= not (a and b);
    outputs(5838) <= not (a and b);
    outputs(5839) <= a;
    outputs(5840) <= b and not a;
    outputs(5841) <= not b;
    outputs(5842) <= a xor b;
    outputs(5843) <= not (a xor b);
    outputs(5844) <= a and b;
    outputs(5845) <= a and not b;
    outputs(5846) <= not b;
    outputs(5847) <= b;
    outputs(5848) <= b and not a;
    outputs(5849) <= a and not b;
    outputs(5850) <= b;
    outputs(5851) <= a xor b;
    outputs(5852) <= a xor b;
    outputs(5853) <= not b or a;
    outputs(5854) <= a and b;
    outputs(5855) <= b;
    outputs(5856) <= not a;
    outputs(5857) <= a;
    outputs(5858) <= a and b;
    outputs(5859) <= not a;
    outputs(5860) <= not (a or b);
    outputs(5861) <= a xor b;
    outputs(5862) <= not (a xor b);
    outputs(5863) <= b and not a;
    outputs(5864) <= not b;
    outputs(5865) <= not (a xor b);
    outputs(5866) <= a;
    outputs(5867) <= a and not b;
    outputs(5868) <= a and not b;
    outputs(5869) <= not (a xor b);
    outputs(5870) <= not (a xor b);
    outputs(5871) <= b and not a;
    outputs(5872) <= b;
    outputs(5873) <= a and b;
    outputs(5874) <= not (a or b);
    outputs(5875) <= not (a and b);
    outputs(5876) <= a and b;
    outputs(5877) <= a xor b;
    outputs(5878) <= a;
    outputs(5879) <= not (a xor b);
    outputs(5880) <= b and not a;
    outputs(5881) <= a and b;
    outputs(5882) <= not (a or b);
    outputs(5883) <= a and not b;
    outputs(5884) <= a;
    outputs(5885) <= not (a or b);
    outputs(5886) <= not (a or b);
    outputs(5887) <= a;
    outputs(5888) <= not (a and b);
    outputs(5889) <= a or b;
    outputs(5890) <= a;
    outputs(5891) <= a and b;
    outputs(5892) <= a and not b;
    outputs(5893) <= not a;
    outputs(5894) <= b;
    outputs(5895) <= a xor b;
    outputs(5896) <= not a;
    outputs(5897) <= a and b;
    outputs(5898) <= a or b;
    outputs(5899) <= a;
    outputs(5900) <= not (a or b);
    outputs(5901) <= a or b;
    outputs(5902) <= a;
    outputs(5903) <= not (a and b);
    outputs(5904) <= a and not b;
    outputs(5905) <= a;
    outputs(5906) <= b;
    outputs(5907) <= not (a xor b);
    outputs(5908) <= a xor b;
    outputs(5909) <= not b;
    outputs(5910) <= not a or b;
    outputs(5911) <= a and b;
    outputs(5912) <= not (a or b);
    outputs(5913) <= not b;
    outputs(5914) <= b;
    outputs(5915) <= b and not a;
    outputs(5916) <= b;
    outputs(5917) <= not b or a;
    outputs(5918) <= a;
    outputs(5919) <= not b;
    outputs(5920) <= not b or a;
    outputs(5921) <= not (a xor b);
    outputs(5922) <= not (a or b);
    outputs(5923) <= b;
    outputs(5924) <= not (a or b);
    outputs(5925) <= a;
    outputs(5926) <= not (a or b);
    outputs(5927) <= b;
    outputs(5928) <= a xor b;
    outputs(5929) <= not (a and b);
    outputs(5930) <= a and not b;
    outputs(5931) <= a and not b;
    outputs(5932) <= a;
    outputs(5933) <= a and not b;
    outputs(5934) <= a and b;
    outputs(5935) <= not (a xor b);
    outputs(5936) <= a xor b;
    outputs(5937) <= b;
    outputs(5938) <= not a;
    outputs(5939) <= b and not a;
    outputs(5940) <= a and b;
    outputs(5941) <= not (a xor b);
    outputs(5942) <= not (a xor b);
    outputs(5943) <= b;
    outputs(5944) <= a;
    outputs(5945) <= not a;
    outputs(5946) <= a or b;
    outputs(5947) <= not a;
    outputs(5948) <= not b;
    outputs(5949) <= a;
    outputs(5950) <= b;
    outputs(5951) <= a and b;
    outputs(5952) <= a;
    outputs(5953) <= b and not a;
    outputs(5954) <= not (a xor b);
    outputs(5955) <= not (a xor b);
    outputs(5956) <= a or b;
    outputs(5957) <= a xor b;
    outputs(5958) <= not b;
    outputs(5959) <= a or b;
    outputs(5960) <= not a;
    outputs(5961) <= b;
    outputs(5962) <= a and not b;
    outputs(5963) <= not b;
    outputs(5964) <= a xor b;
    outputs(5965) <= a xor b;
    outputs(5966) <= b and not a;
    outputs(5967) <= a;
    outputs(5968) <= a and b;
    outputs(5969) <= b;
    outputs(5970) <= not (a or b);
    outputs(5971) <= b;
    outputs(5972) <= not a;
    outputs(5973) <= not (a xor b);
    outputs(5974) <= not (a xor b);
    outputs(5975) <= a xor b;
    outputs(5976) <= a and b;
    outputs(5977) <= not a;
    outputs(5978) <= a and b;
    outputs(5979) <= not (a or b);
    outputs(5980) <= not (a xor b);
    outputs(5981) <= a and b;
    outputs(5982) <= a and not b;
    outputs(5983) <= a;
    outputs(5984) <= not b;
    outputs(5985) <= not a or b;
    outputs(5986) <= not a;
    outputs(5987) <= b;
    outputs(5988) <= not b;
    outputs(5989) <= not b;
    outputs(5990) <= a xor b;
    outputs(5991) <= a;
    outputs(5992) <= a xor b;
    outputs(5993) <= a;
    outputs(5994) <= not b;
    outputs(5995) <= not (a xor b);
    outputs(5996) <= not b or a;
    outputs(5997) <= a;
    outputs(5998) <= a and not b;
    outputs(5999) <= a xor b;
    outputs(6000) <= not a or b;
    outputs(6001) <= not (a or b);
    outputs(6002) <= a xor b;
    outputs(6003) <= not b;
    outputs(6004) <= b;
    outputs(6005) <= not (a or b);
    outputs(6006) <= a;
    outputs(6007) <= not b;
    outputs(6008) <= not b;
    outputs(6009) <= b;
    outputs(6010) <= not a;
    outputs(6011) <= a and not b;
    outputs(6012) <= b and not a;
    outputs(6013) <= a;
    outputs(6014) <= a xor b;
    outputs(6015) <= not a;
    outputs(6016) <= b and not a;
    outputs(6017) <= a and b;
    outputs(6018) <= b;
    outputs(6019) <= a;
    outputs(6020) <= a xor b;
    outputs(6021) <= not (a xor b);
    outputs(6022) <= a and b;
    outputs(6023) <= b and not a;
    outputs(6024) <= a;
    outputs(6025) <= b and not a;
    outputs(6026) <= not a;
    outputs(6027) <= b;
    outputs(6028) <= not b;
    outputs(6029) <= not (a xor b);
    outputs(6030) <= not b;
    outputs(6031) <= a xor b;
    outputs(6032) <= not (a or b);
    outputs(6033) <= not (a or b);
    outputs(6034) <= not b or a;
    outputs(6035) <= a xor b;
    outputs(6036) <= not (a xor b);
    outputs(6037) <= not (a xor b);
    outputs(6038) <= not (a and b);
    outputs(6039) <= b;
    outputs(6040) <= not (a and b);
    outputs(6041) <= not a;
    outputs(6042) <= b and not a;
    outputs(6043) <= not a;
    outputs(6044) <= not (a or b);
    outputs(6045) <= not (a xor b);
    outputs(6046) <= b and not a;
    outputs(6047) <= not b;
    outputs(6048) <= not (a xor b);
    outputs(6049) <= b and not a;
    outputs(6050) <= a and b;
    outputs(6051) <= not (a xor b);
    outputs(6052) <= b;
    outputs(6053) <= not a or b;
    outputs(6054) <= not (a xor b);
    outputs(6055) <= not b;
    outputs(6056) <= not (a or b);
    outputs(6057) <= a xor b;
    outputs(6058) <= not b;
    outputs(6059) <= a xor b;
    outputs(6060) <= a and b;
    outputs(6061) <= a and not b;
    outputs(6062) <= a;
    outputs(6063) <= a xor b;
    outputs(6064) <= not a;
    outputs(6065) <= not (a xor b);
    outputs(6066) <= not b;
    outputs(6067) <= a or b;
    outputs(6068) <= a xor b;
    outputs(6069) <= b;
    outputs(6070) <= a;
    outputs(6071) <= a and b;
    outputs(6072) <= b;
    outputs(6073) <= a;
    outputs(6074) <= not b;
    outputs(6075) <= not (a or b);
    outputs(6076) <= a xor b;
    outputs(6077) <= a;
    outputs(6078) <= not a;
    outputs(6079) <= not a;
    outputs(6080) <= not b or a;
    outputs(6081) <= a;
    outputs(6082) <= not (a or b);
    outputs(6083) <= not b;
    outputs(6084) <= a xor b;
    outputs(6085) <= a;
    outputs(6086) <= a;
    outputs(6087) <= not b;
    outputs(6088) <= not b;
    outputs(6089) <= not b;
    outputs(6090) <= not a;
    outputs(6091) <= b;
    outputs(6092) <= b;
    outputs(6093) <= not (a or b);
    outputs(6094) <= not (a and b);
    outputs(6095) <= a and not b;
    outputs(6096) <= not b;
    outputs(6097) <= a and b;
    outputs(6098) <= not b;
    outputs(6099) <= not b;
    outputs(6100) <= not (a xor b);
    outputs(6101) <= not a;
    outputs(6102) <= not (a or b);
    outputs(6103) <= not (a xor b);
    outputs(6104) <= b;
    outputs(6105) <= not a;
    outputs(6106) <= not (a and b);
    outputs(6107) <= not b;
    outputs(6108) <= a and not b;
    outputs(6109) <= b;
    outputs(6110) <= a or b;
    outputs(6111) <= not a;
    outputs(6112) <= not (a xor b);
    outputs(6113) <= a xor b;
    outputs(6114) <= a xor b;
    outputs(6115) <= b;
    outputs(6116) <= a;
    outputs(6117) <= b and not a;
    outputs(6118) <= a;
    outputs(6119) <= a xor b;
    outputs(6120) <= not b;
    outputs(6121) <= not b;
    outputs(6122) <= not (a or b);
    outputs(6123) <= not a;
    outputs(6124) <= a xor b;
    outputs(6125) <= b and not a;
    outputs(6126) <= a;
    outputs(6127) <= a xor b;
    outputs(6128) <= a xor b;
    outputs(6129) <= not (a xor b);
    outputs(6130) <= not (a or b);
    outputs(6131) <= b and not a;
    outputs(6132) <= not b;
    outputs(6133) <= not b or a;
    outputs(6134) <= a;
    outputs(6135) <= a;
    outputs(6136) <= a;
    outputs(6137) <= a;
    outputs(6138) <= b;
    outputs(6139) <= not (a xor b);
    outputs(6140) <= not a or b;
    outputs(6141) <= b;
    outputs(6142) <= b;
    outputs(6143) <= not b;
    outputs(6144) <= not a;
    outputs(6145) <= a and b;
    outputs(6146) <= a;
    outputs(6147) <= not (a xor b);
    outputs(6148) <= a xor b;
    outputs(6149) <= a xor b;
    outputs(6150) <= not (a xor b);
    outputs(6151) <= not b or a;
    outputs(6152) <= not (a xor b);
    outputs(6153) <= a;
    outputs(6154) <= b;
    outputs(6155) <= not (a xor b);
    outputs(6156) <= not b or a;
    outputs(6157) <= not b or a;
    outputs(6158) <= b and not a;
    outputs(6159) <= b;
    outputs(6160) <= not a;
    outputs(6161) <= not b or a;
    outputs(6162) <= a and b;
    outputs(6163) <= not b;
    outputs(6164) <= a;
    outputs(6165) <= not a or b;
    outputs(6166) <= not (a xor b);
    outputs(6167) <= b;
    outputs(6168) <= b and not a;
    outputs(6169) <= a and not b;
    outputs(6170) <= a;
    outputs(6171) <= a xor b;
    outputs(6172) <= a or b;
    outputs(6173) <= a;
    outputs(6174) <= not a;
    outputs(6175) <= not b;
    outputs(6176) <= not (a xor b);
    outputs(6177) <= a xor b;
    outputs(6178) <= b;
    outputs(6179) <= b;
    outputs(6180) <= not (a xor b);
    outputs(6181) <= not (a or b);
    outputs(6182) <= not b;
    outputs(6183) <= b and not a;
    outputs(6184) <= a xor b;
    outputs(6185) <= b;
    outputs(6186) <= b and not a;
    outputs(6187) <= a;
    outputs(6188) <= not (a xor b);
    outputs(6189) <= a;
    outputs(6190) <= not (a xor b);
    outputs(6191) <= not (a xor b);
    outputs(6192) <= a;
    outputs(6193) <= not b;
    outputs(6194) <= a xor b;
    outputs(6195) <= not b;
    outputs(6196) <= not (a xor b);
    outputs(6197) <= not a or b;
    outputs(6198) <= b and not a;
    outputs(6199) <= not (a and b);
    outputs(6200) <= not (a and b);
    outputs(6201) <= a and not b;
    outputs(6202) <= not (a or b);
    outputs(6203) <= a or b;
    outputs(6204) <= not b or a;
    outputs(6205) <= a xor b;
    outputs(6206) <= not a;
    outputs(6207) <= a;
    outputs(6208) <= not b;
    outputs(6209) <= not (a or b);
    outputs(6210) <= a or b;
    outputs(6211) <= not (a and b);
    outputs(6212) <= not (a or b);
    outputs(6213) <= a;
    outputs(6214) <= a;
    outputs(6215) <= a or b;
    outputs(6216) <= not (a xor b);
    outputs(6217) <= b;
    outputs(6218) <= not (a or b);
    outputs(6219) <= a;
    outputs(6220) <= not b or a;
    outputs(6221) <= not (a xor b);
    outputs(6222) <= not a;
    outputs(6223) <= not b;
    outputs(6224) <= not b or a;
    outputs(6225) <= a;
    outputs(6226) <= a xor b;
    outputs(6227) <= a xor b;
    outputs(6228) <= a;
    outputs(6229) <= b;
    outputs(6230) <= a xor b;
    outputs(6231) <= not a;
    outputs(6232) <= a xor b;
    outputs(6233) <= not a;
    outputs(6234) <= not (a xor b);
    outputs(6235) <= not a;
    outputs(6236) <= not b;
    outputs(6237) <= not b;
    outputs(6238) <= b;
    outputs(6239) <= a;
    outputs(6240) <= a;
    outputs(6241) <= a and not b;
    outputs(6242) <= not (a xor b);
    outputs(6243) <= a xor b;
    outputs(6244) <= a;
    outputs(6245) <= a xor b;
    outputs(6246) <= a xor b;
    outputs(6247) <= not (a xor b);
    outputs(6248) <= not a or b;
    outputs(6249) <= b;
    outputs(6250) <= not b;
    outputs(6251) <= not (a or b);
    outputs(6252) <= not (a xor b);
    outputs(6253) <= a and not b;
    outputs(6254) <= b;
    outputs(6255) <= a xor b;
    outputs(6256) <= not (a xor b);
    outputs(6257) <= not a;
    outputs(6258) <= not (a xor b);
    outputs(6259) <= a and not b;
    outputs(6260) <= not a;
    outputs(6261) <= not a;
    outputs(6262) <= a;
    outputs(6263) <= a xor b;
    outputs(6264) <= not b;
    outputs(6265) <= not b;
    outputs(6266) <= a xor b;
    outputs(6267) <= b and not a;
    outputs(6268) <= a and b;
    outputs(6269) <= b;
    outputs(6270) <= not a or b;
    outputs(6271) <= a;
    outputs(6272) <= a;
    outputs(6273) <= not a or b;
    outputs(6274) <= b;
    outputs(6275) <= not (a or b);
    outputs(6276) <= a xor b;
    outputs(6277) <= a;
    outputs(6278) <= not a;
    outputs(6279) <= b and not a;
    outputs(6280) <= not (a and b);
    outputs(6281) <= not b or a;
    outputs(6282) <= not (a xor b);
    outputs(6283) <= not b;
    outputs(6284) <= not (a xor b);
    outputs(6285) <= not (a xor b);
    outputs(6286) <= not (a and b);
    outputs(6287) <= not (a xor b);
    outputs(6288) <= not a or b;
    outputs(6289) <= b;
    outputs(6290) <= not b;
    outputs(6291) <= a and b;
    outputs(6292) <= not b;
    outputs(6293) <= a xor b;
    outputs(6294) <= a xor b;
    outputs(6295) <= a and b;
    outputs(6296) <= not (a xor b);
    outputs(6297) <= a and b;
    outputs(6298) <= not b;
    outputs(6299) <= a xor b;
    outputs(6300) <= b;
    outputs(6301) <= not a;
    outputs(6302) <= b;
    outputs(6303) <= a or b;
    outputs(6304) <= not (a xor b);
    outputs(6305) <= not (a xor b);
    outputs(6306) <= b;
    outputs(6307) <= a xor b;
    outputs(6308) <= b;
    outputs(6309) <= not (a and b);
    outputs(6310) <= a xor b;
    outputs(6311) <= not b;
    outputs(6312) <= not (a xor b);
    outputs(6313) <= a xor b;
    outputs(6314) <= b;
    outputs(6315) <= not (a xor b);
    outputs(6316) <= not (a xor b);
    outputs(6317) <= not (a xor b);
    outputs(6318) <= a;
    outputs(6319) <= not a or b;
    outputs(6320) <= b;
    outputs(6321) <= not b;
    outputs(6322) <= a and b;
    outputs(6323) <= b and not a;
    outputs(6324) <= not (a xor b);
    outputs(6325) <= not (a xor b);
    outputs(6326) <= a;
    outputs(6327) <= not (a xor b);
    outputs(6328) <= b;
    outputs(6329) <= not b;
    outputs(6330) <= a xor b;
    outputs(6331) <= a and not b;
    outputs(6332) <= a and b;
    outputs(6333) <= b;
    outputs(6334) <= b;
    outputs(6335) <= a;
    outputs(6336) <= not b;
    outputs(6337) <= a xor b;
    outputs(6338) <= not b;
    outputs(6339) <= a xor b;
    outputs(6340) <= not (a xor b);
    outputs(6341) <= not a or b;
    outputs(6342) <= not a;
    outputs(6343) <= not (a and b);
    outputs(6344) <= b;
    outputs(6345) <= not (a or b);
    outputs(6346) <= not a;
    outputs(6347) <= a;
    outputs(6348) <= a and not b;
    outputs(6349) <= b;
    outputs(6350) <= a xor b;
    outputs(6351) <= a xor b;
    outputs(6352) <= b;
    outputs(6353) <= a and not b;
    outputs(6354) <= not b;
    outputs(6355) <= not (a and b);
    outputs(6356) <= not (a xor b);
    outputs(6357) <= a;
    outputs(6358) <= not b;
    outputs(6359) <= not (a and b);
    outputs(6360) <= a and b;
    outputs(6361) <= not (a or b);
    outputs(6362) <= not (a xor b);
    outputs(6363) <= a and b;
    outputs(6364) <= not b;
    outputs(6365) <= a xor b;
    outputs(6366) <= not (a xor b);
    outputs(6367) <= b;
    outputs(6368) <= a and not b;
    outputs(6369) <= not (a xor b);
    outputs(6370) <= not (a xor b);
    outputs(6371) <= not (a xor b);
    outputs(6372) <= a;
    outputs(6373) <= not b or a;
    outputs(6374) <= b;
    outputs(6375) <= not (a xor b);
    outputs(6376) <= a xor b;
    outputs(6377) <= a;
    outputs(6378) <= not (a xor b);
    outputs(6379) <= not (a xor b);
    outputs(6380) <= a;
    outputs(6381) <= b;
    outputs(6382) <= a;
    outputs(6383) <= b;
    outputs(6384) <= a or b;
    outputs(6385) <= a and b;
    outputs(6386) <= not (a and b);
    outputs(6387) <= a or b;
    outputs(6388) <= not b;
    outputs(6389) <= not b or a;
    outputs(6390) <= a xor b;
    outputs(6391) <= not a;
    outputs(6392) <= not a or b;
    outputs(6393) <= not (a or b);
    outputs(6394) <= not (a xor b);
    outputs(6395) <= not (a xor b);
    outputs(6396) <= not (a xor b);
    outputs(6397) <= a;
    outputs(6398) <= b;
    outputs(6399) <= not (a xor b);
    outputs(6400) <= a xor b;
    outputs(6401) <= not b;
    outputs(6402) <= a xor b;
    outputs(6403) <= a xor b;
    outputs(6404) <= a xor b;
    outputs(6405) <= b and not a;
    outputs(6406) <= a;
    outputs(6407) <= a xor b;
    outputs(6408) <= a xor b;
    outputs(6409) <= a and b;
    outputs(6410) <= b;
    outputs(6411) <= a xor b;
    outputs(6412) <= b;
    outputs(6413) <= b;
    outputs(6414) <= not b or a;
    outputs(6415) <= not b or a;
    outputs(6416) <= a or b;
    outputs(6417) <= a and not b;
    outputs(6418) <= not b or a;
    outputs(6419) <= not (a or b);
    outputs(6420) <= not b;
    outputs(6421) <= a;
    outputs(6422) <= not b or a;
    outputs(6423) <= a or b;
    outputs(6424) <= a;
    outputs(6425) <= not (a or b);
    outputs(6426) <= a and not b;
    outputs(6427) <= b;
    outputs(6428) <= not (a xor b);
    outputs(6429) <= not a;
    outputs(6430) <= not a or b;
    outputs(6431) <= not (a and b);
    outputs(6432) <= a and b;
    outputs(6433) <= not b;
    outputs(6434) <= b and not a;
    outputs(6435) <= a and not b;
    outputs(6436) <= a;
    outputs(6437) <= a xor b;
    outputs(6438) <= not (a and b);
    outputs(6439) <= not (a and b);
    outputs(6440) <= b;
    outputs(6441) <= b;
    outputs(6442) <= a;
    outputs(6443) <= not b;
    outputs(6444) <= not (a xor b);
    outputs(6445) <= a;
    outputs(6446) <= not a;
    outputs(6447) <= not (a xor b);
    outputs(6448) <= b and not a;
    outputs(6449) <= not a;
    outputs(6450) <= not b;
    outputs(6451) <= not (a or b);
    outputs(6452) <= a;
    outputs(6453) <= not (a xor b);
    outputs(6454) <= a xor b;
    outputs(6455) <= not a;
    outputs(6456) <= b;
    outputs(6457) <= not a;
    outputs(6458) <= not (a or b);
    outputs(6459) <= not (a or b);
    outputs(6460) <= not b;
    outputs(6461) <= a;
    outputs(6462) <= not (a or b);
    outputs(6463) <= not (a xor b);
    outputs(6464) <= not (a and b);
    outputs(6465) <= a;
    outputs(6466) <= not (a xor b);
    outputs(6467) <= b;
    outputs(6468) <= a and b;
    outputs(6469) <= not a;
    outputs(6470) <= b;
    outputs(6471) <= not (a xor b);
    outputs(6472) <= a;
    outputs(6473) <= not (a xor b);
    outputs(6474) <= not a;
    outputs(6475) <= not a;
    outputs(6476) <= a and not b;
    outputs(6477) <= not b;
    outputs(6478) <= not b;
    outputs(6479) <= not (a xor b);
    outputs(6480) <= not b;
    outputs(6481) <= a and b;
    outputs(6482) <= not (a xor b);
    outputs(6483) <= not a;
    outputs(6484) <= b;
    outputs(6485) <= not b;
    outputs(6486) <= a;
    outputs(6487) <= a and b;
    outputs(6488) <= a xor b;
    outputs(6489) <= b;
    outputs(6490) <= not a;
    outputs(6491) <= a xor b;
    outputs(6492) <= not a;
    outputs(6493) <= a;
    outputs(6494) <= a and not b;
    outputs(6495) <= not b or a;
    outputs(6496) <= b and not a;
    outputs(6497) <= not a or b;
    outputs(6498) <= not (a xor b);
    outputs(6499) <= a;
    outputs(6500) <= not (a xor b);
    outputs(6501) <= not a or b;
    outputs(6502) <= not (a or b);
    outputs(6503) <= a and b;
    outputs(6504) <= b;
    outputs(6505) <= not a;
    outputs(6506) <= a;
    outputs(6507) <= not b;
    outputs(6508) <= not a;
    outputs(6509) <= not b or a;
    outputs(6510) <= not b or a;
    outputs(6511) <= a and b;
    outputs(6512) <= not a;
    outputs(6513) <= a xor b;
    outputs(6514) <= not a or b;
    outputs(6515) <= a;
    outputs(6516) <= b and not a;
    outputs(6517) <= a;
    outputs(6518) <= not b;
    outputs(6519) <= not (a or b);
    outputs(6520) <= b;
    outputs(6521) <= a xor b;
    outputs(6522) <= not a;
    outputs(6523) <= not b;
    outputs(6524) <= not (a and b);
    outputs(6525) <= a or b;
    outputs(6526) <= b;
    outputs(6527) <= a xor b;
    outputs(6528) <= b;
    outputs(6529) <= not (a or b);
    outputs(6530) <= a or b;
    outputs(6531) <= a and b;
    outputs(6532) <= a and b;
    outputs(6533) <= a;
    outputs(6534) <= not (a or b);
    outputs(6535) <= a xor b;
    outputs(6536) <= a or b;
    outputs(6537) <= b;
    outputs(6538) <= b and not a;
    outputs(6539) <= not (a or b);
    outputs(6540) <= a xor b;
    outputs(6541) <= a;
    outputs(6542) <= a or b;
    outputs(6543) <= a and b;
    outputs(6544) <= not a;
    outputs(6545) <= a;
    outputs(6546) <= b and not a;
    outputs(6547) <= a;
    outputs(6548) <= not (a and b);
    outputs(6549) <= not (a xor b);
    outputs(6550) <= a;
    outputs(6551) <= not b or a;
    outputs(6552) <= a;
    outputs(6553) <= not a or b;
    outputs(6554) <= not a;
    outputs(6555) <= b;
    outputs(6556) <= not a;
    outputs(6557) <= not (a xor b);
    outputs(6558) <= a or b;
    outputs(6559) <= a and b;
    outputs(6560) <= b;
    outputs(6561) <= b;
    outputs(6562) <= not b;
    outputs(6563) <= not a;
    outputs(6564) <= not a or b;
    outputs(6565) <= b and not a;
    outputs(6566) <= a or b;
    outputs(6567) <= not b;
    outputs(6568) <= a;
    outputs(6569) <= b;
    outputs(6570) <= a and b;
    outputs(6571) <= not (a xor b);
    outputs(6572) <= a and b;
    outputs(6573) <= not (a or b);
    outputs(6574) <= not a or b;
    outputs(6575) <= not (a xor b);
    outputs(6576) <= not a;
    outputs(6577) <= not (a xor b);
    outputs(6578) <= a;
    outputs(6579) <= not b or a;
    outputs(6580) <= a;
    outputs(6581) <= not (a xor b);
    outputs(6582) <= not (a xor b);
    outputs(6583) <= a xor b;
    outputs(6584) <= not a;
    outputs(6585) <= a xor b;
    outputs(6586) <= not (a and b);
    outputs(6587) <= b;
    outputs(6588) <= b;
    outputs(6589) <= a;
    outputs(6590) <= b;
    outputs(6591) <= not b;
    outputs(6592) <= not b;
    outputs(6593) <= a xor b;
    outputs(6594) <= a;
    outputs(6595) <= not b;
    outputs(6596) <= not (a or b);
    outputs(6597) <= a;
    outputs(6598) <= b;
    outputs(6599) <= a xor b;
    outputs(6600) <= a xor b;
    outputs(6601) <= not (a xor b);
    outputs(6602) <= a and not b;
    outputs(6603) <= a and b;
    outputs(6604) <= not b;
    outputs(6605) <= a and b;
    outputs(6606) <= not a or b;
    outputs(6607) <= b;
    outputs(6608) <= a and not b;
    outputs(6609) <= not b;
    outputs(6610) <= not b;
    outputs(6611) <= not a;
    outputs(6612) <= b and not a;
    outputs(6613) <= b and not a;
    outputs(6614) <= a or b;
    outputs(6615) <= b and not a;
    outputs(6616) <= a and not b;
    outputs(6617) <= not a;
    outputs(6618) <= a;
    outputs(6619) <= not (a and b);
    outputs(6620) <= not (a or b);
    outputs(6621) <= not (a or b);
    outputs(6622) <= not (a and b);
    outputs(6623) <= not a or b;
    outputs(6624) <= not a or b;
    outputs(6625) <= a and b;
    outputs(6626) <= a and not b;
    outputs(6627) <= b and not a;
    outputs(6628) <= a xor b;
    outputs(6629) <= a and b;
    outputs(6630) <= not a;
    outputs(6631) <= a and b;
    outputs(6632) <= b;
    outputs(6633) <= a xor b;
    outputs(6634) <= b;
    outputs(6635) <= a and not b;
    outputs(6636) <= a xor b;
    outputs(6637) <= not b;
    outputs(6638) <= a or b;
    outputs(6639) <= b;
    outputs(6640) <= a and not b;
    outputs(6641) <= not (a and b);
    outputs(6642) <= a and not b;
    outputs(6643) <= not (a xor b);
    outputs(6644) <= b and not a;
    outputs(6645) <= a xor b;
    outputs(6646) <= not (a xor b);
    outputs(6647) <= a xor b;
    outputs(6648) <= not (a xor b);
    outputs(6649) <= not a;
    outputs(6650) <= b and not a;
    outputs(6651) <= not b or a;
    outputs(6652) <= a xor b;
    outputs(6653) <= b;
    outputs(6654) <= not a;
    outputs(6655) <= b;
    outputs(6656) <= not (a or b);
    outputs(6657) <= not (a xor b);
    outputs(6658) <= not (a or b);
    outputs(6659) <= not b;
    outputs(6660) <= not b;
    outputs(6661) <= a and not b;
    outputs(6662) <= not b;
    outputs(6663) <= a xor b;
    outputs(6664) <= b;
    outputs(6665) <= a xor b;
    outputs(6666) <= a and not b;
    outputs(6667) <= a and b;
    outputs(6668) <= not b or a;
    outputs(6669) <= not b;
    outputs(6670) <= b and not a;
    outputs(6671) <= a xor b;
    outputs(6672) <= not a or b;
    outputs(6673) <= not b;
    outputs(6674) <= a;
    outputs(6675) <= a and not b;
    outputs(6676) <= a xor b;
    outputs(6677) <= not b;
    outputs(6678) <= a and not b;
    outputs(6679) <= a xor b;
    outputs(6680) <= not a;
    outputs(6681) <= b and not a;
    outputs(6682) <= not (a or b);
    outputs(6683) <= a;
    outputs(6684) <= b;
    outputs(6685) <= a xor b;
    outputs(6686) <= not (a xor b);
    outputs(6687) <= not (a or b);
    outputs(6688) <= a xor b;
    outputs(6689) <= not (a xor b);
    outputs(6690) <= not (a xor b);
    outputs(6691) <= b;
    outputs(6692) <= a;
    outputs(6693) <= not a;
    outputs(6694) <= a;
    outputs(6695) <= a;
    outputs(6696) <= not a;
    outputs(6697) <= b;
    outputs(6698) <= b and not a;
    outputs(6699) <= a xor b;
    outputs(6700) <= not b;
    outputs(6701) <= a and not b;
    outputs(6702) <= a and b;
    outputs(6703) <= a and b;
    outputs(6704) <= not a or b;
    outputs(6705) <= a xor b;
    outputs(6706) <= not (a xor b);
    outputs(6707) <= not a or b;
    outputs(6708) <= a;
    outputs(6709) <= not (a xor b);
    outputs(6710) <= not b or a;
    outputs(6711) <= not b;
    outputs(6712) <= not (a or b);
    outputs(6713) <= not b;
    outputs(6714) <= a xor b;
    outputs(6715) <= a or b;
    outputs(6716) <= not (a xor b);
    outputs(6717) <= a and b;
    outputs(6718) <= a and not b;
    outputs(6719) <= not (a xor b);
    outputs(6720) <= a;
    outputs(6721) <= a;
    outputs(6722) <= not (a or b);
    outputs(6723) <= b and not a;
    outputs(6724) <= not b;
    outputs(6725) <= a;
    outputs(6726) <= a and not b;
    outputs(6727) <= not (a or b);
    outputs(6728) <= not (a xor b);
    outputs(6729) <= not (a or b);
    outputs(6730) <= not b;
    outputs(6731) <= not a;
    outputs(6732) <= not a;
    outputs(6733) <= a and b;
    outputs(6734) <= a xor b;
    outputs(6735) <= b;
    outputs(6736) <= a xor b;
    outputs(6737) <= not a;
    outputs(6738) <= not a;
    outputs(6739) <= a xor b;
    outputs(6740) <= not (a xor b);
    outputs(6741) <= not (a and b);
    outputs(6742) <= b;
    outputs(6743) <= not b or a;
    outputs(6744) <= a xor b;
    outputs(6745) <= a;
    outputs(6746) <= not (a xor b);
    outputs(6747) <= not a;
    outputs(6748) <= a and not b;
    outputs(6749) <= not b;
    outputs(6750) <= not (a or b);
    outputs(6751) <= b;
    outputs(6752) <= b;
    outputs(6753) <= not b;
    outputs(6754) <= a and not b;
    outputs(6755) <= b and not a;
    outputs(6756) <= a and not b;
    outputs(6757) <= a xor b;
    outputs(6758) <= not (a or b);
    outputs(6759) <= not (a xor b);
    outputs(6760) <= a and b;
    outputs(6761) <= not (a xor b);
    outputs(6762) <= a or b;
    outputs(6763) <= not (a or b);
    outputs(6764) <= not b;
    outputs(6765) <= b and not a;
    outputs(6766) <= a;
    outputs(6767) <= a xor b;
    outputs(6768) <= a and not b;
    outputs(6769) <= b;
    outputs(6770) <= a;
    outputs(6771) <= not (a xor b);
    outputs(6772) <= b;
    outputs(6773) <= a xor b;
    outputs(6774) <= a;
    outputs(6775) <= a;
    outputs(6776) <= b and not a;
    outputs(6777) <= a or b;
    outputs(6778) <= a xor b;
    outputs(6779) <= not a;
    outputs(6780) <= b;
    outputs(6781) <= a xor b;
    outputs(6782) <= not a;
    outputs(6783) <= not (a xor b);
    outputs(6784) <= a xor b;
    outputs(6785) <= not b;
    outputs(6786) <= not (a xor b);
    outputs(6787) <= not (a or b);
    outputs(6788) <= a or b;
    outputs(6789) <= not (a and b);
    outputs(6790) <= b;
    outputs(6791) <= not (a xor b);
    outputs(6792) <= not b;
    outputs(6793) <= a xor b;
    outputs(6794) <= a and not b;
    outputs(6795) <= not b;
    outputs(6796) <= b and not a;
    outputs(6797) <= not a;
    outputs(6798) <= a xor b;
    outputs(6799) <= a;
    outputs(6800) <= not a;
    outputs(6801) <= a and not b;
    outputs(6802) <= not (a and b);
    outputs(6803) <= a and b;
    outputs(6804) <= a xor b;
    outputs(6805) <= not a;
    outputs(6806) <= a xor b;
    outputs(6807) <= not a or b;
    outputs(6808) <= not b;
    outputs(6809) <= not b;
    outputs(6810) <= not b;
    outputs(6811) <= a;
    outputs(6812) <= a or b;
    outputs(6813) <= not a;
    outputs(6814) <= not (a xor b);
    outputs(6815) <= not (a xor b);
    outputs(6816) <= a and b;
    outputs(6817) <= not a;
    outputs(6818) <= b;
    outputs(6819) <= b and not a;
    outputs(6820) <= not (a xor b);
    outputs(6821) <= a xor b;
    outputs(6822) <= not b;
    outputs(6823) <= not (a xor b);
    outputs(6824) <= a;
    outputs(6825) <= not (a xor b);
    outputs(6826) <= a and not b;
    outputs(6827) <= a;
    outputs(6828) <= b;
    outputs(6829) <= not a or b;
    outputs(6830) <= a xor b;
    outputs(6831) <= not b;
    outputs(6832) <= a;
    outputs(6833) <= a and b;
    outputs(6834) <= b and not a;
    outputs(6835) <= a and not b;
    outputs(6836) <= not b or a;
    outputs(6837) <= a or b;
    outputs(6838) <= not a;
    outputs(6839) <= not b;
    outputs(6840) <= a;
    outputs(6841) <= not (a xor b);
    outputs(6842) <= not b;
    outputs(6843) <= a;
    outputs(6844) <= not a;
    outputs(6845) <= not b or a;
    outputs(6846) <= not b or a;
    outputs(6847) <= not (a xor b);
    outputs(6848) <= a xor b;
    outputs(6849) <= not b or a;
    outputs(6850) <= not b or a;
    outputs(6851) <= a xor b;
    outputs(6852) <= not b;
    outputs(6853) <= not (a xor b);
    outputs(6854) <= not (a or b);
    outputs(6855) <= b;
    outputs(6856) <= b and not a;
    outputs(6857) <= a or b;
    outputs(6858) <= not b or a;
    outputs(6859) <= not (a and b);
    outputs(6860) <= b;
    outputs(6861) <= not (a xor b);
    outputs(6862) <= a xor b;
    outputs(6863) <= a and not b;
    outputs(6864) <= b;
    outputs(6865) <= not a;
    outputs(6866) <= a and not b;
    outputs(6867) <= a xor b;
    outputs(6868) <= not a;
    outputs(6869) <= a and not b;
    outputs(6870) <= not a or b;
    outputs(6871) <= a;
    outputs(6872) <= not a;
    outputs(6873) <= not b;
    outputs(6874) <= not (a or b);
    outputs(6875) <= not a or b;
    outputs(6876) <= not b;
    outputs(6877) <= not a or b;
    outputs(6878) <= b;
    outputs(6879) <= not (a xor b);
    outputs(6880) <= not (a and b);
    outputs(6881) <= b and not a;
    outputs(6882) <= not b;
    outputs(6883) <= a xor b;
    outputs(6884) <= not a;
    outputs(6885) <= not a;
    outputs(6886) <= not (a xor b);
    outputs(6887) <= not b or a;
    outputs(6888) <= not (a or b);
    outputs(6889) <= not b or a;
    outputs(6890) <= a;
    outputs(6891) <= a and b;
    outputs(6892) <= not (a or b);
    outputs(6893) <= not b;
    outputs(6894) <= a and b;
    outputs(6895) <= not (a or b);
    outputs(6896) <= not b or a;
    outputs(6897) <= not (a or b);
    outputs(6898) <= not (a or b);
    outputs(6899) <= a;
    outputs(6900) <= a and b;
    outputs(6901) <= b;
    outputs(6902) <= a xor b;
    outputs(6903) <= not b;
    outputs(6904) <= not b or a;
    outputs(6905) <= not a or b;
    outputs(6906) <= b and not a;
    outputs(6907) <= not a;
    outputs(6908) <= a and not b;
    outputs(6909) <= b;
    outputs(6910) <= not (a and b);
    outputs(6911) <= a;
    outputs(6912) <= not a;
    outputs(6913) <= not a or b;
    outputs(6914) <= not b;
    outputs(6915) <= not (a or b);
    outputs(6916) <= not b or a;
    outputs(6917) <= not a;
    outputs(6918) <= a xor b;
    outputs(6919) <= not (a xor b);
    outputs(6920) <= a or b;
    outputs(6921) <= a xor b;
    outputs(6922) <= not a;
    outputs(6923) <= a and b;
    outputs(6924) <= not a;
    outputs(6925) <= a and b;
    outputs(6926) <= not b;
    outputs(6927) <= a xor b;
    outputs(6928) <= a;
    outputs(6929) <= a and b;
    outputs(6930) <= a;
    outputs(6931) <= b and not a;
    outputs(6932) <= a and not b;
    outputs(6933) <= a;
    outputs(6934) <= a and not b;
    outputs(6935) <= a and b;
    outputs(6936) <= a and not b;
    outputs(6937) <= b and not a;
    outputs(6938) <= a and b;
    outputs(6939) <= a or b;
    outputs(6940) <= not (a xor b);
    outputs(6941) <= a;
    outputs(6942) <= b;
    outputs(6943) <= not a;
    outputs(6944) <= a and b;
    outputs(6945) <= not b or a;
    outputs(6946) <= not (a or b);
    outputs(6947) <= not b;
    outputs(6948) <= not a;
    outputs(6949) <= b and not a;
    outputs(6950) <= not b;
    outputs(6951) <= a;
    outputs(6952) <= a xor b;
    outputs(6953) <= a and not b;
    outputs(6954) <= not a;
    outputs(6955) <= a and not b;
    outputs(6956) <= a;
    outputs(6957) <= not a or b;
    outputs(6958) <= a;
    outputs(6959) <= a xor b;
    outputs(6960) <= a or b;
    outputs(6961) <= not (a or b);
    outputs(6962) <= a xor b;
    outputs(6963) <= not b;
    outputs(6964) <= b;
    outputs(6965) <= b and not a;
    outputs(6966) <= b;
    outputs(6967) <= b;
    outputs(6968) <= not b;
    outputs(6969) <= b;
    outputs(6970) <= b and not a;
    outputs(6971) <= a xor b;
    outputs(6972) <= not a;
    outputs(6973) <= a and b;
    outputs(6974) <= not b;
    outputs(6975) <= a and not b;
    outputs(6976) <= not (a or b);
    outputs(6977) <= a and b;
    outputs(6978) <= a;
    outputs(6979) <= not a;
    outputs(6980) <= a xor b;
    outputs(6981) <= not (a or b);
    outputs(6982) <= not a or b;
    outputs(6983) <= a;
    outputs(6984) <= b;
    outputs(6985) <= not (a or b);
    outputs(6986) <= not (a or b);
    outputs(6987) <= a and not b;
    outputs(6988) <= not (a xor b);
    outputs(6989) <= a;
    outputs(6990) <= a and b;
    outputs(6991) <= a xor b;
    outputs(6992) <= not (a or b);
    outputs(6993) <= not (a and b);
    outputs(6994) <= a xor b;
    outputs(6995) <= b and not a;
    outputs(6996) <= not (a xor b);
    outputs(6997) <= a and b;
    outputs(6998) <= not (a or b);
    outputs(6999) <= not (a xor b);
    outputs(7000) <= not b or a;
    outputs(7001) <= not b;
    outputs(7002) <= b and not a;
    outputs(7003) <= not (a xor b);
    outputs(7004) <= not (a xor b);
    outputs(7005) <= a;
    outputs(7006) <= a and b;
    outputs(7007) <= a and b;
    outputs(7008) <= not b or a;
    outputs(7009) <= not (a or b);
    outputs(7010) <= b and not a;
    outputs(7011) <= not a;
    outputs(7012) <= a;
    outputs(7013) <= a and b;
    outputs(7014) <= not (a xor b);
    outputs(7015) <= not (a or b);
    outputs(7016) <= a;
    outputs(7017) <= a and b;
    outputs(7018) <= b and not a;
    outputs(7019) <= not b;
    outputs(7020) <= a and not b;
    outputs(7021) <= not b or a;
    outputs(7022) <= not a;
    outputs(7023) <= not (a xor b);
    outputs(7024) <= a and b;
    outputs(7025) <= a and not b;
    outputs(7026) <= a and not b;
    outputs(7027) <= not (a or b);
    outputs(7028) <= a or b;
    outputs(7029) <= a and b;
    outputs(7030) <= a;
    outputs(7031) <= a and not b;
    outputs(7032) <= not (a xor b);
    outputs(7033) <= not (a or b);
    outputs(7034) <= not a or b;
    outputs(7035) <= a xor b;
    outputs(7036) <= not (a xor b);
    outputs(7037) <= not b or a;
    outputs(7038) <= a and b;
    outputs(7039) <= not (a xor b);
    outputs(7040) <= a xor b;
    outputs(7041) <= not (a xor b);
    outputs(7042) <= b;
    outputs(7043) <= not a;
    outputs(7044) <= b and not a;
    outputs(7045) <= not a;
    outputs(7046) <= b and not a;
    outputs(7047) <= not (a xor b);
    outputs(7048) <= not (a xor b);
    outputs(7049) <= a and not b;
    outputs(7050) <= not a;
    outputs(7051) <= b and not a;
    outputs(7052) <= not (a xor b);
    outputs(7053) <= not b;
    outputs(7054) <= not b;
    outputs(7055) <= b;
    outputs(7056) <= a and b;
    outputs(7057) <= not a;
    outputs(7058) <= a and not b;
    outputs(7059) <= a xor b;
    outputs(7060) <= a xor b;
    outputs(7061) <= b;
    outputs(7062) <= not (a or b);
    outputs(7063) <= b;
    outputs(7064) <= not (a xor b);
    outputs(7065) <= b and not a;
    outputs(7066) <= a and not b;
    outputs(7067) <= not b;
    outputs(7068) <= a and not b;
    outputs(7069) <= not (a xor b);
    outputs(7070) <= b and not a;
    outputs(7071) <= not (a xor b);
    outputs(7072) <= a and b;
    outputs(7073) <= not (a or b);
    outputs(7074) <= a and b;
    outputs(7075) <= b;
    outputs(7076) <= not b or a;
    outputs(7077) <= a;
    outputs(7078) <= a and b;
    outputs(7079) <= a xor b;
    outputs(7080) <= not (a or b);
    outputs(7081) <= not a;
    outputs(7082) <= a xor b;
    outputs(7083) <= not b;
    outputs(7084) <= a and b;
    outputs(7085) <= not (a xor b);
    outputs(7086) <= b;
    outputs(7087) <= not (a xor b);
    outputs(7088) <= not a;
    outputs(7089) <= not b or a;
    outputs(7090) <= b;
    outputs(7091) <= a;
    outputs(7092) <= not b;
    outputs(7093) <= a and b;
    outputs(7094) <= not (a xor b);
    outputs(7095) <= a;
    outputs(7096) <= not (a or b);
    outputs(7097) <= a and not b;
    outputs(7098) <= not (a xor b);
    outputs(7099) <= a and not b;
    outputs(7100) <= b and not a;
    outputs(7101) <= a xor b;
    outputs(7102) <= not (a xor b);
    outputs(7103) <= a and b;
    outputs(7104) <= a and b;
    outputs(7105) <= a and not b;
    outputs(7106) <= b;
    outputs(7107) <= a and b;
    outputs(7108) <= b;
    outputs(7109) <= a;
    outputs(7110) <= not (a and b);
    outputs(7111) <= a and not b;
    outputs(7112) <= not b;
    outputs(7113) <= a;
    outputs(7114) <= not (a xor b);
    outputs(7115) <= a and b;
    outputs(7116) <= b and not a;
    outputs(7117) <= a xor b;
    outputs(7118) <= b;
    outputs(7119) <= not b;
    outputs(7120) <= a and not b;
    outputs(7121) <= not (a xor b);
    outputs(7122) <= not a;
    outputs(7123) <= not (a or b);
    outputs(7124) <= not a;
    outputs(7125) <= not b;
    outputs(7126) <= b;
    outputs(7127) <= not (a or b);
    outputs(7128) <= not b;
    outputs(7129) <= not (a or b);
    outputs(7130) <= a xor b;
    outputs(7131) <= not (a and b);
    outputs(7132) <= not a;
    outputs(7133) <= a;
    outputs(7134) <= a;
    outputs(7135) <= a or b;
    outputs(7136) <= b;
    outputs(7137) <= a;
    outputs(7138) <= not a;
    outputs(7139) <= not b or a;
    outputs(7140) <= b;
    outputs(7141) <= a xor b;
    outputs(7142) <= a xor b;
    outputs(7143) <= a xor b;
    outputs(7144) <= a and not b;
    outputs(7145) <= not (a or b);
    outputs(7146) <= not a;
    outputs(7147) <= b and not a;
    outputs(7148) <= a and not b;
    outputs(7149) <= a and b;
    outputs(7150) <= a and b;
    outputs(7151) <= not a or b;
    outputs(7152) <= a xor b;
    outputs(7153) <= a;
    outputs(7154) <= b and not a;
    outputs(7155) <= b and not a;
    outputs(7156) <= not (a or b);
    outputs(7157) <= not b;
    outputs(7158) <= not b;
    outputs(7159) <= not (a or b);
    outputs(7160) <= a xor b;
    outputs(7161) <= a xor b;
    outputs(7162) <= b and not a;
    outputs(7163) <= not a;
    outputs(7164) <= not b;
    outputs(7165) <= a or b;
    outputs(7166) <= not (a or b);
    outputs(7167) <= not (a xor b);
    outputs(7168) <= not (a or b);
    outputs(7169) <= b;
    outputs(7170) <= b;
    outputs(7171) <= a;
    outputs(7172) <= b;
    outputs(7173) <= not (a xor b);
    outputs(7174) <= b and not a;
    outputs(7175) <= not (a or b);
    outputs(7176) <= not (a or b);
    outputs(7177) <= not (a or b);
    outputs(7178) <= not b;
    outputs(7179) <= b and not a;
    outputs(7180) <= a and b;
    outputs(7181) <= a xor b;
    outputs(7182) <= not (a xor b);
    outputs(7183) <= not (a xor b);
    outputs(7184) <= not b;
    outputs(7185) <= a;
    outputs(7186) <= a xor b;
    outputs(7187) <= not (a xor b);
    outputs(7188) <= a xor b;
    outputs(7189) <= not b;
    outputs(7190) <= a xor b;
    outputs(7191) <= not a;
    outputs(7192) <= a xor b;
    outputs(7193) <= not (a or b);
    outputs(7194) <= a xor b;
    outputs(7195) <= b and not a;
    outputs(7196) <= a and not b;
    outputs(7197) <= not (a or b);
    outputs(7198) <= not a;
    outputs(7199) <= b and not a;
    outputs(7200) <= a and b;
    outputs(7201) <= a and b;
    outputs(7202) <= a and not b;
    outputs(7203) <= not (a xor b);
    outputs(7204) <= a;
    outputs(7205) <= not a;
    outputs(7206) <= not (a or b);
    outputs(7207) <= not b;
    outputs(7208) <= a and not b;
    outputs(7209) <= not b;
    outputs(7210) <= b and not a;
    outputs(7211) <= not (a or b);
    outputs(7212) <= b and not a;
    outputs(7213) <= a and not b;
    outputs(7214) <= not (a and b);
    outputs(7215) <= a xor b;
    outputs(7216) <= not b;
    outputs(7217) <= a and b;
    outputs(7218) <= not (a and b);
    outputs(7219) <= not b;
    outputs(7220) <= a and not b;
    outputs(7221) <= not (a xor b);
    outputs(7222) <= a and not b;
    outputs(7223) <= not (a xor b);
    outputs(7224) <= b;
    outputs(7225) <= not (a xor b);
    outputs(7226) <= not (a xor b);
    outputs(7227) <= a and not b;
    outputs(7228) <= a xor b;
    outputs(7229) <= not a or b;
    outputs(7230) <= not (a xor b);
    outputs(7231) <= b;
    outputs(7232) <= not b;
    outputs(7233) <= not b or a;
    outputs(7234) <= not b;
    outputs(7235) <= not (a or b);
    outputs(7236) <= a xor b;
    outputs(7237) <= not (a or b);
    outputs(7238) <= a or b;
    outputs(7239) <= a xor b;
    outputs(7240) <= a;
    outputs(7241) <= not (a or b);
    outputs(7242) <= not (a xor b);
    outputs(7243) <= not (a or b);
    outputs(7244) <= not (a or b);
    outputs(7245) <= a and not b;
    outputs(7246) <= not (a or b);
    outputs(7247) <= not a;
    outputs(7248) <= b;
    outputs(7249) <= a xor b;
    outputs(7250) <= not b;
    outputs(7251) <= not b;
    outputs(7252) <= b;
    outputs(7253) <= not (a xor b);
    outputs(7254) <= not (a or b);
    outputs(7255) <= not a;
    outputs(7256) <= not (a or b);
    outputs(7257) <= b;
    outputs(7258) <= not b or a;
    outputs(7259) <= a and not b;
    outputs(7260) <= not (a or b);
    outputs(7261) <= a and b;
    outputs(7262) <= b;
    outputs(7263) <= not (a and b);
    outputs(7264) <= not (a xor b);
    outputs(7265) <= a and not b;
    outputs(7266) <= not (a or b);
    outputs(7267) <= a and not b;
    outputs(7268) <= a xor b;
    outputs(7269) <= a and b;
    outputs(7270) <= not (a xor b);
    outputs(7271) <= a and b;
    outputs(7272) <= a and not b;
    outputs(7273) <= not (a xor b);
    outputs(7274) <= not a;
    outputs(7275) <= not a;
    outputs(7276) <= not b;
    outputs(7277) <= a xor b;
    outputs(7278) <= b and not a;
    outputs(7279) <= not (a xor b);
    outputs(7280) <= a;
    outputs(7281) <= a and not b;
    outputs(7282) <= a and not b;
    outputs(7283) <= b and not a;
    outputs(7284) <= not (a or b);
    outputs(7285) <= a and not b;
    outputs(7286) <= a and not b;
    outputs(7287) <= a and not b;
    outputs(7288) <= a or b;
    outputs(7289) <= a;
    outputs(7290) <= not b or a;
    outputs(7291) <= b and not a;
    outputs(7292) <= not (a xor b);
    outputs(7293) <= a and b;
    outputs(7294) <= a xor b;
    outputs(7295) <= not b;
    outputs(7296) <= b and not a;
    outputs(7297) <= not (a xor b);
    outputs(7298) <= a and b;
    outputs(7299) <= not b;
    outputs(7300) <= not (a xor b);
    outputs(7301) <= b and not a;
    outputs(7302) <= a and b;
    outputs(7303) <= a xor b;
    outputs(7304) <= b;
    outputs(7305) <= a and not b;
    outputs(7306) <= b;
    outputs(7307) <= a and not b;
    outputs(7308) <= not (a or b);
    outputs(7309) <= a;
    outputs(7310) <= not b;
    outputs(7311) <= not b;
    outputs(7312) <= a and b;
    outputs(7313) <= a and b;
    outputs(7314) <= not (a xor b);
    outputs(7315) <= b and not a;
    outputs(7316) <= not a;
    outputs(7317) <= not b or a;
    outputs(7318) <= a xor b;
    outputs(7319) <= a and b;
    outputs(7320) <= a and b;
    outputs(7321) <= b;
    outputs(7322) <= b;
    outputs(7323) <= a xor b;
    outputs(7324) <= a xor b;
    outputs(7325) <= b and not a;
    outputs(7326) <= not (a xor b);
    outputs(7327) <= not b;
    outputs(7328) <= a and not b;
    outputs(7329) <= a xor b;
    outputs(7330) <= a;
    outputs(7331) <= not (a or b);
    outputs(7332) <= a;
    outputs(7333) <= not b;
    outputs(7334) <= a and b;
    outputs(7335) <= a xor b;
    outputs(7336) <= a;
    outputs(7337) <= a and not b;
    outputs(7338) <= not (a or b);
    outputs(7339) <= a and not b;
    outputs(7340) <= not (a or b);
    outputs(7341) <= a xor b;
    outputs(7342) <= not a;
    outputs(7343) <= not (a or b);
    outputs(7344) <= b and not a;
    outputs(7345) <= b and not a;
    outputs(7346) <= a and not b;
    outputs(7347) <= a and not b;
    outputs(7348) <= a xor b;
    outputs(7349) <= not a;
    outputs(7350) <= a and not b;
    outputs(7351) <= a and b;
    outputs(7352) <= a and b;
    outputs(7353) <= not (a xor b);
    outputs(7354) <= a and b;
    outputs(7355) <= not a;
    outputs(7356) <= not (a xor b);
    outputs(7357) <= not (a or b);
    outputs(7358) <= not b;
    outputs(7359) <= a and not b;
    outputs(7360) <= a and not b;
    outputs(7361) <= not a;
    outputs(7362) <= not (a xor b);
    outputs(7363) <= not a;
    outputs(7364) <= not a;
    outputs(7365) <= a and b;
    outputs(7366) <= not (a or b);
    outputs(7367) <= b and not a;
    outputs(7368) <= a and not b;
    outputs(7369) <= not (a or b);
    outputs(7370) <= not (a xor b);
    outputs(7371) <= a and not b;
    outputs(7372) <= a xor b;
    outputs(7373) <= b;
    outputs(7374) <= b;
    outputs(7375) <= b and not a;
    outputs(7376) <= a xor b;
    outputs(7377) <= b;
    outputs(7378) <= not b;
    outputs(7379) <= a and b;
    outputs(7380) <= not (a and b);
    outputs(7381) <= a and not b;
    outputs(7382) <= b;
    outputs(7383) <= not (a xor b);
    outputs(7384) <= not a;
    outputs(7385) <= a and b;
    outputs(7386) <= not a;
    outputs(7387) <= a and b;
    outputs(7388) <= not (a xor b);
    outputs(7389) <= not (a xor b);
    outputs(7390) <= a and not b;
    outputs(7391) <= not (a or b);
    outputs(7392) <= not b;
    outputs(7393) <= a xor b;
    outputs(7394) <= not b;
    outputs(7395) <= not (a or b);
    outputs(7396) <= a and b;
    outputs(7397) <= not b or a;
    outputs(7398) <= not (a or b);
    outputs(7399) <= not (a xor b);
    outputs(7400) <= a and not b;
    outputs(7401) <= not b;
    outputs(7402) <= not b;
    outputs(7403) <= not b or a;
    outputs(7404) <= not b;
    outputs(7405) <= b;
    outputs(7406) <= not (a xor b);
    outputs(7407) <= not (a or b);
    outputs(7408) <= a xor b;
    outputs(7409) <= b and not a;
    outputs(7410) <= not (a or b);
    outputs(7411) <= a or b;
    outputs(7412) <= not (a and b);
    outputs(7413) <= a xor b;
    outputs(7414) <= not (a xor b);
    outputs(7415) <= b and not a;
    outputs(7416) <= not (a or b);
    outputs(7417) <= b and not a;
    outputs(7418) <= a and not b;
    outputs(7419) <= a and b;
    outputs(7420) <= b;
    outputs(7421) <= a xor b;
    outputs(7422) <= not (a and b);
    outputs(7423) <= a or b;
    outputs(7424) <= not (a xor b);
    outputs(7425) <= not (a or b);
    outputs(7426) <= not b;
    outputs(7427) <= a and not b;
    outputs(7428) <= a and not b;
    outputs(7429) <= b;
    outputs(7430) <= not a;
    outputs(7431) <= a and b;
    outputs(7432) <= b;
    outputs(7433) <= a;
    outputs(7434) <= not a or b;
    outputs(7435) <= not a or b;
    outputs(7436) <= a and not b;
    outputs(7437) <= not a;
    outputs(7438) <= b and not a;
    outputs(7439) <= not (a xor b);
    outputs(7440) <= a and not b;
    outputs(7441) <= a and b;
    outputs(7442) <= not b;
    outputs(7443) <= a and not b;
    outputs(7444) <= not b;
    outputs(7445) <= a and not b;
    outputs(7446) <= a and b;
    outputs(7447) <= b and not a;
    outputs(7448) <= not (a or b);
    outputs(7449) <= a xor b;
    outputs(7450) <= not (a or b);
    outputs(7451) <= a and b;
    outputs(7452) <= a xor b;
    outputs(7453) <= not a;
    outputs(7454) <= not a;
    outputs(7455) <= not (a xor b);
    outputs(7456) <= b;
    outputs(7457) <= b;
    outputs(7458) <= not b or a;
    outputs(7459) <= a xor b;
    outputs(7460) <= a and b;
    outputs(7461) <= not b;
    outputs(7462) <= not a;
    outputs(7463) <= b and not a;
    outputs(7464) <= a and not b;
    outputs(7465) <= a xor b;
    outputs(7466) <= b and not a;
    outputs(7467) <= a or b;
    outputs(7468) <= a xor b;
    outputs(7469) <= not b;
    outputs(7470) <= not (a xor b);
    outputs(7471) <= b and not a;
    outputs(7472) <= b and not a;
    outputs(7473) <= not (a and b);
    outputs(7474) <= a or b;
    outputs(7475) <= a and b;
    outputs(7476) <= a and b;
    outputs(7477) <= not (a xor b);
    outputs(7478) <= a;
    outputs(7479) <= not (a and b);
    outputs(7480) <= a and not b;
    outputs(7481) <= not a or b;
    outputs(7482) <= not b;
    outputs(7483) <= b and not a;
    outputs(7484) <= not (a xor b);
    outputs(7485) <= a xor b;
    outputs(7486) <= a;
    outputs(7487) <= a;
    outputs(7488) <= not (a or b);
    outputs(7489) <= not b;
    outputs(7490) <= not b;
    outputs(7491) <= not b;
    outputs(7492) <= a and b;
    outputs(7493) <= not a;
    outputs(7494) <= a or b;
    outputs(7495) <= a xor b;
    outputs(7496) <= not (a and b);
    outputs(7497) <= a and not b;
    outputs(7498) <= b and not a;
    outputs(7499) <= a and b;
    outputs(7500) <= a xor b;
    outputs(7501) <= a and not b;
    outputs(7502) <= not (a xor b);
    outputs(7503) <= not (a xor b);
    outputs(7504) <= not (a xor b);
    outputs(7505) <= b and not a;
    outputs(7506) <= b and not a;
    outputs(7507) <= a xor b;
    outputs(7508) <= b and not a;
    outputs(7509) <= a xor b;
    outputs(7510) <= a and b;
    outputs(7511) <= a and not b;
    outputs(7512) <= a and not b;
    outputs(7513) <= not (a xor b);
    outputs(7514) <= a;
    outputs(7515) <= b;
    outputs(7516) <= a;
    outputs(7517) <= not (a and b);
    outputs(7518) <= b and not a;
    outputs(7519) <= not (a xor b);
    outputs(7520) <= not b;
    outputs(7521) <= not (a xor b);
    outputs(7522) <= b;
    outputs(7523) <= b and not a;
    outputs(7524) <= a or b;
    outputs(7525) <= not (a and b);
    outputs(7526) <= a and not b;
    outputs(7527) <= not b;
    outputs(7528) <= b;
    outputs(7529) <= not b;
    outputs(7530) <= not (a and b);
    outputs(7531) <= not a;
    outputs(7532) <= a xor b;
    outputs(7533) <= a and not b;
    outputs(7534) <= a or b;
    outputs(7535) <= a and not b;
    outputs(7536) <= not a or b;
    outputs(7537) <= a and b;
    outputs(7538) <= not a;
    outputs(7539) <= not b or a;
    outputs(7540) <= a and b;
    outputs(7541) <= not b;
    outputs(7542) <= a and not b;
    outputs(7543) <= not b or a;
    outputs(7544) <= a xor b;
    outputs(7545) <= not (a xor b);
    outputs(7546) <= a;
    outputs(7547) <= not (a or b);
    outputs(7548) <= not a;
    outputs(7549) <= not (a xor b);
    outputs(7550) <= a and not b;
    outputs(7551) <= a;
    outputs(7552) <= a and not b;
    outputs(7553) <= b and not a;
    outputs(7554) <= not (a xor b);
    outputs(7555) <= not b;
    outputs(7556) <= a;
    outputs(7557) <= a and not b;
    outputs(7558) <= not (a xor b);
    outputs(7559) <= not a;
    outputs(7560) <= not a or b;
    outputs(7561) <= a;
    outputs(7562) <= a;
    outputs(7563) <= not (a or b);
    outputs(7564) <= a xor b;
    outputs(7565) <= a and not b;
    outputs(7566) <= not b;
    outputs(7567) <= not (a xor b);
    outputs(7568) <= a or b;
    outputs(7569) <= not (a or b);
    outputs(7570) <= a and not b;
    outputs(7571) <= a and b;
    outputs(7572) <= a and b;
    outputs(7573) <= not b;
    outputs(7574) <= b;
    outputs(7575) <= not (a and b);
    outputs(7576) <= not (a xor b);
    outputs(7577) <= not (a xor b);
    outputs(7578) <= not b;
    outputs(7579) <= not b;
    outputs(7580) <= not (a xor b);
    outputs(7581) <= a;
    outputs(7582) <= a xor b;
    outputs(7583) <= not b;
    outputs(7584) <= a and not b;
    outputs(7585) <= a and b;
    outputs(7586) <= b and not a;
    outputs(7587) <= a;
    outputs(7588) <= not (a or b);
    outputs(7589) <= a and not b;
    outputs(7590) <= not b;
    outputs(7591) <= a and b;
    outputs(7592) <= a and b;
    outputs(7593) <= a;
    outputs(7594) <= not b;
    outputs(7595) <= a;
    outputs(7596) <= a xor b;
    outputs(7597) <= a;
    outputs(7598) <= a;
    outputs(7599) <= a and b;
    outputs(7600) <= not b;
    outputs(7601) <= not a or b;
    outputs(7602) <= a;
    outputs(7603) <= a or b;
    outputs(7604) <= not (a xor b);
    outputs(7605) <= not (a xor b);
    outputs(7606) <= a;
    outputs(7607) <= not (a xor b);
    outputs(7608) <= a and not b;
    outputs(7609) <= a xor b;
    outputs(7610) <= b and not a;
    outputs(7611) <= a;
    outputs(7612) <= a;
    outputs(7613) <= not b;
    outputs(7614) <= a;
    outputs(7615) <= not (a xor b);
    outputs(7616) <= not a or b;
    outputs(7617) <= a and not b;
    outputs(7618) <= not (a or b);
    outputs(7619) <= not b;
    outputs(7620) <= a and not b;
    outputs(7621) <= a;
    outputs(7622) <= a xor b;
    outputs(7623) <= b;
    outputs(7624) <= b and not a;
    outputs(7625) <= a;
    outputs(7626) <= b and not a;
    outputs(7627) <= a and b;
    outputs(7628) <= not (a xor b);
    outputs(7629) <= a and b;
    outputs(7630) <= a and b;
    outputs(7631) <= not (a or b);
    outputs(7632) <= a and b;
    outputs(7633) <= a and not b;
    outputs(7634) <= not a;
    outputs(7635) <= b;
    outputs(7636) <= not (a or b);
    outputs(7637) <= a and not b;
    outputs(7638) <= a and b;
    outputs(7639) <= b;
    outputs(7640) <= not (a xor b);
    outputs(7641) <= b;
    outputs(7642) <= not a;
    outputs(7643) <= a and b;
    outputs(7644) <= not b;
    outputs(7645) <= a and not b;
    outputs(7646) <= not a;
    outputs(7647) <= not (a or b);
    outputs(7648) <= not b;
    outputs(7649) <= a and not b;
    outputs(7650) <= not b or a;
    outputs(7651) <= b and not a;
    outputs(7652) <= a;
    outputs(7653) <= a and not b;
    outputs(7654) <= not (a xor b);
    outputs(7655) <= a and b;
    outputs(7656) <= b;
    outputs(7657) <= not b;
    outputs(7658) <= a xor b;
    outputs(7659) <= a;
    outputs(7660) <= a or b;
    outputs(7661) <= b and not a;
    outputs(7662) <= a;
    outputs(7663) <= not a;
    outputs(7664) <= not b;
    outputs(7665) <= not (a xor b);
    outputs(7666) <= b;
    outputs(7667) <= not (a and b);
    outputs(7668) <= b;
    outputs(7669) <= b;
    outputs(7670) <= not (a xor b);
    outputs(7671) <= b and not a;
    outputs(7672) <= b;
    outputs(7673) <= a xor b;
    outputs(7674) <= b and not a;
    outputs(7675) <= not (a or b);
    outputs(7676) <= b;
    outputs(7677) <= not a;
    outputs(7678) <= not a;
    outputs(7679) <= a and b;
end Behavioral;
