library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(5119 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(5119 downto 0);

begin

    layer0_outputs(0) <= inputs(243);
    layer0_outputs(1) <= not(inputs(244));
    layer0_outputs(2) <= (inputs(164)) or (inputs(174));
    layer0_outputs(3) <= not(inputs(184));
    layer0_outputs(4) <= not(inputs(249));
    layer0_outputs(5) <= not((inputs(191)) or (inputs(90)));
    layer0_outputs(6) <= not(inputs(153)) or (inputs(154));
    layer0_outputs(7) <= not(inputs(234));
    layer0_outputs(8) <= not((inputs(127)) or (inputs(194)));
    layer0_outputs(9) <= not(inputs(224));
    layer0_outputs(10) <= not(inputs(23)) or (inputs(181));
    layer0_outputs(11) <= (inputs(76)) or (inputs(126));
    layer0_outputs(12) <= (inputs(143)) or (inputs(34));
    layer0_outputs(13) <= not((inputs(169)) or (inputs(3)));
    layer0_outputs(14) <= not((inputs(52)) xor (inputs(234)));
    layer0_outputs(15) <= not(inputs(20)) or (inputs(217));
    layer0_outputs(16) <= not(inputs(176)) or (inputs(149));
    layer0_outputs(17) <= not((inputs(183)) xor (inputs(44)));
    layer0_outputs(18) <= (inputs(107)) and not (inputs(11));
    layer0_outputs(19) <= inputs(109);
    layer0_outputs(20) <= (inputs(54)) or (inputs(117));
    layer0_outputs(21) <= (inputs(207)) or (inputs(221));
    layer0_outputs(22) <= not((inputs(26)) or (inputs(246)));
    layer0_outputs(23) <= (inputs(9)) or (inputs(96));
    layer0_outputs(24) <= (inputs(99)) and not (inputs(17));
    layer0_outputs(25) <= (inputs(119)) or (inputs(31));
    layer0_outputs(26) <= (inputs(105)) and not (inputs(231));
    layer0_outputs(27) <= (inputs(136)) or (inputs(182));
    layer0_outputs(28) <= (inputs(145)) or (inputs(192));
    layer0_outputs(29) <= (inputs(118)) or (inputs(169));
    layer0_outputs(30) <= not(inputs(105)) or (inputs(69));
    layer0_outputs(31) <= not(inputs(150));
    layer0_outputs(32) <= (inputs(197)) and not (inputs(45));
    layer0_outputs(33) <= not(inputs(45)) or (inputs(197));
    layer0_outputs(34) <= (inputs(252)) or (inputs(178));
    layer0_outputs(35) <= '1';
    layer0_outputs(36) <= not((inputs(196)) xor (inputs(28)));
    layer0_outputs(37) <= not((inputs(206)) or (inputs(209)));
    layer0_outputs(38) <= not((inputs(61)) or (inputs(151)));
    layer0_outputs(39) <= not((inputs(2)) and (inputs(174)));
    layer0_outputs(40) <= not(inputs(8));
    layer0_outputs(41) <= inputs(24);
    layer0_outputs(42) <= inputs(43);
    layer0_outputs(43) <= inputs(98);
    layer0_outputs(44) <= not((inputs(162)) or (inputs(177)));
    layer0_outputs(45) <= not(inputs(148));
    layer0_outputs(46) <= not(inputs(207));
    layer0_outputs(47) <= not(inputs(207)) or (inputs(251));
    layer0_outputs(48) <= not((inputs(166)) or (inputs(196)));
    layer0_outputs(49) <= not((inputs(186)) or (inputs(34)));
    layer0_outputs(50) <= inputs(59);
    layer0_outputs(51) <= not((inputs(85)) or (inputs(74)));
    layer0_outputs(52) <= not((inputs(186)) and (inputs(205)));
    layer0_outputs(53) <= '0';
    layer0_outputs(54) <= not((inputs(19)) or (inputs(46)));
    layer0_outputs(55) <= (inputs(28)) xor (inputs(35));
    layer0_outputs(56) <= not(inputs(7));
    layer0_outputs(57) <= inputs(60);
    layer0_outputs(58) <= (inputs(24)) and not (inputs(207));
    layer0_outputs(59) <= not((inputs(85)) or (inputs(222)));
    layer0_outputs(60) <= inputs(113);
    layer0_outputs(61) <= (inputs(201)) and not (inputs(112));
    layer0_outputs(62) <= not((inputs(132)) or (inputs(138)));
    layer0_outputs(63) <= inputs(177);
    layer0_outputs(64) <= inputs(122);
    layer0_outputs(65) <= inputs(89);
    layer0_outputs(66) <= (inputs(48)) or (inputs(190));
    layer0_outputs(67) <= not((inputs(218)) or (inputs(253)));
    layer0_outputs(68) <= not((inputs(187)) or (inputs(48)));
    layer0_outputs(69) <= not(inputs(36)) or (inputs(128));
    layer0_outputs(70) <= not(inputs(117)) or (inputs(223));
    layer0_outputs(71) <= inputs(89);
    layer0_outputs(72) <= (inputs(194)) and not (inputs(33));
    layer0_outputs(73) <= not((inputs(76)) or (inputs(149)));
    layer0_outputs(74) <= not(inputs(196));
    layer0_outputs(75) <= inputs(242);
    layer0_outputs(76) <= not(inputs(92)) or (inputs(214));
    layer0_outputs(77) <= inputs(230);
    layer0_outputs(78) <= not(inputs(154));
    layer0_outputs(79) <= inputs(214);
    layer0_outputs(80) <= not(inputs(22)) or (inputs(12));
    layer0_outputs(81) <= inputs(42);
    layer0_outputs(82) <= inputs(147);
    layer0_outputs(83) <= inputs(238);
    layer0_outputs(84) <= (inputs(24)) and (inputs(75));
    layer0_outputs(85) <= not(inputs(52));
    layer0_outputs(86) <= not((inputs(114)) xor (inputs(220)));
    layer0_outputs(87) <= (inputs(136)) and not (inputs(18));
    layer0_outputs(88) <= not(inputs(215));
    layer0_outputs(89) <= (inputs(24)) or (inputs(48));
    layer0_outputs(90) <= not((inputs(113)) xor (inputs(211)));
    layer0_outputs(91) <= inputs(85);
    layer0_outputs(92) <= inputs(182);
    layer0_outputs(93) <= (inputs(115)) and not (inputs(219));
    layer0_outputs(94) <= not(inputs(30)) or (inputs(78));
    layer0_outputs(95) <= not(inputs(189)) or (inputs(34));
    layer0_outputs(96) <= (inputs(109)) and not (inputs(135));
    layer0_outputs(97) <= inputs(245);
    layer0_outputs(98) <= inputs(167);
    layer0_outputs(99) <= not(inputs(121));
    layer0_outputs(100) <= not(inputs(66)) or (inputs(237));
    layer0_outputs(101) <= not((inputs(112)) or (inputs(26)));
    layer0_outputs(102) <= not((inputs(239)) or (inputs(198)));
    layer0_outputs(103) <= not(inputs(145));
    layer0_outputs(104) <= (inputs(124)) or (inputs(236));
    layer0_outputs(105) <= not(inputs(139));
    layer0_outputs(106) <= inputs(133);
    layer0_outputs(107) <= (inputs(187)) xor (inputs(235));
    layer0_outputs(108) <= '1';
    layer0_outputs(109) <= (inputs(27)) and not (inputs(13));
    layer0_outputs(110) <= inputs(24);
    layer0_outputs(111) <= (inputs(4)) or (inputs(242));
    layer0_outputs(112) <= inputs(191);
    layer0_outputs(113) <= not((inputs(232)) xor (inputs(169)));
    layer0_outputs(114) <= not((inputs(241)) xor (inputs(209)));
    layer0_outputs(115) <= inputs(230);
    layer0_outputs(116) <= inputs(121);
    layer0_outputs(117) <= not(inputs(212));
    layer0_outputs(118) <= inputs(106);
    layer0_outputs(119) <= not(inputs(42));
    layer0_outputs(120) <= not(inputs(140)) or (inputs(16));
    layer0_outputs(121) <= (inputs(71)) and not (inputs(236));
    layer0_outputs(122) <= not(inputs(133));
    layer0_outputs(123) <= (inputs(232)) xor (inputs(185));
    layer0_outputs(124) <= (inputs(91)) or (inputs(60));
    layer0_outputs(125) <= not(inputs(105));
    layer0_outputs(126) <= not((inputs(208)) xor (inputs(224)));
    layer0_outputs(127) <= inputs(187);
    layer0_outputs(128) <= not((inputs(220)) xor (inputs(250)));
    layer0_outputs(129) <= not((inputs(126)) xor (inputs(124)));
    layer0_outputs(130) <= not(inputs(134));
    layer0_outputs(131) <= not((inputs(81)) or (inputs(24)));
    layer0_outputs(132) <= not((inputs(150)) or (inputs(162)));
    layer0_outputs(133) <= (inputs(88)) and (inputs(0));
    layer0_outputs(134) <= not((inputs(233)) or (inputs(111)));
    layer0_outputs(135) <= not(inputs(238));
    layer0_outputs(136) <= inputs(148);
    layer0_outputs(137) <= not(inputs(26)) or (inputs(246));
    layer0_outputs(138) <= (inputs(170)) and not (inputs(133));
    layer0_outputs(139) <= not(inputs(212)) or (inputs(89));
    layer0_outputs(140) <= not((inputs(48)) or (inputs(5)));
    layer0_outputs(141) <= not((inputs(165)) or (inputs(130)));
    layer0_outputs(142) <= '0';
    layer0_outputs(143) <= (inputs(153)) or (inputs(114));
    layer0_outputs(144) <= (inputs(218)) or (inputs(205));
    layer0_outputs(145) <= (inputs(114)) and not (inputs(94));
    layer0_outputs(146) <= (inputs(40)) or (inputs(172));
    layer0_outputs(147) <= (inputs(224)) or (inputs(236));
    layer0_outputs(148) <= inputs(120);
    layer0_outputs(149) <= inputs(86);
    layer0_outputs(150) <= (inputs(109)) or (inputs(110));
    layer0_outputs(151) <= (inputs(241)) or (inputs(31));
    layer0_outputs(152) <= not((inputs(41)) xor (inputs(112)));
    layer0_outputs(153) <= not(inputs(245));
    layer0_outputs(154) <= not(inputs(218)) or (inputs(49));
    layer0_outputs(155) <= (inputs(202)) or (inputs(12));
    layer0_outputs(156) <= not((inputs(255)) and (inputs(192)));
    layer0_outputs(157) <= '1';
    layer0_outputs(158) <= '1';
    layer0_outputs(159) <= not(inputs(163));
    layer0_outputs(160) <= (inputs(222)) and not (inputs(214));
    layer0_outputs(161) <= not((inputs(94)) or (inputs(241)));
    layer0_outputs(162) <= not((inputs(23)) or (inputs(141)));
    layer0_outputs(163) <= (inputs(117)) and not (inputs(77));
    layer0_outputs(164) <= (inputs(186)) and not (inputs(51));
    layer0_outputs(165) <= not(inputs(126));
    layer0_outputs(166) <= not((inputs(174)) or (inputs(213)));
    layer0_outputs(167) <= not(inputs(55));
    layer0_outputs(168) <= (inputs(59)) xor (inputs(74));
    layer0_outputs(169) <= not(inputs(36)) or (inputs(158));
    layer0_outputs(170) <= (inputs(45)) and (inputs(39));
    layer0_outputs(171) <= not((inputs(48)) and (inputs(207)));
    layer0_outputs(172) <= (inputs(252)) or (inputs(112));
    layer0_outputs(173) <= not((inputs(230)) or (inputs(194)));
    layer0_outputs(174) <= inputs(229);
    layer0_outputs(175) <= inputs(118);
    layer0_outputs(176) <= inputs(157);
    layer0_outputs(177) <= (inputs(24)) and not (inputs(229));
    layer0_outputs(178) <= inputs(25);
    layer0_outputs(179) <= (inputs(108)) or (inputs(200));
    layer0_outputs(180) <= not((inputs(64)) or (inputs(253)));
    layer0_outputs(181) <= (inputs(232)) and not (inputs(113));
    layer0_outputs(182) <= not(inputs(183)) or (inputs(181));
    layer0_outputs(183) <= not((inputs(101)) or (inputs(145)));
    layer0_outputs(184) <= not(inputs(105));
    layer0_outputs(185) <= '1';
    layer0_outputs(186) <= (inputs(127)) or (inputs(124));
    layer0_outputs(187) <= not(inputs(199));
    layer0_outputs(188) <= (inputs(243)) xor (inputs(10));
    layer0_outputs(189) <= (inputs(123)) and not (inputs(145));
    layer0_outputs(190) <= (inputs(50)) or (inputs(5));
    layer0_outputs(191) <= not(inputs(214));
    layer0_outputs(192) <= (inputs(198)) and not (inputs(113));
    layer0_outputs(193) <= not((inputs(74)) or (inputs(61)));
    layer0_outputs(194) <= (inputs(211)) or (inputs(111));
    layer0_outputs(195) <= not((inputs(173)) xor (inputs(123)));
    layer0_outputs(196) <= (inputs(106)) or (inputs(145));
    layer0_outputs(197) <= not((inputs(25)) or (inputs(124)));
    layer0_outputs(198) <= not((inputs(14)) xor (inputs(199)));
    layer0_outputs(199) <= not(inputs(183)) or (inputs(119));
    layer0_outputs(200) <= not(inputs(64));
    layer0_outputs(201) <= inputs(103);
    layer0_outputs(202) <= inputs(210);
    layer0_outputs(203) <= inputs(199);
    layer0_outputs(204) <= not(inputs(38));
    layer0_outputs(205) <= not(inputs(147));
    layer0_outputs(206) <= (inputs(245)) or (inputs(196));
    layer0_outputs(207) <= (inputs(200)) or (inputs(47));
    layer0_outputs(208) <= (inputs(154)) or (inputs(128));
    layer0_outputs(209) <= '0';
    layer0_outputs(210) <= not(inputs(166));
    layer0_outputs(211) <= not((inputs(151)) and (inputs(250)));
    layer0_outputs(212) <= '0';
    layer0_outputs(213) <= not(inputs(70));
    layer0_outputs(214) <= (inputs(65)) and (inputs(1));
    layer0_outputs(215) <= (inputs(120)) xor (inputs(232));
    layer0_outputs(216) <= not(inputs(100));
    layer0_outputs(217) <= inputs(130);
    layer0_outputs(218) <= not(inputs(140));
    layer0_outputs(219) <= (inputs(62)) xor (inputs(81));
    layer0_outputs(220) <= not((inputs(127)) xor (inputs(204)));
    layer0_outputs(221) <= (inputs(60)) or (inputs(65));
    layer0_outputs(222) <= not(inputs(193));
    layer0_outputs(223) <= (inputs(161)) or (inputs(154));
    layer0_outputs(224) <= inputs(95);
    layer0_outputs(225) <= (inputs(37)) xor (inputs(27));
    layer0_outputs(226) <= (inputs(134)) and not (inputs(1));
    layer0_outputs(227) <= (inputs(167)) and not (inputs(240));
    layer0_outputs(228) <= inputs(225);
    layer0_outputs(229) <= not(inputs(174));
    layer0_outputs(230) <= not((inputs(212)) or (inputs(114)));
    layer0_outputs(231) <= (inputs(226)) xor (inputs(251));
    layer0_outputs(232) <= not((inputs(184)) and (inputs(131)));
    layer0_outputs(233) <= not(inputs(7));
    layer0_outputs(234) <= inputs(164);
    layer0_outputs(235) <= inputs(232);
    layer0_outputs(236) <= (inputs(37)) or (inputs(100));
    layer0_outputs(237) <= inputs(195);
    layer0_outputs(238) <= (inputs(115)) and not (inputs(32));
    layer0_outputs(239) <= not(inputs(254)) or (inputs(200));
    layer0_outputs(240) <= (inputs(68)) or (inputs(202));
    layer0_outputs(241) <= (inputs(146)) or (inputs(158));
    layer0_outputs(242) <= '0';
    layer0_outputs(243) <= not(inputs(158));
    layer0_outputs(244) <= (inputs(8)) or (inputs(194));
    layer0_outputs(245) <= not((inputs(141)) xor (inputs(123)));
    layer0_outputs(246) <= not(inputs(87)) or (inputs(126));
    layer0_outputs(247) <= (inputs(41)) and (inputs(153));
    layer0_outputs(248) <= inputs(135);
    layer0_outputs(249) <= not(inputs(196));
    layer0_outputs(250) <= not((inputs(57)) or (inputs(225)));
    layer0_outputs(251) <= not(inputs(239));
    layer0_outputs(252) <= not(inputs(120));
    layer0_outputs(253) <= not(inputs(229));
    layer0_outputs(254) <= inputs(121);
    layer0_outputs(255) <= not(inputs(195)) or (inputs(46));
    layer0_outputs(256) <= not(inputs(118)) or (inputs(19));
    layer0_outputs(257) <= not(inputs(84));
    layer0_outputs(258) <= not((inputs(155)) and (inputs(226)));
    layer0_outputs(259) <= not((inputs(255)) or (inputs(85)));
    layer0_outputs(260) <= not((inputs(15)) or (inputs(147)));
    layer0_outputs(261) <= (inputs(96)) and not (inputs(80));
    layer0_outputs(262) <= (inputs(15)) or (inputs(212));
    layer0_outputs(263) <= (inputs(3)) and not (inputs(26));
    layer0_outputs(264) <= not((inputs(160)) xor (inputs(113)));
    layer0_outputs(265) <= (inputs(222)) or (inputs(139));
    layer0_outputs(266) <= (inputs(175)) and (inputs(113));
    layer0_outputs(267) <= (inputs(75)) and not (inputs(239));
    layer0_outputs(268) <= not((inputs(27)) xor (inputs(158)));
    layer0_outputs(269) <= not(inputs(239)) or (inputs(142));
    layer0_outputs(270) <= (inputs(231)) and not (inputs(60));
    layer0_outputs(271) <= (inputs(104)) and not (inputs(155));
    layer0_outputs(272) <= not((inputs(110)) xor (inputs(220)));
    layer0_outputs(273) <= (inputs(242)) or (inputs(226));
    layer0_outputs(274) <= not((inputs(138)) or (inputs(159)));
    layer0_outputs(275) <= not((inputs(173)) xor (inputs(171)));
    layer0_outputs(276) <= inputs(51);
    layer0_outputs(277) <= not(inputs(211));
    layer0_outputs(278) <= (inputs(62)) or (inputs(28));
    layer0_outputs(279) <= not((inputs(45)) or (inputs(137)));
    layer0_outputs(280) <= not((inputs(147)) or (inputs(145)));
    layer0_outputs(281) <= inputs(183);
    layer0_outputs(282) <= (inputs(114)) or (inputs(63));
    layer0_outputs(283) <= not(inputs(91)) or (inputs(217));
    layer0_outputs(284) <= not(inputs(125)) or (inputs(50));
    layer0_outputs(285) <= not(inputs(109)) or (inputs(47));
    layer0_outputs(286) <= inputs(105);
    layer0_outputs(287) <= inputs(102);
    layer0_outputs(288) <= (inputs(113)) xor (inputs(129));
    layer0_outputs(289) <= not((inputs(161)) and (inputs(64)));
    layer0_outputs(290) <= (inputs(188)) and not (inputs(65));
    layer0_outputs(291) <= (inputs(85)) or (inputs(92));
    layer0_outputs(292) <= not((inputs(121)) or (inputs(105)));
    layer0_outputs(293) <= inputs(164);
    layer0_outputs(294) <= (inputs(187)) and not (inputs(164));
    layer0_outputs(295) <= inputs(37);
    layer0_outputs(296) <= (inputs(88)) xor (inputs(173));
    layer0_outputs(297) <= not(inputs(113));
    layer0_outputs(298) <= (inputs(242)) or (inputs(41));
    layer0_outputs(299) <= not((inputs(158)) or (inputs(145)));
    layer0_outputs(300) <= not(inputs(78));
    layer0_outputs(301) <= not(inputs(42)) or (inputs(229));
    layer0_outputs(302) <= not((inputs(19)) or (inputs(224)));
    layer0_outputs(303) <= (inputs(53)) and not (inputs(223));
    layer0_outputs(304) <= (inputs(25)) or (inputs(63));
    layer0_outputs(305) <= '0';
    layer0_outputs(306) <= not((inputs(22)) or (inputs(232)));
    layer0_outputs(307) <= not(inputs(226));
    layer0_outputs(308) <= inputs(179);
    layer0_outputs(309) <= inputs(100);
    layer0_outputs(310) <= not((inputs(45)) xor (inputs(155)));
    layer0_outputs(311) <= (inputs(245)) or (inputs(178));
    layer0_outputs(312) <= (inputs(193)) and not (inputs(95));
    layer0_outputs(313) <= inputs(55);
    layer0_outputs(314) <= not(inputs(124));
    layer0_outputs(315) <= inputs(125);
    layer0_outputs(316) <= not(inputs(195));
    layer0_outputs(317) <= (inputs(42)) or (inputs(4));
    layer0_outputs(318) <= inputs(141);
    layer0_outputs(319) <= not(inputs(83));
    layer0_outputs(320) <= not(inputs(232));
    layer0_outputs(321) <= not(inputs(146));
    layer0_outputs(322) <= not(inputs(147)) or (inputs(240));
    layer0_outputs(323) <= (inputs(140)) or (inputs(114));
    layer0_outputs(324) <= (inputs(95)) or (inputs(63));
    layer0_outputs(325) <= (inputs(191)) or (inputs(221));
    layer0_outputs(326) <= not(inputs(231)) or (inputs(6));
    layer0_outputs(327) <= not(inputs(85)) or (inputs(176));
    layer0_outputs(328) <= (inputs(121)) or (inputs(104));
    layer0_outputs(329) <= not(inputs(168));
    layer0_outputs(330) <= (inputs(45)) and not (inputs(142));
    layer0_outputs(331) <= (inputs(15)) or (inputs(17));
    layer0_outputs(332) <= not(inputs(30)) or (inputs(211));
    layer0_outputs(333) <= not(inputs(153));
    layer0_outputs(334) <= inputs(210);
    layer0_outputs(335) <= (inputs(59)) or (inputs(148));
    layer0_outputs(336) <= (inputs(223)) and not (inputs(255));
    layer0_outputs(337) <= not(inputs(84));
    layer0_outputs(338) <= not(inputs(91)) or (inputs(44));
    layer0_outputs(339) <= (inputs(133)) and not (inputs(242));
    layer0_outputs(340) <= not(inputs(228));
    layer0_outputs(341) <= not(inputs(247)) or (inputs(112));
    layer0_outputs(342) <= inputs(76);
    layer0_outputs(343) <= (inputs(76)) or (inputs(97));
    layer0_outputs(344) <= inputs(130);
    layer0_outputs(345) <= not((inputs(212)) or (inputs(227)));
    layer0_outputs(346) <= not(inputs(190)) or (inputs(82));
    layer0_outputs(347) <= inputs(141);
    layer0_outputs(348) <= not((inputs(34)) or (inputs(154)));
    layer0_outputs(349) <= (inputs(125)) or (inputs(143));
    layer0_outputs(350) <= not(inputs(41)) or (inputs(199));
    layer0_outputs(351) <= not((inputs(159)) xor (inputs(108)));
    layer0_outputs(352) <= (inputs(179)) or (inputs(97));
    layer0_outputs(353) <= (inputs(199)) and not (inputs(13));
    layer0_outputs(354) <= (inputs(197)) or (inputs(11));
    layer0_outputs(355) <= (inputs(6)) or (inputs(254));
    layer0_outputs(356) <= not(inputs(246)) or (inputs(178));
    layer0_outputs(357) <= not(inputs(236)) or (inputs(35));
    layer0_outputs(358) <= (inputs(98)) or (inputs(210));
    layer0_outputs(359) <= not((inputs(59)) or (inputs(61)));
    layer0_outputs(360) <= inputs(196);
    layer0_outputs(361) <= not(inputs(196));
    layer0_outputs(362) <= (inputs(78)) and (inputs(232));
    layer0_outputs(363) <= not((inputs(207)) xor (inputs(188)));
    layer0_outputs(364) <= not(inputs(198));
    layer0_outputs(365) <= not(inputs(185)) or (inputs(77));
    layer0_outputs(366) <= inputs(106);
    layer0_outputs(367) <= not(inputs(101)) or (inputs(206));
    layer0_outputs(368) <= (inputs(55)) and not (inputs(58));
    layer0_outputs(369) <= inputs(205);
    layer0_outputs(370) <= not(inputs(169));
    layer0_outputs(371) <= (inputs(14)) or (inputs(154));
    layer0_outputs(372) <= not(inputs(247));
    layer0_outputs(373) <= not((inputs(137)) or (inputs(77)));
    layer0_outputs(374) <= not(inputs(235)) or (inputs(114));
    layer0_outputs(375) <= inputs(164);
    layer0_outputs(376) <= not(inputs(223));
    layer0_outputs(377) <= not((inputs(125)) xor (inputs(67)));
    layer0_outputs(378) <= (inputs(66)) xor (inputs(107));
    layer0_outputs(379) <= inputs(151);
    layer0_outputs(380) <= not((inputs(72)) xor (inputs(69)));
    layer0_outputs(381) <= not((inputs(18)) or (inputs(83)));
    layer0_outputs(382) <= inputs(153);
    layer0_outputs(383) <= (inputs(71)) and not (inputs(2));
    layer0_outputs(384) <= (inputs(198)) and not (inputs(73));
    layer0_outputs(385) <= (inputs(27)) and not (inputs(158));
    layer0_outputs(386) <= not(inputs(59)) or (inputs(124));
    layer0_outputs(387) <= not((inputs(113)) or (inputs(133)));
    layer0_outputs(388) <= not(inputs(82)) or (inputs(235));
    layer0_outputs(389) <= (inputs(92)) and not (inputs(143));
    layer0_outputs(390) <= not(inputs(111));
    layer0_outputs(391) <= inputs(106);
    layer0_outputs(392) <= inputs(227);
    layer0_outputs(393) <= (inputs(134)) or (inputs(215));
    layer0_outputs(394) <= (inputs(94)) and not (inputs(126));
    layer0_outputs(395) <= not((inputs(95)) or (inputs(51)));
    layer0_outputs(396) <= not((inputs(22)) or (inputs(254)));
    layer0_outputs(397) <= not(inputs(166));
    layer0_outputs(398) <= not((inputs(251)) or (inputs(179)));
    layer0_outputs(399) <= not((inputs(95)) or (inputs(204)));
    layer0_outputs(400) <= not((inputs(82)) or (inputs(106)));
    layer0_outputs(401) <= inputs(27);
    layer0_outputs(402) <= '0';
    layer0_outputs(403) <= not(inputs(143));
    layer0_outputs(404) <= not(inputs(179));
    layer0_outputs(405) <= inputs(24);
    layer0_outputs(406) <= (inputs(171)) and not (inputs(255));
    layer0_outputs(407) <= not(inputs(193));
    layer0_outputs(408) <= (inputs(169)) and not (inputs(136));
    layer0_outputs(409) <= (inputs(174)) or (inputs(70));
    layer0_outputs(410) <= (inputs(21)) or (inputs(61));
    layer0_outputs(411) <= not((inputs(167)) or (inputs(72)));
    layer0_outputs(412) <= (inputs(168)) and (inputs(172));
    layer0_outputs(413) <= inputs(117);
    layer0_outputs(414) <= not(inputs(103));
    layer0_outputs(415) <= not(inputs(211)) or (inputs(252));
    layer0_outputs(416) <= not(inputs(126));
    layer0_outputs(417) <= not(inputs(224));
    layer0_outputs(418) <= not(inputs(231));
    layer0_outputs(419) <= (inputs(182)) or (inputs(52));
    layer0_outputs(420) <= '1';
    layer0_outputs(421) <= not(inputs(213));
    layer0_outputs(422) <= inputs(60);
    layer0_outputs(423) <= (inputs(229)) or (inputs(220));
    layer0_outputs(424) <= not((inputs(251)) xor (inputs(190)));
    layer0_outputs(425) <= inputs(217);
    layer0_outputs(426) <= (inputs(2)) xor (inputs(46));
    layer0_outputs(427) <= not(inputs(147));
    layer0_outputs(428) <= inputs(244);
    layer0_outputs(429) <= not(inputs(212)) or (inputs(81));
    layer0_outputs(430) <= not(inputs(162)) or (inputs(96));
    layer0_outputs(431) <= not(inputs(180));
    layer0_outputs(432) <= (inputs(26)) and not (inputs(1));
    layer0_outputs(433) <= inputs(78);
    layer0_outputs(434) <= not(inputs(30));
    layer0_outputs(435) <= not((inputs(20)) or (inputs(241)));
    layer0_outputs(436) <= not((inputs(176)) or (inputs(217)));
    layer0_outputs(437) <= not(inputs(221));
    layer0_outputs(438) <= not(inputs(63));
    layer0_outputs(439) <= (inputs(162)) and (inputs(150));
    layer0_outputs(440) <= inputs(120);
    layer0_outputs(441) <= (inputs(209)) or (inputs(217));
    layer0_outputs(442) <= inputs(115);
    layer0_outputs(443) <= not(inputs(150));
    layer0_outputs(444) <= not((inputs(88)) or (inputs(128)));
    layer0_outputs(445) <= (inputs(210)) or (inputs(229));
    layer0_outputs(446) <= not((inputs(187)) xor (inputs(138)));
    layer0_outputs(447) <= (inputs(199)) and not (inputs(154));
    layer0_outputs(448) <= (inputs(122)) or (inputs(182));
    layer0_outputs(449) <= (inputs(122)) xor (inputs(216));
    layer0_outputs(450) <= not(inputs(104)) or (inputs(115));
    layer0_outputs(451) <= '0';
    layer0_outputs(452) <= (inputs(187)) or (inputs(218));
    layer0_outputs(453) <= (inputs(153)) or (inputs(169));
    layer0_outputs(454) <= (inputs(205)) or (inputs(217));
    layer0_outputs(455) <= not((inputs(112)) xor (inputs(225)));
    layer0_outputs(456) <= inputs(221);
    layer0_outputs(457) <= (inputs(217)) and not (inputs(152));
    layer0_outputs(458) <= not(inputs(96));
    layer0_outputs(459) <= not((inputs(135)) or (inputs(130)));
    layer0_outputs(460) <= not((inputs(139)) or (inputs(32)));
    layer0_outputs(461) <= inputs(106);
    layer0_outputs(462) <= not(inputs(28));
    layer0_outputs(463) <= not((inputs(31)) or (inputs(96)));
    layer0_outputs(464) <= (inputs(148)) or (inputs(22));
    layer0_outputs(465) <= not(inputs(190)) or (inputs(195));
    layer0_outputs(466) <= not(inputs(246)) or (inputs(166));
    layer0_outputs(467) <= inputs(38);
    layer0_outputs(468) <= not((inputs(172)) or (inputs(115)));
    layer0_outputs(469) <= not((inputs(162)) or (inputs(128)));
    layer0_outputs(470) <= (inputs(215)) and not (inputs(40));
    layer0_outputs(471) <= (inputs(90)) xor (inputs(35));
    layer0_outputs(472) <= inputs(249);
    layer0_outputs(473) <= not(inputs(248));
    layer0_outputs(474) <= not(inputs(177));
    layer0_outputs(475) <= not(inputs(89)) or (inputs(112));
    layer0_outputs(476) <= (inputs(112)) or (inputs(65));
    layer0_outputs(477) <= not(inputs(119));
    layer0_outputs(478) <= (inputs(212)) and not (inputs(102));
    layer0_outputs(479) <= not((inputs(208)) or (inputs(218)));
    layer0_outputs(480) <= (inputs(91)) or (inputs(3));
    layer0_outputs(481) <= (inputs(135)) and (inputs(89));
    layer0_outputs(482) <= not(inputs(36));
    layer0_outputs(483) <= not(inputs(4));
    layer0_outputs(484) <= inputs(95);
    layer0_outputs(485) <= '1';
    layer0_outputs(486) <= not(inputs(62));
    layer0_outputs(487) <= not(inputs(25)) or (inputs(15));
    layer0_outputs(488) <= (inputs(35)) and not (inputs(82));
    layer0_outputs(489) <= (inputs(59)) and not (inputs(239));
    layer0_outputs(490) <= not(inputs(8));
    layer0_outputs(491) <= not((inputs(52)) xor (inputs(21)));
    layer0_outputs(492) <= not(inputs(152));
    layer0_outputs(493) <= inputs(214);
    layer0_outputs(494) <= '0';
    layer0_outputs(495) <= inputs(76);
    layer0_outputs(496) <= (inputs(66)) or (inputs(124));
    layer0_outputs(497) <= not((inputs(129)) and (inputs(66)));
    layer0_outputs(498) <= not(inputs(215));
    layer0_outputs(499) <= (inputs(11)) xor (inputs(207));
    layer0_outputs(500) <= not((inputs(237)) or (inputs(252)));
    layer0_outputs(501) <= '0';
    layer0_outputs(502) <= not((inputs(76)) or (inputs(14)));
    layer0_outputs(503) <= not(inputs(229));
    layer0_outputs(504) <= (inputs(39)) and not (inputs(232));
    layer0_outputs(505) <= (inputs(51)) or (inputs(129));
    layer0_outputs(506) <= inputs(110);
    layer0_outputs(507) <= not(inputs(100));
    layer0_outputs(508) <= not(inputs(158));
    layer0_outputs(509) <= inputs(200);
    layer0_outputs(510) <= inputs(25);
    layer0_outputs(511) <= (inputs(32)) and not (inputs(182));
    layer0_outputs(512) <= not((inputs(23)) or (inputs(187)));
    layer0_outputs(513) <= not(inputs(174));
    layer0_outputs(514) <= inputs(178);
    layer0_outputs(515) <= not((inputs(207)) xor (inputs(33)));
    layer0_outputs(516) <= inputs(142);
    layer0_outputs(517) <= not((inputs(227)) and (inputs(158)));
    layer0_outputs(518) <= (inputs(52)) or (inputs(71));
    layer0_outputs(519) <= inputs(196);
    layer0_outputs(520) <= (inputs(75)) or (inputs(94));
    layer0_outputs(521) <= (inputs(88)) or (inputs(201));
    layer0_outputs(522) <= (inputs(74)) and not (inputs(51));
    layer0_outputs(523) <= not(inputs(27));
    layer0_outputs(524) <= not((inputs(139)) or (inputs(53)));
    layer0_outputs(525) <= inputs(249);
    layer0_outputs(526) <= inputs(131);
    layer0_outputs(527) <= inputs(224);
    layer0_outputs(528) <= inputs(79);
    layer0_outputs(529) <= inputs(230);
    layer0_outputs(530) <= (inputs(171)) xor (inputs(203));
    layer0_outputs(531) <= not(inputs(78)) or (inputs(239));
    layer0_outputs(532) <= (inputs(142)) or (inputs(73));
    layer0_outputs(533) <= inputs(146);
    layer0_outputs(534) <= (inputs(24)) or (inputs(66));
    layer0_outputs(535) <= not((inputs(109)) and (inputs(176)));
    layer0_outputs(536) <= not(inputs(191));
    layer0_outputs(537) <= not((inputs(46)) or (inputs(109)));
    layer0_outputs(538) <= (inputs(50)) and (inputs(0));
    layer0_outputs(539) <= inputs(150);
    layer0_outputs(540) <= inputs(177);
    layer0_outputs(541) <= not(inputs(98));
    layer0_outputs(542) <= not(inputs(23)) or (inputs(206));
    layer0_outputs(543) <= not((inputs(184)) or (inputs(252)));
    layer0_outputs(544) <= (inputs(233)) or (inputs(194));
    layer0_outputs(545) <= not((inputs(198)) and (inputs(169)));
    layer0_outputs(546) <= (inputs(157)) xor (inputs(142));
    layer0_outputs(547) <= (inputs(42)) and not (inputs(77));
    layer0_outputs(548) <= not(inputs(57)) or (inputs(254));
    layer0_outputs(549) <= not((inputs(133)) or (inputs(77)));
    layer0_outputs(550) <= not(inputs(119));
    layer0_outputs(551) <= (inputs(229)) or (inputs(179));
    layer0_outputs(552) <= (inputs(42)) or (inputs(245));
    layer0_outputs(553) <= (inputs(128)) and not (inputs(255));
    layer0_outputs(554) <= (inputs(11)) or (inputs(39));
    layer0_outputs(555) <= not(inputs(116));
    layer0_outputs(556) <= inputs(56);
    layer0_outputs(557) <= inputs(200);
    layer0_outputs(558) <= not((inputs(125)) or (inputs(43)));
    layer0_outputs(559) <= not((inputs(15)) or (inputs(140)));
    layer0_outputs(560) <= (inputs(219)) or (inputs(190));
    layer0_outputs(561) <= (inputs(218)) and not (inputs(77));
    layer0_outputs(562) <= (inputs(49)) or (inputs(208));
    layer0_outputs(563) <= inputs(206);
    layer0_outputs(564) <= not((inputs(186)) or (inputs(185)));
    layer0_outputs(565) <= (inputs(50)) and not (inputs(159));
    layer0_outputs(566) <= not(inputs(199)) or (inputs(20));
    layer0_outputs(567) <= inputs(28);
    layer0_outputs(568) <= (inputs(139)) xor (inputs(92));
    layer0_outputs(569) <= not((inputs(234)) or (inputs(209)));
    layer0_outputs(570) <= (inputs(91)) or (inputs(66));
    layer0_outputs(571) <= not(inputs(131)) or (inputs(6));
    layer0_outputs(572) <= '0';
    layer0_outputs(573) <= not((inputs(129)) xor (inputs(210)));
    layer0_outputs(574) <= not((inputs(141)) and (inputs(147)));
    layer0_outputs(575) <= not(inputs(44)) or (inputs(192));
    layer0_outputs(576) <= (inputs(200)) or (inputs(18));
    layer0_outputs(577) <= inputs(190);
    layer0_outputs(578) <= not((inputs(100)) or (inputs(132)));
    layer0_outputs(579) <= (inputs(176)) and not (inputs(204));
    layer0_outputs(580) <= not((inputs(66)) or (inputs(59)));
    layer0_outputs(581) <= inputs(66);
    layer0_outputs(582) <= not(inputs(211)) or (inputs(167));
    layer0_outputs(583) <= not((inputs(10)) or (inputs(254)));
    layer0_outputs(584) <= (inputs(70)) and (inputs(10));
    layer0_outputs(585) <= (inputs(9)) and not (inputs(141));
    layer0_outputs(586) <= (inputs(210)) and not (inputs(191));
    layer0_outputs(587) <= inputs(212);
    layer0_outputs(588) <= not(inputs(68)) or (inputs(248));
    layer0_outputs(589) <= not(inputs(91)) or (inputs(130));
    layer0_outputs(590) <= not(inputs(219)) or (inputs(30));
    layer0_outputs(591) <= (inputs(173)) or (inputs(194));
    layer0_outputs(592) <= not((inputs(209)) xor (inputs(164)));
    layer0_outputs(593) <= not(inputs(88)) or (inputs(155));
    layer0_outputs(594) <= (inputs(86)) or (inputs(44));
    layer0_outputs(595) <= (inputs(242)) and not (inputs(226));
    layer0_outputs(596) <= not((inputs(185)) xor (inputs(106)));
    layer0_outputs(597) <= (inputs(221)) and not (inputs(173));
    layer0_outputs(598) <= not((inputs(238)) xor (inputs(47)));
    layer0_outputs(599) <= not(inputs(39));
    layer0_outputs(600) <= (inputs(67)) and not (inputs(77));
    layer0_outputs(601) <= inputs(211);
    layer0_outputs(602) <= not(inputs(183)) or (inputs(221));
    layer0_outputs(603) <= (inputs(218)) and not (inputs(37));
    layer0_outputs(604) <= inputs(40);
    layer0_outputs(605) <= not((inputs(177)) xor (inputs(172)));
    layer0_outputs(606) <= not(inputs(133));
    layer0_outputs(607) <= (inputs(79)) and not (inputs(113));
    layer0_outputs(608) <= not((inputs(243)) or (inputs(253)));
    layer0_outputs(609) <= (inputs(101)) xor (inputs(97));
    layer0_outputs(610) <= not((inputs(93)) xor (inputs(45)));
    layer0_outputs(611) <= not(inputs(228));
    layer0_outputs(612) <= (inputs(104)) or (inputs(136));
    layer0_outputs(613) <= inputs(115);
    layer0_outputs(614) <= (inputs(86)) and not (inputs(93));
    layer0_outputs(615) <= not((inputs(38)) or (inputs(18)));
    layer0_outputs(616) <= (inputs(70)) and not (inputs(236));
    layer0_outputs(617) <= not(inputs(67)) or (inputs(188));
    layer0_outputs(618) <= not(inputs(45)) or (inputs(223));
    layer0_outputs(619) <= not((inputs(208)) xor (inputs(13)));
    layer0_outputs(620) <= (inputs(55)) and not (inputs(99));
    layer0_outputs(621) <= not((inputs(230)) and (inputs(121)));
    layer0_outputs(622) <= not((inputs(236)) and (inputs(121)));
    layer0_outputs(623) <= (inputs(143)) or (inputs(212));
    layer0_outputs(624) <= not(inputs(15)) or (inputs(94));
    layer0_outputs(625) <= (inputs(147)) xor (inputs(12));
    layer0_outputs(626) <= not((inputs(195)) or (inputs(18)));
    layer0_outputs(627) <= (inputs(87)) and not (inputs(190));
    layer0_outputs(628) <= not((inputs(64)) xor (inputs(18)));
    layer0_outputs(629) <= (inputs(76)) or (inputs(42));
    layer0_outputs(630) <= not(inputs(198)) or (inputs(141));
    layer0_outputs(631) <= not(inputs(115));
    layer0_outputs(632) <= not((inputs(227)) or (inputs(82)));
    layer0_outputs(633) <= not((inputs(77)) or (inputs(176)));
    layer0_outputs(634) <= not(inputs(229));
    layer0_outputs(635) <= not(inputs(210));
    layer0_outputs(636) <= (inputs(108)) or (inputs(39));
    layer0_outputs(637) <= not(inputs(21));
    layer0_outputs(638) <= not(inputs(48));
    layer0_outputs(639) <= (inputs(128)) and (inputs(240));
    layer0_outputs(640) <= not((inputs(60)) or (inputs(83)));
    layer0_outputs(641) <= (inputs(129)) or (inputs(120));
    layer0_outputs(642) <= (inputs(99)) or (inputs(81));
    layer0_outputs(643) <= not((inputs(116)) and (inputs(179)));
    layer0_outputs(644) <= not((inputs(180)) or (inputs(191)));
    layer0_outputs(645) <= (inputs(213)) or (inputs(208));
    layer0_outputs(646) <= (inputs(90)) and not (inputs(202));
    layer0_outputs(647) <= (inputs(58)) and not (inputs(46));
    layer0_outputs(648) <= not((inputs(17)) or (inputs(121)));
    layer0_outputs(649) <= inputs(38);
    layer0_outputs(650) <= (inputs(188)) and not (inputs(51));
    layer0_outputs(651) <= not(inputs(230)) or (inputs(91));
    layer0_outputs(652) <= '1';
    layer0_outputs(653) <= (inputs(32)) or (inputs(170));
    layer0_outputs(654) <= (inputs(177)) or (inputs(35));
    layer0_outputs(655) <= inputs(238);
    layer0_outputs(656) <= (inputs(21)) and (inputs(219));
    layer0_outputs(657) <= not(inputs(144)) or (inputs(149));
    layer0_outputs(658) <= inputs(148);
    layer0_outputs(659) <= not(inputs(139)) or (inputs(176));
    layer0_outputs(660) <= (inputs(23)) xor (inputs(194));
    layer0_outputs(661) <= not((inputs(54)) or (inputs(114)));
    layer0_outputs(662) <= inputs(165);
    layer0_outputs(663) <= inputs(76);
    layer0_outputs(664) <= not((inputs(147)) xor (inputs(32)));
    layer0_outputs(665) <= not(inputs(193));
    layer0_outputs(666) <= inputs(83);
    layer0_outputs(667) <= (inputs(144)) and (inputs(142));
    layer0_outputs(668) <= not(inputs(231));
    layer0_outputs(669) <= not(inputs(252));
    layer0_outputs(670) <= not(inputs(167)) or (inputs(25));
    layer0_outputs(671) <= (inputs(222)) or (inputs(27));
    layer0_outputs(672) <= inputs(44);
    layer0_outputs(673) <= (inputs(21)) and not (inputs(13));
    layer0_outputs(674) <= not((inputs(26)) and (inputs(66)));
    layer0_outputs(675) <= not(inputs(68));
    layer0_outputs(676) <= not(inputs(158));
    layer0_outputs(677) <= not(inputs(118));
    layer0_outputs(678) <= not((inputs(217)) or (inputs(127)));
    layer0_outputs(679) <= (inputs(104)) and not (inputs(133));
    layer0_outputs(680) <= not((inputs(14)) or (inputs(242)));
    layer0_outputs(681) <= (inputs(100)) and not (inputs(16));
    layer0_outputs(682) <= (inputs(87)) xor (inputs(60));
    layer0_outputs(683) <= not((inputs(203)) or (inputs(196)));
    layer0_outputs(684) <= not((inputs(3)) or (inputs(210)));
    layer0_outputs(685) <= not((inputs(227)) or (inputs(141)));
    layer0_outputs(686) <= (inputs(95)) or (inputs(22));
    layer0_outputs(687) <= not(inputs(252));
    layer0_outputs(688) <= not((inputs(194)) or (inputs(79)));
    layer0_outputs(689) <= not((inputs(61)) and (inputs(70)));
    layer0_outputs(690) <= inputs(104);
    layer0_outputs(691) <= inputs(9);
    layer0_outputs(692) <= not(inputs(251)) or (inputs(240));
    layer0_outputs(693) <= not(inputs(163));
    layer0_outputs(694) <= not(inputs(156)) or (inputs(28));
    layer0_outputs(695) <= not(inputs(124));
    layer0_outputs(696) <= inputs(164);
    layer0_outputs(697) <= inputs(137);
    layer0_outputs(698) <= not(inputs(244)) or (inputs(78));
    layer0_outputs(699) <= inputs(213);
    layer0_outputs(700) <= not((inputs(15)) or (inputs(137)));
    layer0_outputs(701) <= (inputs(21)) xor (inputs(240));
    layer0_outputs(702) <= not(inputs(127));
    layer0_outputs(703) <= inputs(229);
    layer0_outputs(704) <= not(inputs(89));
    layer0_outputs(705) <= (inputs(164)) and not (inputs(144));
    layer0_outputs(706) <= not((inputs(135)) xor (inputs(196)));
    layer0_outputs(707) <= not((inputs(41)) or (inputs(235)));
    layer0_outputs(708) <= inputs(42);
    layer0_outputs(709) <= inputs(144);
    layer0_outputs(710) <= not(inputs(61)) or (inputs(68));
    layer0_outputs(711) <= not(inputs(108));
    layer0_outputs(712) <= (inputs(235)) and not (inputs(241));
    layer0_outputs(713) <= (inputs(228)) or (inputs(96));
    layer0_outputs(714) <= inputs(232);
    layer0_outputs(715) <= not(inputs(38)) or (inputs(94));
    layer0_outputs(716) <= (inputs(191)) and not (inputs(97));
    layer0_outputs(717) <= (inputs(225)) xor (inputs(112));
    layer0_outputs(718) <= (inputs(154)) and not (inputs(106));
    layer0_outputs(719) <= not(inputs(131)) or (inputs(79));
    layer0_outputs(720) <= not((inputs(59)) xor (inputs(255)));
    layer0_outputs(721) <= not((inputs(120)) or (inputs(63)));
    layer0_outputs(722) <= inputs(4);
    layer0_outputs(723) <= not((inputs(123)) xor (inputs(169)));
    layer0_outputs(724) <= (inputs(250)) xor (inputs(210));
    layer0_outputs(725) <= not((inputs(228)) or (inputs(3)));
    layer0_outputs(726) <= inputs(124);
    layer0_outputs(727) <= not(inputs(92));
    layer0_outputs(728) <= (inputs(181)) and (inputs(57));
    layer0_outputs(729) <= not(inputs(153));
    layer0_outputs(730) <= not(inputs(85));
    layer0_outputs(731) <= (inputs(220)) and not (inputs(81));
    layer0_outputs(732) <= not(inputs(123));
    layer0_outputs(733) <= not((inputs(164)) or (inputs(183)));
    layer0_outputs(734) <= (inputs(212)) or (inputs(244));
    layer0_outputs(735) <= not(inputs(94));
    layer0_outputs(736) <= not(inputs(143));
    layer0_outputs(737) <= (inputs(42)) or (inputs(134));
    layer0_outputs(738) <= '1';
    layer0_outputs(739) <= (inputs(111)) or (inputs(211));
    layer0_outputs(740) <= (inputs(33)) xor (inputs(137));
    layer0_outputs(741) <= (inputs(201)) and not (inputs(245));
    layer0_outputs(742) <= not(inputs(84));
    layer0_outputs(743) <= (inputs(125)) and not (inputs(250));
    layer0_outputs(744) <= (inputs(243)) xor (inputs(176));
    layer0_outputs(745) <= not(inputs(84));
    layer0_outputs(746) <= (inputs(41)) or (inputs(26));
    layer0_outputs(747) <= not((inputs(160)) xor (inputs(116)));
    layer0_outputs(748) <= not(inputs(54));
    layer0_outputs(749) <= not((inputs(20)) and (inputs(167)));
    layer0_outputs(750) <= '1';
    layer0_outputs(751) <= inputs(158);
    layer0_outputs(752) <= not((inputs(183)) and (inputs(71)));
    layer0_outputs(753) <= not((inputs(20)) or (inputs(210)));
    layer0_outputs(754) <= not(inputs(105)) or (inputs(177));
    layer0_outputs(755) <= inputs(1);
    layer0_outputs(756) <= not(inputs(161)) or (inputs(118));
    layer0_outputs(757) <= (inputs(79)) xor (inputs(107));
    layer0_outputs(758) <= (inputs(222)) and not (inputs(31));
    layer0_outputs(759) <= not(inputs(198)) or (inputs(112));
    layer0_outputs(760) <= (inputs(216)) or (inputs(157));
    layer0_outputs(761) <= inputs(36);
    layer0_outputs(762) <= (inputs(22)) and not (inputs(36));
    layer0_outputs(763) <= not((inputs(74)) or (inputs(209)));
    layer0_outputs(764) <= (inputs(27)) and not (inputs(203));
    layer0_outputs(765) <= (inputs(120)) and not (inputs(16));
    layer0_outputs(766) <= not(inputs(102)) or (inputs(111));
    layer0_outputs(767) <= (inputs(201)) or (inputs(195));
    layer0_outputs(768) <= not(inputs(178));
    layer0_outputs(769) <= (inputs(144)) xor (inputs(165));
    layer0_outputs(770) <= '0';
    layer0_outputs(771) <= inputs(182);
    layer0_outputs(772) <= not(inputs(191)) or (inputs(31));
    layer0_outputs(773) <= not(inputs(63)) or (inputs(126));
    layer0_outputs(774) <= not(inputs(125)) or (inputs(255));
    layer0_outputs(775) <= not(inputs(38)) or (inputs(130));
    layer0_outputs(776) <= (inputs(198)) and not (inputs(140));
    layer0_outputs(777) <= not((inputs(243)) xor (inputs(184)));
    layer0_outputs(778) <= not(inputs(75));
    layer0_outputs(779) <= (inputs(95)) or (inputs(11));
    layer0_outputs(780) <= not(inputs(215));
    layer0_outputs(781) <= (inputs(192)) or (inputs(251));
    layer0_outputs(782) <= not((inputs(47)) and (inputs(150)));
    layer0_outputs(783) <= (inputs(74)) and not (inputs(3));
    layer0_outputs(784) <= not(inputs(138));
    layer0_outputs(785) <= not(inputs(84));
    layer0_outputs(786) <= inputs(119);
    layer0_outputs(787) <= not((inputs(137)) or (inputs(192)));
    layer0_outputs(788) <= (inputs(193)) or (inputs(2));
    layer0_outputs(789) <= not(inputs(177));
    layer0_outputs(790) <= inputs(145);
    layer0_outputs(791) <= inputs(139);
    layer0_outputs(792) <= (inputs(58)) and not (inputs(176));
    layer0_outputs(793) <= (inputs(165)) and (inputs(231));
    layer0_outputs(794) <= not(inputs(28)) or (inputs(142));
    layer0_outputs(795) <= not(inputs(244)) or (inputs(131));
    layer0_outputs(796) <= inputs(41);
    layer0_outputs(797) <= not((inputs(173)) or (inputs(214)));
    layer0_outputs(798) <= (inputs(162)) and not (inputs(152));
    layer0_outputs(799) <= (inputs(15)) and not (inputs(224));
    layer0_outputs(800) <= not((inputs(23)) or (inputs(35)));
    layer0_outputs(801) <= not(inputs(33)) or (inputs(81));
    layer0_outputs(802) <= not((inputs(16)) or (inputs(123)));
    layer0_outputs(803) <= not(inputs(136));
    layer0_outputs(804) <= (inputs(105)) and not (inputs(164));
    layer0_outputs(805) <= not(inputs(13));
    layer0_outputs(806) <= (inputs(81)) and not (inputs(16));
    layer0_outputs(807) <= '0';
    layer0_outputs(808) <= not(inputs(232));
    layer0_outputs(809) <= (inputs(227)) or (inputs(205));
    layer0_outputs(810) <= not((inputs(3)) xor (inputs(170)));
    layer0_outputs(811) <= (inputs(245)) and not (inputs(19));
    layer0_outputs(812) <= not(inputs(138));
    layer0_outputs(813) <= not(inputs(52));
    layer0_outputs(814) <= inputs(36);
    layer0_outputs(815) <= not((inputs(7)) or (inputs(179)));
    layer0_outputs(816) <= not(inputs(99)) or (inputs(3));
    layer0_outputs(817) <= not((inputs(196)) and (inputs(230)));
    layer0_outputs(818) <= (inputs(151)) or (inputs(253));
    layer0_outputs(819) <= (inputs(194)) and (inputs(14));
    layer0_outputs(820) <= not((inputs(193)) or (inputs(125)));
    layer0_outputs(821) <= (inputs(224)) or (inputs(22));
    layer0_outputs(822) <= not(inputs(50));
    layer0_outputs(823) <= not(inputs(7)) or (inputs(178));
    layer0_outputs(824) <= not((inputs(244)) or (inputs(189)));
    layer0_outputs(825) <= not(inputs(30));
    layer0_outputs(826) <= (inputs(201)) and not (inputs(145));
    layer0_outputs(827) <= not((inputs(249)) or (inputs(63)));
    layer0_outputs(828) <= not((inputs(236)) and (inputs(200)));
    layer0_outputs(829) <= not(inputs(38));
    layer0_outputs(830) <= (inputs(114)) or (inputs(235));
    layer0_outputs(831) <= (inputs(224)) xor (inputs(117));
    layer0_outputs(832) <= not((inputs(221)) or (inputs(255)));
    layer0_outputs(833) <= inputs(173);
    layer0_outputs(834) <= not(inputs(98)) or (inputs(39));
    layer0_outputs(835) <= not(inputs(202));
    layer0_outputs(836) <= (inputs(100)) or (inputs(53));
    layer0_outputs(837) <= not((inputs(167)) and (inputs(208)));
    layer0_outputs(838) <= (inputs(67)) or (inputs(242));
    layer0_outputs(839) <= inputs(115);
    layer0_outputs(840) <= inputs(164);
    layer0_outputs(841) <= not(inputs(7)) or (inputs(13));
    layer0_outputs(842) <= inputs(86);
    layer0_outputs(843) <= '1';
    layer0_outputs(844) <= not(inputs(192));
    layer0_outputs(845) <= not((inputs(184)) or (inputs(179)));
    layer0_outputs(846) <= not(inputs(75));
    layer0_outputs(847) <= not((inputs(98)) or (inputs(113)));
    layer0_outputs(848) <= not(inputs(222));
    layer0_outputs(849) <= (inputs(248)) xor (inputs(31));
    layer0_outputs(850) <= '0';
    layer0_outputs(851) <= not(inputs(52));
    layer0_outputs(852) <= not(inputs(9));
    layer0_outputs(853) <= (inputs(4)) and not (inputs(235));
    layer0_outputs(854) <= '0';
    layer0_outputs(855) <= (inputs(106)) xor (inputs(223));
    layer0_outputs(856) <= (inputs(181)) and not (inputs(234));
    layer0_outputs(857) <= not(inputs(92));
    layer0_outputs(858) <= inputs(107);
    layer0_outputs(859) <= (inputs(182)) or (inputs(14));
    layer0_outputs(860) <= inputs(133);
    layer0_outputs(861) <= inputs(248);
    layer0_outputs(862) <= inputs(104);
    layer0_outputs(863) <= not(inputs(254));
    layer0_outputs(864) <= not(inputs(76));
    layer0_outputs(865) <= (inputs(119)) xor (inputs(179));
    layer0_outputs(866) <= inputs(123);
    layer0_outputs(867) <= not(inputs(230)) or (inputs(223));
    layer0_outputs(868) <= (inputs(80)) or (inputs(49));
    layer0_outputs(869) <= not(inputs(180)) or (inputs(255));
    layer0_outputs(870) <= not((inputs(3)) or (inputs(157)));
    layer0_outputs(871) <= not(inputs(204));
    layer0_outputs(872) <= not((inputs(30)) xor (inputs(164)));
    layer0_outputs(873) <= not(inputs(128));
    layer0_outputs(874) <= not((inputs(17)) or (inputs(59)));
    layer0_outputs(875) <= not(inputs(41));
    layer0_outputs(876) <= (inputs(178)) or (inputs(216));
    layer0_outputs(877) <= (inputs(113)) or (inputs(30));
    layer0_outputs(878) <= not(inputs(100));
    layer0_outputs(879) <= not(inputs(110));
    layer0_outputs(880) <= inputs(183);
    layer0_outputs(881) <= not(inputs(249));
    layer0_outputs(882) <= (inputs(43)) or (inputs(65));
    layer0_outputs(883) <= not((inputs(111)) and (inputs(90)));
    layer0_outputs(884) <= not(inputs(135)) or (inputs(98));
    layer0_outputs(885) <= not(inputs(143)) or (inputs(172));
    layer0_outputs(886) <= not(inputs(114));
    layer0_outputs(887) <= (inputs(207)) and not (inputs(97));
    layer0_outputs(888) <= not((inputs(207)) xor (inputs(131)));
    layer0_outputs(889) <= (inputs(218)) and not (inputs(121));
    layer0_outputs(890) <= not((inputs(193)) or (inputs(209)));
    layer0_outputs(891) <= not(inputs(234));
    layer0_outputs(892) <= inputs(180);
    layer0_outputs(893) <= inputs(6);
    layer0_outputs(894) <= not((inputs(139)) or (inputs(70)));
    layer0_outputs(895) <= (inputs(223)) and not (inputs(110));
    layer0_outputs(896) <= not((inputs(254)) or (inputs(155)));
    layer0_outputs(897) <= inputs(4);
    layer0_outputs(898) <= not((inputs(129)) xor (inputs(166)));
    layer0_outputs(899) <= not((inputs(172)) or (inputs(144)));
    layer0_outputs(900) <= not(inputs(170));
    layer0_outputs(901) <= (inputs(175)) or (inputs(174));
    layer0_outputs(902) <= not(inputs(246));
    layer0_outputs(903) <= not(inputs(88)) or (inputs(195));
    layer0_outputs(904) <= not(inputs(114));
    layer0_outputs(905) <= (inputs(227)) and not (inputs(112));
    layer0_outputs(906) <= (inputs(75)) or (inputs(92));
    layer0_outputs(907) <= inputs(174);
    layer0_outputs(908) <= inputs(213);
    layer0_outputs(909) <= (inputs(176)) or (inputs(210));
    layer0_outputs(910) <= not((inputs(137)) or (inputs(93)));
    layer0_outputs(911) <= not((inputs(185)) xor (inputs(5)));
    layer0_outputs(912) <= (inputs(197)) xor (inputs(183));
    layer0_outputs(913) <= (inputs(161)) xor (inputs(164));
    layer0_outputs(914) <= (inputs(123)) or (inputs(31));
    layer0_outputs(915) <= (inputs(142)) or (inputs(156));
    layer0_outputs(916) <= not((inputs(1)) xor (inputs(84)));
    layer0_outputs(917) <= not(inputs(230));
    layer0_outputs(918) <= not((inputs(186)) or (inputs(118)));
    layer0_outputs(919) <= not((inputs(82)) or (inputs(114)));
    layer0_outputs(920) <= inputs(38);
    layer0_outputs(921) <= not((inputs(195)) or (inputs(54)));
    layer0_outputs(922) <= not(inputs(16));
    layer0_outputs(923) <= not((inputs(12)) xor (inputs(29)));
    layer0_outputs(924) <= not(inputs(9));
    layer0_outputs(925) <= inputs(105);
    layer0_outputs(926) <= not(inputs(234)) or (inputs(68));
    layer0_outputs(927) <= (inputs(144)) or (inputs(181));
    layer0_outputs(928) <= not(inputs(166)) or (inputs(140));
    layer0_outputs(929) <= not(inputs(212));
    layer0_outputs(930) <= not((inputs(206)) xor (inputs(127)));
    layer0_outputs(931) <= (inputs(107)) or (inputs(58));
    layer0_outputs(932) <= not((inputs(3)) and (inputs(190)));
    layer0_outputs(933) <= inputs(138);
    layer0_outputs(934) <= (inputs(211)) and not (inputs(223));
    layer0_outputs(935) <= (inputs(244)) xor (inputs(203));
    layer0_outputs(936) <= not((inputs(250)) xor (inputs(112)));
    layer0_outputs(937) <= not(inputs(24));
    layer0_outputs(938) <= (inputs(192)) xor (inputs(210));
    layer0_outputs(939) <= not(inputs(196));
    layer0_outputs(940) <= not(inputs(33));
    layer0_outputs(941) <= (inputs(171)) or (inputs(5));
    layer0_outputs(942) <= not(inputs(228)) or (inputs(108));
    layer0_outputs(943) <= inputs(124);
    layer0_outputs(944) <= (inputs(253)) or (inputs(12));
    layer0_outputs(945) <= inputs(24);
    layer0_outputs(946) <= (inputs(45)) or (inputs(203));
    layer0_outputs(947) <= inputs(151);
    layer0_outputs(948) <= (inputs(51)) and not (inputs(18));
    layer0_outputs(949) <= not(inputs(164)) or (inputs(207));
    layer0_outputs(950) <= not((inputs(189)) xor (inputs(155)));
    layer0_outputs(951) <= not(inputs(49)) or (inputs(143));
    layer0_outputs(952) <= not(inputs(118));
    layer0_outputs(953) <= not((inputs(173)) xor (inputs(111)));
    layer0_outputs(954) <= inputs(76);
    layer0_outputs(955) <= (inputs(193)) or (inputs(8));
    layer0_outputs(956) <= not(inputs(145));
    layer0_outputs(957) <= not((inputs(77)) or (inputs(252)));
    layer0_outputs(958) <= inputs(117);
    layer0_outputs(959) <= (inputs(126)) and not (inputs(144));
    layer0_outputs(960) <= inputs(99);
    layer0_outputs(961) <= not((inputs(196)) or (inputs(36)));
    layer0_outputs(962) <= (inputs(220)) or (inputs(190));
    layer0_outputs(963) <= (inputs(43)) or (inputs(19));
    layer0_outputs(964) <= (inputs(187)) or (inputs(144));
    layer0_outputs(965) <= not(inputs(216));
    layer0_outputs(966) <= not((inputs(140)) xor (inputs(34)));
    layer0_outputs(967) <= not(inputs(36));
    layer0_outputs(968) <= not(inputs(174));
    layer0_outputs(969) <= not(inputs(82));
    layer0_outputs(970) <= (inputs(248)) and not (inputs(253));
    layer0_outputs(971) <= inputs(89);
    layer0_outputs(972) <= not(inputs(53));
    layer0_outputs(973) <= not(inputs(249)) or (inputs(57));
    layer0_outputs(974) <= inputs(39);
    layer0_outputs(975) <= inputs(106);
    layer0_outputs(976) <= inputs(87);
    layer0_outputs(977) <= (inputs(124)) or (inputs(101));
    layer0_outputs(978) <= (inputs(128)) or (inputs(146));
    layer0_outputs(979) <= (inputs(41)) and not (inputs(251));
    layer0_outputs(980) <= inputs(192);
    layer0_outputs(981) <= '1';
    layer0_outputs(982) <= inputs(212);
    layer0_outputs(983) <= not(inputs(11)) or (inputs(110));
    layer0_outputs(984) <= not((inputs(178)) or (inputs(214)));
    layer0_outputs(985) <= not(inputs(228));
    layer0_outputs(986) <= inputs(245);
    layer0_outputs(987) <= not((inputs(95)) or (inputs(185)));
    layer0_outputs(988) <= inputs(162);
    layer0_outputs(989) <= not(inputs(28)) or (inputs(234));
    layer0_outputs(990) <= inputs(130);
    layer0_outputs(991) <= not((inputs(145)) or (inputs(144)));
    layer0_outputs(992) <= not((inputs(109)) xor (inputs(29)));
    layer0_outputs(993) <= inputs(180);
    layer0_outputs(994) <= '1';
    layer0_outputs(995) <= not(inputs(147)) or (inputs(166));
    layer0_outputs(996) <= not((inputs(112)) or (inputs(237)));
    layer0_outputs(997) <= not((inputs(186)) or (inputs(118)));
    layer0_outputs(998) <= (inputs(26)) and not (inputs(128));
    layer0_outputs(999) <= not(inputs(45));
    layer0_outputs(1000) <= not((inputs(171)) and (inputs(184)));
    layer0_outputs(1001) <= not(inputs(149)) or (inputs(33));
    layer0_outputs(1002) <= (inputs(252)) xor (inputs(14));
    layer0_outputs(1003) <= inputs(215);
    layer0_outputs(1004) <= not(inputs(246));
    layer0_outputs(1005) <= not(inputs(123));
    layer0_outputs(1006) <= not(inputs(105)) or (inputs(163));
    layer0_outputs(1007) <= (inputs(24)) and not (inputs(18));
    layer0_outputs(1008) <= not((inputs(36)) or (inputs(202)));
    layer0_outputs(1009) <= not((inputs(209)) or (inputs(102)));
    layer0_outputs(1010) <= not(inputs(38)) or (inputs(206));
    layer0_outputs(1011) <= not((inputs(57)) or (inputs(33)));
    layer0_outputs(1012) <= (inputs(152)) xor (inputs(147));
    layer0_outputs(1013) <= inputs(130);
    layer0_outputs(1014) <= (inputs(124)) and not (inputs(37));
    layer0_outputs(1015) <= (inputs(245)) and not (inputs(126));
    layer0_outputs(1016) <= not((inputs(77)) xor (inputs(136)));
    layer0_outputs(1017) <= not(inputs(44));
    layer0_outputs(1018) <= not((inputs(192)) or (inputs(208)));
    layer0_outputs(1019) <= not(inputs(153)) or (inputs(23));
    layer0_outputs(1020) <= not((inputs(5)) or (inputs(117)));
    layer0_outputs(1021) <= (inputs(227)) and not (inputs(91));
    layer0_outputs(1022) <= (inputs(50)) or (inputs(110));
    layer0_outputs(1023) <= inputs(32);
    layer0_outputs(1024) <= inputs(109);
    layer0_outputs(1025) <= (inputs(4)) or (inputs(20));
    layer0_outputs(1026) <= inputs(66);
    layer0_outputs(1027) <= not(inputs(213));
    layer0_outputs(1028) <= not(inputs(222)) or (inputs(50));
    layer0_outputs(1029) <= inputs(129);
    layer0_outputs(1030) <= inputs(246);
    layer0_outputs(1031) <= inputs(15);
    layer0_outputs(1032) <= not(inputs(61));
    layer0_outputs(1033) <= not(inputs(60));
    layer0_outputs(1034) <= (inputs(250)) or (inputs(241));
    layer0_outputs(1035) <= not(inputs(51));
    layer0_outputs(1036) <= not((inputs(204)) or (inputs(65)));
    layer0_outputs(1037) <= not((inputs(145)) and (inputs(67)));
    layer0_outputs(1038) <= not(inputs(16));
    layer0_outputs(1039) <= (inputs(14)) and not (inputs(170));
    layer0_outputs(1040) <= (inputs(163)) and not (inputs(1));
    layer0_outputs(1041) <= not(inputs(120));
    layer0_outputs(1042) <= (inputs(236)) xor (inputs(179));
    layer0_outputs(1043) <= not(inputs(155)) or (inputs(244));
    layer0_outputs(1044) <= not((inputs(171)) or (inputs(221)));
    layer0_outputs(1045) <= not((inputs(133)) or (inputs(165)));
    layer0_outputs(1046) <= not(inputs(200)) or (inputs(85));
    layer0_outputs(1047) <= '0';
    layer0_outputs(1048) <= not((inputs(147)) or (inputs(197)));
    layer0_outputs(1049) <= (inputs(191)) or (inputs(7));
    layer0_outputs(1050) <= inputs(105);
    layer0_outputs(1051) <= (inputs(176)) or (inputs(47));
    layer0_outputs(1052) <= (inputs(228)) and not (inputs(127));
    layer0_outputs(1053) <= (inputs(39)) or (inputs(231));
    layer0_outputs(1054) <= (inputs(244)) or (inputs(77));
    layer0_outputs(1055) <= (inputs(220)) and (inputs(48));
    layer0_outputs(1056) <= inputs(115);
    layer0_outputs(1057) <= (inputs(137)) and not (inputs(210));
    layer0_outputs(1058) <= not(inputs(171));
    layer0_outputs(1059) <= (inputs(148)) xor (inputs(192));
    layer0_outputs(1060) <= inputs(130);
    layer0_outputs(1061) <= (inputs(165)) and (inputs(131));
    layer0_outputs(1062) <= (inputs(240)) or (inputs(155));
    layer0_outputs(1063) <= not(inputs(27)) or (inputs(233));
    layer0_outputs(1064) <= inputs(93);
    layer0_outputs(1065) <= (inputs(183)) xor (inputs(47));
    layer0_outputs(1066) <= (inputs(91)) or (inputs(173));
    layer0_outputs(1067) <= not((inputs(119)) or (inputs(135)));
    layer0_outputs(1068) <= inputs(163);
    layer0_outputs(1069) <= not(inputs(96)) or (inputs(139));
    layer0_outputs(1070) <= not((inputs(206)) or (inputs(241)));
    layer0_outputs(1071) <= (inputs(186)) and not (inputs(197));
    layer0_outputs(1072) <= (inputs(19)) and not (inputs(208));
    layer0_outputs(1073) <= not(inputs(130));
    layer0_outputs(1074) <= not(inputs(195)) or (inputs(113));
    layer0_outputs(1075) <= not((inputs(243)) or (inputs(45)));
    layer0_outputs(1076) <= inputs(182);
    layer0_outputs(1077) <= (inputs(248)) or (inputs(98));
    layer0_outputs(1078) <= not(inputs(116));
    layer0_outputs(1079) <= not((inputs(44)) or (inputs(7)));
    layer0_outputs(1080) <= (inputs(88)) and not (inputs(16));
    layer0_outputs(1081) <= not((inputs(70)) or (inputs(6)));
    layer0_outputs(1082) <= not(inputs(81));
    layer0_outputs(1083) <= not(inputs(132));
    layer0_outputs(1084) <= (inputs(134)) or (inputs(101));
    layer0_outputs(1085) <= (inputs(250)) and not (inputs(201));
    layer0_outputs(1086) <= inputs(216);
    layer0_outputs(1087) <= not(inputs(157));
    layer0_outputs(1088) <= (inputs(80)) xor (inputs(39));
    layer0_outputs(1089) <= (inputs(78)) and not (inputs(173));
    layer0_outputs(1090) <= '1';
    layer0_outputs(1091) <= not(inputs(25));
    layer0_outputs(1092) <= not((inputs(191)) or (inputs(32)));
    layer0_outputs(1093) <= not((inputs(29)) or (inputs(110)));
    layer0_outputs(1094) <= inputs(185);
    layer0_outputs(1095) <= (inputs(91)) and not (inputs(212));
    layer0_outputs(1096) <= (inputs(134)) xor (inputs(151));
    layer0_outputs(1097) <= inputs(235);
    layer0_outputs(1098) <= not(inputs(197)) or (inputs(98));
    layer0_outputs(1099) <= not(inputs(210)) or (inputs(95));
    layer0_outputs(1100) <= not((inputs(79)) and (inputs(239)));
    layer0_outputs(1101) <= not(inputs(108));
    layer0_outputs(1102) <= not(inputs(62));
    layer0_outputs(1103) <= not(inputs(8)) or (inputs(15));
    layer0_outputs(1104) <= inputs(102);
    layer0_outputs(1105) <= (inputs(35)) or (inputs(194));
    layer0_outputs(1106) <= not(inputs(134));
    layer0_outputs(1107) <= (inputs(19)) or (inputs(102));
    layer0_outputs(1108) <= (inputs(6)) and not (inputs(191));
    layer0_outputs(1109) <= not(inputs(62)) or (inputs(239));
    layer0_outputs(1110) <= inputs(178);
    layer0_outputs(1111) <= not(inputs(177));
    layer0_outputs(1112) <= (inputs(160)) and not (inputs(46));
    layer0_outputs(1113) <= inputs(93);
    layer0_outputs(1114) <= (inputs(219)) and not (inputs(248));
    layer0_outputs(1115) <= not((inputs(159)) xor (inputs(238)));
    layer0_outputs(1116) <= (inputs(177)) and (inputs(177));
    layer0_outputs(1117) <= (inputs(195)) or (inputs(6));
    layer0_outputs(1118) <= not(inputs(87));
    layer0_outputs(1119) <= (inputs(154)) and (inputs(166));
    layer0_outputs(1120) <= not(inputs(17)) or (inputs(157));
    layer0_outputs(1121) <= not(inputs(11));
    layer0_outputs(1122) <= not((inputs(124)) or (inputs(123)));
    layer0_outputs(1123) <= not(inputs(175));
    layer0_outputs(1124) <= not(inputs(99));
    layer0_outputs(1125) <= (inputs(80)) xor (inputs(18));
    layer0_outputs(1126) <= (inputs(73)) or (inputs(223));
    layer0_outputs(1127) <= not((inputs(75)) xor (inputs(32)));
    layer0_outputs(1128) <= not(inputs(245));
    layer0_outputs(1129) <= inputs(133);
    layer0_outputs(1130) <= inputs(168);
    layer0_outputs(1131) <= not(inputs(102));
    layer0_outputs(1132) <= (inputs(198)) and (inputs(197));
    layer0_outputs(1133) <= not(inputs(227)) or (inputs(238));
    layer0_outputs(1134) <= (inputs(32)) and not (inputs(64));
    layer0_outputs(1135) <= inputs(82);
    layer0_outputs(1136) <= not(inputs(103)) or (inputs(189));
    layer0_outputs(1137) <= not(inputs(55)) or (inputs(1));
    layer0_outputs(1138) <= not(inputs(60)) or (inputs(107));
    layer0_outputs(1139) <= not((inputs(225)) xor (inputs(200)));
    layer0_outputs(1140) <= not(inputs(105)) or (inputs(22));
    layer0_outputs(1141) <= (inputs(78)) or (inputs(43));
    layer0_outputs(1142) <= not(inputs(54));
    layer0_outputs(1143) <= (inputs(148)) or (inputs(115));
    layer0_outputs(1144) <= not((inputs(156)) or (inputs(140)));
    layer0_outputs(1145) <= not(inputs(158));
    layer0_outputs(1146) <= (inputs(124)) xor (inputs(235));
    layer0_outputs(1147) <= (inputs(248)) xor (inputs(224));
    layer0_outputs(1148) <= not(inputs(248));
    layer0_outputs(1149) <= not((inputs(24)) or (inputs(97)));
    layer0_outputs(1150) <= (inputs(7)) or (inputs(191));
    layer0_outputs(1151) <= inputs(25);
    layer0_outputs(1152) <= not(inputs(48));
    layer0_outputs(1153) <= not(inputs(218));
    layer0_outputs(1154) <= (inputs(76)) and not (inputs(64));
    layer0_outputs(1155) <= not((inputs(89)) or (inputs(152)));
    layer0_outputs(1156) <= not((inputs(152)) or (inputs(67)));
    layer0_outputs(1157) <= inputs(212);
    layer0_outputs(1158) <= not((inputs(199)) and (inputs(57)));
    layer0_outputs(1159) <= (inputs(251)) and (inputs(159));
    layer0_outputs(1160) <= not(inputs(102)) or (inputs(0));
    layer0_outputs(1161) <= not(inputs(136)) or (inputs(25));
    layer0_outputs(1162) <= (inputs(111)) xor (inputs(238));
    layer0_outputs(1163) <= (inputs(224)) or (inputs(196));
    layer0_outputs(1164) <= not(inputs(229));
    layer0_outputs(1165) <= not((inputs(241)) xor (inputs(118)));
    layer0_outputs(1166) <= inputs(146);
    layer0_outputs(1167) <= inputs(88);
    layer0_outputs(1168) <= (inputs(186)) and (inputs(134));
    layer0_outputs(1169) <= inputs(67);
    layer0_outputs(1170) <= not((inputs(82)) or (inputs(52)));
    layer0_outputs(1171) <= not(inputs(56));
    layer0_outputs(1172) <= not((inputs(71)) xor (inputs(102)));
    layer0_outputs(1173) <= inputs(130);
    layer0_outputs(1174) <= inputs(41);
    layer0_outputs(1175) <= (inputs(161)) and not (inputs(166));
    layer0_outputs(1176) <= (inputs(50)) or (inputs(114));
    layer0_outputs(1177) <= inputs(69);
    layer0_outputs(1178) <= not((inputs(34)) xor (inputs(55)));
    layer0_outputs(1179) <= (inputs(228)) or (inputs(181));
    layer0_outputs(1180) <= not(inputs(22));
    layer0_outputs(1181) <= (inputs(56)) and not (inputs(80));
    layer0_outputs(1182) <= (inputs(27)) and not (inputs(149));
    layer0_outputs(1183) <= inputs(87);
    layer0_outputs(1184) <= not((inputs(4)) and (inputs(213)));
    layer0_outputs(1185) <= not(inputs(107)) or (inputs(74));
    layer0_outputs(1186) <= not(inputs(151));
    layer0_outputs(1187) <= (inputs(240)) and (inputs(169));
    layer0_outputs(1188) <= (inputs(2)) or (inputs(209));
    layer0_outputs(1189) <= inputs(149);
    layer0_outputs(1190) <= inputs(165);
    layer0_outputs(1191) <= inputs(164);
    layer0_outputs(1192) <= not(inputs(19));
    layer0_outputs(1193) <= inputs(164);
    layer0_outputs(1194) <= (inputs(2)) or (inputs(123));
    layer0_outputs(1195) <= not(inputs(55)) or (inputs(252));
    layer0_outputs(1196) <= not((inputs(85)) or (inputs(143)));
    layer0_outputs(1197) <= not(inputs(215));
    layer0_outputs(1198) <= (inputs(228)) xor (inputs(56));
    layer0_outputs(1199) <= (inputs(139)) xor (inputs(166));
    layer0_outputs(1200) <= (inputs(71)) and (inputs(231));
    layer0_outputs(1201) <= inputs(170);
    layer0_outputs(1202) <= not(inputs(189)) or (inputs(2));
    layer0_outputs(1203) <= (inputs(161)) and not (inputs(146));
    layer0_outputs(1204) <= not(inputs(129));
    layer0_outputs(1205) <= not((inputs(210)) or (inputs(70)));
    layer0_outputs(1206) <= inputs(28);
    layer0_outputs(1207) <= not((inputs(1)) or (inputs(5)));
    layer0_outputs(1208) <= not(inputs(119)) or (inputs(125));
    layer0_outputs(1209) <= (inputs(174)) xor (inputs(206));
    layer0_outputs(1210) <= (inputs(111)) or (inputs(84));
    layer0_outputs(1211) <= not(inputs(83));
    layer0_outputs(1212) <= inputs(176);
    layer0_outputs(1213) <= not((inputs(107)) and (inputs(147)));
    layer0_outputs(1214) <= (inputs(236)) xor (inputs(123));
    layer0_outputs(1215) <= inputs(146);
    layer0_outputs(1216) <= not((inputs(51)) or (inputs(148)));
    layer0_outputs(1217) <= (inputs(138)) or (inputs(111));
    layer0_outputs(1218) <= (inputs(248)) or (inputs(3));
    layer0_outputs(1219) <= not((inputs(142)) and (inputs(13)));
    layer0_outputs(1220) <= not(inputs(235));
    layer0_outputs(1221) <= inputs(182);
    layer0_outputs(1222) <= not(inputs(149));
    layer0_outputs(1223) <= not((inputs(75)) or (inputs(82)));
    layer0_outputs(1224) <= inputs(231);
    layer0_outputs(1225) <= inputs(36);
    layer0_outputs(1226) <= not(inputs(228));
    layer0_outputs(1227) <= (inputs(33)) and (inputs(127));
    layer0_outputs(1228) <= not(inputs(224)) or (inputs(167));
    layer0_outputs(1229) <= not((inputs(144)) or (inputs(161)));
    layer0_outputs(1230) <= not(inputs(213));
    layer0_outputs(1231) <= inputs(165);
    layer0_outputs(1232) <= inputs(103);
    layer0_outputs(1233) <= not(inputs(129));
    layer0_outputs(1234) <= not(inputs(88));
    layer0_outputs(1235) <= (inputs(175)) and not (inputs(12));
    layer0_outputs(1236) <= (inputs(18)) xor (inputs(80));
    layer0_outputs(1237) <= not((inputs(249)) xor (inputs(235)));
    layer0_outputs(1238) <= (inputs(23)) and not (inputs(144));
    layer0_outputs(1239) <= not((inputs(188)) xor (inputs(234)));
    layer0_outputs(1240) <= not(inputs(88)) or (inputs(113));
    layer0_outputs(1241) <= inputs(100);
    layer0_outputs(1242) <= not(inputs(37));
    layer0_outputs(1243) <= not((inputs(126)) or (inputs(20)));
    layer0_outputs(1244) <= not(inputs(199)) or (inputs(134));
    layer0_outputs(1245) <= inputs(109);
    layer0_outputs(1246) <= not(inputs(227)) or (inputs(39));
    layer0_outputs(1247) <= (inputs(223)) or (inputs(221));
    layer0_outputs(1248) <= (inputs(94)) or (inputs(77));
    layer0_outputs(1249) <= (inputs(181)) or (inputs(163));
    layer0_outputs(1250) <= not((inputs(181)) or (inputs(48)));
    layer0_outputs(1251) <= not(inputs(238)) or (inputs(58));
    layer0_outputs(1252) <= inputs(228);
    layer0_outputs(1253) <= not((inputs(138)) and (inputs(244)));
    layer0_outputs(1254) <= (inputs(36)) and not (inputs(247));
    layer0_outputs(1255) <= (inputs(138)) and not (inputs(1));
    layer0_outputs(1256) <= not((inputs(210)) or (inputs(164)));
    layer0_outputs(1257) <= not((inputs(202)) xor (inputs(200)));
    layer0_outputs(1258) <= (inputs(14)) or (inputs(18));
    layer0_outputs(1259) <= not((inputs(54)) and (inputs(2)));
    layer0_outputs(1260) <= (inputs(74)) and not (inputs(209));
    layer0_outputs(1261) <= inputs(156);
    layer0_outputs(1262) <= (inputs(216)) or (inputs(117));
    layer0_outputs(1263) <= not(inputs(135));
    layer0_outputs(1264) <= not((inputs(174)) or (inputs(104)));
    layer0_outputs(1265) <= not((inputs(57)) or (inputs(30)));
    layer0_outputs(1266) <= not((inputs(53)) and (inputs(60)));
    layer0_outputs(1267) <= not((inputs(36)) or (inputs(163)));
    layer0_outputs(1268) <= not((inputs(206)) or (inputs(17)));
    layer0_outputs(1269) <= inputs(110);
    layer0_outputs(1270) <= not(inputs(119));
    layer0_outputs(1271) <= not((inputs(228)) or (inputs(218)));
    layer0_outputs(1272) <= inputs(168);
    layer0_outputs(1273) <= (inputs(232)) and (inputs(198));
    layer0_outputs(1274) <= '0';
    layer0_outputs(1275) <= (inputs(148)) or (inputs(1));
    layer0_outputs(1276) <= not((inputs(224)) or (inputs(63)));
    layer0_outputs(1277) <= not(inputs(74)) or (inputs(198));
    layer0_outputs(1278) <= not(inputs(61)) or (inputs(237));
    layer0_outputs(1279) <= inputs(45);
    layer0_outputs(1280) <= (inputs(242)) and not (inputs(159));
    layer0_outputs(1281) <= not(inputs(72)) or (inputs(64));
    layer0_outputs(1282) <= not(inputs(63));
    layer0_outputs(1283) <= not(inputs(254));
    layer0_outputs(1284) <= not(inputs(52));
    layer0_outputs(1285) <= inputs(106);
    layer0_outputs(1286) <= not((inputs(87)) or (inputs(176)));
    layer0_outputs(1287) <= (inputs(214)) and not (inputs(223));
    layer0_outputs(1288) <= not((inputs(182)) xor (inputs(170)));
    layer0_outputs(1289) <= not(inputs(1));
    layer0_outputs(1290) <= not(inputs(25)) or (inputs(241));
    layer0_outputs(1291) <= (inputs(5)) xor (inputs(10));
    layer0_outputs(1292) <= inputs(106);
    layer0_outputs(1293) <= not(inputs(36)) or (inputs(114));
    layer0_outputs(1294) <= not(inputs(37));
    layer0_outputs(1295) <= not(inputs(108));
    layer0_outputs(1296) <= inputs(220);
    layer0_outputs(1297) <= (inputs(38)) and not (inputs(17));
    layer0_outputs(1298) <= not((inputs(67)) or (inputs(80)));
    layer0_outputs(1299) <= inputs(147);
    layer0_outputs(1300) <= inputs(76);
    layer0_outputs(1301) <= (inputs(106)) xor (inputs(237));
    layer0_outputs(1302) <= (inputs(15)) xor (inputs(149));
    layer0_outputs(1303) <= '1';
    layer0_outputs(1304) <= (inputs(90)) and (inputs(204));
    layer0_outputs(1305) <= not(inputs(101)) or (inputs(6));
    layer0_outputs(1306) <= (inputs(98)) and not (inputs(67));
    layer0_outputs(1307) <= not(inputs(203)) or (inputs(81));
    layer0_outputs(1308) <= (inputs(78)) xor (inputs(76));
    layer0_outputs(1309) <= inputs(90);
    layer0_outputs(1310) <= not(inputs(135));
    layer0_outputs(1311) <= (inputs(195)) or (inputs(253));
    layer0_outputs(1312) <= (inputs(196)) xor (inputs(169));
    layer0_outputs(1313) <= not((inputs(24)) and (inputs(195)));
    layer0_outputs(1314) <= inputs(72);
    layer0_outputs(1315) <= not(inputs(160)) or (inputs(254));
    layer0_outputs(1316) <= inputs(197);
    layer0_outputs(1317) <= inputs(46);
    layer0_outputs(1318) <= not((inputs(143)) or (inputs(109)));
    layer0_outputs(1319) <= inputs(168);
    layer0_outputs(1320) <= not(inputs(25)) or (inputs(205));
    layer0_outputs(1321) <= not(inputs(25));
    layer0_outputs(1322) <= not((inputs(71)) and (inputs(149)));
    layer0_outputs(1323) <= inputs(101);
    layer0_outputs(1324) <= not((inputs(252)) or (inputs(84)));
    layer0_outputs(1325) <= not(inputs(23));
    layer0_outputs(1326) <= not(inputs(198));
    layer0_outputs(1327) <= not((inputs(184)) xor (inputs(233)));
    layer0_outputs(1328) <= not((inputs(37)) or (inputs(95)));
    layer0_outputs(1329) <= not(inputs(92)) or (inputs(175));
    layer0_outputs(1330) <= (inputs(218)) or (inputs(238));
    layer0_outputs(1331) <= not((inputs(141)) xor (inputs(121)));
    layer0_outputs(1332) <= not((inputs(57)) and (inputs(91)));
    layer0_outputs(1333) <= (inputs(115)) and not (inputs(154));
    layer0_outputs(1334) <= not(inputs(100));
    layer0_outputs(1335) <= inputs(25);
    layer0_outputs(1336) <= inputs(146);
    layer0_outputs(1337) <= not((inputs(102)) or (inputs(13)));
    layer0_outputs(1338) <= not((inputs(17)) and (inputs(199)));
    layer0_outputs(1339) <= (inputs(140)) or (inputs(13));
    layer0_outputs(1340) <= (inputs(119)) and not (inputs(14));
    layer0_outputs(1341) <= (inputs(105)) and not (inputs(145));
    layer0_outputs(1342) <= not((inputs(222)) or (inputs(158)));
    layer0_outputs(1343) <= (inputs(238)) xor (inputs(94));
    layer0_outputs(1344) <= (inputs(26)) or (inputs(241));
    layer0_outputs(1345) <= (inputs(14)) and not (inputs(188));
    layer0_outputs(1346) <= not(inputs(195));
    layer0_outputs(1347) <= inputs(222);
    layer0_outputs(1348) <= inputs(186);
    layer0_outputs(1349) <= inputs(237);
    layer0_outputs(1350) <= (inputs(39)) and not (inputs(255));
    layer0_outputs(1351) <= not(inputs(111));
    layer0_outputs(1352) <= inputs(48);
    layer0_outputs(1353) <= not(inputs(45));
    layer0_outputs(1354) <= inputs(162);
    layer0_outputs(1355) <= not(inputs(122)) or (inputs(48));
    layer0_outputs(1356) <= not((inputs(100)) or (inputs(183)));
    layer0_outputs(1357) <= not((inputs(126)) or (inputs(144)));
    layer0_outputs(1358) <= (inputs(107)) xor (inputs(156));
    layer0_outputs(1359) <= (inputs(192)) xor (inputs(9));
    layer0_outputs(1360) <= not(inputs(156));
    layer0_outputs(1361) <= not((inputs(64)) xor (inputs(150)));
    layer0_outputs(1362) <= not(inputs(117));
    layer0_outputs(1363) <= '0';
    layer0_outputs(1364) <= not(inputs(167));
    layer0_outputs(1365) <= inputs(132);
    layer0_outputs(1366) <= (inputs(217)) and not (inputs(5));
    layer0_outputs(1367) <= not((inputs(231)) and (inputs(58)));
    layer0_outputs(1368) <= (inputs(217)) or (inputs(31));
    layer0_outputs(1369) <= not((inputs(97)) or (inputs(10)));
    layer0_outputs(1370) <= not((inputs(239)) or (inputs(238)));
    layer0_outputs(1371) <= inputs(188);
    layer0_outputs(1372) <= (inputs(65)) and (inputs(32));
    layer0_outputs(1373) <= not(inputs(56));
    layer0_outputs(1374) <= not(inputs(158));
    layer0_outputs(1375) <= inputs(110);
    layer0_outputs(1376) <= inputs(66);
    layer0_outputs(1377) <= not(inputs(119)) or (inputs(19));
    layer0_outputs(1378) <= inputs(135);
    layer0_outputs(1379) <= not((inputs(41)) xor (inputs(57)));
    layer0_outputs(1380) <= (inputs(62)) or (inputs(224));
    layer0_outputs(1381) <= not((inputs(249)) xor (inputs(201)));
    layer0_outputs(1382) <= (inputs(160)) or (inputs(243));
    layer0_outputs(1383) <= (inputs(161)) or (inputs(51));
    layer0_outputs(1384) <= (inputs(87)) and not (inputs(193));
    layer0_outputs(1385) <= not(inputs(109)) or (inputs(128));
    layer0_outputs(1386) <= inputs(226);
    layer0_outputs(1387) <= not(inputs(111)) or (inputs(31));
    layer0_outputs(1388) <= inputs(43);
    layer0_outputs(1389) <= (inputs(168)) and not (inputs(112));
    layer0_outputs(1390) <= not(inputs(147)) or (inputs(188));
    layer0_outputs(1391) <= not(inputs(115));
    layer0_outputs(1392) <= not(inputs(197));
    layer0_outputs(1393) <= not((inputs(68)) or (inputs(53)));
    layer0_outputs(1394) <= (inputs(165)) or (inputs(213));
    layer0_outputs(1395) <= '0';
    layer0_outputs(1396) <= (inputs(37)) or (inputs(223));
    layer0_outputs(1397) <= '1';
    layer0_outputs(1398) <= not((inputs(142)) or (inputs(203)));
    layer0_outputs(1399) <= inputs(112);
    layer0_outputs(1400) <= not(inputs(75)) or (inputs(252));
    layer0_outputs(1401) <= not(inputs(26)) or (inputs(142));
    layer0_outputs(1402) <= not((inputs(243)) xor (inputs(117)));
    layer0_outputs(1403) <= (inputs(69)) or (inputs(233));
    layer0_outputs(1404) <= inputs(93);
    layer0_outputs(1405) <= (inputs(72)) and not (inputs(15));
    layer0_outputs(1406) <= not(inputs(201)) or (inputs(193));
    layer0_outputs(1407) <= not(inputs(138));
    layer0_outputs(1408) <= inputs(25);
    layer0_outputs(1409) <= not(inputs(139)) or (inputs(72));
    layer0_outputs(1410) <= not(inputs(222)) or (inputs(30));
    layer0_outputs(1411) <= not(inputs(109));
    layer0_outputs(1412) <= (inputs(201)) or (inputs(139));
    layer0_outputs(1413) <= (inputs(122)) and not (inputs(169));
    layer0_outputs(1414) <= (inputs(20)) and not (inputs(184));
    layer0_outputs(1415) <= (inputs(62)) and (inputs(241));
    layer0_outputs(1416) <= inputs(193);
    layer0_outputs(1417) <= not(inputs(76));
    layer0_outputs(1418) <= inputs(118);
    layer0_outputs(1419) <= inputs(235);
    layer0_outputs(1420) <= (inputs(132)) or (inputs(234));
    layer0_outputs(1421) <= (inputs(229)) and not (inputs(94));
    layer0_outputs(1422) <= inputs(46);
    layer0_outputs(1423) <= (inputs(202)) and not (inputs(61));
    layer0_outputs(1424) <= not((inputs(79)) xor (inputs(255)));
    layer0_outputs(1425) <= not(inputs(66));
    layer0_outputs(1426) <= not(inputs(180));
    layer0_outputs(1427) <= (inputs(119)) and not (inputs(114));
    layer0_outputs(1428) <= not(inputs(247)) or (inputs(153));
    layer0_outputs(1429) <= (inputs(150)) and not (inputs(73));
    layer0_outputs(1430) <= not((inputs(216)) or (inputs(176)));
    layer0_outputs(1431) <= inputs(192);
    layer0_outputs(1432) <= not((inputs(4)) and (inputs(41)));
    layer0_outputs(1433) <= (inputs(116)) or (inputs(88));
    layer0_outputs(1434) <= (inputs(123)) and not (inputs(113));
    layer0_outputs(1435) <= '1';
    layer0_outputs(1436) <= (inputs(74)) or (inputs(6));
    layer0_outputs(1437) <= not(inputs(249));
    layer0_outputs(1438) <= '0';
    layer0_outputs(1439) <= not(inputs(81));
    layer0_outputs(1440) <= (inputs(184)) or (inputs(253));
    layer0_outputs(1441) <= not((inputs(159)) or (inputs(255)));
    layer0_outputs(1442) <= not((inputs(156)) xor (inputs(47)));
    layer0_outputs(1443) <= (inputs(221)) or (inputs(57));
    layer0_outputs(1444) <= inputs(130);
    layer0_outputs(1445) <= (inputs(74)) and not (inputs(117));
    layer0_outputs(1446) <= not(inputs(181));
    layer0_outputs(1447) <= not(inputs(123));
    layer0_outputs(1448) <= not((inputs(115)) or (inputs(144)));
    layer0_outputs(1449) <= (inputs(14)) and not (inputs(208));
    layer0_outputs(1450) <= (inputs(77)) and not (inputs(236));
    layer0_outputs(1451) <= inputs(113);
    layer0_outputs(1452) <= (inputs(165)) or (inputs(17));
    layer0_outputs(1453) <= not(inputs(41));
    layer0_outputs(1454) <= '0';
    layer0_outputs(1455) <= not((inputs(145)) or (inputs(168)));
    layer0_outputs(1456) <= inputs(85);
    layer0_outputs(1457) <= not(inputs(0)) or (inputs(92));
    layer0_outputs(1458) <= not(inputs(104));
    layer0_outputs(1459) <= inputs(9);
    layer0_outputs(1460) <= not((inputs(232)) and (inputs(59)));
    layer0_outputs(1461) <= not(inputs(42));
    layer0_outputs(1462) <= not(inputs(72));
    layer0_outputs(1463) <= not((inputs(96)) xor (inputs(207)));
    layer0_outputs(1464) <= not(inputs(178));
    layer0_outputs(1465) <= (inputs(53)) xor (inputs(3));
    layer0_outputs(1466) <= not((inputs(78)) or (inputs(67)));
    layer0_outputs(1467) <= (inputs(210)) and not (inputs(84));
    layer0_outputs(1468) <= not(inputs(20));
    layer0_outputs(1469) <= not(inputs(254)) or (inputs(82));
    layer0_outputs(1470) <= not((inputs(101)) or (inputs(212)));
    layer0_outputs(1471) <= (inputs(165)) and (inputs(165));
    layer0_outputs(1472) <= inputs(184);
    layer0_outputs(1473) <= not((inputs(247)) or (inputs(231)));
    layer0_outputs(1474) <= not((inputs(141)) or (inputs(124)));
    layer0_outputs(1475) <= not(inputs(141)) or (inputs(31));
    layer0_outputs(1476) <= (inputs(154)) xor (inputs(124));
    layer0_outputs(1477) <= not(inputs(126)) or (inputs(44));
    layer0_outputs(1478) <= not(inputs(41));
    layer0_outputs(1479) <= inputs(47);
    layer0_outputs(1480) <= (inputs(139)) and (inputs(60));
    layer0_outputs(1481) <= (inputs(195)) or (inputs(207));
    layer0_outputs(1482) <= '0';
    layer0_outputs(1483) <= (inputs(108)) and not (inputs(97));
    layer0_outputs(1484) <= inputs(82);
    layer0_outputs(1485) <= not((inputs(183)) xor (inputs(69)));
    layer0_outputs(1486) <= not((inputs(92)) xor (inputs(74)));
    layer0_outputs(1487) <= not((inputs(36)) or (inputs(237)));
    layer0_outputs(1488) <= inputs(141);
    layer0_outputs(1489) <= (inputs(163)) or (inputs(239));
    layer0_outputs(1490) <= (inputs(151)) and not (inputs(192));
    layer0_outputs(1491) <= not(inputs(165));
    layer0_outputs(1492) <= (inputs(74)) and not (inputs(171));
    layer0_outputs(1493) <= inputs(98);
    layer0_outputs(1494) <= not((inputs(118)) or (inputs(205)));
    layer0_outputs(1495) <= not(inputs(60)) or (inputs(139));
    layer0_outputs(1496) <= inputs(247);
    layer0_outputs(1497) <= not(inputs(14)) or (inputs(59));
    layer0_outputs(1498) <= (inputs(245)) and not (inputs(95));
    layer0_outputs(1499) <= not(inputs(10));
    layer0_outputs(1500) <= not(inputs(123)) or (inputs(10));
    layer0_outputs(1501) <= inputs(228);
    layer0_outputs(1502) <= inputs(38);
    layer0_outputs(1503) <= not((inputs(190)) or (inputs(240)));
    layer0_outputs(1504) <= (inputs(23)) xor (inputs(109));
    layer0_outputs(1505) <= not(inputs(43)) or (inputs(88));
    layer0_outputs(1506) <= (inputs(188)) or (inputs(194));
    layer0_outputs(1507) <= '1';
    layer0_outputs(1508) <= not((inputs(221)) or (inputs(170)));
    layer0_outputs(1509) <= inputs(119);
    layer0_outputs(1510) <= not(inputs(159));
    layer0_outputs(1511) <= '1';
    layer0_outputs(1512) <= not((inputs(4)) or (inputs(63)));
    layer0_outputs(1513) <= (inputs(73)) xor (inputs(37));
    layer0_outputs(1514) <= not(inputs(54)) or (inputs(17));
    layer0_outputs(1515) <= (inputs(64)) or (inputs(24));
    layer0_outputs(1516) <= not((inputs(1)) xor (inputs(238)));
    layer0_outputs(1517) <= inputs(89);
    layer0_outputs(1518) <= inputs(246);
    layer0_outputs(1519) <= not((inputs(135)) xor (inputs(16)));
    layer0_outputs(1520) <= not(inputs(108));
    layer0_outputs(1521) <= inputs(134);
    layer0_outputs(1522) <= not(inputs(177)) or (inputs(226));
    layer0_outputs(1523) <= not(inputs(172));
    layer0_outputs(1524) <= not(inputs(204)) or (inputs(110));
    layer0_outputs(1525) <= inputs(30);
    layer0_outputs(1526) <= not(inputs(44));
    layer0_outputs(1527) <= not(inputs(127)) or (inputs(203));
    layer0_outputs(1528) <= not(inputs(249));
    layer0_outputs(1529) <= (inputs(131)) or (inputs(192));
    layer0_outputs(1530) <= not((inputs(34)) or (inputs(209)));
    layer0_outputs(1531) <= (inputs(122)) and not (inputs(213));
    layer0_outputs(1532) <= not(inputs(88));
    layer0_outputs(1533) <= (inputs(118)) or (inputs(37));
    layer0_outputs(1534) <= (inputs(122)) or (inputs(104));
    layer0_outputs(1535) <= not(inputs(166)) or (inputs(125));
    layer0_outputs(1536) <= (inputs(125)) and not (inputs(110));
    layer0_outputs(1537) <= not(inputs(179));
    layer0_outputs(1538) <= not(inputs(8));
    layer0_outputs(1539) <= '1';
    layer0_outputs(1540) <= (inputs(247)) and not (inputs(75));
    layer0_outputs(1541) <= (inputs(118)) and not (inputs(0));
    layer0_outputs(1542) <= not(inputs(169));
    layer0_outputs(1543) <= not((inputs(30)) or (inputs(154)));
    layer0_outputs(1544) <= inputs(214);
    layer0_outputs(1545) <= inputs(120);
    layer0_outputs(1546) <= not((inputs(145)) or (inputs(99)));
    layer0_outputs(1547) <= inputs(169);
    layer0_outputs(1548) <= not((inputs(199)) and (inputs(122)));
    layer0_outputs(1549) <= inputs(30);
    layer0_outputs(1550) <= (inputs(119)) or (inputs(172));
    layer0_outputs(1551) <= not(inputs(83));
    layer0_outputs(1552) <= (inputs(79)) or (inputs(69));
    layer0_outputs(1553) <= (inputs(213)) or (inputs(209));
    layer0_outputs(1554) <= (inputs(10)) and not (inputs(217));
    layer0_outputs(1555) <= inputs(103);
    layer0_outputs(1556) <= not(inputs(195));
    layer0_outputs(1557) <= (inputs(147)) or (inputs(234));
    layer0_outputs(1558) <= not(inputs(11)) or (inputs(236));
    layer0_outputs(1559) <= (inputs(6)) or (inputs(91));
    layer0_outputs(1560) <= (inputs(160)) xor (inputs(23));
    layer0_outputs(1561) <= (inputs(83)) or (inputs(15));
    layer0_outputs(1562) <= not(inputs(173)) or (inputs(99));
    layer0_outputs(1563) <= not(inputs(117));
    layer0_outputs(1564) <= not((inputs(244)) xor (inputs(195)));
    layer0_outputs(1565) <= not((inputs(202)) xor (inputs(244)));
    layer0_outputs(1566) <= '0';
    layer0_outputs(1567) <= not(inputs(42)) or (inputs(4));
    layer0_outputs(1568) <= inputs(101);
    layer0_outputs(1569) <= not(inputs(131));
    layer0_outputs(1570) <= inputs(57);
    layer0_outputs(1571) <= not(inputs(179));
    layer0_outputs(1572) <= inputs(62);
    layer0_outputs(1573) <= (inputs(192)) and not (inputs(94));
    layer0_outputs(1574) <= not((inputs(108)) xor (inputs(4)));
    layer0_outputs(1575) <= inputs(140);
    layer0_outputs(1576) <= not(inputs(157));
    layer0_outputs(1577) <= (inputs(168)) and not (inputs(49));
    layer0_outputs(1578) <= not(inputs(33)) or (inputs(200));
    layer0_outputs(1579) <= not((inputs(211)) or (inputs(166)));
    layer0_outputs(1580) <= not(inputs(14));
    layer0_outputs(1581) <= (inputs(22)) and not (inputs(148));
    layer0_outputs(1582) <= not((inputs(159)) or (inputs(131)));
    layer0_outputs(1583) <= not(inputs(205));
    layer0_outputs(1584) <= not((inputs(241)) or (inputs(13)));
    layer0_outputs(1585) <= not(inputs(87)) or (inputs(226));
    layer0_outputs(1586) <= (inputs(225)) or (inputs(162));
    layer0_outputs(1587) <= not(inputs(93)) or (inputs(47));
    layer0_outputs(1588) <= inputs(246);
    layer0_outputs(1589) <= (inputs(107)) or (inputs(10));
    layer0_outputs(1590) <= (inputs(128)) and (inputs(67));
    layer0_outputs(1591) <= not(inputs(209));
    layer0_outputs(1592) <= '0';
    layer0_outputs(1593) <= (inputs(197)) and not (inputs(190));
    layer0_outputs(1594) <= inputs(230);
    layer0_outputs(1595) <= inputs(191);
    layer0_outputs(1596) <= inputs(230);
    layer0_outputs(1597) <= not(inputs(89));
    layer0_outputs(1598) <= not((inputs(8)) or (inputs(24)));
    layer0_outputs(1599) <= (inputs(141)) or (inputs(12));
    layer0_outputs(1600) <= (inputs(171)) or (inputs(233));
    layer0_outputs(1601) <= inputs(102);
    layer0_outputs(1602) <= inputs(193);
    layer0_outputs(1603) <= (inputs(17)) or (inputs(197));
    layer0_outputs(1604) <= not(inputs(53));
    layer0_outputs(1605) <= (inputs(12)) or (inputs(157));
    layer0_outputs(1606) <= not(inputs(194));
    layer0_outputs(1607) <= inputs(237);
    layer0_outputs(1608) <= not(inputs(92));
    layer0_outputs(1609) <= not((inputs(142)) and (inputs(224)));
    layer0_outputs(1610) <= not(inputs(237));
    layer0_outputs(1611) <= (inputs(248)) and (inputs(19));
    layer0_outputs(1612) <= (inputs(223)) xor (inputs(249));
    layer0_outputs(1613) <= not(inputs(176));
    layer0_outputs(1614) <= (inputs(103)) and not (inputs(127));
    layer0_outputs(1615) <= inputs(98);
    layer0_outputs(1616) <= not((inputs(53)) or (inputs(111)));
    layer0_outputs(1617) <= not((inputs(254)) or (inputs(179)));
    layer0_outputs(1618) <= (inputs(81)) and not (inputs(158));
    layer0_outputs(1619) <= not(inputs(219)) or (inputs(18));
    layer0_outputs(1620) <= not(inputs(119));
    layer0_outputs(1621) <= (inputs(253)) or (inputs(68));
    layer0_outputs(1622) <= inputs(181);
    layer0_outputs(1623) <= inputs(108);
    layer0_outputs(1624) <= not(inputs(225)) or (inputs(174));
    layer0_outputs(1625) <= not(inputs(155));
    layer0_outputs(1626) <= (inputs(66)) or (inputs(38));
    layer0_outputs(1627) <= inputs(33);
    layer0_outputs(1628) <= not((inputs(226)) or (inputs(246)));
    layer0_outputs(1629) <= (inputs(105)) or (inputs(27));
    layer0_outputs(1630) <= (inputs(183)) and not (inputs(30));
    layer0_outputs(1631) <= not((inputs(64)) xor (inputs(121)));
    layer0_outputs(1632) <= not((inputs(5)) or (inputs(220)));
    layer0_outputs(1633) <= inputs(213);
    layer0_outputs(1634) <= not(inputs(102));
    layer0_outputs(1635) <= not(inputs(0));
    layer0_outputs(1636) <= not(inputs(185));
    layer0_outputs(1637) <= not(inputs(129));
    layer0_outputs(1638) <= (inputs(108)) or (inputs(99));
    layer0_outputs(1639) <= (inputs(141)) or (inputs(122));
    layer0_outputs(1640) <= not(inputs(74)) or (inputs(178));
    layer0_outputs(1641) <= inputs(108);
    layer0_outputs(1642) <= not((inputs(10)) or (inputs(197)));
    layer0_outputs(1643) <= inputs(161);
    layer0_outputs(1644) <= (inputs(121)) or (inputs(148));
    layer0_outputs(1645) <= not((inputs(203)) xor (inputs(148)));
    layer0_outputs(1646) <= inputs(132);
    layer0_outputs(1647) <= not(inputs(72));
    layer0_outputs(1648) <= inputs(162);
    layer0_outputs(1649) <= (inputs(46)) or (inputs(165));
    layer0_outputs(1650) <= (inputs(196)) xor (inputs(61));
    layer0_outputs(1651) <= not((inputs(224)) or (inputs(37)));
    layer0_outputs(1652) <= not((inputs(153)) and (inputs(89)));
    layer0_outputs(1653) <= not(inputs(245));
    layer0_outputs(1654) <= (inputs(76)) or (inputs(109));
    layer0_outputs(1655) <= not((inputs(151)) and (inputs(202)));
    layer0_outputs(1656) <= (inputs(221)) and not (inputs(126));
    layer0_outputs(1657) <= inputs(232);
    layer0_outputs(1658) <= not(inputs(236));
    layer0_outputs(1659) <= (inputs(243)) xor (inputs(123));
    layer0_outputs(1660) <= inputs(167);
    layer0_outputs(1661) <= not(inputs(234));
    layer0_outputs(1662) <= (inputs(150)) and not (inputs(14));
    layer0_outputs(1663) <= not(inputs(85));
    layer0_outputs(1664) <= not(inputs(50)) or (inputs(242));
    layer0_outputs(1665) <= not((inputs(3)) or (inputs(184)));
    layer0_outputs(1666) <= not(inputs(83)) or (inputs(125));
    layer0_outputs(1667) <= (inputs(156)) and not (inputs(255));
    layer0_outputs(1668) <= not((inputs(239)) or (inputs(12)));
    layer0_outputs(1669) <= inputs(60);
    layer0_outputs(1670) <= not(inputs(104)) or (inputs(222));
    layer0_outputs(1671) <= not(inputs(234));
    layer0_outputs(1672) <= (inputs(191)) or (inputs(72));
    layer0_outputs(1673) <= (inputs(183)) or (inputs(2));
    layer0_outputs(1674) <= not(inputs(150));
    layer0_outputs(1675) <= not(inputs(21)) or (inputs(61));
    layer0_outputs(1676) <= (inputs(201)) xor (inputs(214));
    layer0_outputs(1677) <= (inputs(202)) or (inputs(9));
    layer0_outputs(1678) <= not((inputs(17)) and (inputs(13)));
    layer0_outputs(1679) <= not(inputs(24));
    layer0_outputs(1680) <= not((inputs(171)) or (inputs(186)));
    layer0_outputs(1681) <= not((inputs(6)) or (inputs(39)));
    layer0_outputs(1682) <= not(inputs(133));
    layer0_outputs(1683) <= not(inputs(97)) or (inputs(142));
    layer0_outputs(1684) <= inputs(47);
    layer0_outputs(1685) <= '0';
    layer0_outputs(1686) <= not(inputs(15));
    layer0_outputs(1687) <= not(inputs(181));
    layer0_outputs(1688) <= inputs(130);
    layer0_outputs(1689) <= not(inputs(189)) or (inputs(64));
    layer0_outputs(1690) <= not((inputs(220)) xor (inputs(115)));
    layer0_outputs(1691) <= inputs(47);
    layer0_outputs(1692) <= (inputs(166)) and (inputs(6));
    layer0_outputs(1693) <= (inputs(191)) or (inputs(195));
    layer0_outputs(1694) <= '1';
    layer0_outputs(1695) <= (inputs(181)) and not (inputs(12));
    layer0_outputs(1696) <= (inputs(66)) xor (inputs(23));
    layer0_outputs(1697) <= (inputs(221)) or (inputs(242));
    layer0_outputs(1698) <= (inputs(3)) and not (inputs(209));
    layer0_outputs(1699) <= (inputs(220)) and not (inputs(78));
    layer0_outputs(1700) <= inputs(39);
    layer0_outputs(1701) <= (inputs(0)) xor (inputs(184));
    layer0_outputs(1702) <= not(inputs(179)) or (inputs(190));
    layer0_outputs(1703) <= not((inputs(151)) or (inputs(88)));
    layer0_outputs(1704) <= not(inputs(39));
    layer0_outputs(1705) <= not(inputs(178));
    layer0_outputs(1706) <= inputs(167);
    layer0_outputs(1707) <= inputs(147);
    layer0_outputs(1708) <= inputs(106);
    layer0_outputs(1709) <= not(inputs(185)) or (inputs(93));
    layer0_outputs(1710) <= not(inputs(76)) or (inputs(196));
    layer0_outputs(1711) <= inputs(120);
    layer0_outputs(1712) <= (inputs(86)) or (inputs(85));
    layer0_outputs(1713) <= not((inputs(97)) or (inputs(165)));
    layer0_outputs(1714) <= (inputs(104)) or (inputs(142));
    layer0_outputs(1715) <= (inputs(185)) or (inputs(2));
    layer0_outputs(1716) <= inputs(182);
    layer0_outputs(1717) <= not(inputs(90));
    layer0_outputs(1718) <= not(inputs(168));
    layer0_outputs(1719) <= not((inputs(68)) and (inputs(111)));
    layer0_outputs(1720) <= not(inputs(119)) or (inputs(163));
    layer0_outputs(1721) <= (inputs(173)) and (inputs(186));
    layer0_outputs(1722) <= not(inputs(227)) or (inputs(49));
    layer0_outputs(1723) <= '1';
    layer0_outputs(1724) <= (inputs(118)) and not (inputs(19));
    layer0_outputs(1725) <= not(inputs(5));
    layer0_outputs(1726) <= (inputs(216)) and not (inputs(13));
    layer0_outputs(1727) <= '0';
    layer0_outputs(1728) <= not((inputs(112)) or (inputs(83)));
    layer0_outputs(1729) <= not(inputs(172));
    layer0_outputs(1730) <= not((inputs(242)) or (inputs(232)));
    layer0_outputs(1731) <= (inputs(42)) and not (inputs(207));
    layer0_outputs(1732) <= (inputs(236)) and not (inputs(14));
    layer0_outputs(1733) <= (inputs(246)) or (inputs(15));
    layer0_outputs(1734) <= not((inputs(220)) or (inputs(174)));
    layer0_outputs(1735) <= (inputs(179)) or (inputs(181));
    layer0_outputs(1736) <= not(inputs(135)) or (inputs(194));
    layer0_outputs(1737) <= not((inputs(93)) xor (inputs(174)));
    layer0_outputs(1738) <= inputs(11);
    layer0_outputs(1739) <= not(inputs(73)) or (inputs(202));
    layer0_outputs(1740) <= (inputs(232)) and not (inputs(93));
    layer0_outputs(1741) <= not(inputs(227));
    layer0_outputs(1742) <= inputs(170);
    layer0_outputs(1743) <= (inputs(99)) or (inputs(226));
    layer0_outputs(1744) <= inputs(232);
    layer0_outputs(1745) <= not(inputs(73)) or (inputs(148));
    layer0_outputs(1746) <= not(inputs(15));
    layer0_outputs(1747) <= not(inputs(247)) or (inputs(168));
    layer0_outputs(1748) <= not(inputs(152));
    layer0_outputs(1749) <= (inputs(52)) or (inputs(254));
    layer0_outputs(1750) <= not(inputs(228));
    layer0_outputs(1751) <= not((inputs(130)) or (inputs(44)));
    layer0_outputs(1752) <= not((inputs(122)) xor (inputs(154)));
    layer0_outputs(1753) <= not(inputs(8));
    layer0_outputs(1754) <= inputs(246);
    layer0_outputs(1755) <= inputs(159);
    layer0_outputs(1756) <= not((inputs(153)) and (inputs(154)));
    layer0_outputs(1757) <= not((inputs(156)) or (inputs(124)));
    layer0_outputs(1758) <= (inputs(187)) and not (inputs(236));
    layer0_outputs(1759) <= not(inputs(67)) or (inputs(179));
    layer0_outputs(1760) <= inputs(247);
    layer0_outputs(1761) <= not(inputs(153)) or (inputs(228));
    layer0_outputs(1762) <= (inputs(249)) and not (inputs(76));
    layer0_outputs(1763) <= inputs(103);
    layer0_outputs(1764) <= (inputs(180)) and not (inputs(0));
    layer0_outputs(1765) <= (inputs(73)) or (inputs(38));
    layer0_outputs(1766) <= inputs(203);
    layer0_outputs(1767) <= not((inputs(172)) or (inputs(70)));
    layer0_outputs(1768) <= not(inputs(96)) or (inputs(128));
    layer0_outputs(1769) <= '0';
    layer0_outputs(1770) <= inputs(121);
    layer0_outputs(1771) <= not(inputs(59));
    layer0_outputs(1772) <= (inputs(246)) and (inputs(181));
    layer0_outputs(1773) <= inputs(28);
    layer0_outputs(1774) <= (inputs(212)) or (inputs(17));
    layer0_outputs(1775) <= not(inputs(85));
    layer0_outputs(1776) <= not(inputs(113));
    layer0_outputs(1777) <= (inputs(150)) or (inputs(168));
    layer0_outputs(1778) <= (inputs(212)) and not (inputs(33));
    layer0_outputs(1779) <= not(inputs(25));
    layer0_outputs(1780) <= not(inputs(77));
    layer0_outputs(1781) <= (inputs(40)) xor (inputs(56));
    layer0_outputs(1782) <= not(inputs(98));
    layer0_outputs(1783) <= not(inputs(40));
    layer0_outputs(1784) <= (inputs(97)) and not (inputs(95));
    layer0_outputs(1785) <= not((inputs(183)) or (inputs(194)));
    layer0_outputs(1786) <= not(inputs(22));
    layer0_outputs(1787) <= inputs(71);
    layer0_outputs(1788) <= inputs(40);
    layer0_outputs(1789) <= (inputs(43)) or (inputs(111));
    layer0_outputs(1790) <= inputs(51);
    layer0_outputs(1791) <= not(inputs(196));
    layer0_outputs(1792) <= not((inputs(136)) and (inputs(188)));
    layer0_outputs(1793) <= not((inputs(130)) and (inputs(251)));
    layer0_outputs(1794) <= (inputs(7)) or (inputs(180));
    layer0_outputs(1795) <= not((inputs(153)) xor (inputs(123)));
    layer0_outputs(1796) <= not((inputs(207)) or (inputs(5)));
    layer0_outputs(1797) <= inputs(199);
    layer0_outputs(1798) <= inputs(72);
    layer0_outputs(1799) <= inputs(168);
    layer0_outputs(1800) <= not(inputs(205));
    layer0_outputs(1801) <= not(inputs(194));
    layer0_outputs(1802) <= (inputs(91)) or (inputs(61));
    layer0_outputs(1803) <= not((inputs(33)) or (inputs(211)));
    layer0_outputs(1804) <= inputs(218);
    layer0_outputs(1805) <= (inputs(136)) or (inputs(222));
    layer0_outputs(1806) <= '0';
    layer0_outputs(1807) <= (inputs(102)) or (inputs(46));
    layer0_outputs(1808) <= not((inputs(199)) or (inputs(222)));
    layer0_outputs(1809) <= not((inputs(123)) or (inputs(189)));
    layer0_outputs(1810) <= not(inputs(211));
    layer0_outputs(1811) <= (inputs(96)) and not (inputs(161));
    layer0_outputs(1812) <= not(inputs(119));
    layer0_outputs(1813) <= not((inputs(5)) or (inputs(253)));
    layer0_outputs(1814) <= (inputs(84)) or (inputs(83));
    layer0_outputs(1815) <= not((inputs(108)) and (inputs(143)));
    layer0_outputs(1816) <= (inputs(179)) or (inputs(178));
    layer0_outputs(1817) <= (inputs(134)) and not (inputs(41));
    layer0_outputs(1818) <= not((inputs(142)) or (inputs(26)));
    layer0_outputs(1819) <= not(inputs(171)) or (inputs(215));
    layer0_outputs(1820) <= (inputs(166)) and (inputs(201));
    layer0_outputs(1821) <= (inputs(213)) or (inputs(206));
    layer0_outputs(1822) <= inputs(170);
    layer0_outputs(1823) <= (inputs(68)) and not (inputs(244));
    layer0_outputs(1824) <= (inputs(42)) or (inputs(4));
    layer0_outputs(1825) <= not(inputs(146));
    layer0_outputs(1826) <= (inputs(51)) and not (inputs(175));
    layer0_outputs(1827) <= (inputs(228)) or (inputs(160));
    layer0_outputs(1828) <= not((inputs(81)) xor (inputs(83)));
    layer0_outputs(1829) <= not(inputs(142));
    layer0_outputs(1830) <= not((inputs(45)) or (inputs(36)));
    layer0_outputs(1831) <= not(inputs(117));
    layer0_outputs(1832) <= inputs(121);
    layer0_outputs(1833) <= (inputs(3)) xor (inputs(62));
    layer0_outputs(1834) <= not(inputs(197));
    layer0_outputs(1835) <= not((inputs(79)) or (inputs(193)));
    layer0_outputs(1836) <= (inputs(171)) and not (inputs(68));
    layer0_outputs(1837) <= (inputs(160)) xor (inputs(23));
    layer0_outputs(1838) <= not((inputs(18)) or (inputs(224)));
    layer0_outputs(1839) <= (inputs(92)) and not (inputs(145));
    layer0_outputs(1840) <= (inputs(105)) and not (inputs(227));
    layer0_outputs(1841) <= not(inputs(68)) or (inputs(251));
    layer0_outputs(1842) <= not(inputs(45));
    layer0_outputs(1843) <= not(inputs(187));
    layer0_outputs(1844) <= not((inputs(27)) and (inputs(37)));
    layer0_outputs(1845) <= inputs(193);
    layer0_outputs(1846) <= not(inputs(146)) or (inputs(252));
    layer0_outputs(1847) <= not((inputs(54)) or (inputs(57)));
    layer0_outputs(1848) <= not(inputs(7)) or (inputs(160));
    layer0_outputs(1849) <= not((inputs(38)) xor (inputs(7)));
    layer0_outputs(1850) <= (inputs(40)) and not (inputs(220));
    layer0_outputs(1851) <= not(inputs(238));
    layer0_outputs(1852) <= not((inputs(50)) or (inputs(26)));
    layer0_outputs(1853) <= (inputs(101)) or (inputs(99));
    layer0_outputs(1854) <= not((inputs(87)) or (inputs(143)));
    layer0_outputs(1855) <= not(inputs(154)) or (inputs(74));
    layer0_outputs(1856) <= (inputs(168)) or (inputs(97));
    layer0_outputs(1857) <= not(inputs(150));
    layer0_outputs(1858) <= inputs(203);
    layer0_outputs(1859) <= not(inputs(35)) or (inputs(30));
    layer0_outputs(1860) <= (inputs(60)) or (inputs(0));
    layer0_outputs(1861) <= '1';
    layer0_outputs(1862) <= not(inputs(198));
    layer0_outputs(1863) <= not(inputs(83));
    layer0_outputs(1864) <= not(inputs(76)) or (inputs(161));
    layer0_outputs(1865) <= not((inputs(127)) and (inputs(241)));
    layer0_outputs(1866) <= not((inputs(192)) or (inputs(82)));
    layer0_outputs(1867) <= (inputs(127)) or (inputs(1));
    layer0_outputs(1868) <= inputs(39);
    layer0_outputs(1869) <= not(inputs(62));
    layer0_outputs(1870) <= inputs(68);
    layer0_outputs(1871) <= (inputs(158)) or (inputs(213));
    layer0_outputs(1872) <= (inputs(64)) or (inputs(229));
    layer0_outputs(1873) <= not(inputs(36)) or (inputs(79));
    layer0_outputs(1874) <= not(inputs(5));
    layer0_outputs(1875) <= not(inputs(37));
    layer0_outputs(1876) <= (inputs(100)) and not (inputs(28));
    layer0_outputs(1877) <= (inputs(127)) or (inputs(221));
    layer0_outputs(1878) <= not(inputs(101)) or (inputs(238));
    layer0_outputs(1879) <= (inputs(43)) xor (inputs(9));
    layer0_outputs(1880) <= (inputs(135)) and not (inputs(2));
    layer0_outputs(1881) <= (inputs(38)) and not (inputs(201));
    layer0_outputs(1882) <= not(inputs(0));
    layer0_outputs(1883) <= inputs(213);
    layer0_outputs(1884) <= not(inputs(63));
    layer0_outputs(1885) <= inputs(225);
    layer0_outputs(1886) <= not(inputs(51));
    layer0_outputs(1887) <= not((inputs(215)) and (inputs(75)));
    layer0_outputs(1888) <= (inputs(134)) and not (inputs(129));
    layer0_outputs(1889) <= inputs(123);
    layer0_outputs(1890) <= (inputs(182)) or (inputs(149));
    layer0_outputs(1891) <= (inputs(45)) xor (inputs(181));
    layer0_outputs(1892) <= (inputs(4)) or (inputs(32));
    layer0_outputs(1893) <= not(inputs(130));
    layer0_outputs(1894) <= (inputs(211)) or (inputs(236));
    layer0_outputs(1895) <= inputs(149);
    layer0_outputs(1896) <= not((inputs(163)) xor (inputs(172)));
    layer0_outputs(1897) <= not(inputs(52)) or (inputs(179));
    layer0_outputs(1898) <= (inputs(41)) xor (inputs(214));
    layer0_outputs(1899) <= inputs(117);
    layer0_outputs(1900) <= not(inputs(155)) or (inputs(16));
    layer0_outputs(1901) <= inputs(87);
    layer0_outputs(1902) <= '1';
    layer0_outputs(1903) <= (inputs(181)) and not (inputs(190));
    layer0_outputs(1904) <= not((inputs(81)) or (inputs(122)));
    layer0_outputs(1905) <= inputs(132);
    layer0_outputs(1906) <= '1';
    layer0_outputs(1907) <= not(inputs(205)) or (inputs(78));
    layer0_outputs(1908) <= not(inputs(91));
    layer0_outputs(1909) <= (inputs(119)) xor (inputs(155));
    layer0_outputs(1910) <= (inputs(122)) and not (inputs(143));
    layer0_outputs(1911) <= not(inputs(73)) or (inputs(8));
    layer0_outputs(1912) <= not((inputs(219)) or (inputs(156)));
    layer0_outputs(1913) <= not((inputs(145)) or (inputs(88)));
    layer0_outputs(1914) <= not((inputs(146)) or (inputs(216)));
    layer0_outputs(1915) <= inputs(248);
    layer0_outputs(1916) <= (inputs(57)) and not (inputs(174));
    layer0_outputs(1917) <= not((inputs(160)) xor (inputs(131)));
    layer0_outputs(1918) <= not(inputs(159));
    layer0_outputs(1919) <= (inputs(245)) and not (inputs(153));
    layer0_outputs(1920) <= inputs(229);
    layer0_outputs(1921) <= not(inputs(25));
    layer0_outputs(1922) <= inputs(214);
    layer0_outputs(1923) <= not((inputs(46)) or (inputs(158)));
    layer0_outputs(1924) <= not((inputs(148)) or (inputs(237)));
    layer0_outputs(1925) <= (inputs(23)) and not (inputs(241));
    layer0_outputs(1926) <= not(inputs(97));
    layer0_outputs(1927) <= not((inputs(164)) or (inputs(215)));
    layer0_outputs(1928) <= not(inputs(153));
    layer0_outputs(1929) <= inputs(21);
    layer0_outputs(1930) <= not((inputs(172)) and (inputs(121)));
    layer0_outputs(1931) <= not(inputs(215));
    layer0_outputs(1932) <= not((inputs(222)) xor (inputs(139)));
    layer0_outputs(1933) <= not(inputs(208));
    layer0_outputs(1934) <= inputs(182);
    layer0_outputs(1935) <= (inputs(96)) and not (inputs(128));
    layer0_outputs(1936) <= not(inputs(100));
    layer0_outputs(1937) <= not(inputs(101));
    layer0_outputs(1938) <= not((inputs(203)) or (inputs(185)));
    layer0_outputs(1939) <= not(inputs(243));
    layer0_outputs(1940) <= (inputs(243)) xor (inputs(113));
    layer0_outputs(1941) <= not((inputs(231)) or (inputs(177)));
    layer0_outputs(1942) <= not(inputs(39));
    layer0_outputs(1943) <= '1';
    layer0_outputs(1944) <= not(inputs(101));
    layer0_outputs(1945) <= not((inputs(107)) xor (inputs(1)));
    layer0_outputs(1946) <= '1';
    layer0_outputs(1947) <= (inputs(164)) xor (inputs(133));
    layer0_outputs(1948) <= (inputs(49)) or (inputs(157));
    layer0_outputs(1949) <= (inputs(9)) or (inputs(159));
    layer0_outputs(1950) <= inputs(153);
    layer0_outputs(1951) <= inputs(161);
    layer0_outputs(1952) <= (inputs(253)) or (inputs(78));
    layer0_outputs(1953) <= (inputs(150)) and not (inputs(140));
    layer0_outputs(1954) <= not(inputs(117));
    layer0_outputs(1955) <= (inputs(123)) or (inputs(30));
    layer0_outputs(1956) <= (inputs(151)) or (inputs(110));
    layer0_outputs(1957) <= not(inputs(87));
    layer0_outputs(1958) <= (inputs(206)) or (inputs(128));
    layer0_outputs(1959) <= (inputs(162)) or (inputs(13));
    layer0_outputs(1960) <= not(inputs(9)) or (inputs(238));
    layer0_outputs(1961) <= (inputs(153)) or (inputs(250));
    layer0_outputs(1962) <= (inputs(12)) or (inputs(248));
    layer0_outputs(1963) <= (inputs(3)) or (inputs(50));
    layer0_outputs(1964) <= not(inputs(100));
    layer0_outputs(1965) <= inputs(122);
    layer0_outputs(1966) <= inputs(220);
    layer0_outputs(1967) <= not(inputs(77));
    layer0_outputs(1968) <= not(inputs(233)) or (inputs(30));
    layer0_outputs(1969) <= (inputs(237)) and (inputs(47));
    layer0_outputs(1970) <= not((inputs(72)) xor (inputs(31)));
    layer0_outputs(1971) <= not((inputs(79)) or (inputs(58)));
    layer0_outputs(1972) <= inputs(124);
    layer0_outputs(1973) <= (inputs(23)) and not (inputs(82));
    layer0_outputs(1974) <= not(inputs(156));
    layer0_outputs(1975) <= (inputs(14)) or (inputs(26));
    layer0_outputs(1976) <= not(inputs(227)) or (inputs(164));
    layer0_outputs(1977) <= not(inputs(215));
    layer0_outputs(1978) <= (inputs(70)) xor (inputs(86));
    layer0_outputs(1979) <= (inputs(247)) and not (inputs(209));
    layer0_outputs(1980) <= inputs(151);
    layer0_outputs(1981) <= inputs(94);
    layer0_outputs(1982) <= (inputs(176)) and not (inputs(142));
    layer0_outputs(1983) <= not((inputs(74)) or (inputs(130)));
    layer0_outputs(1984) <= not(inputs(109));
    layer0_outputs(1985) <= inputs(101);
    layer0_outputs(1986) <= not(inputs(91));
    layer0_outputs(1987) <= not((inputs(203)) or (inputs(97)));
    layer0_outputs(1988) <= not(inputs(61));
    layer0_outputs(1989) <= not(inputs(84));
    layer0_outputs(1990) <= '1';
    layer0_outputs(1991) <= not(inputs(211)) or (inputs(31));
    layer0_outputs(1992) <= inputs(92);
    layer0_outputs(1993) <= (inputs(65)) and (inputs(160));
    layer0_outputs(1994) <= (inputs(180)) and not (inputs(155));
    layer0_outputs(1995) <= not(inputs(245));
    layer0_outputs(1996) <= inputs(121);
    layer0_outputs(1997) <= (inputs(206)) or (inputs(190));
    layer0_outputs(1998) <= (inputs(84)) or (inputs(193));
    layer0_outputs(1999) <= inputs(173);
    layer0_outputs(2000) <= not((inputs(173)) or (inputs(84)));
    layer0_outputs(2001) <= '0';
    layer0_outputs(2002) <= not((inputs(8)) xor (inputs(223)));
    layer0_outputs(2003) <= not(inputs(131));
    layer0_outputs(2004) <= (inputs(116)) and not (inputs(243));
    layer0_outputs(2005) <= (inputs(109)) and not (inputs(30));
    layer0_outputs(2006) <= (inputs(180)) and not (inputs(241));
    layer0_outputs(2007) <= (inputs(204)) and not (inputs(99));
    layer0_outputs(2008) <= inputs(18);
    layer0_outputs(2009) <= inputs(118);
    layer0_outputs(2010) <= not(inputs(84));
    layer0_outputs(2011) <= not(inputs(80)) or (inputs(69));
    layer0_outputs(2012) <= inputs(57);
    layer0_outputs(2013) <= (inputs(93)) and not (inputs(245));
    layer0_outputs(2014) <= not(inputs(162));
    layer0_outputs(2015) <= '1';
    layer0_outputs(2016) <= (inputs(22)) and not (inputs(238));
    layer0_outputs(2017) <= (inputs(19)) and not (inputs(192));
    layer0_outputs(2018) <= (inputs(75)) and not (inputs(57));
    layer0_outputs(2019) <= not((inputs(87)) xor (inputs(212)));
    layer0_outputs(2020) <= '0';
    layer0_outputs(2021) <= not(inputs(103)) or (inputs(249));
    layer0_outputs(2022) <= not((inputs(169)) xor (inputs(218)));
    layer0_outputs(2023) <= inputs(89);
    layer0_outputs(2024) <= (inputs(31)) or (inputs(242));
    layer0_outputs(2025) <= not((inputs(42)) or (inputs(240)));
    layer0_outputs(2026) <= inputs(35);
    layer0_outputs(2027) <= (inputs(98)) and not (inputs(94));
    layer0_outputs(2028) <= not((inputs(201)) or (inputs(181)));
    layer0_outputs(2029) <= not((inputs(69)) xor (inputs(5)));
    layer0_outputs(2030) <= not((inputs(45)) or (inputs(50)));
    layer0_outputs(2031) <= (inputs(143)) or (inputs(153));
    layer0_outputs(2032) <= inputs(206);
    layer0_outputs(2033) <= not(inputs(184));
    layer0_outputs(2034) <= inputs(88);
    layer0_outputs(2035) <= not(inputs(228)) or (inputs(129));
    layer0_outputs(2036) <= not(inputs(150));
    layer0_outputs(2037) <= (inputs(169)) and not (inputs(187));
    layer0_outputs(2038) <= (inputs(229)) or (inputs(197));
    layer0_outputs(2039) <= (inputs(174)) or (inputs(114));
    layer0_outputs(2040) <= not(inputs(95));
    layer0_outputs(2041) <= (inputs(116)) xor (inputs(66));
    layer0_outputs(2042) <= not(inputs(152));
    layer0_outputs(2043) <= not(inputs(102)) or (inputs(186));
    layer0_outputs(2044) <= inputs(211);
    layer0_outputs(2045) <= not(inputs(200));
    layer0_outputs(2046) <= not((inputs(200)) xor (inputs(95)));
    layer0_outputs(2047) <= (inputs(77)) or (inputs(94));
    layer0_outputs(2048) <= not(inputs(40)) or (inputs(209));
    layer0_outputs(2049) <= (inputs(55)) and not (inputs(95));
    layer0_outputs(2050) <= not(inputs(131));
    layer0_outputs(2051) <= inputs(222);
    layer0_outputs(2052) <= not(inputs(72)) or (inputs(128));
    layer0_outputs(2053) <= not(inputs(94)) or (inputs(48));
    layer0_outputs(2054) <= not(inputs(245)) or (inputs(119));
    layer0_outputs(2055) <= not((inputs(223)) or (inputs(185)));
    layer0_outputs(2056) <= not((inputs(12)) or (inputs(119)));
    layer0_outputs(2057) <= inputs(232);
    layer0_outputs(2058) <= (inputs(236)) or (inputs(223));
    layer0_outputs(2059) <= (inputs(127)) or (inputs(36));
    layer0_outputs(2060) <= inputs(70);
    layer0_outputs(2061) <= (inputs(166)) or (inputs(68));
    layer0_outputs(2062) <= (inputs(175)) and not (inputs(207));
    layer0_outputs(2063) <= inputs(118);
    layer0_outputs(2064) <= not(inputs(255));
    layer0_outputs(2065) <= not((inputs(186)) and (inputs(54)));
    layer0_outputs(2066) <= not(inputs(216));
    layer0_outputs(2067) <= (inputs(3)) and not (inputs(47));
    layer0_outputs(2068) <= inputs(211);
    layer0_outputs(2069) <= (inputs(116)) xor (inputs(113));
    layer0_outputs(2070) <= not(inputs(79));
    layer0_outputs(2071) <= not((inputs(139)) or (inputs(173)));
    layer0_outputs(2072) <= not(inputs(18)) or (inputs(191));
    layer0_outputs(2073) <= not(inputs(166));
    layer0_outputs(2074) <= inputs(9);
    layer0_outputs(2075) <= not(inputs(99)) or (inputs(88));
    layer0_outputs(2076) <= not((inputs(241)) or (inputs(138)));
    layer0_outputs(2077) <= inputs(91);
    layer0_outputs(2078) <= (inputs(82)) xor (inputs(37));
    layer0_outputs(2079) <= (inputs(188)) or (inputs(161));
    layer0_outputs(2080) <= inputs(220);
    layer0_outputs(2081) <= (inputs(160)) and not (inputs(188));
    layer0_outputs(2082) <= not(inputs(252));
    layer0_outputs(2083) <= '1';
    layer0_outputs(2084) <= (inputs(102)) and not (inputs(33));
    layer0_outputs(2085) <= not(inputs(120)) or (inputs(182));
    layer0_outputs(2086) <= not((inputs(226)) or (inputs(163)));
    layer0_outputs(2087) <= not(inputs(226)) or (inputs(163));
    layer0_outputs(2088) <= (inputs(113)) or (inputs(154));
    layer0_outputs(2089) <= not(inputs(220));
    layer0_outputs(2090) <= '0';
    layer0_outputs(2091) <= not(inputs(126));
    layer0_outputs(2092) <= not(inputs(179));
    layer0_outputs(2093) <= inputs(163);
    layer0_outputs(2094) <= not(inputs(86));
    layer0_outputs(2095) <= (inputs(37)) or (inputs(131));
    layer0_outputs(2096) <= (inputs(47)) or (inputs(0));
    layer0_outputs(2097) <= '1';
    layer0_outputs(2098) <= not((inputs(245)) or (inputs(180)));
    layer0_outputs(2099) <= (inputs(113)) or (inputs(180));
    layer0_outputs(2100) <= (inputs(141)) xor (inputs(107));
    layer0_outputs(2101) <= inputs(38);
    layer0_outputs(2102) <= not((inputs(97)) xor (inputs(35)));
    layer0_outputs(2103) <= not((inputs(110)) or (inputs(46)));
    layer0_outputs(2104) <= not(inputs(221)) or (inputs(83));
    layer0_outputs(2105) <= '1';
    layer0_outputs(2106) <= not(inputs(103)) or (inputs(217));
    layer0_outputs(2107) <= inputs(79);
    layer0_outputs(2108) <= not((inputs(73)) or (inputs(207)));
    layer0_outputs(2109) <= not((inputs(62)) or (inputs(8)));
    layer0_outputs(2110) <= inputs(95);
    layer0_outputs(2111) <= inputs(59);
    layer0_outputs(2112) <= not(inputs(199)) or (inputs(53));
    layer0_outputs(2113) <= inputs(186);
    layer0_outputs(2114) <= (inputs(100)) or (inputs(188));
    layer0_outputs(2115) <= '0';
    layer0_outputs(2116) <= not(inputs(140));
    layer0_outputs(2117) <= not(inputs(146)) or (inputs(152));
    layer0_outputs(2118) <= (inputs(33)) and (inputs(31));
    layer0_outputs(2119) <= not(inputs(81)) or (inputs(93));
    layer0_outputs(2120) <= (inputs(94)) and not (inputs(240));
    layer0_outputs(2121) <= not(inputs(221));
    layer0_outputs(2122) <= not(inputs(181));
    layer0_outputs(2123) <= not(inputs(247));
    layer0_outputs(2124) <= (inputs(212)) xor (inputs(175));
    layer0_outputs(2125) <= inputs(128);
    layer0_outputs(2126) <= not(inputs(8)) or (inputs(19));
    layer0_outputs(2127) <= not(inputs(243));
    layer0_outputs(2128) <= inputs(58);
    layer0_outputs(2129) <= inputs(60);
    layer0_outputs(2130) <= not((inputs(5)) or (inputs(17)));
    layer0_outputs(2131) <= not(inputs(85));
    layer0_outputs(2132) <= (inputs(101)) and not (inputs(160));
    layer0_outputs(2133) <= (inputs(167)) or (inputs(178));
    layer0_outputs(2134) <= inputs(81);
    layer0_outputs(2135) <= not(inputs(39));
    layer0_outputs(2136) <= inputs(230);
    layer0_outputs(2137) <= not((inputs(198)) or (inputs(0)));
    layer0_outputs(2138) <= not(inputs(26)) or (inputs(89));
    layer0_outputs(2139) <= (inputs(2)) and (inputs(35));
    layer0_outputs(2140) <= (inputs(68)) or (inputs(193));
    layer0_outputs(2141) <= inputs(230);
    layer0_outputs(2142) <= not((inputs(89)) or (inputs(205)));
    layer0_outputs(2143) <= not((inputs(19)) or (inputs(21)));
    layer0_outputs(2144) <= (inputs(212)) and not (inputs(169));
    layer0_outputs(2145) <= not(inputs(176));
    layer0_outputs(2146) <= not((inputs(27)) xor (inputs(6)));
    layer0_outputs(2147) <= (inputs(181)) xor (inputs(90));
    layer0_outputs(2148) <= not(inputs(90));
    layer0_outputs(2149) <= (inputs(81)) and not (inputs(159));
    layer0_outputs(2150) <= not(inputs(131));
    layer0_outputs(2151) <= not(inputs(223));
    layer0_outputs(2152) <= not(inputs(67)) or (inputs(51));
    layer0_outputs(2153) <= not((inputs(41)) or (inputs(113)));
    layer0_outputs(2154) <= '0';
    layer0_outputs(2155) <= not(inputs(181));
    layer0_outputs(2156) <= not((inputs(19)) or (inputs(208)));
    layer0_outputs(2157) <= (inputs(132)) and not (inputs(73));
    layer0_outputs(2158) <= not(inputs(91));
    layer0_outputs(2159) <= inputs(75);
    layer0_outputs(2160) <= (inputs(56)) and not (inputs(19));
    layer0_outputs(2161) <= not((inputs(33)) or (inputs(139)));
    layer0_outputs(2162) <= not((inputs(222)) or (inputs(92)));
    layer0_outputs(2163) <= (inputs(81)) or (inputs(203));
    layer0_outputs(2164) <= inputs(81);
    layer0_outputs(2165) <= not((inputs(91)) or (inputs(93)));
    layer0_outputs(2166) <= not(inputs(247)) or (inputs(155));
    layer0_outputs(2167) <= not(inputs(13));
    layer0_outputs(2168) <= not((inputs(230)) and (inputs(121)));
    layer0_outputs(2169) <= (inputs(55)) and not (inputs(200));
    layer0_outputs(2170) <= inputs(234);
    layer0_outputs(2171) <= '0';
    layer0_outputs(2172) <= not((inputs(162)) or (inputs(246)));
    layer0_outputs(2173) <= (inputs(106)) and not (inputs(143));
    layer0_outputs(2174) <= (inputs(150)) and not (inputs(116));
    layer0_outputs(2175) <= not((inputs(33)) or (inputs(129)));
    layer0_outputs(2176) <= inputs(180);
    layer0_outputs(2177) <= not(inputs(183)) or (inputs(48));
    layer0_outputs(2178) <= not(inputs(90));
    layer0_outputs(2179) <= (inputs(35)) xor (inputs(236));
    layer0_outputs(2180) <= not(inputs(242));
    layer0_outputs(2181) <= not(inputs(52));
    layer0_outputs(2182) <= not(inputs(112));
    layer0_outputs(2183) <= (inputs(189)) or (inputs(85));
    layer0_outputs(2184) <= not((inputs(104)) or (inputs(92)));
    layer0_outputs(2185) <= not(inputs(230)) or (inputs(108));
    layer0_outputs(2186) <= (inputs(106)) or (inputs(105));
    layer0_outputs(2187) <= not(inputs(210));
    layer0_outputs(2188) <= (inputs(62)) and (inputs(56));
    layer0_outputs(2189) <= not(inputs(133));
    layer0_outputs(2190) <= not(inputs(89));
    layer0_outputs(2191) <= not((inputs(192)) or (inputs(169)));
    layer0_outputs(2192) <= '0';
    layer0_outputs(2193) <= not(inputs(235));
    layer0_outputs(2194) <= not(inputs(29));
    layer0_outputs(2195) <= not((inputs(84)) or (inputs(0)));
    layer0_outputs(2196) <= '1';
    layer0_outputs(2197) <= (inputs(27)) or (inputs(48));
    layer0_outputs(2198) <= inputs(221);
    layer0_outputs(2199) <= (inputs(49)) xor (inputs(15));
    layer0_outputs(2200) <= '0';
    layer0_outputs(2201) <= (inputs(87)) or (inputs(214));
    layer0_outputs(2202) <= inputs(87);
    layer0_outputs(2203) <= inputs(44);
    layer0_outputs(2204) <= (inputs(196)) and not (inputs(254));
    layer0_outputs(2205) <= (inputs(145)) or (inputs(95));
    layer0_outputs(2206) <= not((inputs(176)) or (inputs(192)));
    layer0_outputs(2207) <= not((inputs(68)) or (inputs(207)));
    layer0_outputs(2208) <= not((inputs(209)) or (inputs(229)));
    layer0_outputs(2209) <= not(inputs(74));
    layer0_outputs(2210) <= not((inputs(115)) and (inputs(134)));
    layer0_outputs(2211) <= inputs(152);
    layer0_outputs(2212) <= (inputs(11)) and not (inputs(202));
    layer0_outputs(2213) <= (inputs(156)) or (inputs(172));
    layer0_outputs(2214) <= not(inputs(168)) or (inputs(126));
    layer0_outputs(2215) <= (inputs(82)) and not (inputs(233));
    layer0_outputs(2216) <= (inputs(65)) or (inputs(214));
    layer0_outputs(2217) <= (inputs(180)) xor (inputs(112));
    layer0_outputs(2218) <= not(inputs(116));
    layer0_outputs(2219) <= (inputs(81)) xor (inputs(52));
    layer0_outputs(2220) <= inputs(228);
    layer0_outputs(2221) <= (inputs(125)) or (inputs(93));
    layer0_outputs(2222) <= (inputs(19)) or (inputs(2));
    layer0_outputs(2223) <= not(inputs(135));
    layer0_outputs(2224) <= not((inputs(200)) xor (inputs(14)));
    layer0_outputs(2225) <= (inputs(38)) and not (inputs(219));
    layer0_outputs(2226) <= (inputs(218)) or (inputs(205));
    layer0_outputs(2227) <= inputs(165);
    layer0_outputs(2228) <= inputs(124);
    layer0_outputs(2229) <= not((inputs(177)) or (inputs(214)));
    layer0_outputs(2230) <= '1';
    layer0_outputs(2231) <= (inputs(92)) or (inputs(111));
    layer0_outputs(2232) <= not((inputs(205)) xor (inputs(216)));
    layer0_outputs(2233) <= not(inputs(178));
    layer0_outputs(2234) <= (inputs(187)) or (inputs(3));
    layer0_outputs(2235) <= not((inputs(35)) or (inputs(172)));
    layer0_outputs(2236) <= inputs(138);
    layer0_outputs(2237) <= '0';
    layer0_outputs(2238) <= (inputs(189)) or (inputs(175));
    layer0_outputs(2239) <= inputs(246);
    layer0_outputs(2240) <= (inputs(72)) and (inputs(174));
    layer0_outputs(2241) <= inputs(231);
    layer0_outputs(2242) <= (inputs(236)) or (inputs(51));
    layer0_outputs(2243) <= not((inputs(208)) or (inputs(32)));
    layer0_outputs(2244) <= inputs(185);
    layer0_outputs(2245) <= '0';
    layer0_outputs(2246) <= not(inputs(32)) or (inputs(239));
    layer0_outputs(2247) <= inputs(233);
    layer0_outputs(2248) <= not(inputs(52)) or (inputs(241));
    layer0_outputs(2249) <= not(inputs(22)) or (inputs(31));
    layer0_outputs(2250) <= (inputs(149)) and (inputs(229));
    layer0_outputs(2251) <= not((inputs(37)) or (inputs(33)));
    layer0_outputs(2252) <= not(inputs(135)) or (inputs(191));
    layer0_outputs(2253) <= inputs(248);
    layer0_outputs(2254) <= '0';
    layer0_outputs(2255) <= not((inputs(128)) or (inputs(244)));
    layer0_outputs(2256) <= (inputs(64)) or (inputs(112));
    layer0_outputs(2257) <= not(inputs(124));
    layer0_outputs(2258) <= (inputs(147)) and not (inputs(3));
    layer0_outputs(2259) <= not(inputs(181));
    layer0_outputs(2260) <= (inputs(62)) or (inputs(69));
    layer0_outputs(2261) <= inputs(132);
    layer0_outputs(2262) <= inputs(84);
    layer0_outputs(2263) <= (inputs(146)) or (inputs(146));
    layer0_outputs(2264) <= (inputs(16)) and (inputs(128));
    layer0_outputs(2265) <= (inputs(143)) or (inputs(112));
    layer0_outputs(2266) <= not((inputs(111)) or (inputs(10)));
    layer0_outputs(2267) <= (inputs(180)) or (inputs(251));
    layer0_outputs(2268) <= (inputs(105)) and not (inputs(206));
    layer0_outputs(2269) <= not((inputs(82)) xor (inputs(28)));
    layer0_outputs(2270) <= (inputs(49)) or (inputs(38));
    layer0_outputs(2271) <= inputs(89);
    layer0_outputs(2272) <= not(inputs(233)) or (inputs(13));
    layer0_outputs(2273) <= inputs(34);
    layer0_outputs(2274) <= (inputs(182)) and not (inputs(189));
    layer0_outputs(2275) <= inputs(227);
    layer0_outputs(2276) <= not((inputs(34)) and (inputs(4)));
    layer0_outputs(2277) <= (inputs(242)) xor (inputs(232));
    layer0_outputs(2278) <= (inputs(111)) or (inputs(88));
    layer0_outputs(2279) <= not(inputs(41));
    layer0_outputs(2280) <= not(inputs(68));
    layer0_outputs(2281) <= not(inputs(24));
    layer0_outputs(2282) <= inputs(25);
    layer0_outputs(2283) <= (inputs(64)) xor (inputs(156));
    layer0_outputs(2284) <= inputs(232);
    layer0_outputs(2285) <= (inputs(255)) xor (inputs(88));
    layer0_outputs(2286) <= not((inputs(0)) xor (inputs(107)));
    layer0_outputs(2287) <= inputs(171);
    layer0_outputs(2288) <= not(inputs(107));
    layer0_outputs(2289) <= (inputs(80)) or (inputs(215));
    layer0_outputs(2290) <= (inputs(241)) and not (inputs(121));
    layer0_outputs(2291) <= not(inputs(27)) or (inputs(189));
    layer0_outputs(2292) <= inputs(6);
    layer0_outputs(2293) <= not((inputs(159)) or (inputs(175)));
    layer0_outputs(2294) <= (inputs(128)) xor (inputs(195));
    layer0_outputs(2295) <= (inputs(218)) and not (inputs(153));
    layer0_outputs(2296) <= not((inputs(248)) xor (inputs(231)));
    layer0_outputs(2297) <= not(inputs(228));
    layer0_outputs(2298) <= (inputs(3)) and not (inputs(160));
    layer0_outputs(2299) <= (inputs(67)) or (inputs(187));
    layer0_outputs(2300) <= not((inputs(247)) or (inputs(195)));
    layer0_outputs(2301) <= (inputs(230)) and not (inputs(90));
    layer0_outputs(2302) <= not((inputs(125)) or (inputs(26)));
    layer0_outputs(2303) <= (inputs(159)) or (inputs(129));
    layer0_outputs(2304) <= (inputs(164)) or (inputs(166));
    layer0_outputs(2305) <= (inputs(98)) or (inputs(210));
    layer0_outputs(2306) <= not(inputs(85));
    layer0_outputs(2307) <= inputs(88);
    layer0_outputs(2308) <= inputs(133);
    layer0_outputs(2309) <= inputs(193);
    layer0_outputs(2310) <= inputs(153);
    layer0_outputs(2311) <= not(inputs(69));
    layer0_outputs(2312) <= not((inputs(218)) and (inputs(27)));
    layer0_outputs(2313) <= (inputs(10)) and not (inputs(19));
    layer0_outputs(2314) <= not(inputs(136)) or (inputs(96));
    layer0_outputs(2315) <= (inputs(61)) xor (inputs(67));
    layer0_outputs(2316) <= not((inputs(250)) xor (inputs(63)));
    layer0_outputs(2317) <= not(inputs(247)) or (inputs(94));
    layer0_outputs(2318) <= not((inputs(10)) and (inputs(8)));
    layer0_outputs(2319) <= not(inputs(29));
    layer0_outputs(2320) <= (inputs(126)) or (inputs(12));
    layer0_outputs(2321) <= not((inputs(69)) and (inputs(217)));
    layer0_outputs(2322) <= not(inputs(59)) or (inputs(191));
    layer0_outputs(2323) <= inputs(83);
    layer0_outputs(2324) <= (inputs(188)) or (inputs(4));
    layer0_outputs(2325) <= '1';
    layer0_outputs(2326) <= (inputs(198)) or (inputs(238));
    layer0_outputs(2327) <= not((inputs(150)) or (inputs(161)));
    layer0_outputs(2328) <= (inputs(22)) or (inputs(110));
    layer0_outputs(2329) <= (inputs(120)) and not (inputs(176));
    layer0_outputs(2330) <= not((inputs(129)) or (inputs(103)));
    layer0_outputs(2331) <= (inputs(38)) and not (inputs(253));
    layer0_outputs(2332) <= not(inputs(167));
    layer0_outputs(2333) <= not((inputs(194)) or (inputs(86)));
    layer0_outputs(2334) <= (inputs(59)) xor (inputs(245));
    layer0_outputs(2335) <= not(inputs(115));
    layer0_outputs(2336) <= (inputs(121)) xor (inputs(128));
    layer0_outputs(2337) <= inputs(90);
    layer0_outputs(2338) <= not((inputs(125)) xor (inputs(122)));
    layer0_outputs(2339) <= (inputs(118)) or (inputs(108));
    layer0_outputs(2340) <= not(inputs(152));
    layer0_outputs(2341) <= (inputs(50)) and not (inputs(145));
    layer0_outputs(2342) <= inputs(183);
    layer0_outputs(2343) <= (inputs(66)) or (inputs(198));
    layer0_outputs(2344) <= (inputs(222)) xor (inputs(69));
    layer0_outputs(2345) <= inputs(235);
    layer0_outputs(2346) <= not(inputs(40)) or (inputs(239));
    layer0_outputs(2347) <= not((inputs(95)) xor (inputs(75)));
    layer0_outputs(2348) <= not(inputs(193)) or (inputs(112));
    layer0_outputs(2349) <= not((inputs(11)) and (inputs(72)));
    layer0_outputs(2350) <= inputs(210);
    layer0_outputs(2351) <= (inputs(229)) and not (inputs(102));
    layer0_outputs(2352) <= (inputs(237)) or (inputs(82));
    layer0_outputs(2353) <= not(inputs(163)) or (inputs(63));
    layer0_outputs(2354) <= not((inputs(202)) and (inputs(202)));
    layer0_outputs(2355) <= not(inputs(133));
    layer0_outputs(2356) <= inputs(67);
    layer0_outputs(2357) <= not(inputs(183));
    layer0_outputs(2358) <= not(inputs(139)) or (inputs(225));
    layer0_outputs(2359) <= not((inputs(166)) or (inputs(152)));
    layer0_outputs(2360) <= not(inputs(99));
    layer0_outputs(2361) <= '0';
    layer0_outputs(2362) <= not((inputs(242)) or (inputs(176)));
    layer0_outputs(2363) <= (inputs(162)) or (inputs(65));
    layer0_outputs(2364) <= (inputs(12)) xor (inputs(6));
    layer0_outputs(2365) <= (inputs(228)) or (inputs(37));
    layer0_outputs(2366) <= inputs(103);
    layer0_outputs(2367) <= inputs(245);
    layer0_outputs(2368) <= not((inputs(45)) xor (inputs(207)));
    layer0_outputs(2369) <= inputs(34);
    layer0_outputs(2370) <= not((inputs(231)) and (inputs(120)));
    layer0_outputs(2371) <= not(inputs(33)) or (inputs(197));
    layer0_outputs(2372) <= inputs(208);
    layer0_outputs(2373) <= not((inputs(54)) or (inputs(62)));
    layer0_outputs(2374) <= (inputs(212)) xor (inputs(40));
    layer0_outputs(2375) <= (inputs(29)) and (inputs(38));
    layer0_outputs(2376) <= not(inputs(246));
    layer0_outputs(2377) <= not(inputs(27));
    layer0_outputs(2378) <= '0';
    layer0_outputs(2379) <= not((inputs(148)) or (inputs(166)));
    layer0_outputs(2380) <= not((inputs(32)) xor (inputs(210)));
    layer0_outputs(2381) <= not(inputs(44)) or (inputs(191));
    layer0_outputs(2382) <= not((inputs(80)) or (inputs(84)));
    layer0_outputs(2383) <= inputs(144);
    layer0_outputs(2384) <= inputs(113);
    layer0_outputs(2385) <= not((inputs(130)) or (inputs(185)));
    layer0_outputs(2386) <= (inputs(194)) xor (inputs(149));
    layer0_outputs(2387) <= (inputs(247)) and not (inputs(253));
    layer0_outputs(2388) <= (inputs(192)) or (inputs(219));
    layer0_outputs(2389) <= (inputs(128)) or (inputs(122));
    layer0_outputs(2390) <= inputs(250);
    layer0_outputs(2391) <= (inputs(174)) or (inputs(20));
    layer0_outputs(2392) <= not(inputs(215)) or (inputs(2));
    layer0_outputs(2393) <= inputs(147);
    layer0_outputs(2394) <= (inputs(209)) or (inputs(116));
    layer0_outputs(2395) <= (inputs(113)) or (inputs(248));
    layer0_outputs(2396) <= not((inputs(218)) xor (inputs(188)));
    layer0_outputs(2397) <= not((inputs(51)) or (inputs(10)));
    layer0_outputs(2398) <= not((inputs(97)) or (inputs(192)));
    layer0_outputs(2399) <= not((inputs(167)) or (inputs(255)));
    layer0_outputs(2400) <= '0';
    layer0_outputs(2401) <= (inputs(68)) xor (inputs(50));
    layer0_outputs(2402) <= inputs(162);
    layer0_outputs(2403) <= (inputs(132)) and not (inputs(20));
    layer0_outputs(2404) <= not(inputs(39));
    layer0_outputs(2405) <= not((inputs(23)) or (inputs(47)));
    layer0_outputs(2406) <= not((inputs(13)) or (inputs(86)));
    layer0_outputs(2407) <= inputs(133);
    layer0_outputs(2408) <= not(inputs(75)) or (inputs(151));
    layer0_outputs(2409) <= (inputs(71)) or (inputs(81));
    layer0_outputs(2410) <= not(inputs(100)) or (inputs(225));
    layer0_outputs(2411) <= (inputs(160)) and not (inputs(145));
    layer0_outputs(2412) <= not(inputs(171)) or (inputs(93));
    layer0_outputs(2413) <= (inputs(232)) and (inputs(123));
    layer0_outputs(2414) <= not((inputs(188)) xor (inputs(63)));
    layer0_outputs(2415) <= not((inputs(241)) or (inputs(183)));
    layer0_outputs(2416) <= not(inputs(10));
    layer0_outputs(2417) <= inputs(163);
    layer0_outputs(2418) <= not(inputs(230)) or (inputs(116));
    layer0_outputs(2419) <= (inputs(252)) and not (inputs(102));
    layer0_outputs(2420) <= (inputs(79)) or (inputs(9));
    layer0_outputs(2421) <= not(inputs(201));
    layer0_outputs(2422) <= not(inputs(93));
    layer0_outputs(2423) <= inputs(83);
    layer0_outputs(2424) <= '0';
    layer0_outputs(2425) <= inputs(130);
    layer0_outputs(2426) <= (inputs(241)) or (inputs(228));
    layer0_outputs(2427) <= inputs(20);
    layer0_outputs(2428) <= not(inputs(57)) or (inputs(175));
    layer0_outputs(2429) <= not(inputs(20)) or (inputs(189));
    layer0_outputs(2430) <= not(inputs(104));
    layer0_outputs(2431) <= (inputs(128)) or (inputs(82));
    layer0_outputs(2432) <= inputs(249);
    layer0_outputs(2433) <= not((inputs(155)) and (inputs(53)));
    layer0_outputs(2434) <= inputs(20);
    layer0_outputs(2435) <= '1';
    layer0_outputs(2436) <= not(inputs(219));
    layer0_outputs(2437) <= not(inputs(253));
    layer0_outputs(2438) <= not(inputs(19)) or (inputs(15));
    layer0_outputs(2439) <= not(inputs(234));
    layer0_outputs(2440) <= (inputs(171)) xor (inputs(191));
    layer0_outputs(2441) <= not(inputs(83));
    layer0_outputs(2442) <= not(inputs(235));
    layer0_outputs(2443) <= not(inputs(215));
    layer0_outputs(2444) <= (inputs(133)) and not (inputs(141));
    layer0_outputs(2445) <= (inputs(231)) and not (inputs(72));
    layer0_outputs(2446) <= not((inputs(34)) or (inputs(71)));
    layer0_outputs(2447) <= not(inputs(1)) or (inputs(163));
    layer0_outputs(2448) <= inputs(229);
    layer0_outputs(2449) <= inputs(245);
    layer0_outputs(2450) <= not(inputs(154)) or (inputs(202));
    layer0_outputs(2451) <= inputs(91);
    layer0_outputs(2452) <= not((inputs(25)) or (inputs(252)));
    layer0_outputs(2453) <= inputs(98);
    layer0_outputs(2454) <= not(inputs(166)) or (inputs(128));
    layer0_outputs(2455) <= inputs(229);
    layer0_outputs(2456) <= not(inputs(114));
    layer0_outputs(2457) <= '0';
    layer0_outputs(2458) <= '0';
    layer0_outputs(2459) <= not(inputs(195));
    layer0_outputs(2460) <= not(inputs(135)) or (inputs(191));
    layer0_outputs(2461) <= inputs(94);
    layer0_outputs(2462) <= inputs(213);
    layer0_outputs(2463) <= (inputs(120)) or (inputs(239));
    layer0_outputs(2464) <= not(inputs(32));
    layer0_outputs(2465) <= (inputs(122)) xor (inputs(60));
    layer0_outputs(2466) <= not(inputs(162));
    layer0_outputs(2467) <= not((inputs(255)) or (inputs(236)));
    layer0_outputs(2468) <= inputs(117);
    layer0_outputs(2469) <= inputs(179);
    layer0_outputs(2470) <= inputs(197);
    layer0_outputs(2471) <= not(inputs(183)) or (inputs(45));
    layer0_outputs(2472) <= not(inputs(84));
    layer0_outputs(2473) <= not(inputs(103)) or (inputs(163));
    layer0_outputs(2474) <= not(inputs(242)) or (inputs(18));
    layer0_outputs(2475) <= (inputs(66)) and not (inputs(145));
    layer0_outputs(2476) <= (inputs(133)) and not (inputs(46));
    layer0_outputs(2477) <= not(inputs(130));
    layer0_outputs(2478) <= (inputs(85)) and not (inputs(192));
    layer0_outputs(2479) <= inputs(40);
    layer0_outputs(2480) <= not((inputs(188)) and (inputs(243)));
    layer0_outputs(2481) <= (inputs(22)) and not (inputs(233));
    layer0_outputs(2482) <= not((inputs(229)) or (inputs(117)));
    layer0_outputs(2483) <= (inputs(243)) or (inputs(5));
    layer0_outputs(2484) <= (inputs(8)) or (inputs(45));
    layer0_outputs(2485) <= inputs(35);
    layer0_outputs(2486) <= (inputs(59)) or (inputs(107));
    layer0_outputs(2487) <= not((inputs(190)) or (inputs(178)));
    layer0_outputs(2488) <= (inputs(161)) or (inputs(230));
    layer0_outputs(2489) <= not(inputs(241));
    layer0_outputs(2490) <= (inputs(144)) or (inputs(84));
    layer0_outputs(2491) <= not((inputs(152)) or (inputs(180)));
    layer0_outputs(2492) <= not((inputs(222)) or (inputs(184)));
    layer0_outputs(2493) <= not(inputs(101)) or (inputs(253));
    layer0_outputs(2494) <= inputs(17);
    layer0_outputs(2495) <= inputs(87);
    layer0_outputs(2496) <= not(inputs(122)) or (inputs(221));
    layer0_outputs(2497) <= not(inputs(230)) or (inputs(17));
    layer0_outputs(2498) <= not(inputs(83));
    layer0_outputs(2499) <= '0';
    layer0_outputs(2500) <= inputs(86);
    layer0_outputs(2501) <= not(inputs(251)) or (inputs(14));
    layer0_outputs(2502) <= inputs(25);
    layer0_outputs(2503) <= not((inputs(35)) xor (inputs(26)));
    layer0_outputs(2504) <= not(inputs(234));
    layer0_outputs(2505) <= inputs(69);
    layer0_outputs(2506) <= not(inputs(193)) or (inputs(76));
    layer0_outputs(2507) <= not(inputs(110));
    layer0_outputs(2508) <= (inputs(192)) xor (inputs(235));
    layer0_outputs(2509) <= (inputs(182)) or (inputs(4));
    layer0_outputs(2510) <= not(inputs(50));
    layer0_outputs(2511) <= '0';
    layer0_outputs(2512) <= not(inputs(47)) or (inputs(6));
    layer0_outputs(2513) <= not(inputs(9)) or (inputs(222));
    layer0_outputs(2514) <= not(inputs(65));
    layer0_outputs(2515) <= inputs(99);
    layer0_outputs(2516) <= not(inputs(213));
    layer0_outputs(2517) <= inputs(103);
    layer0_outputs(2518) <= (inputs(0)) or (inputs(34));
    layer0_outputs(2519) <= inputs(241);
    layer0_outputs(2520) <= '1';
    layer0_outputs(2521) <= '1';
    layer0_outputs(2522) <= (inputs(210)) and not (inputs(128));
    layer0_outputs(2523) <= not((inputs(43)) xor (inputs(18)));
    layer0_outputs(2524) <= not((inputs(86)) or (inputs(127)));
    layer0_outputs(2525) <= (inputs(171)) or (inputs(212));
    layer0_outputs(2526) <= inputs(226);
    layer0_outputs(2527) <= inputs(230);
    layer0_outputs(2528) <= inputs(211);
    layer0_outputs(2529) <= not((inputs(33)) xor (inputs(49)));
    layer0_outputs(2530) <= not((inputs(217)) or (inputs(167)));
    layer0_outputs(2531) <= not((inputs(53)) or (inputs(173)));
    layer0_outputs(2532) <= not((inputs(135)) xor (inputs(166)));
    layer0_outputs(2533) <= not((inputs(231)) or (inputs(118)));
    layer0_outputs(2534) <= (inputs(58)) and (inputs(48));
    layer0_outputs(2535) <= not(inputs(101));
    layer0_outputs(2536) <= not(inputs(128)) or (inputs(47));
    layer0_outputs(2537) <= (inputs(220)) or (inputs(141));
    layer0_outputs(2538) <= (inputs(84)) or (inputs(164));
    layer0_outputs(2539) <= not(inputs(100));
    layer0_outputs(2540) <= (inputs(10)) or (inputs(51));
    layer0_outputs(2541) <= not(inputs(12)) or (inputs(228));
    layer0_outputs(2542) <= (inputs(244)) xor (inputs(249));
    layer0_outputs(2543) <= not(inputs(184));
    layer0_outputs(2544) <= (inputs(216)) xor (inputs(197));
    layer0_outputs(2545) <= (inputs(116)) or (inputs(34));
    layer0_outputs(2546) <= not(inputs(87)) or (inputs(253));
    layer0_outputs(2547) <= not((inputs(124)) or (inputs(28)));
    layer0_outputs(2548) <= inputs(211);
    layer0_outputs(2549) <= inputs(250);
    layer0_outputs(2550) <= inputs(213);
    layer0_outputs(2551) <= not((inputs(69)) or (inputs(39)));
    layer0_outputs(2552) <= not((inputs(174)) and (inputs(204)));
    layer0_outputs(2553) <= not(inputs(11));
    layer0_outputs(2554) <= not((inputs(86)) or (inputs(140)));
    layer0_outputs(2555) <= not((inputs(236)) xor (inputs(10)));
    layer0_outputs(2556) <= not(inputs(117));
    layer0_outputs(2557) <= '0';
    layer0_outputs(2558) <= not(inputs(51)) or (inputs(51));
    layer0_outputs(2559) <= '1';
    layer0_outputs(2560) <= (inputs(118)) xor (inputs(189));
    layer0_outputs(2561) <= (inputs(165)) xor (inputs(182));
    layer0_outputs(2562) <= not((inputs(214)) xor (inputs(246)));
    layer0_outputs(2563) <= (inputs(136)) or (inputs(169));
    layer0_outputs(2564) <= inputs(122);
    layer0_outputs(2565) <= not(inputs(79));
    layer0_outputs(2566) <= not(inputs(27));
    layer0_outputs(2567) <= inputs(153);
    layer0_outputs(2568) <= (inputs(130)) or (inputs(141));
    layer0_outputs(2569) <= not((inputs(125)) and (inputs(162)));
    layer0_outputs(2570) <= inputs(23);
    layer0_outputs(2571) <= not(inputs(180)) or (inputs(35));
    layer0_outputs(2572) <= not(inputs(144));
    layer0_outputs(2573) <= not(inputs(5));
    layer0_outputs(2574) <= (inputs(95)) and not (inputs(11));
    layer0_outputs(2575) <= not((inputs(68)) xor (inputs(24)));
    layer0_outputs(2576) <= not(inputs(123)) or (inputs(246));
    layer0_outputs(2577) <= (inputs(209)) or (inputs(86));
    layer0_outputs(2578) <= not(inputs(55)) or (inputs(50));
    layer0_outputs(2579) <= not(inputs(193));
    layer0_outputs(2580) <= not(inputs(167)) or (inputs(88));
    layer0_outputs(2581) <= (inputs(185)) or (inputs(98));
    layer0_outputs(2582) <= not(inputs(233)) or (inputs(61));
    layer0_outputs(2583) <= not(inputs(124)) or (inputs(58));
    layer0_outputs(2584) <= (inputs(46)) or (inputs(7));
    layer0_outputs(2585) <= not((inputs(118)) or (inputs(114)));
    layer0_outputs(2586) <= (inputs(24)) and not (inputs(116));
    layer0_outputs(2587) <= not((inputs(39)) xor (inputs(159)));
    layer0_outputs(2588) <= (inputs(4)) xor (inputs(0));
    layer0_outputs(2589) <= not(inputs(101));
    layer0_outputs(2590) <= not(inputs(90)) or (inputs(190));
    layer0_outputs(2591) <= (inputs(136)) xor (inputs(224));
    layer0_outputs(2592) <= inputs(183);
    layer0_outputs(2593) <= (inputs(164)) and not (inputs(224));
    layer0_outputs(2594) <= not((inputs(71)) xor (inputs(25)));
    layer0_outputs(2595) <= not(inputs(230));
    layer0_outputs(2596) <= (inputs(101)) or (inputs(82));
    layer0_outputs(2597) <= not((inputs(252)) or (inputs(14)));
    layer0_outputs(2598) <= (inputs(72)) and not (inputs(139));
    layer0_outputs(2599) <= not((inputs(47)) xor (inputs(234)));
    layer0_outputs(2600) <= (inputs(150)) or (inputs(241));
    layer0_outputs(2601) <= not((inputs(220)) or (inputs(197)));
    layer0_outputs(2602) <= (inputs(27)) and not (inputs(141));
    layer0_outputs(2603) <= (inputs(213)) or (inputs(180));
    layer0_outputs(2604) <= not((inputs(252)) xor (inputs(219)));
    layer0_outputs(2605) <= not(inputs(86));
    layer0_outputs(2606) <= not(inputs(116)) or (inputs(10));
    layer0_outputs(2607) <= not((inputs(37)) and (inputs(22)));
    layer0_outputs(2608) <= not(inputs(37));
    layer0_outputs(2609) <= (inputs(60)) and not (inputs(201));
    layer0_outputs(2610) <= (inputs(205)) and not (inputs(148));
    layer0_outputs(2611) <= inputs(100);
    layer0_outputs(2612) <= (inputs(237)) or (inputs(72));
    layer0_outputs(2613) <= not((inputs(219)) xor (inputs(216)));
    layer0_outputs(2614) <= not(inputs(19));
    layer0_outputs(2615) <= (inputs(138)) and not (inputs(178));
    layer0_outputs(2616) <= not(inputs(28));
    layer0_outputs(2617) <= not(inputs(119));
    layer0_outputs(2618) <= not(inputs(145)) or (inputs(208));
    layer0_outputs(2619) <= (inputs(81)) or (inputs(76));
    layer0_outputs(2620) <= not(inputs(168)) or (inputs(116));
    layer0_outputs(2621) <= inputs(19);
    layer0_outputs(2622) <= (inputs(88)) xor (inputs(139));
    layer0_outputs(2623) <= (inputs(39)) xor (inputs(62));
    layer0_outputs(2624) <= (inputs(48)) and not (inputs(251));
    layer0_outputs(2625) <= inputs(215);
    layer0_outputs(2626) <= not((inputs(187)) or (inputs(159)));
    layer0_outputs(2627) <= not(inputs(87)) or (inputs(181));
    layer0_outputs(2628) <= not(inputs(54));
    layer0_outputs(2629) <= not(inputs(213));
    layer0_outputs(2630) <= not(inputs(189));
    layer0_outputs(2631) <= not(inputs(64)) or (inputs(28));
    layer0_outputs(2632) <= (inputs(144)) and not (inputs(7));
    layer0_outputs(2633) <= inputs(246);
    layer0_outputs(2634) <= inputs(23);
    layer0_outputs(2635) <= not((inputs(148)) or (inputs(88)));
    layer0_outputs(2636) <= inputs(99);
    layer0_outputs(2637) <= not((inputs(219)) or (inputs(110)));
    layer0_outputs(2638) <= not(inputs(255)) or (inputs(254));
    layer0_outputs(2639) <= inputs(23);
    layer0_outputs(2640) <= inputs(228);
    layer0_outputs(2641) <= not(inputs(26));
    layer0_outputs(2642) <= not(inputs(74)) or (inputs(206));
    layer0_outputs(2643) <= not(inputs(204));
    layer0_outputs(2644) <= inputs(152);
    layer0_outputs(2645) <= not(inputs(147)) or (inputs(148));
    layer0_outputs(2646) <= not(inputs(163));
    layer0_outputs(2647) <= '1';
    layer0_outputs(2648) <= inputs(221);
    layer0_outputs(2649) <= not((inputs(20)) or (inputs(54)));
    layer0_outputs(2650) <= inputs(234);
    layer0_outputs(2651) <= (inputs(106)) xor (inputs(204));
    layer0_outputs(2652) <= (inputs(149)) and not (inputs(63));
    layer0_outputs(2653) <= not(inputs(87));
    layer0_outputs(2654) <= not(inputs(75));
    layer0_outputs(2655) <= not((inputs(223)) or (inputs(229)));
    layer0_outputs(2656) <= (inputs(117)) and not (inputs(72));
    layer0_outputs(2657) <= not(inputs(168)) or (inputs(99));
    layer0_outputs(2658) <= inputs(246);
    layer0_outputs(2659) <= (inputs(47)) or (inputs(34));
    layer0_outputs(2660) <= '0';
    layer0_outputs(2661) <= not(inputs(177)) or (inputs(112));
    layer0_outputs(2662) <= (inputs(195)) or (inputs(141));
    layer0_outputs(2663) <= not(inputs(21)) or (inputs(200));
    layer0_outputs(2664) <= inputs(156);
    layer0_outputs(2665) <= not(inputs(193));
    layer0_outputs(2666) <= inputs(203);
    layer0_outputs(2667) <= not(inputs(165)) or (inputs(97));
    layer0_outputs(2668) <= (inputs(11)) and not (inputs(238));
    layer0_outputs(2669) <= not(inputs(188));
    layer0_outputs(2670) <= (inputs(38)) or (inputs(97));
    layer0_outputs(2671) <= (inputs(227)) and (inputs(202));
    layer0_outputs(2672) <= (inputs(69)) and not (inputs(20));
    layer0_outputs(2673) <= not(inputs(10));
    layer0_outputs(2674) <= not((inputs(72)) xor (inputs(61)));
    layer0_outputs(2675) <= not(inputs(119));
    layer0_outputs(2676) <= not((inputs(160)) or (inputs(208)));
    layer0_outputs(2677) <= not(inputs(182)) or (inputs(37));
    layer0_outputs(2678) <= inputs(87);
    layer0_outputs(2679) <= not((inputs(111)) or (inputs(112)));
    layer0_outputs(2680) <= (inputs(116)) and not (inputs(156));
    layer0_outputs(2681) <= not(inputs(94));
    layer0_outputs(2682) <= (inputs(181)) or (inputs(33));
    layer0_outputs(2683) <= not(inputs(60));
    layer0_outputs(2684) <= not((inputs(14)) or (inputs(99)));
    layer0_outputs(2685) <= not(inputs(189)) or (inputs(63));
    layer0_outputs(2686) <= inputs(26);
    layer0_outputs(2687) <= inputs(210);
    layer0_outputs(2688) <= not(inputs(27)) or (inputs(242));
    layer0_outputs(2689) <= (inputs(76)) or (inputs(139));
    layer0_outputs(2690) <= (inputs(218)) and not (inputs(130));
    layer0_outputs(2691) <= (inputs(161)) and not (inputs(47));
    layer0_outputs(2692) <= (inputs(186)) xor (inputs(235));
    layer0_outputs(2693) <= not(inputs(153));
    layer0_outputs(2694) <= not(inputs(203));
    layer0_outputs(2695) <= inputs(84);
    layer0_outputs(2696) <= (inputs(97)) xor (inputs(177));
    layer0_outputs(2697) <= not((inputs(168)) or (inputs(46)));
    layer0_outputs(2698) <= inputs(92);
    layer0_outputs(2699) <= not((inputs(126)) xor (inputs(217)));
    layer0_outputs(2700) <= (inputs(172)) or (inputs(147));
    layer0_outputs(2701) <= (inputs(101)) or (inputs(114));
    layer0_outputs(2702) <= (inputs(191)) or (inputs(141));
    layer0_outputs(2703) <= (inputs(72)) and not (inputs(62));
    layer0_outputs(2704) <= not(inputs(152)) or (inputs(131));
    layer0_outputs(2705) <= (inputs(114)) or (inputs(192));
    layer0_outputs(2706) <= (inputs(228)) and not (inputs(35));
    layer0_outputs(2707) <= not((inputs(175)) and (inputs(241)));
    layer0_outputs(2708) <= (inputs(145)) and not (inputs(80));
    layer0_outputs(2709) <= not(inputs(26)) or (inputs(186));
    layer0_outputs(2710) <= not((inputs(193)) xor (inputs(172)));
    layer0_outputs(2711) <= not((inputs(34)) or (inputs(9)));
    layer0_outputs(2712) <= not(inputs(44));
    layer0_outputs(2713) <= not(inputs(25));
    layer0_outputs(2714) <= (inputs(203)) or (inputs(137));
    layer0_outputs(2715) <= not(inputs(149));
    layer0_outputs(2716) <= not((inputs(191)) or (inputs(38)));
    layer0_outputs(2717) <= (inputs(230)) or (inputs(190));
    layer0_outputs(2718) <= not((inputs(135)) or (inputs(214)));
    layer0_outputs(2719) <= inputs(126);
    layer0_outputs(2720) <= '1';
    layer0_outputs(2721) <= (inputs(106)) and not (inputs(103));
    layer0_outputs(2722) <= (inputs(85)) or (inputs(203));
    layer0_outputs(2723) <= not((inputs(225)) or (inputs(19)));
    layer0_outputs(2724) <= not(inputs(116));
    layer0_outputs(2725) <= not((inputs(126)) or (inputs(18)));
    layer0_outputs(2726) <= '1';
    layer0_outputs(2727) <= not(inputs(42));
    layer0_outputs(2728) <= (inputs(188)) and not (inputs(88));
    layer0_outputs(2729) <= inputs(183);
    layer0_outputs(2730) <= (inputs(94)) or (inputs(130));
    layer0_outputs(2731) <= not((inputs(30)) xor (inputs(242)));
    layer0_outputs(2732) <= not((inputs(33)) xor (inputs(70)));
    layer0_outputs(2733) <= not((inputs(54)) or (inputs(4)));
    layer0_outputs(2734) <= not((inputs(233)) xor (inputs(255)));
    layer0_outputs(2735) <= not((inputs(11)) or (inputs(139)));
    layer0_outputs(2736) <= not(inputs(136));
    layer0_outputs(2737) <= inputs(137);
    layer0_outputs(2738) <= '1';
    layer0_outputs(2739) <= (inputs(14)) or (inputs(190));
    layer0_outputs(2740) <= not(inputs(101)) or (inputs(190));
    layer0_outputs(2741) <= not(inputs(215));
    layer0_outputs(2742) <= inputs(145);
    layer0_outputs(2743) <= inputs(247);
    layer0_outputs(2744) <= inputs(116);
    layer0_outputs(2745) <= not(inputs(173)) or (inputs(76));
    layer0_outputs(2746) <= not((inputs(129)) xor (inputs(100)));
    layer0_outputs(2747) <= inputs(174);
    layer0_outputs(2748) <= inputs(73);
    layer0_outputs(2749) <= not(inputs(227));
    layer0_outputs(2750) <= (inputs(247)) and not (inputs(6));
    layer0_outputs(2751) <= (inputs(56)) and not (inputs(111));
    layer0_outputs(2752) <= not(inputs(9));
    layer0_outputs(2753) <= inputs(180);
    layer0_outputs(2754) <= not(inputs(183));
    layer0_outputs(2755) <= (inputs(234)) xor (inputs(195));
    layer0_outputs(2756) <= not(inputs(210)) or (inputs(14));
    layer0_outputs(2757) <= not((inputs(236)) or (inputs(218)));
    layer0_outputs(2758) <= (inputs(180)) or (inputs(176));
    layer0_outputs(2759) <= (inputs(7)) or (inputs(76));
    layer0_outputs(2760) <= (inputs(61)) or (inputs(90));
    layer0_outputs(2761) <= '0';
    layer0_outputs(2762) <= (inputs(138)) and not (inputs(234));
    layer0_outputs(2763) <= (inputs(118)) xor (inputs(3));
    layer0_outputs(2764) <= not((inputs(133)) xor (inputs(50)));
    layer0_outputs(2765) <= not((inputs(226)) or (inputs(34)));
    layer0_outputs(2766) <= (inputs(34)) or (inputs(119));
    layer0_outputs(2767) <= not(inputs(204)) or (inputs(63));
    layer0_outputs(2768) <= not((inputs(122)) or (inputs(28)));
    layer0_outputs(2769) <= not(inputs(103)) or (inputs(93));
    layer0_outputs(2770) <= not((inputs(115)) or (inputs(236)));
    layer0_outputs(2771) <= (inputs(84)) or (inputs(253));
    layer0_outputs(2772) <= (inputs(98)) or (inputs(103));
    layer0_outputs(2773) <= (inputs(95)) or (inputs(207));
    layer0_outputs(2774) <= not(inputs(105));
    layer0_outputs(2775) <= inputs(148);
    layer0_outputs(2776) <= inputs(247);
    layer0_outputs(2777) <= inputs(181);
    layer0_outputs(2778) <= not((inputs(233)) xor (inputs(184)));
    layer0_outputs(2779) <= '0';
    layer0_outputs(2780) <= not((inputs(38)) or (inputs(96)));
    layer0_outputs(2781) <= not(inputs(225));
    layer0_outputs(2782) <= inputs(221);
    layer0_outputs(2783) <= (inputs(27)) and (inputs(53));
    layer0_outputs(2784) <= inputs(119);
    layer0_outputs(2785) <= not(inputs(169));
    layer0_outputs(2786) <= not((inputs(36)) and (inputs(200)));
    layer0_outputs(2787) <= not(inputs(203));
    layer0_outputs(2788) <= (inputs(8)) and not (inputs(7));
    layer0_outputs(2789) <= not(inputs(234)) or (inputs(72));
    layer0_outputs(2790) <= not(inputs(152)) or (inputs(114));
    layer0_outputs(2791) <= (inputs(127)) or (inputs(140));
    layer0_outputs(2792) <= not(inputs(174));
    layer0_outputs(2793) <= (inputs(94)) and not (inputs(40));
    layer0_outputs(2794) <= '1';
    layer0_outputs(2795) <= '1';
    layer0_outputs(2796) <= not((inputs(92)) xor (inputs(49)));
    layer0_outputs(2797) <= not(inputs(114));
    layer0_outputs(2798) <= inputs(179);
    layer0_outputs(2799) <= (inputs(135)) and not (inputs(6));
    layer0_outputs(2800) <= not(inputs(251)) or (inputs(62));
    layer0_outputs(2801) <= (inputs(88)) and not (inputs(22));
    layer0_outputs(2802) <= inputs(106);
    layer0_outputs(2803) <= (inputs(203)) xor (inputs(209));
    layer0_outputs(2804) <= inputs(162);
    layer0_outputs(2805) <= inputs(55);
    layer0_outputs(2806) <= not((inputs(178)) or (inputs(145)));
    layer0_outputs(2807) <= (inputs(9)) and not (inputs(208));
    layer0_outputs(2808) <= (inputs(132)) and not (inputs(108));
    layer0_outputs(2809) <= not(inputs(177));
    layer0_outputs(2810) <= (inputs(217)) or (inputs(31));
    layer0_outputs(2811) <= not((inputs(71)) or (inputs(177)));
    layer0_outputs(2812) <= not(inputs(177));
    layer0_outputs(2813) <= inputs(213);
    layer0_outputs(2814) <= (inputs(251)) and (inputs(192));
    layer0_outputs(2815) <= (inputs(208)) and not (inputs(68));
    layer0_outputs(2816) <= not((inputs(146)) or (inputs(51)));
    layer0_outputs(2817) <= not(inputs(165));
    layer0_outputs(2818) <= not(inputs(139));
    layer0_outputs(2819) <= inputs(186);
    layer0_outputs(2820) <= inputs(146);
    layer0_outputs(2821) <= inputs(99);
    layer0_outputs(2822) <= (inputs(34)) and (inputs(168));
    layer0_outputs(2823) <= inputs(24);
    layer0_outputs(2824) <= inputs(183);
    layer0_outputs(2825) <= not((inputs(89)) or (inputs(120)));
    layer0_outputs(2826) <= inputs(131);
    layer0_outputs(2827) <= not(inputs(136)) or (inputs(127));
    layer0_outputs(2828) <= not(inputs(191));
    layer0_outputs(2829) <= not(inputs(87)) or (inputs(174));
    layer0_outputs(2830) <= (inputs(38)) and not (inputs(159));
    layer0_outputs(2831) <= not(inputs(20));
    layer0_outputs(2832) <= not(inputs(11)) or (inputs(220));
    layer0_outputs(2833) <= not((inputs(239)) xor (inputs(115)));
    layer0_outputs(2834) <= not(inputs(155));
    layer0_outputs(2835) <= not((inputs(231)) and (inputs(172)));
    layer0_outputs(2836) <= not(inputs(147));
    layer0_outputs(2837) <= inputs(162);
    layer0_outputs(2838) <= (inputs(77)) and not (inputs(130));
    layer0_outputs(2839) <= inputs(151);
    layer0_outputs(2840) <= inputs(210);
    layer0_outputs(2841) <= (inputs(118)) and not (inputs(112));
    layer0_outputs(2842) <= not(inputs(198));
    layer0_outputs(2843) <= (inputs(64)) or (inputs(35));
    layer0_outputs(2844) <= not(inputs(90));
    layer0_outputs(2845) <= (inputs(165)) xor (inputs(0));
    layer0_outputs(2846) <= not((inputs(192)) or (inputs(110)));
    layer0_outputs(2847) <= inputs(180);
    layer0_outputs(2848) <= (inputs(228)) or (inputs(66));
    layer0_outputs(2849) <= not((inputs(83)) xor (inputs(191)));
    layer0_outputs(2850) <= not((inputs(79)) or (inputs(221)));
    layer0_outputs(2851) <= not((inputs(33)) and (inputs(192)));
    layer0_outputs(2852) <= inputs(135);
    layer0_outputs(2853) <= not(inputs(243));
    layer0_outputs(2854) <= not(inputs(58));
    layer0_outputs(2855) <= (inputs(62)) xor (inputs(96));
    layer0_outputs(2856) <= '0';
    layer0_outputs(2857) <= not(inputs(25)) or (inputs(246));
    layer0_outputs(2858) <= (inputs(70)) or (inputs(69));
    layer0_outputs(2859) <= not(inputs(146));
    layer0_outputs(2860) <= (inputs(36)) or (inputs(52));
    layer0_outputs(2861) <= not(inputs(178)) or (inputs(248));
    layer0_outputs(2862) <= not((inputs(167)) or (inputs(104)));
    layer0_outputs(2863) <= (inputs(142)) or (inputs(172));
    layer0_outputs(2864) <= not(inputs(229));
    layer0_outputs(2865) <= not(inputs(9)) or (inputs(113));
    layer0_outputs(2866) <= not((inputs(4)) xor (inputs(135)));
    layer0_outputs(2867) <= (inputs(48)) and (inputs(239));
    layer0_outputs(2868) <= (inputs(12)) and (inputs(16));
    layer0_outputs(2869) <= inputs(242);
    layer0_outputs(2870) <= not(inputs(187));
    layer0_outputs(2871) <= (inputs(153)) and not (inputs(189));
    layer0_outputs(2872) <= not(inputs(83));
    layer0_outputs(2873) <= inputs(62);
    layer0_outputs(2874) <= (inputs(101)) and not (inputs(239));
    layer0_outputs(2875) <= (inputs(164)) or (inputs(179));
    layer0_outputs(2876) <= not(inputs(162));
    layer0_outputs(2877) <= not((inputs(176)) or (inputs(164)));
    layer0_outputs(2878) <= inputs(129);
    layer0_outputs(2879) <= not(inputs(178));
    layer0_outputs(2880) <= (inputs(187)) xor (inputs(138));
    layer0_outputs(2881) <= inputs(25);
    layer0_outputs(2882) <= inputs(230);
    layer0_outputs(2883) <= inputs(24);
    layer0_outputs(2884) <= inputs(29);
    layer0_outputs(2885) <= not(inputs(22));
    layer0_outputs(2886) <= (inputs(167)) or (inputs(151));
    layer0_outputs(2887) <= (inputs(24)) or (inputs(5));
    layer0_outputs(2888) <= inputs(121);
    layer0_outputs(2889) <= (inputs(160)) xor (inputs(176));
    layer0_outputs(2890) <= (inputs(128)) and not (inputs(47));
    layer0_outputs(2891) <= not(inputs(170));
    layer0_outputs(2892) <= (inputs(86)) and not (inputs(57));
    layer0_outputs(2893) <= not(inputs(162)) or (inputs(192));
    layer0_outputs(2894) <= not(inputs(229));
    layer0_outputs(2895) <= not((inputs(55)) xor (inputs(43)));
    layer0_outputs(2896) <= (inputs(253)) and not (inputs(78));
    layer0_outputs(2897) <= inputs(73);
    layer0_outputs(2898) <= not(inputs(198));
    layer0_outputs(2899) <= not(inputs(51));
    layer0_outputs(2900) <= not(inputs(9)) or (inputs(227));
    layer0_outputs(2901) <= inputs(7);
    layer0_outputs(2902) <= (inputs(136)) and not (inputs(234));
    layer0_outputs(2903) <= not((inputs(156)) or (inputs(31)));
    layer0_outputs(2904) <= not((inputs(8)) or (inputs(113)));
    layer0_outputs(2905) <= (inputs(23)) or (inputs(51));
    layer0_outputs(2906) <= not(inputs(136)) or (inputs(48));
    layer0_outputs(2907) <= (inputs(112)) and not (inputs(36));
    layer0_outputs(2908) <= inputs(244);
    layer0_outputs(2909) <= not((inputs(241)) xor (inputs(72)));
    layer0_outputs(2910) <= not(inputs(152));
    layer0_outputs(2911) <= inputs(227);
    layer0_outputs(2912) <= not(inputs(171));
    layer0_outputs(2913) <= (inputs(132)) or (inputs(101));
    layer0_outputs(2914) <= (inputs(6)) or (inputs(164));
    layer0_outputs(2915) <= not((inputs(111)) xor (inputs(181)));
    layer0_outputs(2916) <= not(inputs(104));
    layer0_outputs(2917) <= inputs(147);
    layer0_outputs(2918) <= not(inputs(254));
    layer0_outputs(2919) <= inputs(68);
    layer0_outputs(2920) <= not(inputs(72));
    layer0_outputs(2921) <= (inputs(200)) and not (inputs(134));
    layer0_outputs(2922) <= '1';
    layer0_outputs(2923) <= not(inputs(105));
    layer0_outputs(2924) <= not(inputs(111));
    layer0_outputs(2925) <= not(inputs(227));
    layer0_outputs(2926) <= not(inputs(150));
    layer0_outputs(2927) <= '1';
    layer0_outputs(2928) <= inputs(229);
    layer0_outputs(2929) <= (inputs(247)) xor (inputs(216));
    layer0_outputs(2930) <= not(inputs(97));
    layer0_outputs(2931) <= not(inputs(18));
    layer0_outputs(2932) <= (inputs(204)) and not (inputs(109));
    layer0_outputs(2933) <= not((inputs(237)) or (inputs(157)));
    layer0_outputs(2934) <= not((inputs(80)) or (inputs(132)));
    layer0_outputs(2935) <= (inputs(226)) and not (inputs(1));
    layer0_outputs(2936) <= inputs(102);
    layer0_outputs(2937) <= not(inputs(38));
    layer0_outputs(2938) <= not(inputs(203));
    layer0_outputs(2939) <= not(inputs(164)) or (inputs(172));
    layer0_outputs(2940) <= (inputs(237)) or (inputs(30));
    layer0_outputs(2941) <= not((inputs(171)) xor (inputs(175)));
    layer0_outputs(2942) <= inputs(52);
    layer0_outputs(2943) <= (inputs(233)) and not (inputs(126));
    layer0_outputs(2944) <= (inputs(203)) and (inputs(96));
    layer0_outputs(2945) <= (inputs(78)) xor (inputs(11));
    layer0_outputs(2946) <= (inputs(163)) and not (inputs(44));
    layer0_outputs(2947) <= (inputs(5)) xor (inputs(143));
    layer0_outputs(2948) <= (inputs(54)) or (inputs(80));
    layer0_outputs(2949) <= not((inputs(50)) and (inputs(235)));
    layer0_outputs(2950) <= inputs(151);
    layer0_outputs(2951) <= inputs(167);
    layer0_outputs(2952) <= not((inputs(66)) xor (inputs(202)));
    layer0_outputs(2953) <= (inputs(29)) xor (inputs(255));
    layer0_outputs(2954) <= not(inputs(248)) or (inputs(248));
    layer0_outputs(2955) <= (inputs(73)) and not (inputs(171));
    layer0_outputs(2956) <= inputs(40);
    layer0_outputs(2957) <= inputs(6);
    layer0_outputs(2958) <= not(inputs(174));
    layer0_outputs(2959) <= (inputs(11)) or (inputs(187));
    layer0_outputs(2960) <= (inputs(143)) and not (inputs(157));
    layer0_outputs(2961) <= not(inputs(123));
    layer0_outputs(2962) <= (inputs(73)) xor (inputs(194));
    layer0_outputs(2963) <= not((inputs(230)) and (inputs(217)));
    layer0_outputs(2964) <= inputs(194);
    layer0_outputs(2965) <= not((inputs(161)) and (inputs(253)));
    layer0_outputs(2966) <= inputs(116);
    layer0_outputs(2967) <= inputs(55);
    layer0_outputs(2968) <= not((inputs(105)) xor (inputs(152)));
    layer0_outputs(2969) <= not((inputs(29)) xor (inputs(248)));
    layer0_outputs(2970) <= (inputs(253)) or (inputs(183));
    layer0_outputs(2971) <= (inputs(157)) or (inputs(99));
    layer0_outputs(2972) <= (inputs(23)) and not (inputs(30));
    layer0_outputs(2973) <= inputs(6);
    layer0_outputs(2974) <= not((inputs(29)) or (inputs(51)));
    layer0_outputs(2975) <= (inputs(188)) or (inputs(207));
    layer0_outputs(2976) <= (inputs(92)) and not (inputs(254));
    layer0_outputs(2977) <= not((inputs(237)) or (inputs(160)));
    layer0_outputs(2978) <= (inputs(56)) or (inputs(159));
    layer0_outputs(2979) <= not(inputs(140)) or (inputs(48));
    layer0_outputs(2980) <= not((inputs(189)) or (inputs(233)));
    layer0_outputs(2981) <= not(inputs(175)) or (inputs(3));
    layer0_outputs(2982) <= not((inputs(16)) xor (inputs(221)));
    layer0_outputs(2983) <= (inputs(77)) or (inputs(48));
    layer0_outputs(2984) <= not(inputs(232));
    layer0_outputs(2985) <= (inputs(79)) xor (inputs(2));
    layer0_outputs(2986) <= not(inputs(37));
    layer0_outputs(2987) <= inputs(127);
    layer0_outputs(2988) <= not(inputs(178));
    layer0_outputs(2989) <= not((inputs(11)) or (inputs(56)));
    layer0_outputs(2990) <= not((inputs(255)) or (inputs(159)));
    layer0_outputs(2991) <= inputs(120);
    layer0_outputs(2992) <= not(inputs(25));
    layer0_outputs(2993) <= not((inputs(212)) or (inputs(172)));
    layer0_outputs(2994) <= (inputs(104)) and not (inputs(50));
    layer0_outputs(2995) <= (inputs(218)) or (inputs(97));
    layer0_outputs(2996) <= not(inputs(86)) or (inputs(242));
    layer0_outputs(2997) <= not(inputs(156));
    layer0_outputs(2998) <= (inputs(134)) or (inputs(134));
    layer0_outputs(2999) <= (inputs(128)) xor (inputs(119));
    layer0_outputs(3000) <= inputs(118);
    layer0_outputs(3001) <= not(inputs(69)) or (inputs(12));
    layer0_outputs(3002) <= not(inputs(219));
    layer0_outputs(3003) <= '1';
    layer0_outputs(3004) <= inputs(230);
    layer0_outputs(3005) <= (inputs(29)) xor (inputs(93));
    layer0_outputs(3006) <= not(inputs(229));
    layer0_outputs(3007) <= (inputs(146)) and not (inputs(64));
    layer0_outputs(3008) <= (inputs(52)) or (inputs(112));
    layer0_outputs(3009) <= not((inputs(55)) or (inputs(93)));
    layer0_outputs(3010) <= not(inputs(94));
    layer0_outputs(3011) <= (inputs(26)) and not (inputs(206));
    layer0_outputs(3012) <= inputs(238);
    layer0_outputs(3013) <= not(inputs(136)) or (inputs(47));
    layer0_outputs(3014) <= not(inputs(194)) or (inputs(223));
    layer0_outputs(3015) <= not(inputs(146));
    layer0_outputs(3016) <= '0';
    layer0_outputs(3017) <= (inputs(182)) or (inputs(177));
    layer0_outputs(3018) <= not(inputs(233));
    layer0_outputs(3019) <= (inputs(87)) or (inputs(92));
    layer0_outputs(3020) <= not(inputs(209));
    layer0_outputs(3021) <= (inputs(232)) and not (inputs(33));
    layer0_outputs(3022) <= not((inputs(149)) or (inputs(6)));
    layer0_outputs(3023) <= (inputs(56)) xor (inputs(222));
    layer0_outputs(3024) <= (inputs(208)) and (inputs(165));
    layer0_outputs(3025) <= inputs(166);
    layer0_outputs(3026) <= not(inputs(104)) or (inputs(22));
    layer0_outputs(3027) <= (inputs(254)) or (inputs(157));
    layer0_outputs(3028) <= not(inputs(166)) or (inputs(238));
    layer0_outputs(3029) <= not((inputs(126)) or (inputs(49)));
    layer0_outputs(3030) <= not(inputs(137));
    layer0_outputs(3031) <= (inputs(196)) and not (inputs(109));
    layer0_outputs(3032) <= not(inputs(159)) or (inputs(61));
    layer0_outputs(3033) <= inputs(22);
    layer0_outputs(3034) <= (inputs(40)) and not (inputs(239));
    layer0_outputs(3035) <= (inputs(69)) or (inputs(30));
    layer0_outputs(3036) <= not(inputs(29)) or (inputs(76));
    layer0_outputs(3037) <= (inputs(95)) and not (inputs(222));
    layer0_outputs(3038) <= (inputs(116)) or (inputs(244));
    layer0_outputs(3039) <= not(inputs(122)) or (inputs(81));
    layer0_outputs(3040) <= not((inputs(83)) or (inputs(94)));
    layer0_outputs(3041) <= inputs(233);
    layer0_outputs(3042) <= (inputs(68)) and not (inputs(49));
    layer0_outputs(3043) <= not(inputs(108));
    layer0_outputs(3044) <= (inputs(138)) or (inputs(22));
    layer0_outputs(3045) <= (inputs(162)) and not (inputs(94));
    layer0_outputs(3046) <= inputs(233);
    layer0_outputs(3047) <= (inputs(122)) and (inputs(151));
    layer0_outputs(3048) <= not((inputs(69)) or (inputs(142)));
    layer0_outputs(3049) <= not(inputs(218)) or (inputs(40));
    layer0_outputs(3050) <= not(inputs(44));
    layer0_outputs(3051) <= (inputs(115)) or (inputs(114));
    layer0_outputs(3052) <= not((inputs(86)) and (inputs(207)));
    layer0_outputs(3053) <= (inputs(26)) xor (inputs(223));
    layer0_outputs(3054) <= not(inputs(121)) or (inputs(144));
    layer0_outputs(3055) <= (inputs(96)) xor (inputs(81));
    layer0_outputs(3056) <= (inputs(193)) or (inputs(162));
    layer0_outputs(3057) <= not((inputs(157)) and (inputs(172)));
    layer0_outputs(3058) <= inputs(85);
    layer0_outputs(3059) <= '1';
    layer0_outputs(3060) <= (inputs(107)) or (inputs(46));
    layer0_outputs(3061) <= inputs(157);
    layer0_outputs(3062) <= not((inputs(64)) or (inputs(198)));
    layer0_outputs(3063) <= (inputs(235)) xor (inputs(130));
    layer0_outputs(3064) <= (inputs(49)) and not (inputs(47));
    layer0_outputs(3065) <= not((inputs(180)) or (inputs(187)));
    layer0_outputs(3066) <= inputs(232);
    layer0_outputs(3067) <= (inputs(106)) and not (inputs(48));
    layer0_outputs(3068) <= not(inputs(173));
    layer0_outputs(3069) <= (inputs(240)) or (inputs(129));
    layer0_outputs(3070) <= not((inputs(143)) xor (inputs(156)));
    layer0_outputs(3071) <= (inputs(3)) or (inputs(35));
    layer0_outputs(3072) <= inputs(196);
    layer0_outputs(3073) <= (inputs(179)) or (inputs(215));
    layer0_outputs(3074) <= inputs(117);
    layer0_outputs(3075) <= not((inputs(4)) or (inputs(2)));
    layer0_outputs(3076) <= '1';
    layer0_outputs(3077) <= (inputs(31)) and (inputs(197));
    layer0_outputs(3078) <= inputs(43);
    layer0_outputs(3079) <= not(inputs(82));
    layer0_outputs(3080) <= inputs(25);
    layer0_outputs(3081) <= not(inputs(243)) or (inputs(240));
    layer0_outputs(3082) <= inputs(197);
    layer0_outputs(3083) <= inputs(233);
    layer0_outputs(3084) <= not(inputs(44));
    layer0_outputs(3085) <= not(inputs(149));
    layer0_outputs(3086) <= inputs(120);
    layer0_outputs(3087) <= (inputs(69)) or (inputs(45));
    layer0_outputs(3088) <= not((inputs(53)) and (inputs(29)));
    layer0_outputs(3089) <= not(inputs(167));
    layer0_outputs(3090) <= (inputs(62)) and (inputs(90));
    layer0_outputs(3091) <= (inputs(123)) xor (inputs(189));
    layer0_outputs(3092) <= inputs(147);
    layer0_outputs(3093) <= not(inputs(144)) or (inputs(55));
    layer0_outputs(3094) <= not(inputs(167)) or (inputs(160));
    layer0_outputs(3095) <= (inputs(235)) or (inputs(198));
    layer0_outputs(3096) <= (inputs(84)) or (inputs(163));
    layer0_outputs(3097) <= (inputs(168)) and not (inputs(31));
    layer0_outputs(3098) <= inputs(179);
    layer0_outputs(3099) <= not(inputs(216));
    layer0_outputs(3100) <= (inputs(49)) or (inputs(33));
    layer0_outputs(3101) <= (inputs(225)) and not (inputs(61));
    layer0_outputs(3102) <= not(inputs(28));
    layer0_outputs(3103) <= not(inputs(189));
    layer0_outputs(3104) <= (inputs(134)) xor (inputs(184));
    layer0_outputs(3105) <= inputs(103);
    layer0_outputs(3106) <= not((inputs(42)) or (inputs(42)));
    layer0_outputs(3107) <= inputs(205);
    layer0_outputs(3108) <= not((inputs(101)) or (inputs(116)));
    layer0_outputs(3109) <= inputs(71);
    layer0_outputs(3110) <= not(inputs(187));
    layer0_outputs(3111) <= (inputs(230)) and not (inputs(98));
    layer0_outputs(3112) <= inputs(115);
    layer0_outputs(3113) <= not(inputs(150));
    layer0_outputs(3114) <= (inputs(151)) or (inputs(183));
    layer0_outputs(3115) <= (inputs(123)) and (inputs(66));
    layer0_outputs(3116) <= not(inputs(139));
    layer0_outputs(3117) <= not(inputs(45)) or (inputs(105));
    layer0_outputs(3118) <= not(inputs(220)) or (inputs(66));
    layer0_outputs(3119) <= not(inputs(86));
    layer0_outputs(3120) <= not((inputs(5)) or (inputs(188)));
    layer0_outputs(3121) <= (inputs(100)) and not (inputs(100));
    layer0_outputs(3122) <= inputs(163);
    layer0_outputs(3123) <= not((inputs(143)) xor (inputs(77)));
    layer0_outputs(3124) <= (inputs(159)) xor (inputs(221));
    layer0_outputs(3125) <= (inputs(246)) and not (inputs(7));
    layer0_outputs(3126) <= not(inputs(137)) or (inputs(16));
    layer0_outputs(3127) <= (inputs(24)) and not (inputs(218));
    layer0_outputs(3128) <= not(inputs(222));
    layer0_outputs(3129) <= not((inputs(28)) or (inputs(171)));
    layer0_outputs(3130) <= (inputs(21)) xor (inputs(193));
    layer0_outputs(3131) <= (inputs(145)) and not (inputs(45));
    layer0_outputs(3132) <= not(inputs(106));
    layer0_outputs(3133) <= (inputs(37)) and not (inputs(53));
    layer0_outputs(3134) <= not(inputs(101));
    layer0_outputs(3135) <= not(inputs(179));
    layer0_outputs(3136) <= not((inputs(255)) or (inputs(108)));
    layer0_outputs(3137) <= not(inputs(120)) or (inputs(203));
    layer0_outputs(3138) <= not(inputs(148));
    layer0_outputs(3139) <= not(inputs(28)) or (inputs(234));
    layer0_outputs(3140) <= not(inputs(85));
    layer0_outputs(3141) <= not((inputs(122)) xor (inputs(172)));
    layer0_outputs(3142) <= not(inputs(207));
    layer0_outputs(3143) <= not((inputs(14)) or (inputs(196)));
    layer0_outputs(3144) <= not((inputs(38)) xor (inputs(1)));
    layer0_outputs(3145) <= inputs(8);
    layer0_outputs(3146) <= not(inputs(1));
    layer0_outputs(3147) <= not(inputs(171)) or (inputs(65));
    layer0_outputs(3148) <= not(inputs(22)) or (inputs(222));
    layer0_outputs(3149) <= (inputs(122)) and not (inputs(203));
    layer0_outputs(3150) <= (inputs(165)) and not (inputs(214));
    layer0_outputs(3151) <= inputs(170);
    layer0_outputs(3152) <= (inputs(82)) or (inputs(29));
    layer0_outputs(3153) <= not(inputs(94)) or (inputs(139));
    layer0_outputs(3154) <= not(inputs(104));
    layer0_outputs(3155) <= not(inputs(182));
    layer0_outputs(3156) <= (inputs(128)) xor (inputs(165));
    layer0_outputs(3157) <= not(inputs(164));
    layer0_outputs(3158) <= not(inputs(225)) or (inputs(159));
    layer0_outputs(3159) <= (inputs(31)) xor (inputs(254));
    layer0_outputs(3160) <= not((inputs(117)) or (inputs(130)));
    layer0_outputs(3161) <= inputs(97);
    layer0_outputs(3162) <= (inputs(165)) and not (inputs(254));
    layer0_outputs(3163) <= not(inputs(140)) or (inputs(63));
    layer0_outputs(3164) <= (inputs(90)) and not (inputs(19));
    layer0_outputs(3165) <= (inputs(52)) and not (inputs(178));
    layer0_outputs(3166) <= not((inputs(225)) or (inputs(140)));
    layer0_outputs(3167) <= not(inputs(72));
    layer0_outputs(3168) <= (inputs(1)) and not (inputs(240));
    layer0_outputs(3169) <= (inputs(232)) and (inputs(21));
    layer0_outputs(3170) <= not(inputs(2)) or (inputs(192));
    layer0_outputs(3171) <= not(inputs(7));
    layer0_outputs(3172) <= (inputs(17)) or (inputs(208));
    layer0_outputs(3173) <= not((inputs(9)) xor (inputs(7)));
    layer0_outputs(3174) <= (inputs(38)) and not (inputs(209));
    layer0_outputs(3175) <= (inputs(49)) or (inputs(40));
    layer0_outputs(3176) <= (inputs(75)) and not (inputs(189));
    layer0_outputs(3177) <= not((inputs(1)) or (inputs(15)));
    layer0_outputs(3178) <= not(inputs(121));
    layer0_outputs(3179) <= not(inputs(82)) or (inputs(161));
    layer0_outputs(3180) <= not((inputs(169)) or (inputs(223)));
    layer0_outputs(3181) <= inputs(148);
    layer0_outputs(3182) <= not(inputs(102));
    layer0_outputs(3183) <= (inputs(249)) xor (inputs(243));
    layer0_outputs(3184) <= not(inputs(105));
    layer0_outputs(3185) <= inputs(114);
    layer0_outputs(3186) <= (inputs(170)) or (inputs(213));
    layer0_outputs(3187) <= (inputs(186)) and not (inputs(46));
    layer0_outputs(3188) <= inputs(247);
    layer0_outputs(3189) <= not(inputs(229));
    layer0_outputs(3190) <= not(inputs(209)) or (inputs(129));
    layer0_outputs(3191) <= not(inputs(170));
    layer0_outputs(3192) <= inputs(187);
    layer0_outputs(3193) <= inputs(175);
    layer0_outputs(3194) <= inputs(94);
    layer0_outputs(3195) <= inputs(98);
    layer0_outputs(3196) <= not((inputs(241)) xor (inputs(68)));
    layer0_outputs(3197) <= inputs(85);
    layer0_outputs(3198) <= (inputs(146)) and not (inputs(32));
    layer0_outputs(3199) <= (inputs(160)) or (inputs(180));
    layer0_outputs(3200) <= inputs(246);
    layer0_outputs(3201) <= (inputs(89)) and not (inputs(85));
    layer0_outputs(3202) <= (inputs(120)) and not (inputs(145));
    layer0_outputs(3203) <= not((inputs(29)) xor (inputs(190)));
    layer0_outputs(3204) <= not(inputs(21)) or (inputs(176));
    layer0_outputs(3205) <= (inputs(217)) and not (inputs(54));
    layer0_outputs(3206) <= inputs(98);
    layer0_outputs(3207) <= not(inputs(152));
    layer0_outputs(3208) <= (inputs(132)) or (inputs(175));
    layer0_outputs(3209) <= not(inputs(33)) or (inputs(193));
    layer0_outputs(3210) <= (inputs(47)) and not (inputs(13));
    layer0_outputs(3211) <= not(inputs(238));
    layer0_outputs(3212) <= not((inputs(194)) or (inputs(101)));
    layer0_outputs(3213) <= inputs(21);
    layer0_outputs(3214) <= inputs(228);
    layer0_outputs(3215) <= not(inputs(109));
    layer0_outputs(3216) <= (inputs(48)) xor (inputs(22));
    layer0_outputs(3217) <= not(inputs(228));
    layer0_outputs(3218) <= not(inputs(38)) or (inputs(8));
    layer0_outputs(3219) <= not((inputs(102)) xor (inputs(235)));
    layer0_outputs(3220) <= not(inputs(26));
    layer0_outputs(3221) <= (inputs(123)) or (inputs(243));
    layer0_outputs(3222) <= (inputs(88)) and not (inputs(18));
    layer0_outputs(3223) <= not((inputs(240)) or (inputs(89)));
    layer0_outputs(3224) <= (inputs(236)) or (inputs(189));
    layer0_outputs(3225) <= inputs(67);
    layer0_outputs(3226) <= not(inputs(26)) or (inputs(24));
    layer0_outputs(3227) <= inputs(67);
    layer0_outputs(3228) <= inputs(232);
    layer0_outputs(3229) <= (inputs(118)) and not (inputs(241));
    layer0_outputs(3230) <= not(inputs(123)) or (inputs(138));
    layer0_outputs(3231) <= (inputs(162)) and not (inputs(252));
    layer0_outputs(3232) <= not(inputs(194));
    layer0_outputs(3233) <= (inputs(87)) xor (inputs(208));
    layer0_outputs(3234) <= not(inputs(30)) or (inputs(65));
    layer0_outputs(3235) <= not((inputs(132)) or (inputs(89)));
    layer0_outputs(3236) <= (inputs(132)) and not (inputs(223));
    layer0_outputs(3237) <= (inputs(183)) or (inputs(166));
    layer0_outputs(3238) <= (inputs(73)) and not (inputs(252));
    layer0_outputs(3239) <= (inputs(123)) or (inputs(77));
    layer0_outputs(3240) <= (inputs(209)) and not (inputs(251));
    layer0_outputs(3241) <= not(inputs(119)) or (inputs(201));
    layer0_outputs(3242) <= not(inputs(83));
    layer0_outputs(3243) <= inputs(202);
    layer0_outputs(3244) <= (inputs(197)) and not (inputs(240));
    layer0_outputs(3245) <= not(inputs(250));
    layer0_outputs(3246) <= not(inputs(85));
    layer0_outputs(3247) <= not(inputs(106));
    layer0_outputs(3248) <= not((inputs(83)) xor (inputs(111)));
    layer0_outputs(3249) <= not(inputs(195));
    layer0_outputs(3250) <= not(inputs(106)) or (inputs(71));
    layer0_outputs(3251) <= (inputs(167)) and (inputs(89));
    layer0_outputs(3252) <= not((inputs(234)) and (inputs(169)));
    layer0_outputs(3253) <= (inputs(43)) or (inputs(52));
    layer0_outputs(3254) <= not(inputs(99)) or (inputs(229));
    layer0_outputs(3255) <= inputs(133);
    layer0_outputs(3256) <= not((inputs(252)) or (inputs(49)));
    layer0_outputs(3257) <= inputs(103);
    layer0_outputs(3258) <= (inputs(103)) xor (inputs(134));
    layer0_outputs(3259) <= (inputs(174)) or (inputs(56));
    layer0_outputs(3260) <= (inputs(18)) or (inputs(12));
    layer0_outputs(3261) <= not(inputs(94));
    layer0_outputs(3262) <= not(inputs(52)) or (inputs(223));
    layer0_outputs(3263) <= not(inputs(4)) or (inputs(142));
    layer0_outputs(3264) <= not(inputs(182)) or (inputs(58));
    layer0_outputs(3265) <= not(inputs(9)) or (inputs(31));
    layer0_outputs(3266) <= not(inputs(168)) or (inputs(254));
    layer0_outputs(3267) <= inputs(174);
    layer0_outputs(3268) <= (inputs(53)) and not (inputs(187));
    layer0_outputs(3269) <= inputs(73);
    layer0_outputs(3270) <= not((inputs(150)) or (inputs(163)));
    layer0_outputs(3271) <= '0';
    layer0_outputs(3272) <= not(inputs(229));
    layer0_outputs(3273) <= not((inputs(242)) or (inputs(160)));
    layer0_outputs(3274) <= (inputs(237)) and (inputs(109));
    layer0_outputs(3275) <= not(inputs(118));
    layer0_outputs(3276) <= not(inputs(77));
    layer0_outputs(3277) <= (inputs(248)) or (inputs(142));
    layer0_outputs(3278) <= inputs(94);
    layer0_outputs(3279) <= inputs(180);
    layer0_outputs(3280) <= '1';
    layer0_outputs(3281) <= not((inputs(69)) or (inputs(30)));
    layer0_outputs(3282) <= inputs(203);
    layer0_outputs(3283) <= not(inputs(116));
    layer0_outputs(3284) <= not((inputs(74)) xor (inputs(26)));
    layer0_outputs(3285) <= not((inputs(89)) and (inputs(90)));
    layer0_outputs(3286) <= not((inputs(255)) xor (inputs(135)));
    layer0_outputs(3287) <= not((inputs(159)) xor (inputs(8)));
    layer0_outputs(3288) <= inputs(48);
    layer0_outputs(3289) <= (inputs(11)) or (inputs(140));
    layer0_outputs(3290) <= (inputs(229)) and (inputs(233));
    layer0_outputs(3291) <= not(inputs(115)) or (inputs(11));
    layer0_outputs(3292) <= not(inputs(18)) or (inputs(13));
    layer0_outputs(3293) <= not((inputs(82)) xor (inputs(243)));
    layer0_outputs(3294) <= inputs(226);
    layer0_outputs(3295) <= not((inputs(162)) or (inputs(213)));
    layer0_outputs(3296) <= not((inputs(92)) xor (inputs(89)));
    layer0_outputs(3297) <= not(inputs(137));
    layer0_outputs(3298) <= (inputs(205)) and not (inputs(81));
    layer0_outputs(3299) <= not((inputs(101)) or (inputs(117)));
    layer0_outputs(3300) <= (inputs(67)) and not (inputs(125));
    layer0_outputs(3301) <= (inputs(4)) and not (inputs(47));
    layer0_outputs(3302) <= not(inputs(237));
    layer0_outputs(3303) <= not(inputs(182));
    layer0_outputs(3304) <= not(inputs(202));
    layer0_outputs(3305) <= inputs(90);
    layer0_outputs(3306) <= (inputs(127)) and not (inputs(32));
    layer0_outputs(3307) <= inputs(56);
    layer0_outputs(3308) <= '1';
    layer0_outputs(3309) <= not((inputs(64)) xor (inputs(20)));
    layer0_outputs(3310) <= '0';
    layer0_outputs(3311) <= (inputs(221)) and (inputs(226));
    layer0_outputs(3312) <= '1';
    layer0_outputs(3313) <= (inputs(9)) xor (inputs(40));
    layer0_outputs(3314) <= (inputs(214)) and not (inputs(237));
    layer0_outputs(3315) <= (inputs(246)) and not (inputs(51));
    layer0_outputs(3316) <= '1';
    layer0_outputs(3317) <= not((inputs(219)) xor (inputs(146)));
    layer0_outputs(3318) <= (inputs(176)) and not (inputs(0));
    layer0_outputs(3319) <= inputs(5);
    layer0_outputs(3320) <= inputs(65);
    layer0_outputs(3321) <= (inputs(175)) or (inputs(219));
    layer0_outputs(3322) <= (inputs(246)) and not (inputs(51));
    layer0_outputs(3323) <= (inputs(164)) or (inputs(232));
    layer0_outputs(3324) <= not(inputs(125));
    layer0_outputs(3325) <= inputs(169);
    layer0_outputs(3326) <= (inputs(242)) or (inputs(22));
    layer0_outputs(3327) <= (inputs(40)) and not (inputs(119));
    layer0_outputs(3328) <= not(inputs(222));
    layer0_outputs(3329) <= not((inputs(37)) or (inputs(214)));
    layer0_outputs(3330) <= '0';
    layer0_outputs(3331) <= not((inputs(74)) or (inputs(142)));
    layer0_outputs(3332) <= not(inputs(88)) or (inputs(53));
    layer0_outputs(3333) <= not(inputs(90)) or (inputs(214));
    layer0_outputs(3334) <= (inputs(139)) and not (inputs(231));
    layer0_outputs(3335) <= not(inputs(216)) or (inputs(169));
    layer0_outputs(3336) <= not(inputs(211)) or (inputs(167));
    layer0_outputs(3337) <= not((inputs(34)) or (inputs(15)));
    layer0_outputs(3338) <= not(inputs(134));
    layer0_outputs(3339) <= not(inputs(10)) or (inputs(162));
    layer0_outputs(3340) <= (inputs(191)) or (inputs(125));
    layer0_outputs(3341) <= not(inputs(80));
    layer0_outputs(3342) <= not(inputs(93));
    layer0_outputs(3343) <= not(inputs(120));
    layer0_outputs(3344) <= not(inputs(98));
    layer0_outputs(3345) <= (inputs(173)) or (inputs(180));
    layer0_outputs(3346) <= not((inputs(188)) or (inputs(190)));
    layer0_outputs(3347) <= (inputs(185)) and not (inputs(108));
    layer0_outputs(3348) <= not(inputs(109)) or (inputs(149));
    layer0_outputs(3349) <= not(inputs(147));
    layer0_outputs(3350) <= (inputs(252)) and (inputs(63));
    layer0_outputs(3351) <= (inputs(44)) and not (inputs(197));
    layer0_outputs(3352) <= (inputs(85)) and not (inputs(241));
    layer0_outputs(3353) <= (inputs(155)) or (inputs(128));
    layer0_outputs(3354) <= inputs(158);
    layer0_outputs(3355) <= inputs(60);
    layer0_outputs(3356) <= (inputs(13)) and not (inputs(208));
    layer0_outputs(3357) <= not((inputs(96)) and (inputs(84)));
    layer0_outputs(3358) <= (inputs(22)) or (inputs(225));
    layer0_outputs(3359) <= not((inputs(110)) or (inputs(191)));
    layer0_outputs(3360) <= inputs(75);
    layer0_outputs(3361) <= '0';
    layer0_outputs(3362) <= inputs(107);
    layer0_outputs(3363) <= inputs(26);
    layer0_outputs(3364) <= not((inputs(177)) or (inputs(164)));
    layer0_outputs(3365) <= not((inputs(207)) or (inputs(77)));
    layer0_outputs(3366) <= (inputs(182)) or (inputs(14));
    layer0_outputs(3367) <= (inputs(103)) xor (inputs(10));
    layer0_outputs(3368) <= not(inputs(108));
    layer0_outputs(3369) <= (inputs(143)) xor (inputs(134));
    layer0_outputs(3370) <= not(inputs(21)) or (inputs(240));
    layer0_outputs(3371) <= not((inputs(39)) or (inputs(99)));
    layer0_outputs(3372) <= inputs(113);
    layer0_outputs(3373) <= (inputs(245)) and not (inputs(31));
    layer0_outputs(3374) <= (inputs(195)) or (inputs(173));
    layer0_outputs(3375) <= (inputs(158)) xor (inputs(171));
    layer0_outputs(3376) <= inputs(186);
    layer0_outputs(3377) <= not(inputs(176));
    layer0_outputs(3378) <= '1';
    layer0_outputs(3379) <= (inputs(153)) or (inputs(224));
    layer0_outputs(3380) <= not((inputs(224)) xor (inputs(2)));
    layer0_outputs(3381) <= not((inputs(65)) or (inputs(39)));
    layer0_outputs(3382) <= inputs(151);
    layer0_outputs(3383) <= not((inputs(132)) or (inputs(231)));
    layer0_outputs(3384) <= not(inputs(201)) or (inputs(45));
    layer0_outputs(3385) <= (inputs(104)) or (inputs(80));
    layer0_outputs(3386) <= (inputs(24)) and not (inputs(225));
    layer0_outputs(3387) <= inputs(211);
    layer0_outputs(3388) <= not(inputs(178)) or (inputs(222));
    layer0_outputs(3389) <= not((inputs(214)) or (inputs(33)));
    layer0_outputs(3390) <= (inputs(235)) or (inputs(180));
    layer0_outputs(3391) <= not(inputs(26));
    layer0_outputs(3392) <= (inputs(9)) and not (inputs(141));
    layer0_outputs(3393) <= not(inputs(231)) or (inputs(62));
    layer0_outputs(3394) <= inputs(77);
    layer0_outputs(3395) <= not(inputs(154)) or (inputs(111));
    layer0_outputs(3396) <= not(inputs(136)) or (inputs(73));
    layer0_outputs(3397) <= (inputs(72)) and not (inputs(137));
    layer0_outputs(3398) <= inputs(148);
    layer0_outputs(3399) <= '0';
    layer0_outputs(3400) <= not(inputs(212)) or (inputs(115));
    layer0_outputs(3401) <= inputs(35);
    layer0_outputs(3402) <= not(inputs(220)) or (inputs(16));
    layer0_outputs(3403) <= (inputs(71)) and not (inputs(142));
    layer0_outputs(3404) <= not((inputs(206)) xor (inputs(85)));
    layer0_outputs(3405) <= not((inputs(63)) or (inputs(226)));
    layer0_outputs(3406) <= (inputs(119)) and not (inputs(30));
    layer0_outputs(3407) <= not(inputs(42)) or (inputs(129));
    layer0_outputs(3408) <= not(inputs(83));
    layer0_outputs(3409) <= not(inputs(70)) or (inputs(157));
    layer0_outputs(3410) <= not(inputs(162));
    layer0_outputs(3411) <= (inputs(23)) and (inputs(75));
    layer0_outputs(3412) <= not(inputs(129));
    layer0_outputs(3413) <= not(inputs(56));
    layer0_outputs(3414) <= not(inputs(13));
    layer0_outputs(3415) <= not(inputs(41));
    layer0_outputs(3416) <= inputs(156);
    layer0_outputs(3417) <= not(inputs(138));
    layer0_outputs(3418) <= not(inputs(115));
    layer0_outputs(3419) <= inputs(228);
    layer0_outputs(3420) <= inputs(245);
    layer0_outputs(3421) <= not((inputs(236)) or (inputs(181)));
    layer0_outputs(3422) <= (inputs(2)) or (inputs(188));
    layer0_outputs(3423) <= not(inputs(31));
    layer0_outputs(3424) <= not(inputs(158));
    layer0_outputs(3425) <= inputs(161);
    layer0_outputs(3426) <= not(inputs(42));
    layer0_outputs(3427) <= '1';
    layer0_outputs(3428) <= inputs(131);
    layer0_outputs(3429) <= inputs(44);
    layer0_outputs(3430) <= (inputs(231)) and (inputs(26));
    layer0_outputs(3431) <= inputs(23);
    layer0_outputs(3432) <= not(inputs(252));
    layer0_outputs(3433) <= inputs(134);
    layer0_outputs(3434) <= (inputs(173)) or (inputs(97));
    layer0_outputs(3435) <= not(inputs(7));
    layer0_outputs(3436) <= inputs(104);
    layer0_outputs(3437) <= not((inputs(207)) or (inputs(230)));
    layer0_outputs(3438) <= (inputs(35)) or (inputs(49));
    layer0_outputs(3439) <= (inputs(96)) and not (inputs(52));
    layer0_outputs(3440) <= (inputs(22)) xor (inputs(93));
    layer0_outputs(3441) <= inputs(84);
    layer0_outputs(3442) <= inputs(22);
    layer0_outputs(3443) <= not(inputs(211)) or (inputs(218));
    layer0_outputs(3444) <= not(inputs(145));
    layer0_outputs(3445) <= not(inputs(82));
    layer0_outputs(3446) <= (inputs(212)) and not (inputs(241));
    layer0_outputs(3447) <= inputs(209);
    layer0_outputs(3448) <= not((inputs(12)) xor (inputs(194)));
    layer0_outputs(3449) <= not(inputs(197));
    layer0_outputs(3450) <= (inputs(203)) and not (inputs(108));
    layer0_outputs(3451) <= not(inputs(120));
    layer0_outputs(3452) <= (inputs(71)) and not (inputs(67));
    layer0_outputs(3453) <= inputs(76);
    layer0_outputs(3454) <= not((inputs(91)) or (inputs(108)));
    layer0_outputs(3455) <= (inputs(7)) and not (inputs(184));
    layer0_outputs(3456) <= not(inputs(61)) or (inputs(249));
    layer0_outputs(3457) <= not(inputs(222));
    layer0_outputs(3458) <= (inputs(71)) and not (inputs(110));
    layer0_outputs(3459) <= not((inputs(194)) xor (inputs(181)));
    layer0_outputs(3460) <= (inputs(174)) or (inputs(173));
    layer0_outputs(3461) <= inputs(144);
    layer0_outputs(3462) <= inputs(224);
    layer0_outputs(3463) <= inputs(24);
    layer0_outputs(3464) <= '1';
    layer0_outputs(3465) <= not((inputs(250)) or (inputs(249)));
    layer0_outputs(3466) <= inputs(167);
    layer0_outputs(3467) <= inputs(193);
    layer0_outputs(3468) <= not(inputs(208));
    layer0_outputs(3469) <= not(inputs(43)) or (inputs(25));
    layer0_outputs(3470) <= not((inputs(100)) or (inputs(131)));
    layer0_outputs(3471) <= not((inputs(80)) or (inputs(150)));
    layer0_outputs(3472) <= not(inputs(18));
    layer0_outputs(3473) <= inputs(88);
    layer0_outputs(3474) <= not(inputs(194)) or (inputs(68));
    layer0_outputs(3475) <= not((inputs(94)) or (inputs(240)));
    layer0_outputs(3476) <= (inputs(132)) or (inputs(198));
    layer0_outputs(3477) <= (inputs(92)) and not (inputs(46));
    layer0_outputs(3478) <= inputs(63);
    layer0_outputs(3479) <= inputs(223);
    layer0_outputs(3480) <= (inputs(218)) and not (inputs(77));
    layer0_outputs(3481) <= not(inputs(132));
    layer0_outputs(3482) <= inputs(103);
    layer0_outputs(3483) <= (inputs(132)) xor (inputs(146));
    layer0_outputs(3484) <= (inputs(118)) and not (inputs(65));
    layer0_outputs(3485) <= '1';
    layer0_outputs(3486) <= not(inputs(129));
    layer0_outputs(3487) <= (inputs(197)) or (inputs(115));
    layer0_outputs(3488) <= inputs(18);
    layer0_outputs(3489) <= inputs(90);
    layer0_outputs(3490) <= (inputs(16)) xor (inputs(63));
    layer0_outputs(3491) <= not(inputs(170)) or (inputs(29));
    layer0_outputs(3492) <= not(inputs(121)) or (inputs(70));
    layer0_outputs(3493) <= not((inputs(60)) or (inputs(15)));
    layer0_outputs(3494) <= '0';
    layer0_outputs(3495) <= not(inputs(32));
    layer0_outputs(3496) <= not((inputs(64)) xor (inputs(188)));
    layer0_outputs(3497) <= not(inputs(195));
    layer0_outputs(3498) <= inputs(78);
    layer0_outputs(3499) <= inputs(247);
    layer0_outputs(3500) <= not(inputs(22));
    layer0_outputs(3501) <= inputs(166);
    layer0_outputs(3502) <= (inputs(161)) and (inputs(254));
    layer0_outputs(3503) <= not((inputs(23)) or (inputs(187)));
    layer0_outputs(3504) <= (inputs(68)) and not (inputs(219));
    layer0_outputs(3505) <= not((inputs(160)) or (inputs(179)));
    layer0_outputs(3506) <= '1';
    layer0_outputs(3507) <= (inputs(167)) and not (inputs(187));
    layer0_outputs(3508) <= inputs(236);
    layer0_outputs(3509) <= not((inputs(75)) and (inputs(71)));
    layer0_outputs(3510) <= inputs(130);
    layer0_outputs(3511) <= not(inputs(59)) or (inputs(182));
    layer0_outputs(3512) <= not(inputs(73)) or (inputs(166));
    layer0_outputs(3513) <= not(inputs(214)) or (inputs(114));
    layer0_outputs(3514) <= inputs(187);
    layer0_outputs(3515) <= (inputs(74)) or (inputs(16));
    layer0_outputs(3516) <= inputs(176);
    layer0_outputs(3517) <= not(inputs(86));
    layer0_outputs(3518) <= (inputs(89)) and not (inputs(192));
    layer0_outputs(3519) <= inputs(116);
    layer0_outputs(3520) <= (inputs(37)) and not (inputs(204));
    layer0_outputs(3521) <= inputs(197);
    layer0_outputs(3522) <= inputs(230);
    layer0_outputs(3523) <= inputs(37);
    layer0_outputs(3524) <= inputs(216);
    layer0_outputs(3525) <= not((inputs(3)) or (inputs(171)));
    layer0_outputs(3526) <= (inputs(173)) and not (inputs(16));
    layer0_outputs(3527) <= not((inputs(118)) or (inputs(155)));
    layer0_outputs(3528) <= inputs(77);
    layer0_outputs(3529) <= not(inputs(170)) or (inputs(183));
    layer0_outputs(3530) <= (inputs(77)) and not (inputs(89));
    layer0_outputs(3531) <= '0';
    layer0_outputs(3532) <= (inputs(196)) and not (inputs(19));
    layer0_outputs(3533) <= (inputs(39)) and not (inputs(92));
    layer0_outputs(3534) <= (inputs(13)) and not (inputs(35));
    layer0_outputs(3535) <= inputs(192);
    layer0_outputs(3536) <= not(inputs(187));
    layer0_outputs(3537) <= inputs(154);
    layer0_outputs(3538) <= not(inputs(230));
    layer0_outputs(3539) <= inputs(246);
    layer0_outputs(3540) <= (inputs(21)) or (inputs(34));
    layer0_outputs(3541) <= not(inputs(204)) or (inputs(34));
    layer0_outputs(3542) <= (inputs(15)) and not (inputs(185));
    layer0_outputs(3543) <= not((inputs(112)) or (inputs(248)));
    layer0_outputs(3544) <= not((inputs(125)) xor (inputs(64)));
    layer0_outputs(3545) <= inputs(1);
    layer0_outputs(3546) <= '1';
    layer0_outputs(3547) <= (inputs(192)) and (inputs(212));
    layer0_outputs(3548) <= not((inputs(175)) or (inputs(218)));
    layer0_outputs(3549) <= not(inputs(129));
    layer0_outputs(3550) <= not(inputs(189)) or (inputs(208));
    layer0_outputs(3551) <= inputs(97);
    layer0_outputs(3552) <= not(inputs(149)) or (inputs(19));
    layer0_outputs(3553) <= (inputs(1)) and not (inputs(127));
    layer0_outputs(3554) <= not(inputs(141));
    layer0_outputs(3555) <= not((inputs(190)) or (inputs(206)));
    layer0_outputs(3556) <= not((inputs(221)) or (inputs(177)));
    layer0_outputs(3557) <= (inputs(153)) and not (inputs(102));
    layer0_outputs(3558) <= not(inputs(91)) or (inputs(219));
    layer0_outputs(3559) <= (inputs(205)) and not (inputs(14));
    layer0_outputs(3560) <= (inputs(10)) and not (inputs(70));
    layer0_outputs(3561) <= not((inputs(253)) or (inputs(212)));
    layer0_outputs(3562) <= inputs(121);
    layer0_outputs(3563) <= not((inputs(127)) or (inputs(177)));
    layer0_outputs(3564) <= not((inputs(152)) and (inputs(121)));
    layer0_outputs(3565) <= not(inputs(56)) or (inputs(26));
    layer0_outputs(3566) <= (inputs(244)) and not (inputs(106));
    layer0_outputs(3567) <= inputs(230);
    layer0_outputs(3568) <= (inputs(251)) and not (inputs(55));
    layer0_outputs(3569) <= not(inputs(4));
    layer0_outputs(3570) <= not((inputs(239)) or (inputs(110)));
    layer0_outputs(3571) <= not((inputs(225)) or (inputs(31)));
    layer0_outputs(3572) <= (inputs(246)) xor (inputs(208));
    layer0_outputs(3573) <= inputs(212);
    layer0_outputs(3574) <= (inputs(253)) or (inputs(24));
    layer0_outputs(3575) <= not(inputs(252));
    layer0_outputs(3576) <= inputs(235);
    layer0_outputs(3577) <= not((inputs(239)) or (inputs(23)));
    layer0_outputs(3578) <= (inputs(197)) and not (inputs(142));
    layer0_outputs(3579) <= not(inputs(42)) or (inputs(18));
    layer0_outputs(3580) <= inputs(62);
    layer0_outputs(3581) <= not(inputs(240)) or (inputs(85));
    layer0_outputs(3582) <= inputs(40);
    layer0_outputs(3583) <= (inputs(252)) or (inputs(239));
    layer0_outputs(3584) <= inputs(198);
    layer0_outputs(3585) <= (inputs(18)) or (inputs(223));
    layer0_outputs(3586) <= not(inputs(151));
    layer0_outputs(3587) <= not((inputs(174)) xor (inputs(221)));
    layer0_outputs(3588) <= (inputs(243)) xor (inputs(48));
    layer0_outputs(3589) <= not((inputs(25)) or (inputs(48)));
    layer0_outputs(3590) <= (inputs(231)) and not (inputs(112));
    layer0_outputs(3591) <= not(inputs(46));
    layer0_outputs(3592) <= not((inputs(186)) xor (inputs(193)));
    layer0_outputs(3593) <= not(inputs(26));
    layer0_outputs(3594) <= (inputs(178)) or (inputs(213));
    layer0_outputs(3595) <= '1';
    layer0_outputs(3596) <= not(inputs(132)) or (inputs(16));
    layer0_outputs(3597) <= not((inputs(206)) or (inputs(77)));
    layer0_outputs(3598) <= (inputs(238)) xor (inputs(249));
    layer0_outputs(3599) <= not((inputs(27)) or (inputs(56)));
    layer0_outputs(3600) <= inputs(140);
    layer0_outputs(3601) <= not(inputs(20)) or (inputs(114));
    layer0_outputs(3602) <= (inputs(10)) or (inputs(178));
    layer0_outputs(3603) <= not((inputs(62)) xor (inputs(255)));
    layer0_outputs(3604) <= inputs(98);
    layer0_outputs(3605) <= (inputs(100)) and not (inputs(235));
    layer0_outputs(3606) <= (inputs(250)) or (inputs(169));
    layer0_outputs(3607) <= '0';
    layer0_outputs(3608) <= not(inputs(16));
    layer0_outputs(3609) <= not((inputs(89)) xor (inputs(182)));
    layer0_outputs(3610) <= not(inputs(78));
    layer0_outputs(3611) <= (inputs(215)) and not (inputs(86));
    layer0_outputs(3612) <= not(inputs(140)) or (inputs(254));
    layer0_outputs(3613) <= (inputs(72)) and not (inputs(44));
    layer0_outputs(3614) <= (inputs(109)) and not (inputs(209));
    layer0_outputs(3615) <= not(inputs(74));
    layer0_outputs(3616) <= not(inputs(124)) or (inputs(80));
    layer0_outputs(3617) <= '0';
    layer0_outputs(3618) <= inputs(41);
    layer0_outputs(3619) <= '0';
    layer0_outputs(3620) <= not(inputs(187)) or (inputs(223));
    layer0_outputs(3621) <= (inputs(40)) and not (inputs(236));
    layer0_outputs(3622) <= inputs(70);
    layer0_outputs(3623) <= (inputs(67)) and not (inputs(1));
    layer0_outputs(3624) <= inputs(102);
    layer0_outputs(3625) <= inputs(22);
    layer0_outputs(3626) <= not(inputs(144));
    layer0_outputs(3627) <= not(inputs(232));
    layer0_outputs(3628) <= not((inputs(49)) or (inputs(67)));
    layer0_outputs(3629) <= (inputs(27)) and not (inputs(189));
    layer0_outputs(3630) <= not(inputs(83));
    layer0_outputs(3631) <= (inputs(158)) or (inputs(202));
    layer0_outputs(3632) <= not(inputs(189)) or (inputs(147));
    layer0_outputs(3633) <= not((inputs(101)) or (inputs(147)));
    layer0_outputs(3634) <= inputs(173);
    layer0_outputs(3635) <= inputs(147);
    layer0_outputs(3636) <= (inputs(212)) xor (inputs(90));
    layer0_outputs(3637) <= not((inputs(105)) and (inputs(82)));
    layer0_outputs(3638) <= inputs(49);
    layer0_outputs(3639) <= not((inputs(106)) xor (inputs(172)));
    layer0_outputs(3640) <= (inputs(0)) or (inputs(20));
    layer0_outputs(3641) <= not((inputs(238)) xor (inputs(139)));
    layer0_outputs(3642) <= inputs(209);
    layer0_outputs(3643) <= (inputs(241)) xor (inputs(17));
    layer0_outputs(3644) <= not(inputs(178));
    layer0_outputs(3645) <= not(inputs(175)) or (inputs(154));
    layer0_outputs(3646) <= not((inputs(130)) or (inputs(113)));
    layer0_outputs(3647) <= inputs(180);
    layer0_outputs(3648) <= not(inputs(242));
    layer0_outputs(3649) <= inputs(219);
    layer0_outputs(3650) <= (inputs(0)) and not (inputs(119));
    layer0_outputs(3651) <= not(inputs(157));
    layer0_outputs(3652) <= (inputs(46)) or (inputs(128));
    layer0_outputs(3653) <= not((inputs(87)) and (inputs(31)));
    layer0_outputs(3654) <= (inputs(202)) and not (inputs(232));
    layer0_outputs(3655) <= not(inputs(206));
    layer0_outputs(3656) <= inputs(155);
    layer0_outputs(3657) <= not((inputs(110)) or (inputs(3)));
    layer0_outputs(3658) <= not(inputs(253)) or (inputs(104));
    layer0_outputs(3659) <= (inputs(154)) or (inputs(118));
    layer0_outputs(3660) <= not((inputs(2)) xor (inputs(255)));
    layer0_outputs(3661) <= not(inputs(142));
    layer0_outputs(3662) <= not((inputs(131)) and (inputs(44)));
    layer0_outputs(3663) <= not(inputs(167));
    layer0_outputs(3664) <= inputs(97);
    layer0_outputs(3665) <= not(inputs(217));
    layer0_outputs(3666) <= not(inputs(205)) or (inputs(14));
    layer0_outputs(3667) <= not((inputs(57)) xor (inputs(13)));
    layer0_outputs(3668) <= inputs(140);
    layer0_outputs(3669) <= not(inputs(177)) or (inputs(74));
    layer0_outputs(3670) <= not(inputs(249));
    layer0_outputs(3671) <= (inputs(183)) or (inputs(174));
    layer0_outputs(3672) <= not(inputs(190));
    layer0_outputs(3673) <= (inputs(253)) and not (inputs(14));
    layer0_outputs(3674) <= (inputs(251)) and (inputs(205));
    layer0_outputs(3675) <= not((inputs(175)) or (inputs(216)));
    layer0_outputs(3676) <= inputs(78);
    layer0_outputs(3677) <= (inputs(28)) and not (inputs(56));
    layer0_outputs(3678) <= not(inputs(115));
    layer0_outputs(3679) <= (inputs(187)) and not (inputs(239));
    layer0_outputs(3680) <= not((inputs(92)) or (inputs(80)));
    layer0_outputs(3681) <= not(inputs(133));
    layer0_outputs(3682) <= not((inputs(23)) or (inputs(190)));
    layer0_outputs(3683) <= (inputs(208)) or (inputs(188));
    layer0_outputs(3684) <= not(inputs(103));
    layer0_outputs(3685) <= not(inputs(47));
    layer0_outputs(3686) <= not((inputs(194)) or (inputs(186)));
    layer0_outputs(3687) <= not(inputs(71));
    layer0_outputs(3688) <= not((inputs(64)) or (inputs(7)));
    layer0_outputs(3689) <= not((inputs(210)) xor (inputs(240)));
    layer0_outputs(3690) <= not(inputs(91));
    layer0_outputs(3691) <= not(inputs(19)) or (inputs(113));
    layer0_outputs(3692) <= (inputs(170)) or (inputs(253));
    layer0_outputs(3693) <= inputs(104);
    layer0_outputs(3694) <= inputs(140);
    layer0_outputs(3695) <= not(inputs(55));
    layer0_outputs(3696) <= inputs(166);
    layer0_outputs(3697) <= not(inputs(28)) or (inputs(235));
    layer0_outputs(3698) <= inputs(23);
    layer0_outputs(3699) <= inputs(108);
    layer0_outputs(3700) <= inputs(135);
    layer0_outputs(3701) <= inputs(181);
    layer0_outputs(3702) <= (inputs(29)) and not (inputs(175));
    layer0_outputs(3703) <= not(inputs(137)) or (inputs(130));
    layer0_outputs(3704) <= not(inputs(84));
    layer0_outputs(3705) <= (inputs(202)) or (inputs(255));
    layer0_outputs(3706) <= (inputs(16)) or (inputs(130));
    layer0_outputs(3707) <= not((inputs(232)) or (inputs(4)));
    layer0_outputs(3708) <= (inputs(164)) xor (inputs(145));
    layer0_outputs(3709) <= inputs(104);
    layer0_outputs(3710) <= not((inputs(39)) or (inputs(95)));
    layer0_outputs(3711) <= (inputs(40)) and (inputs(114));
    layer0_outputs(3712) <= inputs(158);
    layer0_outputs(3713) <= not((inputs(126)) and (inputs(240)));
    layer0_outputs(3714) <= (inputs(142)) or (inputs(21));
    layer0_outputs(3715) <= not(inputs(184)) or (inputs(144));
    layer0_outputs(3716) <= inputs(107);
    layer0_outputs(3717) <= (inputs(108)) or (inputs(58));
    layer0_outputs(3718) <= inputs(127);
    layer0_outputs(3719) <= (inputs(87)) or (inputs(209));
    layer0_outputs(3720) <= (inputs(7)) and not (inputs(114));
    layer0_outputs(3721) <= inputs(110);
    layer0_outputs(3722) <= (inputs(79)) or (inputs(39));
    layer0_outputs(3723) <= not(inputs(28)) or (inputs(35));
    layer0_outputs(3724) <= not((inputs(240)) or (inputs(206)));
    layer0_outputs(3725) <= inputs(179);
    layer0_outputs(3726) <= (inputs(106)) and not (inputs(253));
    layer0_outputs(3727) <= (inputs(5)) or (inputs(90));
    layer0_outputs(3728) <= (inputs(47)) or (inputs(93));
    layer0_outputs(3729) <= (inputs(211)) or (inputs(228));
    layer0_outputs(3730) <= not(inputs(153));
    layer0_outputs(3731) <= inputs(105);
    layer0_outputs(3732) <= not(inputs(248));
    layer0_outputs(3733) <= not((inputs(102)) or (inputs(21)));
    layer0_outputs(3734) <= (inputs(180)) or (inputs(227));
    layer0_outputs(3735) <= inputs(48);
    layer0_outputs(3736) <= (inputs(97)) and not (inputs(97));
    layer0_outputs(3737) <= not(inputs(186));
    layer0_outputs(3738) <= (inputs(56)) and not (inputs(250));
    layer0_outputs(3739) <= inputs(181);
    layer0_outputs(3740) <= (inputs(81)) and not (inputs(240));
    layer0_outputs(3741) <= inputs(57);
    layer0_outputs(3742) <= not(inputs(53));
    layer0_outputs(3743) <= not(inputs(27)) or (inputs(157));
    layer0_outputs(3744) <= (inputs(126)) or (inputs(151));
    layer0_outputs(3745) <= not(inputs(43));
    layer0_outputs(3746) <= inputs(106);
    layer0_outputs(3747) <= (inputs(169)) or (inputs(161));
    layer0_outputs(3748) <= (inputs(213)) or (inputs(32));
    layer0_outputs(3749) <= not(inputs(60)) or (inputs(100));
    layer0_outputs(3750) <= (inputs(90)) xor (inputs(138));
    layer0_outputs(3751) <= (inputs(215)) or (inputs(211));
    layer0_outputs(3752) <= inputs(24);
    layer0_outputs(3753) <= not((inputs(112)) xor (inputs(244)));
    layer0_outputs(3754) <= '1';
    layer0_outputs(3755) <= (inputs(159)) or (inputs(78));
    layer0_outputs(3756) <= '1';
    layer0_outputs(3757) <= not((inputs(91)) xor (inputs(190)));
    layer0_outputs(3758) <= inputs(211);
    layer0_outputs(3759) <= not(inputs(135)) or (inputs(160));
    layer0_outputs(3760) <= inputs(19);
    layer0_outputs(3761) <= (inputs(158)) or (inputs(12));
    layer0_outputs(3762) <= '0';
    layer0_outputs(3763) <= not((inputs(229)) or (inputs(34)));
    layer0_outputs(3764) <= (inputs(111)) or (inputs(122));
    layer0_outputs(3765) <= (inputs(138)) and not (inputs(21));
    layer0_outputs(3766) <= not(inputs(145));
    layer0_outputs(3767) <= not(inputs(83)) or (inputs(193));
    layer0_outputs(3768) <= inputs(196);
    layer0_outputs(3769) <= not((inputs(72)) xor (inputs(128)));
    layer0_outputs(3770) <= (inputs(43)) and not (inputs(199));
    layer0_outputs(3771) <= not(inputs(215));
    layer0_outputs(3772) <= not(inputs(100));
    layer0_outputs(3773) <= (inputs(96)) or (inputs(101));
    layer0_outputs(3774) <= not((inputs(196)) xor (inputs(137)));
    layer0_outputs(3775) <= not(inputs(72)) or (inputs(95));
    layer0_outputs(3776) <= not(inputs(169));
    layer0_outputs(3777) <= not((inputs(51)) or (inputs(146)));
    layer0_outputs(3778) <= not(inputs(174));
    layer0_outputs(3779) <= not((inputs(109)) xor (inputs(81)));
    layer0_outputs(3780) <= not(inputs(31)) or (inputs(92));
    layer0_outputs(3781) <= (inputs(89)) or (inputs(243));
    layer0_outputs(3782) <= not(inputs(105));
    layer0_outputs(3783) <= '1';
    layer0_outputs(3784) <= inputs(145);
    layer0_outputs(3785) <= not((inputs(183)) or (inputs(167)));
    layer0_outputs(3786) <= not((inputs(59)) or (inputs(6)));
    layer0_outputs(3787) <= (inputs(245)) or (inputs(102));
    layer0_outputs(3788) <= not((inputs(204)) and (inputs(216)));
    layer0_outputs(3789) <= not(inputs(213));
    layer0_outputs(3790) <= not(inputs(163));
    layer0_outputs(3791) <= not((inputs(210)) or (inputs(0)));
    layer0_outputs(3792) <= (inputs(235)) or (inputs(159));
    layer0_outputs(3793) <= not(inputs(171));
    layer0_outputs(3794) <= not(inputs(195));
    layer0_outputs(3795) <= not((inputs(227)) or (inputs(71)));
    layer0_outputs(3796) <= not((inputs(2)) and (inputs(199)));
    layer0_outputs(3797) <= inputs(84);
    layer0_outputs(3798) <= not(inputs(169));
    layer0_outputs(3799) <= (inputs(43)) and not (inputs(99));
    layer0_outputs(3800) <= not((inputs(157)) or (inputs(140)));
    layer0_outputs(3801) <= not((inputs(107)) or (inputs(17)));
    layer0_outputs(3802) <= not(inputs(93));
    layer0_outputs(3803) <= not(inputs(166));
    layer0_outputs(3804) <= (inputs(118)) or (inputs(150));
    layer0_outputs(3805) <= not((inputs(70)) or (inputs(127)));
    layer0_outputs(3806) <= not(inputs(57));
    layer0_outputs(3807) <= not((inputs(17)) xor (inputs(95)));
    layer0_outputs(3808) <= (inputs(251)) or (inputs(149));
    layer0_outputs(3809) <= (inputs(225)) or (inputs(11));
    layer0_outputs(3810) <= not(inputs(214));
    layer0_outputs(3811) <= not((inputs(80)) or (inputs(84)));
    layer0_outputs(3812) <= not(inputs(247));
    layer0_outputs(3813) <= inputs(89);
    layer0_outputs(3814) <= not(inputs(35));
    layer0_outputs(3815) <= (inputs(233)) xor (inputs(111));
    layer0_outputs(3816) <= not((inputs(30)) or (inputs(151)));
    layer0_outputs(3817) <= '0';
    layer0_outputs(3818) <= inputs(77);
    layer0_outputs(3819) <= (inputs(140)) or (inputs(66));
    layer0_outputs(3820) <= inputs(67);
    layer0_outputs(3821) <= not(inputs(247));
    layer0_outputs(3822) <= (inputs(204)) or (inputs(165));
    layer0_outputs(3823) <= not((inputs(60)) xor (inputs(223)));
    layer0_outputs(3824) <= not((inputs(117)) or (inputs(143)));
    layer0_outputs(3825) <= (inputs(250)) and not (inputs(177));
    layer0_outputs(3826) <= (inputs(4)) or (inputs(149));
    layer0_outputs(3827) <= (inputs(190)) xor (inputs(49));
    layer0_outputs(3828) <= (inputs(123)) or (inputs(8));
    layer0_outputs(3829) <= not((inputs(45)) or (inputs(52)));
    layer0_outputs(3830) <= inputs(138);
    layer0_outputs(3831) <= not((inputs(160)) or (inputs(148)));
    layer0_outputs(3832) <= inputs(227);
    layer0_outputs(3833) <= '1';
    layer0_outputs(3834) <= not((inputs(196)) or (inputs(212)));
    layer0_outputs(3835) <= (inputs(96)) or (inputs(102));
    layer0_outputs(3836) <= not(inputs(93)) or (inputs(134));
    layer0_outputs(3837) <= (inputs(116)) and not (inputs(72));
    layer0_outputs(3838) <= not(inputs(135));
    layer0_outputs(3839) <= inputs(217);
    layer0_outputs(3840) <= not((inputs(59)) xor (inputs(38)));
    layer0_outputs(3841) <= not(inputs(217)) or (inputs(223));
    layer0_outputs(3842) <= (inputs(136)) xor (inputs(109));
    layer0_outputs(3843) <= not(inputs(253)) or (inputs(160));
    layer0_outputs(3844) <= not(inputs(37)) or (inputs(40));
    layer0_outputs(3845) <= not(inputs(176));
    layer0_outputs(3846) <= not((inputs(241)) or (inputs(245)));
    layer0_outputs(3847) <= not(inputs(217));
    layer0_outputs(3848) <= inputs(244);
    layer0_outputs(3849) <= (inputs(146)) and not (inputs(73));
    layer0_outputs(3850) <= not((inputs(197)) xor (inputs(96)));
    layer0_outputs(3851) <= not((inputs(188)) or (inputs(203)));
    layer0_outputs(3852) <= not(inputs(118));
    layer0_outputs(3853) <= inputs(206);
    layer0_outputs(3854) <= not(inputs(57)) or (inputs(52));
    layer0_outputs(3855) <= not(inputs(195)) or (inputs(13));
    layer0_outputs(3856) <= not(inputs(211));
    layer0_outputs(3857) <= (inputs(32)) or (inputs(247));
    layer0_outputs(3858) <= '0';
    layer0_outputs(3859) <= not((inputs(225)) xor (inputs(195)));
    layer0_outputs(3860) <= not((inputs(219)) xor (inputs(186)));
    layer0_outputs(3861) <= not((inputs(128)) xor (inputs(84)));
    layer0_outputs(3862) <= not((inputs(47)) or (inputs(22)));
    layer0_outputs(3863) <= not((inputs(228)) xor (inputs(198)));
    layer0_outputs(3864) <= not((inputs(204)) or (inputs(244)));
    layer0_outputs(3865) <= inputs(61);
    layer0_outputs(3866) <= (inputs(65)) and not (inputs(13));
    layer0_outputs(3867) <= not(inputs(156));
    layer0_outputs(3868) <= inputs(141);
    layer0_outputs(3869) <= not((inputs(6)) or (inputs(43)));
    layer0_outputs(3870) <= (inputs(236)) xor (inputs(131));
    layer0_outputs(3871) <= '1';
    layer0_outputs(3872) <= not(inputs(142)) or (inputs(94));
    layer0_outputs(3873) <= not((inputs(9)) or (inputs(170)));
    layer0_outputs(3874) <= inputs(216);
    layer0_outputs(3875) <= inputs(24);
    layer0_outputs(3876) <= not((inputs(63)) or (inputs(83)));
    layer0_outputs(3877) <= not(inputs(201));
    layer0_outputs(3878) <= not(inputs(172));
    layer0_outputs(3879) <= not(inputs(70));
    layer0_outputs(3880) <= not((inputs(141)) and (inputs(120)));
    layer0_outputs(3881) <= (inputs(107)) xor (inputs(226));
    layer0_outputs(3882) <= (inputs(219)) xor (inputs(80));
    layer0_outputs(3883) <= not((inputs(206)) and (inputs(4)));
    layer0_outputs(3884) <= (inputs(19)) or (inputs(28));
    layer0_outputs(3885) <= not(inputs(60));
    layer0_outputs(3886) <= inputs(164);
    layer0_outputs(3887) <= (inputs(66)) xor (inputs(49));
    layer0_outputs(3888) <= not((inputs(46)) or (inputs(234)));
    layer0_outputs(3889) <= inputs(194);
    layer0_outputs(3890) <= not(inputs(160));
    layer0_outputs(3891) <= (inputs(207)) or (inputs(85));
    layer0_outputs(3892) <= inputs(8);
    layer0_outputs(3893) <= inputs(237);
    layer0_outputs(3894) <= not(inputs(9));
    layer0_outputs(3895) <= not(inputs(124));
    layer0_outputs(3896) <= (inputs(178)) and not (inputs(209));
    layer0_outputs(3897) <= not(inputs(148));
    layer0_outputs(3898) <= (inputs(87)) or (inputs(252));
    layer0_outputs(3899) <= (inputs(100)) and not (inputs(240));
    layer0_outputs(3900) <= not((inputs(19)) or (inputs(243)));
    layer0_outputs(3901) <= inputs(23);
    layer0_outputs(3902) <= not(inputs(212));
    layer0_outputs(3903) <= inputs(145);
    layer0_outputs(3904) <= not((inputs(3)) or (inputs(179)));
    layer0_outputs(3905) <= not((inputs(43)) or (inputs(110)));
    layer0_outputs(3906) <= (inputs(117)) and not (inputs(179));
    layer0_outputs(3907) <= not(inputs(243));
    layer0_outputs(3908) <= not(inputs(248));
    layer0_outputs(3909) <= (inputs(135)) and not (inputs(54));
    layer0_outputs(3910) <= not((inputs(202)) or (inputs(1)));
    layer0_outputs(3911) <= not((inputs(95)) xor (inputs(17)));
    layer0_outputs(3912) <= not((inputs(252)) or (inputs(208)));
    layer0_outputs(3913) <= not(inputs(82));
    layer0_outputs(3914) <= not(inputs(201)) or (inputs(16));
    layer0_outputs(3915) <= inputs(133);
    layer0_outputs(3916) <= not((inputs(65)) and (inputs(140)));
    layer0_outputs(3917) <= not(inputs(127)) or (inputs(13));
    layer0_outputs(3918) <= not(inputs(196)) or (inputs(6));
    layer0_outputs(3919) <= not((inputs(252)) or (inputs(137)));
    layer0_outputs(3920) <= (inputs(71)) or (inputs(25));
    layer0_outputs(3921) <= not(inputs(79)) or (inputs(250));
    layer0_outputs(3922) <= not((inputs(122)) or (inputs(119)));
    layer0_outputs(3923) <= not(inputs(173));
    layer0_outputs(3924) <= not((inputs(123)) or (inputs(69)));
    layer0_outputs(3925) <= inputs(130);
    layer0_outputs(3926) <= not(inputs(70)) or (inputs(221));
    layer0_outputs(3927) <= not((inputs(77)) or (inputs(53)));
    layer0_outputs(3928) <= (inputs(53)) or (inputs(108));
    layer0_outputs(3929) <= not(inputs(141));
    layer0_outputs(3930) <= not(inputs(234));
    layer0_outputs(3931) <= (inputs(133)) xor (inputs(160));
    layer0_outputs(3932) <= inputs(98);
    layer0_outputs(3933) <= (inputs(249)) xor (inputs(185));
    layer0_outputs(3934) <= not(inputs(131)) or (inputs(218));
    layer0_outputs(3935) <= not(inputs(9)) or (inputs(181));
    layer0_outputs(3936) <= inputs(250);
    layer0_outputs(3937) <= not(inputs(229));
    layer0_outputs(3938) <= not((inputs(233)) and (inputs(248)));
    layer0_outputs(3939) <= (inputs(103)) and not (inputs(86));
    layer0_outputs(3940) <= not((inputs(203)) or (inputs(187)));
    layer0_outputs(3941) <= not((inputs(58)) or (inputs(111)));
    layer0_outputs(3942) <= not((inputs(208)) or (inputs(160)));
    layer0_outputs(3943) <= (inputs(115)) or (inputs(146));
    layer0_outputs(3944) <= not((inputs(28)) or (inputs(95)));
    layer0_outputs(3945) <= (inputs(249)) and not (inputs(237));
    layer0_outputs(3946) <= not((inputs(145)) xor (inputs(180)));
    layer0_outputs(3947) <= (inputs(220)) and not (inputs(186));
    layer0_outputs(3948) <= (inputs(235)) xor (inputs(216));
    layer0_outputs(3949) <= not((inputs(66)) and (inputs(235)));
    layer0_outputs(3950) <= not((inputs(13)) or (inputs(145)));
    layer0_outputs(3951) <= inputs(36);
    layer0_outputs(3952) <= not((inputs(226)) or (inputs(24)));
    layer0_outputs(3953) <= not(inputs(54));
    layer0_outputs(3954) <= inputs(200);
    layer0_outputs(3955) <= not(inputs(179));
    layer0_outputs(3956) <= (inputs(69)) or (inputs(71));
    layer0_outputs(3957) <= not(inputs(182));
    layer0_outputs(3958) <= (inputs(235)) or (inputs(199));
    layer0_outputs(3959) <= (inputs(117)) and not (inputs(67));
    layer0_outputs(3960) <= inputs(163);
    layer0_outputs(3961) <= (inputs(226)) or (inputs(15));
    layer0_outputs(3962) <= (inputs(50)) or (inputs(249));
    layer0_outputs(3963) <= (inputs(62)) and not (inputs(237));
    layer0_outputs(3964) <= inputs(180);
    layer0_outputs(3965) <= inputs(190);
    layer0_outputs(3966) <= (inputs(207)) xor (inputs(2));
    layer0_outputs(3967) <= not(inputs(144));
    layer0_outputs(3968) <= inputs(122);
    layer0_outputs(3969) <= inputs(15);
    layer0_outputs(3970) <= not(inputs(54));
    layer0_outputs(3971) <= not(inputs(248));
    layer0_outputs(3972) <= (inputs(133)) and not (inputs(64));
    layer0_outputs(3973) <= inputs(42);
    layer0_outputs(3974) <= not((inputs(6)) or (inputs(10)));
    layer0_outputs(3975) <= (inputs(102)) xor (inputs(149));
    layer0_outputs(3976) <= inputs(60);
    layer0_outputs(3977) <= inputs(224);
    layer0_outputs(3978) <= inputs(50);
    layer0_outputs(3979) <= inputs(63);
    layer0_outputs(3980) <= inputs(75);
    layer0_outputs(3981) <= not(inputs(169));
    layer0_outputs(3982) <= not((inputs(108)) or (inputs(109)));
    layer0_outputs(3983) <= not(inputs(105));
    layer0_outputs(3984) <= not((inputs(219)) xor (inputs(208)));
    layer0_outputs(3985) <= (inputs(225)) or (inputs(161));
    layer0_outputs(3986) <= not(inputs(212));
    layer0_outputs(3987) <= (inputs(133)) and not (inputs(126));
    layer0_outputs(3988) <= (inputs(133)) and not (inputs(110));
    layer0_outputs(3989) <= inputs(94);
    layer0_outputs(3990) <= not(inputs(20)) or (inputs(222));
    layer0_outputs(3991) <= (inputs(107)) xor (inputs(15));
    layer0_outputs(3992) <= inputs(248);
    layer0_outputs(3993) <= (inputs(205)) and not (inputs(10));
    layer0_outputs(3994) <= not((inputs(208)) and (inputs(0)));
    layer0_outputs(3995) <= not(inputs(149));
    layer0_outputs(3996) <= not(inputs(164)) or (inputs(132));
    layer0_outputs(3997) <= (inputs(242)) xor (inputs(63));
    layer0_outputs(3998) <= (inputs(120)) or (inputs(4));
    layer0_outputs(3999) <= not((inputs(161)) or (inputs(64)));
    layer0_outputs(4000) <= not(inputs(154)) or (inputs(121));
    layer0_outputs(4001) <= not(inputs(147));
    layer0_outputs(4002) <= not((inputs(79)) or (inputs(252)));
    layer0_outputs(4003) <= (inputs(59)) and not (inputs(216));
    layer0_outputs(4004) <= not((inputs(42)) or (inputs(103)));
    layer0_outputs(4005) <= (inputs(96)) xor (inputs(130));
    layer0_outputs(4006) <= (inputs(106)) xor (inputs(173));
    layer0_outputs(4007) <= not(inputs(238));
    layer0_outputs(4008) <= not(inputs(61)) or (inputs(14));
    layer0_outputs(4009) <= inputs(137);
    layer0_outputs(4010) <= not((inputs(100)) and (inputs(131)));
    layer0_outputs(4011) <= not(inputs(147));
    layer0_outputs(4012) <= inputs(162);
    layer0_outputs(4013) <= (inputs(236)) or (inputs(80));
    layer0_outputs(4014) <= not(inputs(59));
    layer0_outputs(4015) <= (inputs(114)) and not (inputs(146));
    layer0_outputs(4016) <= (inputs(61)) or (inputs(59));
    layer0_outputs(4017) <= (inputs(75)) xor (inputs(207));
    layer0_outputs(4018) <= (inputs(71)) and not (inputs(106));
    layer0_outputs(4019) <= (inputs(248)) or (inputs(127));
    layer0_outputs(4020) <= not((inputs(9)) or (inputs(213)));
    layer0_outputs(4021) <= not(inputs(116)) or (inputs(2));
    layer0_outputs(4022) <= (inputs(19)) or (inputs(33));
    layer0_outputs(4023) <= inputs(36);
    layer0_outputs(4024) <= inputs(110);
    layer0_outputs(4025) <= not(inputs(49)) or (inputs(249));
    layer0_outputs(4026) <= not((inputs(164)) or (inputs(169)));
    layer0_outputs(4027) <= inputs(69);
    layer0_outputs(4028) <= (inputs(253)) and not (inputs(175));
    layer0_outputs(4029) <= not((inputs(120)) xor (inputs(255)));
    layer0_outputs(4030) <= (inputs(246)) and not (inputs(39));
    layer0_outputs(4031) <= not((inputs(58)) or (inputs(44)));
    layer0_outputs(4032) <= inputs(141);
    layer0_outputs(4033) <= (inputs(117)) and not (inputs(80));
    layer0_outputs(4034) <= not((inputs(50)) or (inputs(255)));
    layer0_outputs(4035) <= not((inputs(49)) or (inputs(7)));
    layer0_outputs(4036) <= not(inputs(169)) or (inputs(90));
    layer0_outputs(4037) <= (inputs(64)) or (inputs(197));
    layer0_outputs(4038) <= not(inputs(247));
    layer0_outputs(4039) <= not(inputs(218)) or (inputs(95));
    layer0_outputs(4040) <= inputs(146);
    layer0_outputs(4041) <= not(inputs(230));
    layer0_outputs(4042) <= not(inputs(7));
    layer0_outputs(4043) <= not(inputs(67));
    layer0_outputs(4044) <= '1';
    layer0_outputs(4045) <= (inputs(56)) xor (inputs(54));
    layer0_outputs(4046) <= not((inputs(211)) or (inputs(247)));
    layer0_outputs(4047) <= '1';
    layer0_outputs(4048) <= not(inputs(197)) or (inputs(188));
    layer0_outputs(4049) <= not(inputs(99)) or (inputs(78));
    layer0_outputs(4050) <= (inputs(74)) or (inputs(2));
    layer0_outputs(4051) <= (inputs(78)) or (inputs(33));
    layer0_outputs(4052) <= (inputs(219)) or (inputs(111));
    layer0_outputs(4053) <= not(inputs(107));
    layer0_outputs(4054) <= (inputs(90)) and not (inputs(193));
    layer0_outputs(4055) <= inputs(224);
    layer0_outputs(4056) <= (inputs(203)) and not (inputs(125));
    layer0_outputs(4057) <= not(inputs(202));
    layer0_outputs(4058) <= not(inputs(154)) or (inputs(27));
    layer0_outputs(4059) <= not(inputs(238));
    layer0_outputs(4060) <= '1';
    layer0_outputs(4061) <= (inputs(176)) or (inputs(203));
    layer0_outputs(4062) <= not(inputs(89));
    layer0_outputs(4063) <= inputs(232);
    layer0_outputs(4064) <= not(inputs(56));
    layer0_outputs(4065) <= (inputs(209)) or (inputs(59));
    layer0_outputs(4066) <= (inputs(247)) or (inputs(195));
    layer0_outputs(4067) <= inputs(59);
    layer0_outputs(4068) <= not(inputs(91));
    layer0_outputs(4069) <= not(inputs(245)) or (inputs(125));
    layer0_outputs(4070) <= not(inputs(71));
    layer0_outputs(4071) <= inputs(205);
    layer0_outputs(4072) <= (inputs(205)) and not (inputs(166));
    layer0_outputs(4073) <= (inputs(184)) xor (inputs(185));
    layer0_outputs(4074) <= not(inputs(137)) or (inputs(175));
    layer0_outputs(4075) <= inputs(12);
    layer0_outputs(4076) <= inputs(135);
    layer0_outputs(4077) <= not(inputs(45));
    layer0_outputs(4078) <= (inputs(136)) and not (inputs(71));
    layer0_outputs(4079) <= (inputs(100)) or (inputs(108));
    layer0_outputs(4080) <= (inputs(191)) or (inputs(185));
    layer0_outputs(4081) <= not((inputs(89)) or (inputs(62)));
    layer0_outputs(4082) <= not((inputs(165)) or (inputs(32)));
    layer0_outputs(4083) <= (inputs(8)) xor (inputs(240));
    layer0_outputs(4084) <= (inputs(83)) or (inputs(158));
    layer0_outputs(4085) <= (inputs(80)) xor (inputs(224));
    layer0_outputs(4086) <= not((inputs(194)) and (inputs(110)));
    layer0_outputs(4087) <= not((inputs(179)) xor (inputs(90)));
    layer0_outputs(4088) <= not(inputs(92)) or (inputs(185));
    layer0_outputs(4089) <= (inputs(178)) or (inputs(121));
    layer0_outputs(4090) <= not((inputs(218)) xor (inputs(227)));
    layer0_outputs(4091) <= not(inputs(85));
    layer0_outputs(4092) <= not(inputs(71));
    layer0_outputs(4093) <= not(inputs(53)) or (inputs(162));
    layer0_outputs(4094) <= (inputs(222)) or (inputs(238));
    layer0_outputs(4095) <= (inputs(57)) xor (inputs(0));
    layer0_outputs(4096) <= not(inputs(39));
    layer0_outputs(4097) <= not(inputs(104)) or (inputs(198));
    layer0_outputs(4098) <= not(inputs(107));
    layer0_outputs(4099) <= (inputs(210)) xor (inputs(195));
    layer0_outputs(4100) <= '1';
    layer0_outputs(4101) <= not(inputs(41)) or (inputs(180));
    layer0_outputs(4102) <= (inputs(75)) or (inputs(205));
    layer0_outputs(4103) <= (inputs(252)) or (inputs(144));
    layer0_outputs(4104) <= (inputs(76)) xor (inputs(225));
    layer0_outputs(4105) <= not(inputs(26));
    layer0_outputs(4106) <= (inputs(53)) and not (inputs(157));
    layer0_outputs(4107) <= not(inputs(174)) or (inputs(32));
    layer0_outputs(4108) <= (inputs(88)) or (inputs(212));
    layer0_outputs(4109) <= (inputs(186)) and not (inputs(49));
    layer0_outputs(4110) <= inputs(62);
    layer0_outputs(4111) <= not((inputs(172)) or (inputs(93)));
    layer0_outputs(4112) <= '0';
    layer0_outputs(4113) <= not(inputs(51));
    layer0_outputs(4114) <= not((inputs(20)) and (inputs(22)));
    layer0_outputs(4115) <= (inputs(184)) or (inputs(205));
    layer0_outputs(4116) <= inputs(233);
    layer0_outputs(4117) <= inputs(122);
    layer0_outputs(4118) <= (inputs(36)) or (inputs(128));
    layer0_outputs(4119) <= '0';
    layer0_outputs(4120) <= inputs(97);
    layer0_outputs(4121) <= inputs(230);
    layer0_outputs(4122) <= not(inputs(170));
    layer0_outputs(4123) <= not((inputs(99)) or (inputs(70)));
    layer0_outputs(4124) <= not(inputs(112)) or (inputs(206));
    layer0_outputs(4125) <= (inputs(231)) and not (inputs(151));
    layer0_outputs(4126) <= inputs(149);
    layer0_outputs(4127) <= (inputs(163)) or (inputs(158));
    layer0_outputs(4128) <= '1';
    layer0_outputs(4129) <= not(inputs(131));
    layer0_outputs(4130) <= not(inputs(27));
    layer0_outputs(4131) <= inputs(231);
    layer0_outputs(4132) <= not(inputs(217)) or (inputs(161));
    layer0_outputs(4133) <= not(inputs(122));
    layer0_outputs(4134) <= inputs(233);
    layer0_outputs(4135) <= (inputs(28)) and (inputs(228));
    layer0_outputs(4136) <= inputs(231);
    layer0_outputs(4137) <= inputs(27);
    layer0_outputs(4138) <= not(inputs(58)) or (inputs(177));
    layer0_outputs(4139) <= not((inputs(42)) and (inputs(167)));
    layer0_outputs(4140) <= (inputs(24)) xor (inputs(255));
    layer0_outputs(4141) <= '0';
    layer0_outputs(4142) <= not(inputs(28)) or (inputs(150));
    layer0_outputs(4143) <= not(inputs(8)) or (inputs(91));
    layer0_outputs(4144) <= inputs(25);
    layer0_outputs(4145) <= inputs(147);
    layer0_outputs(4146) <= not((inputs(135)) and (inputs(51)));
    layer0_outputs(4147) <= not(inputs(2));
    layer0_outputs(4148) <= not(inputs(174));
    layer0_outputs(4149) <= inputs(63);
    layer0_outputs(4150) <= (inputs(79)) and not (inputs(107));
    layer0_outputs(4151) <= not(inputs(70));
    layer0_outputs(4152) <= (inputs(191)) or (inputs(238));
    layer0_outputs(4153) <= not(inputs(178));
    layer0_outputs(4154) <= (inputs(99)) and not (inputs(124));
    layer0_outputs(4155) <= (inputs(236)) or (inputs(170));
    layer0_outputs(4156) <= '0';
    layer0_outputs(4157) <= (inputs(176)) xor (inputs(6));
    layer0_outputs(4158) <= (inputs(90)) or (inputs(51));
    layer0_outputs(4159) <= (inputs(217)) or (inputs(254));
    layer0_outputs(4160) <= inputs(237);
    layer0_outputs(4161) <= inputs(100);
    layer0_outputs(4162) <= (inputs(151)) and not (inputs(173));
    layer0_outputs(4163) <= (inputs(207)) and not (inputs(63));
    layer0_outputs(4164) <= (inputs(148)) or (inputs(149));
    layer0_outputs(4165) <= not(inputs(126)) or (inputs(153));
    layer0_outputs(4166) <= not((inputs(206)) or (inputs(220)));
    layer0_outputs(4167) <= not(inputs(40)) or (inputs(96));
    layer0_outputs(4168) <= not((inputs(206)) or (inputs(37)));
    layer0_outputs(4169) <= not((inputs(84)) or (inputs(117)));
    layer0_outputs(4170) <= not(inputs(29)) or (inputs(239));
    layer0_outputs(4171) <= not((inputs(94)) or (inputs(217)));
    layer0_outputs(4172) <= not((inputs(96)) or (inputs(247)));
    layer0_outputs(4173) <= (inputs(10)) and not (inputs(111));
    layer0_outputs(4174) <= (inputs(227)) xor (inputs(0));
    layer0_outputs(4175) <= (inputs(152)) and (inputs(125));
    layer0_outputs(4176) <= not(inputs(178));
    layer0_outputs(4177) <= inputs(157);
    layer0_outputs(4178) <= not((inputs(190)) xor (inputs(55)));
    layer0_outputs(4179) <= inputs(194);
    layer0_outputs(4180) <= '1';
    layer0_outputs(4181) <= not((inputs(211)) or (inputs(98)));
    layer0_outputs(4182) <= (inputs(102)) xor (inputs(149));
    layer0_outputs(4183) <= inputs(103);
    layer0_outputs(4184) <= not(inputs(216)) or (inputs(41));
    layer0_outputs(4185) <= not((inputs(24)) xor (inputs(63)));
    layer0_outputs(4186) <= (inputs(248)) or (inputs(144));
    layer0_outputs(4187) <= not(inputs(189));
    layer0_outputs(4188) <= not(inputs(68));
    layer0_outputs(4189) <= not(inputs(106)) or (inputs(34));
    layer0_outputs(4190) <= (inputs(228)) and (inputs(144));
    layer0_outputs(4191) <= (inputs(5)) or (inputs(207));
    layer0_outputs(4192) <= not(inputs(103));
    layer0_outputs(4193) <= (inputs(248)) or (inputs(97));
    layer0_outputs(4194) <= (inputs(200)) or (inputs(151));
    layer0_outputs(4195) <= not(inputs(6));
    layer0_outputs(4196) <= not(inputs(23)) or (inputs(18));
    layer0_outputs(4197) <= (inputs(196)) xor (inputs(211));
    layer0_outputs(4198) <= not(inputs(143)) or (inputs(166));
    layer0_outputs(4199) <= (inputs(98)) or (inputs(115));
    layer0_outputs(4200) <= not(inputs(121)) or (inputs(184));
    layer0_outputs(4201) <= (inputs(136)) and not (inputs(109));
    layer0_outputs(4202) <= inputs(65);
    layer0_outputs(4203) <= (inputs(35)) or (inputs(229));
    layer0_outputs(4204) <= not((inputs(67)) or (inputs(24)));
    layer0_outputs(4205) <= not((inputs(104)) xor (inputs(111)));
    layer0_outputs(4206) <= inputs(83);
    layer0_outputs(4207) <= not(inputs(126));
    layer0_outputs(4208) <= (inputs(178)) or (inputs(90));
    layer0_outputs(4209) <= (inputs(53)) and (inputs(61));
    layer0_outputs(4210) <= not(inputs(73));
    layer0_outputs(4211) <= inputs(119);
    layer0_outputs(4212) <= not(inputs(94));
    layer0_outputs(4213) <= (inputs(61)) and not (inputs(88));
    layer0_outputs(4214) <= not((inputs(111)) or (inputs(31)));
    layer0_outputs(4215) <= (inputs(231)) xor (inputs(58));
    layer0_outputs(4216) <= not((inputs(88)) xor (inputs(188)));
    layer0_outputs(4217) <= not(inputs(132));
    layer0_outputs(4218) <= inputs(121);
    layer0_outputs(4219) <= (inputs(172)) and (inputs(44));
    layer0_outputs(4220) <= (inputs(118)) and not (inputs(194));
    layer0_outputs(4221) <= (inputs(161)) xor (inputs(189));
    layer0_outputs(4222) <= (inputs(219)) and not (inputs(49));
    layer0_outputs(4223) <= (inputs(93)) xor (inputs(117));
    layer0_outputs(4224) <= not(inputs(91)) or (inputs(204));
    layer0_outputs(4225) <= not(inputs(54));
    layer0_outputs(4226) <= not(inputs(55)) or (inputs(76));
    layer0_outputs(4227) <= (inputs(255)) or (inputs(137));
    layer0_outputs(4228) <= (inputs(161)) and not (inputs(48));
    layer0_outputs(4229) <= inputs(91);
    layer0_outputs(4230) <= inputs(75);
    layer0_outputs(4231) <= not(inputs(29)) or (inputs(182));
    layer0_outputs(4232) <= not((inputs(150)) xor (inputs(135)));
    layer0_outputs(4233) <= (inputs(9)) or (inputs(59));
    layer0_outputs(4234) <= inputs(18);
    layer0_outputs(4235) <= not(inputs(165));
    layer0_outputs(4236) <= not((inputs(107)) or (inputs(176)));
    layer0_outputs(4237) <= (inputs(228)) and not (inputs(143));
    layer0_outputs(4238) <= inputs(85);
    layer0_outputs(4239) <= (inputs(208)) or (inputs(196));
    layer0_outputs(4240) <= not((inputs(5)) or (inputs(141)));
    layer0_outputs(4241) <= '0';
    layer0_outputs(4242) <= not((inputs(174)) and (inputs(126)));
    layer0_outputs(4243) <= not(inputs(24));
    layer0_outputs(4244) <= '0';
    layer0_outputs(4245) <= (inputs(156)) and (inputs(78));
    layer0_outputs(4246) <= not(inputs(25));
    layer0_outputs(4247) <= inputs(79);
    layer0_outputs(4248) <= inputs(20);
    layer0_outputs(4249) <= inputs(29);
    layer0_outputs(4250) <= (inputs(84)) or (inputs(178));
    layer0_outputs(4251) <= (inputs(16)) or (inputs(79));
    layer0_outputs(4252) <= (inputs(117)) and not (inputs(162));
    layer0_outputs(4253) <= not((inputs(45)) and (inputs(91)));
    layer0_outputs(4254) <= not((inputs(209)) or (inputs(12)));
    layer0_outputs(4255) <= not(inputs(27));
    layer0_outputs(4256) <= not(inputs(27));
    layer0_outputs(4257) <= (inputs(215)) and not (inputs(33));
    layer0_outputs(4258) <= not(inputs(197)) or (inputs(118));
    layer0_outputs(4259) <= (inputs(133)) or (inputs(129));
    layer0_outputs(4260) <= (inputs(182)) or (inputs(179));
    layer0_outputs(4261) <= inputs(246);
    layer0_outputs(4262) <= not((inputs(46)) or (inputs(50)));
    layer0_outputs(4263) <= not(inputs(163));
    layer0_outputs(4264) <= (inputs(80)) or (inputs(60));
    layer0_outputs(4265) <= (inputs(238)) or (inputs(189));
    layer0_outputs(4266) <= inputs(33);
    layer0_outputs(4267) <= not((inputs(125)) and (inputs(216)));
    layer0_outputs(4268) <= not(inputs(122)) or (inputs(15));
    layer0_outputs(4269) <= (inputs(207)) xor (inputs(159));
    layer0_outputs(4270) <= inputs(116);
    layer0_outputs(4271) <= (inputs(143)) xor (inputs(104));
    layer0_outputs(4272) <= not((inputs(219)) or (inputs(138)));
    layer0_outputs(4273) <= not(inputs(171));
    layer0_outputs(4274) <= (inputs(248)) xor (inputs(80));
    layer0_outputs(4275) <= inputs(8);
    layer0_outputs(4276) <= inputs(184);
    layer0_outputs(4277) <= not(inputs(121));
    layer0_outputs(4278) <= not(inputs(42));
    layer0_outputs(4279) <= not(inputs(134)) or (inputs(144));
    layer0_outputs(4280) <= inputs(68);
    layer0_outputs(4281) <= (inputs(214)) or (inputs(150));
    layer0_outputs(4282) <= not((inputs(38)) or (inputs(201)));
    layer0_outputs(4283) <= inputs(250);
    layer0_outputs(4284) <= not(inputs(182));
    layer0_outputs(4285) <= not((inputs(91)) xor (inputs(64)));
    layer0_outputs(4286) <= not(inputs(64)) or (inputs(13));
    layer0_outputs(4287) <= not(inputs(58));
    layer0_outputs(4288) <= not(inputs(218)) or (inputs(120));
    layer0_outputs(4289) <= not(inputs(34)) or (inputs(66));
    layer0_outputs(4290) <= inputs(118);
    layer0_outputs(4291) <= not((inputs(39)) and (inputs(75)));
    layer0_outputs(4292) <= (inputs(37)) and not (inputs(158));
    layer0_outputs(4293) <= not(inputs(43));
    layer0_outputs(4294) <= not(inputs(8)) or (inputs(152));
    layer0_outputs(4295) <= not(inputs(129));
    layer0_outputs(4296) <= not(inputs(152));
    layer0_outputs(4297) <= (inputs(133)) or (inputs(240));
    layer0_outputs(4298) <= (inputs(103)) and not (inputs(166));
    layer0_outputs(4299) <= not(inputs(247));
    layer0_outputs(4300) <= inputs(120);
    layer0_outputs(4301) <= inputs(226);
    layer0_outputs(4302) <= not(inputs(83));
    layer0_outputs(4303) <= not(inputs(135));
    layer0_outputs(4304) <= not(inputs(140));
    layer0_outputs(4305) <= not(inputs(43)) or (inputs(231));
    layer0_outputs(4306) <= not(inputs(236));
    layer0_outputs(4307) <= (inputs(165)) or (inputs(47));
    layer0_outputs(4308) <= (inputs(117)) or (inputs(197));
    layer0_outputs(4309) <= not(inputs(114));
    layer0_outputs(4310) <= not((inputs(209)) or (inputs(238)));
    layer0_outputs(4311) <= (inputs(191)) and not (inputs(221));
    layer0_outputs(4312) <= not((inputs(249)) and (inputs(183)));
    layer0_outputs(4313) <= not((inputs(56)) and (inputs(110)));
    layer0_outputs(4314) <= (inputs(162)) or (inputs(238));
    layer0_outputs(4315) <= (inputs(146)) and not (inputs(225));
    layer0_outputs(4316) <= inputs(67);
    layer0_outputs(4317) <= inputs(125);
    layer0_outputs(4318) <= inputs(86);
    layer0_outputs(4319) <= '0';
    layer0_outputs(4320) <= not(inputs(117)) or (inputs(8));
    layer0_outputs(4321) <= (inputs(16)) and (inputs(150));
    layer0_outputs(4322) <= not((inputs(148)) xor (inputs(167)));
    layer0_outputs(4323) <= not(inputs(41));
    layer0_outputs(4324) <= not(inputs(45)) or (inputs(109));
    layer0_outputs(4325) <= (inputs(218)) and not (inputs(152));
    layer0_outputs(4326) <= (inputs(113)) or (inputs(110));
    layer0_outputs(4327) <= (inputs(152)) and not (inputs(20));
    layer0_outputs(4328) <= inputs(81);
    layer0_outputs(4329) <= not(inputs(255)) or (inputs(220));
    layer0_outputs(4330) <= (inputs(72)) xor (inputs(4));
    layer0_outputs(4331) <= inputs(30);
    layer0_outputs(4332) <= (inputs(57)) or (inputs(242));
    layer0_outputs(4333) <= inputs(90);
    layer0_outputs(4334) <= not(inputs(120)) or (inputs(170));
    layer0_outputs(4335) <= (inputs(219)) or (inputs(31));
    layer0_outputs(4336) <= (inputs(116)) and not (inputs(237));
    layer0_outputs(4337) <= inputs(21);
    layer0_outputs(4338) <= (inputs(12)) and (inputs(37));
    layer0_outputs(4339) <= (inputs(254)) or (inputs(150));
    layer0_outputs(4340) <= not(inputs(135)) or (inputs(224));
    layer0_outputs(4341) <= not(inputs(85));
    layer0_outputs(4342) <= (inputs(4)) and not (inputs(190));
    layer0_outputs(4343) <= (inputs(231)) and not (inputs(173));
    layer0_outputs(4344) <= inputs(157);
    layer0_outputs(4345) <= not((inputs(102)) or (inputs(193)));
    layer0_outputs(4346) <= not(inputs(53));
    layer0_outputs(4347) <= inputs(236);
    layer0_outputs(4348) <= '1';
    layer0_outputs(4349) <= inputs(245);
    layer0_outputs(4350) <= (inputs(201)) and (inputs(246));
    layer0_outputs(4351) <= inputs(216);
    layer0_outputs(4352) <= not(inputs(120)) or (inputs(20));
    layer0_outputs(4353) <= (inputs(116)) and not (inputs(242));
    layer0_outputs(4354) <= not(inputs(63)) or (inputs(123));
    layer0_outputs(4355) <= not(inputs(86));
    layer0_outputs(4356) <= not(inputs(179));
    layer0_outputs(4357) <= inputs(177);
    layer0_outputs(4358) <= (inputs(28)) and not (inputs(72));
    layer0_outputs(4359) <= not((inputs(126)) or (inputs(163)));
    layer0_outputs(4360) <= (inputs(105)) and not (inputs(237));
    layer0_outputs(4361) <= not((inputs(90)) or (inputs(76)));
    layer0_outputs(4362) <= inputs(100);
    layer0_outputs(4363) <= not(inputs(65));
    layer0_outputs(4364) <= not((inputs(229)) or (inputs(222)));
    layer0_outputs(4365) <= not((inputs(227)) or (inputs(224)));
    layer0_outputs(4366) <= (inputs(29)) and not (inputs(48));
    layer0_outputs(4367) <= '0';
    layer0_outputs(4368) <= not((inputs(31)) or (inputs(213)));
    layer0_outputs(4369) <= not(inputs(229)) or (inputs(19));
    layer0_outputs(4370) <= (inputs(227)) or (inputs(169));
    layer0_outputs(4371) <= (inputs(81)) or (inputs(128));
    layer0_outputs(4372) <= inputs(194);
    layer0_outputs(4373) <= not(inputs(37));
    layer0_outputs(4374) <= (inputs(36)) and (inputs(160));
    layer0_outputs(4375) <= not((inputs(62)) or (inputs(171)));
    layer0_outputs(4376) <= (inputs(223)) and not (inputs(15));
    layer0_outputs(4377) <= (inputs(47)) or (inputs(226));
    layer0_outputs(4378) <= not((inputs(144)) or (inputs(172)));
    layer0_outputs(4379) <= not(inputs(99));
    layer0_outputs(4380) <= (inputs(214)) xor (inputs(6));
    layer0_outputs(4381) <= not(inputs(80)) or (inputs(65));
    layer0_outputs(4382) <= not((inputs(26)) or (inputs(17)));
    layer0_outputs(4383) <= not(inputs(9));
    layer0_outputs(4384) <= not(inputs(73)) or (inputs(22));
    layer0_outputs(4385) <= not(inputs(113));
    layer0_outputs(4386) <= not(inputs(248));
    layer0_outputs(4387) <= (inputs(32)) or (inputs(23));
    layer0_outputs(4388) <= not((inputs(161)) or (inputs(245)));
    layer0_outputs(4389) <= (inputs(21)) and not (inputs(70));
    layer0_outputs(4390) <= inputs(105);
    layer0_outputs(4391) <= not(inputs(74));
    layer0_outputs(4392) <= not(inputs(179));
    layer0_outputs(4393) <= inputs(151);
    layer0_outputs(4394) <= not((inputs(21)) and (inputs(51)));
    layer0_outputs(4395) <= (inputs(201)) and not (inputs(64));
    layer0_outputs(4396) <= not(inputs(158)) or (inputs(196));
    layer0_outputs(4397) <= not(inputs(106));
    layer0_outputs(4398) <= not((inputs(178)) xor (inputs(62)));
    layer0_outputs(4399) <= not((inputs(59)) xor (inputs(225)));
    layer0_outputs(4400) <= not((inputs(72)) or (inputs(230)));
    layer0_outputs(4401) <= not(inputs(76));
    layer0_outputs(4402) <= not(inputs(218)) or (inputs(66));
    layer0_outputs(4403) <= (inputs(231)) and not (inputs(59));
    layer0_outputs(4404) <= (inputs(148)) or (inputs(133));
    layer0_outputs(4405) <= not(inputs(151));
    layer0_outputs(4406) <= (inputs(105)) and not (inputs(36));
    layer0_outputs(4407) <= (inputs(120)) and not (inputs(254));
    layer0_outputs(4408) <= not((inputs(197)) and (inputs(186)));
    layer0_outputs(4409) <= not(inputs(41)) or (inputs(32));
    layer0_outputs(4410) <= not(inputs(60));
    layer0_outputs(4411) <= '1';
    layer0_outputs(4412) <= not(inputs(167));
    layer0_outputs(4413) <= inputs(15);
    layer0_outputs(4414) <= (inputs(151)) and not (inputs(61));
    layer0_outputs(4415) <= (inputs(123)) and not (inputs(192));
    layer0_outputs(4416) <= not(inputs(196)) or (inputs(155));
    layer0_outputs(4417) <= (inputs(162)) or (inputs(39));
    layer0_outputs(4418) <= (inputs(115)) or (inputs(52));
    layer0_outputs(4419) <= not(inputs(248)) or (inputs(95));
    layer0_outputs(4420) <= not(inputs(41));
    layer0_outputs(4421) <= not((inputs(16)) or (inputs(93)));
    layer0_outputs(4422) <= not((inputs(173)) or (inputs(126)));
    layer0_outputs(4423) <= inputs(85);
    layer0_outputs(4424) <= not(inputs(28));
    layer0_outputs(4425) <= not((inputs(189)) xor (inputs(104)));
    layer0_outputs(4426) <= not(inputs(196)) or (inputs(62));
    layer0_outputs(4427) <= (inputs(136)) and not (inputs(210));
    layer0_outputs(4428) <= not((inputs(253)) or (inputs(152)));
    layer0_outputs(4429) <= not(inputs(137)) or (inputs(254));
    layer0_outputs(4430) <= not(inputs(239));
    layer0_outputs(4431) <= not((inputs(143)) or (inputs(92)));
    layer0_outputs(4432) <= (inputs(22)) and not (inputs(236));
    layer0_outputs(4433) <= '0';
    layer0_outputs(4434) <= (inputs(44)) or (inputs(239));
    layer0_outputs(4435) <= not(inputs(150)) or (inputs(54));
    layer0_outputs(4436) <= inputs(24);
    layer0_outputs(4437) <= (inputs(28)) and not (inputs(147));
    layer0_outputs(4438) <= (inputs(232)) and not (inputs(95));
    layer0_outputs(4439) <= not(inputs(116)) or (inputs(95));
    layer0_outputs(4440) <= not(inputs(246));
    layer0_outputs(4441) <= not(inputs(56));
    layer0_outputs(4442) <= (inputs(252)) or (inputs(82));
    layer0_outputs(4443) <= not(inputs(114));
    layer0_outputs(4444) <= (inputs(153)) or (inputs(192));
    layer0_outputs(4445) <= not((inputs(97)) or (inputs(96)));
    layer0_outputs(4446) <= (inputs(142)) and not (inputs(2));
    layer0_outputs(4447) <= not(inputs(246));
    layer0_outputs(4448) <= (inputs(149)) and (inputs(189));
    layer0_outputs(4449) <= inputs(83);
    layer0_outputs(4450) <= not(inputs(247)) or (inputs(16));
    layer0_outputs(4451) <= not((inputs(41)) xor (inputs(72)));
    layer0_outputs(4452) <= not((inputs(161)) or (inputs(53)));
    layer0_outputs(4453) <= not(inputs(122)) or (inputs(239));
    layer0_outputs(4454) <= not((inputs(72)) xor (inputs(80)));
    layer0_outputs(4455) <= inputs(162);
    layer0_outputs(4456) <= '1';
    layer0_outputs(4457) <= inputs(144);
    layer0_outputs(4458) <= not(inputs(219));
    layer0_outputs(4459) <= '1';
    layer0_outputs(4460) <= not(inputs(189));
    layer0_outputs(4461) <= (inputs(171)) or (inputs(188));
    layer0_outputs(4462) <= inputs(161);
    layer0_outputs(4463) <= not(inputs(36));
    layer0_outputs(4464) <= (inputs(20)) and not (inputs(251));
    layer0_outputs(4465) <= not(inputs(121));
    layer0_outputs(4466) <= (inputs(100)) and not (inputs(239));
    layer0_outputs(4467) <= (inputs(56)) xor (inputs(114));
    layer0_outputs(4468) <= inputs(62);
    layer0_outputs(4469) <= inputs(118);
    layer0_outputs(4470) <= not(inputs(137)) or (inputs(180));
    layer0_outputs(4471) <= inputs(178);
    layer0_outputs(4472) <= not((inputs(16)) xor (inputs(153)));
    layer0_outputs(4473) <= not(inputs(165));
    layer0_outputs(4474) <= '1';
    layer0_outputs(4475) <= (inputs(241)) or (inputs(220));
    layer0_outputs(4476) <= not(inputs(215));
    layer0_outputs(4477) <= not((inputs(131)) xor (inputs(175)));
    layer0_outputs(4478) <= not(inputs(216));
    layer0_outputs(4479) <= not(inputs(244)) or (inputs(7));
    layer0_outputs(4480) <= not((inputs(5)) or (inputs(64)));
    layer0_outputs(4481) <= inputs(39);
    layer0_outputs(4482) <= not(inputs(203));
    layer0_outputs(4483) <= not((inputs(79)) or (inputs(45)));
    layer0_outputs(4484) <= not((inputs(219)) or (inputs(228)));
    layer0_outputs(4485) <= not(inputs(215)) or (inputs(14));
    layer0_outputs(4486) <= not((inputs(2)) or (inputs(41)));
    layer0_outputs(4487) <= (inputs(170)) and not (inputs(17));
    layer0_outputs(4488) <= not((inputs(150)) xor (inputs(120)));
    layer0_outputs(4489) <= (inputs(187)) and not (inputs(1));
    layer0_outputs(4490) <= inputs(20);
    layer0_outputs(4491) <= (inputs(181)) and not (inputs(13));
    layer0_outputs(4492) <= not(inputs(84));
    layer0_outputs(4493) <= inputs(213);
    layer0_outputs(4494) <= not(inputs(252));
    layer0_outputs(4495) <= '1';
    layer0_outputs(4496) <= (inputs(21)) or (inputs(45));
    layer0_outputs(4497) <= not(inputs(146));
    layer0_outputs(4498) <= not(inputs(237)) or (inputs(208));
    layer0_outputs(4499) <= inputs(100);
    layer0_outputs(4500) <= not((inputs(233)) or (inputs(132)));
    layer0_outputs(4501) <= (inputs(183)) and not (inputs(118));
    layer0_outputs(4502) <= not(inputs(21));
    layer0_outputs(4503) <= not(inputs(237));
    layer0_outputs(4504) <= (inputs(188)) or (inputs(145));
    layer0_outputs(4505) <= (inputs(228)) or (inputs(205));
    layer0_outputs(4506) <= not(inputs(168));
    layer0_outputs(4507) <= inputs(52);
    layer0_outputs(4508) <= inputs(247);
    layer0_outputs(4509) <= not(inputs(248));
    layer0_outputs(4510) <= (inputs(37)) and not (inputs(206));
    layer0_outputs(4511) <= (inputs(56)) or (inputs(172));
    layer0_outputs(4512) <= (inputs(161)) and not (inputs(254));
    layer0_outputs(4513) <= not(inputs(168)) or (inputs(161));
    layer0_outputs(4514) <= not((inputs(57)) or (inputs(34)));
    layer0_outputs(4515) <= (inputs(120)) and not (inputs(145));
    layer0_outputs(4516) <= not(inputs(145)) or (inputs(191));
    layer0_outputs(4517) <= inputs(7);
    layer0_outputs(4518) <= (inputs(198)) or (inputs(75));
    layer0_outputs(4519) <= inputs(85);
    layer0_outputs(4520) <= inputs(157);
    layer0_outputs(4521) <= inputs(229);
    layer0_outputs(4522) <= (inputs(34)) or (inputs(225));
    layer0_outputs(4523) <= inputs(187);
    layer0_outputs(4524) <= inputs(136);
    layer0_outputs(4525) <= not(inputs(69));
    layer0_outputs(4526) <= not((inputs(148)) or (inputs(190)));
    layer0_outputs(4527) <= not(inputs(106)) or (inputs(177));
    layer0_outputs(4528) <= (inputs(133)) and not (inputs(179));
    layer0_outputs(4529) <= inputs(47);
    layer0_outputs(4530) <= not(inputs(210));
    layer0_outputs(4531) <= not(inputs(154)) or (inputs(1));
    layer0_outputs(4532) <= not((inputs(157)) and (inputs(105)));
    layer0_outputs(4533) <= (inputs(115)) or (inputs(253));
    layer0_outputs(4534) <= not((inputs(10)) and (inputs(38)));
    layer0_outputs(4535) <= inputs(115);
    layer0_outputs(4536) <= inputs(202);
    layer0_outputs(4537) <= (inputs(198)) and not (inputs(206));
    layer0_outputs(4538) <= not((inputs(70)) or (inputs(211)));
    layer0_outputs(4539) <= not((inputs(204)) xor (inputs(124)));
    layer0_outputs(4540) <= not((inputs(231)) or (inputs(209)));
    layer0_outputs(4541) <= not((inputs(27)) or (inputs(61)));
    layer0_outputs(4542) <= (inputs(239)) or (inputs(148));
    layer0_outputs(4543) <= (inputs(236)) and not (inputs(4));
    layer0_outputs(4544) <= inputs(167);
    layer0_outputs(4545) <= not(inputs(182)) or (inputs(120));
    layer0_outputs(4546) <= not(inputs(152)) or (inputs(185));
    layer0_outputs(4547) <= (inputs(98)) or (inputs(104));
    layer0_outputs(4548) <= not(inputs(132));
    layer0_outputs(4549) <= (inputs(98)) and not (inputs(74));
    layer0_outputs(4550) <= not((inputs(204)) or (inputs(213)));
    layer0_outputs(4551) <= inputs(150);
    layer0_outputs(4552) <= not(inputs(166));
    layer0_outputs(4553) <= '0';
    layer0_outputs(4554) <= (inputs(92)) and not (inputs(142));
    layer0_outputs(4555) <= not((inputs(99)) xor (inputs(86)));
    layer0_outputs(4556) <= inputs(66);
    layer0_outputs(4557) <= not(inputs(68));
    layer0_outputs(4558) <= not(inputs(97));
    layer0_outputs(4559) <= inputs(112);
    layer0_outputs(4560) <= (inputs(139)) and (inputs(132));
    layer0_outputs(4561) <= not(inputs(114));
    layer0_outputs(4562) <= inputs(56);
    layer0_outputs(4563) <= '0';
    layer0_outputs(4564) <= (inputs(69)) and (inputs(25));
    layer0_outputs(4565) <= (inputs(132)) or (inputs(247));
    layer0_outputs(4566) <= '1';
    layer0_outputs(4567) <= inputs(186);
    layer0_outputs(4568) <= not(inputs(66));
    layer0_outputs(4569) <= (inputs(177)) xor (inputs(76));
    layer0_outputs(4570) <= not((inputs(244)) or (inputs(64)));
    layer0_outputs(4571) <= not((inputs(44)) or (inputs(7)));
    layer0_outputs(4572) <= (inputs(43)) or (inputs(67));
    layer0_outputs(4573) <= (inputs(232)) and not (inputs(193));
    layer0_outputs(4574) <= not(inputs(146)) or (inputs(43));
    layer0_outputs(4575) <= not(inputs(23));
    layer0_outputs(4576) <= (inputs(46)) or (inputs(119));
    layer0_outputs(4577) <= '0';
    layer0_outputs(4578) <= not(inputs(82));
    layer0_outputs(4579) <= not((inputs(214)) and (inputs(0)));
    layer0_outputs(4580) <= inputs(9);
    layer0_outputs(4581) <= (inputs(224)) or (inputs(45));
    layer0_outputs(4582) <= not(inputs(193));
    layer0_outputs(4583) <= inputs(116);
    layer0_outputs(4584) <= (inputs(29)) and not (inputs(81));
    layer0_outputs(4585) <= not((inputs(212)) or (inputs(68)));
    layer0_outputs(4586) <= not(inputs(188)) or (inputs(111));
    layer0_outputs(4587) <= (inputs(198)) or (inputs(125));
    layer0_outputs(4588) <= (inputs(65)) or (inputs(220));
    layer0_outputs(4589) <= (inputs(77)) or (inputs(163));
    layer0_outputs(4590) <= inputs(182);
    layer0_outputs(4591) <= (inputs(190)) and (inputs(105));
    layer0_outputs(4592) <= not(inputs(233));
    layer0_outputs(4593) <= not(inputs(164));
    layer0_outputs(4594) <= not(inputs(154)) or (inputs(102));
    layer0_outputs(4595) <= not(inputs(105)) or (inputs(99));
    layer0_outputs(4596) <= not(inputs(10)) or (inputs(144));
    layer0_outputs(4597) <= (inputs(244)) xor (inputs(55));
    layer0_outputs(4598) <= not(inputs(172));
    layer0_outputs(4599) <= not(inputs(143));
    layer0_outputs(4600) <= (inputs(58)) or (inputs(125));
    layer0_outputs(4601) <= inputs(115);
    layer0_outputs(4602) <= (inputs(20)) and not (inputs(8));
    layer0_outputs(4603) <= (inputs(163)) and (inputs(140));
    layer0_outputs(4604) <= inputs(150);
    layer0_outputs(4605) <= inputs(237);
    layer0_outputs(4606) <= not((inputs(39)) or (inputs(36)));
    layer0_outputs(4607) <= not(inputs(123));
    layer0_outputs(4608) <= not(inputs(104));
    layer0_outputs(4609) <= not((inputs(69)) xor (inputs(49)));
    layer0_outputs(4610) <= not((inputs(231)) or (inputs(202)));
    layer0_outputs(4611) <= (inputs(62)) and not (inputs(164));
    layer0_outputs(4612) <= not(inputs(103));
    layer0_outputs(4613) <= '0';
    layer0_outputs(4614) <= (inputs(106)) or (inputs(51));
    layer0_outputs(4615) <= not((inputs(239)) or (inputs(217)));
    layer0_outputs(4616) <= not(inputs(138)) or (inputs(222));
    layer0_outputs(4617) <= not(inputs(99));
    layer0_outputs(4618) <= inputs(199);
    layer0_outputs(4619) <= not(inputs(245)) or (inputs(252));
    layer0_outputs(4620) <= '0';
    layer0_outputs(4621) <= not(inputs(109)) or (inputs(203));
    layer0_outputs(4622) <= inputs(137);
    layer0_outputs(4623) <= not(inputs(67));
    layer0_outputs(4624) <= not(inputs(93));
    layer0_outputs(4625) <= not((inputs(172)) xor (inputs(220)));
    layer0_outputs(4626) <= inputs(217);
    layer0_outputs(4627) <= inputs(220);
    layer0_outputs(4628) <= (inputs(165)) and (inputs(231));
    layer0_outputs(4629) <= (inputs(130)) or (inputs(154));
    layer0_outputs(4630) <= not(inputs(20)) or (inputs(177));
    layer0_outputs(4631) <= (inputs(30)) and not (inputs(158));
    layer0_outputs(4632) <= (inputs(185)) or (inputs(240));
    layer0_outputs(4633) <= inputs(191);
    layer0_outputs(4634) <= not((inputs(35)) or (inputs(252)));
    layer0_outputs(4635) <= (inputs(151)) and not (inputs(26));
    layer0_outputs(4636) <= (inputs(123)) or (inputs(35));
    layer0_outputs(4637) <= not(inputs(105));
    layer0_outputs(4638) <= not(inputs(172));
    layer0_outputs(4639) <= (inputs(131)) and not (inputs(119));
    layer0_outputs(4640) <= (inputs(156)) and not (inputs(236));
    layer0_outputs(4641) <= (inputs(22)) and not (inputs(131));
    layer0_outputs(4642) <= not(inputs(226)) or (inputs(96));
    layer0_outputs(4643) <= inputs(26);
    layer0_outputs(4644) <= not(inputs(108));
    layer0_outputs(4645) <= not(inputs(104));
    layer0_outputs(4646) <= not((inputs(146)) xor (inputs(134)));
    layer0_outputs(4647) <= not(inputs(107)) or (inputs(205));
    layer0_outputs(4648) <= inputs(160);
    layer0_outputs(4649) <= inputs(232);
    layer0_outputs(4650) <= not(inputs(45));
    layer0_outputs(4651) <= inputs(183);
    layer0_outputs(4652) <= inputs(110);
    layer0_outputs(4653) <= inputs(253);
    layer0_outputs(4654) <= not((inputs(116)) or (inputs(100)));
    layer0_outputs(4655) <= not(inputs(237));
    layer0_outputs(4656) <= not(inputs(89));
    layer0_outputs(4657) <= not((inputs(36)) or (inputs(15)));
    layer0_outputs(4658) <= (inputs(25)) and (inputs(116));
    layer0_outputs(4659) <= (inputs(51)) or (inputs(91));
    layer0_outputs(4660) <= (inputs(156)) or (inputs(177));
    layer0_outputs(4661) <= not((inputs(220)) or (inputs(95)));
    layer0_outputs(4662) <= not((inputs(84)) or (inputs(29)));
    layer0_outputs(4663) <= (inputs(87)) and not (inputs(135));
    layer0_outputs(4664) <= (inputs(35)) or (inputs(55));
    layer0_outputs(4665) <= not(inputs(168));
    layer0_outputs(4666) <= (inputs(217)) and not (inputs(15));
    layer0_outputs(4667) <= not(inputs(161));
    layer0_outputs(4668) <= (inputs(141)) and not (inputs(65));
    layer0_outputs(4669) <= (inputs(40)) and not (inputs(146));
    layer0_outputs(4670) <= (inputs(33)) or (inputs(196));
    layer0_outputs(4671) <= not(inputs(15));
    layer0_outputs(4672) <= not((inputs(177)) or (inputs(21)));
    layer0_outputs(4673) <= not(inputs(101));
    layer0_outputs(4674) <= (inputs(227)) and not (inputs(31));
    layer0_outputs(4675) <= not(inputs(210));
    layer0_outputs(4676) <= not(inputs(81)) or (inputs(95));
    layer0_outputs(4677) <= (inputs(235)) or (inputs(217));
    layer0_outputs(4678) <= not(inputs(166));
    layer0_outputs(4679) <= inputs(90);
    layer0_outputs(4680) <= not(inputs(17));
    layer0_outputs(4681) <= not((inputs(35)) or (inputs(46)));
    layer0_outputs(4682) <= inputs(204);
    layer0_outputs(4683) <= not((inputs(8)) or (inputs(78)));
    layer0_outputs(4684) <= not((inputs(47)) or (inputs(78)));
    layer0_outputs(4685) <= not(inputs(27)) or (inputs(114));
    layer0_outputs(4686) <= not(inputs(55));
    layer0_outputs(4687) <= not(inputs(197));
    layer0_outputs(4688) <= not(inputs(122)) or (inputs(229));
    layer0_outputs(4689) <= (inputs(136)) and not (inputs(125));
    layer0_outputs(4690) <= inputs(119);
    layer0_outputs(4691) <= inputs(136);
    layer0_outputs(4692) <= not(inputs(45)) or (inputs(204));
    layer0_outputs(4693) <= inputs(222);
    layer0_outputs(4694) <= not((inputs(99)) xor (inputs(117)));
    layer0_outputs(4695) <= inputs(177);
    layer0_outputs(4696) <= not(inputs(224)) or (inputs(251));
    layer0_outputs(4697) <= not((inputs(160)) xor (inputs(204)));
    layer0_outputs(4698) <= (inputs(199)) or (inputs(252));
    layer0_outputs(4699) <= (inputs(191)) or (inputs(71));
    layer0_outputs(4700) <= (inputs(167)) and not (inputs(100));
    layer0_outputs(4701) <= (inputs(169)) and not (inputs(46));
    layer0_outputs(4702) <= (inputs(120)) and (inputs(104));
    layer0_outputs(4703) <= (inputs(110)) or (inputs(144));
    layer0_outputs(4704) <= not(inputs(146));
    layer0_outputs(4705) <= inputs(151);
    layer0_outputs(4706) <= (inputs(93)) or (inputs(7));
    layer0_outputs(4707) <= (inputs(70)) or (inputs(85));
    layer0_outputs(4708) <= (inputs(101)) and not (inputs(206));
    layer0_outputs(4709) <= (inputs(148)) xor (inputs(158));
    layer0_outputs(4710) <= (inputs(198)) and not (inputs(143));
    layer0_outputs(4711) <= not(inputs(55));
    layer0_outputs(4712) <= (inputs(170)) and not (inputs(50));
    layer0_outputs(4713) <= not(inputs(75)) or (inputs(175));
    layer0_outputs(4714) <= (inputs(206)) and not (inputs(111));
    layer0_outputs(4715) <= inputs(148);
    layer0_outputs(4716) <= inputs(179);
    layer0_outputs(4717) <= inputs(0);
    layer0_outputs(4718) <= not((inputs(207)) xor (inputs(11)));
    layer0_outputs(4719) <= not(inputs(228)) or (inputs(78));
    layer0_outputs(4720) <= not((inputs(217)) or (inputs(223)));
    layer0_outputs(4721) <= (inputs(243)) and (inputs(234));
    layer0_outputs(4722) <= not((inputs(43)) or (inputs(45)));
    layer0_outputs(4723) <= not((inputs(191)) or (inputs(231)));
    layer0_outputs(4724) <= not(inputs(27)) or (inputs(239));
    layer0_outputs(4725) <= not(inputs(8));
    layer0_outputs(4726) <= not((inputs(204)) and (inputs(104)));
    layer0_outputs(4727) <= (inputs(38)) or (inputs(92));
    layer0_outputs(4728) <= not(inputs(210)) or (inputs(30));
    layer0_outputs(4729) <= (inputs(15)) or (inputs(56));
    layer0_outputs(4730) <= not(inputs(204));
    layer0_outputs(4731) <= (inputs(246)) or (inputs(29));
    layer0_outputs(4732) <= (inputs(205)) or (inputs(191));
    layer0_outputs(4733) <= (inputs(2)) and not (inputs(222));
    layer0_outputs(4734) <= not((inputs(146)) or (inputs(86)));
    layer0_outputs(4735) <= (inputs(17)) or (inputs(129));
    layer0_outputs(4736) <= not(inputs(175));
    layer0_outputs(4737) <= inputs(9);
    layer0_outputs(4738) <= '1';
    layer0_outputs(4739) <= (inputs(225)) and not (inputs(131));
    layer0_outputs(4740) <= (inputs(88)) and (inputs(98));
    layer0_outputs(4741) <= not(inputs(76));
    layer0_outputs(4742) <= '0';
    layer0_outputs(4743) <= inputs(131);
    layer0_outputs(4744) <= not((inputs(142)) and (inputs(136)));
    layer0_outputs(4745) <= inputs(60);
    layer0_outputs(4746) <= (inputs(180)) or (inputs(104));
    layer0_outputs(4747) <= '0';
    layer0_outputs(4748) <= inputs(98);
    layer0_outputs(4749) <= (inputs(52)) xor (inputs(186));
    layer0_outputs(4750) <= (inputs(36)) or (inputs(218));
    layer0_outputs(4751) <= (inputs(90)) xor (inputs(138));
    layer0_outputs(4752) <= (inputs(158)) or (inputs(205));
    layer0_outputs(4753) <= (inputs(65)) and not (inputs(97));
    layer0_outputs(4754) <= '0';
    layer0_outputs(4755) <= not((inputs(189)) xor (inputs(124)));
    layer0_outputs(4756) <= not((inputs(181)) or (inputs(202)));
    layer0_outputs(4757) <= not(inputs(149));
    layer0_outputs(4758) <= not(inputs(252));
    layer0_outputs(4759) <= not(inputs(85));
    layer0_outputs(4760) <= (inputs(8)) and (inputs(30));
    layer0_outputs(4761) <= (inputs(131)) xor (inputs(21));
    layer0_outputs(4762) <= not(inputs(90));
    layer0_outputs(4763) <= (inputs(183)) and (inputs(74));
    layer0_outputs(4764) <= not((inputs(190)) or (inputs(129)));
    layer0_outputs(4765) <= (inputs(170)) or (inputs(100));
    layer0_outputs(4766) <= (inputs(104)) and not (inputs(109));
    layer0_outputs(4767) <= inputs(76);
    layer0_outputs(4768) <= (inputs(109)) and not (inputs(35));
    layer0_outputs(4769) <= not(inputs(73));
    layer0_outputs(4770) <= (inputs(134)) and not (inputs(17));
    layer0_outputs(4771) <= not(inputs(117)) or (inputs(73));
    layer0_outputs(4772) <= (inputs(163)) or (inputs(187));
    layer0_outputs(4773) <= (inputs(250)) and (inputs(157));
    layer0_outputs(4774) <= inputs(59);
    layer0_outputs(4775) <= not(inputs(119));
    layer0_outputs(4776) <= (inputs(71)) and not (inputs(103));
    layer0_outputs(4777) <= inputs(210);
    layer0_outputs(4778) <= not((inputs(230)) or (inputs(194)));
    layer0_outputs(4779) <= (inputs(135)) and not (inputs(53));
    layer0_outputs(4780) <= inputs(154);
    layer0_outputs(4781) <= not((inputs(174)) or (inputs(194)));
    layer0_outputs(4782) <= not(inputs(171));
    layer0_outputs(4783) <= (inputs(174)) or (inputs(192));
    layer0_outputs(4784) <= (inputs(157)) or (inputs(163));
    layer0_outputs(4785) <= not((inputs(69)) xor (inputs(238)));
    layer0_outputs(4786) <= '0';
    layer0_outputs(4787) <= not(inputs(170));
    layer0_outputs(4788) <= not(inputs(119)) or (inputs(155));
    layer0_outputs(4789) <= (inputs(118)) or (inputs(208));
    layer0_outputs(4790) <= not((inputs(207)) xor (inputs(7)));
    layer0_outputs(4791) <= (inputs(230)) and not (inputs(31));
    layer0_outputs(4792) <= inputs(140);
    layer0_outputs(4793) <= (inputs(32)) xor (inputs(76));
    layer0_outputs(4794) <= (inputs(104)) and not (inputs(160));
    layer0_outputs(4795) <= (inputs(13)) and not (inputs(87));
    layer0_outputs(4796) <= (inputs(80)) xor (inputs(165));
    layer0_outputs(4797) <= inputs(103);
    layer0_outputs(4798) <= not(inputs(215));
    layer0_outputs(4799) <= not((inputs(173)) or (inputs(206)));
    layer0_outputs(4800) <= not(inputs(217));
    layer0_outputs(4801) <= inputs(163);
    layer0_outputs(4802) <= not(inputs(180));
    layer0_outputs(4803) <= (inputs(82)) and not (inputs(148));
    layer0_outputs(4804) <= (inputs(199)) or (inputs(165));
    layer0_outputs(4805) <= not((inputs(55)) or (inputs(94)));
    layer0_outputs(4806) <= (inputs(191)) or (inputs(244));
    layer0_outputs(4807) <= not(inputs(166));
    layer0_outputs(4808) <= not(inputs(100));
    layer0_outputs(4809) <= not((inputs(17)) or (inputs(148)));
    layer0_outputs(4810) <= not(inputs(130));
    layer0_outputs(4811) <= (inputs(237)) and not (inputs(201));
    layer0_outputs(4812) <= inputs(93);
    layer0_outputs(4813) <= not((inputs(19)) or (inputs(122)));
    layer0_outputs(4814) <= not(inputs(78)) or (inputs(66));
    layer0_outputs(4815) <= not((inputs(157)) and (inputs(78)));
    layer0_outputs(4816) <= not(inputs(186));
    layer0_outputs(4817) <= '1';
    layer0_outputs(4818) <= not(inputs(178));
    layer0_outputs(4819) <= (inputs(186)) or (inputs(156));
    layer0_outputs(4820) <= (inputs(55)) and not (inputs(137));
    layer0_outputs(4821) <= not(inputs(73)) or (inputs(87));
    layer0_outputs(4822) <= not(inputs(198)) or (inputs(17));
    layer0_outputs(4823) <= inputs(80);
    layer0_outputs(4824) <= not(inputs(181)) or (inputs(79));
    layer0_outputs(4825) <= (inputs(27)) or (inputs(159));
    layer0_outputs(4826) <= inputs(247);
    layer0_outputs(4827) <= not(inputs(83));
    layer0_outputs(4828) <= not(inputs(210));
    layer0_outputs(4829) <= not(inputs(75)) or (inputs(1));
    layer0_outputs(4830) <= not(inputs(146));
    layer0_outputs(4831) <= inputs(154);
    layer0_outputs(4832) <= not(inputs(195));
    layer0_outputs(4833) <= not(inputs(90));
    layer0_outputs(4834) <= inputs(212);
    layer0_outputs(4835) <= (inputs(129)) or (inputs(98));
    layer0_outputs(4836) <= not(inputs(21)) or (inputs(82));
    layer0_outputs(4837) <= not((inputs(78)) and (inputs(167)));
    layer0_outputs(4838) <= not(inputs(254));
    layer0_outputs(4839) <= not(inputs(24));
    layer0_outputs(4840) <= inputs(106);
    layer0_outputs(4841) <= inputs(247);
    layer0_outputs(4842) <= not(inputs(58));
    layer0_outputs(4843) <= not(inputs(108));
    layer0_outputs(4844) <= not(inputs(172)) or (inputs(32));
    layer0_outputs(4845) <= (inputs(1)) and (inputs(13));
    layer0_outputs(4846) <= not(inputs(184));
    layer0_outputs(4847) <= inputs(120);
    layer0_outputs(4848) <= (inputs(203)) or (inputs(21));
    layer0_outputs(4849) <= not(inputs(231)) or (inputs(83));
    layer0_outputs(4850) <= (inputs(184)) and not (inputs(91));
    layer0_outputs(4851) <= inputs(131);
    layer0_outputs(4852) <= inputs(192);
    layer0_outputs(4853) <= not(inputs(14));
    layer0_outputs(4854) <= inputs(103);
    layer0_outputs(4855) <= (inputs(42)) or (inputs(83));
    layer0_outputs(4856) <= not(inputs(149));
    layer0_outputs(4857) <= not((inputs(176)) or (inputs(186)));
    layer0_outputs(4858) <= not(inputs(170));
    layer0_outputs(4859) <= (inputs(116)) or (inputs(68));
    layer0_outputs(4860) <= (inputs(234)) or (inputs(16));
    layer0_outputs(4861) <= not((inputs(214)) or (inputs(176)));
    layer0_outputs(4862) <= inputs(68);
    layer0_outputs(4863) <= not(inputs(230));
    layer0_outputs(4864) <= not(inputs(239));
    layer0_outputs(4865) <= inputs(170);
    layer0_outputs(4866) <= not((inputs(226)) or (inputs(188)));
    layer0_outputs(4867) <= not(inputs(4)) or (inputs(109));
    layer0_outputs(4868) <= (inputs(87)) and not (inputs(126));
    layer0_outputs(4869) <= not(inputs(212));
    layer0_outputs(4870) <= not(inputs(44));
    layer0_outputs(4871) <= '0';
    layer0_outputs(4872) <= not((inputs(79)) or (inputs(227)));
    layer0_outputs(4873) <= not((inputs(189)) xor (inputs(19)));
    layer0_outputs(4874) <= inputs(163);
    layer0_outputs(4875) <= not(inputs(227));
    layer0_outputs(4876) <= not(inputs(244));
    layer0_outputs(4877) <= not(inputs(165));
    layer0_outputs(4878) <= not(inputs(67)) or (inputs(102));
    layer0_outputs(4879) <= not(inputs(61)) or (inputs(142));
    layer0_outputs(4880) <= (inputs(17)) and (inputs(17));
    layer0_outputs(4881) <= not((inputs(96)) xor (inputs(192)));
    layer0_outputs(4882) <= not(inputs(204)) or (inputs(253));
    layer0_outputs(4883) <= not((inputs(95)) xor (inputs(29)));
    layer0_outputs(4884) <= inputs(199);
    layer0_outputs(4885) <= (inputs(61)) and not (inputs(205));
    layer0_outputs(4886) <= inputs(114);
    layer0_outputs(4887) <= not(inputs(106));
    layer0_outputs(4888) <= inputs(136);
    layer0_outputs(4889) <= not((inputs(122)) or (inputs(114)));
    layer0_outputs(4890) <= (inputs(199)) and not (inputs(64));
    layer0_outputs(4891) <= not((inputs(11)) or (inputs(250)));
    layer0_outputs(4892) <= inputs(245);
    layer0_outputs(4893) <= not((inputs(91)) xor (inputs(126)));
    layer0_outputs(4894) <= (inputs(105)) and (inputs(166));
    layer0_outputs(4895) <= (inputs(160)) or (inputs(171));
    layer0_outputs(4896) <= not((inputs(222)) or (inputs(112)));
    layer0_outputs(4897) <= '1';
    layer0_outputs(4898) <= not(inputs(20));
    layer0_outputs(4899) <= not(inputs(110));
    layer0_outputs(4900) <= not((inputs(156)) xor (inputs(17)));
    layer0_outputs(4901) <= '1';
    layer0_outputs(4902) <= (inputs(95)) xor (inputs(32));
    layer0_outputs(4903) <= (inputs(196)) and not (inputs(86));
    layer0_outputs(4904) <= inputs(42);
    layer0_outputs(4905) <= not((inputs(110)) or (inputs(198)));
    layer0_outputs(4906) <= not((inputs(21)) or (inputs(238)));
    layer0_outputs(4907) <= not((inputs(204)) or (inputs(92)));
    layer0_outputs(4908) <= not(inputs(115)) or (inputs(19));
    layer0_outputs(4909) <= not(inputs(83)) or (inputs(112));
    layer0_outputs(4910) <= inputs(120);
    layer0_outputs(4911) <= (inputs(97)) or (inputs(67));
    layer0_outputs(4912) <= not(inputs(203));
    layer0_outputs(4913) <= not((inputs(145)) xor (inputs(129)));
    layer0_outputs(4914) <= (inputs(119)) and (inputs(40));
    layer0_outputs(4915) <= (inputs(154)) or (inputs(245));
    layer0_outputs(4916) <= (inputs(88)) and not (inputs(18));
    layer0_outputs(4917) <= '0';
    layer0_outputs(4918) <= '1';
    layer0_outputs(4919) <= not((inputs(202)) or (inputs(243)));
    layer0_outputs(4920) <= not((inputs(136)) xor (inputs(143)));
    layer0_outputs(4921) <= not(inputs(118));
    layer0_outputs(4922) <= inputs(103);
    layer0_outputs(4923) <= inputs(77);
    layer0_outputs(4924) <= (inputs(146)) or (inputs(107));
    layer0_outputs(4925) <= (inputs(69)) xor (inputs(190));
    layer0_outputs(4926) <= inputs(246);
    layer0_outputs(4927) <= not((inputs(92)) or (inputs(53)));
    layer0_outputs(4928) <= inputs(37);
    layer0_outputs(4929) <= not(inputs(225)) or (inputs(112));
    layer0_outputs(4930) <= (inputs(205)) or (inputs(172));
    layer0_outputs(4931) <= not(inputs(113));
    layer0_outputs(4932) <= inputs(59);
    layer0_outputs(4933) <= inputs(216);
    layer0_outputs(4934) <= not(inputs(138));
    layer0_outputs(4935) <= inputs(133);
    layer0_outputs(4936) <= (inputs(16)) xor (inputs(63));
    layer0_outputs(4937) <= not(inputs(144));
    layer0_outputs(4938) <= (inputs(53)) and not (inputs(31));
    layer0_outputs(4939) <= '0';
    layer0_outputs(4940) <= (inputs(155)) or (inputs(32));
    layer0_outputs(4941) <= not((inputs(180)) or (inputs(200)));
    layer0_outputs(4942) <= not((inputs(112)) or (inputs(217)));
    layer0_outputs(4943) <= (inputs(162)) or (inputs(70));
    layer0_outputs(4944) <= not(inputs(25));
    layer0_outputs(4945) <= not(inputs(89));
    layer0_outputs(4946) <= not(inputs(153)) or (inputs(8));
    layer0_outputs(4947) <= not((inputs(125)) or (inputs(74)));
    layer0_outputs(4948) <= not(inputs(146)) or (inputs(153));
    layer0_outputs(4949) <= (inputs(216)) and not (inputs(111));
    layer0_outputs(4950) <= (inputs(18)) or (inputs(17));
    layer0_outputs(4951) <= inputs(182);
    layer0_outputs(4952) <= (inputs(69)) and not (inputs(29));
    layer0_outputs(4953) <= not(inputs(198)) or (inputs(131));
    layer0_outputs(4954) <= not((inputs(34)) xor (inputs(160)));
    layer0_outputs(4955) <= inputs(234);
    layer0_outputs(4956) <= not((inputs(192)) or (inputs(104)));
    layer0_outputs(4957) <= not(inputs(188));
    layer0_outputs(4958) <= (inputs(51)) or (inputs(66));
    layer0_outputs(4959) <= (inputs(163)) and not (inputs(151));
    layer0_outputs(4960) <= not(inputs(46));
    layer0_outputs(4961) <= not(inputs(110));
    layer0_outputs(4962) <= inputs(116);
    layer0_outputs(4963) <= '0';
    layer0_outputs(4964) <= inputs(8);
    layer0_outputs(4965) <= (inputs(3)) xor (inputs(93));
    layer0_outputs(4966) <= (inputs(224)) or (inputs(113));
    layer0_outputs(4967) <= not(inputs(245));
    layer0_outputs(4968) <= not((inputs(113)) or (inputs(43)));
    layer0_outputs(4969) <= not((inputs(202)) or (inputs(158)));
    layer0_outputs(4970) <= not((inputs(43)) and (inputs(234)));
    layer0_outputs(4971) <= inputs(137);
    layer0_outputs(4972) <= (inputs(150)) and not (inputs(78));
    layer0_outputs(4973) <= inputs(28);
    layer0_outputs(4974) <= not(inputs(136)) or (inputs(163));
    layer0_outputs(4975) <= not(inputs(121)) or (inputs(88));
    layer0_outputs(4976) <= inputs(86);
    layer0_outputs(4977) <= inputs(68);
    layer0_outputs(4978) <= inputs(89);
    layer0_outputs(4979) <= (inputs(8)) and not (inputs(254));
    layer0_outputs(4980) <= not(inputs(199)) or (inputs(158));
    layer0_outputs(4981) <= inputs(112);
    layer0_outputs(4982) <= not(inputs(215));
    layer0_outputs(4983) <= (inputs(117)) and not (inputs(143));
    layer0_outputs(4984) <= '1';
    layer0_outputs(4985) <= not(inputs(88));
    layer0_outputs(4986) <= not(inputs(25));
    layer0_outputs(4987) <= inputs(68);
    layer0_outputs(4988) <= not(inputs(195));
    layer0_outputs(4989) <= not(inputs(67));
    layer0_outputs(4990) <= (inputs(181)) and (inputs(81));
    layer0_outputs(4991) <= (inputs(128)) or (inputs(124));
    layer0_outputs(4992) <= (inputs(70)) and not (inputs(5));
    layer0_outputs(4993) <= not(inputs(222));
    layer0_outputs(4994) <= not(inputs(9)) or (inputs(3));
    layer0_outputs(4995) <= (inputs(61)) and not (inputs(127));
    layer0_outputs(4996) <= not((inputs(94)) or (inputs(156)));
    layer0_outputs(4997) <= (inputs(213)) and not (inputs(73));
    layer0_outputs(4998) <= '1';
    layer0_outputs(4999) <= not((inputs(93)) or (inputs(107)));
    layer0_outputs(5000) <= not((inputs(99)) or (inputs(199)));
    layer0_outputs(5001) <= inputs(164);
    layer0_outputs(5002) <= not((inputs(151)) and (inputs(102)));
    layer0_outputs(5003) <= (inputs(248)) or (inputs(202));
    layer0_outputs(5004) <= inputs(180);
    layer0_outputs(5005) <= inputs(127);
    layer0_outputs(5006) <= '1';
    layer0_outputs(5007) <= not(inputs(97));
    layer0_outputs(5008) <= not(inputs(211));
    layer0_outputs(5009) <= (inputs(74)) xor (inputs(233));
    layer0_outputs(5010) <= (inputs(37)) xor (inputs(55));
    layer0_outputs(5011) <= inputs(21);
    layer0_outputs(5012) <= not(inputs(102));
    layer0_outputs(5013) <= not(inputs(41));
    layer0_outputs(5014) <= inputs(10);
    layer0_outputs(5015) <= (inputs(83)) or (inputs(197));
    layer0_outputs(5016) <= not((inputs(36)) or (inputs(44)));
    layer0_outputs(5017) <= (inputs(68)) or (inputs(115));
    layer0_outputs(5018) <= inputs(230);
    layer0_outputs(5019) <= not(inputs(230));
    layer0_outputs(5020) <= not(inputs(122));
    layer0_outputs(5021) <= not(inputs(80)) or (inputs(175));
    layer0_outputs(5022) <= '0';
    layer0_outputs(5023) <= not(inputs(127));
    layer0_outputs(5024) <= (inputs(138)) and not (inputs(20));
    layer0_outputs(5025) <= not((inputs(201)) or (inputs(33)));
    layer0_outputs(5026) <= inputs(90);
    layer0_outputs(5027) <= (inputs(105)) or (inputs(147));
    layer0_outputs(5028) <= inputs(58);
    layer0_outputs(5029) <= (inputs(56)) and not (inputs(205));
    layer0_outputs(5030) <= inputs(75);
    layer0_outputs(5031) <= not(inputs(213));
    layer0_outputs(5032) <= inputs(231);
    layer0_outputs(5033) <= (inputs(65)) or (inputs(178));
    layer0_outputs(5034) <= inputs(163);
    layer0_outputs(5035) <= not((inputs(244)) or (inputs(218)));
    layer0_outputs(5036) <= (inputs(54)) and not (inputs(127));
    layer0_outputs(5037) <= (inputs(118)) and not (inputs(94));
    layer0_outputs(5038) <= inputs(117);
    layer0_outputs(5039) <= inputs(117);
    layer0_outputs(5040) <= inputs(172);
    layer0_outputs(5041) <= (inputs(113)) xor (inputs(134));
    layer0_outputs(5042) <= not(inputs(229));
    layer0_outputs(5043) <= inputs(8);
    layer0_outputs(5044) <= inputs(177);
    layer0_outputs(5045) <= inputs(165);
    layer0_outputs(5046) <= (inputs(157)) or (inputs(226));
    layer0_outputs(5047) <= not(inputs(193));
    layer0_outputs(5048) <= (inputs(132)) or (inputs(132));
    layer0_outputs(5049) <= not(inputs(219));
    layer0_outputs(5050) <= inputs(65);
    layer0_outputs(5051) <= not(inputs(225));
    layer0_outputs(5052) <= not(inputs(248)) or (inputs(16));
    layer0_outputs(5053) <= not((inputs(253)) or (inputs(116)));
    layer0_outputs(5054) <= not((inputs(175)) or (inputs(6)));
    layer0_outputs(5055) <= not(inputs(203));
    layer0_outputs(5056) <= '1';
    layer0_outputs(5057) <= not(inputs(71)) or (inputs(108));
    layer0_outputs(5058) <= not(inputs(167)) or (inputs(188));
    layer0_outputs(5059) <= inputs(20);
    layer0_outputs(5060) <= (inputs(7)) and not (inputs(13));
    layer0_outputs(5061) <= (inputs(243)) or (inputs(207));
    layer0_outputs(5062) <= not(inputs(139)) or (inputs(231));
    layer0_outputs(5063) <= not(inputs(139)) or (inputs(65));
    layer0_outputs(5064) <= not(inputs(201));
    layer0_outputs(5065) <= not((inputs(239)) or (inputs(74)));
    layer0_outputs(5066) <= not((inputs(246)) xor (inputs(44)));
    layer0_outputs(5067) <= not((inputs(36)) or (inputs(19)));
    layer0_outputs(5068) <= not((inputs(138)) or (inputs(76)));
    layer0_outputs(5069) <= inputs(68);
    layer0_outputs(5070) <= not(inputs(41));
    layer0_outputs(5071) <= (inputs(74)) or (inputs(149));
    layer0_outputs(5072) <= not(inputs(233)) or (inputs(4));
    layer0_outputs(5073) <= not((inputs(250)) xor (inputs(1)));
    layer0_outputs(5074) <= (inputs(40)) and not (inputs(54));
    layer0_outputs(5075) <= (inputs(43)) and not (inputs(117));
    layer0_outputs(5076) <= not(inputs(57));
    layer0_outputs(5077) <= not((inputs(172)) xor (inputs(107)));
    layer0_outputs(5078) <= not(inputs(138));
    layer0_outputs(5079) <= not(inputs(99));
    layer0_outputs(5080) <= (inputs(234)) or (inputs(144));
    layer0_outputs(5081) <= (inputs(34)) or (inputs(49));
    layer0_outputs(5082) <= not((inputs(166)) xor (inputs(213)));
    layer0_outputs(5083) <= not(inputs(8));
    layer0_outputs(5084) <= (inputs(235)) or (inputs(150));
    layer0_outputs(5085) <= inputs(3);
    layer0_outputs(5086) <= (inputs(143)) and not (inputs(40));
    layer0_outputs(5087) <= inputs(89);
    layer0_outputs(5088) <= not((inputs(160)) or (inputs(246)));
    layer0_outputs(5089) <= not(inputs(133)) or (inputs(196));
    layer0_outputs(5090) <= (inputs(82)) and not (inputs(182));
    layer0_outputs(5091) <= not(inputs(130)) or (inputs(19));
    layer0_outputs(5092) <= (inputs(252)) and not (inputs(138));
    layer0_outputs(5093) <= not(inputs(202)) or (inputs(4));
    layer0_outputs(5094) <= not(inputs(87)) or (inputs(95));
    layer0_outputs(5095) <= not((inputs(172)) or (inputs(170)));
    layer0_outputs(5096) <= not(inputs(126));
    layer0_outputs(5097) <= not(inputs(102));
    layer0_outputs(5098) <= (inputs(156)) xor (inputs(205));
    layer0_outputs(5099) <= (inputs(171)) or (inputs(63));
    layer0_outputs(5100) <= not((inputs(147)) or (inputs(127)));
    layer0_outputs(5101) <= (inputs(96)) and not (inputs(198));
    layer0_outputs(5102) <= (inputs(223)) or (inputs(101));
    layer0_outputs(5103) <= inputs(76);
    layer0_outputs(5104) <= inputs(210);
    layer0_outputs(5105) <= not(inputs(129));
    layer0_outputs(5106) <= (inputs(22)) and not (inputs(114));
    layer0_outputs(5107) <= inputs(37);
    layer0_outputs(5108) <= inputs(214);
    layer0_outputs(5109) <= not((inputs(242)) or (inputs(239)));
    layer0_outputs(5110) <= not((inputs(255)) xor (inputs(98)));
    layer0_outputs(5111) <= (inputs(254)) or (inputs(101));
    layer0_outputs(5112) <= (inputs(183)) xor (inputs(229));
    layer0_outputs(5113) <= (inputs(32)) and not (inputs(12));
    layer0_outputs(5114) <= (inputs(36)) xor (inputs(54));
    layer0_outputs(5115) <= (inputs(86)) or (inputs(184));
    layer0_outputs(5116) <= not(inputs(209));
    layer0_outputs(5117) <= inputs(151);
    layer0_outputs(5118) <= inputs(100);
    layer0_outputs(5119) <= (inputs(52)) or (inputs(172));
    outputs(0) <= not((layer0_outputs(2813)) xor (layer0_outputs(4579)));
    outputs(1) <= layer0_outputs(3785);
    outputs(2) <= not(layer0_outputs(1470));
    outputs(3) <= not(layer0_outputs(1195));
    outputs(4) <= (layer0_outputs(3994)) or (layer0_outputs(2935));
    outputs(5) <= layer0_outputs(342);
    outputs(6) <= not(layer0_outputs(3404)) or (layer0_outputs(724));
    outputs(7) <= not(layer0_outputs(4847));
    outputs(8) <= (layer0_outputs(3371)) xor (layer0_outputs(1925));
    outputs(9) <= not(layer0_outputs(2809));
    outputs(10) <= not(layer0_outputs(4988));
    outputs(11) <= not(layer0_outputs(1964));
    outputs(12) <= not(layer0_outputs(2014));
    outputs(13) <= layer0_outputs(1643);
    outputs(14) <= not(layer0_outputs(2714));
    outputs(15) <= not(layer0_outputs(3557));
    outputs(16) <= layer0_outputs(543);
    outputs(17) <= layer0_outputs(4233);
    outputs(18) <= not(layer0_outputs(4602));
    outputs(19) <= not((layer0_outputs(1814)) xor (layer0_outputs(1160)));
    outputs(20) <= layer0_outputs(1270);
    outputs(21) <= layer0_outputs(586);
    outputs(22) <= not(layer0_outputs(3401));
    outputs(23) <= layer0_outputs(4906);
    outputs(24) <= layer0_outputs(3522);
    outputs(25) <= layer0_outputs(3380);
    outputs(26) <= not((layer0_outputs(4048)) and (layer0_outputs(4469)));
    outputs(27) <= (layer0_outputs(2873)) or (layer0_outputs(4959));
    outputs(28) <= (layer0_outputs(922)) or (layer0_outputs(3514));
    outputs(29) <= (layer0_outputs(3223)) and not (layer0_outputs(4524));
    outputs(30) <= layer0_outputs(2697);
    outputs(31) <= not(layer0_outputs(4339));
    outputs(32) <= layer0_outputs(1154);
    outputs(33) <= not((layer0_outputs(3388)) and (layer0_outputs(4576)));
    outputs(34) <= not((layer0_outputs(1537)) or (layer0_outputs(4863)));
    outputs(35) <= not((layer0_outputs(4068)) and (layer0_outputs(1390)));
    outputs(36) <= not((layer0_outputs(2997)) and (layer0_outputs(968)));
    outputs(37) <= not(layer0_outputs(4107));
    outputs(38) <= layer0_outputs(4446);
    outputs(39) <= (layer0_outputs(656)) xor (layer0_outputs(3898));
    outputs(40) <= (layer0_outputs(3608)) xor (layer0_outputs(3598));
    outputs(41) <= (layer0_outputs(244)) and not (layer0_outputs(1847));
    outputs(42) <= layer0_outputs(4743);
    outputs(43) <= not(layer0_outputs(816));
    outputs(44) <= not(layer0_outputs(248));
    outputs(45) <= (layer0_outputs(1404)) and not (layer0_outputs(3159));
    outputs(46) <= (layer0_outputs(2169)) or (layer0_outputs(4663));
    outputs(47) <= layer0_outputs(2044);
    outputs(48) <= layer0_outputs(760);
    outputs(49) <= (layer0_outputs(623)) and not (layer0_outputs(895));
    outputs(50) <= not(layer0_outputs(27));
    outputs(51) <= layer0_outputs(2136);
    outputs(52) <= layer0_outputs(1269);
    outputs(53) <= not(layer0_outputs(1474));
    outputs(54) <= not(layer0_outputs(4561));
    outputs(55) <= not(layer0_outputs(1521));
    outputs(56) <= not(layer0_outputs(1567));
    outputs(57) <= (layer0_outputs(2277)) and (layer0_outputs(302));
    outputs(58) <= layer0_outputs(1166);
    outputs(59) <= not(layer0_outputs(2970));
    outputs(60) <= not(layer0_outputs(2644));
    outputs(61) <= not(layer0_outputs(4971));
    outputs(62) <= layer0_outputs(3631);
    outputs(63) <= not((layer0_outputs(3780)) xor (layer0_outputs(1632)));
    outputs(64) <= layer0_outputs(3075);
    outputs(65) <= (layer0_outputs(476)) xor (layer0_outputs(2678));
    outputs(66) <= not(layer0_outputs(2098));
    outputs(67) <= layer0_outputs(709);
    outputs(68) <= not((layer0_outputs(3382)) xor (layer0_outputs(2199)));
    outputs(69) <= layer0_outputs(2161);
    outputs(70) <= not((layer0_outputs(3024)) xor (layer0_outputs(4605)));
    outputs(71) <= (layer0_outputs(1336)) and not (layer0_outputs(1825));
    outputs(72) <= layer0_outputs(2858);
    outputs(73) <= (layer0_outputs(16)) xor (layer0_outputs(2286));
    outputs(74) <= not(layer0_outputs(404));
    outputs(75) <= (layer0_outputs(4681)) and (layer0_outputs(2971));
    outputs(76) <= (layer0_outputs(1500)) and not (layer0_outputs(1125));
    outputs(77) <= not(layer0_outputs(1318));
    outputs(78) <= not((layer0_outputs(1822)) and (layer0_outputs(966)));
    outputs(79) <= (layer0_outputs(4328)) xor (layer0_outputs(1059));
    outputs(80) <= not(layer0_outputs(4899));
    outputs(81) <= layer0_outputs(491);
    outputs(82) <= not(layer0_outputs(1582));
    outputs(83) <= (layer0_outputs(3451)) and not (layer0_outputs(950));
    outputs(84) <= layer0_outputs(4966);
    outputs(85) <= (layer0_outputs(3666)) xor (layer0_outputs(3793));
    outputs(86) <= (layer0_outputs(1396)) xor (layer0_outputs(2981));
    outputs(87) <= layer0_outputs(700);
    outputs(88) <= not((layer0_outputs(1511)) xor (layer0_outputs(4480)));
    outputs(89) <= layer0_outputs(4708);
    outputs(90) <= layer0_outputs(3679);
    outputs(91) <= (layer0_outputs(3451)) and not (layer0_outputs(3210));
    outputs(92) <= (layer0_outputs(3461)) or (layer0_outputs(4603));
    outputs(93) <= layer0_outputs(2875);
    outputs(94) <= not(layer0_outputs(4922)) or (layer0_outputs(5044));
    outputs(95) <= layer0_outputs(4512);
    outputs(96) <= (layer0_outputs(4025)) and not (layer0_outputs(447));
    outputs(97) <= not(layer0_outputs(3968));
    outputs(98) <= not((layer0_outputs(1834)) and (layer0_outputs(3856)));
    outputs(99) <= not(layer0_outputs(2737));
    outputs(100) <= not(layer0_outputs(2518));
    outputs(101) <= not(layer0_outputs(736)) or (layer0_outputs(4063));
    outputs(102) <= layer0_outputs(2798);
    outputs(103) <= not((layer0_outputs(861)) xor (layer0_outputs(3753)));
    outputs(104) <= layer0_outputs(4405);
    outputs(105) <= layer0_outputs(2143);
    outputs(106) <= not(layer0_outputs(2321));
    outputs(107) <= layer0_outputs(798);
    outputs(108) <= not(layer0_outputs(5117));
    outputs(109) <= not(layer0_outputs(1076));
    outputs(110) <= layer0_outputs(3498);
    outputs(111) <= not(layer0_outputs(4779)) or (layer0_outputs(2265));
    outputs(112) <= not(layer0_outputs(4441));
    outputs(113) <= not(layer0_outputs(4241));
    outputs(114) <= not((layer0_outputs(4198)) xor (layer0_outputs(3694)));
    outputs(115) <= not(layer0_outputs(3662));
    outputs(116) <= (layer0_outputs(4864)) and not (layer0_outputs(448));
    outputs(117) <= layer0_outputs(298);
    outputs(118) <= not(layer0_outputs(4805));
    outputs(119) <= layer0_outputs(1808);
    outputs(120) <= not((layer0_outputs(3366)) or (layer0_outputs(1167)));
    outputs(121) <= (layer0_outputs(2384)) and not (layer0_outputs(2940));
    outputs(122) <= layer0_outputs(437);
    outputs(123) <= layer0_outputs(2753);
    outputs(124) <= not((layer0_outputs(2133)) xor (layer0_outputs(358)));
    outputs(125) <= (layer0_outputs(2370)) or (layer0_outputs(4190));
    outputs(126) <= layer0_outputs(4052);
    outputs(127) <= not(layer0_outputs(879));
    outputs(128) <= not((layer0_outputs(3897)) or (layer0_outputs(868)));
    outputs(129) <= not(layer0_outputs(3884));
    outputs(130) <= layer0_outputs(739);
    outputs(131) <= layer0_outputs(784);
    outputs(132) <= not((layer0_outputs(113)) and (layer0_outputs(285)));
    outputs(133) <= (layer0_outputs(561)) xor (layer0_outputs(3796));
    outputs(134) <= not(layer0_outputs(4539));
    outputs(135) <= (layer0_outputs(530)) or (layer0_outputs(4652));
    outputs(136) <= layer0_outputs(550);
    outputs(137) <= not(layer0_outputs(1534));
    outputs(138) <= (layer0_outputs(4059)) and not (layer0_outputs(1285));
    outputs(139) <= (layer0_outputs(2855)) or (layer0_outputs(3676));
    outputs(140) <= not(layer0_outputs(1412));
    outputs(141) <= (layer0_outputs(3337)) and (layer0_outputs(3034));
    outputs(142) <= (layer0_outputs(669)) and not (layer0_outputs(1805));
    outputs(143) <= (layer0_outputs(4987)) or (layer0_outputs(3038));
    outputs(144) <= (layer0_outputs(5052)) xor (layer0_outputs(4642));
    outputs(145) <= not((layer0_outputs(2650)) xor (layer0_outputs(3873)));
    outputs(146) <= not((layer0_outputs(2222)) or (layer0_outputs(820)));
    outputs(147) <= not(layer0_outputs(4739));
    outputs(148) <= not(layer0_outputs(5088));
    outputs(149) <= not(layer0_outputs(1866));
    outputs(150) <= (layer0_outputs(297)) xor (layer0_outputs(1122));
    outputs(151) <= not((layer0_outputs(3834)) and (layer0_outputs(407)));
    outputs(152) <= (layer0_outputs(4179)) and not (layer0_outputs(4160));
    outputs(153) <= not(layer0_outputs(5037));
    outputs(154) <= not(layer0_outputs(4388));
    outputs(155) <= layer0_outputs(3078);
    outputs(156) <= (layer0_outputs(1594)) and (layer0_outputs(4506));
    outputs(157) <= (layer0_outputs(487)) xor (layer0_outputs(1180));
    outputs(158) <= not((layer0_outputs(281)) xor (layer0_outputs(271)));
    outputs(159) <= not(layer0_outputs(4409));
    outputs(160) <= layer0_outputs(2076);
    outputs(161) <= not(layer0_outputs(1771));
    outputs(162) <= layer0_outputs(4470);
    outputs(163) <= layer0_outputs(4199);
    outputs(164) <= not(layer0_outputs(2364)) or (layer0_outputs(732));
    outputs(165) <= not(layer0_outputs(2477));
    outputs(166) <= not((layer0_outputs(4857)) or (layer0_outputs(1091)));
    outputs(167) <= not((layer0_outputs(3707)) and (layer0_outputs(4619)));
    outputs(168) <= (layer0_outputs(596)) and (layer0_outputs(3922));
    outputs(169) <= not((layer0_outputs(455)) and (layer0_outputs(944)));
    outputs(170) <= (layer0_outputs(4141)) or (layer0_outputs(2730));
    outputs(171) <= (layer0_outputs(1703)) and not (layer0_outputs(384));
    outputs(172) <= not(layer0_outputs(4171));
    outputs(173) <= not(layer0_outputs(345));
    outputs(174) <= not((layer0_outputs(4392)) xor (layer0_outputs(2154)));
    outputs(175) <= (layer0_outputs(2210)) and (layer0_outputs(1143));
    outputs(176) <= layer0_outputs(5020);
    outputs(177) <= not(layer0_outputs(3750));
    outputs(178) <= not(layer0_outputs(2569)) or (layer0_outputs(647));
    outputs(179) <= layer0_outputs(2976);
    outputs(180) <= not(layer0_outputs(359));
    outputs(181) <= (layer0_outputs(2620)) and (layer0_outputs(2931));
    outputs(182) <= not((layer0_outputs(3512)) and (layer0_outputs(3095)));
    outputs(183) <= layer0_outputs(3931);
    outputs(184) <= (layer0_outputs(72)) and not (layer0_outputs(4487));
    outputs(185) <= (layer0_outputs(796)) or (layer0_outputs(717));
    outputs(186) <= layer0_outputs(4849);
    outputs(187) <= (layer0_outputs(3608)) and not (layer0_outputs(3659));
    outputs(188) <= (layer0_outputs(3252)) and not (layer0_outputs(2329));
    outputs(189) <= not(layer0_outputs(2886));
    outputs(190) <= not(layer0_outputs(379));
    outputs(191) <= not(layer0_outputs(2894));
    outputs(192) <= (layer0_outputs(1686)) xor (layer0_outputs(3673));
    outputs(193) <= not(layer0_outputs(4900));
    outputs(194) <= not(layer0_outputs(3497));
    outputs(195) <= layer0_outputs(30);
    outputs(196) <= (layer0_outputs(4895)) and not (layer0_outputs(3508));
    outputs(197) <= not(layer0_outputs(872));
    outputs(198) <= not(layer0_outputs(3879)) or (layer0_outputs(3738));
    outputs(199) <= (layer0_outputs(3981)) and not (layer0_outputs(1509));
    outputs(200) <= not(layer0_outputs(3549));
    outputs(201) <= layer0_outputs(790);
    outputs(202) <= not(layer0_outputs(2626));
    outputs(203) <= layer0_outputs(3308);
    outputs(204) <= not(layer0_outputs(166));
    outputs(205) <= not((layer0_outputs(3224)) and (layer0_outputs(3777)));
    outputs(206) <= (layer0_outputs(3465)) or (layer0_outputs(1415));
    outputs(207) <= (layer0_outputs(1764)) xor (layer0_outputs(3542));
    outputs(208) <= layer0_outputs(520);
    outputs(209) <= (layer0_outputs(1299)) and not (layer0_outputs(3902));
    outputs(210) <= (layer0_outputs(745)) xor (layer0_outputs(4394));
    outputs(211) <= not(layer0_outputs(3232));
    outputs(212) <= not(layer0_outputs(1391));
    outputs(213) <= (layer0_outputs(2287)) and not (layer0_outputs(1305));
    outputs(214) <= (layer0_outputs(588)) and not (layer0_outputs(4175));
    outputs(215) <= (layer0_outputs(2426)) and not (layer0_outputs(3366));
    outputs(216) <= not(layer0_outputs(2153));
    outputs(217) <= not(layer0_outputs(995));
    outputs(218) <= not(layer0_outputs(693));
    outputs(219) <= not(layer0_outputs(3104));
    outputs(220) <= layer0_outputs(2486);
    outputs(221) <= (layer0_outputs(2919)) and not (layer0_outputs(1779));
    outputs(222) <= not((layer0_outputs(1320)) and (layer0_outputs(95)));
    outputs(223) <= not(layer0_outputs(116));
    outputs(224) <= not(layer0_outputs(415));
    outputs(225) <= (layer0_outputs(1542)) and not (layer0_outputs(539));
    outputs(226) <= layer0_outputs(2462);
    outputs(227) <= not((layer0_outputs(1918)) and (layer0_outputs(4694)));
    outputs(228) <= (layer0_outputs(2926)) and not (layer0_outputs(2186));
    outputs(229) <= layer0_outputs(115);
    outputs(230) <= not(layer0_outputs(4604));
    outputs(231) <= not(layer0_outputs(995));
    outputs(232) <= (layer0_outputs(1304)) xor (layer0_outputs(1467));
    outputs(233) <= (layer0_outputs(1518)) and not (layer0_outputs(3936));
    outputs(234) <= not((layer0_outputs(3336)) xor (layer0_outputs(1047)));
    outputs(235) <= (layer0_outputs(2301)) or (layer0_outputs(3711));
    outputs(236) <= (layer0_outputs(907)) xor (layer0_outputs(1589));
    outputs(237) <= not(layer0_outputs(4540));
    outputs(238) <= not((layer0_outputs(3496)) and (layer0_outputs(4070)));
    outputs(239) <= layer0_outputs(2880);
    outputs(240) <= not(layer0_outputs(1799));
    outputs(241) <= not(layer0_outputs(2422));
    outputs(242) <= (layer0_outputs(1641)) or (layer0_outputs(1245));
    outputs(243) <= not(layer0_outputs(3009));
    outputs(244) <= not(layer0_outputs(283)) or (layer0_outputs(3721));
    outputs(245) <= not(layer0_outputs(1230));
    outputs(246) <= layer0_outputs(4991);
    outputs(247) <= layer0_outputs(4727);
    outputs(248) <= layer0_outputs(979);
    outputs(249) <= layer0_outputs(1155);
    outputs(250) <= layer0_outputs(4296);
    outputs(251) <= not((layer0_outputs(4369)) or (layer0_outputs(4410)));
    outputs(252) <= layer0_outputs(2844);
    outputs(253) <= layer0_outputs(587);
    outputs(254) <= (layer0_outputs(2421)) xor (layer0_outputs(2196));
    outputs(255) <= (layer0_outputs(2616)) or (layer0_outputs(1488));
    outputs(256) <= layer0_outputs(217);
    outputs(257) <= not(layer0_outputs(626));
    outputs(258) <= not(layer0_outputs(1460));
    outputs(259) <= not((layer0_outputs(2996)) xor (layer0_outputs(4824)));
    outputs(260) <= not(layer0_outputs(1461));
    outputs(261) <= layer0_outputs(1731);
    outputs(262) <= not(layer0_outputs(4359));
    outputs(263) <= not((layer0_outputs(4458)) xor (layer0_outputs(1348)));
    outputs(264) <= not(layer0_outputs(2482));
    outputs(265) <= not(layer0_outputs(2951));
    outputs(266) <= (layer0_outputs(4036)) and not (layer0_outputs(4723));
    outputs(267) <= not(layer0_outputs(2053));
    outputs(268) <= layer0_outputs(3194);
    outputs(269) <= layer0_outputs(3989);
    outputs(270) <= layer0_outputs(3980);
    outputs(271) <= not((layer0_outputs(402)) or (layer0_outputs(2117)));
    outputs(272) <= layer0_outputs(1981);
    outputs(273) <= not(layer0_outputs(4910));
    outputs(274) <= not(layer0_outputs(4211)) or (layer0_outputs(484));
    outputs(275) <= layer0_outputs(619);
    outputs(276) <= not(layer0_outputs(1577));
    outputs(277) <= layer0_outputs(2012);
    outputs(278) <= (layer0_outputs(550)) and (layer0_outputs(4546));
    outputs(279) <= (layer0_outputs(2700)) and not (layer0_outputs(2621));
    outputs(280) <= not(layer0_outputs(1254));
    outputs(281) <= (layer0_outputs(3414)) and not (layer0_outputs(2524));
    outputs(282) <= not((layer0_outputs(4697)) xor (layer0_outputs(2455)));
    outputs(283) <= not((layer0_outputs(5119)) xor (layer0_outputs(1508)));
    outputs(284) <= (layer0_outputs(3361)) xor (layer0_outputs(3487));
    outputs(285) <= not(layer0_outputs(3048));
    outputs(286) <= not(layer0_outputs(868));
    outputs(287) <= not((layer0_outputs(1829)) or (layer0_outputs(3159)));
    outputs(288) <= layer0_outputs(3925);
    outputs(289) <= (layer0_outputs(1176)) and not (layer0_outputs(2166));
    outputs(290) <= layer0_outputs(477);
    outputs(291) <= not(layer0_outputs(1917));
    outputs(292) <= layer0_outputs(1669);
    outputs(293) <= layer0_outputs(1928);
    outputs(294) <= not(layer0_outputs(4844)) or (layer0_outputs(3227));
    outputs(295) <= layer0_outputs(3526);
    outputs(296) <= not(layer0_outputs(4948));
    outputs(297) <= layer0_outputs(4521);
    outputs(298) <= not((layer0_outputs(1587)) and (layer0_outputs(4194)));
    outputs(299) <= not(layer0_outputs(817)) or (layer0_outputs(4820));
    outputs(300) <= not(layer0_outputs(51)) or (layer0_outputs(303));
    outputs(301) <= not(layer0_outputs(4868));
    outputs(302) <= (layer0_outputs(4008)) xor (layer0_outputs(432));
    outputs(303) <= layer0_outputs(3722);
    outputs(304) <= not(layer0_outputs(4497));
    outputs(305) <= not((layer0_outputs(1829)) and (layer0_outputs(535)));
    outputs(306) <= not(layer0_outputs(1233));
    outputs(307) <= not((layer0_outputs(2507)) and (layer0_outputs(4713)));
    outputs(308) <= not((layer0_outputs(1349)) or (layer0_outputs(4375)));
    outputs(309) <= (layer0_outputs(1581)) xor (layer0_outputs(2981));
    outputs(310) <= not(layer0_outputs(774));
    outputs(311) <= layer0_outputs(1175);
    outputs(312) <= (layer0_outputs(2073)) and (layer0_outputs(332));
    outputs(313) <= layer0_outputs(4813);
    outputs(314) <= not(layer0_outputs(2562));
    outputs(315) <= layer0_outputs(3452);
    outputs(316) <= layer0_outputs(1220);
    outputs(317) <= layer0_outputs(4934);
    outputs(318) <= not(layer0_outputs(2605));
    outputs(319) <= (layer0_outputs(3235)) and not (layer0_outputs(2032));
    outputs(320) <= (layer0_outputs(3601)) and (layer0_outputs(1186));
    outputs(321) <= layer0_outputs(1175);
    outputs(322) <= not(layer0_outputs(1783));
    outputs(323) <= not(layer0_outputs(3677)) or (layer0_outputs(2755));
    outputs(324) <= not(layer0_outputs(2884)) or (layer0_outputs(4806));
    outputs(325) <= not(layer0_outputs(1229)) or (layer0_outputs(2917));
    outputs(326) <= not((layer0_outputs(3545)) xor (layer0_outputs(4475)));
    outputs(327) <= not(layer0_outputs(3466));
    outputs(328) <= layer0_outputs(784);
    outputs(329) <= layer0_outputs(3816);
    outputs(330) <= layer0_outputs(4660);
    outputs(331) <= layer0_outputs(4066);
    outputs(332) <= not((layer0_outputs(3536)) xor (layer0_outputs(1612)));
    outputs(333) <= (layer0_outputs(3706)) and not (layer0_outputs(2135));
    outputs(334) <= layer0_outputs(2769);
    outputs(335) <= not(layer0_outputs(5093));
    outputs(336) <= (layer0_outputs(3427)) and not (layer0_outputs(2050));
    outputs(337) <= (layer0_outputs(311)) or (layer0_outputs(4583));
    outputs(338) <= not(layer0_outputs(1101)) or (layer0_outputs(2057));
    outputs(339) <= (layer0_outputs(2394)) or (layer0_outputs(4380));
    outputs(340) <= not(layer0_outputs(1127));
    outputs(341) <= layer0_outputs(4801);
    outputs(342) <= not((layer0_outputs(4760)) or (layer0_outputs(3335)));
    outputs(343) <= not(layer0_outputs(173));
    outputs(344) <= (layer0_outputs(3513)) xor (layer0_outputs(958));
    outputs(345) <= layer0_outputs(2862);
    outputs(346) <= not(layer0_outputs(2824));
    outputs(347) <= not(layer0_outputs(3579));
    outputs(348) <= (layer0_outputs(1083)) xor (layer0_outputs(4561));
    outputs(349) <= layer0_outputs(1077);
    outputs(350) <= not(layer0_outputs(4816)) or (layer0_outputs(484));
    outputs(351) <= not(layer0_outputs(2279));
    outputs(352) <= not(layer0_outputs(1428));
    outputs(353) <= layer0_outputs(3425);
    outputs(354) <= (layer0_outputs(1415)) or (layer0_outputs(1173));
    outputs(355) <= layer0_outputs(1263);
    outputs(356) <= layer0_outputs(1173);
    outputs(357) <= (layer0_outputs(3285)) and (layer0_outputs(1066));
    outputs(358) <= not(layer0_outputs(3620));
    outputs(359) <= not((layer0_outputs(3471)) xor (layer0_outputs(1289)));
    outputs(360) <= layer0_outputs(4709);
    outputs(361) <= layer0_outputs(2332);
    outputs(362) <= not(layer0_outputs(1272));
    outputs(363) <= not(layer0_outputs(2498));
    outputs(364) <= (layer0_outputs(3)) and not (layer0_outputs(4447));
    outputs(365) <= not(layer0_outputs(1832));
    outputs(366) <= (layer0_outputs(2736)) and not (layer0_outputs(1996));
    outputs(367) <= not(layer0_outputs(3563));
    outputs(368) <= layer0_outputs(3039);
    outputs(369) <= not(layer0_outputs(3280)) or (layer0_outputs(292));
    outputs(370) <= not(layer0_outputs(2746)) or (layer0_outputs(2453));
    outputs(371) <= not(layer0_outputs(612));
    outputs(372) <= (layer0_outputs(1578)) and (layer0_outputs(3178));
    outputs(373) <= (layer0_outputs(981)) and not (layer0_outputs(582));
    outputs(374) <= not(layer0_outputs(4327));
    outputs(375) <= not(layer0_outputs(1167)) or (layer0_outputs(2213));
    outputs(376) <= not(layer0_outputs(2681));
    outputs(377) <= not(layer0_outputs(4544));
    outputs(378) <= (layer0_outputs(83)) xor (layer0_outputs(475));
    outputs(379) <= (layer0_outputs(3244)) or (layer0_outputs(1450));
    outputs(380) <= not(layer0_outputs(3043));
    outputs(381) <= (layer0_outputs(343)) or (layer0_outputs(4846));
    outputs(382) <= not(layer0_outputs(4500));
    outputs(383) <= (layer0_outputs(1641)) and not (layer0_outputs(2172));
    outputs(384) <= layer0_outputs(115);
    outputs(385) <= layer0_outputs(2042);
    outputs(386) <= not(layer0_outputs(3855));
    outputs(387) <= not(layer0_outputs(2493)) or (layer0_outputs(2583));
    outputs(388) <= layer0_outputs(3741);
    outputs(389) <= (layer0_outputs(1260)) and not (layer0_outputs(154));
    outputs(390) <= not(layer0_outputs(4961));
    outputs(391) <= (layer0_outputs(2387)) and not (layer0_outputs(3869));
    outputs(392) <= layer0_outputs(2142);
    outputs(393) <= not(layer0_outputs(98));
    outputs(394) <= layer0_outputs(1816);
    outputs(395) <= (layer0_outputs(5086)) or (layer0_outputs(3387));
    outputs(396) <= layer0_outputs(1333);
    outputs(397) <= (layer0_outputs(2632)) or (layer0_outputs(2367));
    outputs(398) <= not((layer0_outputs(730)) and (layer0_outputs(3550)));
    outputs(399) <= not((layer0_outputs(4276)) and (layer0_outputs(3671)));
    outputs(400) <= layer0_outputs(1519);
    outputs(401) <= (layer0_outputs(1998)) and (layer0_outputs(4082));
    outputs(402) <= layer0_outputs(2528);
    outputs(403) <= not(layer0_outputs(1846)) or (layer0_outputs(1029));
    outputs(404) <= not(layer0_outputs(4335)) or (layer0_outputs(2890));
    outputs(405) <= (layer0_outputs(1688)) or (layer0_outputs(2100));
    outputs(406) <= (layer0_outputs(1185)) and not (layer0_outputs(371));
    outputs(407) <= layer0_outputs(2295);
    outputs(408) <= not(layer0_outputs(2050));
    outputs(409) <= not(layer0_outputs(3562));
    outputs(410) <= layer0_outputs(3663);
    outputs(411) <= not(layer0_outputs(3153));
    outputs(412) <= not(layer0_outputs(3015)) or (layer0_outputs(234));
    outputs(413) <= not(layer0_outputs(321));
    outputs(414) <= (layer0_outputs(3286)) or (layer0_outputs(4747));
    outputs(415) <= layer0_outputs(4552);
    outputs(416) <= layer0_outputs(596);
    outputs(417) <= (layer0_outputs(2586)) xor (layer0_outputs(660));
    outputs(418) <= not((layer0_outputs(2123)) and (layer0_outputs(890)));
    outputs(419) <= not(layer0_outputs(3540));
    outputs(420) <= not(layer0_outputs(29));
    outputs(421) <= (layer0_outputs(315)) and (layer0_outputs(674));
    outputs(422) <= layer0_outputs(2396);
    outputs(423) <= not((layer0_outputs(4785)) or (layer0_outputs(4013)));
    outputs(424) <= not(layer0_outputs(3802));
    outputs(425) <= not(layer0_outputs(1130));
    outputs(426) <= not(layer0_outputs(2679));
    outputs(427) <= not(layer0_outputs(1847));
    outputs(428) <= not(layer0_outputs(129));
    outputs(429) <= not(layer0_outputs(3014));
    outputs(430) <= layer0_outputs(383);
    outputs(431) <= layer0_outputs(3463);
    outputs(432) <= layer0_outputs(31);
    outputs(433) <= (layer0_outputs(1328)) xor (layer0_outputs(4025));
    outputs(434) <= not(layer0_outputs(3349)) or (layer0_outputs(460));
    outputs(435) <= not((layer0_outputs(4632)) xor (layer0_outputs(2656)));
    outputs(436) <= not((layer0_outputs(2468)) xor (layer0_outputs(4395)));
    outputs(437) <= not(layer0_outputs(3501));
    outputs(438) <= layer0_outputs(3327);
    outputs(439) <= (layer0_outputs(743)) or (layer0_outputs(1443));
    outputs(440) <= not(layer0_outputs(2338));
    outputs(441) <= (layer0_outputs(1860)) and not (layer0_outputs(3830));
    outputs(442) <= not(layer0_outputs(720));
    outputs(443) <= layer0_outputs(519);
    outputs(444) <= not((layer0_outputs(3290)) xor (layer0_outputs(989)));
    outputs(445) <= (layer0_outputs(4791)) and (layer0_outputs(302));
    outputs(446) <= layer0_outputs(4812);
    outputs(447) <= not(layer0_outputs(531));
    outputs(448) <= not(layer0_outputs(372));
    outputs(449) <= layer0_outputs(1165);
    outputs(450) <= layer0_outputs(978);
    outputs(451) <= layer0_outputs(3903);
    outputs(452) <= not(layer0_outputs(2232));
    outputs(453) <= (layer0_outputs(5038)) xor (layer0_outputs(4541));
    outputs(454) <= not(layer0_outputs(2952)) or (layer0_outputs(3328));
    outputs(455) <= (layer0_outputs(3919)) and (layer0_outputs(4630));
    outputs(456) <= not((layer0_outputs(3079)) xor (layer0_outputs(4601)));
    outputs(457) <= not(layer0_outputs(1984));
    outputs(458) <= layer0_outputs(715);
    outputs(459) <= layer0_outputs(3338);
    outputs(460) <= layer0_outputs(3416);
    outputs(461) <= (layer0_outputs(2241)) and (layer0_outputs(2723));
    outputs(462) <= not(layer0_outputs(4165));
    outputs(463) <= layer0_outputs(1208);
    outputs(464) <= not(layer0_outputs(243)) or (layer0_outputs(5034));
    outputs(465) <= not((layer0_outputs(4576)) and (layer0_outputs(4207)));
    outputs(466) <= layer0_outputs(4758);
    outputs(467) <= layer0_outputs(4645);
    outputs(468) <= not(layer0_outputs(2595));
    outputs(469) <= not(layer0_outputs(1332)) or (layer0_outputs(1274));
    outputs(470) <= layer0_outputs(836);
    outputs(471) <= layer0_outputs(236);
    outputs(472) <= (layer0_outputs(4428)) and (layer0_outputs(2104));
    outputs(473) <= layer0_outputs(1310);
    outputs(474) <= layer0_outputs(3355);
    outputs(475) <= (layer0_outputs(2099)) and (layer0_outputs(2693));
    outputs(476) <= layer0_outputs(186);
    outputs(477) <= not((layer0_outputs(350)) and (layer0_outputs(3704)));
    outputs(478) <= not(layer0_outputs(4302));
    outputs(479) <= not((layer0_outputs(1321)) xor (layer0_outputs(188)));
    outputs(480) <= not((layer0_outputs(726)) xor (layer0_outputs(1145)));
    outputs(481) <= not(layer0_outputs(2563));
    outputs(482) <= not(layer0_outputs(2008));
    outputs(483) <= not((layer0_outputs(4871)) xor (layer0_outputs(4624)));
    outputs(484) <= not(layer0_outputs(466));
    outputs(485) <= not((layer0_outputs(2836)) or (layer0_outputs(4624)));
    outputs(486) <= not((layer0_outputs(4780)) or (layer0_outputs(574)));
    outputs(487) <= not(layer0_outputs(4622));
    outputs(488) <= not((layer0_outputs(2854)) and (layer0_outputs(3444)));
    outputs(489) <= not(layer0_outputs(3401));
    outputs(490) <= not(layer0_outputs(1614));
    outputs(491) <= (layer0_outputs(2488)) and not (layer0_outputs(1947));
    outputs(492) <= (layer0_outputs(2113)) xor (layer0_outputs(3282));
    outputs(493) <= layer0_outputs(1718);
    outputs(494) <= layer0_outputs(3785);
    outputs(495) <= layer0_outputs(1827);
    outputs(496) <= not((layer0_outputs(696)) xor (layer0_outputs(229)));
    outputs(497) <= (layer0_outputs(1141)) and not (layer0_outputs(3150));
    outputs(498) <= layer0_outputs(2967);
    outputs(499) <= layer0_outputs(506);
    outputs(500) <= not(layer0_outputs(4358));
    outputs(501) <= layer0_outputs(4462);
    outputs(502) <= not(layer0_outputs(4751));
    outputs(503) <= layer0_outputs(3477);
    outputs(504) <= layer0_outputs(4639);
    outputs(505) <= not(layer0_outputs(3651));
    outputs(506) <= layer0_outputs(4277);
    outputs(507) <= not((layer0_outputs(597)) or (layer0_outputs(2549)));
    outputs(508) <= not(layer0_outputs(756));
    outputs(509) <= layer0_outputs(2415);
    outputs(510) <= not(layer0_outputs(1510));
    outputs(511) <= layer0_outputs(347);
    outputs(512) <= layer0_outputs(1779);
    outputs(513) <= (layer0_outputs(3291)) and not (layer0_outputs(2434));
    outputs(514) <= (layer0_outputs(2152)) and not (layer0_outputs(2677));
    outputs(515) <= (layer0_outputs(4204)) and not (layer0_outputs(2198));
    outputs(516) <= (layer0_outputs(2312)) and not (layer0_outputs(4352));
    outputs(517) <= not(layer0_outputs(2657));
    outputs(518) <= not((layer0_outputs(1833)) or (layer0_outputs(3625)));
    outputs(519) <= layer0_outputs(2598);
    outputs(520) <= layer0_outputs(2740);
    outputs(521) <= (layer0_outputs(707)) xor (layer0_outputs(1079));
    outputs(522) <= not((layer0_outputs(425)) or (layer0_outputs(1741)));
    outputs(523) <= (layer0_outputs(4876)) and (layer0_outputs(2102));
    outputs(524) <= (layer0_outputs(2961)) and (layer0_outputs(22));
    outputs(525) <= (layer0_outputs(503)) and not (layer0_outputs(671));
    outputs(526) <= not((layer0_outputs(3926)) or (layer0_outputs(4184)));
    outputs(527) <= not(layer0_outputs(3703));
    outputs(528) <= not(layer0_outputs(660));
    outputs(529) <= (layer0_outputs(1710)) and not (layer0_outputs(477));
    outputs(530) <= (layer0_outputs(2797)) and not (layer0_outputs(2238));
    outputs(531) <= (layer0_outputs(3763)) and not (layer0_outputs(5085));
    outputs(532) <= (layer0_outputs(148)) and (layer0_outputs(4378));
    outputs(533) <= not((layer0_outputs(4984)) or (layer0_outputs(4328)));
    outputs(534) <= (layer0_outputs(2681)) and (layer0_outputs(3356));
    outputs(535) <= (layer0_outputs(2618)) and not (layer0_outputs(1943));
    outputs(536) <= (layer0_outputs(4722)) and not (layer0_outputs(324));
    outputs(537) <= (layer0_outputs(3383)) and not (layer0_outputs(3618));
    outputs(538) <= (layer0_outputs(2551)) and not (layer0_outputs(29));
    outputs(539) <= (layer0_outputs(47)) and not (layer0_outputs(3026));
    outputs(540) <= (layer0_outputs(592)) and not (layer0_outputs(1245));
    outputs(541) <= not((layer0_outputs(2197)) or (layer0_outputs(2730)));
    outputs(542) <= not(layer0_outputs(3071));
    outputs(543) <= layer0_outputs(1044);
    outputs(544) <= (layer0_outputs(2055)) and not (layer0_outputs(3795));
    outputs(545) <= not((layer0_outputs(149)) or (layer0_outputs(4750)));
    outputs(546) <= (layer0_outputs(3108)) and not (layer0_outputs(2242));
    outputs(547) <= (layer0_outputs(33)) and not (layer0_outputs(2394));
    outputs(548) <= (layer0_outputs(1604)) xor (layer0_outputs(4337));
    outputs(549) <= layer0_outputs(2156);
    outputs(550) <= not((layer0_outputs(936)) or (layer0_outputs(2093)));
    outputs(551) <= (layer0_outputs(1924)) and not (layer0_outputs(2636));
    outputs(552) <= not(layer0_outputs(1234));
    outputs(553) <= (layer0_outputs(632)) and not (layer0_outputs(568));
    outputs(554) <= layer0_outputs(4534);
    outputs(555) <= not((layer0_outputs(2525)) or (layer0_outputs(3963)));
    outputs(556) <= (layer0_outputs(918)) and not (layer0_outputs(2427));
    outputs(557) <= (layer0_outputs(2716)) and not (layer0_outputs(630));
    outputs(558) <= not((layer0_outputs(1898)) or (layer0_outputs(3972)));
    outputs(559) <= not((layer0_outputs(282)) or (layer0_outputs(1275)));
    outputs(560) <= (layer0_outputs(1516)) and not (layer0_outputs(2234));
    outputs(561) <= (layer0_outputs(1001)) and not (layer0_outputs(2826));
    outputs(562) <= (layer0_outputs(2374)) and not (layer0_outputs(1119));
    outputs(563) <= layer0_outputs(3733);
    outputs(564) <= layer0_outputs(183);
    outputs(565) <= (layer0_outputs(3578)) xor (layer0_outputs(985));
    outputs(566) <= layer0_outputs(1879);
    outputs(567) <= not((layer0_outputs(2244)) or (layer0_outputs(4052)));
    outputs(568) <= layer0_outputs(3048);
    outputs(569) <= (layer0_outputs(197)) and (layer0_outputs(3999));
    outputs(570) <= not(layer0_outputs(2674));
    outputs(571) <= (layer0_outputs(258)) and not (layer0_outputs(5058));
    outputs(572) <= not((layer0_outputs(2183)) or (layer0_outputs(2662)));
    outputs(573) <= (layer0_outputs(152)) and not (layer0_outputs(2874));
    outputs(574) <= (layer0_outputs(1315)) and not (layer0_outputs(2486));
    outputs(575) <= (layer0_outputs(4146)) and not (layer0_outputs(2906));
    outputs(576) <= (layer0_outputs(3491)) and (layer0_outputs(1122));
    outputs(577) <= not((layer0_outputs(3490)) or (layer0_outputs(3828)));
    outputs(578) <= (layer0_outputs(3473)) and not (layer0_outputs(1281));
    outputs(579) <= not(layer0_outputs(496));
    outputs(580) <= layer0_outputs(62);
    outputs(581) <= (layer0_outputs(1393)) and not (layer0_outputs(946));
    outputs(582) <= (layer0_outputs(4655)) and (layer0_outputs(268));
    outputs(583) <= not((layer0_outputs(1212)) or (layer0_outputs(4127)));
    outputs(584) <= (layer0_outputs(691)) and not (layer0_outputs(2920));
    outputs(585) <= not((layer0_outputs(3506)) or (layer0_outputs(3809)));
    outputs(586) <= layer0_outputs(3365);
    outputs(587) <= (layer0_outputs(1149)) and (layer0_outputs(165));
    outputs(588) <= '0';
    outputs(589) <= (layer0_outputs(2661)) and (layer0_outputs(4790));
    outputs(590) <= not((layer0_outputs(1649)) or (layer0_outputs(2651)));
    outputs(591) <= layer0_outputs(3097);
    outputs(592) <= (layer0_outputs(3445)) and (layer0_outputs(2778));
    outputs(593) <= (layer0_outputs(2398)) and (layer0_outputs(1298));
    outputs(594) <= (layer0_outputs(2519)) and not (layer0_outputs(2817));
    outputs(595) <= not((layer0_outputs(2574)) or (layer0_outputs(3928)));
    outputs(596) <= (layer0_outputs(4927)) and (layer0_outputs(1582));
    outputs(597) <= (layer0_outputs(4087)) and not (layer0_outputs(1179));
    outputs(598) <= (layer0_outputs(4467)) and (layer0_outputs(340));
    outputs(599) <= not((layer0_outputs(2315)) or (layer0_outputs(2004)));
    outputs(600) <= (layer0_outputs(3180)) and (layer0_outputs(1780));
    outputs(601) <= (layer0_outputs(2930)) and not (layer0_outputs(2502));
    outputs(602) <= (layer0_outputs(203)) xor (layer0_outputs(3832));
    outputs(603) <= (layer0_outputs(5082)) and not (layer0_outputs(3516));
    outputs(604) <= (layer0_outputs(490)) and not (layer0_outputs(1383));
    outputs(605) <= not((layer0_outputs(1348)) or (layer0_outputs(2056)));
    outputs(606) <= layer0_outputs(3191);
    outputs(607) <= (layer0_outputs(2816)) and not (layer0_outputs(897));
    outputs(608) <= layer0_outputs(1216);
    outputs(609) <= not(layer0_outputs(3564));
    outputs(610) <= (layer0_outputs(2464)) and not (layer0_outputs(2741));
    outputs(611) <= (layer0_outputs(4558)) and not (layer0_outputs(1720));
    outputs(612) <= (layer0_outputs(14)) and (layer0_outputs(2405));
    outputs(613) <= (layer0_outputs(4809)) and not (layer0_outputs(552));
    outputs(614) <= (layer0_outputs(525)) and not (layer0_outputs(3076));
    outputs(615) <= not((layer0_outputs(3636)) or (layer0_outputs(1892)));
    outputs(616) <= (layer0_outputs(3511)) and not (layer0_outputs(1807));
    outputs(617) <= not((layer0_outputs(3302)) xor (layer0_outputs(2912)));
    outputs(618) <= not(layer0_outputs(4404));
    outputs(619) <= (layer0_outputs(3678)) and (layer0_outputs(815));
    outputs(620) <= not((layer0_outputs(2545)) or (layer0_outputs(962)));
    outputs(621) <= (layer0_outputs(153)) and not (layer0_outputs(2659));
    outputs(622) <= (layer0_outputs(2001)) and not (layer0_outputs(171));
    outputs(623) <= (layer0_outputs(2693)) and not (layer0_outputs(1858));
    outputs(624) <= not(layer0_outputs(4608));
    outputs(625) <= (layer0_outputs(813)) and (layer0_outputs(2235));
    outputs(626) <= layer0_outputs(2165);
    outputs(627) <= (layer0_outputs(4968)) and (layer0_outputs(1737));
    outputs(628) <= (layer0_outputs(2655)) and not (layer0_outputs(4513));
    outputs(629) <= not((layer0_outputs(906)) or (layer0_outputs(2734)));
    outputs(630) <= (layer0_outputs(3359)) and (layer0_outputs(44));
    outputs(631) <= (layer0_outputs(3824)) and (layer0_outputs(569));
    outputs(632) <= (layer0_outputs(1050)) and not (layer0_outputs(4699));
    outputs(633) <= (layer0_outputs(3749)) and not (layer0_outputs(2966));
    outputs(634) <= (layer0_outputs(1268)) and not (layer0_outputs(2705));
    outputs(635) <= (layer0_outputs(4236)) xor (layer0_outputs(3077));
    outputs(636) <= not(layer0_outputs(2866));
    outputs(637) <= (layer0_outputs(2229)) and (layer0_outputs(1486));
    outputs(638) <= (layer0_outputs(259)) xor (layer0_outputs(104));
    outputs(639) <= (layer0_outputs(3136)) and not (layer0_outputs(2183));
    outputs(640) <= not(layer0_outputs(602));
    outputs(641) <= layer0_outputs(4393);
    outputs(642) <= layer0_outputs(2801);
    outputs(643) <= layer0_outputs(5022);
    outputs(644) <= (layer0_outputs(4271)) and not (layer0_outputs(4911));
    outputs(645) <= (layer0_outputs(4399)) and not (layer0_outputs(4504));
    outputs(646) <= (layer0_outputs(2628)) and not (layer0_outputs(3492));
    outputs(647) <= (layer0_outputs(4585)) and (layer0_outputs(628));
    outputs(648) <= (layer0_outputs(4797)) and not (layer0_outputs(4322));
    outputs(649) <= (layer0_outputs(1307)) and (layer0_outputs(3299));
    outputs(650) <= (layer0_outputs(3525)) and not (layer0_outputs(2829));
    outputs(651) <= not((layer0_outputs(1485)) or (layer0_outputs(602)));
    outputs(652) <= (layer0_outputs(1642)) and not (layer0_outputs(1919));
    outputs(653) <= not((layer0_outputs(4615)) or (layer0_outputs(2214)));
    outputs(654) <= (layer0_outputs(1256)) and (layer0_outputs(3845));
    outputs(655) <= (layer0_outputs(98)) and (layer0_outputs(2138));
    outputs(656) <= not((layer0_outputs(1640)) and (layer0_outputs(4070)));
    outputs(657) <= not((layer0_outputs(4095)) or (layer0_outputs(1040)));
    outputs(658) <= (layer0_outputs(2799)) and (layer0_outputs(1081));
    outputs(659) <= not((layer0_outputs(318)) or (layer0_outputs(4110)));
    outputs(660) <= not(layer0_outputs(3343));
    outputs(661) <= (layer0_outputs(4148)) and not (layer0_outputs(3255));
    outputs(662) <= not(layer0_outputs(211));
    outputs(663) <= not(layer0_outputs(464));
    outputs(664) <= (layer0_outputs(4401)) and not (layer0_outputs(3508));
    outputs(665) <= not((layer0_outputs(3826)) or (layer0_outputs(1046)));
    outputs(666) <= (layer0_outputs(4568)) and not (layer0_outputs(3948));
    outputs(667) <= not((layer0_outputs(1621)) or (layer0_outputs(791)));
    outputs(668) <= not((layer0_outputs(5032)) or (layer0_outputs(2253)));
    outputs(669) <= not((layer0_outputs(1592)) or (layer0_outputs(2489)));
    outputs(670) <= not(layer0_outputs(20));
    outputs(671) <= layer0_outputs(3085);
    outputs(672) <= (layer0_outputs(870)) and not (layer0_outputs(4326));
    outputs(673) <= layer0_outputs(337);
    outputs(674) <= not((layer0_outputs(3371)) xor (layer0_outputs(3877)));
    outputs(675) <= (layer0_outputs(4638)) and not (layer0_outputs(4080));
    outputs(676) <= not(layer0_outputs(670));
    outputs(677) <= (layer0_outputs(4360)) and not (layer0_outputs(3035));
    outputs(678) <= '0';
    outputs(679) <= (layer0_outputs(1327)) and (layer0_outputs(2846));
    outputs(680) <= (layer0_outputs(2833)) and not (layer0_outputs(2702));
    outputs(681) <= (layer0_outputs(2329)) and not (layer0_outputs(2303));
    outputs(682) <= not(layer0_outputs(4612));
    outputs(683) <= (layer0_outputs(682)) and (layer0_outputs(1666));
    outputs(684) <= (layer0_outputs(3860)) and (layer0_outputs(2992));
    outputs(685) <= not(layer0_outputs(1638));
    outputs(686) <= (layer0_outputs(4584)) xor (layer0_outputs(4403));
    outputs(687) <= (layer0_outputs(4156)) and (layer0_outputs(299));
    outputs(688) <= not(layer0_outputs(2909));
    outputs(689) <= (layer0_outputs(2986)) xor (layer0_outputs(3622));
    outputs(690) <= not((layer0_outputs(4695)) or (layer0_outputs(3289)));
    outputs(691) <= '0';
    outputs(692) <= (layer0_outputs(4057)) and not (layer0_outputs(2361));
    outputs(693) <= (layer0_outputs(4108)) and not (layer0_outputs(3044));
    outputs(694) <= (layer0_outputs(460)) and not (layer0_outputs(2596));
    outputs(695) <= (layer0_outputs(2194)) and not (layer0_outputs(2205));
    outputs(696) <= (layer0_outputs(1142)) and not (layer0_outputs(2638));
    outputs(697) <= (layer0_outputs(4201)) and (layer0_outputs(3370));
    outputs(698) <= layer0_outputs(3104);
    outputs(699) <= (layer0_outputs(4894)) and not (layer0_outputs(1161));
    outputs(700) <= not((layer0_outputs(4084)) or (layer0_outputs(548)));
    outputs(701) <= (layer0_outputs(2178)) and (layer0_outputs(1543));
    outputs(702) <= not((layer0_outputs(2887)) or (layer0_outputs(958)));
    outputs(703) <= (layer0_outputs(1283)) and not (layer0_outputs(505));
    outputs(704) <= (layer0_outputs(911)) and not (layer0_outputs(4865));
    outputs(705) <= (layer0_outputs(3272)) and not (layer0_outputs(3487));
    outputs(706) <= (layer0_outputs(1207)) and (layer0_outputs(1266));
    outputs(707) <= not((layer0_outputs(4592)) or (layer0_outputs(4600)));
    outputs(708) <= not(layer0_outputs(3358));
    outputs(709) <= layer0_outputs(195);
    outputs(710) <= (layer0_outputs(3825)) and not (layer0_outputs(1154));
    outputs(711) <= (layer0_outputs(1849)) and (layer0_outputs(2831));
    outputs(712) <= not((layer0_outputs(1758)) or (layer0_outputs(3819)));
    outputs(713) <= not((layer0_outputs(3573)) xor (layer0_outputs(1195)));
    outputs(714) <= (layer0_outputs(69)) and (layer0_outputs(3709));
    outputs(715) <= (layer0_outputs(688)) and not (layer0_outputs(12));
    outputs(716) <= not((layer0_outputs(855)) xor (layer0_outputs(267)));
    outputs(717) <= (layer0_outputs(2633)) and not (layer0_outputs(4815));
    outputs(718) <= not(layer0_outputs(2324));
    outputs(719) <= not((layer0_outputs(3374)) or (layer0_outputs(2448)));
    outputs(720) <= not((layer0_outputs(4656)) or (layer0_outputs(2221)));
    outputs(721) <= not((layer0_outputs(4454)) or (layer0_outputs(2)));
    outputs(722) <= (layer0_outputs(763)) and (layer0_outputs(1391));
    outputs(723) <= not((layer0_outputs(3870)) or (layer0_outputs(3008)));
    outputs(724) <= not((layer0_outputs(2707)) or (layer0_outputs(4485)));
    outputs(725) <= (layer0_outputs(1520)) and (layer0_outputs(1841));
    outputs(726) <= not((layer0_outputs(2807)) or (layer0_outputs(2695)));
    outputs(727) <= (layer0_outputs(231)) and (layer0_outputs(3731));
    outputs(728) <= not((layer0_outputs(3685)) or (layer0_outputs(3510)));
    outputs(729) <= layer0_outputs(2511);
    outputs(730) <= (layer0_outputs(2449)) and (layer0_outputs(3249));
    outputs(731) <= (layer0_outputs(2162)) and not (layer0_outputs(964));
    outputs(732) <= (layer0_outputs(2870)) and not (layer0_outputs(439));
    outputs(733) <= not(layer0_outputs(3241));
    outputs(734) <= not((layer0_outputs(2686)) or (layer0_outputs(1732)));
    outputs(735) <= (layer0_outputs(2861)) and not (layer0_outputs(3750));
    outputs(736) <= (layer0_outputs(8)) and (layer0_outputs(5019));
    outputs(737) <= not(layer0_outputs(909));
    outputs(738) <= not(layer0_outputs(2059));
    outputs(739) <= (layer0_outputs(2531)) and (layer0_outputs(2986));
    outputs(740) <= (layer0_outputs(1448)) and not (layer0_outputs(4819));
    outputs(741) <= (layer0_outputs(3814)) and (layer0_outputs(742));
    outputs(742) <= (layer0_outputs(2040)) and not (layer0_outputs(2926));
    outputs(743) <= (layer0_outputs(1928)) and not (layer0_outputs(1529));
    outputs(744) <= not((layer0_outputs(1107)) or (layer0_outputs(3208)));
    outputs(745) <= (layer0_outputs(1159)) and (layer0_outputs(1446));
    outputs(746) <= not(layer0_outputs(2860));
    outputs(747) <= (layer0_outputs(3496)) and (layer0_outputs(4272));
    outputs(748) <= not(layer0_outputs(2883));
    outputs(749) <= '0';
    outputs(750) <= not((layer0_outputs(4849)) xor (layer0_outputs(1894)));
    outputs(751) <= (layer0_outputs(1327)) and (layer0_outputs(3777));
    outputs(752) <= not((layer0_outputs(3989)) or (layer0_outputs(2722)));
    outputs(753) <= not((layer0_outputs(3279)) or (layer0_outputs(717)));
    outputs(754) <= (layer0_outputs(2606)) and (layer0_outputs(3022));
    outputs(755) <= not(layer0_outputs(1911));
    outputs(756) <= not((layer0_outputs(2597)) or (layer0_outputs(993)));
    outputs(757) <= not(layer0_outputs(1748));
    outputs(758) <= (layer0_outputs(4383)) and not (layer0_outputs(3708));
    outputs(759) <= (layer0_outputs(2977)) and (layer0_outputs(2191));
    outputs(760) <= (layer0_outputs(4766)) and not (layer0_outputs(2363));
    outputs(761) <= not((layer0_outputs(1804)) or (layer0_outputs(4703)));
    outputs(762) <= not((layer0_outputs(892)) xor (layer0_outputs(262)));
    outputs(763) <= (layer0_outputs(4634)) and (layer0_outputs(4123));
    outputs(764) <= (layer0_outputs(314)) and not (layer0_outputs(2942));
    outputs(765) <= (layer0_outputs(8)) and (layer0_outputs(2715));
    outputs(766) <= layer0_outputs(3527);
    outputs(767) <= not((layer0_outputs(1408)) or (layer0_outputs(1650)));
    outputs(768) <= not(layer0_outputs(836));
    outputs(769) <= (layer0_outputs(3651)) and not (layer0_outputs(4220));
    outputs(770) <= (layer0_outputs(4409)) and not (layer0_outputs(315));
    outputs(771) <= (layer0_outputs(74)) and not (layer0_outputs(1975));
    outputs(772) <= '0';
    outputs(773) <= (layer0_outputs(545)) and not (layer0_outputs(1929));
    outputs(774) <= (layer0_outputs(341)) and not (layer0_outputs(102));
    outputs(775) <= (layer0_outputs(2934)) and not (layer0_outputs(3760));
    outputs(776) <= (layer0_outputs(4967)) and not (layer0_outputs(453));
    outputs(777) <= (layer0_outputs(2175)) and (layer0_outputs(2333));
    outputs(778) <= (layer0_outputs(3382)) and not (layer0_outputs(2019));
    outputs(779) <= not(layer0_outputs(584));
    outputs(780) <= (layer0_outputs(1262)) xor (layer0_outputs(4308));
    outputs(781) <= (layer0_outputs(3368)) and (layer0_outputs(4650));
    outputs(782) <= (layer0_outputs(2852)) or (layer0_outputs(4367));
    outputs(783) <= layer0_outputs(1008);
    outputs(784) <= (layer0_outputs(2572)) and not (layer0_outputs(4727));
    outputs(785) <= (layer0_outputs(3918)) and not (layer0_outputs(422));
    outputs(786) <= layer0_outputs(2109);
    outputs(787) <= not(layer0_outputs(1939)) or (layer0_outputs(1706));
    outputs(788) <= (layer0_outputs(468)) and not (layer0_outputs(4765));
    outputs(789) <= not((layer0_outputs(4860)) or (layer0_outputs(198)));
    outputs(790) <= (layer0_outputs(4700)) and not (layer0_outputs(840));
    outputs(791) <= (layer0_outputs(2029)) and not (layer0_outputs(4471));
    outputs(792) <= layer0_outputs(4575);
    outputs(793) <= (layer0_outputs(1878)) and (layer0_outputs(4899));
    outputs(794) <= not((layer0_outputs(1891)) or (layer0_outputs(4446)));
    outputs(795) <= (layer0_outputs(5110)) and (layer0_outputs(36));
    outputs(796) <= not(layer0_outputs(3434));
    outputs(797) <= (layer0_outputs(3259)) and not (layer0_outputs(2825));
    outputs(798) <= (layer0_outputs(3942)) and not (layer0_outputs(2718));
    outputs(799) <= not((layer0_outputs(2365)) xor (layer0_outputs(3393)));
    outputs(800) <= (layer0_outputs(2553)) and not (layer0_outputs(2473));
    outputs(801) <= '0';
    outputs(802) <= not((layer0_outputs(2311)) xor (layer0_outputs(140)));
    outputs(803) <= (layer0_outputs(2251)) and (layer0_outputs(2665));
    outputs(804) <= (layer0_outputs(1759)) and not (layer0_outputs(1136));
    outputs(805) <= not((layer0_outputs(4715)) or (layer0_outputs(2478)));
    outputs(806) <= not((layer0_outputs(4130)) xor (layer0_outputs(2915)));
    outputs(807) <= (layer0_outputs(559)) and (layer0_outputs(2994));
    outputs(808) <= (layer0_outputs(849)) xor (layer0_outputs(3739));
    outputs(809) <= (layer0_outputs(1574)) and not (layer0_outputs(3808));
    outputs(810) <= not((layer0_outputs(2508)) or (layer0_outputs(182)));
    outputs(811) <= (layer0_outputs(3563)) and not (layer0_outputs(884));
    outputs(812) <= (layer0_outputs(4779)) and not (layer0_outputs(5086));
    outputs(813) <= not((layer0_outputs(1914)) xor (layer0_outputs(739)));
    outputs(814) <= not((layer0_outputs(960)) or (layer0_outputs(1781)));
    outputs(815) <= (layer0_outputs(1196)) and not (layer0_outputs(3483));
    outputs(816) <= (layer0_outputs(400)) and (layer0_outputs(348));
    outputs(817) <= (layer0_outputs(3246)) and (layer0_outputs(2796));
    outputs(818) <= (layer0_outputs(4986)) and not (layer0_outputs(1174));
    outputs(819) <= (layer0_outputs(2416)) and not (layer0_outputs(2041));
    outputs(820) <= not((layer0_outputs(4145)) or (layer0_outputs(1465)));
    outputs(821) <= (layer0_outputs(2354)) and (layer0_outputs(4286));
    outputs(822) <= layer0_outputs(4900);
    outputs(823) <= layer0_outputs(1012);
    outputs(824) <= (layer0_outputs(4597)) and not (layer0_outputs(1168));
    outputs(825) <= not((layer0_outputs(1189)) xor (layer0_outputs(2699)));
    outputs(826) <= layer0_outputs(1045);
    outputs(827) <= not((layer0_outputs(2619)) xor (layer0_outputs(3005)));
    outputs(828) <= (layer0_outputs(4364)) xor (layer0_outputs(4614));
    outputs(829) <= (layer0_outputs(113)) and not (layer0_outputs(250));
    outputs(830) <= layer0_outputs(379);
    outputs(831) <= not(layer0_outputs(761));
    outputs(832) <= layer0_outputs(1324);
    outputs(833) <= (layer0_outputs(573)) and not (layer0_outputs(3094));
    outputs(834) <= not((layer0_outputs(4099)) or (layer0_outputs(276)));
    outputs(835) <= (layer0_outputs(947)) and (layer0_outputs(2757));
    outputs(836) <= not((layer0_outputs(3266)) or (layer0_outputs(2239)));
    outputs(837) <= (layer0_outputs(4257)) and not (layer0_outputs(3652));
    outputs(838) <= not((layer0_outputs(2106)) or (layer0_outputs(3241)));
    outputs(839) <= not((layer0_outputs(402)) or (layer0_outputs(4793)));
    outputs(840) <= layer0_outputs(139);
    outputs(841) <= '0';
    outputs(842) <= (layer0_outputs(1830)) and (layer0_outputs(2703));
    outputs(843) <= (layer0_outputs(4100)) and not (layer0_outputs(4977));
    outputs(844) <= (layer0_outputs(3468)) and (layer0_outputs(3860));
    outputs(845) <= (layer0_outputs(2195)) and (layer0_outputs(4176));
    outputs(846) <= (layer0_outputs(3609)) and not (layer0_outputs(1790));
    outputs(847) <= not(layer0_outputs(2689));
    outputs(848) <= not((layer0_outputs(2221)) or (layer0_outputs(4926)));
    outputs(849) <= (layer0_outputs(3878)) and not (layer0_outputs(4735));
    outputs(850) <= (layer0_outputs(728)) and not (layer0_outputs(575));
    outputs(851) <= (layer0_outputs(1325)) xor (layer0_outputs(1762));
    outputs(852) <= (layer0_outputs(2206)) and not (layer0_outputs(4677));
    outputs(853) <= layer0_outputs(950);
    outputs(854) <= (layer0_outputs(640)) and (layer0_outputs(3405));
    outputs(855) <= (layer0_outputs(870)) and not (layer0_outputs(2657));
    outputs(856) <= (layer0_outputs(1181)) and not (layer0_outputs(3173));
    outputs(857) <= not((layer0_outputs(3063)) or (layer0_outputs(2052)));
    outputs(858) <= (layer0_outputs(1848)) and not (layer0_outputs(846));
    outputs(859) <= (layer0_outputs(85)) and (layer0_outputs(2318));
    outputs(860) <= (layer0_outputs(2274)) or (layer0_outputs(2432));
    outputs(861) <= not((layer0_outputs(4483)) xor (layer0_outputs(1181)));
    outputs(862) <= not(layer0_outputs(30));
    outputs(863) <= (layer0_outputs(3829)) and not (layer0_outputs(288));
    outputs(864) <= not((layer0_outputs(1244)) or (layer0_outputs(4707)));
    outputs(865) <= (layer0_outputs(2396)) and not (layer0_outputs(4265));
    outputs(866) <= not((layer0_outputs(3082)) xor (layer0_outputs(4437)));
    outputs(867) <= layer0_outputs(3696);
    outputs(868) <= (layer0_outputs(2248)) and not (layer0_outputs(3325));
    outputs(869) <= not((layer0_outputs(1624)) xor (layer0_outputs(2805)));
    outputs(870) <= layer0_outputs(4778);
    outputs(871) <= (layer0_outputs(4757)) and (layer0_outputs(3171));
    outputs(872) <= not(layer0_outputs(1151));
    outputs(873) <= not((layer0_outputs(4581)) or (layer0_outputs(217)));
    outputs(874) <= (layer0_outputs(2405)) and (layer0_outputs(471));
    outputs(875) <= (layer0_outputs(801)) and not (layer0_outputs(4696));
    outputs(876) <= layer0_outputs(2414);
    outputs(877) <= (layer0_outputs(1185)) and not (layer0_outputs(1025));
    outputs(878) <= (layer0_outputs(1472)) and not (layer0_outputs(2417));
    outputs(879) <= (layer0_outputs(2293)) and not (layer0_outputs(2959));
    outputs(880) <= layer0_outputs(661);
    outputs(881) <= (layer0_outputs(787)) and (layer0_outputs(224));
    outputs(882) <= (layer0_outputs(3588)) and (layer0_outputs(204));
    outputs(883) <= (layer0_outputs(1312)) and not (layer0_outputs(450));
    outputs(884) <= not((layer0_outputs(2959)) or (layer0_outputs(4536)));
    outputs(885) <= (layer0_outputs(3503)) and not (layer0_outputs(3007));
    outputs(886) <= (layer0_outputs(3481)) and not (layer0_outputs(4280));
    outputs(887) <= (layer0_outputs(2591)) and (layer0_outputs(1974));
    outputs(888) <= not((layer0_outputs(159)) or (layer0_outputs(2349)));
    outputs(889) <= (layer0_outputs(3110)) and not (layer0_outputs(3759));
    outputs(890) <= (layer0_outputs(2768)) and not (layer0_outputs(579));
    outputs(891) <= (layer0_outputs(944)) and not (layer0_outputs(3336));
    outputs(892) <= (layer0_outputs(274)) and (layer0_outputs(4327));
    outputs(893) <= (layer0_outputs(68)) and not (layer0_outputs(4186));
    outputs(894) <= (layer0_outputs(2630)) and (layer0_outputs(820));
    outputs(895) <= layer0_outputs(2554);
    outputs(896) <= not((layer0_outputs(1718)) or (layer0_outputs(4232)));
    outputs(897) <= (layer0_outputs(3867)) and (layer0_outputs(22));
    outputs(898) <= (layer0_outputs(1463)) and not (layer0_outputs(3258));
    outputs(899) <= (layer0_outputs(4431)) and (layer0_outputs(3544));
    outputs(900) <= (layer0_outputs(2554)) and not (layer0_outputs(1129));
    outputs(901) <= layer0_outputs(3554);
    outputs(902) <= not(layer0_outputs(2692));
    outputs(903) <= (layer0_outputs(4026)) and not (layer0_outputs(2485));
    outputs(904) <= not((layer0_outputs(4187)) and (layer0_outputs(1529)));
    outputs(905) <= layer0_outputs(2023);
    outputs(906) <= not((layer0_outputs(3460)) or (layer0_outputs(1177)));
    outputs(907) <= (layer0_outputs(2724)) and not (layer0_outputs(716));
    outputs(908) <= not(layer0_outputs(3332));
    outputs(909) <= not(layer0_outputs(4565));
    outputs(910) <= not(layer0_outputs(2177)) or (layer0_outputs(4553));
    outputs(911) <= (layer0_outputs(834)) and (layer0_outputs(3589));
    outputs(912) <= not(layer0_outputs(593));
    outputs(913) <= not(layer0_outputs(2147));
    outputs(914) <= not((layer0_outputs(1947)) or (layer0_outputs(360)));
    outputs(915) <= not((layer0_outputs(708)) or (layer0_outputs(1139)));
    outputs(916) <= (layer0_outputs(938)) xor (layer0_outputs(573));
    outputs(917) <= not(layer0_outputs(4953));
    outputs(918) <= not((layer0_outputs(170)) or (layer0_outputs(84)));
    outputs(919) <= (layer0_outputs(1976)) and not (layer0_outputs(2704));
    outputs(920) <= (layer0_outputs(2877)) and not (layer0_outputs(3285));
    outputs(921) <= (layer0_outputs(3242)) and (layer0_outputs(886));
    outputs(922) <= '0';
    outputs(923) <= not(layer0_outputs(686));
    outputs(924) <= not((layer0_outputs(2297)) or (layer0_outputs(2428)));
    outputs(925) <= (layer0_outputs(469)) and not (layer0_outputs(352));
    outputs(926) <= layer0_outputs(121);
    outputs(927) <= (layer0_outputs(3935)) and not (layer0_outputs(2793));
    outputs(928) <= not(layer0_outputs(3216));
    outputs(929) <= (layer0_outputs(2978)) and not (layer0_outputs(4752));
    outputs(930) <= layer0_outputs(1734);
    outputs(931) <= layer0_outputs(1020);
    outputs(932) <= (layer0_outputs(3251)) and (layer0_outputs(1598));
    outputs(933) <= (layer0_outputs(723)) and not (layer0_outputs(4104));
    outputs(934) <= (layer0_outputs(90)) and (layer0_outputs(606));
    outputs(935) <= not((layer0_outputs(182)) or (layer0_outputs(2066)));
    outputs(936) <= (layer0_outputs(5068)) and not (layer0_outputs(24));
    outputs(937) <= (layer0_outputs(1082)) and not (layer0_outputs(3253));
    outputs(938) <= (layer0_outputs(3116)) and not (layer0_outputs(788));
    outputs(939) <= not((layer0_outputs(776)) xor (layer0_outputs(3004)));
    outputs(940) <= not((layer0_outputs(1359)) or (layer0_outputs(1151)));
    outputs(941) <= '0';
    outputs(942) <= layer0_outputs(4129);
    outputs(943) <= not(layer0_outputs(1246));
    outputs(944) <= (layer0_outputs(2512)) and not (layer0_outputs(3523));
    outputs(945) <= (layer0_outputs(1141)) xor (layer0_outputs(1535));
    outputs(946) <= (layer0_outputs(1378)) and not (layer0_outputs(2164));
    outputs(947) <= (layer0_outputs(792)) and (layer0_outputs(2020));
    outputs(948) <= (layer0_outputs(1034)) and not (layer0_outputs(174));
    outputs(949) <= (layer0_outputs(1835)) and (layer0_outputs(622));
    outputs(950) <= not((layer0_outputs(1970)) or (layer0_outputs(3870)));
    outputs(951) <= (layer0_outputs(2257)) and not (layer0_outputs(2567));
    outputs(952) <= (layer0_outputs(4330)) and not (layer0_outputs(3983));
    outputs(953) <= layer0_outputs(2144);
    outputs(954) <= not(layer0_outputs(240));
    outputs(955) <= (layer0_outputs(1369)) and (layer0_outputs(4782));
    outputs(956) <= (layer0_outputs(376)) and not (layer0_outputs(3773));
    outputs(957) <= (layer0_outputs(1587)) and not (layer0_outputs(146));
    outputs(958) <= (layer0_outputs(5105)) and (layer0_outputs(1509));
    outputs(959) <= (layer0_outputs(725)) and (layer0_outputs(3974));
    outputs(960) <= (layer0_outputs(4356)) and not (layer0_outputs(2369));
    outputs(961) <= not((layer0_outputs(1807)) or (layer0_outputs(2063)));
    outputs(962) <= layer0_outputs(1183);
    outputs(963) <= not(layer0_outputs(3313));
    outputs(964) <= not(layer0_outputs(1735));
    outputs(965) <= (layer0_outputs(4882)) and (layer0_outputs(474));
    outputs(966) <= not(layer0_outputs(5119));
    outputs(967) <= (layer0_outputs(976)) and not (layer0_outputs(470));
    outputs(968) <= (layer0_outputs(4042)) and (layer0_outputs(2994));
    outputs(969) <= (layer0_outputs(3603)) and not (layer0_outputs(1948));
    outputs(970) <= layer0_outputs(569);
    outputs(971) <= not((layer0_outputs(3715)) or (layer0_outputs(3195)));
    outputs(972) <= not((layer0_outputs(2352)) or (layer0_outputs(1306)));
    outputs(973) <= not((layer0_outputs(4084)) or (layer0_outputs(3590)));
    outputs(974) <= (layer0_outputs(2572)) and not (layer0_outputs(4334));
    outputs(975) <= not(layer0_outputs(831));
    outputs(976) <= (layer0_outputs(3544)) and not (layer0_outputs(4573));
    outputs(977) <= (layer0_outputs(558)) and not (layer0_outputs(2971));
    outputs(978) <= (layer0_outputs(880)) and not (layer0_outputs(903));
    outputs(979) <= (layer0_outputs(2899)) and not (layer0_outputs(1212));
    outputs(980) <= (layer0_outputs(5089)) and (layer0_outputs(1904));
    outputs(981) <= not((layer0_outputs(1742)) or (layer0_outputs(3028)));
    outputs(982) <= layer0_outputs(2535);
    outputs(983) <= (layer0_outputs(3171)) and (layer0_outputs(966));
    outputs(984) <= (layer0_outputs(2669)) and (layer0_outputs(1616));
    outputs(985) <= not((layer0_outputs(492)) or (layer0_outputs(371)));
    outputs(986) <= (layer0_outputs(4189)) xor (layer0_outputs(4855));
    outputs(987) <= (layer0_outputs(1751)) and (layer0_outputs(5062));
    outputs(988) <= (layer0_outputs(1569)) and (layer0_outputs(5055));
    outputs(989) <= '0';
    outputs(990) <= (layer0_outputs(3672)) and not (layer0_outputs(2215));
    outputs(991) <= (layer0_outputs(598)) and not (layer0_outputs(3434));
    outputs(992) <= '0';
    outputs(993) <= not((layer0_outputs(3293)) xor (layer0_outputs(3524)));
    outputs(994) <= (layer0_outputs(4787)) and not (layer0_outputs(4902));
    outputs(995) <= not((layer0_outputs(4859)) or (layer0_outputs(2005)));
    outputs(996) <= (layer0_outputs(3807)) and not (layer0_outputs(2078));
    outputs(997) <= (layer0_outputs(3834)) and not (layer0_outputs(4936));
    outputs(998) <= not(layer0_outputs(2714));
    outputs(999) <= (layer0_outputs(2513)) and not (layer0_outputs(3236));
    outputs(1000) <= (layer0_outputs(1374)) and not (layer0_outputs(4061));
    outputs(1001) <= (layer0_outputs(3503)) and not (layer0_outputs(189));
    outputs(1002) <= not((layer0_outputs(737)) or (layer0_outputs(645)));
    outputs(1003) <= (layer0_outputs(3638)) and not (layer0_outputs(5091));
    outputs(1004) <= (layer0_outputs(2709)) and not (layer0_outputs(1643));
    outputs(1005) <= (layer0_outputs(462)) xor (layer0_outputs(643));
    outputs(1006) <= (layer0_outputs(2816)) and (layer0_outputs(3507));
    outputs(1007) <= layer0_outputs(4540);
    outputs(1008) <= not((layer0_outputs(3318)) or (layer0_outputs(1749)));
    outputs(1009) <= (layer0_outputs(4166)) and not (layer0_outputs(2430));
    outputs(1010) <= not((layer0_outputs(731)) or (layer0_outputs(1629)));
    outputs(1011) <= layer0_outputs(1334);
    outputs(1012) <= (layer0_outputs(3876)) and not (layer0_outputs(3210));
    outputs(1013) <= not((layer0_outputs(4285)) xor (layer0_outputs(644)));
    outputs(1014) <= not((layer0_outputs(4979)) xor (layer0_outputs(4602)));
    outputs(1015) <= (layer0_outputs(3733)) and (layer0_outputs(4346));
    outputs(1016) <= layer0_outputs(2544);
    outputs(1017) <= not((layer0_outputs(1166)) or (layer0_outputs(2079)));
    outputs(1018) <= (layer0_outputs(4256)) and not (layer0_outputs(1247));
    outputs(1019) <= (layer0_outputs(2333)) and not (layer0_outputs(4314));
    outputs(1020) <= (layer0_outputs(4111)) and (layer0_outputs(4684));
    outputs(1021) <= not((layer0_outputs(3985)) or (layer0_outputs(4022)));
    outputs(1022) <= layer0_outputs(2000);
    outputs(1023) <= (layer0_outputs(3511)) and (layer0_outputs(4477));
    outputs(1024) <= not(layer0_outputs(1610));
    outputs(1025) <= not(layer0_outputs(1325));
    outputs(1026) <= not((layer0_outputs(4019)) or (layer0_outputs(2154)));
    outputs(1027) <= not(layer0_outputs(430));
    outputs(1028) <= (layer0_outputs(1188)) or (layer0_outputs(2419));
    outputs(1029) <= (layer0_outputs(1094)) and (layer0_outputs(4303));
    outputs(1030) <= layer0_outputs(2426);
    outputs(1031) <= (layer0_outputs(1828)) and not (layer0_outputs(3421));
    outputs(1032) <= (layer0_outputs(3102)) and not (layer0_outputs(1399));
    outputs(1033) <= layer0_outputs(3649);
    outputs(1034) <= not(layer0_outputs(1851)) or (layer0_outputs(2975));
    outputs(1035) <= (layer0_outputs(3226)) and (layer0_outputs(4386));
    outputs(1036) <= layer0_outputs(4305);
    outputs(1037) <= not((layer0_outputs(2763)) and (layer0_outputs(3669)));
    outputs(1038) <= layer0_outputs(4239);
    outputs(1039) <= layer0_outputs(61);
    outputs(1040) <= (layer0_outputs(1771)) and not (layer0_outputs(3439));
    outputs(1041) <= not(layer0_outputs(4756));
    outputs(1042) <= layer0_outputs(66);
    outputs(1043) <= layer0_outputs(3808);
    outputs(1044) <= (layer0_outputs(1620)) and (layer0_outputs(3554));
    outputs(1045) <= layer0_outputs(597);
    outputs(1046) <= not((layer0_outputs(67)) and (layer0_outputs(4825)));
    outputs(1047) <= not(layer0_outputs(567));
    outputs(1048) <= layer0_outputs(2496);
    outputs(1049) <= layer0_outputs(5100);
    outputs(1050) <= not(layer0_outputs(1323));
    outputs(1051) <= not(layer0_outputs(3601));
    outputs(1052) <= not(layer0_outputs(2772));
    outputs(1053) <= (layer0_outputs(1222)) xor (layer0_outputs(1749));
    outputs(1054) <= not((layer0_outputs(3849)) xor (layer0_outputs(1031)));
    outputs(1055) <= not((layer0_outputs(1852)) and (layer0_outputs(4411)));
    outputs(1056) <= layer0_outputs(980);
    outputs(1057) <= not((layer0_outputs(2334)) and (layer0_outputs(1855)));
    outputs(1058) <= (layer0_outputs(2908)) or (layer0_outputs(4651));
    outputs(1059) <= not(layer0_outputs(2615));
    outputs(1060) <= not(layer0_outputs(364));
    outputs(1061) <= (layer0_outputs(1121)) or (layer0_outputs(2956));
    outputs(1062) <= not((layer0_outputs(5109)) and (layer0_outputs(3575)));
    outputs(1063) <= not(layer0_outputs(397));
    outputs(1064) <= not(layer0_outputs(2459)) or (layer0_outputs(2911));
    outputs(1065) <= not(layer0_outputs(4552));
    outputs(1066) <= not(layer0_outputs(4406));
    outputs(1067) <= not(layer0_outputs(491));
    outputs(1068) <= (layer0_outputs(439)) or (layer0_outputs(2141));
    outputs(1069) <= layer0_outputs(2167);
    outputs(1070) <= layer0_outputs(3704);
    outputs(1071) <= not((layer0_outputs(1899)) or (layer0_outputs(2212)));
    outputs(1072) <= layer0_outputs(1716);
    outputs(1073) <= not(layer0_outputs(644));
    outputs(1074) <= layer0_outputs(3419);
    outputs(1075) <= not(layer0_outputs(1991));
    outputs(1076) <= not(layer0_outputs(2121));
    outputs(1077) <= layer0_outputs(4448);
    outputs(1078) <= not(layer0_outputs(3561));
    outputs(1079) <= not(layer0_outputs(1765)) or (layer0_outputs(2345));
    outputs(1080) <= not(layer0_outputs(4872));
    outputs(1081) <= layer0_outputs(785);
    outputs(1082) <= layer0_outputs(1125);
    outputs(1083) <= not(layer0_outputs(2243));
    outputs(1084) <= (layer0_outputs(3292)) xor (layer0_outputs(1409));
    outputs(1085) <= layer0_outputs(2690);
    outputs(1086) <= not(layer0_outputs(287));
    outputs(1087) <= layer0_outputs(3469);
    outputs(1088) <= layer0_outputs(2603);
    outputs(1089) <= layer0_outputs(1442);
    outputs(1090) <= not(layer0_outputs(307));
    outputs(1091) <= layer0_outputs(3012);
    outputs(1092) <= not((layer0_outputs(1600)) xor (layer0_outputs(973)));
    outputs(1093) <= not(layer0_outputs(3648)) or (layer0_outputs(2304));
    outputs(1094) <= not(layer0_outputs(5008));
    outputs(1095) <= not(layer0_outputs(4416));
    outputs(1096) <= not(layer0_outputs(4390));
    outputs(1097) <= layer0_outputs(1132);
    outputs(1098) <= layer0_outputs(1311);
    outputs(1099) <= (layer0_outputs(4674)) and (layer0_outputs(3913));
    outputs(1100) <= (layer0_outputs(3990)) xor (layer0_outputs(2584));
    outputs(1101) <= not(layer0_outputs(3206));
    outputs(1102) <= layer0_outputs(4931);
    outputs(1103) <= (layer0_outputs(4207)) and (layer0_outputs(659));
    outputs(1104) <= layer0_outputs(3124);
    outputs(1105) <= not(layer0_outputs(1675));
    outputs(1106) <= not(layer0_outputs(2155));
    outputs(1107) <= layer0_outputs(2269);
    outputs(1108) <= not(layer0_outputs(2579)) or (layer0_outputs(4739));
    outputs(1109) <= (layer0_outputs(4343)) xor (layer0_outputs(4276));
    outputs(1110) <= not((layer0_outputs(7)) xor (layer0_outputs(3965)));
    outputs(1111) <= layer0_outputs(1157);
    outputs(1112) <= not(layer0_outputs(3737));
    outputs(1113) <= (layer0_outputs(3977)) or (layer0_outputs(2067));
    outputs(1114) <= not((layer0_outputs(2265)) or (layer0_outputs(914)));
    outputs(1115) <= (layer0_outputs(1398)) xor (layer0_outputs(1968));
    outputs(1116) <= not(layer0_outputs(3770));
    outputs(1117) <= layer0_outputs(1136);
    outputs(1118) <= layer0_outputs(2950);
    outputs(1119) <= (layer0_outputs(1566)) xor (layer0_outputs(2758));
    outputs(1120) <= not((layer0_outputs(128)) and (layer0_outputs(832)));
    outputs(1121) <= layer0_outputs(3182);
    outputs(1122) <= (layer0_outputs(2734)) xor (layer0_outputs(3973));
    outputs(1123) <= not(layer0_outputs(3474));
    outputs(1124) <= layer0_outputs(101);
    outputs(1125) <= not(layer0_outputs(4708));
    outputs(1126) <= not(layer0_outputs(1899));
    outputs(1127) <= not(layer0_outputs(1733));
    outputs(1128) <= (layer0_outputs(146)) and not (layer0_outputs(2125));
    outputs(1129) <= (layer0_outputs(1085)) xor (layer0_outputs(5098));
    outputs(1130) <= layer0_outputs(2526);
    outputs(1131) <= not(layer0_outputs(429));
    outputs(1132) <= not((layer0_outputs(3979)) and (layer0_outputs(1809)));
    outputs(1133) <= (layer0_outputs(821)) xor (layer0_outputs(3740));
    outputs(1134) <= (layer0_outputs(297)) and not (layer0_outputs(4794));
    outputs(1135) <= (layer0_outputs(3818)) xor (layer0_outputs(1756));
    outputs(1136) <= (layer0_outputs(3624)) xor (layer0_outputs(885));
    outputs(1137) <= layer0_outputs(4010);
    outputs(1138) <= layer0_outputs(3307);
    outputs(1139) <= layer0_outputs(4674);
    outputs(1140) <= (layer0_outputs(4777)) xor (layer0_outputs(4190));
    outputs(1141) <= (layer0_outputs(657)) and not (layer0_outputs(2453));
    outputs(1142) <= not((layer0_outputs(1550)) and (layer0_outputs(4570)));
    outputs(1143) <= layer0_outputs(4065);
    outputs(1144) <= not(layer0_outputs(3555));
    outputs(1145) <= not(layer0_outputs(3161));
    outputs(1146) <= not(layer0_outputs(2945));
    outputs(1147) <= (layer0_outputs(1472)) and not (layer0_outputs(4482));
    outputs(1148) <= not(layer0_outputs(2620)) or (layer0_outputs(1994));
    outputs(1149) <= (layer0_outputs(2972)) and not (layer0_outputs(121));
    outputs(1150) <= not(layer0_outputs(2587));
    outputs(1151) <= layer0_outputs(3661);
    outputs(1152) <= (layer0_outputs(2813)) or (layer0_outputs(4946));
    outputs(1153) <= layer0_outputs(3772);
    outputs(1154) <= not(layer0_outputs(2701));
    outputs(1155) <= layer0_outputs(2113);
    outputs(1156) <= not((layer0_outputs(727)) xor (layer0_outputs(4248)));
    outputs(1157) <= not((layer0_outputs(199)) or (layer0_outputs(60)));
    outputs(1158) <= not((layer0_outputs(3066)) and (layer0_outputs(2127)));
    outputs(1159) <= not(layer0_outputs(489));
    outputs(1160) <= layer0_outputs(880);
    outputs(1161) <= layer0_outputs(4578);
    outputs(1162) <= not(layer0_outputs(37));
    outputs(1163) <= not(layer0_outputs(2685)) or (layer0_outputs(2914));
    outputs(1164) <= not((layer0_outputs(4881)) and (layer0_outputs(4478)));
    outputs(1165) <= layer0_outputs(3881);
    outputs(1166) <= layer0_outputs(1821);
    outputs(1167) <= not(layer0_outputs(3820)) or (layer0_outputs(4850));
    outputs(1168) <= not((layer0_outputs(4215)) and (layer0_outputs(3907)));
    outputs(1169) <= not(layer0_outputs(1239)) or (layer0_outputs(312));
    outputs(1170) <= (layer0_outputs(1374)) and not (layer0_outputs(1979));
    outputs(1171) <= layer0_outputs(3025);
    outputs(1172) <= (layer0_outputs(747)) and not (layer0_outputs(3674));
    outputs(1173) <= (layer0_outputs(5011)) or (layer0_outputs(803));
    outputs(1174) <= not(layer0_outputs(316));
    outputs(1175) <= not(layer0_outputs(1048));
    outputs(1176) <= not(layer0_outputs(1965)) or (layer0_outputs(2342));
    outputs(1177) <= (layer0_outputs(778)) or (layer0_outputs(1262));
    outputs(1178) <= not((layer0_outputs(1853)) xor (layer0_outputs(3090)));
    outputs(1179) <= not(layer0_outputs(1617));
    outputs(1180) <= (layer0_outputs(1776)) and not (layer0_outputs(2868));
    outputs(1181) <= not(layer0_outputs(4898));
    outputs(1182) <= not(layer0_outputs(424));
    outputs(1183) <= not((layer0_outputs(3668)) and (layer0_outputs(73)));
    outputs(1184) <= not((layer0_outputs(2998)) xor (layer0_outputs(3510)));
    outputs(1185) <= layer0_outputs(2381);
    outputs(1186) <= not(layer0_outputs(4362));
    outputs(1187) <= not(layer0_outputs(3847));
    outputs(1188) <= layer0_outputs(2010);
    outputs(1189) <= (layer0_outputs(1583)) xor (layer0_outputs(926));
    outputs(1190) <= not((layer0_outputs(1313)) and (layer0_outputs(2467)));
    outputs(1191) <= not(layer0_outputs(3273)) or (layer0_outputs(1355));
    outputs(1192) <= layer0_outputs(3017);
    outputs(1193) <= not(layer0_outputs(2885));
    outputs(1194) <= not(layer0_outputs(1601));
    outputs(1195) <= layer0_outputs(2319);
    outputs(1196) <= layer0_outputs(744);
    outputs(1197) <= not((layer0_outputs(3735)) xor (layer0_outputs(4868)));
    outputs(1198) <= (layer0_outputs(4445)) and not (layer0_outputs(3505));
    outputs(1199) <= layer0_outputs(3543);
    outputs(1200) <= (layer0_outputs(63)) or (layer0_outputs(137));
    outputs(1201) <= layer0_outputs(2174);
    outputs(1202) <= (layer0_outputs(1389)) and not (layer0_outputs(765));
    outputs(1203) <= layer0_outputs(878);
    outputs(1204) <= (layer0_outputs(103)) and (layer0_outputs(3579));
    outputs(1205) <= not(layer0_outputs(3587));
    outputs(1206) <= not((layer0_outputs(2230)) xor (layer0_outputs(2819)));
    outputs(1207) <= layer0_outputs(580);
    outputs(1208) <= not((layer0_outputs(2543)) or (layer0_outputs(1008)));
    outputs(1209) <= not(layer0_outputs(3020));
    outputs(1210) <= not(layer0_outputs(4296));
    outputs(1211) <= layer0_outputs(5081);
    outputs(1212) <= not(layer0_outputs(2082)) or (layer0_outputs(32));
    outputs(1213) <= not(layer0_outputs(46)) or (layer0_outputs(4693));
    outputs(1214) <= not(layer0_outputs(333)) or (layer0_outputs(4444));
    outputs(1215) <= layer0_outputs(4853);
    outputs(1216) <= layer0_outputs(1462);
    outputs(1217) <= not(layer0_outputs(3263)) or (layer0_outputs(444));
    outputs(1218) <= layer0_outputs(4448);
    outputs(1219) <= not(layer0_outputs(4015));
    outputs(1220) <= layer0_outputs(2666);
    outputs(1221) <= layer0_outputs(1389);
    outputs(1222) <= not(layer0_outputs(344));
    outputs(1223) <= layer0_outputs(4937);
    outputs(1224) <= not((layer0_outputs(3193)) xor (layer0_outputs(2104)));
    outputs(1225) <= layer0_outputs(3697);
    outputs(1226) <= not(layer0_outputs(2438)) or (layer0_outputs(3853));
    outputs(1227) <= layer0_outputs(319);
    outputs(1228) <= (layer0_outputs(1337)) and (layer0_outputs(3630));
    outputs(1229) <= layer0_outputs(4632);
    outputs(1230) <= not((layer0_outputs(2084)) or (layer0_outputs(4193)));
    outputs(1231) <= layer0_outputs(2914);
    outputs(1232) <= layer0_outputs(3391);
    outputs(1233) <= not(layer0_outputs(5009)) or (layer0_outputs(4085));
    outputs(1234) <= (layer0_outputs(4610)) xor (layer0_outputs(1281));
    outputs(1235) <= layer0_outputs(767);
    outputs(1236) <= not(layer0_outputs(1714));
    outputs(1237) <= not((layer0_outputs(2143)) xor (layer0_outputs(3225)));
    outputs(1238) <= layer0_outputs(3139);
    outputs(1239) <= not(layer0_outputs(4426)) or (layer0_outputs(3398));
    outputs(1240) <= not(layer0_outputs(4186));
    outputs(1241) <= (layer0_outputs(1775)) and not (layer0_outputs(4885));
    outputs(1242) <= (layer0_outputs(2051)) or (layer0_outputs(675));
    outputs(1243) <= (layer0_outputs(4673)) and not (layer0_outputs(177));
    outputs(1244) <= not(layer0_outputs(1972));
    outputs(1245) <= not(layer0_outputs(2191));
    outputs(1246) <= (layer0_outputs(4618)) and not (layer0_outputs(4760));
    outputs(1247) <= not(layer0_outputs(1464)) or (layer0_outputs(2252));
    outputs(1248) <= layer0_outputs(4242);
    outputs(1249) <= not((layer0_outputs(4494)) and (layer0_outputs(4530)));
    outputs(1250) <= not((layer0_outputs(4159)) xor (layer0_outputs(3116)));
    outputs(1251) <= (layer0_outputs(654)) or (layer0_outputs(3278));
    outputs(1252) <= not(layer0_outputs(4873)) or (layer0_outputs(408));
    outputs(1253) <= not(layer0_outputs(3724));
    outputs(1254) <= not(layer0_outputs(2701));
    outputs(1255) <= not(layer0_outputs(2723)) or (layer0_outputs(3684));
    outputs(1256) <= (layer0_outputs(534)) and (layer0_outputs(2182));
    outputs(1257) <= layer0_outputs(2007);
    outputs(1258) <= (layer0_outputs(4612)) or (layer0_outputs(3438));
    outputs(1259) <= (layer0_outputs(3509)) and not (layer0_outputs(4981));
    outputs(1260) <= layer0_outputs(2969);
    outputs(1261) <= not(layer0_outputs(2466));
    outputs(1262) <= not((layer0_outputs(2812)) and (layer0_outputs(1513)));
    outputs(1263) <= (layer0_outputs(1736)) and (layer0_outputs(1630));
    outputs(1264) <= not(layer0_outputs(2164)) or (layer0_outputs(3766));
    outputs(1265) <= not(layer0_outputs(2532));
    outputs(1266) <= (layer0_outputs(2349)) and (layer0_outputs(2835));
    outputs(1267) <= not(layer0_outputs(614));
    outputs(1268) <= not(layer0_outputs(2821));
    outputs(1269) <= (layer0_outputs(1820)) or (layer0_outputs(876));
    outputs(1270) <= not((layer0_outputs(424)) and (layer0_outputs(3211)));
    outputs(1271) <= (layer0_outputs(2843)) or (layer0_outputs(3133));
    outputs(1272) <= not((layer0_outputs(1737)) and (layer0_outputs(4821)));
    outputs(1273) <= layer0_outputs(4662);
    outputs(1274) <= not(layer0_outputs(681));
    outputs(1275) <= not(layer0_outputs(2063));
    outputs(1276) <= (layer0_outputs(1303)) and not (layer0_outputs(4977));
    outputs(1277) <= layer0_outputs(555);
    outputs(1278) <= not(layer0_outputs(2643)) or (layer0_outputs(4627));
    outputs(1279) <= not((layer0_outputs(981)) and (layer0_outputs(1636)));
    outputs(1280) <= not(layer0_outputs(1665));
    outputs(1281) <= layer0_outputs(3418);
    outputs(1282) <= (layer0_outputs(1911)) and not (layer0_outputs(2383));
    outputs(1283) <= layer0_outputs(3172);
    outputs(1284) <= layer0_outputs(3379);
    outputs(1285) <= layer0_outputs(4604);
    outputs(1286) <= layer0_outputs(380);
    outputs(1287) <= not(layer0_outputs(215)) or (layer0_outputs(3574));
    outputs(1288) <= layer0_outputs(653);
    outputs(1289) <= not((layer0_outputs(4125)) and (layer0_outputs(161)));
    outputs(1290) <= (layer0_outputs(179)) and (layer0_outputs(826));
    outputs(1291) <= layer0_outputs(1311);
    outputs(1292) <= layer0_outputs(1394);
    outputs(1293) <= not(layer0_outputs(4460)) or (layer0_outputs(5097));
    outputs(1294) <= (layer0_outputs(1103)) xor (layer0_outputs(5032));
    outputs(1295) <= (layer0_outputs(1726)) and (layer0_outputs(881));
    outputs(1296) <= not(layer0_outputs(500));
    outputs(1297) <= layer0_outputs(3692);
    outputs(1298) <= not(layer0_outputs(822)) or (layer0_outputs(2094));
    outputs(1299) <= layer0_outputs(989);
    outputs(1300) <= (layer0_outputs(3748)) and (layer0_outputs(497));
    outputs(1301) <= (layer0_outputs(4889)) and not (layer0_outputs(163));
    outputs(1302) <= not(layer0_outputs(1345));
    outputs(1303) <= (layer0_outputs(3044)) xor (layer0_outputs(2139));
    outputs(1304) <= layer0_outputs(4384);
    outputs(1305) <= not(layer0_outputs(3912));
    outputs(1306) <= (layer0_outputs(728)) or (layer0_outputs(705));
    outputs(1307) <= layer0_outputs(192);
    outputs(1308) <= not(layer0_outputs(4655));
    outputs(1309) <= not(layer0_outputs(2754)) or (layer0_outputs(2839));
    outputs(1310) <= not(layer0_outputs(4841));
    outputs(1311) <= layer0_outputs(4692);
    outputs(1312) <= not((layer0_outputs(1098)) and (layer0_outputs(45)));
    outputs(1313) <= layer0_outputs(293);
    outputs(1314) <= not((layer0_outputs(303)) xor (layer0_outputs(875)));
    outputs(1315) <= not((layer0_outputs(1588)) xor (layer0_outputs(4526)));
    outputs(1316) <= (layer0_outputs(3654)) or (layer0_outputs(4028));
    outputs(1317) <= (layer0_outputs(1209)) or (layer0_outputs(4768));
    outputs(1318) <= (layer0_outputs(2179)) or (layer0_outputs(2524));
    outputs(1319) <= (layer0_outputs(4775)) and not (layer0_outputs(4344));
    outputs(1320) <= not(layer0_outputs(4122)) or (layer0_outputs(781));
    outputs(1321) <= not((layer0_outputs(4594)) and (layer0_outputs(1803)));
    outputs(1322) <= layer0_outputs(1330);
    outputs(1323) <= not(layer0_outputs(4158)) or (layer0_outputs(32));
    outputs(1324) <= layer0_outputs(4056);
    outputs(1325) <= layer0_outputs(4619);
    outputs(1326) <= not((layer0_outputs(4954)) and (layer0_outputs(396)));
    outputs(1327) <= not(layer0_outputs(1658));
    outputs(1328) <= layer0_outputs(1751);
    outputs(1329) <= not(layer0_outputs(5037));
    outputs(1330) <= not(layer0_outputs(4658));
    outputs(1331) <= layer0_outputs(3685);
    outputs(1332) <= layer0_outputs(2044);
    outputs(1333) <= not((layer0_outputs(4679)) xor (layer0_outputs(3525)));
    outputs(1334) <= not(layer0_outputs(1261));
    outputs(1335) <= not(layer0_outputs(1370)) or (layer0_outputs(478));
    outputs(1336) <= not((layer0_outputs(1433)) or (layer0_outputs(2263)));
    outputs(1337) <= not((layer0_outputs(420)) and (layer0_outputs(3561)));
    outputs(1338) <= layer0_outputs(2847);
    outputs(1339) <= not(layer0_outputs(3190)) or (layer0_outputs(1854));
    outputs(1340) <= (layer0_outputs(1576)) and (layer0_outputs(876));
    outputs(1341) <= (layer0_outputs(3070)) and (layer0_outputs(3396));
    outputs(1342) <= layer0_outputs(576);
    outputs(1343) <= not((layer0_outputs(2861)) and (layer0_outputs(3581)));
    outputs(1344) <= layer0_outputs(3237);
    outputs(1345) <= not(layer0_outputs(1060));
    outputs(1346) <= not(layer0_outputs(3996));
    outputs(1347) <= layer0_outputs(1467);
    outputs(1348) <= not(layer0_outputs(4678));
    outputs(1349) <= not(layer0_outputs(442));
    outputs(1350) <= not((layer0_outputs(3400)) or (layer0_outputs(2384)));
    outputs(1351) <= not(layer0_outputs(1996)) or (layer0_outputs(1818));
    outputs(1352) <= not(layer0_outputs(4944)) or (layer0_outputs(1971));
    outputs(1353) <= not((layer0_outputs(3112)) or (layer0_outputs(1879)));
    outputs(1354) <= layer0_outputs(2687);
    outputs(1355) <= not((layer0_outputs(553)) or (layer0_outputs(2259)));
    outputs(1356) <= (layer0_outputs(4386)) and (layer0_outputs(4384));
    outputs(1357) <= not((layer0_outputs(4336)) or (layer0_outputs(2323)));
    outputs(1358) <= layer0_outputs(4501);
    outputs(1359) <= layer0_outputs(4806);
    outputs(1360) <= layer0_outputs(4155);
    outputs(1361) <= layer0_outputs(2058);
    outputs(1362) <= layer0_outputs(4670);
    outputs(1363) <= layer0_outputs(1695);
    outputs(1364) <= not(layer0_outputs(1608));
    outputs(1365) <= not((layer0_outputs(3005)) or (layer0_outputs(4851)));
    outputs(1366) <= not((layer0_outputs(4236)) and (layer0_outputs(2421)));
    outputs(1367) <= (layer0_outputs(4385)) and not (layer0_outputs(74));
    outputs(1368) <= (layer0_outputs(3340)) and not (layer0_outputs(2564));
    outputs(1369) <= layer0_outputs(3517);
    outputs(1370) <= not(layer0_outputs(2661)) or (layer0_outputs(3827));
    outputs(1371) <= layer0_outputs(5004);
    outputs(1372) <= (layer0_outputs(263)) or (layer0_outputs(3566));
    outputs(1373) <= layer0_outputs(1231);
    outputs(1374) <= not(layer0_outputs(665)) or (layer0_outputs(3235));
    outputs(1375) <= (layer0_outputs(667)) xor (layer0_outputs(1878));
    outputs(1376) <= not(layer0_outputs(2781));
    outputs(1377) <= not(layer0_outputs(2403));
    outputs(1378) <= layer0_outputs(4590);
    outputs(1379) <= layer0_outputs(1934);
    outputs(1380) <= not(layer0_outputs(1180)) or (layer0_outputs(4461));
    outputs(1381) <= layer0_outputs(2360);
    outputs(1382) <= not((layer0_outputs(406)) xor (layer0_outputs(1667)));
    outputs(1383) <= layer0_outputs(1481);
    outputs(1384) <= not(layer0_outputs(4991));
    outputs(1385) <= (layer0_outputs(4569)) or (layer0_outputs(2032));
    outputs(1386) <= (layer0_outputs(3643)) or (layer0_outputs(1973));
    outputs(1387) <= (layer0_outputs(3397)) xor (layer0_outputs(4788));
    outputs(1388) <= not(layer0_outputs(3035));
    outputs(1389) <= not((layer0_outputs(3716)) and (layer0_outputs(3267)));
    outputs(1390) <= not(layer0_outputs(512));
    outputs(1391) <= layer0_outputs(2216);
    outputs(1392) <= (layer0_outputs(2742)) xor (layer0_outputs(4488));
    outputs(1393) <= not(layer0_outputs(80));
    outputs(1394) <= (layer0_outputs(4081)) and not (layer0_outputs(2096));
    outputs(1395) <= not((layer0_outputs(3128)) and (layer0_outputs(568)));
    outputs(1396) <= not(layer0_outputs(3644));
    outputs(1397) <= not(layer0_outputs(374)) or (layer0_outputs(3121));
    outputs(1398) <= not(layer0_outputs(4545));
    outputs(1399) <= (layer0_outputs(4550)) xor (layer0_outputs(1439));
    outputs(1400) <= not(layer0_outputs(2521)) or (layer0_outputs(310));
    outputs(1401) <= not((layer0_outputs(3302)) and (layer0_outputs(2506)));
    outputs(1402) <= not(layer0_outputs(2913)) or (layer0_outputs(2782));
    outputs(1403) <= not(layer0_outputs(4809)) or (layer0_outputs(3768));
    outputs(1404) <= not(layer0_outputs(1712));
    outputs(1405) <= not(layer0_outputs(2863));
    outputs(1406) <= layer0_outputs(3242);
    outputs(1407) <= (layer0_outputs(845)) xor (layer0_outputs(2738));
    outputs(1408) <= layer0_outputs(3134);
    outputs(1409) <= not(layer0_outputs(642));
    outputs(1410) <= not(layer0_outputs(2036));
    outputs(1411) <= (layer0_outputs(1547)) or (layer0_outputs(1798));
    outputs(1412) <= not(layer0_outputs(3910));
    outputs(1413) <= layer0_outputs(1966);
    outputs(1414) <= layer0_outputs(4636);
    outputs(1415) <= not(layer0_outputs(2988));
    outputs(1416) <= not((layer0_outputs(4423)) or (layer0_outputs(3372)));
    outputs(1417) <= (layer0_outputs(4555)) and (layer0_outputs(3275));
    outputs(1418) <= not((layer0_outputs(2599)) and (layer0_outputs(3317)));
    outputs(1419) <= not((layer0_outputs(1413)) or (layer0_outputs(2999)));
    outputs(1420) <= not(layer0_outputs(3354));
    outputs(1421) <= not(layer0_outputs(1493));
    outputs(1422) <= not(layer0_outputs(3794));
    outputs(1423) <= (layer0_outputs(1715)) or (layer0_outputs(5092));
    outputs(1424) <= (layer0_outputs(1440)) and (layer0_outputs(4170));
    outputs(1425) <= layer0_outputs(3169);
    outputs(1426) <= not(layer0_outputs(1813));
    outputs(1427) <= layer0_outputs(658);
    outputs(1428) <= layer0_outputs(2007);
    outputs(1429) <= not(layer0_outputs(4407));
    outputs(1430) <= not(layer0_outputs(1403)) or (layer0_outputs(3246));
    outputs(1431) <= (layer0_outputs(916)) and (layer0_outputs(2330));
    outputs(1432) <= not(layer0_outputs(1426)) or (layer0_outputs(2372));
    outputs(1433) <= not(layer0_outputs(3105));
    outputs(1434) <= not(layer0_outputs(4672));
    outputs(1435) <= layer0_outputs(3160);
    outputs(1436) <= not(layer0_outputs(88));
    outputs(1437) <= not(layer0_outputs(915));
    outputs(1438) <= not(layer0_outputs(4857));
    outputs(1439) <= not(layer0_outputs(3851));
    outputs(1440) <= not(layer0_outputs(3900)) or (layer0_outputs(3535));
    outputs(1441) <= layer0_outputs(1569);
    outputs(1442) <= layer0_outputs(2469);
    outputs(1443) <= (layer0_outputs(34)) or (layer0_outputs(456));
    outputs(1444) <= not(layer0_outputs(2750));
    outputs(1445) <= not(layer0_outputs(2575));
    outputs(1446) <= not(layer0_outputs(4802));
    outputs(1447) <= layer0_outputs(4710);
    outputs(1448) <= (layer0_outputs(4650)) and not (layer0_outputs(2877));
    outputs(1449) <= not(layer0_outputs(2629));
    outputs(1450) <= not((layer0_outputs(1458)) xor (layer0_outputs(3489)));
    outputs(1451) <= not(layer0_outputs(2308));
    outputs(1452) <= not(layer0_outputs(1665));
    outputs(1453) <= not((layer0_outputs(2079)) xor (layer0_outputs(490)));
    outputs(1454) <= layer0_outputs(334);
    outputs(1455) <= (layer0_outputs(1073)) and not (layer0_outputs(2874));
    outputs(1456) <= layer0_outputs(1146);
    outputs(1457) <= not((layer0_outputs(522)) and (layer0_outputs(4758)));
    outputs(1458) <= not(layer0_outputs(4286)) or (layer0_outputs(2522));
    outputs(1459) <= not(layer0_outputs(3384));
    outputs(1460) <= not((layer0_outputs(2504)) or (layer0_outputs(2060)));
    outputs(1461) <= (layer0_outputs(2166)) and (layer0_outputs(4518));
    outputs(1462) <= not((layer0_outputs(4050)) xor (layer0_outputs(3568)));
    outputs(1463) <= (layer0_outputs(1519)) and (layer0_outputs(1083));
    outputs(1464) <= layer0_outputs(2335);
    outputs(1465) <= not(layer0_outputs(4719));
    outputs(1466) <= layer0_outputs(4417);
    outputs(1467) <= not(layer0_outputs(4220));
    outputs(1468) <= not(layer0_outputs(44)) or (layer0_outputs(894));
    outputs(1469) <= (layer0_outputs(2688)) and not (layer0_outputs(4315));
    outputs(1470) <= layer0_outputs(952);
    outputs(1471) <= not((layer0_outputs(3346)) and (layer0_outputs(1092)));
    outputs(1472) <= not(layer0_outputs(309));
    outputs(1473) <= not(layer0_outputs(3899));
    outputs(1474) <= not(layer0_outputs(1256));
    outputs(1475) <= not(layer0_outputs(733));
    outputs(1476) <= layer0_outputs(4562);
    outputs(1477) <= not(layer0_outputs(2491)) or (layer0_outputs(1132));
    outputs(1478) <= layer0_outputs(4332);
    outputs(1479) <= not(layer0_outputs(2828)) or (layer0_outputs(3681));
    outputs(1480) <= not(layer0_outputs(1615));
    outputs(1481) <= not(layer0_outputs(4258));
    outputs(1482) <= not(layer0_outputs(2454));
    outputs(1483) <= not(layer0_outputs(4535));
    outputs(1484) <= not((layer0_outputs(135)) and (layer0_outputs(839)));
    outputs(1485) <= (layer0_outputs(3626)) and not (layer0_outputs(3972));
    outputs(1486) <= not((layer0_outputs(5064)) and (layer0_outputs(2193)));
    outputs(1487) <= not(layer0_outputs(1555));
    outputs(1488) <= not(layer0_outputs(4696)) or (layer0_outputs(1295));
    outputs(1489) <= not((layer0_outputs(2655)) and (layer0_outputs(4273)));
    outputs(1490) <= not(layer0_outputs(2695));
    outputs(1491) <= not(layer0_outputs(2086)) or (layer0_outputs(4522));
    outputs(1492) <= not(layer0_outputs(4183));
    outputs(1493) <= not(layer0_outputs(965)) or (layer0_outputs(3122));
    outputs(1494) <= layer0_outputs(2376);
    outputs(1495) <= layer0_outputs(4351);
    outputs(1496) <= (layer0_outputs(1997)) and not (layer0_outputs(43));
    outputs(1497) <= not(layer0_outputs(2743));
    outputs(1498) <= not((layer0_outputs(2439)) xor (layer0_outputs(563)));
    outputs(1499) <= layer0_outputs(3734);
    outputs(1500) <= layer0_outputs(5001);
    outputs(1501) <= not((layer0_outputs(2918)) and (layer0_outputs(2389)));
    outputs(1502) <= (layer0_outputs(2687)) and (layer0_outputs(3920));
    outputs(1503) <= (layer0_outputs(3705)) and not (layer0_outputs(667));
    outputs(1504) <= not(layer0_outputs(1104));
    outputs(1505) <= not(layer0_outputs(1606));
    outputs(1506) <= (layer0_outputs(4309)) and not (layer0_outputs(1605));
    outputs(1507) <= layer0_outputs(4414);
    outputs(1508) <= layer0_outputs(4810);
    outputs(1509) <= layer0_outputs(1701);
    outputs(1510) <= not((layer0_outputs(2347)) xor (layer0_outputs(4887)));
    outputs(1511) <= not((layer0_outputs(3075)) and (layer0_outputs(1534)));
    outputs(1512) <= not(layer0_outputs(4476));
    outputs(1513) <= not(layer0_outputs(4962));
    outputs(1514) <= not(layer0_outputs(2260));
    outputs(1515) <= layer0_outputs(4094);
    outputs(1516) <= not(layer0_outputs(3381));
    outputs(1517) <= not(layer0_outputs(1285)) or (layer0_outputs(864));
    outputs(1518) <= (layer0_outputs(459)) or (layer0_outputs(1223));
    outputs(1519) <= layer0_outputs(1720);
    outputs(1520) <= not((layer0_outputs(3080)) xor (layer0_outputs(4600)));
    outputs(1521) <= not((layer0_outputs(1254)) xor (layer0_outputs(3320)));
    outputs(1522) <= (layer0_outputs(1558)) and (layer0_outputs(1501));
    outputs(1523) <= not(layer0_outputs(1095));
    outputs(1524) <= layer0_outputs(4260);
    outputs(1525) <= layer0_outputs(4646);
    outputs(1526) <= not(layer0_outputs(3389));
    outputs(1527) <= layer0_outputs(4192);
    outputs(1528) <= layer0_outputs(2309);
    outputs(1529) <= layer0_outputs(2740);
    outputs(1530) <= not((layer0_outputs(3029)) and (layer0_outputs(3659)));
    outputs(1531) <= layer0_outputs(4915);
    outputs(1532) <= not(layer0_outputs(140));
    outputs(1533) <= not(layer0_outputs(4572)) or (layer0_outputs(2372));
    outputs(1534) <= (layer0_outputs(4194)) or (layer0_outputs(2290));
    outputs(1535) <= not(layer0_outputs(1568));
    outputs(1536) <= layer0_outputs(4300);
    outputs(1537) <= layer0_outputs(4211);
    outputs(1538) <= (layer0_outputs(4355)) and (layer0_outputs(2170));
    outputs(1539) <= not(layer0_outputs(4912));
    outputs(1540) <= layer0_outputs(4263);
    outputs(1541) <= (layer0_outputs(2629)) xor (layer0_outputs(3580));
    outputs(1542) <= not(layer0_outputs(1221));
    outputs(1543) <= not((layer0_outputs(4689)) xor (layer0_outputs(2923)));
    outputs(1544) <= (layer0_outputs(329)) and (layer0_outputs(4117));
    outputs(1545) <= not(layer0_outputs(2071));
    outputs(1546) <= not(layer0_outputs(4200));
    outputs(1547) <= layer0_outputs(3726);
    outputs(1548) <= (layer0_outputs(2472)) and not (layer0_outputs(4836));
    outputs(1549) <= layer0_outputs(865);
    outputs(1550) <= not(layer0_outputs(3932));
    outputs(1551) <= layer0_outputs(3216);
    outputs(1552) <= not((layer0_outputs(3880)) and (layer0_outputs(1676)));
    outputs(1553) <= (layer0_outputs(2271)) and (layer0_outputs(1324));
    outputs(1554) <= (layer0_outputs(393)) and (layer0_outputs(3509));
    outputs(1555) <= (layer0_outputs(3196)) and not (layer0_outputs(4592));
    outputs(1556) <= (layer0_outputs(4939)) xor (layer0_outputs(3813));
    outputs(1557) <= (layer0_outputs(2364)) and not (layer0_outputs(1002));
    outputs(1558) <= not(layer0_outputs(279)) or (layer0_outputs(3947));
    outputs(1559) <= (layer0_outputs(5007)) xor (layer0_outputs(2419));
    outputs(1560) <= not((layer0_outputs(1457)) xor (layer0_outputs(3646)));
    outputs(1561) <= layer0_outputs(4568);
    outputs(1562) <= not(layer0_outputs(1026));
    outputs(1563) <= (layer0_outputs(2698)) or (layer0_outputs(3850));
    outputs(1564) <= layer0_outputs(2717);
    outputs(1565) <= not(layer0_outputs(4957)) or (layer0_outputs(3728));
    outputs(1566) <= not(layer0_outputs(1843));
    outputs(1567) <= layer0_outputs(2817);
    outputs(1568) <= layer0_outputs(2420);
    outputs(1569) <= (layer0_outputs(3062)) and (layer0_outputs(4049));
    outputs(1570) <= (layer0_outputs(1382)) xor (layer0_outputs(1732));
    outputs(1571) <= not((layer0_outputs(4486)) or (layer0_outputs(2168)));
    outputs(1572) <= (layer0_outputs(4810)) and not (layer0_outputs(4485));
    outputs(1573) <= not(layer0_outputs(827)) or (layer0_outputs(3322));
    outputs(1574) <= (layer0_outputs(387)) and (layer0_outputs(2514));
    outputs(1575) <= not(layer0_outputs(4886));
    outputs(1576) <= not(layer0_outputs(4294));
    outputs(1577) <= layer0_outputs(4704);
    outputs(1578) <= layer0_outputs(804);
    outputs(1579) <= layer0_outputs(55);
    outputs(1580) <= not(layer0_outputs(2916));
    outputs(1581) <= not(layer0_outputs(4608));
    outputs(1582) <= not((layer0_outputs(3370)) xor (layer0_outputs(389)));
    outputs(1583) <= not((layer0_outputs(2137)) xor (layer0_outputs(2882)));
    outputs(1584) <= (layer0_outputs(4579)) xor (layer0_outputs(3956));
    outputs(1585) <= not((layer0_outputs(23)) and (layer0_outputs(1750)));
    outputs(1586) <= not(layer0_outputs(2963)) or (layer0_outputs(3455));
    outputs(1587) <= (layer0_outputs(4208)) and not (layer0_outputs(3114));
    outputs(1588) <= layer0_outputs(2075);
    outputs(1589) <= not((layer0_outputs(506)) or (layer0_outputs(4062)));
    outputs(1590) <= (layer0_outputs(979)) and not (layer0_outputs(1603));
    outputs(1591) <= not(layer0_outputs(4132));
    outputs(1592) <= not((layer0_outputs(4880)) xor (layer0_outputs(4960)));
    outputs(1593) <= (layer0_outputs(4098)) xor (layer0_outputs(3868));
    outputs(1594) <= not(layer0_outputs(3632));
    outputs(1595) <= layer0_outputs(4452);
    outputs(1596) <= not((layer0_outputs(3203)) or (layer0_outputs(3092)));
    outputs(1597) <= (layer0_outputs(2178)) xor (layer0_outputs(246));
    outputs(1598) <= layer0_outputs(1364);
    outputs(1599) <= layer0_outputs(4473);
    outputs(1600) <= not(layer0_outputs(1523));
    outputs(1601) <= not(layer0_outputs(4716));
    outputs(1602) <= not((layer0_outputs(4324)) xor (layer0_outputs(18)));
    outputs(1603) <= not(layer0_outputs(1923));
    outputs(1604) <= (layer0_outputs(1767)) xor (layer0_outputs(33));
    outputs(1605) <= layer0_outputs(746);
    outputs(1606) <= not(layer0_outputs(1365));
    outputs(1607) <= (layer0_outputs(1862)) and not (layer0_outputs(1323));
    outputs(1608) <= not(layer0_outputs(4429));
    outputs(1609) <= (layer0_outputs(5027)) and not (layer0_outputs(1039));
    outputs(1610) <= (layer0_outputs(1326)) xor (layer0_outputs(4698));
    outputs(1611) <= layer0_outputs(5099);
    outputs(1612) <= not(layer0_outputs(2916));
    outputs(1613) <= (layer0_outputs(4525)) and not (layer0_outputs(4963));
    outputs(1614) <= (layer0_outputs(4980)) and not (layer0_outputs(3042));
    outputs(1615) <= not(layer0_outputs(10));
    outputs(1616) <= not(layer0_outputs(1930));
    outputs(1617) <= (layer0_outputs(1030)) and not (layer0_outputs(4318));
    outputs(1618) <= not(layer0_outputs(802));
    outputs(1619) <= not(layer0_outputs(1856));
    outputs(1620) <= not(layer0_outputs(1191));
    outputs(1621) <= not(layer0_outputs(1458));
    outputs(1622) <= not(layer0_outputs(4118));
    outputs(1623) <= (layer0_outputs(4418)) xor (layer0_outputs(3756));
    outputs(1624) <= not(layer0_outputs(435));
    outputs(1625) <= not((layer0_outputs(2794)) xor (layer0_outputs(3534)));
    outputs(1626) <= layer0_outputs(813);
    outputs(1627) <= layer0_outputs(1063);
    outputs(1628) <= not(layer0_outputs(1912));
    outputs(1629) <= not(layer0_outputs(721));
    outputs(1630) <= layer0_outputs(1833);
    outputs(1631) <= layer0_outputs(4072);
    outputs(1632) <= not(layer0_outputs(3501));
    outputs(1633) <= not((layer0_outputs(3356)) or (layer0_outputs(2683)));
    outputs(1634) <= (layer0_outputs(4771)) and (layer0_outputs(3948));
    outputs(1635) <= not(layer0_outputs(723)) or (layer0_outputs(673));
    outputs(1636) <= not(layer0_outputs(797));
    outputs(1637) <= (layer0_outputs(4634)) xor (layer0_outputs(2967));
    outputs(1638) <= not(layer0_outputs(4449));
    outputs(1639) <= (layer0_outputs(4076)) xor (layer0_outputs(4553));
    outputs(1640) <= not(layer0_outputs(3398));
    outputs(1641) <= layer0_outputs(921);
    outputs(1642) <= layer0_outputs(1485);
    outputs(1643) <= layer0_outputs(1049);
    outputs(1644) <= not((layer0_outputs(1240)) or (layer0_outputs(1319)));
    outputs(1645) <= not(layer0_outputs(1447));
    outputs(1646) <= not(layer0_outputs(3120));
    outputs(1647) <= not(layer0_outputs(3578));
    outputs(1648) <= (layer0_outputs(4923)) and not (layer0_outputs(3127));
    outputs(1649) <= not(layer0_outputs(2778));
    outputs(1650) <= not(layer0_outputs(4240));
    outputs(1651) <= layer0_outputs(862);
    outputs(1652) <= layer0_outputs(65);
    outputs(1653) <= layer0_outputs(3772);
    outputs(1654) <= (layer0_outputs(1015)) and not (layer0_outputs(3072));
    outputs(1655) <= layer0_outputs(3818);
    outputs(1656) <= not(layer0_outputs(3801));
    outputs(1657) <= not(layer0_outputs(1253));
    outputs(1658) <= (layer0_outputs(4191)) and not (layer0_outputs(3978));
    outputs(1659) <= layer0_outputs(5000);
    outputs(1660) <= not(layer0_outputs(1143));
    outputs(1661) <= not((layer0_outputs(339)) or (layer0_outputs(2343)));
    outputs(1662) <= not(layer0_outputs(3051));
    outputs(1663) <= (layer0_outputs(2956)) and not (layer0_outputs(4285));
    outputs(1664) <= not(layer0_outputs(926)) or (layer0_outputs(3977));
    outputs(1665) <= not(layer0_outputs(3189)) or (layer0_outputs(1979));
    outputs(1666) <= (layer0_outputs(1377)) xor (layer0_outputs(4092));
    outputs(1667) <= layer0_outputs(4558);
    outputs(1668) <= (layer0_outputs(3712)) or (layer0_outputs(178));
    outputs(1669) <= (layer0_outputs(196)) and not (layer0_outputs(1264));
    outputs(1670) <= layer0_outputs(3559);
    outputs(1671) <= (layer0_outputs(3422)) and not (layer0_outputs(4507));
    outputs(1672) <= layer0_outputs(1785);
    outputs(1673) <= not(layer0_outputs(1410)) or (layer0_outputs(2964));
    outputs(1674) <= not((layer0_outputs(4000)) xor (layer0_outputs(1497)));
    outputs(1675) <= (layer0_outputs(2137)) and (layer0_outputs(2780));
    outputs(1676) <= (layer0_outputs(748)) and not (layer0_outputs(2002));
    outputs(1677) <= (layer0_outputs(1842)) xor (layer0_outputs(1118));
    outputs(1678) <= (layer0_outputs(3959)) xor (layer0_outputs(2696));
    outputs(1679) <= layer0_outputs(1924);
    outputs(1680) <= not(layer0_outputs(419));
    outputs(1681) <= layer0_outputs(2859);
    outputs(1682) <= layer0_outputs(122);
    outputs(1683) <= layer0_outputs(3124);
    outputs(1684) <= layer0_outputs(1218);
    outputs(1685) <= not(layer0_outputs(4726)) or (layer0_outputs(2929));
    outputs(1686) <= not(layer0_outputs(4519));
    outputs(1687) <= (layer0_outputs(1599)) and not (layer0_outputs(589));
    outputs(1688) <= (layer0_outputs(3177)) xor (layer0_outputs(2153));
    outputs(1689) <= not(layer0_outputs(2060));
    outputs(1690) <= layer0_outputs(833);
    outputs(1691) <= not((layer0_outputs(773)) and (layer0_outputs(3971)));
    outputs(1692) <= layer0_outputs(84);
    outputs(1693) <= not(layer0_outputs(2835));
    outputs(1694) <= not(layer0_outputs(4483));
    outputs(1695) <= layer0_outputs(2141);
    outputs(1696) <= (layer0_outputs(2435)) xor (layer0_outputs(4653));
    outputs(1697) <= not((layer0_outputs(4888)) xor (layer0_outputs(5041)));
    outputs(1698) <= not(layer0_outputs(4907));
    outputs(1699) <= not(layer0_outputs(2892));
    outputs(1700) <= not((layer0_outputs(1570)) xor (layer0_outputs(1228)));
    outputs(1701) <= (layer0_outputs(2791)) and not (layer0_outputs(382));
    outputs(1702) <= layer0_outputs(2284);
    outputs(1703) <= not((layer0_outputs(976)) xor (layer0_outputs(5059)));
    outputs(1704) <= (layer0_outputs(500)) and not (layer0_outputs(2031));
    outputs(1705) <= layer0_outputs(1476);
    outputs(1706) <= not(layer0_outputs(4465));
    outputs(1707) <= (layer0_outputs(4856)) and (layer0_outputs(157));
    outputs(1708) <= (layer0_outputs(87)) xor (layer0_outputs(2023));
    outputs(1709) <= not((layer0_outputs(4453)) xor (layer0_outputs(1095)));
    outputs(1710) <= not(layer0_outputs(2168));
    outputs(1711) <= layer0_outputs(176);
    outputs(1712) <= (layer0_outputs(630)) and not (layer0_outputs(4754));
    outputs(1713) <= layer0_outputs(3188);
    outputs(1714) <= (layer0_outputs(45)) and (layer0_outputs(3262));
    outputs(1715) <= (layer0_outputs(1233)) xor (layer0_outputs(2037));
    outputs(1716) <= not(layer0_outputs(5015));
    outputs(1717) <= layer0_outputs(1498);
    outputs(1718) <= not(layer0_outputs(4804));
    outputs(1719) <= (layer0_outputs(4640)) or (layer0_outputs(595));
    outputs(1720) <= layer0_outputs(4766);
    outputs(1721) <= (layer0_outputs(4626)) xor (layer0_outputs(472));
    outputs(1722) <= (layer0_outputs(1015)) and (layer0_outputs(2842));
    outputs(1723) <= layer0_outputs(4176);
    outputs(1724) <= not(layer0_outputs(4635));
    outputs(1725) <= (layer0_outputs(4555)) and (layer0_outputs(916));
    outputs(1726) <= not(layer0_outputs(4862));
    outputs(1727) <= (layer0_outputs(1663)) and (layer0_outputs(1766));
    outputs(1728) <= layer0_outputs(1427);
    outputs(1729) <= not(layer0_outputs(548));
    outputs(1730) <= layer0_outputs(25);
    outputs(1731) <= layer0_outputs(71);
    outputs(1732) <= not(layer0_outputs(1792));
    outputs(1733) <= not(layer0_outputs(2004));
    outputs(1734) <= layer0_outputs(4102);
    outputs(1735) <= not((layer0_outputs(4720)) or (layer0_outputs(4371)));
    outputs(1736) <= not((layer0_outputs(2675)) or (layer0_outputs(1119)));
    outputs(1737) <= layer0_outputs(3155);
    outputs(1738) <= (layer0_outputs(4515)) and not (layer0_outputs(2611));
    outputs(1739) <= not((layer0_outputs(859)) xor (layer0_outputs(655)));
    outputs(1740) <= (layer0_outputs(972)) and not (layer0_outputs(4272));
    outputs(1741) <= (layer0_outputs(4946)) and not (layer0_outputs(1717));
    outputs(1742) <= not(layer0_outputs(1660));
    outputs(1743) <= not(layer0_outputs(1662));
    outputs(1744) <= layer0_outputs(3284);
    outputs(1745) <= not(layer0_outputs(2314));
    outputs(1746) <= (layer0_outputs(4827)) and not (layer0_outputs(5115));
    outputs(1747) <= not((layer0_outputs(4796)) or (layer0_outputs(5)));
    outputs(1748) <= layer0_outputs(1054);
    outputs(1749) <= (layer0_outputs(3430)) xor (layer0_outputs(2322));
    outputs(1750) <= (layer0_outputs(762)) or (layer0_outputs(3535));
    outputs(1751) <= (layer0_outputs(4295)) and (layer0_outputs(673));
    outputs(1752) <= not((layer0_outputs(99)) or (layer0_outputs(581)));
    outputs(1753) <= (layer0_outputs(2785)) and not (layer0_outputs(1407));
    outputs(1754) <= not(layer0_outputs(3604));
    outputs(1755) <= layer0_outputs(1150);
    outputs(1756) <= layer0_outputs(1546);
    outputs(1757) <= not(layer0_outputs(2274));
    outputs(1758) <= layer0_outputs(4557);
    outputs(1759) <= not((layer0_outputs(2436)) and (layer0_outputs(1286)));
    outputs(1760) <= not(layer0_outputs(3684));
    outputs(1761) <= not(layer0_outputs(1622));
    outputs(1762) <= not((layer0_outputs(9)) xor (layer0_outputs(2743)));
    outputs(1763) <= layer0_outputs(3953);
    outputs(1764) <= layer0_outputs(4078);
    outputs(1765) <= (layer0_outputs(2233)) and not (layer0_outputs(1853));
    outputs(1766) <= not(layer0_outputs(4542));
    outputs(1767) <= not(layer0_outputs(1109));
    outputs(1768) <= not(layer0_outputs(3476));
    outputs(1769) <= not((layer0_outputs(4976)) xor (layer0_outputs(4601)));
    outputs(1770) <= not(layer0_outputs(2818));
    outputs(1771) <= not(layer0_outputs(2980));
    outputs(1772) <= not((layer0_outputs(2139)) xor (layer0_outputs(1799)));
    outputs(1773) <= not(layer0_outputs(1593));
    outputs(1774) <= not(layer0_outputs(220));
    outputs(1775) <= not((layer0_outputs(3938)) or (layer0_outputs(1215)));
    outputs(1776) <= not(layer0_outputs(1379));
    outputs(1777) <= layer0_outputs(3406);
    outputs(1778) <= layer0_outputs(3770);
    outputs(1779) <= not(layer0_outputs(3943));
    outputs(1780) <= not(layer0_outputs(1597)) or (layer0_outputs(2385));
    outputs(1781) <= not(layer0_outputs(4817)) or (layer0_outputs(4831));
    outputs(1782) <= (layer0_outputs(3572)) and (layer0_outputs(3431));
    outputs(1783) <= not(layer0_outputs(3335));
    outputs(1784) <= not(layer0_outputs(1817));
    outputs(1785) <= not(layer0_outputs(4400));
    outputs(1786) <= (layer0_outputs(1637)) and not (layer0_outputs(859));
    outputs(1787) <= layer0_outputs(816);
    outputs(1788) <= layer0_outputs(3482);
    outputs(1789) <= (layer0_outputs(2082)) and not (layer0_outputs(4564));
    outputs(1790) <= layer0_outputs(5026);
    outputs(1791) <= layer0_outputs(423);
    outputs(1792) <= not(layer0_outputs(4164));
    outputs(1793) <= not(layer0_outputs(1757));
    outputs(1794) <= not(layer0_outputs(2941));
    outputs(1795) <= not((layer0_outputs(4559)) xor (layer0_outputs(968)));
    outputs(1796) <= (layer0_outputs(1549)) and not (layer0_outputs(3339));
    outputs(1797) <= not(layer0_outputs(1133));
    outputs(1798) <= layer0_outputs(1082);
    outputs(1799) <= not((layer0_outputs(4690)) xor (layer0_outputs(4456)));
    outputs(1800) <= not(layer0_outputs(1215));
    outputs(1801) <= (layer0_outputs(2887)) and not (layer0_outputs(685));
    outputs(1802) <= layer0_outputs(4412);
    outputs(1803) <= layer0_outputs(552);
    outputs(1804) <= not(layer0_outputs(1087));
    outputs(1805) <= not((layer0_outputs(3517)) xor (layer0_outputs(4454)));
    outputs(1806) <= (layer0_outputs(1837)) and not (layer0_outputs(363));
    outputs(1807) <= (layer0_outputs(3731)) and (layer0_outputs(1559));
    outputs(1808) <= (layer0_outputs(2732)) and not (layer0_outputs(5010));
    outputs(1809) <= not((layer0_outputs(5017)) or (layer0_outputs(4556)));
    outputs(1810) <= not(layer0_outputs(4103));
    outputs(1811) <= (layer0_outputs(4044)) and (layer0_outputs(5113));
    outputs(1812) <= layer0_outputs(4841);
    outputs(1813) <= not(layer0_outputs(1730));
    outputs(1814) <= layer0_outputs(3933);
    outputs(1815) <= not((layer0_outputs(4917)) or (layer0_outputs(776)));
    outputs(1816) <= not(layer0_outputs(2250));
    outputs(1817) <= not(layer0_outputs(642));
    outputs(1818) <= (layer0_outputs(1705)) and not (layer0_outputs(4510));
    outputs(1819) <= not(layer0_outputs(3612));
    outputs(1820) <= layer0_outputs(1356);
    outputs(1821) <= layer0_outputs(1491);
    outputs(1822) <= layer0_outputs(2045);
    outputs(1823) <= (layer0_outputs(320)) xor (layer0_outputs(657));
    outputs(1824) <= not((layer0_outputs(2917)) or (layer0_outputs(3055)));
    outputs(1825) <= layer0_outputs(4523);
    outputs(1826) <= not(layer0_outputs(136));
    outputs(1827) <= layer0_outputs(2985);
    outputs(1828) <= (layer0_outputs(4302)) and not (layer0_outputs(3858));
    outputs(1829) <= not(layer0_outputs(1660));
    outputs(1830) <= layer0_outputs(3742);
    outputs(1831) <= (layer0_outputs(3528)) xor (layer0_outputs(4424));
    outputs(1832) <= not(layer0_outputs(4039));
    outputs(1833) <= not((layer0_outputs(1747)) and (layer0_outputs(418)));
    outputs(1834) <= layer0_outputs(2353);
    outputs(1835) <= not(layer0_outputs(4542));
    outputs(1836) <= (layer0_outputs(2512)) and not (layer0_outputs(4187));
    outputs(1837) <= layer0_outputs(4910);
    outputs(1838) <= not(layer0_outputs(3974));
    outputs(1839) <= (layer0_outputs(939)) and not (layer0_outputs(4012));
    outputs(1840) <= not(layer0_outputs(952));
    outputs(1841) <= not(layer0_outputs(3888));
    outputs(1842) <= not((layer0_outputs(1501)) xor (layer0_outputs(3855)));
    outputs(1843) <= layer0_outputs(4188);
    outputs(1844) <= not(layer0_outputs(2217));
    outputs(1845) <= not(layer0_outputs(1190));
    outputs(1846) <= layer0_outputs(2484);
    outputs(1847) <= layer0_outputs(111);
    outputs(1848) <= not(layer0_outputs(4595));
    outputs(1849) <= (layer0_outputs(3066)) and (layer0_outputs(747));
    outputs(1850) <= layer0_outputs(945);
    outputs(1851) <= not(layer0_outputs(2296));
    outputs(1852) <= layer0_outputs(4290);
    outputs(1853) <= (layer0_outputs(2856)) or (layer0_outputs(2882));
    outputs(1854) <= not(layer0_outputs(3551));
    outputs(1855) <= not((layer0_outputs(4770)) xor (layer0_outputs(4104)));
    outputs(1856) <= layer0_outputs(4218);
    outputs(1857) <= layer0_outputs(792);
    outputs(1858) <= not(layer0_outputs(1812)) or (layer0_outputs(4218));
    outputs(1859) <= not(layer0_outputs(1461));
    outputs(1860) <= not(layer0_outputs(5115));
    outputs(1861) <= (layer0_outputs(560)) or (layer0_outputs(1097));
    outputs(1862) <= layer0_outputs(703);
    outputs(1863) <= layer0_outputs(2584);
    outputs(1864) <= not((layer0_outputs(1895)) or (layer0_outputs(2987)));
    outputs(1865) <= not(layer0_outputs(917));
    outputs(1866) <= (layer0_outputs(4021)) and not (layer0_outputs(2294));
    outputs(1867) <= not(layer0_outputs(2749));
    outputs(1868) <= (layer0_outputs(3207)) and not (layer0_outputs(1484));
    outputs(1869) <= layer0_outputs(3067);
    outputs(1870) <= layer0_outputs(4995);
    outputs(1871) <= layer0_outputs(3844);
    outputs(1872) <= not((layer0_outputs(3109)) xor (layer0_outputs(4118)));
    outputs(1873) <= not(layer0_outputs(648));
    outputs(1874) <= not(layer0_outputs(1004));
    outputs(1875) <= (layer0_outputs(3780)) and not (layer0_outputs(1106));
    outputs(1876) <= layer0_outputs(2324);
    outputs(1877) <= layer0_outputs(1035);
    outputs(1878) <= layer0_outputs(1545);
    outputs(1879) <= not((layer0_outputs(4731)) xor (layer0_outputs(1801)));
    outputs(1880) <= (layer0_outputs(3068)) xor (layer0_outputs(3377));
    outputs(1881) <= layer0_outputs(3588);
    outputs(1882) <= layer0_outputs(2802);
    outputs(1883) <= layer0_outputs(1858);
    outputs(1884) <= (layer0_outputs(4153)) and not (layer0_outputs(1849));
    outputs(1885) <= not((layer0_outputs(168)) or (layer0_outputs(4537)));
    outputs(1886) <= layer0_outputs(992);
    outputs(1887) <= not(layer0_outputs(5118));
    outputs(1888) <= (layer0_outputs(2360)) and not (layer0_outputs(3532));
    outputs(1889) <= layer0_outputs(4914);
    outputs(1890) <= layer0_outputs(4203);
    outputs(1891) <= not(layer0_outputs(2380));
    outputs(1892) <= layer0_outputs(2754);
    outputs(1893) <= not(layer0_outputs(1706));
    outputs(1894) <= layer0_outputs(107);
    outputs(1895) <= (layer0_outputs(701)) and (layer0_outputs(1776));
    outputs(1896) <= layer0_outputs(1775);
    outputs(1897) <= layer0_outputs(426);
    outputs(1898) <= layer0_outputs(3926);
    outputs(1899) <= (layer0_outputs(3861)) and not (layer0_outputs(5013));
    outputs(1900) <= (layer0_outputs(1025)) and not (layer0_outputs(4710));
    outputs(1901) <= (layer0_outputs(4017)) and (layer0_outputs(3646));
    outputs(1902) <= not(layer0_outputs(1524));
    outputs(1903) <= not(layer0_outputs(769));
    outputs(1904) <= (layer0_outputs(4188)) xor (layer0_outputs(4202));
    outputs(1905) <= not((layer0_outputs(2567)) xor (layer0_outputs(3039)));
    outputs(1906) <= not((layer0_outputs(704)) or (layer0_outputs(1354)));
    outputs(1907) <= not((layer0_outputs(4244)) xor (layer0_outputs(2968)));
    outputs(1908) <= not((layer0_outputs(3584)) or (layer0_outputs(282)));
    outputs(1909) <= layer0_outputs(2899);
    outputs(1910) <= layer0_outputs(189);
    outputs(1911) <= not((layer0_outputs(1960)) xor (layer0_outputs(4283)));
    outputs(1912) <= (layer0_outputs(4972)) xor (layer0_outputs(2852));
    outputs(1913) <= not((layer0_outputs(223)) xor (layer0_outputs(1087)));
    outputs(1914) <= layer0_outputs(1702);
    outputs(1915) <= not(layer0_outputs(4035));
    outputs(1916) <= layer0_outputs(4805);
    outputs(1917) <= not((layer0_outputs(4316)) or (layer0_outputs(3696)));
    outputs(1918) <= not(layer0_outputs(4053)) or (layer0_outputs(2648));
    outputs(1919) <= not(layer0_outputs(227));
    outputs(1920) <= (layer0_outputs(4827)) and (layer0_outputs(571));
    outputs(1921) <= layer0_outputs(1178);
    outputs(1922) <= not(layer0_outputs(2490));
    outputs(1923) <= layer0_outputs(3140);
    outputs(1924) <= (layer0_outputs(1989)) and not (layer0_outputs(275));
    outputs(1925) <= layer0_outputs(2379);
    outputs(1926) <= (layer0_outputs(1770)) and (layer0_outputs(4940));
    outputs(1927) <= layer0_outputs(4949);
    outputs(1928) <= layer0_outputs(697);
    outputs(1929) <= layer0_outputs(4492);
    outputs(1930) <= layer0_outputs(3138);
    outputs(1931) <= not(layer0_outputs(2190));
    outputs(1932) <= not(layer0_outputs(1526)) or (layer0_outputs(3350));
    outputs(1933) <= (layer0_outputs(1640)) xor (layer0_outputs(300));
    outputs(1934) <= layer0_outputs(4363);
    outputs(1935) <= layer0_outputs(3440);
    outputs(1936) <= (layer0_outputs(3644)) xor (layer0_outputs(2140));
    outputs(1937) <= layer0_outputs(3322);
    outputs(1938) <= layer0_outputs(901);
    outputs(1939) <= (layer0_outputs(286)) and (layer0_outputs(322));
    outputs(1940) <= layer0_outputs(4941);
    outputs(1941) <= layer0_outputs(2181);
    outputs(1942) <= layer0_outputs(2073);
    outputs(1943) <= (layer0_outputs(1693)) xor (layer0_outputs(734));
    outputs(1944) <= not(layer0_outputs(4316));
    outputs(1945) <= not((layer0_outputs(1380)) xor (layer0_outputs(3672)));
    outputs(1946) <= not((layer0_outputs(4869)) or (layer0_outputs(5078)));
    outputs(1947) <= not((layer0_outputs(4013)) or (layer0_outputs(2503)));
    outputs(1948) <= layer0_outputs(3939);
    outputs(1949) <= not(layer0_outputs(4575));
    outputs(1950) <= not(layer0_outputs(7));
    outputs(1951) <= not(layer0_outputs(418));
    outputs(1952) <= (layer0_outputs(1944)) and not (layer0_outputs(4935));
    outputs(1953) <= (layer0_outputs(2930)) and not (layer0_outputs(2756));
    outputs(1954) <= layer0_outputs(1594);
    outputs(1955) <= not((layer0_outputs(4958)) or (layer0_outputs(4951)));
    outputs(1956) <= (layer0_outputs(405)) and not (layer0_outputs(4027));
    outputs(1957) <= not(layer0_outputs(1930));
    outputs(1958) <= (layer0_outputs(3284)) and not (layer0_outputs(1068));
    outputs(1959) <= not(layer0_outputs(2070)) or (layer0_outputs(369));
    outputs(1960) <= (layer0_outputs(4389)) and (layer0_outputs(4832));
    outputs(1961) <= layer0_outputs(3140);
    outputs(1962) <= not(layer0_outputs(4449));
    outputs(1963) <= layer0_outputs(656);
    outputs(1964) <= not((layer0_outputs(2118)) xor (layer0_outputs(2061)));
    outputs(1965) <= not(layer0_outputs(621));
    outputs(1966) <= not(layer0_outputs(4031));
    outputs(1967) <= (layer0_outputs(1142)) and not (layer0_outputs(276));
    outputs(1968) <= layer0_outputs(3277);
    outputs(1969) <= (layer0_outputs(3448)) and (layer0_outputs(680));
    outputs(1970) <= (layer0_outputs(1283)) and not (layer0_outputs(442));
    outputs(1971) <= not(layer0_outputs(1006));
    outputs(1972) <= layer0_outputs(975);
    outputs(1973) <= layer0_outputs(280);
    outputs(1974) <= not(layer0_outputs(840));
    outputs(1975) <= (layer0_outputs(1857)) and not (layer0_outputs(3507));
    outputs(1976) <= not(layer0_outputs(1562));
    outputs(1977) <= (layer0_outputs(1782)) and not (layer0_outputs(2326));
    outputs(1978) <= (layer0_outputs(4636)) and not (layer0_outputs(4040));
    outputs(1979) <= layer0_outputs(3714);
    outputs(1980) <= layer0_outputs(2702);
    outputs(1981) <= layer0_outputs(4223);
    outputs(1982) <= (layer0_outputs(2857)) and (layer0_outputs(4173));
    outputs(1983) <= not(layer0_outputs(3417));
    outputs(1984) <= (layer0_outputs(2131)) and not (layer0_outputs(4705));
    outputs(1985) <= layer0_outputs(4848);
    outputs(1986) <= not(layer0_outputs(4814));
    outputs(1987) <= not((layer0_outputs(3450)) xor (layer0_outputs(1357)));
    outputs(1988) <= layer0_outputs(2441);
    outputs(1989) <= not((layer0_outputs(3960)) or (layer0_outputs(3862)));
    outputs(1990) <= (layer0_outputs(888)) and (layer0_outputs(294));
    outputs(1991) <= layer0_outputs(1999);
    outputs(1992) <= (layer0_outputs(2224)) or (layer0_outputs(1952));
    outputs(1993) <= (layer0_outputs(4244)) or (layer0_outputs(1314));
    outputs(1994) <= layer0_outputs(4965);
    outputs(1995) <= not((layer0_outputs(4898)) xor (layer0_outputs(1279)));
    outputs(1996) <= (layer0_outputs(210)) and not (layer0_outputs(3531));
    outputs(1997) <= layer0_outputs(1713);
    outputs(1998) <= (layer0_outputs(3135)) and not (layer0_outputs(1));
    outputs(1999) <= layer0_outputs(2339);
    outputs(2000) <= not((layer0_outputs(2127)) and (layer0_outputs(4345)));
    outputs(2001) <= layer0_outputs(4011);
    outputs(2002) <= not((layer0_outputs(3636)) xor (layer0_outputs(3310)));
    outputs(2003) <= (layer0_outputs(4659)) xor (layer0_outputs(3009));
    outputs(2004) <= layer0_outputs(4110);
    outputs(2005) <= not(layer0_outputs(1475));
    outputs(2006) <= not(layer0_outputs(1864));
    outputs(2007) <= not(layer0_outputs(3070));
    outputs(2008) <= not((layer0_outputs(3778)) and (layer0_outputs(2158)));
    outputs(2009) <= not(layer0_outputs(4424)) or (layer0_outputs(987));
    outputs(2010) <= layer0_outputs(1156);
    outputs(2011) <= layer0_outputs(3212);
    outputs(2012) <= (layer0_outputs(4818)) xor (layer0_outputs(447));
    outputs(2013) <= not(layer0_outputs(2103)) or (layer0_outputs(2033));
    outputs(2014) <= layer0_outputs(3470);
    outputs(2015) <= layer0_outputs(1965);
    outputs(2016) <= layer0_outputs(3086);
    outputs(2017) <= not(layer0_outputs(1653));
    outputs(2018) <= layer0_outputs(4517);
    outputs(2019) <= not(layer0_outputs(1058));
    outputs(2020) <= layer0_outputs(1309);
    outputs(2021) <= (layer0_outputs(2488)) xor (layer0_outputs(4018));
    outputs(2022) <= '0';
    outputs(2023) <= layer0_outputs(3326);
    outputs(2024) <= (layer0_outputs(3041)) and (layer0_outputs(4941));
    outputs(2025) <= not(layer0_outputs(2830)) or (layer0_outputs(516));
    outputs(2026) <= layer0_outputs(3781);
    outputs(2027) <= not(layer0_outputs(818));
    outputs(2028) <= not(layer0_outputs(621));
    outputs(2029) <= not((layer0_outputs(4618)) or (layer0_outputs(3320)));
    outputs(2030) <= not((layer0_outputs(666)) or (layer0_outputs(4314)));
    outputs(2031) <= layer0_outputs(5074);
    outputs(2032) <= not(layer0_outputs(4820));
    outputs(2033) <= not(layer0_outputs(3851));
    outputs(2034) <= not(layer0_outputs(1681));
    outputs(2035) <= not((layer0_outputs(1722)) and (layer0_outputs(2792)));
    outputs(2036) <= not((layer0_outputs(3888)) or (layer0_outputs(352)));
    outputs(2037) <= not(layer0_outputs(3247));
    outputs(2038) <= not(layer0_outputs(536)) or (layer0_outputs(1086));
    outputs(2039) <= not(layer0_outputs(3403));
    outputs(2040) <= not(layer0_outputs(4206));
    outputs(2041) <= not(layer0_outputs(274));
    outputs(2042) <= (layer0_outputs(1886)) and (layer0_outputs(1414));
    outputs(2043) <= layer0_outputs(1821);
    outputs(2044) <= (layer0_outputs(2776)) and not (layer0_outputs(5055));
    outputs(2045) <= not(layer0_outputs(1302));
    outputs(2046) <= not(layer0_outputs(5095));
    outputs(2047) <= (layer0_outputs(4258)) and (layer0_outputs(4654));
    outputs(2048) <= layer0_outputs(3161);
    outputs(2049) <= not(layer0_outputs(825));
    outputs(2050) <= layer0_outputs(1128);
    outputs(2051) <= (layer0_outputs(3268)) and (layer0_outputs(2631));
    outputs(2052) <= (layer0_outputs(2266)) and not (layer0_outputs(3141));
    outputs(2053) <= (layer0_outputs(2762)) and not (layer0_outputs(4536));
    outputs(2054) <= layer0_outputs(479);
    outputs(2055) <= not((layer0_outputs(714)) or (layer0_outputs(3397)));
    outputs(2056) <= layer0_outputs(4041);
    outputs(2057) <= not(layer0_outputs(1610));
    outputs(2058) <= not(layer0_outputs(5020));
    outputs(2059) <= not((layer0_outputs(5073)) xor (layer0_outputs(419)));
    outputs(2060) <= (layer0_outputs(523)) and (layer0_outputs(2514));
    outputs(2061) <= not(layer0_outputs(1553));
    outputs(2062) <= not(layer0_outputs(1409));
    outputs(2063) <= layer0_outputs(3099);
    outputs(2064) <= not(layer0_outputs(5079));
    outputs(2065) <= not(layer0_outputs(578));
    outputs(2066) <= layer0_outputs(145);
    outputs(2067) <= not((layer0_outputs(825)) and (layer0_outputs(2543)));
    outputs(2068) <= layer0_outputs(4861);
    outputs(2069) <= not(layer0_outputs(1700)) or (layer0_outputs(1013));
    outputs(2070) <= not((layer0_outputs(779)) xor (layer0_outputs(4431)));
    outputs(2071) <= layer0_outputs(3909);
    outputs(2072) <= not(layer0_outputs(1697));
    outputs(2073) <= not(layer0_outputs(998)) or (layer0_outputs(214));
    outputs(2074) <= layer0_outputs(2109);
    outputs(2075) <= layer0_outputs(4195);
    outputs(2076) <= not(layer0_outputs(4329)) or (layer0_outputs(3195));
    outputs(2077) <= not((layer0_outputs(2576)) and (layer0_outputs(2064)));
    outputs(2078) <= not(layer0_outputs(2675));
    outputs(2079) <= (layer0_outputs(4596)) and (layer0_outputs(891));
    outputs(2080) <= (layer0_outputs(4982)) and (layer0_outputs(4415));
    outputs(2081) <= layer0_outputs(841);
    outputs(2082) <= (layer0_outputs(3654)) and not (layer0_outputs(3294));
    outputs(2083) <= not(layer0_outputs(4662));
    outputs(2084) <= not(layer0_outputs(97));
    outputs(2085) <= not((layer0_outputs(1248)) xor (layer0_outputs(1790)));
    outputs(2086) <= (layer0_outputs(710)) and not (layer0_outputs(359));
    outputs(2087) <= layer0_outputs(1646);
    outputs(2088) <= layer0_outputs(684);
    outputs(2089) <= (layer0_outputs(3555)) and (layer0_outputs(890));
    outputs(2090) <= not(layer0_outputs(4058));
    outputs(2091) <= (layer0_outputs(1955)) and not (layer0_outputs(5044));
    outputs(2092) <= layer0_outputs(1453);
    outputs(2093) <= not((layer0_outputs(2038)) and (layer0_outputs(904)));
    outputs(2094) <= layer0_outputs(4836);
    outputs(2095) <= not(layer0_outputs(1416));
    outputs(2096) <= (layer0_outputs(2982)) and (layer0_outputs(2745));
    outputs(2097) <= layer0_outputs(143);
    outputs(2098) <= not((layer0_outputs(3136)) or (layer0_outputs(4192)));
    outputs(2099) <= layer0_outputs(4114);
    outputs(2100) <= not((layer0_outputs(1788)) or (layer0_outputs(2491)));
    outputs(2101) <= not(layer0_outputs(1782));
    outputs(2102) <= layer0_outputs(3405);
    outputs(2103) <= not(layer0_outputs(1917));
    outputs(2104) <= layer0_outputs(3657);
    outputs(2105) <= layer0_outputs(91);
    outputs(2106) <= layer0_outputs(2802);
    outputs(2107) <= layer0_outputs(2865);
    outputs(2108) <= not(layer0_outputs(2074));
    outputs(2109) <= layer0_outputs(4533);
    outputs(2110) <= (layer0_outputs(5034)) and not (layer0_outputs(2856));
    outputs(2111) <= not((layer0_outputs(385)) or (layer0_outputs(3643)));
    outputs(2112) <= not(layer0_outputs(4562));
    outputs(2113) <= not((layer0_outputs(2784)) xor (layer0_outputs(3955)));
    outputs(2114) <= (layer0_outputs(1342)) and (layer0_outputs(4969));
    outputs(2115) <= (layer0_outputs(2786)) and not (layer0_outputs(4024));
    outputs(2116) <= (layer0_outputs(1153)) and not (layer0_outputs(1857));
    outputs(2117) <= not(layer0_outputs(228));
    outputs(2118) <= layer0_outputs(2208);
    outputs(2119) <= not(layer0_outputs(3594));
    outputs(2120) <= layer0_outputs(2386);
    outputs(2121) <= not(layer0_outputs(894));
    outputs(2122) <= (layer0_outputs(2446)) and not (layer0_outputs(1949));
    outputs(2123) <= layer0_outputs(2261);
    outputs(2124) <= (layer0_outputs(2808)) and not (layer0_outputs(4374));
    outputs(2125) <= (layer0_outputs(3850)) and not (layer0_outputs(4633));
    outputs(2126) <= layer0_outputs(361);
    outputs(2127) <= layer0_outputs(240);
    outputs(2128) <= not((layer0_outputs(190)) xor (layer0_outputs(2691)));
    outputs(2129) <= layer0_outputs(2992);
    outputs(2130) <= (layer0_outputs(4183)) and (layer0_outputs(4267));
    outputs(2131) <= layer0_outputs(436);
    outputs(2132) <= layer0_outputs(3096);
    outputs(2133) <= not(layer0_outputs(4189));
    outputs(2134) <= (layer0_outputs(2433)) and not (layer0_outputs(1006));
    outputs(2135) <= not(layer0_outputs(2973));
    outputs(2136) <= not(layer0_outputs(3698));
    outputs(2137) <= layer0_outputs(498);
    outputs(2138) <= layer0_outputs(3956);
    outputs(2139) <= layer0_outputs(2775);
    outputs(2140) <= not((layer0_outputs(3638)) xor (layer0_outputs(3477)));
    outputs(2141) <= layer0_outputs(2601);
    outputs(2142) <= not((layer0_outputs(507)) and (layer0_outputs(321)));
    outputs(2143) <= layer0_outputs(1074);
    outputs(2144) <= not(layer0_outputs(4224)) or (layer0_outputs(3274));
    outputs(2145) <= not(layer0_outputs(5060));
    outputs(2146) <= layer0_outputs(1743);
    outputs(2147) <= not(layer0_outputs(2182)) or (layer0_outputs(1786));
    outputs(2148) <= (layer0_outputs(2637)) and not (layer0_outputs(577));
    outputs(2149) <= (layer0_outputs(951)) xor (layer0_outputs(2987));
    outputs(2150) <= not(layer0_outputs(4481));
    outputs(2151) <= not((layer0_outputs(2430)) and (layer0_outputs(5002)));
    outputs(2152) <= (layer0_outputs(4468)) xor (layer0_outputs(1860));
    outputs(2153) <= layer0_outputs(1531);
    outputs(2154) <= not((layer0_outputs(3995)) or (layer0_outputs(4732)));
    outputs(2155) <= layer0_outputs(306);
    outputs(2156) <= not(layer0_outputs(4149));
    outputs(2157) <= not(layer0_outputs(313));
    outputs(2158) <= not(layer0_outputs(1861)) or (layer0_outputs(3537));
    outputs(2159) <= not((layer0_outputs(955)) or (layer0_outputs(604)));
    outputs(2160) <= layer0_outputs(1859);
    outputs(2161) <= (layer0_outputs(3415)) and not (layer0_outputs(2110));
    outputs(2162) <= not(layer0_outputs(4616));
    outputs(2163) <= layer0_outputs(2984);
    outputs(2164) <= not(layer0_outputs(778)) or (layer0_outputs(1024));
    outputs(2165) <= not(layer0_outputs(4284)) or (layer0_outputs(860));
    outputs(2166) <= (layer0_outputs(2478)) or (layer0_outputs(4635));
    outputs(2167) <= (layer0_outputs(3970)) and not (layer0_outputs(2903));
    outputs(2168) <= not(layer0_outputs(2359));
    outputs(2169) <= not(layer0_outputs(4825));
    outputs(2170) <= (layer0_outputs(4534)) xor (layer0_outputs(214));
    outputs(2171) <= layer0_outputs(3699);
    outputs(2172) <= layer0_outputs(4463);
    outputs(2173) <= not((layer0_outputs(1901)) or (layer0_outputs(499)));
    outputs(2174) <= not(layer0_outputs(2365));
    outputs(2175) <= not((layer0_outputs(3761)) xor (layer0_outputs(2559)));
    outputs(2176) <= not(layer0_outputs(3344)) or (layer0_outputs(2262));
    outputs(2177) <= not(layer0_outputs(4217));
    outputs(2178) <= layer0_outputs(2249);
    outputs(2179) <= not(layer0_outputs(2873));
    outputs(2180) <= not(layer0_outputs(445));
    outputs(2181) <= layer0_outputs(4769);
    outputs(2182) <= not(layer0_outputs(3767));
    outputs(2183) <= layer0_outputs(4819);
    outputs(2184) <= (layer0_outputs(415)) and (layer0_outputs(4105));
    outputs(2185) <= not((layer0_outputs(192)) or (layer0_outputs(2288)));
    outputs(2186) <= layer0_outputs(5114);
    outputs(2187) <= layer0_outputs(2563);
    outputs(2188) <= (layer0_outputs(497)) xor (layer0_outputs(159));
    outputs(2189) <= (layer0_outputs(1835)) and not (layer0_outputs(1994));
    outputs(2190) <= (layer0_outputs(1074)) and not (layer0_outputs(2218));
    outputs(2191) <= not(layer0_outputs(3297));
    outputs(2192) <= (layer0_outputs(1255)) and not (layer0_outputs(766));
    outputs(2193) <= (layer0_outputs(2673)) and (layer0_outputs(272));
    outputs(2194) <= layer0_outputs(272);
    outputs(2195) <= not(layer0_outputs(631));
    outputs(2196) <= layer0_outputs(1272);
    outputs(2197) <= layer0_outputs(3428);
    outputs(2198) <= not((layer0_outputs(623)) xor (layer0_outputs(4563)));
    outputs(2199) <= not(layer0_outputs(686));
    outputs(2200) <= not(layer0_outputs(4136));
    outputs(2201) <= (layer0_outputs(3743)) and not (layer0_outputs(373));
    outputs(2202) <= (layer0_outputs(598)) and not (layer0_outputs(1932));
    outputs(2203) <= not((layer0_outputs(5089)) and (layer0_outputs(2667)));
    outputs(2204) <= not(layer0_outputs(237));
    outputs(2205) <= not(layer0_outputs(292));
    outputs(2206) <= (layer0_outputs(2609)) and not (layer0_outputs(357));
    outputs(2207) <= (layer0_outputs(1939)) and not (layer0_outputs(4870));
    outputs(2208) <= not(layer0_outputs(3073));
    outputs(2209) <= (layer0_outputs(634)) and not (layer0_outputs(4776));
    outputs(2210) <= not(layer0_outputs(1593));
    outputs(2211) <= not(layer0_outputs(691));
    outputs(2212) <= not(layer0_outputs(3160));
    outputs(2213) <= layer0_outputs(1621);
    outputs(2214) <= not(layer0_outputs(2583));
    outputs(2215) <= (layer0_outputs(2955)) or (layer0_outputs(3502));
    outputs(2216) <= (layer0_outputs(4420)) and not (layer0_outputs(4492));
    outputs(2217) <= not(layer0_outputs(5063));
    outputs(2218) <= (layer0_outputs(106)) and not (layer0_outputs(3279));
    outputs(2219) <= layer0_outputs(3915);
    outputs(2220) <= (layer0_outputs(613)) and not (layer0_outputs(3582));
    outputs(2221) <= not(layer0_outputs(1140));
    outputs(2222) <= layer0_outputs(3353);
    outputs(2223) <= not(layer0_outputs(1117));
    outputs(2224) <= layer0_outputs(4971);
    outputs(2225) <= (layer0_outputs(3969)) or (layer0_outputs(2401));
    outputs(2226) <= layer0_outputs(1171);
    outputs(2227) <= not((layer0_outputs(4055)) or (layer0_outputs(59)));
    outputs(2228) <= not((layer0_outputs(2799)) xor (layer0_outputs(1705)));
    outputs(2229) <= not(layer0_outputs(3637)) or (layer0_outputs(2652));
    outputs(2230) <= (layer0_outputs(3716)) and not (layer0_outputs(3462));
    outputs(2231) <= (layer0_outputs(1099)) and not (layer0_outputs(122));
    outputs(2232) <= not((layer0_outputs(3625)) or (layer0_outputs(4626)));
    outputs(2233) <= (layer0_outputs(254)) and not (layer0_outputs(2226));
    outputs(2234) <= layer0_outputs(925);
    outputs(2235) <= layer0_outputs(2310);
    outputs(2236) <= layer0_outputs(2966);
    outputs(2237) <= not(layer0_outputs(445));
    outputs(2238) <= not(layer0_outputs(2964));
    outputs(2239) <= (layer0_outputs(3591)) and (layer0_outputs(399));
    outputs(2240) <= not(layer0_outputs(304));
    outputs(2241) <= layer0_outputs(605);
    outputs(2242) <= layer0_outputs(4042);
    outputs(2243) <= (layer0_outputs(2159)) xor (layer0_outputs(2748));
    outputs(2244) <= not(layer0_outputs(4443));
    outputs(2245) <= not(layer0_outputs(1756)) or (layer0_outputs(1210));
    outputs(2246) <= not(layer0_outputs(969));
    outputs(2247) <= (layer0_outputs(1499)) and (layer0_outputs(2468));
    outputs(2248) <= not(layer0_outputs(3420));
    outputs(2249) <= layer0_outputs(3665);
    outputs(2250) <= not(layer0_outputs(649));
    outputs(2251) <= not(layer0_outputs(2576));
    outputs(2252) <= layer0_outputs(1444);
    outputs(2253) <= (layer0_outputs(3287)) and not (layer0_outputs(194));
    outputs(2254) <= not(layer0_outputs(3857));
    outputs(2255) <= not((layer0_outputs(1989)) and (layer0_outputs(3094)));
    outputs(2256) <= (layer0_outputs(2787)) and (layer0_outputs(4718));
    outputs(2257) <= not(layer0_outputs(4439));
    outputs(2258) <= (layer0_outputs(3931)) or (layer0_outputs(2134));
    outputs(2259) <= not(layer0_outputs(3431));
    outputs(2260) <= (layer0_outputs(1120)) and not (layer0_outputs(4737));
    outputs(2261) <= (layer0_outputs(2529)) and not (layer0_outputs(2659));
    outputs(2262) <= not(layer0_outputs(354));
    outputs(2263) <= not(layer0_outputs(4377)) or (layer0_outputs(2919));
    outputs(2264) <= layer0_outputs(3682);
    outputs(2265) <= not(layer0_outputs(2358));
    outputs(2266) <= (layer0_outputs(3599)) and not (layer0_outputs(3247));
    outputs(2267) <= not((layer0_outputs(4395)) or (layer0_outputs(2120)));
    outputs(2268) <= (layer0_outputs(3890)) and (layer0_outputs(1260));
    outputs(2269) <= layer0_outputs(1704);
    outputs(2270) <= layer0_outputs(613);
    outputs(2271) <= not(layer0_outputs(2654));
    outputs(2272) <= not(layer0_outputs(1116));
    outputs(2273) <= not(layer0_outputs(3521));
    outputs(2274) <= (layer0_outputs(1392)) and not (layer0_outputs(235));
    outputs(2275) <= layer0_outputs(3251);
    outputs(2276) <= (layer0_outputs(2777)) xor (layer0_outputs(2853));
    outputs(2277) <= layer0_outputs(4799);
    outputs(2278) <= not((layer0_outputs(1036)) xor (layer0_outputs(3493)));
    outputs(2279) <= (layer0_outputs(3197)) and not (layer0_outputs(3922));
    outputs(2280) <= (layer0_outputs(1619)) and (layer0_outputs(4993));
    outputs(2281) <= not((layer0_outputs(3498)) or (layer0_outputs(194)));
    outputs(2282) <= layer0_outputs(204);
    outputs(2283) <= layer0_outputs(2765);
    outputs(2284) <= not(layer0_outputs(2833));
    outputs(2285) <= (layer0_outputs(1090)) and not (layer0_outputs(4295));
    outputs(2286) <= (layer0_outputs(3426)) xor (layer0_outputs(1417));
    outputs(2287) <= layer0_outputs(759);
    outputs(2288) <= not((layer0_outputs(4097)) or (layer0_outputs(2250)));
    outputs(2289) <= not(layer0_outputs(923));
    outputs(2290) <= layer0_outputs(249);
    outputs(2291) <= (layer0_outputs(986)) xor (layer0_outputs(1229));
    outputs(2292) <= layer0_outputs(2752);
    outputs(2293) <= not(layer0_outputs(1067));
    outputs(2294) <= not(layer0_outputs(1656));
    outputs(2295) <= layer0_outputs(1490);
    outputs(2296) <= not((layer0_outputs(4666)) or (layer0_outputs(75)));
    outputs(2297) <= not(layer0_outputs(3690));
    outputs(2298) <= not(layer0_outputs(2479));
    outputs(2299) <= not(layer0_outputs(79));
    outputs(2300) <= (layer0_outputs(2527)) xor (layer0_outputs(1768));
    outputs(2301) <= (layer0_outputs(513)) and not (layer0_outputs(2220));
    outputs(2302) <= layer0_outputs(1747);
    outputs(2303) <= not((layer0_outputs(2979)) or (layer0_outputs(2427)));
    outputs(2304) <= (layer0_outputs(80)) and (layer0_outputs(2716));
    outputs(2305) <= not((layer0_outputs(353)) or (layer0_outputs(4376)));
    outputs(2306) <= not(layer0_outputs(617));
    outputs(2307) <= layer0_outputs(635);
    outputs(2308) <= (layer0_outputs(3330)) or (layer0_outputs(3167));
    outputs(2309) <= not((layer0_outputs(5061)) or (layer0_outputs(2805)));
    outputs(2310) <= not((layer0_outputs(4645)) or (layer0_outputs(1755)));
    outputs(2311) <= (layer0_outputs(117)) and (layer0_outputs(4096));
    outputs(2312) <= not((layer0_outputs(2049)) or (layer0_outputs(5104)));
    outputs(2313) <= layer0_outputs(1803);
    outputs(2314) <= layer0_outputs(1770);
    outputs(2315) <= not((layer0_outputs(4169)) or (layer0_outputs(1684)));
    outputs(2316) <= not(layer0_outputs(2410));
    outputs(2317) <= (layer0_outputs(3497)) and (layer0_outputs(4953));
    outputs(2318) <= not(layer0_outputs(3283));
    outputs(2319) <= not((layer0_outputs(4241)) xor (layer0_outputs(2928)));
    outputs(2320) <= layer0_outputs(1840);
    outputs(2321) <= not(layer0_outputs(4516));
    outputs(2322) <= not(layer0_outputs(1196));
    outputs(2323) <= layer0_outputs(3334);
    outputs(2324) <= not(layer0_outputs(2588)) or (layer0_outputs(4938));
    outputs(2325) <= (layer0_outputs(4064)) and not (layer0_outputs(1147));
    outputs(2326) <= not((layer0_outputs(3729)) or (layer0_outputs(2355)));
    outputs(2327) <= (layer0_outputs(1653)) and not (layer0_outputs(2096));
    outputs(2328) <= not(layer0_outputs(1765));
    outputs(2329) <= (layer0_outputs(2831)) and not (layer0_outputs(4108));
    outputs(2330) <= not((layer0_outputs(2559)) xor (layer0_outputs(3585)));
    outputs(2331) <= layer0_outputs(4686);
    outputs(2332) <= (layer0_outputs(1921)) and not (layer0_outputs(3439));
    outputs(2333) <= not(layer0_outputs(216));
    outputs(2334) <= not(layer0_outputs(3934));
    outputs(2335) <= layer0_outputs(4336);
    outputs(2336) <= not(layer0_outputs(4617));
    outputs(2337) <= (layer0_outputs(3329)) xor (layer0_outputs(4763));
    outputs(2338) <= layer0_outputs(3593);
    outputs(2339) <= layer0_outputs(2132);
    outputs(2340) <= not(layer0_outputs(3683));
    outputs(2341) <= not((layer0_outputs(4903)) or (layer0_outputs(591)));
    outputs(2342) <= layer0_outputs(3692);
    outputs(2343) <= layer0_outputs(1832);
    outputs(2344) <= layer0_outputs(1014);
    outputs(2345) <= layer0_outputs(4038);
    outputs(2346) <= (layer0_outputs(3732)) and (layer0_outputs(3084));
    outputs(2347) <= not((layer0_outputs(661)) or (layer0_outputs(354)));
    outputs(2348) <= (layer0_outputs(3)) xor (layer0_outputs(1586));
    outputs(2349) <= not((layer0_outputs(577)) or (layer0_outputs(5097)));
    outputs(2350) <= layer0_outputs(1536);
    outputs(2351) <= layer0_outputs(436);
    outputs(2352) <= (layer0_outputs(3666)) and not (layer0_outputs(70));
    outputs(2353) <= not(layer0_outputs(2602));
    outputs(2354) <= (layer0_outputs(2989)) and not (layer0_outputs(1915));
    outputs(2355) <= (layer0_outputs(2065)) and not (layer0_outputs(244));
    outputs(2356) <= (layer0_outputs(4996)) and (layer0_outputs(4078));
    outputs(2357) <= layer0_outputs(2644);
    outputs(2358) <= layer0_outputs(1791);
    outputs(2359) <= (layer0_outputs(233)) and not (layer0_outputs(4311));
    outputs(2360) <= not(layer0_outputs(2706));
    outputs(2361) <= layer0_outputs(3074);
    outputs(2362) <= not(layer0_outputs(1787));
    outputs(2363) <= not(layer0_outputs(4197));
    outputs(2364) <= not(layer0_outputs(112));
    outputs(2365) <= layer0_outputs(82);
    outputs(2366) <= layer0_outputs(705);
    outputs(2367) <= layer0_outputs(4020);
    outputs(2368) <= not(layer0_outputs(1359));
    outputs(2369) <= (layer0_outputs(2354)) and not (layer0_outputs(3303));
    outputs(2370) <= (layer0_outputs(1639)) xor (layer0_outputs(1227));
    outputs(2371) <= not(layer0_outputs(2639));
    outputs(2372) <= not(layer0_outputs(2218));
    outputs(2373) <= not((layer0_outputs(1193)) xor (layer0_outputs(4093)));
    outputs(2374) <= layer0_outputs(977);
    outputs(2375) <= not(layer0_outputs(3730));
    outputs(2376) <= layer0_outputs(3764);
    outputs(2377) <= not(layer0_outputs(3259));
    outputs(2378) <= (layer0_outputs(1202)) and (layer0_outputs(3837));
    outputs(2379) <= layer0_outputs(829);
    outputs(2380) <= (layer0_outputs(56)) and (layer0_outputs(4859));
    outputs(2381) <= (layer0_outputs(1387)) and (layer0_outputs(4457));
    outputs(2382) <= not(layer0_outputs(3533));
    outputs(2383) <= not(layer0_outputs(1926));
    outputs(2384) <= not((layer0_outputs(1155)) or (layer0_outputs(1573)));
    outputs(2385) <= layer0_outputs(2991);
    outputs(2386) <= (layer0_outputs(2416)) and not (layer0_outputs(392));
    outputs(2387) <= not((layer0_outputs(2483)) xor (layer0_outputs(4037)));
    outputs(2388) <= not(layer0_outputs(974));
    outputs(2389) <= layer0_outputs(4451);
    outputs(2390) <= layer0_outputs(2820);
    outputs(2391) <= (layer0_outputs(4162)) and not (layer0_outputs(4301));
    outputs(2392) <= not(layer0_outputs(333));
    outputs(2393) <= not(layer0_outputs(4580));
    outputs(2394) <= not(layer0_outputs(3572));
    outputs(2395) <= not(layer0_outputs(834));
    outputs(2396) <= (layer0_outputs(93)) and not (layer0_outputs(1051));
    outputs(2397) <= not(layer0_outputs(4481));
    outputs(2398) <= not(layer0_outputs(70)) or (layer0_outputs(1456));
    outputs(2399) <= not(layer0_outputs(1344));
    outputs(2400) <= not(layer0_outputs(1949));
    outputs(2401) <= not(layer0_outputs(556));
    outputs(2402) <= not(layer0_outputs(905));
    outputs(2403) <= not((layer0_outputs(518)) and (layer0_outputs(2234)));
    outputs(2404) <= not((layer0_outputs(3984)) xor (layer0_outputs(4306)));
    outputs(2405) <= not((layer0_outputs(900)) and (layer0_outputs(5046)));
    outputs(2406) <= layer0_outputs(2894);
    outputs(2407) <= not((layer0_outputs(2051)) or (layer0_outputs(4253)));
    outputs(2408) <= not(layer0_outputs(367));
    outputs(2409) <= layer0_outputs(3562);
    outputs(2410) <= not(layer0_outputs(2498));
    outputs(2411) <= layer0_outputs(2425);
    outputs(2412) <= layer0_outputs(1241);
    outputs(2413) <= (layer0_outputs(4897)) and (layer0_outputs(1011));
    outputs(2414) <= not(layer0_outputs(5007));
    outputs(2415) <= not((layer0_outputs(257)) or (layer0_outputs(4826)));
    outputs(2416) <= (layer0_outputs(2645)) xor (layer0_outputs(86));
    outputs(2417) <= layer0_outputs(1556);
    outputs(2418) <= not((layer0_outputs(1738)) or (layer0_outputs(3798)));
    outputs(2419) <= (layer0_outputs(1429)) or (layer0_outputs(4917));
    outputs(2420) <= not(layer0_outputs(308));
    outputs(2421) <= (layer0_outputs(1309)) and not (layer0_outputs(1023));
    outputs(2422) <= not(layer0_outputs(1053));
    outputs(2423) <= (layer0_outputs(689)) and not (layer0_outputs(734));
    outputs(2424) <= not(layer0_outputs(4379));
    outputs(2425) <= (layer0_outputs(2504)) and (layer0_outputs(3052));
    outputs(2426) <= layer0_outputs(2362);
    outputs(2427) <= (layer0_outputs(843)) xor (layer0_outputs(1305));
    outputs(2428) <= not(layer0_outputs(3111));
    outputs(2429) <= layer0_outputs(3894);
    outputs(2430) <= (layer0_outputs(2424)) xor (layer0_outputs(2664));
    outputs(2431) <= (layer0_outputs(4008)) and not (layer0_outputs(4947));
    outputs(2432) <= not(layer0_outputs(1929));
    outputs(2433) <= not(layer0_outputs(510));
    outputs(2434) <= layer0_outputs(2088);
    outputs(2435) <= not(layer0_outputs(467));
    outputs(2436) <= (layer0_outputs(3998)) and (layer0_outputs(5017));
    outputs(2437) <= not(layer0_outputs(2385));
    outputs(2438) <= (layer0_outputs(4103)) and not (layer0_outputs(2801));
    outputs(2439) <= layer0_outputs(2538);
    outputs(2440) <= (layer0_outputs(2463)) and not (layer0_outputs(2872));
    outputs(2441) <= layer0_outputs(4206);
    outputs(2442) <= not(layer0_outputs(1042));
    outputs(2443) <= layer0_outputs(3541);
    outputs(2444) <= not((layer0_outputs(1163)) or (layer0_outputs(4436)));
    outputs(2445) <= not(layer0_outputs(41));
    outputs(2446) <= layer0_outputs(3773);
    outputs(2447) <= layer0_outputs(1783);
    outputs(2448) <= not(layer0_outputs(1904));
    outputs(2449) <= not((layer0_outputs(1620)) and (layer0_outputs(2748)));
    outputs(2450) <= layer0_outputs(3352);
    outputs(2451) <= not(layer0_outputs(3030));
    outputs(2452) <= layer0_outputs(4781);
    outputs(2453) <= layer0_outputs(1250);
    outputs(2454) <= layer0_outputs(4259);
    outputs(2455) <= not(layer0_outputs(814)) or (layer0_outputs(4422));
    outputs(2456) <= layer0_outputs(293);
    outputs(2457) <= not((layer0_outputs(3119)) xor (layer0_outputs(2708)));
    outputs(2458) <= not((layer0_outputs(927)) xor (layer0_outputs(546)));
    outputs(2459) <= layer0_outputs(361);
    outputs(2460) <= not(layer0_outputs(3880)) or (layer0_outputs(4761));
    outputs(2461) <= not(layer0_outputs(1500));
    outputs(2462) <= not(layer0_outputs(719));
    outputs(2463) <= layer0_outputs(3810);
    outputs(2464) <= layer0_outputs(4799);
    outputs(2465) <= layer0_outputs(4243);
    outputs(2466) <= not((layer0_outputs(3924)) or (layer0_outputs(2947)));
    outputs(2467) <= not(layer0_outputs(4443));
    outputs(2468) <= (layer0_outputs(2850)) and not (layer0_outputs(3098));
    outputs(2469) <= not((layer0_outputs(1116)) or (layer0_outputs(2590)));
    outputs(2470) <= layer0_outputs(3006);
    outputs(2471) <= (layer0_outputs(4872)) and not (layer0_outputs(5043));
    outputs(2472) <= (layer0_outputs(2035)) and not (layer0_outputs(4497));
    outputs(2473) <= (layer0_outputs(1895)) and not (layer0_outputs(360));
    outputs(2474) <= layer0_outputs(3045);
    outputs(2475) <= (layer0_outputs(4736)) and not (layer0_outputs(3294));
    outputs(2476) <= not(layer0_outputs(2387));
    outputs(2477) <= not(layer0_outputs(1677));
    outputs(2478) <= not(layer0_outputs(1893));
    outputs(2479) <= (layer0_outputs(3106)) and not (layer0_outputs(53));
    outputs(2480) <= layer0_outputs(4675);
    outputs(2481) <= not(layer0_outputs(1427));
    outputs(2482) <= (layer0_outputs(3846)) and not (layer0_outputs(3454));
    outputs(2483) <= not(layer0_outputs(3214));
    outputs(2484) <= not(layer0_outputs(3463));
    outputs(2485) <= layer0_outputs(4382);
    outputs(2486) <= (layer0_outputs(498)) and not (layer0_outputs(3522));
    outputs(2487) <= (layer0_outputs(1401)) and not (layer0_outputs(394));
    outputs(2488) <= (layer0_outputs(2676)) and not (layer0_outputs(2606));
    outputs(2489) <= layer0_outputs(1725);
    outputs(2490) <= layer0_outputs(2713);
    outputs(2491) <= not(layer0_outputs(1633));
    outputs(2492) <= not(layer0_outputs(519));
    outputs(2493) <= (layer0_outputs(1055)) xor (layer0_outputs(3917));
    outputs(2494) <= not(layer0_outputs(2848));
    outputs(2495) <= (layer0_outputs(3316)) and (layer0_outputs(526));
    outputs(2496) <= (layer0_outputs(1530)) or (layer0_outputs(2593));
    outputs(2497) <= not(layer0_outputs(4934));
    outputs(2498) <= not(layer0_outputs(5011)) or (layer0_outputs(53));
    outputs(2499) <= (layer0_outputs(1339)) and (layer0_outputs(4478));
    outputs(2500) <= (layer0_outputs(795)) and not (layer0_outputs(2883));
    outputs(2501) <= layer0_outputs(4246);
    outputs(2502) <= not((layer0_outputs(1070)) xor (layer0_outputs(3341)));
    outputs(2503) <= not(layer0_outputs(2150));
    outputs(2504) <= not((layer0_outputs(2770)) or (layer0_outputs(3590)));
    outputs(2505) <= not((layer0_outputs(3630)) and (layer0_outputs(2071)));
    outputs(2506) <= not((layer0_outputs(3755)) or (layer0_outputs(2148)));
    outputs(2507) <= (layer0_outputs(2628)) xor (layer0_outputs(1150));
    outputs(2508) <= not((layer0_outputs(3806)) xor (layer0_outputs(3464)));
    outputs(2509) <= (layer0_outputs(4840)) and not (layer0_outputs(4051));
    outputs(2510) <= layer0_outputs(3605);
    outputs(2511) <= not((layer0_outputs(1131)) and (layer0_outputs(105)));
    outputs(2512) <= layer0_outputs(118);
    outputs(2513) <= layer0_outputs(3941);
    outputs(2514) <= (layer0_outputs(3229)) and (layer0_outputs(3103));
    outputs(2515) <= not(layer0_outputs(878));
    outputs(2516) <= not(layer0_outputs(1922));
    outputs(2517) <= not(layer0_outputs(1019));
    outputs(2518) <= not((layer0_outputs(4754)) or (layer0_outputs(2823)));
    outputs(2519) <= (layer0_outputs(438)) and not (layer0_outputs(3277));
    outputs(2520) <= not(layer0_outputs(3326));
    outputs(2521) <= (layer0_outputs(1299)) and (layer0_outputs(1609));
    outputs(2522) <= layer0_outputs(4054);
    outputs(2523) <= layer0_outputs(4418);
    outputs(2524) <= layer0_outputs(4749);
    outputs(2525) <= (layer0_outputs(277)) and not (layer0_outputs(2239));
    outputs(2526) <= (layer0_outputs(5009)) xor (layer0_outputs(4102));
    outputs(2527) <= not(layer0_outputs(1983));
    outputs(2528) <= not(layer0_outputs(1700));
    outputs(2529) <= not(layer0_outputs(2036)) or (layer0_outputs(92));
    outputs(2530) <= layer0_outputs(3952);
    outputs(2531) <= not(layer0_outputs(3408));
    outputs(2532) <= layer0_outputs(2594);
    outputs(2533) <= (layer0_outputs(4891)) or (layer0_outputs(1536));
    outputs(2534) <= (layer0_outputs(2980)) and (layer0_outputs(5057));
    outputs(2535) <= layer0_outputs(2227);
    outputs(2536) <= not(layer0_outputs(1633));
    outputs(2537) <= (layer0_outputs(2362)) and not (layer0_outputs(919));
    outputs(2538) <= layer0_outputs(2300);
    outputs(2539) <= not(layer0_outputs(4320));
    outputs(2540) <= layer0_outputs(4033);
    outputs(2541) <= (layer0_outputs(3449)) and not (layer0_outputs(3108));
    outputs(2542) <= (layer0_outputs(5071)) and (layer0_outputs(3597));
    outputs(2543) <= layer0_outputs(1189);
    outputs(2544) <= layer0_outputs(2913);
    outputs(2545) <= not(layer0_outputs(1252));
    outputs(2546) <= layer0_outputs(1796);
    outputs(2547) <= (layer0_outputs(3556)) and not (layer0_outputs(144));
    outputs(2548) <= (layer0_outputs(91)) or (layer0_outputs(1193));
    outputs(2549) <= (layer0_outputs(4980)) and not (layer0_outputs(3705));
    outputs(2550) <= not(layer0_outputs(2455));
    outputs(2551) <= not(layer0_outputs(5033));
    outputs(2552) <= (layer0_outputs(417)) and not (layer0_outputs(3454));
    outputs(2553) <= (layer0_outputs(681)) and not (layer0_outputs(228));
    outputs(2554) <= layer0_outputs(3765);
    outputs(2555) <= (layer0_outputs(2622)) and (layer0_outputs(4582));
    outputs(2556) <= (layer0_outputs(1753)) and not (layer0_outputs(78));
    outputs(2557) <= not(layer0_outputs(1837));
    outputs(2558) <= not(layer0_outputs(699));
    outputs(2559) <= layer0_outputs(933);
    outputs(2560) <= not(layer0_outputs(1211));
    outputs(2561) <= not(layer0_outputs(4767));
    outputs(2562) <= (layer0_outputs(1585)) xor (layer0_outputs(57));
    outputs(2563) <= not(layer0_outputs(41));
    outputs(2564) <= (layer0_outputs(4442)) or (layer0_outputs(1051));
    outputs(2565) <= not(layer0_outputs(3448));
    outputs(2566) <= not((layer0_outputs(672)) xor (layer0_outputs(1774)));
    outputs(2567) <= layer0_outputs(431);
    outputs(2568) <= not((layer0_outputs(2578)) and (layer0_outputs(213)));
    outputs(2569) <= not((layer0_outputs(1515)) xor (layer0_outputs(4521)));
    outputs(2570) <= layer0_outputs(2654);
    outputs(2571) <= not((layer0_outputs(2077)) or (layer0_outputs(2957)));
    outputs(2572) <= layer0_outputs(2515);
    outputs(2573) <= (layer0_outputs(4790)) and not (layer0_outputs(3111));
    outputs(2574) <= not(layer0_outputs(1531));
    outputs(2575) <= not(layer0_outputs(4954)) or (layer0_outputs(4669));
    outputs(2576) <= not(layer0_outputs(2737));
    outputs(2577) <= (layer0_outputs(1873)) xor (layer0_outputs(1138));
    outputs(2578) <= layer0_outputs(1982);
    outputs(2579) <= not(layer0_outputs(1795));
    outputs(2580) <= layer0_outputs(614);
    outputs(2581) <= not(layer0_outputs(2205));
    outputs(2582) <= (layer0_outputs(3768)) xor (layer0_outputs(2540));
    outputs(2583) <= not((layer0_outputs(4376)) or (layer0_outputs(753)));
    outputs(2584) <= (layer0_outputs(4665)) and not (layer0_outputs(4544));
    outputs(2585) <= layer0_outputs(3349);
    outputs(2586) <= (layer0_outputs(1157)) and (layer0_outputs(4001));
    outputs(2587) <= (layer0_outputs(4862)) or (layer0_outputs(1968));
    outputs(2588) <= (layer0_outputs(123)) and not (layer0_outputs(349));
    outputs(2589) <= not(layer0_outputs(148)) or (layer0_outputs(4914));
    outputs(2590) <= (layer0_outputs(903)) and not (layer0_outputs(310));
    outputs(2591) <= (layer0_outputs(736)) and not (layer0_outputs(3841));
    outputs(2592) <= not(layer0_outputs(1956));
    outputs(2593) <= layer0_outputs(3946);
    outputs(2594) <= not(layer0_outputs(1792)) or (layer0_outputs(3997));
    outputs(2595) <= layer0_outputs(351);
    outputs(2596) <= not(layer0_outputs(4587));
    outputs(2597) <= (layer0_outputs(1584)) xor (layer0_outputs(1158));
    outputs(2598) <= (layer0_outputs(128)) and not (layer0_outputs(2791));
    outputs(2599) <= layer0_outputs(2165);
    outputs(2600) <= layer0_outputs(2375);
    outputs(2601) <= not(layer0_outputs(2582));
    outputs(2602) <= not(layer0_outputs(1673)) or (layer0_outputs(2116));
    outputs(2603) <= (layer0_outputs(4565)) and not (layer0_outputs(793));
    outputs(2604) <= not((layer0_outputs(1419)) xor (layer0_outputs(3992)));
    outputs(2605) <= (layer0_outputs(3757)) or (layer0_outputs(1258));
    outputs(2606) <= not(layer0_outputs(1096));
    outputs(2607) <= not(layer0_outputs(1214));
    outputs(2608) <= not((layer0_outputs(481)) or (layer0_outputs(4164)));
    outputs(2609) <= not(layer0_outputs(1276));
    outputs(2610) <= not(layer0_outputs(3876));
    outputs(2611) <= layer0_outputs(5100);
    outputs(2612) <= not(layer0_outputs(4281));
    outputs(2613) <= not(layer0_outputs(2012)) or (layer0_outputs(4259));
    outputs(2614) <= (layer0_outputs(4364)) xor (layer0_outputs(2270));
    outputs(2615) <= not(layer0_outputs(1634));
    outputs(2616) <= layer0_outputs(4528);
    outputs(2617) <= not(layer0_outputs(2973));
    outputs(2618) <= not((layer0_outputs(2228)) or (layer0_outputs(18)));
    outputs(2619) <= not((layer0_outputs(225)) and (layer0_outputs(923)));
    outputs(2620) <= not(layer0_outputs(2731));
    outputs(2621) <= not(layer0_outputs(2306));
    outputs(2622) <= layer0_outputs(1084);
    outputs(2623) <= not((layer0_outputs(4230)) or (layer0_outputs(124)));
    outputs(2624) <= not((layer0_outputs(3413)) xor (layer0_outputs(4140)));
    outputs(2625) <= (layer0_outputs(2202)) or (layer0_outputs(5065));
    outputs(2626) <= not((layer0_outputs(4191)) xor (layer0_outputs(3892)));
    outputs(2627) <= not(layer0_outputs(3701));
    outputs(2628) <= not((layer0_outputs(2810)) xor (layer0_outputs(4109)));
    outputs(2629) <= not(layer0_outputs(4142));
    outputs(2630) <= not(layer0_outputs(4185));
    outputs(2631) <= (layer0_outputs(2457)) xor (layer0_outputs(3180));
    outputs(2632) <= not(layer0_outputs(4232));
    outputs(2633) <= (layer0_outputs(991)) and not (layer0_outputs(1730));
    outputs(2634) <= not((layer0_outputs(1533)) xor (layer0_outputs(185)));
    outputs(2635) <= not(layer0_outputs(1462)) or (layer0_outputs(4137));
    outputs(2636) <= layer0_outputs(2895);
    outputs(2637) <= layer0_outputs(1913);
    outputs(2638) <= not((layer0_outputs(4004)) xor (layer0_outputs(3864)));
    outputs(2639) <= layer0_outputs(3835);
    outputs(2640) <= not((layer0_outputs(4226)) and (layer0_outputs(1777)));
    outputs(2641) <= layer0_outputs(2327);
    outputs(2642) <= not((layer0_outputs(4047)) xor (layer0_outputs(5112)));
    outputs(2643) <= not((layer0_outputs(3151)) or (layer0_outputs(1257)));
    outputs(2644) <= layer0_outputs(1105);
    outputs(2645) <= not(layer0_outputs(913));
    outputs(2646) <= layer0_outputs(4769);
    outputs(2647) <= not(layer0_outputs(4123)) or (layer0_outputs(4462));
    outputs(2648) <= (layer0_outputs(1237)) and (layer0_outputs(1725));
    outputs(2649) <= (layer0_outputs(1422)) or (layer0_outputs(2690));
    outputs(2650) <= not(layer0_outputs(3811));
    outputs(2651) <= (layer0_outputs(1761)) and (layer0_outputs(3691));
    outputs(2652) <= (layer0_outputs(618)) xor (layer0_outputs(4047));
    outputs(2653) <= not(layer0_outputs(743));
    outputs(2654) <= (layer0_outputs(3257)) and (layer0_outputs(2445));
    outputs(2655) <= not(layer0_outputs(4254));
    outputs(2656) <= not((layer0_outputs(946)) xor (layer0_outputs(395)));
    outputs(2657) <= not(layer0_outputs(3423)) or (layer0_outputs(3403));
    outputs(2658) <= layer0_outputs(4893);
    outputs(2659) <= (layer0_outputs(251)) xor (layer0_outputs(5094));
    outputs(2660) <= not(layer0_outputs(4151));
    outputs(2661) <= (layer0_outputs(3137)) and (layer0_outputs(2331));
    outputs(2662) <= layer0_outputs(1525);
    outputs(2663) <= not(layer0_outputs(4341));
    outputs(2664) <= not((layer0_outputs(160)) xor (layer0_outputs(4006)));
    outputs(2665) <= not(layer0_outputs(5053));
    outputs(2666) <= layer0_outputs(2423);
    outputs(2667) <= not(layer0_outputs(3221)) or (layer0_outputs(242));
    outputs(2668) <= layer0_outputs(1000);
    outputs(2669) <= not(layer0_outputs(4083));
    outputs(2670) <= not(layer0_outputs(611)) or (layer0_outputs(908));
    outputs(2671) <= not(layer0_outputs(1300));
    outputs(2672) <= layer0_outputs(586);
    outputs(2673) <= not(layer0_outputs(2719));
    outputs(2674) <= layer0_outputs(2124);
    outputs(2675) <= (layer0_outputs(4372)) and not (layer0_outputs(1024));
    outputs(2676) <= not((layer0_outputs(4786)) or (layer0_outputs(2651)));
    outputs(2677) <= layer0_outputs(2910);
    outputs(2678) <= layer0_outputs(846);
    outputs(2679) <= (layer0_outputs(1416)) or (layer0_outputs(2508));
    outputs(2680) <= not((layer0_outputs(325)) xor (layer0_outputs(2564)));
    outputs(2681) <= (layer0_outputs(163)) xor (layer0_outputs(2495));
    outputs(2682) <= (layer0_outputs(2444)) and not (layer0_outputs(1721));
    outputs(2683) <= (layer0_outputs(2496)) and (layer0_outputs(1753));
    outputs(2684) <= not(layer0_outputs(3721));
    outputs(2685) <= not(layer0_outputs(4700)) or (layer0_outputs(5048));
    outputs(2686) <= (layer0_outputs(4044)) xor (layer0_outputs(1728));
    outputs(2687) <= not(layer0_outputs(387));
    outputs(2688) <= not((layer0_outputs(676)) xor (layer0_outputs(3758)));
    outputs(2689) <= (layer0_outputs(3468)) xor (layer0_outputs(4672));
    outputs(2690) <= not(layer0_outputs(1841));
    outputs(2691) <= not(layer0_outputs(4034)) or (layer0_outputs(2146));
    outputs(2692) <= not(layer0_outputs(3938));
    outputs(2693) <= not((layer0_outputs(3418)) and (layer0_outputs(3190)));
    outputs(2694) <= (layer0_outputs(1244)) and not (layer0_outputs(1714));
    outputs(2695) <= layer0_outputs(2315);
    outputs(2696) <= not(layer0_outputs(541));
    outputs(2697) <= not((layer0_outputs(203)) or (layer0_outputs(1950)));
    outputs(2698) <= not(layer0_outputs(2493));
    outputs(2699) <= (layer0_outputs(2780)) xor (layer0_outputs(4915));
    outputs(2700) <= not(layer0_outputs(3201));
    outputs(2701) <= not(layer0_outputs(696));
    outputs(2702) <= not(layer0_outputs(1379));
    outputs(2703) <= layer0_outputs(3467);
    outputs(2704) <= (layer0_outputs(1602)) xor (layer0_outputs(270));
    outputs(2705) <= (layer0_outputs(1073)) and not (layer0_outputs(1944));
    outputs(2706) <= not((layer0_outputs(3900)) xor (layer0_outputs(4472)));
    outputs(2707) <= layer0_outputs(2357);
    outputs(2708) <= not((layer0_outputs(3131)) or (layer0_outputs(2698)));
    outputs(2709) <= not((layer0_outputs(1900)) xor (layer0_outputs(3054)));
    outputs(2710) <= not((layer0_outputs(2617)) xor (layer0_outputs(2886)));
    outputs(2711) <= layer0_outputs(4925);
    outputs(2712) <= not(layer0_outputs(1909));
    outputs(2713) <= not(layer0_outputs(2688));
    outputs(2714) <= layer0_outputs(4252);
    outputs(2715) <= (layer0_outputs(1632)) and not (layer0_outputs(5060));
    outputs(2716) <= not((layer0_outputs(4419)) xor (layer0_outputs(5029)));
    outputs(2717) <= (layer0_outputs(879)) and not (layer0_outputs(1205));
    outputs(2718) <= not((layer0_outputs(4871)) xor (layer0_outputs(2000)));
    outputs(2719) <= not(layer0_outputs(2509));
    outputs(2720) <= not(layer0_outputs(663));
    outputs(2721) <= not(layer0_outputs(4488));
    outputs(2722) <= (layer0_outputs(5112)) and not (layer0_outputs(11));
    outputs(2723) <= (layer0_outputs(932)) xor (layer0_outputs(246));
    outputs(2724) <= (layer0_outputs(4905)) and not (layer0_outputs(1663));
    outputs(2725) <= not((layer0_outputs(2888)) or (layer0_outputs(631)));
    outputs(2726) <= layer0_outputs(1945);
    outputs(2727) <= not((layer0_outputs(1496)) xor (layer0_outputs(4665)));
    outputs(2728) <= not((layer0_outputs(744)) xor (layer0_outputs(3949)));
    outputs(2729) <= not(layer0_outputs(4668));
    outputs(2730) <= not(layer0_outputs(2280));
    outputs(2731) <= not(layer0_outputs(3960));
    outputs(2732) <= layer0_outputs(2375);
    outputs(2733) <= (layer0_outputs(1032)) and not (layer0_outputs(1767));
    outputs(2734) <= not(layer0_outputs(264));
    outputs(2735) <= (layer0_outputs(2471)) and not (layer0_outputs(3635));
    outputs(2736) <= layer0_outputs(2790);
    outputs(2737) <= not(layer0_outputs(3158)) or (layer0_outputs(4549));
    outputs(2738) <= not(layer0_outputs(1613)) or (layer0_outputs(3492));
    outputs(2739) <= not(layer0_outputs(3647));
    outputs(2740) <= (layer0_outputs(2308)) xor (layer0_outputs(2500));
    outputs(2741) <= layer0_outputs(3911);
    outputs(2742) <= not(layer0_outputs(3840));
    outputs(2743) <= not((layer0_outputs(105)) xor (layer0_outputs(169)));
    outputs(2744) <= not(layer0_outputs(2022));
    outputs(2745) <= (layer0_outputs(4807)) and (layer0_outputs(702));
    outputs(2746) <= not(layer0_outputs(5027));
    outputs(2747) <= (layer0_outputs(4547)) and not (layer0_outputs(2957));
    outputs(2748) <= not((layer0_outputs(885)) xor (layer0_outputs(4287)));
    outputs(2749) <= layer0_outputs(4237);
    outputs(2750) <= layer0_outputs(1243);
    outputs(2751) <= not(layer0_outputs(4185));
    outputs(2752) <= (layer0_outputs(877)) and (layer0_outputs(1967));
    outputs(2753) <= layer0_outputs(2876);
    outputs(2754) <= not((layer0_outputs(798)) xor (layer0_outputs(1480)));
    outputs(2755) <= not(layer0_outputs(3557));
    outputs(2756) <= (layer0_outputs(2163)) and (layer0_outputs(1225));
    outputs(2757) <= not(layer0_outputs(1191));
    outputs(2758) <= not(layer0_outputs(2011)) or (layer0_outputs(2640));
    outputs(2759) <= not(layer0_outputs(2382));
    outputs(2760) <= (layer0_outputs(5054)) and not (layer0_outputs(116));
    outputs(2761) <= not(layer0_outputs(2406));
    outputs(2762) <= layer0_outputs(73);
    outputs(2763) <= (layer0_outputs(17)) and (layer0_outputs(141));
    outputs(2764) <= not(layer0_outputs(355)) or (layer0_outputs(4588));
    outputs(2765) <= layer0_outputs(1056);
    outputs(2766) <= layer0_outputs(1736);
    outputs(2767) <= (layer0_outputs(358)) and not (layer0_outputs(2719));
    outputs(2768) <= not(layer0_outputs(2539));
    outputs(2769) <= not(layer0_outputs(4768));
    outputs(2770) <= not((layer0_outputs(4361)) xor (layer0_outputs(2958)));
    outputs(2771) <= layer0_outputs(4421);
    outputs(2772) <= layer0_outputs(3264);
    outputs(2773) <= layer0_outputs(3152);
    outputs(2774) <= (layer0_outputs(3313)) and (layer0_outputs(13));
    outputs(2775) <= (layer0_outputs(132)) and (layer0_outputs(4011));
    outputs(2776) <= (layer0_outputs(934)) and not (layer0_outputs(1867));
    outputs(2777) <= not(layer0_outputs(741));
    outputs(2778) <= layer0_outputs(1908);
    outputs(2779) <= not(layer0_outputs(4427)) or (layer0_outputs(4099));
    outputs(2780) <= (layer0_outputs(5054)) xor (layer0_outputs(2811));
    outputs(2781) <= not((layer0_outputs(1798)) xor (layer0_outputs(1300)));
    outputs(2782) <= not(layer0_outputs(4676));
    outputs(2783) <= layer0_outputs(1364);
    outputs(2784) <= (layer0_outputs(600)) or (layer0_outputs(2557));
    outputs(2785) <= (layer0_outputs(4146)) and not (layer0_outputs(42));
    outputs(2786) <= not((layer0_outputs(335)) or (layer0_outputs(3097)));
    outputs(2787) <= (layer0_outputs(1635)) and not (layer0_outputs(646));
    outputs(2788) <= (layer0_outputs(4054)) xor (layer0_outputs(351));
    outputs(2789) <= not((layer0_outputs(2795)) xor (layer0_outputs(219)));
    outputs(2790) <= layer0_outputs(3270);
    outputs(2791) <= (layer0_outputs(3843)) and not (layer0_outputs(3466));
    outputs(2792) <= (layer0_outputs(4208)) xor (layer0_outputs(1854));
    outputs(2793) <= layer0_outputs(165);
    outputs(2794) <= not((layer0_outputs(3193)) or (layer0_outputs(862)));
    outputs(2795) <= layer0_outputs(2027);
    outputs(2796) <= (layer0_outputs(3906)) and (layer0_outputs(2155));
    outputs(2797) <= (layer0_outputs(641)) xor (layer0_outputs(4720));
    outputs(2798) <= (layer0_outputs(4884)) xor (layer0_outputs(5056));
    outputs(2799) <= not((layer0_outputs(486)) xor (layer0_outputs(4075)));
    outputs(2800) <= (layer0_outputs(465)) xor (layer0_outputs(1877));
    outputs(2801) <= (layer0_outputs(4120)) or (layer0_outputs(2069));
    outputs(2802) <= not(layer0_outputs(2540)) or (layer0_outputs(3300));
    outputs(2803) <= not((layer0_outputs(4567)) xor (layer0_outputs(3323)));
    outputs(2804) <= not(layer0_outputs(2280)) or (layer0_outputs(3500));
    outputs(2805) <= layer0_outputs(1560);
    outputs(2806) <= not((layer0_outputs(4695)) xor (layer0_outputs(1583)));
    outputs(2807) <= not(layer0_outputs(4160));
    outputs(2808) <= layer0_outputs(1266);
    outputs(2809) <= layer0_outputs(2808);
    outputs(2810) <= (layer0_outputs(4069)) xor (layer0_outputs(3957));
    outputs(2811) <= layer0_outputs(2889);
    outputs(2812) <= layer0_outputs(3372);
    outputs(2813) <= not(layer0_outputs(26));
    outputs(2814) <= not(layer0_outputs(1217));
    outputs(2815) <= not(layer0_outputs(1580)) or (layer0_outputs(2517));
    outputs(2816) <= not((layer0_outputs(2402)) xor (layer0_outputs(2482)));
    outputs(2817) <= not(layer0_outputs(463));
    outputs(2818) <= layer0_outputs(1920);
    outputs(2819) <= not(layer0_outputs(1897));
    outputs(2820) <= not(layer0_outputs(4255));
    outputs(2821) <= not((layer0_outputs(3550)) and (layer0_outputs(1696)));
    outputs(2822) <= not(layer0_outputs(2337));
    outputs(2823) <= not(layer0_outputs(2845));
    outputs(2824) <= not((layer0_outputs(821)) xor (layer0_outputs(3499)));
    outputs(2825) <= (layer0_outputs(3228)) xor (layer0_outputs(3391));
    outputs(2826) <= layer0_outputs(2667);
    outputs(2827) <= not((layer0_outputs(2962)) or (layer0_outputs(1769)));
    outputs(2828) <= layer0_outputs(373);
    outputs(2829) <= not(layer0_outputs(3117)) or (layer0_outputs(1455));
    outputs(2830) <= not(layer0_outputs(1489));
    outputs(2831) <= (layer0_outputs(1351)) and not (layer0_outputs(3678));
    outputs(2832) <= layer0_outputs(3068);
    outputs(2833) <= (layer0_outputs(2216)) and not (layer0_outputs(4963));
    outputs(2834) <= (layer0_outputs(3616)) and not (layer0_outputs(2901));
    outputs(2835) <= layer0_outputs(711);
    outputs(2836) <= not((layer0_outputs(1836)) or (layer0_outputs(919)));
    outputs(2837) <= not((layer0_outputs(4715)) or (layer0_outputs(2047)));
    outputs(2838) <= layer0_outputs(3519);
    outputs(2839) <= (layer0_outputs(3610)) xor (layer0_outputs(1373));
    outputs(2840) <= not((layer0_outputs(2389)) or (layer0_outputs(2292)));
    outputs(2841) <= not(layer0_outputs(1696));
    outputs(2842) <= not((layer0_outputs(1271)) xor (layer0_outputs(1284)));
    outputs(2843) <= (layer0_outputs(1916)) xor (layer0_outputs(3687));
    outputs(2844) <= not(layer0_outputs(4894));
    outputs(2845) <= not(layer0_outputs(434));
    outputs(2846) <= not(layer0_outputs(1772));
    outputs(2847) <= not(layer0_outputs(4888)) or (layer0_outputs(25));
    outputs(2848) <= (layer0_outputs(4068)) and not (layer0_outputs(4916));
    outputs(2849) <= not(layer0_outputs(3909));
    outputs(2850) <= not(layer0_outputs(1794));
    outputs(2851) <= not(layer0_outputs(2838));
    outputs(2852) <= (layer0_outputs(3368)) and not (layer0_outputs(1269));
    outputs(2853) <= not((layer0_outputs(3091)) or (layer0_outputs(305)));
    outputs(2854) <= not((layer0_outputs(1762)) xor (layer0_outputs(16)));
    outputs(2855) <= not(layer0_outputs(1337));
    outputs(2856) <= (layer0_outputs(1715)) xor (layer0_outputs(2170));
    outputs(2857) <= not(layer0_outputs(2035)) or (layer0_outputs(4776));
    outputs(2858) <= (layer0_outputs(1639)) xor (layer0_outputs(3844));
    outputs(2859) <= layer0_outputs(4331);
    outputs(2860) <= (layer0_outputs(4359)) and (layer0_outputs(1120));
    outputs(2861) <= (layer0_outputs(2892)) and not (layer0_outputs(1114));
    outputs(2862) <= not(layer0_outputs(4354));
    outputs(2863) <= not(layer0_outputs(1844));
    outputs(2864) <= not(layer0_outputs(3281));
    outputs(2865) <= not((layer0_outputs(308)) or (layer0_outputs(2451)));
    outputs(2866) <= layer0_outputs(4527);
    outputs(2867) <= (layer0_outputs(344)) and not (layer0_outputs(1759));
    outputs(2868) <= layer0_outputs(987);
    outputs(2869) <= (layer0_outputs(2865)) and (layer0_outputs(2891));
    outputs(2870) <= (layer0_outputs(1203)) and (layer0_outputs(346));
    outputs(2871) <= layer0_outputs(3250);
    outputs(2872) <= not(layer0_outputs(5045));
    outputs(2873) <= layer0_outputs(49);
    outputs(2874) <= (layer0_outputs(1576)) and not (layer0_outputs(3613));
    outputs(2875) <= not(layer0_outputs(3036));
    outputs(2876) <= not(layer0_outputs(2085));
    outputs(2877) <= (layer0_outputs(3261)) and not (layer0_outputs(1275));
    outputs(2878) <= layer0_outputs(334);
    outputs(2879) <= layer0_outputs(4338);
    outputs(2880) <= not((layer0_outputs(1673)) or (layer0_outputs(2346)));
    outputs(2881) <= not((layer0_outputs(5042)) or (layer0_outputs(4024)));
    outputs(2882) <= layer0_outputs(1561);
    outputs(2883) <= not(layer0_outputs(2278));
    outputs(2884) <= layer0_outputs(3010);
    outputs(2885) <= not(layer0_outputs(2306)) or (layer0_outputs(4773));
    outputs(2886) <= (layer0_outputs(770)) xor (layer0_outputs(1814));
    outputs(2887) <= not((layer0_outputs(2433)) and (layer0_outputs(4379)));
    outputs(2888) <= not((layer0_outputs(4851)) xor (layer0_outputs(414)));
    outputs(2889) <= layer0_outputs(956);
    outputs(2890) <= layer0_outputs(1411);
    outputs(2891) <= not((layer0_outputs(2691)) or (layer0_outputs(4778)));
    outputs(2892) <= not(layer0_outputs(296));
    outputs(2893) <= not((layer0_outputs(1134)) and (layer0_outputs(1338)));
    outputs(2894) <= (layer0_outputs(210)) and not (layer0_outputs(3583));
    outputs(2895) <= not(layer0_outputs(1716));
    outputs(2896) <= (layer0_outputs(3472)) xor (layer0_outputs(2773));
    outputs(2897) <= (layer0_outputs(4340)) xor (layer0_outputs(2921));
    outputs(2898) <= (layer0_outputs(4261)) xor (layer0_outputs(5108));
    outputs(2899) <= not(layer0_outputs(1873));
    outputs(2900) <= (layer0_outputs(735)) and not (layer0_outputs(4590));
    outputs(2901) <= layer0_outputs(329);
    outputs(2902) <= layer0_outputs(2188);
    outputs(2903) <= not(layer0_outputs(1634));
    outputs(2904) <= layer0_outputs(4353);
    outputs(2905) <= not(layer0_outputs(2710));
    outputs(2906) <= not(layer0_outputs(2921));
    outputs(2907) <= not((layer0_outputs(3660)) and (layer0_outputs(4451)));
    outputs(2908) <= (layer0_outputs(3331)) or (layer0_outputs(1573));
    outputs(2909) <= not(layer0_outputs(1654));
    outputs(2910) <= (layer0_outputs(1422)) and (layer0_outputs(1883));
    outputs(2911) <= layer0_outputs(1561);
    outputs(2912) <= not((layer0_outputs(495)) or (layer0_outputs(3283)));
    outputs(2913) <= not(layer0_outputs(453));
    outputs(2914) <= not((layer0_outputs(4159)) xor (layer0_outputs(1502)));
    outputs(2915) <= (layer0_outputs(1282)) xor (layer0_outputs(4231));
    outputs(2916) <= not(layer0_outputs(1358));
    outputs(2917) <= layer0_outputs(123);
    outputs(2918) <= not((layer0_outputs(3908)) xor (layer0_outputs(3652)));
    outputs(2919) <= layer0_outputs(3873);
    outputs(2920) <= layer0_outputs(4391);
    outputs(2921) <= (layer0_outputs(411)) xor (layer0_outputs(11));
    outputs(2922) <= not((layer0_outputs(3553)) or (layer0_outputs(1308)));
    outputs(2923) <= (layer0_outputs(1367)) and not (layer0_outputs(4543));
    outputs(2924) <= layer0_outputs(4421);
    outputs(2925) <= not(layer0_outputs(1334)) or (layer0_outputs(2858));
    outputs(2926) <= not((layer0_outputs(218)) xor (layer0_outputs(1874)));
    outputs(2927) <= layer0_outputs(861);
    outputs(2928) <= not((layer0_outputs(678)) xor (layer0_outputs(5066)));
    outputs(2929) <= not((layer0_outputs(3304)) xor (layer0_outputs(2906)));
    outputs(2930) <= (layer0_outputs(4829)) and not (layer0_outputs(1172));
    outputs(2931) <= layer0_outputs(2466);
    outputs(2932) <= not((layer0_outputs(4132)) xor (layer0_outputs(824)));
    outputs(2933) <= not(layer0_outputs(458)) or (layer0_outputs(2049));
    outputs(2934) <= not((layer0_outputs(1957)) xor (layer0_outputs(3782)));
    outputs(2935) <= layer0_outputs(4396);
    outputs(2936) <= not((layer0_outputs(2944)) xor (layer0_outputs(2373)));
    outputs(2937) <= layer0_outputs(4215);
    outputs(2938) <= layer0_outputs(1493);
    outputs(2939) <= not((layer0_outputs(860)) xor (layer0_outputs(3119)));
    outputs(2940) <= (layer0_outputs(1670)) and (layer0_outputs(777));
    outputs(2941) <= not(layer0_outputs(523)) or (layer0_outputs(4133));
    outputs(2942) <= (layer0_outputs(3110)) and not (layer0_outputs(3859));
    outputs(2943) <= (layer0_outputs(928)) and not (layer0_outputs(1286));
    outputs(2944) <= not(layer0_outputs(1036));
    outputs(2945) <= (layer0_outputs(266)) or (layer0_outputs(450));
    outputs(2946) <= not((layer0_outputs(126)) and (layer0_outputs(1035)));
    outputs(2947) <= (layer0_outputs(312)) or (layer0_outputs(1021));
    outputs(2948) <= not(layer0_outputs(4045));
    outputs(2949) <= layer0_outputs(3766);
    outputs(2950) <= (layer0_outputs(601)) xor (layer0_outputs(5061));
    outputs(2951) <= not(layer0_outputs(730));
    outputs(2952) <= (layer0_outputs(3215)) and (layer0_outputs(1123));
    outputs(2953) <= (layer0_outputs(262)) and not (layer0_outputs(2030));
    outputs(2954) <= not((layer0_outputs(4265)) xor (layer0_outputs(1224)));
    outputs(2955) <= not(layer0_outputs(3764));
    outputs(2956) <= (layer0_outputs(492)) xor (layer0_outputs(1405));
    outputs(2957) <= not((layer0_outputs(2119)) and (layer0_outputs(3299)));
    outputs(2958) <= not((layer0_outputs(4668)) or (layer0_outputs(1651)));
    outputs(2959) <= layer0_outputs(4999);
    outputs(2960) <= layer0_outputs(2388);
    outputs(2961) <= not(layer0_outputs(2539));
    outputs(2962) <= not((layer0_outputs(4985)) xor (layer0_outputs(4922)));
    outputs(2963) <= (layer0_outputs(1612)) xor (layer0_outputs(399));
    outputs(2964) <= (layer0_outputs(3809)) and not (layer0_outputs(2497));
    outputs(2965) <= (layer0_outputs(3615)) and (layer0_outputs(4270));
    outputs(2966) <= layer0_outputs(2275);
    outputs(2967) <= not(layer0_outputs(4623)) or (layer0_outputs(2889));
    outputs(2968) <= not((layer0_outputs(4896)) xor (layer0_outputs(3130)));
    outputs(2969) <= not((layer0_outputs(64)) xor (layer0_outputs(4792)));
    outputs(2970) <= layer0_outputs(4135);
    outputs(2971) <= layer0_outputs(284);
    outputs(2972) <= layer0_outputs(1420);
    outputs(2973) <= not(layer0_outputs(3725));
    outputs(2974) <= (layer0_outputs(575)) xor (layer0_outputs(1384));
    outputs(2975) <= layer0_outputs(1717);
    outputs(2976) <= layer0_outputs(4284);
    outputs(2977) <= (layer0_outputs(2527)) and not (layer0_outputs(1863));
    outputs(2978) <= not((layer0_outputs(3269)) or (layer0_outputs(4229)));
    outputs(2979) <= not(layer0_outputs(847));
    outputs(2980) <= not((layer0_outputs(3443)) and (layer0_outputs(1564)));
    outputs(2981) <= (layer0_outputs(4625)) and (layer0_outputs(4425));
    outputs(2982) <= layer0_outputs(4133);
    outputs(2983) <= not((layer0_outputs(2264)) xor (layer0_outputs(1952)));
    outputs(2984) <= layer0_outputs(5062);
    outputs(2985) <= (layer0_outputs(1331)) xor (layer0_outputs(4831));
    outputs(2986) <= not((layer0_outputs(1805)) or (layer0_outputs(3784)));
    outputs(2987) <= not(layer0_outputs(1964));
    outputs(2988) <= (layer0_outputs(4117)) xor (layer0_outputs(4009));
    outputs(2989) <= not(layer0_outputs(3744));
    outputs(2990) <= not(layer0_outputs(532)) or (layer0_outputs(1681));
    outputs(2991) <= layer0_outputs(4330);
    outputs(2992) <= not(layer0_outputs(2546));
    outputs(2993) <= not(layer0_outputs(653));
    outputs(2994) <= not((layer0_outputs(3069)) xor (layer0_outputs(676)));
    outputs(2995) <= not(layer0_outputs(3198));
    outputs(2996) <= not((layer0_outputs(3103)) xor (layer0_outputs(4304)));
    outputs(2997) <= not(layer0_outputs(2297)) or (layer0_outputs(4725));
    outputs(2998) <= (layer0_outputs(356)) xor (layer0_outputs(2328));
    outputs(2999) <= (layer0_outputs(65)) xor (layer0_outputs(2422));
    outputs(3000) <= layer0_outputs(3639);
    outputs(3001) <= layer0_outputs(3130);
    outputs(3002) <= layer0_outputs(4688);
    outputs(3003) <= (layer0_outputs(4210)) and not (layer0_outputs(3945));
    outputs(3004) <= layer0_outputs(4795);
    outputs(3005) <= layer0_outputs(4757);
    outputs(3006) <= layer0_outputs(1052);
    outputs(3007) <= (layer0_outputs(4661)) xor (layer0_outputs(3825));
    outputs(3008) <= not(layer0_outputs(2764));
    outputs(3009) <= not((layer0_outputs(539)) and (layer0_outputs(2732)));
    outputs(3010) <= not((layer0_outputs(134)) xor (layer0_outputs(4813)));
    outputs(3011) <= (layer0_outputs(2990)) and (layer0_outputs(1687));
    outputs(3012) <= not(layer0_outputs(4407));
    outputs(3013) <= layer0_outputs(2744);
    outputs(3014) <= not(layer0_outputs(3755));
    outputs(3015) <= (layer0_outputs(3296)) and not (layer0_outputs(133));
    outputs(3016) <= not(layer0_outputs(773));
    outputs(3017) <= not(layer0_outputs(1470));
    outputs(3018) <= not((layer0_outputs(382)) or (layer0_outputs(1170)));
    outputs(3019) <= not((layer0_outputs(4687)) xor (layer0_outputs(2712)));
    outputs(3020) <= layer0_outputs(2674);
    outputs(3021) <= not(layer0_outputs(3156));
    outputs(3022) <= not(layer0_outputs(3708));
    outputs(3023) <= layer0_outputs(3533);
    outputs(3024) <= not((layer0_outputs(4301)) xor (layer0_outputs(1701)));
    outputs(3025) <= not(layer0_outputs(1124));
    outputs(3026) <= not((layer0_outputs(3886)) or (layer0_outputs(4245)));
    outputs(3027) <= not((layer0_outputs(4797)) xor (layer0_outputs(1647)));
    outputs(3028) <= not((layer0_outputs(1504)) xor (layer0_outputs(89)));
    outputs(3029) <= (layer0_outputs(416)) and not (layer0_outputs(4317));
    outputs(3030) <= layer0_outputs(3185);
    outputs(3031) <= not(layer0_outputs(794));
    outputs(3032) <= not(layer0_outputs(2304));
    outputs(3033) <= (layer0_outputs(1045)) xor (layer0_outputs(252));
    outputs(3034) <= layer0_outputs(3215);
    outputs(3035) <= not(layer0_outputs(4924));
    outputs(3036) <= layer0_outputs(2635);
    outputs(3037) <= (layer0_outputs(560)) xor (layer0_outputs(1538));
    outputs(3038) <= layer0_outputs(593);
    outputs(3039) <= not(layer0_outputs(769));
    outputs(3040) <= not((layer0_outputs(1183)) xor (layer0_outputs(3362)));
    outputs(3041) <= not(layer0_outputs(4705));
    outputs(3042) <= not((layer0_outputs(4551)) or (layer0_outputs(4105)));
    outputs(3043) <= layer0_outputs(4398);
    outputs(3044) <= (layer0_outputs(4144)) xor (layer0_outputs(4204));
    outputs(3045) <= not(layer0_outputs(3723)) or (layer0_outputs(4154));
    outputs(3046) <= not(layer0_outputs(651));
    outputs(3047) <= not((layer0_outputs(5092)) or (layer0_outputs(196)));
    outputs(3048) <= layer0_outputs(4886);
    outputs(3049) <= (layer0_outputs(300)) xor (layer0_outputs(3593));
    outputs(3050) <= not(layer0_outputs(19));
    outputs(3051) <= not(layer0_outputs(2185)) or (layer0_outputs(4221));
    outputs(3052) <= (layer0_outputs(4625)) and not (layer0_outputs(2762));
    outputs(3053) <= layer0_outputs(1019);
    outputs(3054) <= (layer0_outputs(167)) xor (layer0_outputs(2121));
    outputs(3055) <= (layer0_outputs(4438)) or (layer0_outputs(2855));
    outputs(3056) <= not(layer0_outputs(2968));
    outputs(3057) <= not(layer0_outputs(2872));
    outputs(3058) <= layer0_outputs(4423);
    outputs(3059) <= (layer0_outputs(4960)) xor (layer0_outputs(258));
    outputs(3060) <= (layer0_outputs(1047)) xor (layer0_outputs(1885));
    outputs(3061) <= not(layer0_outputs(3647));
    outputs(3062) <= not(layer0_outputs(4930)) or (layer0_outputs(88));
    outputs(3063) <= not(layer0_outputs(1604));
    outputs(3064) <= not((layer0_outputs(3278)) or (layer0_outputs(4902)));
    outputs(3065) <= not((layer0_outputs(5077)) xor (layer0_outputs(289)));
    outputs(3066) <= layer0_outputs(3157);
    outputs(3067) <= not(layer0_outputs(4341));
    outputs(3068) <= (layer0_outputs(3226)) and (layer0_outputs(2596));
    outputs(3069) <= (layer0_outputs(1294)) xor (layer0_outputs(474));
    outputs(3070) <= not(layer0_outputs(1956));
    outputs(3071) <= not(layer0_outputs(3411));
    outputs(3072) <= (layer0_outputs(1353)) and (layer0_outputs(99));
    outputs(3073) <= not(layer0_outputs(4824));
    outputs(3074) <= (layer0_outputs(4663)) or (layer0_outputs(4997));
    outputs(3075) <= layer0_outputs(2593);
    outputs(3076) <= not(layer0_outputs(3394));
    outputs(3077) <= layer0_outputs(2227);
    outputs(3078) <= not((layer0_outputs(3988)) xor (layer0_outputs(851)));
    outputs(3079) <= not((layer0_outputs(4767)) or (layer0_outputs(4689)));
    outputs(3080) <= not(layer0_outputs(1560));
    outputs(3081) <= not((layer0_outputs(4740)) or (layer0_outputs(4958)));
    outputs(3082) <= not((layer0_outputs(1618)) or (layer0_outputs(2580)));
    outputs(3083) <= not((layer0_outputs(2041)) xor (layer0_outputs(1234)));
    outputs(3084) <= not(layer0_outputs(3670));
    outputs(3085) <= not(layer0_outputs(4095)) or (layer0_outputs(4349));
    outputs(3086) <= not((layer0_outputs(4419)) or (layer0_outputs(3505)));
    outputs(3087) <= not(layer0_outputs(3393));
    outputs(3088) <= not(layer0_outputs(2910));
    outputs(3089) <= layer0_outputs(1883);
    outputs(3090) <= not(layer0_outputs(726)) or (layer0_outputs(901));
    outputs(3091) <= layer0_outputs(1971);
    outputs(3092) <= layer0_outputs(3204);
    outputs(3093) <= (layer0_outputs(2307)) xor (layer0_outputs(156));
    outputs(3094) <= not(layer0_outputs(221));
    outputs(3095) <= (layer0_outputs(1259)) and (layer0_outputs(4842));
    outputs(3096) <= not(layer0_outputs(1637));
    outputs(3097) <= not(layer0_outputs(3089));
    outputs(3098) <= layer0_outputs(1986);
    outputs(3099) <= not(layer0_outputs(1232));
    outputs(3100) <= layer0_outputs(3276);
    outputs(3101) <= not(layer0_outputs(3918));
    outputs(3102) <= not(layer0_outputs(2897));
    outputs(3103) <= not(layer0_outputs(942));
    outputs(3104) <= (layer0_outputs(1268)) xor (layer0_outputs(2431));
    outputs(3105) <= not(layer0_outputs(1144));
    outputs(3106) <= layer0_outputs(1353);
    outputs(3107) <= not(layer0_outputs(953)) or (layer0_outputs(3945));
    outputs(3108) <= not(layer0_outputs(4875));
    outputs(3109) <= (layer0_outputs(2924)) xor (layer0_outputs(3746));
    outputs(3110) <= (layer0_outputs(1894)) and (layer0_outputs(1478));
    outputs(3111) <= not(layer0_outputs(4932));
    outputs(3112) <= (layer0_outputs(4505)) or (layer0_outputs(1371));
    outputs(3113) <= not(layer0_outputs(2969));
    outputs(3114) <= not((layer0_outputs(1713)) or (layer0_outputs(2983)));
    outputs(3115) <= layer0_outputs(127);
    outputs(3116) <= (layer0_outputs(2469)) and not (layer0_outputs(4484));
    outputs(3117) <= layer0_outputs(1822);
    outputs(3118) <= layer0_outputs(206);
    outputs(3119) <= not((layer0_outputs(1340)) or (layer0_outputs(3481)));
    outputs(3120) <= layer0_outputs(3874);
    outputs(3121) <= not(layer0_outputs(3596));
    outputs(3122) <= not((layer0_outputs(1494)) or (layer0_outputs(3462)));
    outputs(3123) <= (layer0_outputs(3944)) and not (layer0_outputs(2481));
    outputs(3124) <= layer0_outputs(4403);
    outputs(3125) <= not(layer0_outputs(1202)) or (layer0_outputs(4080));
    outputs(3126) <= layer0_outputs(1421);
    outputs(3127) <= layer0_outputs(4956);
    outputs(3128) <= (layer0_outputs(2125)) or (layer0_outputs(3759));
    outputs(3129) <= layer0_outputs(2449);
    outputs(3130) <= layer0_outputs(2560);
    outputs(3131) <= (layer0_outputs(2578)) xor (layer0_outputs(3582));
    outputs(3132) <= layer0_outputs(1265);
    outputs(3133) <= layer0_outputs(599);
    outputs(3134) <= (layer0_outputs(3807)) and (layer0_outputs(4796));
    outputs(3135) <= not(layer0_outputs(3118));
    outputs(3136) <= not((layer0_outputs(1568)) xor (layer0_outputs(4049)));
    outputs(3137) <= not(layer0_outputs(893));
    outputs(3138) <= layer0_outputs(4629);
    outputs(3139) <= (layer0_outputs(3691)) and not (layer0_outputs(4015));
    outputs(3140) <= not(layer0_outputs(4912));
    outputs(3141) <= (layer0_outputs(2825)) and not (layer0_outputs(858));
    outputs(3142) <= not(layer0_outputs(3824));
    outputs(3143) <= not(layer0_outputs(81));
    outputs(3144) <= not(layer0_outputs(317));
    outputs(3145) <= not((layer0_outputs(4369)) or (layer0_outputs(2078)));
    outputs(3146) <= layer0_outputs(4081);
    outputs(3147) <= layer0_outputs(77);
    outputs(3148) <= (layer0_outputs(2087)) and not (layer0_outputs(4003));
    outputs(3149) <= layer0_outputs(3237);
    outputs(3150) <= not(layer0_outputs(3155));
    outputs(3151) <= layer0_outputs(2395);
    outputs(3152) <= (layer0_outputs(637)) and not (layer0_outputs(1308));
    outputs(3153) <= layer0_outputs(250);
    outputs(3154) <= layer0_outputs(857);
    outputs(3155) <= layer0_outputs(5001);
    outputs(3156) <= (layer0_outputs(805)) and not (layer0_outputs(3100));
    outputs(3157) <= layer0_outputs(2658);
    outputs(3158) <= not(layer0_outputs(5103));
    outputs(3159) <= not((layer0_outputs(4266)) or (layer0_outputs(3730)));
    outputs(3160) <= not(layer0_outputs(4704)) or (layer0_outputs(2452));
    outputs(3161) <= not((layer0_outputs(3239)) or (layer0_outputs(3998)));
    outputs(3162) <= layer0_outputs(1540);
    outputs(3163) <= not((layer0_outputs(1982)) xor (layer0_outputs(3135)));
    outputs(3164) <= not((layer0_outputs(1350)) or (layer0_outputs(3698)));
    outputs(3165) <= not(layer0_outputs(2988));
    outputs(3166) <= (layer0_outputs(227)) and not (layer0_outputs(5035));
    outputs(3167) <= layer0_outputs(3512);
    outputs(3168) <= not(layer0_outputs(2516));
    outputs(3169) <= layer0_outputs(2002);
    outputs(3170) <= (layer0_outputs(3894)) and (layer0_outputs(4525));
    outputs(3171) <= (layer0_outputs(1328)) and (layer0_outputs(1631));
    outputs(3172) <= not((layer0_outputs(1926)) xor (layer0_outputs(1201)));
    outputs(3173) <= (layer0_outputs(1276)) and not (layer0_outputs(3976));
    outputs(3174) <= layer0_outputs(4649);
    outputs(3175) <= layer0_outputs(1129);
    outputs(3176) <= (layer0_outputs(2631)) xor (layer0_outputs(3157));
    outputs(3177) <= layer0_outputs(2943);
    outputs(3178) <= not(layer0_outputs(2766));
    outputs(3179) <= not((layer0_outputs(3202)) or (layer0_outputs(761)));
    outputs(3180) <= not((layer0_outputs(4247)) or (layer0_outputs(2843)));
    outputs(3181) <= (layer0_outputs(2440)) and not (layer0_outputs(4413));
    outputs(3182) <= not(layer0_outputs(2111));
    outputs(3183) <= layer0_outputs(4741);
    outputs(3184) <= not((layer0_outputs(5019)) and (layer0_outputs(2604)));
    outputs(3185) <= not(layer0_outputs(2497));
    outputs(3186) <= layer0_outputs(3125);
    outputs(3187) <= layer0_outputs(1394);
    outputs(3188) <= layer0_outputs(775);
    outputs(3189) <= not(layer0_outputs(5072));
    outputs(3190) <= not(layer0_outputs(4800));
    outputs(3191) <= (layer0_outputs(1937)) xor (layer0_outputs(1850));
    outputs(3192) <= not(layer0_outputs(4299));
    outputs(3193) <= not(layer0_outputs(3249));
    outputs(3194) <= not((layer0_outputs(3031)) xor (layer0_outputs(5056)));
    outputs(3195) <= not((layer0_outputs(4021)) or (layer0_outputs(3623)));
    outputs(3196) <= not(layer0_outputs(4016));
    outputs(3197) <= layer0_outputs(4639);
    outputs(3198) <= layer0_outputs(377);
    outputs(3199) <= layer0_outputs(4177);
    outputs(3200) <= layer0_outputs(1040);
    outputs(3201) <= (layer0_outputs(1988)) and not (layer0_outputs(5103));
    outputs(3202) <= layer0_outputs(4030);
    outputs(3203) <= layer0_outputs(514);
    outputs(3204) <= not(layer0_outputs(517));
    outputs(3205) <= not(layer0_outputs(370)) or (layer0_outputs(72));
    outputs(3206) <= layer0_outputs(1961);
    outputs(3207) <= not(layer0_outputs(3089)) or (layer0_outputs(3635));
    outputs(3208) <= (layer0_outputs(149)) xor (layer0_outputs(1397));
    outputs(3209) <= not(layer0_outputs(1589));
    outputs(3210) <= layer0_outputs(2432);
    outputs(3211) <= layer0_outputs(754);
    outputs(3212) <= not(layer0_outputs(139));
    outputs(3213) <= not(layer0_outputs(963));
    outputs(3214) <= not(layer0_outputs(3011));
    outputs(3215) <= not((layer0_outputs(3458)) xor (layer0_outputs(4976)));
    outputs(3216) <= layer0_outputs(3710);
    outputs(3217) <= layer0_outputs(1102);
    outputs(3218) <= not((layer0_outputs(3253)) xor (layer0_outputs(4529)));
    outputs(3219) <= layer0_outputs(1086);
    outputs(3220) <= (layer0_outputs(3419)) and not (layer0_outputs(1227));
    outputs(3221) <= not(layer0_outputs(1406)) or (layer0_outputs(1013));
    outputs(3222) <= not(layer0_outputs(255));
    outputs(3223) <= not((layer0_outputs(1356)) and (layer0_outputs(810)));
    outputs(3224) <= not((layer0_outputs(4585)) or (layer0_outputs(1064)));
    outputs(3225) <= layer0_outputs(3577);
    outputs(3226) <= not(layer0_outputs(57));
    outputs(3227) <= not((layer0_outputs(2240)) or (layer0_outputs(4273)));
    outputs(3228) <= not(layer0_outputs(3518));
    outputs(3229) <= not((layer0_outputs(3455)) or (layer0_outputs(4402)));
    outputs(3230) <= not((layer0_outputs(4333)) or (layer0_outputs(3699)));
    outputs(3231) <= (layer0_outputs(1436)) xor (layer0_outputs(4853));
    outputs(3232) <= layer0_outputs(3125);
    outputs(3233) <= layer0_outputs(4951);
    outputs(3234) <= (layer0_outputs(4212)) and not (layer0_outputs(3980));
    outputs(3235) <= not((layer0_outputs(2128)) or (layer0_outputs(4643)));
    outputs(3236) <= not((layer0_outputs(4422)) xor (layer0_outputs(2084)));
    outputs(3237) <= (layer0_outputs(2106)) and (layer0_outputs(3220));
    outputs(3238) <= layer0_outputs(4833);
    outputs(3239) <= (layer0_outputs(4984)) and not (layer0_outputs(4706));
    outputs(3240) <= (layer0_outputs(3365)) and not (layer0_outputs(4041));
    outputs(3241) <= (layer0_outputs(993)) and not (layer0_outputs(4641));
    outputs(3242) <= layer0_outputs(1780);
    outputs(3243) <= not(layer0_outputs(746));
    outputs(3244) <= not(layer0_outputs(3957));
    outputs(3245) <= not((layer0_outputs(4126)) xor (layer0_outputs(381)));
    outputs(3246) <= (layer0_outputs(1764)) and (layer0_outputs(864));
    outputs(3247) <= not(layer0_outputs(4885));
    outputs(3248) <= not(layer0_outputs(3821));
    outputs(3249) <= layer0_outputs(1201);
    outputs(3250) <= layer0_outputs(1316);
    outputs(3251) <= not(layer0_outputs(3264));
    outputs(3252) <= layer0_outputs(2776);
    outputs(3253) <= not((layer0_outputs(3079)) and (layer0_outputs(965)));
    outputs(3254) <= layer0_outputs(4535);
    outputs(3255) <= (layer0_outputs(3290)) and not (layer0_outputs(3762));
    outputs(3256) <= layer0_outputs(3688);
    outputs(3257) <= not(layer0_outputs(4));
    outputs(3258) <= (layer0_outputs(1235)) or (layer0_outputs(1804));
    outputs(3259) <= (layer0_outputs(1052)) and not (layer0_outputs(620));
    outputs(3260) <= layer0_outputs(615);
    outputs(3261) <= not(layer0_outputs(4840));
    outputs(3262) <= (layer0_outputs(502)) and (layer0_outputs(4097));
    outputs(3263) <= not((layer0_outputs(1918)) and (layer0_outputs(3303)));
    outputs(3264) <= not(layer0_outputs(3033));
    outputs(3265) <= layer0_outputs(1740);
    outputs(3266) <= layer0_outputs(3021);
    outputs(3267) <= layer0_outputs(4222);
    outputs(3268) <= not((layer0_outputs(1162)) xor (layer0_outputs(2024)));
    outputs(3269) <= not((layer0_outputs(2197)) or (layer0_outputs(2985)));
    outputs(3270) <= (layer0_outputs(184)) and (layer0_outputs(2318));
    outputs(3271) <= not((layer0_outputs(3093)) xor (layer0_outputs(3458)));
    outputs(3272) <= not((layer0_outputs(4978)) or (layer0_outputs(4311)));
    outputs(3273) <= not((layer0_outputs(5049)) or (layer0_outputs(2461)));
    outputs(3274) <= not(layer0_outputs(2595));
    outputs(3275) <= layer0_outputs(1489);
    outputs(3276) <= layer0_outputs(3184);
    outputs(3277) <= not(layer0_outputs(2905));
    outputs(3278) <= not((layer0_outputs(1584)) xor (layer0_outputs(4027)));
    outputs(3279) <= (layer0_outputs(2854)) and not (layer0_outputs(1352));
    outputs(3280) <= layer0_outputs(2338);
    outputs(3281) <= not((layer0_outputs(3357)) xor (layer0_outputs(2592)));
    outputs(3282) <= layer0_outputs(802);
    outputs(3283) <= (layer0_outputs(4167)) and (layer0_outputs(3179));
    outputs(3284) <= layer0_outputs(633);
    outputs(3285) <= not(layer0_outputs(4832));
    outputs(3286) <= not((layer0_outputs(1607)) or (layer0_outputs(3771)));
    outputs(3287) <= not(layer0_outputs(4440));
    outputs(3288) <= layer0_outputs(4660);
    outputs(3289) <= layer0_outputs(3435);
    outputs(3290) <= (layer0_outputs(4262)) and (layer0_outputs(2866));
    outputs(3291) <= (layer0_outputs(2747)) and not (layer0_outputs(2298));
    outputs(3292) <= not(layer0_outputs(421));
    outputs(3293) <= not((layer0_outputs(695)) xor (layer0_outputs(2252)));
    outputs(3294) <= (layer0_outputs(1875)) and not (layer0_outputs(4942));
    outputs(3295) <= (layer0_outputs(3615)) and not (layer0_outputs(3560));
    outputs(3296) <= (layer0_outputs(3450)) or (layer0_outputs(4374));
    outputs(3297) <= (layer0_outputs(236)) xor (layer0_outputs(719));
    outputs(3298) <= (layer0_outputs(143)) and not (layer0_outputs(154));
    outputs(3299) <= (layer0_outputs(1624)) and not (layer0_outputs(4230));
    outputs(3300) <= layer0_outputs(3823);
    outputs(3301) <= layer0_outputs(92);
    outputs(3302) <= (layer0_outputs(3742)) and not (layer0_outputs(150));
    outputs(3303) <= layer0_outputs(3739);
    outputs(3304) <= (layer0_outputs(2798)) and (layer0_outputs(3475));
    outputs(3305) <= (layer0_outputs(4801)) and (layer0_outputs(4682));
    outputs(3306) <= not(layer0_outputs(2353));
    outputs(3307) <= (layer0_outputs(760)) and (layer0_outputs(2102));
    outputs(3308) <= (layer0_outputs(4139)) and not (layer0_outputs(199));
    outputs(3309) <= not(layer0_outputs(3728));
    outputs(3310) <= layer0_outputs(4870);
    outputs(3311) <= layer0_outputs(2837);
    outputs(3312) <= not(layer0_outputs(1335));
    outputs(3313) <= not(layer0_outputs(1459));
    outputs(3314) <= not(layer0_outputs(4412));
    outputs(3315) <= not(layer0_outputs(1126)) or (layer0_outputs(524));
    outputs(3316) <= not((layer0_outputs(3182)) xor (layer0_outputs(5057)));
    outputs(3317) <= not(layer0_outputs(299)) or (layer0_outputs(4225));
    outputs(3318) <= not(layer0_outputs(2571));
    outputs(3319) <= layer0_outputs(4933);
    outputs(3320) <= not(layer0_outputs(4782));
    outputs(3321) <= layer0_outputs(4131);
    outputs(3322) <= layer0_outputs(3205);
    outputs(3323) <= (layer0_outputs(4019)) and (layer0_outputs(3690));
    outputs(3324) <= layer0_outputs(4772);
    outputs(3325) <= not(layer0_outputs(1912)) or (layer0_outputs(266));
    outputs(3326) <= (layer0_outputs(561)) and not (layer0_outputs(4163));
    outputs(3327) <= (layer0_outputs(2847)) and (layer0_outputs(4578));
    outputs(3328) <= layer0_outputs(3896);
    outputs(3329) <= layer0_outputs(1657);
    outputs(3330) <= (layer0_outputs(2009)) xor (layer0_outputs(3552));
    outputs(3331) <= not((layer0_outputs(2928)) xor (layer0_outputs(1432)));
    outputs(3332) <= (layer0_outputs(4821)) and (layer0_outputs(4649));
    outputs(3333) <= (layer0_outputs(2258)) and (layer0_outputs(4961));
    outputs(3334) <= (layer0_outputs(4240)) or (layer0_outputs(533));
    outputs(3335) <= layer0_outputs(2220);
    outputs(3336) <= layer0_outputs(1423);
    outputs(3337) <= layer0_outputs(3885);
    outputs(3338) <= (layer0_outputs(395)) and not (layer0_outputs(3385));
    outputs(3339) <= not(layer0_outputs(2150)) or (layer0_outputs(2207));
    outputs(3340) <= (layer0_outputs(4480)) and (layer0_outputs(2537));
    outputs(3341) <= layer0_outputs(2750);
    outputs(3342) <= not(layer0_outputs(3037));
    outputs(3343) <= not(layer0_outputs(1565));
    outputs(3344) <= layer0_outputs(3649);
    outputs(3345) <= (layer0_outputs(1897)) and not (layer0_outputs(2300));
    outputs(3346) <= not(layer0_outputs(50));
    outputs(3347) <= (layer0_outputs(4179)) or (layer0_outputs(4142));
    outputs(3348) <= (layer0_outputs(2147)) and not (layer0_outputs(4067));
    outputs(3349) <= layer0_outputs(1630);
    outputs(3350) <= not(layer0_outputs(3410));
    outputs(3351) <= not((layer0_outputs(1868)) and (layer0_outputs(427)));
    outputs(3352) <= layer0_outputs(2995);
    outputs(3353) <= layer0_outputs(720);
    outputs(3354) <= (layer0_outputs(844)) and not (layer0_outputs(1317));
    outputs(3355) <= not(layer0_outputs(1446));
    outputs(3356) <= not(layer0_outputs(2203));
    outputs(3357) <= layer0_outputs(4444);
    outputs(3358) <= not(layer0_outputs(4846));
    outputs(3359) <= (layer0_outputs(3486)) xor (layer0_outputs(4908));
    outputs(3360) <= (layer0_outputs(161)) and (layer0_outputs(2083));
    outputs(3361) <= not(layer0_outputs(3049));
    outputs(3362) <= (layer0_outputs(1484)) xor (layer0_outputs(4865));
    outputs(3363) <= (layer0_outputs(1574)) and (layer0_outputs(4666));
    outputs(3364) <= layer0_outputs(1079);
    outputs(3365) <= not(layer0_outputs(1623));
    outputs(3366) <= layer0_outputs(3050);
    outputs(3367) <= (layer0_outputs(4774)) xor (layer0_outputs(3754));
    outputs(3368) <= not(layer0_outputs(2414));
    outputs(3369) <= layer0_outputs(2025);
    outputs(3370) <= not((layer0_outputs(2323)) or (layer0_outputs(1001)));
    outputs(3371) <= not(layer0_outputs(780));
    outputs(3372) <= layer0_outputs(2093);
    outputs(3373) <= not(layer0_outputs(2696));
    outputs(3374) <= not(layer0_outputs(4631)) or (layer0_outputs(3074));
    outputs(3375) <= layer0_outputs(4722);
    outputs(3376) <= (layer0_outputs(4537)) or (layer0_outputs(174));
    outputs(3377) <= not((layer0_outputs(426)) or (layer0_outputs(1572)));
    outputs(3378) <= (layer0_outputs(3256)) and not (layer0_outputs(1078));
    outputs(3379) <= (layer0_outputs(3162)) or (layer0_outputs(325));
    outputs(3380) <= layer0_outputs(529);
    outputs(3381) <= layer0_outputs(412);
    outputs(3382) <= not(layer0_outputs(2759));
    outputs(3383) <= not(layer0_outputs(4050));
    outputs(3384) <= not((layer0_outputs(835)) or (layer0_outputs(948)));
    outputs(3385) <= not((layer0_outputs(1525)) or (layer0_outputs(2379)));
    outputs(3386) <= not((layer0_outputs(4094)) or (layer0_outputs(4028)));
    outputs(3387) <= layer0_outputs(4571);
    outputs(3388) <= not((layer0_outputs(1209)) xor (layer0_outputs(3961)));
    outputs(3389) <= not((layer0_outputs(4429)) xor (layer0_outputs(3166)));
    outputs(3390) <= not(layer0_outputs(2783));
    outputs(3391) <= not(layer0_outputs(3686)) or (layer0_outputs(1742));
    outputs(3392) <= layer0_outputs(208);
    outputs(3393) <= (layer0_outputs(2310)) and not (layer0_outputs(585));
    outputs(3394) <= not((layer0_outputs(3478)) or (layer0_outputs(2159)));
    outputs(3395) <= not((layer0_outputs(1280)) or (layer0_outputs(4510)));
    outputs(3396) <= not(layer0_outputs(89));
    outputs(3397) <= not(layer0_outputs(679));
    outputs(3398) <= layer0_outputs(2706);
    outputs(3399) <= not(layer0_outputs(1579));
    outputs(3400) <= not(layer0_outputs(954));
    outputs(3401) <= not(layer0_outputs(2521)) or (layer0_outputs(833));
    outputs(3402) <= not((layer0_outputs(2760)) or (layer0_outputs(4432)));
    outputs(3403) <= not((layer0_outputs(3727)) or (layer0_outputs(3100)));
    outputs(3404) <= not(layer0_outputs(3491)) or (layer0_outputs(97));
    outputs(3405) <= (layer0_outputs(1259)) and not (layer0_outputs(1661));
    outputs(3406) <= not((layer0_outputs(3010)) xor (layer0_outputs(3146)));
    outputs(3407) <= (layer0_outputs(767)) and (layer0_outputs(4814));
    outputs(3408) <= not((layer0_outputs(5021)) xor (layer0_outputs(337)));
    outputs(3409) <= not(layer0_outputs(527));
    outputs(3410) <= layer0_outputs(957);
    outputs(3411) <= not((layer0_outputs(692)) and (layer0_outputs(4531)));
    outputs(3412) <= (layer0_outputs(142)) xor (layer0_outputs(3674));
    outputs(3413) <= not((layer0_outputs(1528)) and (layer0_outputs(4479)));
    outputs(3414) <= not(layer0_outputs(814)) or (layer0_outputs(2402));
    outputs(3415) <= (layer0_outputs(4692)) and not (layer0_outputs(4023));
    outputs(3416) <= (layer0_outputs(220)) xor (layer0_outputs(772));
    outputs(3417) <= not((layer0_outputs(3819)) xor (layer0_outputs(440)));
    outputs(3418) <= not(layer0_outputs(520));
    outputs(3419) <= not(layer0_outputs(3908));
    outputs(3420) <= layer0_outputs(2774);
    outputs(3421) <= layer0_outputs(1003);
    outputs(3422) <= layer0_outputs(493);
    outputs(3423) <= (layer0_outputs(1219)) and not (layer0_outputs(4435));
    outputs(3424) <= not(layer0_outputs(3950));
    outputs(3425) <= (layer0_outputs(1760)) and not (layer0_outputs(5030));
    outputs(3426) <= not(layer0_outputs(882));
    outputs(3427) <= not(layer0_outputs(2864));
    outputs(3428) <= (layer0_outputs(5099)) or (layer0_outputs(1959));
    outputs(3429) <= (layer0_outputs(2641)) and not (layer0_outputs(3367));
    outputs(3430) <= (layer0_outputs(793)) or (layer0_outputs(4004));
    outputs(3431) <= (layer0_outputs(3990)) and not (layer0_outputs(326));
    outputs(3432) <= (layer0_outputs(2974)) and not (layer0_outputs(4298));
    outputs(3433) <= not(layer0_outputs(422));
    outputs(3434) <= (layer0_outputs(1516)) and not (layer0_outputs(1900));
    outputs(3435) <= not(layer0_outputs(2436));
    outputs(3436) <= (layer0_outputs(537)) and (layer0_outputs(1093));
    outputs(3437) <= layer0_outputs(4465);
    outputs(3438) <= not((layer0_outputs(5105)) xor (layer0_outputs(4466)));
    outputs(3439) <= (layer0_outputs(1318)) and not (layer0_outputs(1343));
    outputs(3440) <= (layer0_outputs(4246)) or (layer0_outputs(1302));
    outputs(3441) <= (layer0_outputs(2918)) and not (layer0_outputs(3358));
    outputs(3442) <= not(layer0_outputs(4973));
    outputs(3443) <= not(layer0_outputs(2784));
    outputs(3444) <= not(layer0_outputs(1197)) or (layer0_outputs(3107));
    outputs(3445) <= not(layer0_outputs(931));
    outputs(3446) <= not(layer0_outputs(1661));
    outputs(3447) <= (layer0_outputs(5016)) and (layer0_outputs(3255));
    outputs(3448) <= not(layer0_outputs(4802));
    outputs(3449) <= (layer0_outputs(4120)) xor (layer0_outputs(4968));
    outputs(3450) <= (layer0_outputs(417)) and not (layer0_outputs(2077));
    outputs(3451) <= layer0_outputs(1366);
    outputs(3452) <= (layer0_outputs(4012)) xor (layer0_outputs(1231));
    outputs(3453) <= layer0_outputs(587);
    outputs(3454) <= not((layer0_outputs(2212)) or (layer0_outputs(3024)));
    outputs(3455) <= (layer0_outputs(1739)) and not (layer0_outputs(4869));
    outputs(3456) <= (layer0_outputs(314)) and (layer0_outputs(4974));
    outputs(3457) <= not(layer0_outputs(1153));
    outputs(3458) <= (layer0_outputs(4410)) and not (layer0_outputs(708));
    outputs(3459) <= (layer0_outputs(1506)) and (layer0_outputs(4681));
    outputs(3460) <= (layer0_outputs(4277)) and not (layer0_outputs(528));
    outputs(3461) <= not(layer0_outputs(3442));
    outputs(3462) <= not(layer0_outputs(3176));
    outputs(3463) <= not(layer0_outputs(4450));
    outputs(3464) <= layer0_outputs(988);
    outputs(3465) <= not(layer0_outputs(4574)) or (layer0_outputs(3321));
    outputs(3466) <= layer0_outputs(583);
    outputs(3467) <= layer0_outputs(3228);
    outputs(3468) <= not(layer0_outputs(3258));
    outputs(3469) <= layer0_outputs(4260);
    outputs(3470) <= layer0_outputs(3446);
    outputs(3471) <= not(layer0_outputs(1206));
    outputs(3472) <= (layer0_outputs(2624)) xor (layer0_outputs(1526));
    outputs(3473) <= layer0_outputs(2796);
    outputs(3474) <= (layer0_outputs(818)) xor (layer0_outputs(1012));
    outputs(3475) <= (layer0_outputs(454)) and (layer0_outputs(4114));
    outputs(3476) <= not((layer0_outputs(3504)) or (layer0_outputs(1552)));
    outputs(3477) <= not(layer0_outputs(2123));
    outputs(3478) <= not(layer0_outputs(2173));
    outputs(3479) <= layer0_outputs(4874);
    outputs(3480) <= layer0_outputs(3941);
    outputs(3481) <= not((layer0_outputs(4129)) and (layer0_outputs(2463)));
    outputs(3482) <= not((layer0_outputs(4702)) or (layer0_outputs(4581)));
    outputs(3483) <= not(layer0_outputs(2893));
    outputs(3484) <= not(layer0_outputs(3875));
    outputs(3485) <= not((layer0_outputs(3060)) or (layer0_outputs(2122)));
    outputs(3486) <= (layer0_outputs(1049)) xor (layer0_outputs(463));
    outputs(3487) <= not(layer0_outputs(4882));
    outputs(3488) <= not(layer0_outputs(3346));
    outputs(3489) <= not(layer0_outputs(2789));
    outputs(3490) <= (layer0_outputs(3935)) and not (layer0_outputs(2443));
    outputs(3491) <= (layer0_outputs(2056)) or (layer0_outputs(4032));
    outputs(3492) <= not(layer0_outputs(4458));
    outputs(3493) <= not((layer0_outputs(4426)) or (layer0_outputs(1431)));
    outputs(3494) <= (layer0_outputs(3628)) and not (layer0_outputs(4026));
    outputs(3495) <= (layer0_outputs(3597)) xor (layer0_outputs(579));
    outputs(3496) <= (layer0_outputs(1608)) and not (layer0_outputs(4342));
    outputs(3497) <= (layer0_outputs(2612)) xor (layer0_outputs(256));
    outputs(3498) <= (layer0_outputs(1686)) and not (layer0_outputs(1108));
    outputs(3499) <= not((layer0_outputs(858)) and (layer0_outputs(455)));
    outputs(3500) <= (layer0_outputs(4606)) and (layer0_outputs(1424));
    outputs(3501) <= not((layer0_outputs(3920)) xor (layer0_outputs(1200)));
    outputs(3502) <= not((layer0_outputs(3165)) or (layer0_outputs(2721)));
    outputs(3503) <= layer0_outputs(4651);
    outputs(3504) <= (layer0_outputs(4101)) and (layer0_outputs(1915));
    outputs(3505) <= layer0_outputs(3751);
    outputs(3506) <= layer0_outputs(2006);
    outputs(3507) <= not((layer0_outputs(700)) xor (layer0_outputs(1711)));
    outputs(3508) <= (layer0_outputs(838)) xor (layer0_outputs(3263));
    outputs(3509) <= (layer0_outputs(1236)) xor (layer0_outputs(5051));
    outputs(3510) <= (layer0_outputs(3569)) and not (layer0_outputs(2090));
    outputs(3511) <= not((layer0_outputs(2476)) xor (layer0_outputs(2809)));
    outputs(3512) <= not((layer0_outputs(4595)) xor (layer0_outputs(3230)));
    outputs(3513) <= (layer0_outputs(1740)) and (layer0_outputs(2538));
    outputs(3514) <= layer0_outputs(978);
    outputs(3515) <= not((layer0_outputs(3541)) or (layer0_outputs(1347)));
    outputs(3516) <= layer0_outputs(1284);
    outputs(3517) <= not(layer0_outputs(1455));
    outputs(3518) <= layer0_outputs(650);
    outputs(3519) <= (layer0_outputs(1758)) or (layer0_outputs(3832));
    outputs(3520) <= not(layer0_outputs(342));
    outputs(3521) <= (layer0_outputs(82)) and not (layer0_outputs(3212));
    outputs(3522) <= (layer0_outputs(3154)) and (layer0_outputs(1287));
    outputs(3523) <= not(layer0_outputs(3813));
    outputs(3524) <= not((layer0_outputs(4248)) and (layer0_outputs(3861)));
    outputs(3525) <= not((layer0_outputs(928)) xor (layer0_outputs(4784)));
    outputs(3526) <= layer0_outputs(3192);
    outputs(3527) <= layer0_outputs(4228);
    outputs(3528) <= (layer0_outputs(336)) xor (layer0_outputs(662));
    outputs(3529) <= not((layer0_outputs(1773)) or (layer0_outputs(5052)));
    outputs(3530) <= layer0_outputs(1273);
    outputs(3531) <= not(layer0_outputs(779));
    outputs(3532) <= not(layer0_outputs(3174));
    outputs(3533) <= not(layer0_outputs(2341));
    outputs(3534) <= not(layer0_outputs(1655));
    outputs(3535) <= layer0_outputs(2727);
    outputs(3536) <= not((layer0_outputs(3978)) or (layer0_outputs(366)));
    outputs(3537) <= layer0_outputs(1319);
    outputs(3538) <= not(layer0_outputs(2881));
    outputs(3539) <= (layer0_outputs(2407)) and (layer0_outputs(1875));
    outputs(3540) <= not(layer0_outputs(3865));
    outputs(3541) <= (layer0_outputs(4519)) or (layer0_outputs(4949));
    outputs(3542) <= layer0_outputs(2649);
    outputs(3543) <= not((layer0_outputs(562)) or (layer0_outputs(2619)));
    outputs(3544) <= not(layer0_outputs(345));
    outputs(3545) <= not(layer0_outputs(2745));
    outputs(3546) <= not(layer0_outputs(4706));
    outputs(3547) <= not(layer0_outputs(3891)) or (layer0_outputs(5076));
    outputs(3548) <= not(layer0_outputs(1752));
    outputs(3549) <= not(layer0_outputs(2282));
    outputs(3550) <= layer0_outputs(4294);
    outputs(3551) <= layer0_outputs(4892);
    outputs(3552) <= (layer0_outputs(4086)) and (layer0_outputs(709));
    outputs(3553) <= (layer0_outputs(3267)) or (layer0_outputs(3236));
    outputs(3554) <= (layer0_outputs(180)) and (layer0_outputs(1544));
    outputs(3555) <= (layer0_outputs(909)) or (layer0_outputs(4783));
    outputs(3556) <= not((layer0_outputs(1490)) xor (layer0_outputs(740)));
    outputs(3557) <= (layer0_outputs(933)) and (layer0_outputs(3464));
    outputs(3558) <= not(layer0_outputs(328));
    outputs(3559) <= not(layer0_outputs(4172));
    outputs(3560) <= (layer0_outputs(3905)) and (layer0_outputs(4843));
    outputs(3561) <= not(layer0_outputs(4292));
    outputs(3562) <= (layer0_outputs(2717)) and (layer0_outputs(4864));
    outputs(3563) <= not((layer0_outputs(1562)) and (layer0_outputs(4830)));
    outputs(3564) <= not(layer0_outputs(3189));
    outputs(3565) <= not(layer0_outputs(370));
    outputs(3566) <= (layer0_outputs(54)) and not (layer0_outputs(3709));
    outputs(3567) <= (layer0_outputs(4920)) or (layer0_outputs(1591));
    outputs(3568) <= (layer0_outputs(3862)) and not (layer0_outputs(4526));
    outputs(3569) <= not((layer0_outputs(4169)) xor (layer0_outputs(2134)));
    outputs(3570) <= (layer0_outputs(1491)) xor (layer0_outputs(3913));
    outputs(3571) <= (layer0_outputs(3662)) and not (layer0_outputs(1802));
    outputs(3572) <= (layer0_outputs(1778)) and not (layer0_outputs(26));
    outputs(3573) <= layer0_outputs(4698);
    outputs(3574) <= not(layer0_outputs(2517));
    outputs(3575) <= (layer0_outputs(4683)) and (layer0_outputs(2663));
    outputs(3576) <= layer0_outputs(982);
    outputs(3577) <= (layer0_outputs(1890)) or (layer0_outputs(5033));
    outputs(3578) <= not(layer0_outputs(3305));
    outputs(3579) <= layer0_outputs(2367);
    outputs(3580) <= (layer0_outputs(801)) and not (layer0_outputs(1388));
    outputs(3581) <= layer0_outputs(2319);
    outputs(3582) <= (layer0_outputs(2085)) and not (layer0_outputs(1517));
    outputs(3583) <= layer0_outputs(2194);
    outputs(3584) <= (layer0_outputs(277)) and (layer0_outputs(2255));
    outputs(3585) <= not(layer0_outputs(1288));
    outputs(3586) <= (layer0_outputs(1709)) and not (layer0_outputs(21));
    outputs(3587) <= not((layer0_outputs(4131)) or (layer0_outputs(4256)));
    outputs(3588) <= (layer0_outputs(3523)) and not (layer0_outputs(4943));
    outputs(3589) <= (layer0_outputs(4172)) and not (layer0_outputs(462));
    outputs(3590) <= layer0_outputs(912);
    outputs(3591) <= not(layer0_outputs(2322));
    outputs(3592) <= (layer0_outputs(3875)) and not (layer0_outputs(751));
    outputs(3593) <= (layer0_outputs(1350)) and not (layer0_outputs(2305));
    outputs(3594) <= (layer0_outputs(3442)) and not (layer0_outputs(3181));
    outputs(3595) <= layer0_outputs(2273);
    outputs(3596) <= (layer0_outputs(466)) and not (layer0_outputs(5045));
    outputs(3597) <= (layer0_outputs(2474)) and (layer0_outputs(2604));
    outputs(3598) <= layer0_outputs(1362);
    outputs(3599) <= not(layer0_outputs(4014));
    outputs(3600) <= (layer0_outputs(4957)) and (layer0_outputs(58));
    outputs(3601) <= (layer0_outputs(403)) and not (layer0_outputs(1385));
    outputs(3602) <= layer0_outputs(2320);
    outputs(3603) <= layer0_outputs(651);
    outputs(3604) <= not((layer0_outputs(1744)) or (layer0_outputs(3762)));
    outputs(3605) <= (layer0_outputs(259)) and (layer0_outputs(4734));
    outputs(3606) <= not(layer0_outputs(3218));
    outputs(3607) <= (layer0_outputs(1494)) and (layer0_outputs(3424));
    outputs(3608) <= layer0_outputs(1907);
    outputs(3609) <= layer0_outputs(3951);
    outputs(3610) <= not(layer0_outputs(4121));
    outputs(3611) <= not(layer0_outputs(2989));
    outputs(3612) <= (layer0_outputs(469)) and (layer0_outputs(701));
    outputs(3613) <= (layer0_outputs(1652)) and not (layer0_outputs(3374));
    outputs(3614) <= not(layer0_outputs(2072));
    outputs(3615) <= not(layer0_outputs(1998));
    outputs(3616) <= (layer0_outputs(3778)) and (layer0_outputs(578));
    outputs(3617) <= layer0_outputs(2442);
    outputs(3618) <= not(layer0_outputs(4406));
    outputs(3619) <= not((layer0_outputs(2440)) and (layer0_outputs(3276)));
    outputs(3620) <= (layer0_outputs(3847)) and not (layer0_outputs(1330));
    outputs(3621) <= layer0_outputs(5107);
    outputs(3622) <= (layer0_outputs(902)) xor (layer0_outputs(3115));
    outputs(3623) <= layer0_outputs(1824);
    outputs(3624) <= (layer0_outputs(1199)) and not (layer0_outputs(4804));
    outputs(3625) <= not(layer0_outputs(1075));
    outputs(3626) <= layer0_outputs(5106);
    outputs(3627) <= (layer0_outputs(2905)) and not (layer0_outputs(4966));
    outputs(3628) <= not((layer0_outputs(2142)) xor (layer0_outputs(1186)));
    outputs(3629) <= (layer0_outputs(4546)) xor (layer0_outputs(1578));
    outputs(3630) <= (layer0_outputs(1617)) and (layer0_outputs(1937));
    outputs(3631) <= not(layer0_outputs(3381));
    outputs(3632) <= not(layer0_outputs(1097));
    outputs(3633) <= (layer0_outputs(3432)) and not (layer0_outputs(2821));
    outputs(3634) <= layer0_outputs(4761);
    outputs(3635) <= layer0_outputs(4249);
    outputs(3636) <= not(layer0_outputs(2804));
    outputs(3637) <= (layer0_outputs(1655)) and not (layer0_outputs(4085));
    outputs(3638) <= layer0_outputs(170);
    outputs(3639) <= (layer0_outputs(764)) and not (layer0_outputs(3947));
    outputs(3640) <= layer0_outputs(5028);
    outputs(3641) <= (layer0_outputs(4863)) and (layer0_outputs(251));
    outputs(3642) <= (layer0_outputs(1893)) and (layer0_outputs(3675));
    outputs(3643) <= (layer0_outputs(275)) and (layer0_outputs(3897));
    outputs(3644) <= (layer0_outputs(2850)) and not (layer0_outputs(3197));
    outputs(3645) <= (layer0_outputs(1682)) and (layer0_outputs(2983));
    outputs(3646) <= not(layer0_outputs(3385));
    outputs(3647) <= not(layer0_outputs(2725));
    outputs(3648) <= layer0_outputs(3629);
    outputs(3649) <= not((layer0_outputs(4647)) or (layer0_outputs(2157)));
    outputs(3650) <= not((layer0_outputs(1871)) or (layer0_outputs(3198)));
    outputs(3651) <= not(layer0_outputs(612));
    outputs(3652) <= not((layer0_outputs(3098)) and (layer0_outputs(1038)));
    outputs(3653) <= (layer0_outputs(2189)) and (layer0_outputs(3165));
    outputs(3654) <= not(layer0_outputs(4616));
    outputs(3655) <= layer0_outputs(4408);
    outputs(3656) <= (layer0_outputs(4736)) and not (layer0_outputs(865));
    outputs(3657) <= (layer0_outputs(886)) and not (layer0_outputs(530));
    outputs(3658) <= (layer0_outputs(3995)) and not (layer0_outputs(3436));
    outputs(3659) <= not((layer0_outputs(4199)) or (layer0_outputs(5003)));
    outputs(3660) <= (layer0_outputs(4310)) and not (layer0_outputs(811));
    outputs(3661) <= layer0_outputs(1072);
    outputs(3662) <= (layer0_outputs(3842)) and not (layer0_outputs(2713));
    outputs(3663) <= not(layer0_outputs(3348)) or (layer0_outputs(3997));
    outputs(3664) <= not(layer0_outputs(5108));
    outputs(3665) <= (layer0_outputs(2532)) and (layer0_outputs(1464));
    outputs(3666) <= not((layer0_outputs(1743)) xor (layer0_outputs(2099)));
    outputs(3667) <= not(layer0_outputs(4257));
    outputs(3668) <= layer0_outputs(4654);
    outputs(3669) <= layer0_outputs(4432);
    outputs(3670) <= (layer0_outputs(2412)) and not (layer0_outputs(2039));
    outputs(3671) <= not(layer0_outputs(4947));
    outputs(3672) <= not((layer0_outputs(599)) or (layer0_outputs(1699)));
    outputs(3673) <= layer0_outputs(1022);
    outputs(3674) <= (layer0_outputs(130)) and not (layer0_outputs(2247));
    outputs(3675) <= not(layer0_outputs(3500));
    outputs(3676) <= not((layer0_outputs(1845)) or (layer0_outputs(2614)));
    outputs(3677) <= layer0_outputs(2838);
    outputs(3678) <= (layer0_outputs(4238)) xor (layer0_outputs(4181));
    outputs(3679) <= (layer0_outputs(2331)) or (layer0_outputs(1698));
    outputs(3680) <= layer0_outputs(4828);
    outputs(3681) <= (layer0_outputs(2811)) and (layer0_outputs(2467));
    outputs(3682) <= layer0_outputs(1941);
    outputs(3683) <= layer0_outputs(2298);
    outputs(3684) <= (layer0_outputs(564)) and (layer0_outputs(2144));
    outputs(3685) <= layer0_outputs(2341);
    outputs(3686) <= not(layer0_outputs(2103));
    outputs(3687) <= not(layer0_outputs(193));
    outputs(3688) <= layer0_outputs(1995);
    outputs(3689) <= not((layer0_outputs(4935)) or (layer0_outputs(544)));
    outputs(3690) <= not((layer0_outputs(542)) or (layer0_outputs(3516)));
    outputs(3691) <= (layer0_outputs(1788)) and (layer0_outputs(3871));
    outputs(3692) <= (layer0_outputs(3288)) and not (layer0_outputs(4491));
    outputs(3693) <= not(layer0_outputs(4685));
    outputs(3694) <= layer0_outputs(1279);
    outputs(3695) <= not(layer0_outputs(3929));
    outputs(3696) <= (layer0_outputs(3078)) and not (layer0_outputs(4225));
    outputs(3697) <= not(layer0_outputs(1512));
    outputs(3698) <= not(layer0_outputs(1242)) or (layer0_outputs(2013));
    outputs(3699) <= not((layer0_outputs(3345)) or (layer0_outputs(4693)));
    outputs(3700) <= not((layer0_outputs(1296)) or (layer0_outputs(781)));
    outputs(3701) <= not((layer0_outputs(3927)) or (layer0_outputs(4221)));
    outputs(3702) <= not((layer0_outputs(4621)) and (layer0_outputs(1874)));
    outputs(3703) <= not((layer0_outputs(2343)) or (layer0_outputs(3822)));
    outputs(3704) <= not((layer0_outputs(2636)) or (layer0_outputs(1724)));
    outputs(3705) <= (layer0_outputs(1800)) and not (layer0_outputs(3745));
    outputs(3706) <= not(layer0_outputs(3480));
    outputs(3707) <= not(layer0_outputs(2608));
    outputs(3708) <= (layer0_outputs(2585)) and not (layer0_outputs(396));
    outputs(3709) <= not(layer0_outputs(483)) or (layer0_outputs(3351));
    outputs(3710) <= (layer0_outputs(3536)) and not (layer0_outputs(655));
    outputs(3711) <= layer0_outputs(4389);
    outputs(3712) <= not(layer0_outputs(1555));
    outputs(3713) <= not(layer0_outputs(1816));
    outputs(3714) <= layer0_outputs(59);
    outputs(3715) <= (layer0_outputs(4059)) and (layer0_outputs(3386));
    outputs(3716) <= not(layer0_outputs(3472));
    outputs(3717) <= not((layer0_outputs(3352)) or (layer0_outputs(1595)));
    outputs(3718) <= not(layer0_outputs(3591));
    outputs(3719) <= (layer0_outputs(2984)) and not (layer0_outputs(368));
    outputs(3720) <= (layer0_outputs(2800)) and not (layer0_outputs(1386));
    outputs(3721) <= (layer0_outputs(2830)) and not (layer0_outputs(1429));
    outputs(3722) <= layer0_outputs(918);
    outputs(3723) <= (layer0_outputs(114)) and not (layer0_outputs(2768));
    outputs(3724) <= layer0_outputs(1088);
    outputs(3725) <= (layer0_outputs(3940)) and not (layer0_outputs(164));
    outputs(3726) <= layer0_outputs(1098);
    outputs(3727) <= not(layer0_outputs(1871));
    outputs(3728) <= not(layer0_outputs(4815)) or (layer0_outputs(4234));
    outputs(3729) <= not((layer0_outputs(4644)) or (layer0_outputs(3893)));
    outputs(3730) <= (layer0_outputs(2064)) and not (layer0_outputs(524));
    outputs(3731) <= not(layer0_outputs(1600));
    outputs(3732) <= not(layer0_outputs(4289));
    outputs(3733) <= (layer0_outputs(3633)) and not (layer0_outputs(2826));
    outputs(3734) <= (layer0_outputs(4830)) and (layer0_outputs(253));
    outputs(3735) <= not(layer0_outputs(3056));
    outputs(3736) <= not(layer0_outputs(3624));
    outputs(3737) <= (layer0_outputs(2382)) and not (layer0_outputs(3604));
    outputs(3738) <= layer0_outputs(1027);
    outputs(3739) <= (layer0_outputs(1784)) xor (layer0_outputs(3914));
    outputs(3740) <= (layer0_outputs(636)) and not (layer0_outputs(3693));
    outputs(3741) <= not(layer0_outputs(169));
    outputs(3742) <= not(layer0_outputs(1923)) or (layer0_outputs(2849));
    outputs(3743) <= (layer0_outputs(1907)) and not (layer0_outputs(2869));
    outputs(3744) <= not((layer0_outputs(3318)) or (layer0_outputs(645)));
    outputs(3745) <= not(layer0_outputs(988));
    outputs(3746) <= (layer0_outputs(2891)) xor (layer0_outputs(265));
    outputs(3747) <= not(layer0_outputs(3420));
    outputs(3748) <= not(layer0_outputs(2733));
    outputs(3749) <= layer0_outputs(1581);
    outputs(3750) <= layer0_outputs(1072);
    outputs(3751) <= layer0_outputs(647);
    outputs(3752) <= (layer0_outputs(2556)) and not (layer0_outputs(3200));
    outputs(3753) <= not((layer0_outputs(2990)) xor (layer0_outputs(3951)));
    outputs(3754) <= (layer0_outputs(2501)) and (layer0_outputs(4309));
    outputs(3755) <= not((layer0_outputs(689)) and (layer0_outputs(291)));
    outputs(3756) <= not(layer0_outputs(4349));
    outputs(3757) <= not((layer0_outputs(1521)) or (layer0_outputs(3452)));
    outputs(3758) <= not(layer0_outputs(1905)) or (layer0_outputs(3168));
    outputs(3759) <= not(layer0_outputs(3407));
    outputs(3760) <= not(layer0_outputs(4093));
    outputs(3761) <= not(layer0_outputs(967));
    outputs(3762) <= not(layer0_outputs(1417));
    outputs(3763) <= (layer0_outputs(1164)) and not (layer0_outputs(2366));
    outputs(3764) <= not((layer0_outputs(5053)) xor (layer0_outputs(39)));
    outputs(3765) <= not((layer0_outputs(4250)) or (layer0_outputs(2381)));
    outputs(3766) <= not(layer0_outputs(2080));
    outputs(3767) <= not(layer0_outputs(4281));
    outputs(3768) <= not(layer0_outputs(2573));
    outputs(3769) <= not(layer0_outputs(2464)) or (layer0_outputs(3618));
    outputs(3770) <= (layer0_outputs(2721)) and (layer0_outputs(555));
    outputs(3771) <= not(layer0_outputs(4373));
    outputs(3772) <= not(layer0_outputs(5067));
    outputs(3773) <= layer0_outputs(1208);
    outputs(3774) <= not(layer0_outputs(4250));
    outputs(3775) <= (layer0_outputs(3338)) and not (layer0_outputs(1395));
    outputs(3776) <= (layer0_outputs(3404)) and (layer0_outputs(808));
    outputs(3777) <= not((layer0_outputs(392)) or (layer0_outputs(990)));
    outputs(3778) <= layer0_outputs(1473);
    outputs(3779) <= not(layer0_outputs(2709)) or (layer0_outputs(2129));
    outputs(3780) <= not(layer0_outputs(3749));
    outputs(3781) <= layer0_outputs(1789);
    outputs(3782) <= (layer0_outputs(931)) and not (layer0_outputs(3007));
    outputs(3783) <= layer0_outputs(1729);
    outputs(3784) <= not(layer0_outputs(2703));
    outputs(3785) <= not((layer0_outputs(1983)) xor (layer0_outputs(3061)));
    outputs(3786) <= (layer0_outputs(1619)) and not (layer0_outputs(1017));
    outputs(3787) <= not((layer0_outputs(380)) xor (layer0_outputs(4113)));
    outputs(3788) <= (layer0_outputs(481)) xor (layer0_outputs(1113));
    outputs(3789) <= not(layer0_outputs(1038)) or (layer0_outputs(278));
    outputs(3790) <= layer0_outputs(488);
    outputs(3791) <= (layer0_outputs(1963)) and not (layer0_outputs(4318));
    outputs(3792) <= (layer0_outputs(768)) and not (layer0_outputs(2495));
    outputs(3793) <= layer0_outputs(4137);
    outputs(3794) <= layer0_outputs(3689);
    outputs(3795) <= (layer0_outputs(2015)) xor (layer0_outputs(3206));
    outputs(3796) <= layer0_outputs(4729);
    outputs(3797) <= not((layer0_outputs(3758)) or (layer0_outputs(4556)));
    outputs(3798) <= not((layer0_outputs(3467)) or (layer0_outputs(4541)));
    outputs(3799) <= not((layer0_outputs(3052)) xor (layer0_outputs(2518)));
    outputs(3800) <= (layer0_outputs(2925)) and (layer0_outputs(2881));
    outputs(3801) <= not((layer0_outputs(2030)) and (layer0_outputs(3581)));
    outputs(3802) <= not((layer0_outputs(1495)) or (layer0_outputs(60)));
    outputs(3803) <= (layer0_outputs(2494)) or (layer0_outputs(3033));
    outputs(3804) <= (layer0_outputs(2976)) and (layer0_outputs(429));
    outputs(3805) <= (layer0_outputs(1645)) and not (layer0_outputs(4420));
    outputs(3806) <= (layer0_outputs(2481)) or (layer0_outputs(331));
    outputs(3807) <= not((layer0_outputs(393)) or (layer0_outputs(375)));
    outputs(3808) <= (layer0_outputs(1961)) and not (layer0_outputs(2735));
    outputs(3809) <= not(layer0_outputs(3954));
    outputs(3810) <= (layer0_outputs(1048)) and not (layer0_outputs(4372));
    outputs(3811) <= not(layer0_outputs(3218));
    outputs(3812) <= layer0_outputs(3530);
    outputs(3813) <= layer0_outputs(4484);
    outputs(3814) <= (layer0_outputs(4430)) and (layer0_outputs(5059));
    outputs(3815) <= layer0_outputs(2485);
    outputs(3816) <= not(layer0_outputs(3558));
    outputs(3817) <= not(layer0_outputs(4271));
    outputs(3818) <= not(layer0_outputs(2616));
    outputs(3819) <= not((layer0_outputs(294)) or (layer0_outputs(3139)));
    outputs(3820) <= (layer0_outputs(1683)) and (layer0_outputs(3295));
    outputs(3821) <= not((layer0_outputs(4274)) or (layer0_outputs(2267)));
    outputs(3822) <= not((layer0_outputs(1296)) or (layer0_outputs(1405)));
    outputs(3823) <= (layer0_outputs(2888)) xor (layer0_outputs(5031));
    outputs(3824) <= not(layer0_outputs(713));
    outputs(3825) <= (layer0_outputs(643)) and not (layer0_outputs(2429));
    outputs(3826) <= layer0_outputs(198);
    outputs(3827) <= layer0_outputs(1342);
    outputs(3828) <= (layer0_outputs(4320)) and not (layer0_outputs(1187));
    outputs(3829) <= (layer0_outputs(930)) and not (layer0_outputs(1400));
    outputs(3830) <= layer0_outputs(468);
    outputs(3831) <= not((layer0_outputs(4952)) or (layer0_outputs(2642)));
    outputs(3832) <= not((layer0_outputs(2417)) or (layer0_outputs(3792)));
    outputs(3833) <= not((layer0_outputs(2742)) or (layer0_outputs(24)));
    outputs(3834) <= layer0_outputs(2653);
    outputs(3835) <= layer0_outputs(3552);
    outputs(3836) <= not(layer0_outputs(3333));
    outputs(3837) <= (layer0_outputs(3394)) xor (layer0_outputs(4360));
    outputs(3838) <= not((layer0_outputs(3240)) or (layer0_outputs(206)));
    outputs(3839) <= not(layer0_outputs(2840));
    outputs(3840) <= (layer0_outputs(3606)) xor (layer0_outputs(120));
    outputs(3841) <= layer0_outputs(2653);
    outputs(3842) <= (layer0_outputs(1692)) or (layer0_outputs(4950));
    outputs(3843) <= not(layer0_outputs(301)) or (layer0_outputs(1089));
    outputs(3844) <= (layer0_outputs(1606)) and (layer0_outputs(590));
    outputs(3845) <= not(layer0_outputs(3787));
    outputs(3846) <= (layer0_outputs(4490)) and (layer0_outputs(1298));
    outputs(3847) <= (layer0_outputs(1124)) and (layer0_outputs(954));
    outputs(3848) <= not(layer0_outputs(4916));
    outputs(3849) <= (layer0_outputs(2958)) and not (layer0_outputs(3631));
    outputs(3850) <= (layer0_outputs(280)) and (layer0_outputs(401));
    outputs(3851) <= (layer0_outputs(4043)) and not (layer0_outputs(2885));
    outputs(3852) <= not((layer0_outputs(2388)) or (layer0_outputs(4350)));
    outputs(3853) <= layer0_outputs(632);
    outputs(3854) <= (layer0_outputs(867)) or (layer0_outputs(1938));
    outputs(3855) <= not((layer0_outputs(558)) or (layer0_outputs(1935)));
    outputs(3856) <= layer0_outputs(1977);
    outputs(3857) <= not((layer0_outputs(2399)) xor (layer0_outputs(3789)));
    outputs(3858) <= (layer0_outputs(3085)) xor (layer0_outputs(2962));
    outputs(3859) <= not((layer0_outputs(1615)) and (layer0_outputs(4339)));
    outputs(3860) <= not(layer0_outputs(4630));
    outputs(3861) <= layer0_outputs(2017);
    outputs(3862) <= not(layer0_outputs(2650));
    outputs(3863) <= (layer0_outputs(4385)) and (layer0_outputs(2827));
    outputs(3864) <= (layer0_outputs(1451)) xor (layer0_outputs(2094));
    outputs(3865) <= not((layer0_outputs(1541)) or (layer0_outputs(874)));
    outputs(3866) <= layer0_outputs(4723);
    outputs(3867) <= not(layer0_outputs(830));
    outputs(3868) <= (layer0_outputs(2933)) and (layer0_outputs(899));
    outputs(3869) <= not(layer0_outputs(2547));
    outputs(3870) <= layer0_outputs(2533);
    outputs(3871) <= (layer0_outputs(1)) and (layer0_outputs(4611));
    outputs(3872) <= (layer0_outputs(100)) xor (layer0_outputs(3148));
    outputs(3873) <= (layer0_outputs(2246)) xor (layer0_outputs(3027));
    outputs(3874) <= layer0_outputs(3859);
    outputs(3875) <= (layer0_outputs(5082)) and not (layer0_outputs(3083));
    outputs(3876) <= not((layer0_outputs(4387)) xor (layer0_outputs(3445)));
    outputs(3877) <= not((layer0_outputs(4037)) xor (layer0_outputs(2271)));
    outputs(3878) <= (layer0_outputs(3020)) and (layer0_outputs(4213));
    outputs(3879) <= not((layer0_outputs(1590)) or (layer0_outputs(482)));
    outputs(3880) <= (layer0_outputs(4460)) and not (layer0_outputs(3569));
    outputs(3881) <= (layer0_outputs(832)) and not (layer0_outputs(2788));
    outputs(3882) <= (layer0_outputs(3999)) and not (layer0_outputs(3493));
    outputs(3883) <= (layer0_outputs(444)) and not (layer0_outputs(1540));
    outputs(3884) <= (layer0_outputs(4656)) xor (layer0_outputs(4833));
    outputs(3885) <= layer0_outputs(2602);
    outputs(3886) <= layer0_outputs(4017);
    outputs(3887) <= not(layer0_outputs(1763));
    outputs(3888) <= not((layer0_outputs(4362)) or (layer0_outputs(283)));
    outputs(3889) <= (layer0_outputs(3488)) and (layer0_outputs(3637));
    outputs(3890) <= (layer0_outputs(5042)) and not (layer0_outputs(3476));
    outputs(3891) <= not((layer0_outputs(3936)) or (layer0_outputs(1699)));
    outputs(3892) <= not(layer0_outputs(77));
    outputs(3893) <= not(layer0_outputs(2818)) or (layer0_outputs(1430));
    outputs(3894) <= (layer0_outputs(3062)) and (layer0_outputs(1815));
    outputs(3895) <= (layer0_outputs(1205)) and (layer0_outputs(2016));
    outputs(3896) <= layer0_outputs(2273);
    outputs(3897) <= not((layer0_outputs(1688)) or (layer0_outputs(3224)));
    outputs(3898) <= (layer0_outputs(1889)) and not (layer0_outputs(5046));
    outputs(3899) <= (layer0_outputs(1099)) xor (layer0_outputs(2307));
    outputs(3900) <= (layer0_outputs(3176)) and (layer0_outputs(844));
    outputs(3901) <= not(layer0_outputs(238));
    outputs(3902) <= (layer0_outputs(4896)) and (layer0_outputs(996));
    outputs(3903) <= not((layer0_outputs(4404)) or (layer0_outputs(1820)));
    outputs(3904) <= not(layer0_outputs(2114));
    outputs(3905) <= (layer0_outputs(2569)) and not (layer0_outputs(2386));
    outputs(3906) <= not((layer0_outputs(2302)) or (layer0_outputs(758)));
    outputs(3907) <= not(layer0_outputs(2857));
    outputs(3908) <= (layer0_outputs(3864)) and not (layer0_outputs(4783));
    outputs(3909) <= not(layer0_outputs(3499));
    outputs(3910) <= (layer0_outputs(3099)) and not (layer0_outputs(4224));
    outputs(3911) <= not(layer0_outputs(446));
    outputs(3912) <= (layer0_outputs(1274)) or (layer0_outputs(2617));
    outputs(3913) <= (layer0_outputs(4500)) and not (layer0_outputs(4040));
    outputs(3914) <= (layer0_outputs(4184)) and not (layer0_outputs(3433));
    outputs(3915) <= not(layer0_outputs(1386));
    outputs(3916) <= (layer0_outputs(5072)) and not (layer0_outputs(1021));
    outputs(3917) <= layer0_outputs(3402);
    outputs(3918) <= layer0_outputs(1825);
    outputs(3919) <= layer0_outputs(4593);
    outputs(3920) <= not((layer0_outputs(3000)) or (layer0_outputs(4491)));
    outputs(3921) <= layer0_outputs(1174);
    outputs(3922) <= (layer0_outputs(5051)) and not (layer0_outputs(1901));
    outputs(3923) <= not(layer0_outputs(2009));
    outputs(3924) <= (layer0_outputs(4664)) and not (layer0_outputs(1080));
    outputs(3925) <= not((layer0_outputs(1913)) xor (layer0_outputs(606)));
    outputs(3926) <= layer0_outputs(3213);
    outputs(3927) <= (layer0_outputs(4598)) and (layer0_outputs(4464));
    outputs(3928) <= layer0_outputs(4213);
    outputs(3929) <= (layer0_outputs(2812)) and not (layer0_outputs(4325));
    outputs(3930) <= not((layer0_outputs(1016)) or (layer0_outputs(2771)));
    outputs(3931) <= not(layer0_outputs(4438));
    outputs(3932) <= not((layer0_outputs(4442)) xor (layer0_outputs(1371)));
    outputs(3933) <= layer0_outputs(4876);
    outputs(3934) <= layer0_outputs(2767);
    outputs(3935) <= not(layer0_outputs(1586));
    outputs(3936) <= not(layer0_outputs(3204));
    outputs(3937) <= not(layer0_outputs(1468));
    outputs(3938) <= layer0_outputs(4904);
    outputs(3939) <= not(layer0_outputs(1852));
    outputs(3940) <= layer0_outputs(997);
    outputs(3941) <= not(layer0_outputs(1080));
    outputs(3942) <= not(layer0_outputs(3345));
    outputs(3943) <= layer0_outputs(706);
    outputs(3944) <= not((layer0_outputs(5080)) and (layer0_outputs(3529)));
    outputs(3945) <= (layer0_outputs(4548)) and not (layer0_outputs(800));
    outputs(3946) <= not((layer0_outputs(2550)) or (layer0_outputs(4591)));
    outputs(3947) <= not(layer0_outputs(5018));
    outputs(3948) <= layer0_outputs(278);
    outputs(3949) <= (layer0_outputs(1161)) and not (layer0_outputs(967));
    outputs(3950) <= not(layer0_outputs(2705));
    outputs(3951) <= not(layer0_outputs(521));
    outputs(3952) <= not(layer0_outputs(1880));
    outputs(3953) <= (layer0_outputs(480)) and (layer0_outputs(4494));
    outputs(3954) <= not(layer0_outputs(2058));
    outputs(3955) <= (layer0_outputs(4764)) and not (layer0_outputs(5068));
    outputs(3956) <= layer0_outputs(398);
    outputs(3957) <= layer0_outputs(1009);
    outputs(3958) <= layer0_outputs(4392);
    outputs(3959) <= not(layer0_outputs(5084));
    outputs(3960) <= not((layer0_outputs(219)) or (layer0_outputs(2975)));
    outputs(3961) <= not((layer0_outputs(4955)) or (layer0_outputs(1055)));
    outputs(3962) <= layer0_outputs(256);
    outputs(3963) <= (layer0_outputs(2059)) and (layer0_outputs(2101));
    outputs(3964) <= (layer0_outputs(3548)) and not (layer0_outputs(2747));
    outputs(3965) <= (layer0_outputs(4163)) and not (layer0_outputs(1117));
    outputs(3966) <= (layer0_outputs(1204)) and not (layer0_outputs(2610));
    outputs(3967) <= (layer0_outputs(4969)) or (layer0_outputs(1483));
    outputs(3968) <= not(layer0_outputs(3456));
    outputs(3969) <= (layer0_outputs(1563)) and not (layer0_outputs(162));
    outputs(3970) <= not(layer0_outputs(542));
    outputs(3971) <= (layer0_outputs(4530)) and not (layer0_outputs(3837));
    outputs(3972) <= (layer0_outputs(3154)) and (layer0_outputs(2086));
    outputs(3973) <= not(layer0_outputs(659));
    outputs(3974) <= (layer0_outputs(608)) and not (layer0_outputs(1958));
    outputs(3975) <= (layer0_outputs(191)) and not (layer0_outputs(4826));
    outputs(3976) <= (layer0_outputs(1065)) and not (layer0_outputs(1347));
    outputs(3977) <= not((layer0_outputs(2878)) or (layer0_outputs(1588)));
    outputs(3978) <= (layer0_outputs(1867)) xor (layer0_outputs(2751));
    outputs(3979) <= (layer0_outputs(3788)) and not (layer0_outputs(5070));
    outputs(3980) <= layer0_outputs(4437);
    outputs(3981) <= (layer0_outputs(991)) and (layer0_outputs(2185));
    outputs(3982) <= (layer0_outputs(2328)) and not (layer0_outputs(2157));
    outputs(3983) <= not(layer0_outputs(4278));
    outputs(3984) <= (layer0_outputs(254)) xor (layer0_outputs(2898));
    outputs(3985) <= (layer0_outputs(3378)) xor (layer0_outputs(641));
    outputs(3986) <= layer0_outputs(2757);
    outputs(3987) <= not((layer0_outputs(1495)) xor (layer0_outputs(1071)));
    outputs(3988) <= (layer0_outputs(1850)) or (layer0_outputs(4321));
    outputs(3989) <= (layer0_outputs(973)) and not (layer0_outputs(268));
    outputs(3990) <= layer0_outputs(3717);
    outputs(3991) <= (layer0_outputs(629)) and not (layer0_outputs(4493));
    outputs(3992) <= not(layer0_outputs(486));
    outputs(3993) <= layer0_outputs(4994);
    outputs(3994) <= not(layer0_outputs(5104));
    outputs(3995) <= (layer0_outputs(3793)) and (layer0_outputs(1238));
    outputs(3996) <= layer0_outputs(2864);
    outputs(3997) <= layer0_outputs(4378);
    outputs(3998) <= not((layer0_outputs(1707)) or (layer0_outputs(3084)));
    outputs(3999) <= not(layer0_outputs(4347));
    outputs(4000) <= not((layer0_outputs(3407)) or (layer0_outputs(2575)));
    outputs(4001) <= not(layer0_outputs(1844));
    outputs(4002) <= not(layer0_outputs(3038));
    outputs(4003) <= (layer0_outputs(4771)) and not (layer0_outputs(1985));
    outputs(4004) <= (layer0_outputs(1752)) and not (layer0_outputs(4152));
    outputs(4005) <= not(layer0_outputs(452));
    outputs(4006) <= (layer0_outputs(1936)) and (layer0_outputs(808));
    outputs(4007) <= (layer0_outputs(4753)) or (layer0_outputs(3515));
    outputs(4008) <= (layer0_outputs(554)) and not (layer0_outputs(1420));
    outputs(4009) <= (layer0_outputs(3907)) xor (layer0_outputs(927));
    outputs(4010) <= layer0_outputs(3986);
    outputs(4011) <= layer0_outputs(5075);
    outputs(4012) <= layer0_outputs(427);
    outputs(4013) <= not((layer0_outputs(2718)) xor (layer0_outputs(4128)));
    outputs(4014) <= (layer0_outputs(1441)) and not (layer0_outputs(413));
    outputs(4015) <= layer0_outputs(1182);
    outputs(4016) <= (layer0_outputs(1448)) and not (layer0_outputs(83));
    outputs(4017) <= not((layer0_outputs(3209)) and (layer0_outputs(39)));
    outputs(4018) <= (layer0_outputs(3018)) and not (layer0_outputs(1836));
    outputs(4019) <= layer0_outputs(5047);
    outputs(4020) <= (layer0_outputs(3520)) and (layer0_outputs(2487));
    outputs(4021) <= (layer0_outputs(4503)) and not (layer0_outputs(2261));
    outputs(4022) <= not(layer0_outputs(4116));
    outputs(4023) <= (layer0_outputs(459)) and not (layer0_outputs(3369));
    outputs(4024) <= not((layer0_outputs(332)) and (layer0_outputs(4167)));
    outputs(4025) <= (layer0_outputs(1194)) and (layer0_outputs(2601));
    outputs(4026) <= layer0_outputs(4866);
    outputs(4027) <= not(layer0_outputs(1207));
    outputs(4028) <= layer0_outputs(3011);
    outputs(4029) <= layer0_outputs(4464);
    outputs(4030) <= not((layer0_outputs(2066)) xor (layer0_outputs(1460)));
    outputs(4031) <= (layer0_outputs(4440)) and not (layer0_outputs(3589));
    outputs(4032) <= not((layer0_outputs(1950)) xor (layer0_outputs(1819)));
    outputs(4033) <= (layer0_outputs(5012)) and not (layer0_outputs(937));
    outputs(4034) <= not((layer0_outputs(809)) or (layer0_outputs(1321)));
    outputs(4035) <= not(layer0_outputs(5111));
    outputs(4036) <= (layer0_outputs(2954)) and not (layer0_outputs(5102));
    outputs(4037) <= layer0_outputs(5107);
    outputs(4038) <= (layer0_outputs(2145)) and not (layer0_outputs(2344));
    outputs(4039) <= not(layer0_outputs(3823));
    outputs(4040) <= not(layer0_outputs(690));
    outputs(4041) <= (layer0_outputs(4235)) and not (layer0_outputs(1002));
    outputs(4042) <= not(layer0_outputs(2633));
    outputs(4043) <= not(layer0_outputs(1010));
    outputs(4044) <= not((layer0_outputs(305)) xor (layer0_outputs(3816)));
    outputs(4045) <= layer0_outputs(3621);
    outputs(4046) <= not(layer0_outputs(3112));
    outputs(4047) <= (layer0_outputs(4675)) and not (layer0_outputs(2390));
    outputs(4048) <= not(layer0_outputs(4489));
    outputs(4049) <= (layer0_outputs(847)) and not (layer0_outputs(2135));
    outputs(4050) <= layer0_outputs(3702);
    outputs(4051) <= layer0_outputs(3232);
    outputs(4052) <= not(layer0_outputs(1922));
    outputs(4053) <= (layer0_outputs(3003)) and (layer0_outputs(2222));
    outputs(4054) <= (layer0_outputs(3217)) and not (layer0_outputs(1693));
    outputs(4055) <= not(layer0_outputs(4298));
    outputs(4056) <= (layer0_outputs(242)) or (layer0_outputs(3640));
    outputs(4057) <= not(layer0_outputs(4657)) or (layer0_outputs(3545));
    outputs(4058) <= not((layer0_outputs(3170)) and (layer0_outputs(2408)));
    outputs(4059) <= (layer0_outputs(1896)) and (layer0_outputs(4877));
    outputs(4060) <= (layer0_outputs(1131)) and (layer0_outputs(135));
    outputs(4061) <= not((layer0_outputs(850)) or (layer0_outputs(2140)));
    outputs(4062) <= not((layer0_outputs(2226)) or (layer0_outputs(3306)));
    outputs(4063) <= not(layer0_outputs(2366));
    outputs(4064) <= not(layer0_outputs(628));
    outputs(4065) <= layer0_outputs(3006);
    outputs(4066) <= layer0_outputs(3760);
    outputs(4067) <= (layer0_outputs(3621)) and (layer0_outputs(3444));
    outputs(4068) <= (layer0_outputs(3341)) and not (layer0_outputs(1505));
    outputs(4069) <= (layer0_outputs(654)) and (layer0_outputs(2412));
    outputs(4070) <= layer0_outputs(1938);
    outputs(4071) <= layer0_outputs(1680);
    outputs(4072) <= not(layer0_outputs(637));
    outputs(4073) <= (layer0_outputs(346)) and not (layer0_outputs(562));
    outputs(4074) <= layer0_outputs(4673);
    outputs(4075) <= not(layer0_outputs(2548));
    outputs(4076) <= not(layer0_outputs(711)) or (layer0_outputs(646));
    outputs(4077) <= not((layer0_outputs(2936)) or (layer0_outputs(4508)));
    outputs(4078) <= not(layer0_outputs(2201));
    outputs(4079) <= (layer0_outputs(202)) xor (layer0_outputs(3142));
    outputs(4080) <= (layer0_outputs(3252)) and (layer0_outputs(1709));
    outputs(4081) <= not(layer0_outputs(4287));
    outputs(4082) <= layer0_outputs(488);
    outputs(4083) <= not(layer0_outputs(3836));
    outputs(4084) <= layer0_outputs(2626);
    outputs(4085) <= (layer0_outputs(1204)) and not (layer0_outputs(493));
    outputs(4086) <= not((layer0_outputs(1951)) or (layer0_outputs(3123)));
    outputs(4087) <= (layer0_outputs(1684)) or (layer0_outputs(3991));
    outputs(4088) <= not(layer0_outputs(2735));
    outputs(4089) <= (layer0_outputs(2087)) and not (layer0_outputs(1905));
    outputs(4090) <= not(layer0_outputs(2425));
    outputs(4091) <= not((layer0_outputs(803)) xor (layer0_outputs(1094)));
    outputs(4092) <= layer0_outputs(3327);
    outputs(4093) <= (layer0_outputs(205)) and not (layer0_outputs(3906));
    outputs(4094) <= not((layer0_outputs(2600)) xor (layer0_outputs(4300)));
    outputs(4095) <= layer0_outputs(2533);
    outputs(4096) <= layer0_outputs(4638);
    outputs(4097) <= not(layer0_outputs(1710)) or (layer0_outputs(3693));
    outputs(4098) <= (layer0_outputs(3441)) or (layer0_outputs(3854));
    outputs(4099) <= not(layer0_outputs(1703));
    outputs(4100) <= layer0_outputs(4197);
    outputs(4101) <= not(layer0_outputs(3126)) or (layer0_outputs(3147));
    outputs(4102) <= layer0_outputs(3181);
    outputs(4103) <= not((layer0_outputs(2251)) and (layer0_outputs(741)));
    outputs(4104) <= (layer0_outputs(1345)) xor (layer0_outputs(4039));
    outputs(4105) <= layer0_outputs(2561);
    outputs(4106) <= not(layer0_outputs(2272));
    outputs(4107) <= not(layer0_outputs(869));
    outputs(4108) <= (layer0_outputs(1602)) xor (layer0_outputs(3576));
    outputs(4109) <= (layer0_outputs(3856)) and not (layer0_outputs(4415));
    outputs(4110) <= not(layer0_outputs(3286)) or (layer0_outputs(627));
    outputs(4111) <= not(layer0_outputs(4018));
    outputs(4112) <= layer0_outputs(94);
    outputs(4113) <= layer0_outputs(2841);
    outputs(4114) <= not(layer0_outputs(1884)) or (layer0_outputs(2409));
    outputs(4115) <= layer0_outputs(3436);
    outputs(4116) <= layer0_outputs(4923);
    outputs(4117) <= layer0_outputs(3641);
    outputs(4118) <= not(layer0_outputs(4453)) or (layer0_outputs(4181));
    outputs(4119) <= (layer0_outputs(2018)) xor (layer0_outputs(4990));
    outputs(4120) <= not(layer0_outputs(4921));
    outputs(4121) <= not(layer0_outputs(4043)) or (layer0_outputs(1459));
    outputs(4122) <= not(layer0_outputs(1163)) or (layer0_outputs(5013));
    outputs(4123) <= (layer0_outputs(3877)) and not (layer0_outputs(2411));
    outputs(4124) <= not(layer0_outputs(610)) or (layer0_outputs(1629));
    outputs(4125) <= not(layer0_outputs(1565));
    outputs(4126) <= (layer0_outputs(433)) or (layer0_outputs(5069));
    outputs(4127) <= not(layer0_outputs(4035));
    outputs(4128) <= layer0_outputs(609);
    outputs(4129) <= layer0_outputs(1237);
    outputs(4130) <= (layer0_outputs(3395)) or (layer0_outputs(1757));
    outputs(4131) <= (layer0_outputs(2339)) or (layer0_outputs(201));
    outputs(4132) <= not(layer0_outputs(398));
    outputs(4133) <= layer0_outputs(3433);
    outputs(4134) <= not((layer0_outputs(2665)) and (layer0_outputs(3871)));
    outputs(4135) <= layer0_outputs(110);
    outputs(4136) <= not(layer0_outputs(1257));
    outputs(4137) <= not(layer0_outputs(3138));
    outputs(4138) <= not(layer0_outputs(817));
    outputs(4139) <= not(layer0_outputs(4685));
    outputs(4140) <= not(layer0_outputs(1250));
    outputs(4141) <= not(layer0_outputs(1261));
    outputs(4142) <= layer0_outputs(3202);
    outputs(4143) <= not(layer0_outputs(2736));
    outputs(4144) <= not(layer0_outputs(1605));
    outputs(4145) <= (layer0_outputs(2739)) xor (layer0_outputs(1683));
    outputs(4146) <= (layer0_outputs(2682)) and (layer0_outputs(740));
    outputs(4147) <= layer0_outputs(2848);
    outputs(4148) <= (layer0_outputs(2950)) and not (layer0_outputs(3354));
    outputs(4149) <= (layer0_outputs(3915)) or (layer0_outputs(4365));
    outputs(4150) <= not(layer0_outputs(37)) or (layer0_outputs(4745));
    outputs(4151) <= not(layer0_outputs(4091)) or (layer0_outputs(2465));
    outputs(4152) <= not(layer0_outputs(3944)) or (layer0_outputs(1158));
    outputs(4153) <= not(layer0_outputs(830)) or (layer0_outputs(4620));
    outputs(4154) <= not((layer0_outputs(2869)) and (layer0_outputs(3446)));
    outputs(4155) <= not(layer0_outputs(1138)) or (layer0_outputs(3866));
    outputs(4156) <= layer0_outputs(2407);
    outputs(4157) <= (layer0_outputs(129)) and not (layer0_outputs(4447));
    outputs(4158) <= (layer0_outputs(1596)) and (layer0_outputs(232));
    outputs(4159) <= not(layer0_outputs(2510)) or (layer0_outputs(4854));
    outputs(4160) <= not(layer0_outputs(3459));
    outputs(4161) <= (layer0_outputs(2534)) xor (layer0_outputs(1523));
    outputs(4162) <= layer0_outputs(3962);
    outputs(4163) <= layer0_outputs(2766);
    outputs(4164) <= layer0_outputs(3170);
    outputs(4165) <= (layer0_outputs(2373)) xor (layer0_outputs(1831));
    outputs(4166) <= (layer0_outputs(3230)) and (layer0_outputs(5036));
    outputs(4167) <= (layer0_outputs(3324)) and (layer0_outputs(1668));
    outputs(4168) <= not((layer0_outputs(912)) xor (layer0_outputs(3713)));
    outputs(4169) <= layer0_outputs(1985);
    outputs(4170) <= layer0_outputs(2174);
    outputs(4171) <= layer0_outputs(2658);
    outputs(4172) <= not(layer0_outputs(2332));
    outputs(4173) <= not((layer0_outputs(5015)) xor (layer0_outputs(2236)));
    outputs(4174) <= not(layer0_outputs(1728)) or (layer0_outputs(87));
    outputs(4175) <= not((layer0_outputs(2635)) and (layer0_outputs(914)));
    outputs(4176) <= layer0_outputs(3047);
    outputs(4177) <= layer0_outputs(2026);
    outputs(4178) <= not((layer0_outputs(4749)) xor (layer0_outputs(2278)));
    outputs(4179) <= not(layer0_outputs(5075)) or (layer0_outputs(2623));
    outputs(4180) <= not(layer0_outputs(2974));
    outputs(4181) <= not(layer0_outputs(4388)) or (layer0_outputs(607));
    outputs(4182) <= not(layer0_outputs(2316)) or (layer0_outputs(2006));
    outputs(4183) <= layer0_outputs(2401);
    outputs(4184) <= layer0_outputs(1760);
    outputs(4185) <= (layer0_outputs(4913)) xor (layer0_outputs(3425));
    outputs(4186) <= (layer0_outputs(2253)) and not (layer0_outputs(1148));
    outputs(4187) <= not((layer0_outputs(729)) xor (layer0_outputs(5039)));
    outputs(4188) <= layer0_outputs(4943);
    outputs(4189) <= (layer0_outputs(4398)) xor (layer0_outputs(2492));
    outputs(4190) <= not(layer0_outputs(4254));
    outputs(4191) <= (layer0_outputs(4728)) xor (layer0_outputs(4566));
    outputs(4192) <= not((layer0_outputs(252)) or (layer0_outputs(2890)));
    outputs(4193) <= layer0_outputs(4772);
    outputs(4194) <= not((layer0_outputs(4325)) or (layer0_outputs(4835)));
    outputs(4195) <= (layer0_outputs(908)) xor (layer0_outputs(2156));
    outputs(4196) <= not(layer0_outputs(688)) or (layer0_outputs(882));
    outputs(4197) <= layer0_outputs(1826);
    outputs(4198) <= not(layer0_outputs(2715)) or (layer0_outputs(2132));
    outputs(4199) <= not(layer0_outputs(668)) or (layer0_outputs(3839));
    outputs(4200) <= not(layer0_outputs(2351)) or (layer0_outputs(3426));
    outputs(4201) <= layer0_outputs(3987);
    outputs(4202) <= (layer0_outputs(2048)) and not (layer0_outputs(3238));
    outputs(4203) <= (layer0_outputs(3657)) and not (layer0_outputs(4467));
    outputs(4204) <= layer0_outputs(1135);
    outputs(4205) <= (layer0_outputs(1962)) and not (layer0_outputs(3069));
    outputs(4206) <= (layer0_outputs(1763)) and not (layer0_outputs(1290));
    outputs(4207) <= (layer0_outputs(1644)) and not (layer0_outputs(3868));
    outputs(4208) <= not(layer0_outputs(40));
    outputs(4209) <= layer0_outputs(226);
    outputs(4210) <= not(layer0_outputs(749)) or (layer0_outputs(4000));
    outputs(4211) <= (layer0_outputs(842)) and not (layer0_outputs(4743));
    outputs(4212) <= layer0_outputs(124);
    outputs(4213) <= (layer0_outputs(1932)) xor (layer0_outputs(3037));
    outputs(4214) <= (layer0_outputs(1463)) and (layer0_outputs(947));
    outputs(4215) <= layer0_outputs(2929);
    outputs(4216) <= not((layer0_outputs(1672)) or (layer0_outputs(3761)));
    outputs(4217) <= not((layer0_outputs(3689)) and (layer0_outputs(580)));
    outputs(4218) <= not((layer0_outputs(4061)) xor (layer0_outputs(4622)));
    outputs(4219) <= layer0_outputs(970);
    outputs(4220) <= not(layer0_outputs(2605)) or (layer0_outputs(1376));
    outputs(4221) <= not(layer0_outputs(857));
    outputs(4222) <= not(layer0_outputs(2710));
    outputs(4223) <= not(layer0_outputs(2589));
    outputs(4224) <= layer0_outputs(3800);
    outputs(4225) <= (layer0_outputs(4229)) or (layer0_outputs(2268));
    outputs(4226) <= layer0_outputs(2112);
    outputs(4227) <= not(layer0_outputs(722));
    outputs(4228) <= not(layer0_outputs(4502)) or (layer0_outputs(4237));
    outputs(4229) <= (layer0_outputs(4599)) and not (layer0_outputs(869));
    outputs(4230) <= layer0_outputs(3183);
    outputs(4231) <= (layer0_outputs(2977)) and not (layer0_outputs(2160));
    outputs(4232) <= (layer0_outputs(434)) xor (layer0_outputs(69));
    outputs(4233) <= not(layer0_outputs(356));
    outputs(4234) <= layer0_outputs(1888);
    outputs(4235) <= not(layer0_outputs(3018)) or (layer0_outputs(1745));
    outputs(4236) <= layer0_outputs(2260);
    outputs(4237) <= not((layer0_outputs(2819)) xor (layer0_outputs(4875)));
    outputs(4238) <= (layer0_outputs(1890)) or (layer0_outputs(658));
    outputs(4239) <= (layer0_outputs(525)) or (layer0_outputs(3147));
    outputs(4240) <= not(layer0_outputs(386)) or (layer0_outputs(1648));
    outputs(4241) <= (layer0_outputs(1800)) and not (layer0_outputs(531));
    outputs(4242) <= not(layer0_outputs(1172));
    outputs(4243) <= layer0_outputs(855);
    outputs(4244) <= not(layer0_outputs(2207));
    outputs(4245) <= layer0_outputs(685);
    outputs(4246) <= not(layer0_outputs(2927)) or (layer0_outputs(2247));
    outputs(4247) <= (layer0_outputs(3106)) or (layer0_outputs(317));
    outputs(4248) <= not((layer0_outputs(2294)) xor (layer0_outputs(2031)));
    outputs(4249) <= not(layer0_outputs(1437)) or (layer0_outputs(3240));
    outputs(4250) <= not(layer0_outputs(1645));
    outputs(4251) <= (layer0_outputs(697)) xor (layer0_outputs(2393));
    outputs(4252) <= layer0_outputs(1104);
    outputs(4253) <= not(layer0_outputs(1062));
    outputs(4254) <= layer0_outputs(4709);
    outputs(4255) <= not(layer0_outputs(852));
    outputs(4256) <= not(layer0_outputs(4346));
    outputs(4257) <= not((layer0_outputs(620)) and (layer0_outputs(4335)));
    outputs(4258) <= not(layer0_outputs(4077)) or (layer0_outputs(1066));
    outputs(4259) <= layer0_outputs(1469);
    outputs(4260) <= (layer0_outputs(2993)) xor (layer0_outputs(4368));
    outputs(4261) <= not(layer0_outputs(3416));
    outputs(4262) <= layer0_outputs(3567);
    outputs(4263) <= layer0_outputs(3225);
    outputs(4264) <= not(layer0_outputs(2138)) or (layer0_outputs(712));
    outputs(4265) <= layer0_outputs(1301);
    outputs(4266) <= layer0_outputs(1418);
    outputs(4267) <= layer0_outputs(4517);
    outputs(4268) <= not(layer0_outputs(2671));
    outputs(4269) <= not(layer0_outputs(3040));
    outputs(4270) <= not((layer0_outputs(1312)) or (layer0_outputs(323)));
    outputs(4271) <= (layer0_outputs(1093)) xor (layer0_outputs(4391));
    outputs(4272) <= not((layer0_outputs(4303)) and (layer0_outputs(3003)));
    outputs(4273) <= layer0_outputs(2484);
    outputs(4274) <= (layer0_outputs(2853)) xor (layer0_outputs(3120));
    outputs(4275) <= (layer0_outputs(2092)) xor (layer0_outputs(4166));
    outputs(4276) <= not(layer0_outputs(2878));
    outputs(4277) <= layer0_outputs(4547);
    outputs(4278) <= not((layer0_outputs(4279)) xor (layer0_outputs(451)));
    outputs(4279) <= (layer0_outputs(3073)) or (layer0_outputs(4134));
    outputs(4280) <= not(layer0_outputs(3955)) or (layer0_outputs(1903));
    outputs(4281) <= (layer0_outputs(3424)) and not (layer0_outputs(1164));
    outputs(4282) <= not((layer0_outputs(2037)) xor (layer0_outputs(1778)));
    outputs(4283) <= layer0_outputs(410);
    outputs(4284) <= layer0_outputs(4691);
    outputs(4285) <= not((layer0_outputs(3333)) and (layer0_outputs(1999)));
    outputs(4286) <= (layer0_outputs(1357)) and (layer0_outputs(2731));
    outputs(4287) <= not(layer0_outputs(1067));
    outputs(4288) <= (layer0_outputs(4304)) and not (layer0_outputs(145));
    outputs(4289) <= (layer0_outputs(4591)) or (layer0_outputs(1809));
    outputs(4290) <= (layer0_outputs(3129)) xor (layer0_outputs(1384));
    outputs(4291) <= (layer0_outputs(871)) xor (layer0_outputs(4538));
    outputs(4292) <= (layer0_outputs(3840)) and not (layer0_outputs(3266));
    outputs(4293) <= (layer0_outputs(1408)) and (layer0_outputs(1105));
    outputs(4294) <= layer0_outputs(375);
    outputs(4295) <= not(layer0_outputs(3821));
    outputs(4296) <= layer0_outputs(1826);
    outputs(4297) <= layer0_outputs(5091);
    outputs(4298) <= not((layer0_outputs(1707)) xor (layer0_outputs(3214)));
    outputs(4299) <= (layer0_outputs(2634)) and not (layer0_outputs(785));
    outputs(4300) <= not(layer0_outputs(2555));
    outputs(4301) <= (layer0_outputs(3400)) and (layer0_outputs(4430));
    outputs(4302) <= not(layer0_outputs(5088));
    outputs(4303) <= (layer0_outputs(58)) or (layer0_outputs(3200));
    outputs(4304) <= (layer0_outputs(5023)) and (layer0_outputs(1410));
    outputs(4305) <= (layer0_outputs(1973)) and (layer0_outputs(195));
    outputs(4306) <= layer0_outputs(1601);
    outputs(4307) <= not(layer0_outputs(3131));
    outputs(4308) <= not(layer0_outputs(2571));
    outputs(4309) <= (layer0_outputs(4138)) or (layer0_outputs(1438));
    outputs(4310) <= layer0_outputs(1676);
    outputs(4311) <= (layer0_outputs(1772)) or (layer0_outputs(1304));
    outputs(4312) <= (layer0_outputs(3392)) or (layer0_outputs(63));
    outputs(4313) <= not(layer0_outputs(3586));
    outputs(4314) <= (layer0_outputs(261)) xor (layer0_outputs(3457));
    outputs(4315) <= (layer0_outputs(703)) and not (layer0_outputs(4803));
    outputs(4316) <= (layer0_outputs(4847)) and (layer0_outputs(2542));
    outputs(4317) <= layer0_outputs(4288);
    outputs(4318) <= (layer0_outputs(2461)) or (layer0_outputs(3156));
    outputs(4319) <= not((layer0_outputs(197)) xor (layer0_outputs(1238)));
    outputs(4320) <= not((layer0_outputs(4684)) and (layer0_outputs(4759)));
    outputs(4321) <= not(layer0_outputs(443));
    outputs(4322) <= (layer0_outputs(2725)) and not (layer0_outputs(881));
    outputs(4323) <= layer0_outputs(1288);
    outputs(4324) <= (layer0_outputs(938)) or (layer0_outputs(1980));
    outputs(4325) <= (layer0_outputs(3482)) or (layer0_outputs(856));
    outputs(4326) <= not(layer0_outputs(241));
    outputs(4327) <= (layer0_outputs(42)) xor (layer0_outputs(298));
    outputs(4328) <= (layer0_outputs(2022)) and not (layer0_outputs(1449));
    outputs(4329) <= not((layer0_outputs(2804)) xor (layer0_outputs(1542)));
    outputs(4330) <= (layer0_outputs(2492)) xor (layer0_outputs(601));
    outputs(4331) <= not((layer0_outputs(557)) and (layer0_outputs(4724)));
    outputs(4332) <= (layer0_outputs(6)) xor (layer0_outputs(4139));
    outputs(4333) <= not(layer0_outputs(2043));
    outputs(4334) <= layer0_outputs(330);
    outputs(4335) <= layer0_outputs(175);
    outputs(4336) <= not(layer0_outputs(1320));
    outputs(4337) <= layer0_outputs(786);
    outputs(4338) <= not(layer0_outputs(822)) or (layer0_outputs(446));
    outputs(4339) <= not(layer0_outputs(3065)) or (layer0_outputs(3447));
    outputs(4340) <= not(layer0_outputs(2259)) or (layer0_outputs(495));
    outputs(4341) <= not(layer0_outputs(4587));
    outputs(4342) <= not(layer0_outputs(522)) or (layer0_outputs(383));
    outputs(4343) <= not(layer0_outputs(4584)) or (layer0_outputs(0));
    outputs(4344) <= not((layer0_outputs(3788)) xor (layer0_outputs(2840)));
    outputs(4345) <= not(layer0_outputs(951)) or (layer0_outputs(3720));
    outputs(4346) <= not(layer0_outputs(2711));
    outputs(4347) <= not((layer0_outputs(1377)) or (layer0_outputs(131)));
    outputs(4348) <= layer0_outputs(1870);
    outputs(4349) <= (layer0_outputs(2133)) and (layer0_outputs(1418));
    outputs(4350) <= not((layer0_outputs(867)) xor (layer0_outputs(3656)));
    outputs(4351) <= not(layer0_outputs(4090));
    outputs(4352) <= layer0_outputs(2057);
    outputs(4353) <= not(layer0_outputs(4570));
    outputs(4354) <= not((layer0_outputs(1571)) xor (layer0_outputs(28)));
    outputs(4355) <= not(layer0_outputs(3275));
    outputs(4356) <= layer0_outputs(1974);
    outputs(4357) <= (layer0_outputs(873)) and (layer0_outputs(585));
    outputs(4358) <= layer0_outputs(2591);
    outputs(4359) <= not(layer0_outputs(3706));
    outputs(4360) <= not((layer0_outputs(1473)) or (layer0_outputs(290)));
    outputs(4361) <= not(layer0_outputs(4502)) or (layer0_outputs(835));
    outputs(4362) <= layer0_outputs(1050);
    outputs(4363) <= not(layer0_outputs(377));
    outputs(4364) <= not(layer0_outputs(3134));
    outputs(4365) <= (layer0_outputs(4216)) or (layer0_outputs(609));
    outputs(4366) <= not(layer0_outputs(4683)) or (layer0_outputs(110));
    outputs(4367) <= not(layer0_outputs(397));
    outputs(4368) <= not(layer0_outputs(5002));
    outputs(4369) <= (layer0_outputs(3412)) and not (layer0_outputs(2403));
    outputs(4370) <= (layer0_outputs(4661)) xor (layer0_outputs(3790));
    outputs(4371) <= not(layer0_outputs(1513)) or (layer0_outputs(4659));
    outputs(4372) <= layer0_outputs(3700);
    outputs(4373) <= not((layer0_outputs(93)) xor (layer0_outputs(4520)));
    outputs(4374) <= (layer0_outputs(4228)) or (layer0_outputs(3648));
    outputs(4375) <= (layer0_outputs(2101)) and not (layer0_outputs(3584));
    outputs(4376) <= not((layer0_outputs(4029)) xor (layer0_outputs(2285)));
    outputs(4377) <= (layer0_outputs(2870)) and not (layer0_outputs(2027));
    outputs(4378) <= layer0_outputs(4690);
    outputs(4379) <= not(layer0_outputs(1575));
    outputs(4380) <= layer0_outputs(888);
    outputs(4381) <= layer0_outputs(3323);
    outputs(4382) <= layer0_outputs(3719);
    outputs(4383) <= (layer0_outputs(2999)) and not (layer0_outputs(4613));
    outputs(4384) <= layer0_outputs(600);
    outputs(4385) <= layer0_outputs(2577);
    outputs(4386) <= not(layer0_outputs(5085));
    outputs(4387) <= (layer0_outputs(4983)) and (layer0_outputs(1110));
    outputs(4388) <= not((layer0_outputs(3680)) xor (layer0_outputs(3351)));
    outputs(4389) <= layer0_outputs(2755);
    outputs(4390) <= (layer0_outputs(1287)) or (layer0_outputs(2965));
    outputs(4391) <= (layer0_outputs(4233)) and not (layer0_outputs(215));
    outputs(4392) <= not(layer0_outputs(1954));
    outputs(4393) <= not(layer0_outputs(2347));
    outputs(4394) <= (layer0_outputs(239)) and not (layer0_outputs(650));
    outputs(4395) <= (layer0_outputs(1548)) and (layer0_outputs(1925));
    outputs(4396) <= not(layer0_outputs(4670)) or (layer0_outputs(2787));
    outputs(4397) <= not(layer0_outputs(1674));
    outputs(4398) <= layer0_outputs(4387);
    outputs(4399) <= not(layer0_outputs(2568));
    outputs(4400) <= (layer0_outputs(4203)) and not (layer0_outputs(3718));
    outputs(4401) <= (layer0_outputs(1089)) or (layer0_outputs(1481));
    outputs(4402) <= layer0_outputs(52);
    outputs(4403) <= layer0_outputs(1545);
    outputs(4404) <= not(layer0_outputs(1551));
    outputs(4405) <= not((layer0_outputs(1547)) xor (layer0_outputs(999)));
    outputs(4406) <= (layer0_outputs(4064)) or (layer0_outputs(2884));
    outputs(4407) <= not(layer0_outputs(4775));
    outputs(4408) <= layer0_outputs(3774);
    outputs(4409) <= layer0_outputs(231);
    outputs(4410) <= layer0_outputs(1335);
    outputs(4411) <= not((layer0_outputs(3667)) xor (layer0_outputs(4445)));
    outputs(4412) <= layer0_outputs(4469);
    outputs(4413) <= not(layer0_outputs(1887));
    outputs(4414) <= layer0_outputs(3599);
    outputs(4415) <= not((layer0_outputs(2410)) xor (layer0_outputs(1487)));
    outputs(4416) <= (layer0_outputs(2256)) xor (layer0_outputs(690));
    outputs(4417) <= layer0_outputs(3057);
    outputs(4418) <= not((layer0_outputs(3166)) xor (layer0_outputs(4573)));
    outputs(4419) <= (layer0_outputs(4908)) and not (layer0_outputs(2790));
    outputs(4420) <= layer0_outputs(849);
    outputs(4421) <= not(layer0_outputs(2039));
    outputs(4422) <= not((layer0_outputs(791)) and (layer0_outputs(3153)));
    outputs(4423) <= not(layer0_outputs(3841)) or (layer0_outputs(1885));
    outputs(4424) <= (layer0_outputs(1078)) xor (layer0_outputs(3013));
    outputs(4425) <= not((layer0_outputs(2955)) xor (layer0_outputs(3178)));
    outputs(4426) <= (layer0_outputs(4539)) and (layer0_outputs(4124));
    outputs(4427) <= not(layer0_outputs(1081));
    outputs(4428) <= layer0_outputs(472);
    outputs(4429) <= (layer0_outputs(4999)) xor (layer0_outputs(4051));
    outputs(4430) <= layer0_outputs(1953);
    outputs(4431) <= (layer0_outputs(616)) xor (layer0_outputs(340));
    outputs(4432) <= (layer0_outputs(3474)) and not (layer0_outputs(1972));
    outputs(4433) <= not(layer0_outputs(155));
    outputs(4434) <= (layer0_outputs(4005)) xor (layer0_outputs(2371));
    outputs(4435) <= not(layer0_outputs(1222));
    outputs(4436) <= not(layer0_outputs(889));
    outputs(4437) <= (layer0_outputs(2176)) and (layer0_outputs(3890));
    outputs(4438) <= not(layer0_outputs(733));
    outputs(4439) <= (layer0_outputs(1976)) and not (layer0_outputs(3287));
    outputs(4440) <= not((layer0_outputs(1967)) and (layer0_outputs(2010)));
    outputs(4441) <= not(layer0_outputs(2340)) or (layer0_outputs(4928));
    outputs(4442) <= not((layer0_outputs(4877)) or (layer0_outputs(1941)));
    outputs(4443) <= not((layer0_outputs(3265)) and (layer0_outputs(4291)));
    outputs(4444) <= not((layer0_outputs(1650)) xor (layer0_outputs(376)));
    outputs(4445) <= not(layer0_outputs(4262));
    outputs(4446) <= layer0_outputs(4925);
    outputs(4447) <= not(layer0_outputs(1033));
    outputs(4448) <= layer0_outputs(4628);
    outputs(4449) <= (layer0_outputs(3528)) and not (layer0_outputs(4845));
    outputs(4450) <= (layer0_outputs(1152)) xor (layer0_outputs(2608));
    outputs(4451) <= not((layer0_outputs(961)) and (layer0_outputs(3088)));
    outputs(4452) <= (layer0_outputs(3025)) xor (layer0_outputs(1482));
    outputs(4453) <= not(layer0_outputs(3113));
    outputs(4454) <= layer0_outputs(3324);
    outputs(4455) <= layer0_outputs(1662);
    outputs(4456) <= not((layer0_outputs(5024)) or (layer0_outputs(4997)));
    outputs(4457) <= not(layer0_outputs(3471));
    outputs(4458) <= not(layer0_outputs(745)) or (layer0_outputs(2895));
    outputs(4459) <= not(layer0_outputs(475)) or (layer0_outputs(2834));
    outputs(4460) <= not((layer0_outputs(2896)) xor (layer0_outputs(949)));
    outputs(4461) <= not((layer0_outputs(2130)) xor (layer0_outputs(2282)));
    outputs(4462) <= layer0_outputs(178);
    outputs(4463) <= (layer0_outputs(95)) and (layer0_outputs(1044));
    outputs(4464) <= layer0_outputs(3363);
    outputs(4465) <= not(layer0_outputs(2711)) or (layer0_outputs(2586));
    outputs(4466) <= not(layer0_outputs(4032));
    outputs(4467) <= layer0_outputs(4874);
    outputs(4468) <= layer0_outputs(892);
    outputs(4469) <= layer0_outputs(1340);
    outputs(4470) <= not((layer0_outputs(3331)) xor (layer0_outputs(1934)));
    outputs(4471) <= (layer0_outputs(348)) or (layer0_outputs(3300));
    outputs(4472) <= not((layer0_outputs(2172)) and (layer0_outputs(4355)));
    outputs(4473) <= layer0_outputs(1456);
    outputs(4474) <= not(layer0_outputs(4509));
    outputs(4475) <= not((layer0_outputs(3838)) or (layer0_outputs(1431)));
    outputs(4476) <= (layer0_outputs(3422)) xor (layer0_outputs(4842));
    outputs(4477) <= not((layer0_outputs(2677)) xor (layer0_outputs(86)));
    outputs(4478) <= layer0_outputs(1855);
    outputs(4479) <= (layer0_outputs(4764)) and not (layer0_outputs(3519));
    outputs(4480) <= not(layer0_outputs(2510)) or (layer0_outputs(3057));
    outputs(4481) <= not(layer0_outputs(3609));
    outputs(4482) <= layer0_outputs(1522);
    outputs(4483) <= not((layer0_outputs(3927)) or (layer0_outputs(4071)));
    outputs(4484) <= (layer0_outputs(566)) xor (layer0_outputs(260));
    outputs(4485) <= (layer0_outputs(3378)) or (layer0_outputs(5003));
    outputs(4486) <= not(layer0_outputs(1466)) or (layer0_outputs(1147));
    outputs(4487) <= not(layer0_outputs(917));
    outputs(4488) <= not(layer0_outputs(2846)) or (layer0_outputs(3141));
    outputs(4489) <= (layer0_outputs(1597)) xor (layer0_outputs(4762));
    outputs(4490) <= not(layer0_outputs(547)) or (layer0_outputs(2108));
    outputs(4491) <= (layer0_outputs(2045)) xor (layer0_outputs(111));
    outputs(4492) <= not((layer0_outputs(4737)) xor (layer0_outputs(4214)));
    outputs(4493) <= not((layer0_outputs(2223)) xor (layer0_outputs(4321)));
    outputs(4494) <= layer0_outputs(1404);
    outputs(4495) <= not(layer0_outputs(2314));
    outputs(4496) <= (layer0_outputs(1690)) and not (layer0_outputs(1702));
    outputs(4497) <= layer0_outputs(229);
    outputs(4498) <= not((layer0_outputs(3091)) or (layer0_outputs(4986)));
    outputs(4499) <= not((layer0_outputs(1862)) xor (layer0_outputs(1130)));
    outputs(4500) <= not(layer0_outputs(1437));
    outputs(4501) <= layer0_outputs(515);
    outputs(4502) <= not((layer0_outputs(549)) or (layer0_outputs(634)));
    outputs(4503) <= (layer0_outputs(4560)) xor (layer0_outputs(243));
    outputs(4504) <= layer0_outputs(1232);
    outputs(4505) <= (layer0_outputs(4755)) and not (layer0_outputs(193));
    outputs(4506) <= not(layer0_outputs(289)) or (layer0_outputs(3889));
    outputs(4507) <= layer0_outputs(1508);
    outputs(4508) <= not((layer0_outputs(2289)) xor (layer0_outputs(1636)));
    outputs(4509) <= layer0_outputs(1754);
    outputs(4510) <= layer0_outputs(1378);
    outputs(4511) <= (layer0_outputs(267)) or (layer0_outputs(1307));
    outputs(4512) <= not((layer0_outputs(4807)) and (layer0_outputs(3911)));
    outputs(4513) <= layer0_outputs(3800);
    outputs(4514) <= not(layer0_outputs(257)) or (layer0_outputs(2938));
    outputs(4515) <= (layer0_outputs(412)) xor (layer0_outputs(1447));
    outputs(4516) <= not((layer0_outputs(4975)) xor (layer0_outputs(3799)));
    outputs(4517) <= not(layer0_outputs(4548));
    outputs(4518) <= layer0_outputs(4089);
    outputs(4519) <= (layer0_outputs(2879)) xor (layer0_outputs(3605));
    outputs(4520) <= not(layer0_outputs(176));
    outputs(4521) <= not(layer0_outputs(2325)) or (layer0_outputs(433));
    outputs(4522) <= not((layer0_outputs(3573)) and (layer0_outputs(4397)));
    outputs(4523) <= not(layer0_outputs(4463));
    outputs(4524) <= (layer0_outputs(3086)) and not (layer0_outputs(306));
    outputs(4525) <= (layer0_outputs(3409)) xor (layer0_outputs(3602));
    outputs(4526) <= not(layer0_outputs(3364));
    outputs(4527) <= not(layer0_outputs(3470)) or (layer0_outputs(2908));
    outputs(4528) <= not((layer0_outputs(50)) xor (layer0_outputs(732)));
    outputs(4529) <= (layer0_outputs(665)) xor (layer0_outputs(3767));
    outputs(4530) <= (layer0_outputs(291)) and not (layer0_outputs(5098));
    outputs(4531) <= not(layer0_outputs(4909));
    outputs(4532) <= (layer0_outputs(4750)) or (layer0_outputs(3774));
    outputs(4533) <= not(layer0_outputs(775));
    outputs(4534) <= not(layer0_outputs(1830));
    outputs(4535) <= not(layer0_outputs(2114));
    outputs(4536) <= not(layer0_outputs(4373));
    outputs(4537) <= not((layer0_outputs(2565)) and (layer0_outputs(200)));
    outputs(4538) <= not(layer0_outputs(943)) or (layer0_outputs(1981));
    outputs(4539) <= (layer0_outputs(3722)) xor (layer0_outputs(3169));
    outputs(4540) <= layer0_outputs(1931);
    outputs(4541) <= not((layer0_outputs(2302)) and (layer0_outputs(2286)));
    outputs(4542) <= layer0_outputs(2979);
    outputs(4543) <= (layer0_outputs(3227)) and not (layer0_outputs(279));
    outputs(4544) <= not((layer0_outputs(1482)) xor (layer0_outputs(2454)));
    outputs(4545) <= layer0_outputs(662);
    outputs(4546) <= (layer0_outputs(3387)) xor (layer0_outputs(75));
    outputs(4547) <= layer0_outputs(1690);
    outputs(4548) <= layer0_outputs(810);
    outputs(4549) <= not(layer0_outputs(4088));
    outputs(4550) <= not(layer0_outputs(4834));
    outputs(4551) <= not(layer0_outputs(414));
    outputs(4552) <= (layer0_outputs(4157)) and (layer0_outputs(2676));
    outputs(4553) <= not(layer0_outputs(56)) or (layer0_outputs(724));
    outputs(4554) <= layer0_outputs(1365);
    outputs(4555) <= (layer0_outputs(582)) and (layer0_outputs(4393));
    outputs(4556) <= not((layer0_outputs(3376)) xor (layer0_outputs(4427)));
    outputs(4557) <= layer0_outputs(2257);
    outputs(4558) <= (layer0_outputs(2991)) and not (layer0_outputs(3633));
    outputs(4559) <= not(layer0_outputs(1682));
    outputs(4560) <= (layer0_outputs(1351)) and not (layer0_outputs(1671));
    outputs(4561) <= layer0_outputs(3058);
    outputs(4562) <= not(layer0_outputs(2295));
    outputs(4563) <= not(layer0_outputs(3383)) or (layer0_outputs(935));
    outputs(4564) <= (layer0_outputs(461)) and not (layer0_outputs(3937));
    outputs(4565) <= not(layer0_outputs(2939));
    outputs(4566) <= not(layer0_outputs(3592));
    outputs(4567) <= (layer0_outputs(3735)) or (layer0_outputs(4589));
    outputs(4568) <= layer0_outputs(3183);
    outputs(4569) <= (layer0_outputs(1903)) xor (layer0_outputs(4714));
    outputs(4570) <= (layer0_outputs(3532)) and (layer0_outputs(3414));
    outputs(4571) <= not(layer0_outputs(640));
    outputs(4572) <= layer0_outputs(2656);
    outputs(4573) <= layer0_outputs(2075);
    outputs(4574) <= (layer0_outputs(4524)) and not (layer0_outputs(3051));
    outputs(4575) <= not((layer0_outputs(1112)) and (layer0_outputs(3256)));
    outputs(4576) <= layer0_outputs(4058);
    outputs(4577) <= not(layer0_outputs(4001));
    outputs(4578) <= not(layer0_outputs(553));
    outputs(4579) <= (layer0_outputs(1802)) and not (layer0_outputs(183));
    outputs(4580) <= not(layer0_outputs(3811));
    outputs(4581) <= (layer0_outputs(1407)) xor (layer0_outputs(3460));
    outputs(4582) <= not((layer0_outputs(1358)) and (layer0_outputs(837)));
    outputs(4583) <= not((layer0_outputs(2684)) xor (layer0_outputs(1708)));
    outputs(4584) <= (layer0_outputs(3295)) xor (layer0_outputs(799));
    outputs(4585) <= not((layer0_outputs(3019)) xor (layer0_outputs(1101)));
    outputs(4586) <= not((layer0_outputs(2348)) xor (layer0_outputs(4883)));
    outputs(4587) <= not(layer0_outputs(2370));
    outputs(4588) <= layer0_outputs(584);
    outputs(4589) <= not(layer0_outputs(1106));
    outputs(4590) <= not(layer0_outputs(3107));
    outputs(4591) <= layer0_outputs(2003);
    outputs(4592) <= not(layer0_outputs(3753)) or (layer0_outputs(4010));
    outputs(4593) <= not(layer0_outputs(404));
    outputs(4594) <= not(layer0_outputs(1235));
    outputs(4595) <= (layer0_outputs(932)) xor (layer0_outputs(2513));
    outputs(4596) <= not((layer0_outputs(1443)) xor (layer0_outputs(4353)));
    outputs(4597) <= (layer0_outputs(1265)) or (layer0_outputs(181));
    outputs(4598) <= not((layer0_outputs(3901)) xor (layer0_outputs(4929)));
    outputs(4599) <= (layer0_outputs(1450)) and (layer0_outputs(508));
    outputs(4600) <= not(layer0_outputs(1666)) or (layer0_outputs(2176));
    outputs(4601) <= not(layer0_outputs(372)) or (layer0_outputs(4073));
    outputs(4602) <= not((layer0_outputs(1214)) xor (layer0_outputs(4150)));
    outputs(4603) <= layer0_outputs(1541);
    outputs(4604) <= layer0_outputs(3489);
    outputs(4605) <= not((layer0_outputs(38)) or (layer0_outputs(766)));
    outputs(4606) <= not((layer0_outputs(4195)) and (layer0_outputs(2615)));
    outputs(4607) <= not(layer0_outputs(1213)) or (layer0_outputs(2948));
    outputs(4608) <= (layer0_outputs(2358)) xor (layer0_outputs(4143));
    outputs(4609) <= (layer0_outputs(2741)) and (layer0_outputs(1341));
    outputs(4610) <= not((layer0_outputs(3395)) xor (layer0_outputs(1856)));
    outputs(4611) <= layer0_outputs(3127);
    outputs(4612) <= (layer0_outputs(4569)) and (layer0_outputs(4324));
    outputs(4613) <= layer0_outputs(3943);
    outputs(4614) <= not((layer0_outputs(338)) and (layer0_outputs(425)));
    outputs(4615) <= (layer0_outputs(4901)) and not (layer0_outputs(2210));
    outputs(4616) <= (layer0_outputs(341)) and not (layer0_outputs(1354));
    outputs(4617) <= not((layer0_outputs(3679)) or (layer0_outputs(3822)));
    outputs(4618) <= layer0_outputs(2225);
    outputs(4619) <= not((layer0_outputs(5118)) xor (layer0_outputs(3029)));
    outputs(4620) <= (layer0_outputs(2942)) and (layer0_outputs(953));
    outputs(4621) <= not((layer0_outputs(1091)) or (layer0_outputs(4072)));
    outputs(4622) <= (layer0_outputs(710)) and (layer0_outputs(971));
    outputs(4623) <= layer0_outputs(432);
    outputs(4624) <= not(layer0_outputs(2758));
    outputs(4625) <= layer0_outputs(1241);
    outputs(4626) <= (layer0_outputs(5096)) and not (layer0_outputs(1649));
    outputs(4627) <= (layer0_outputs(2580)) and not (layer0_outputs(3046));
    outputs(4628) <= (layer0_outputs(1678)) xor (layer0_outputs(5083));
    outputs(4629) <= not(layer0_outputs(1329));
    outputs(4630) <= layer0_outputs(2901);
    outputs(4631) <= not(layer0_outputs(4725));
    outputs(4632) <= not(layer0_outputs(3082));
    outputs(4633) <= layer0_outputs(4402);
    outputs(4634) <= not(layer0_outputs(137));
    outputs(4635) <= (layer0_outputs(3664)) and not (layer0_outputs(980));
    outputs(4636) <= not(layer0_outputs(4343));
    outputs(4637) <= (layer0_outputs(5111)) and not (layer0_outputs(3488));
    outputs(4638) <= not((layer0_outputs(2201)) and (layer0_outputs(972)));
    outputs(4639) <= (layer0_outputs(1477)) and not (layer0_outputs(1959));
    outputs(4640) <= layer0_outputs(2475);
    outputs(4641) <= (layer0_outputs(1559)) and (layer0_outputs(929));
    outputs(4642) <= layer0_outputs(4365);
    outputs(4643) <= layer0_outputs(4964);
    outputs(4644) <= not((layer0_outputs(2820)) xor (layer0_outputs(1471)));
    outputs(4645) <= (layer0_outputs(2573)) and not (layer0_outputs(478));
    outputs(4646) <= not(layer0_outputs(1549));
    outputs(4647) <= layer0_outputs(504);
    outputs(4648) <= not((layer0_outputs(2107)) or (layer0_outputs(3260)));
    outputs(4649) <= (layer0_outputs(3986)) and not (layer0_outputs(3650));
    outputs(4650) <= not(layer0_outputs(4527));
    outputs(4651) <= not(layer0_outputs(852));
    outputs(4652) <= not(layer0_outputs(1869)) or (layer0_outputs(2490));
    outputs(4653) <= (layer0_outputs(4800)) and (layer0_outputs(1995));
    outputs(4654) <= not((layer0_outputs(2350)) or (layer0_outputs(718)));
    outputs(4655) <= not(layer0_outputs(3558));
    outputs(4656) <= layer0_outputs(3863);
    outputs(4657) <= not(layer0_outputs(1921));
    outputs(4658) <= not((layer0_outputs(2204)) or (layer0_outputs(3677)));
    outputs(4659) <= not(layer0_outputs(551));
    outputs(4660) <= not(layer0_outputs(3782));
    outputs(4661) <= not(layer0_outputs(2131));
    outputs(4662) <= not((layer0_outputs(2535)) xor (layer0_outputs(1168)));
    outputs(4663) <= (layer0_outputs(2337)) and not (layer0_outputs(2907));
    outputs(4664) <= layer0_outputs(1838);
    outputs(4665) <= not(layer0_outputs(3567));
    outputs(4666) <= (layer0_outputs(2948)) and not (layer0_outputs(3137));
    outputs(4667) <= (layer0_outputs(920)) and not (layer0_outputs(4752));
    outputs(4668) <= not(layer0_outputs(5080));
    outputs(4669) <= (layer0_outputs(1027)) and not (layer0_outputs(715));
    outputs(4670) <= not((layer0_outputs(2213)) or (layer0_outputs(5004)));
    outputs(4671) <= not(layer0_outputs(441));
    outputs(4672) <= (layer0_outputs(1381)) and not (layer0_outputs(3083));
    outputs(4673) <= not((layer0_outputs(1492)) xor (layer0_outputs(3916)));
    outputs(4674) <= (layer0_outputs(3665)) and (layer0_outputs(971));
    outputs(4675) <= not((layer0_outputs(4897)) and (layer0_outputs(714)));
    outputs(4676) <= (layer0_outputs(2670)) and not (layer0_outputs(2932));
    outputs(4677) <= not(layer0_outputs(1563));
    outputs(4678) <= layer0_outputs(4938);
    outputs(4679) <= (layer0_outputs(3355)) xor (layer0_outputs(3617));
    outputs(4680) <= not(layer0_outputs(2692));
    outputs(4681) <= not(layer0_outputs(1452));
    outputs(4682) <= layer0_outputs(977);
    outputs(4683) <= (layer0_outputs(3087)) and not (layer0_outputs(2290));
    outputs(4684) <= not((layer0_outputs(554)) xor (layer0_outputs(1891)));
    outputs(4685) <= (layer0_outputs(1628)) and not (layer0_outputs(2458));
    outputs(4686) <= not(layer0_outputs(2288));
    outputs(4687) <= not((layer0_outputs(3827)) or (layer0_outputs(1945)));
    outputs(4688) <= layer0_outputs(391);
    outputs(4689) <= layer0_outputs(2098);
    outputs(4690) <= layer0_outputs(891);
    outputs(4691) <= not(layer0_outputs(1382));
    outputs(4692) <= not((layer0_outputs(3034)) xor (layer0_outputs(241)));
    outputs(4693) <= not(layer0_outputs(2900));
    outputs(4694) <= (layer0_outputs(4149)) xor (layer0_outputs(559));
    outputs(4695) <= layer0_outputs(3222);
    outputs(4696) <= not((layer0_outputs(2557)) or (layer0_outputs(823)));
    outputs(4697) <= (layer0_outputs(2487)) and not (layer0_outputs(527));
    outputs(4698) <= not((layer0_outputs(718)) or (layer0_outputs(4839)));
    outputs(4699) <= layer0_outputs(4518);
    outputs(4700) <= not(layer0_outputs(3043));
    outputs(4701) <= not((layer0_outputs(2738)) xor (layer0_outputs(4144)));
    outputs(4702) <= layer0_outputs(1992);
    outputs(4703) <= not(layer0_outputs(1179));
    outputs(4704) <= layer0_outputs(3019);
    outputs(4705) <= (layer0_outputs(2091)) and not (layer0_outputs(4930));
    outputs(4706) <= not((layer0_outputs(4168)) xor (layer0_outputs(2169)));
    outputs(4707) <= not(layer0_outputs(4357));
    outputs(4708) <= (layer0_outputs(2645)) and not (layer0_outputs(1368));
    outputs(4709) <= (layer0_outputs(1887)) and (layer0_outputs(3377));
    outputs(4710) <= not((layer0_outputs(4066)) or (layer0_outputs(1362)));
    outputs(4711) <= (layer0_outputs(668)) and not (layer0_outputs(1023));
    outputs(4712) <= not((layer0_outputs(1114)) xor (layer0_outputs(4993)));
    outputs(4713) <= layer0_outputs(872);
    outputs(4714) <= (layer0_outputs(2173)) and not (layer0_outputs(3315));
    outputs(4715) <= not(layer0_outputs(1848));
    outputs(4716) <= not((layer0_outputs(420)) and (layer0_outputs(1647)));
    outputs(4717) <= (layer0_outputs(4835)) or (layer0_outputs(4182));
    outputs(4718) <= (layer0_outputs(1810)) and not (layer0_outputs(4174));
    outputs(4719) <= (layer0_outputs(3340)) xor (layer0_outputs(545));
    outputs(4720) <= not((layer0_outputs(327)) xor (layer0_outputs(104)));
    outputs(4721) <= not(layer0_outputs(2241));
    outputs(4722) <= layer0_outputs(2262);
    outputs(4723) <= (layer0_outputs(4744)) and (layer0_outputs(3229));
    outputs(4724) <= (layer0_outputs(2368)) xor (layer0_outputs(3885));
    outputs(4725) <= layer0_outputs(4280);
    outputs(4726) <= layer0_outputs(2925);
    outputs(4727) <= not((layer0_outputs(786)) xor (layer0_outputs(5038)));
    outputs(4728) <= not(layer0_outputs(1745));
    outputs(4729) <= not(layer0_outputs(3701));
    outputs(4730) <= (layer0_outputs(54)) and (layer0_outputs(156));
    outputs(4731) <= (layer0_outputs(940)) and not (layer0_outputs(4397));
    outputs(4732) <= not(layer0_outputs(2068));
    outputs(4733) <= not((layer0_outputs(3040)) or (layer0_outputs(4127)));
    outputs(4734) <= layer0_outputs(4476);
    outputs(4735) <= not(layer0_outputs(4022));
    outputs(4736) <= not((layer0_outputs(589)) and (layer0_outputs(4878)));
    outputs(4737) <= (layer0_outputs(3686)) and not (layer0_outputs(4116));
    outputs(4738) <= (layer0_outputs(4147)) and (layer0_outputs(1914));
    outputs(4739) <= layer0_outputs(389);
    outputs(4740) <= layer0_outputs(4794);
    outputs(4741) <= not((layer0_outputs(3321)) or (layer0_outputs(2188)));
    outputs(4742) <= not(layer0_outputs(400));
    outputs(4743) <= layer0_outputs(3627);
    outputs(4744) <= (layer0_outputs(3830)) and not (layer0_outputs(2849));
    outputs(4745) <= layer0_outputs(839);
    outputs(4746) <= layer0_outputs(1889);
    outputs(4747) <= not((layer0_outputs(66)) or (layer0_outputs(3031)));
    outputs(4748) <= not(layer0_outputs(4677));
    outputs(4749) <= (layer0_outputs(3732)) and (layer0_outputs(2376));
    outputs(4750) <= not(layer0_outputs(1100)) or (layer0_outputs(3881));
    outputs(4751) <= not(layer0_outputs(4607));
    outputs(4752) <= not(layer0_outputs(3004));
    outputs(4753) <= (layer0_outputs(421)) and not (layer0_outputs(21));
    outputs(4754) <= not((layer0_outputs(1277)) and (layer0_outputs(4100)));
    outputs(4755) <= layer0_outputs(3820);
    outputs(4756) <= layer0_outputs(4614);
    outputs(4757) <= not(layer0_outputs(1946)) or (layer0_outputs(2530));
    outputs(4758) <= layer0_outputs(906);
    outputs(4759) <= layer0_outputs(3087);
    outputs(4760) <= not((layer0_outputs(3966)) or (layer0_outputs(4115)));
    outputs(4761) <= (layer0_outputs(4472)) and not (layer0_outputs(4498));
    outputs(4762) <= not(layer0_outputs(1498)) or (layer0_outputs(4171));
    outputs(4763) <= not(layer0_outputs(3815));
    outputs(4764) <= not(layer0_outputs(1423));
    outputs(4765) <= not((layer0_outputs(3021)) or (layer0_outputs(4721)));
    outputs(4766) <= not(layer0_outputs(1496));
    outputs(4767) <= not((layer0_outputs(2934)) or (layer0_outputs(4293)));
    outputs(4768) <= (layer0_outputs(2529)) and not (layer0_outputs(151));
    outputs(4769) <= (layer0_outputs(3513)) and (layer0_outputs(3968));
    outputs(4770) <= not(layer0_outputs(5018));
    outputs(4771) <= not(layer0_outputs(1425)) or (layer0_outputs(4812));
    outputs(4772) <= layer0_outputs(3174);
    outputs(4773) <= (layer0_outputs(3065)) and not (layer0_outputs(3853));
    outputs(4774) <= layer0_outputs(2502);
    outputs(4775) <= layer0_outputs(3437);
    outputs(4776) <= not(layer0_outputs(3223));
    outputs(4777) <= not(layer0_outputs(3254));
    outputs(4778) <= not(layer0_outputs(85));
    outputs(4779) <= layer0_outputs(683);
    outputs(4780) <= not((layer0_outputs(1813)) xor (layer0_outputs(4574)));
    outputs(4781) <= (layer0_outputs(1028)) and not (layer0_outputs(2932));
    outputs(4782) <= not(layer0_outputs(735));
    outputs(4783) <= not(layer0_outputs(3390));
    outputs(4784) <= not(layer0_outputs(28));
    outputs(4785) <= (layer0_outputs(2054)) and (layer0_outputs(3901));
    outputs(4786) <= not((layer0_outputs(3529)) or (layer0_outputs(1595)));
    outputs(4787) <= not((layer0_outputs(290)) or (layer0_outputs(4155)));
    outputs(4788) <= (layer0_outputs(1933)) and not (layer0_outputs(2662));
    outputs(4789) <= layer0_outputs(4227);
    outputs(4790) <= not((layer0_outputs(2700)) or (layer0_outputs(1951)));
    outputs(4791) <= (layer0_outputs(3002)) and not (layer0_outputs(3966));
    outputs(4792) <= not(layer0_outputs(3953)) or (layer0_outputs(4883));
    outputs(4793) <= not(layer0_outputs(3220));
    outputs(4794) <= not((layer0_outputs(2081)) or (layer0_outputs(1733)));
    outputs(4795) <= not(layer0_outputs(1211));
    outputs(4796) <= (layer0_outputs(1689)) and not (layer0_outputs(237));
    outputs(4797) <= not(layer0_outputs(4994));
    outputs(4798) <= (layer0_outputs(1148)) and (layer0_outputs(945));
    outputs(4799) <= (layer0_outputs(1888)) xor (layer0_outputs(4858));
    outputs(4800) <= layer0_outputs(48);
    outputs(4801) <= not(layer0_outputs(2136));
    outputs(4802) <= (layer0_outputs(4988)) and not (layer0_outputs(4196));
    outputs(4803) <= (layer0_outputs(1503)) and not (layer0_outputs(4307));
    outputs(4804) <= not((layer0_outputs(1942)) or (layer0_outputs(731)));
    outputs(4805) <= not((layer0_outputs(4694)) xor (layer0_outputs(2744)));
    outputs(4806) <= (layer0_outputs(1810)) and not (layer0_outputs(4637));
    outputs(4807) <= not(layer0_outputs(4889));
    outputs(4808) <= layer0_outputs(2902);
    outputs(4809) <= (layer0_outputs(2014)) and not (layer0_outputs(3985));
    outputs(4810) <= not((layer0_outputs(1060)) xor (layer0_outputs(1766)));
    outputs(4811) <= not(layer0_outputs(1863));
    outputs(4812) <= not(layer0_outputs(2267));
    outputs(4813) <= layer0_outputs(961);
    outputs(4814) <= (layer0_outputs(2359)) and not (layer0_outputs(3668));
    outputs(4815) <= not(layer0_outputs(4644));
    outputs(4816) <= not(layer0_outputs(301));
    outputs(4817) <= not((layer0_outputs(3741)) or (layer0_outputs(4955)));
    outputs(4818) <= not(layer0_outputs(4351));
    outputs(4819) <= (layer0_outputs(1801)) and (layer0_outputs(391));
    outputs(4820) <= not((layer0_outputs(1200)) or (layer0_outputs(482)));
    outputs(4821) <= (layer0_outputs(1554)) and (layer0_outputs(1512));
    outputs(4822) <= layer0_outputs(343);
    outputs(4823) <= (layer0_outputs(405)) and (layer0_outputs(2451));
    outputs(4824) <= layer0_outputs(4090);
    outputs(4825) <= layer0_outputs(764);
    outputs(4826) <= layer0_outputs(173);
    outputs(4827) <= not((layer0_outputs(3265)) or (layer0_outputs(5029)));
    outputs(4828) <= not((layer0_outputs(245)) or (layer0_outputs(3072)));
    outputs(4829) <= layer0_outputs(925);
    outputs(4830) <= not(layer0_outputs(1603));
    outputs(4831) <= not(layer0_outputs(3095));
    outputs(4832) <= not(layer0_outputs(910));
    outputs(4833) <= not(layer0_outputs(2625));
    outputs(4834) <= not((layer0_outputs(3319)) or (layer0_outputs(2283)));
    outputs(4835) <= (layer0_outputs(3413)) and not (layer0_outputs(2309));
    outputs(4836) <= (layer0_outputs(249)) and not (layer0_outputs(1744));
    outputs(4837) <= (layer0_outputs(3118)) and (layer0_outputs(4036));
    outputs(4838) <= layer0_outputs(4079);
    outputs(4839) <= not(layer0_outputs(4688));
    outputs(4840) <= layer0_outputs(2599);
    outputs(4841) <= not((layer0_outputs(2978)) or (layer0_outputs(887)));
    outputs(4842) <= not(layer0_outputs(996));
    outputs(4843) <= (layer0_outputs(150)) and (layer0_outputs(385));
    outputs(4844) <= not(layer0_outputs(1218));
    outputs(4845) <= not(layer0_outputs(4843));
    outputs(4846) <= layer0_outputs(1271);
    outputs(4847) <= (layer0_outputs(4765)) and not (layer0_outputs(2522));
    outputs(4848) <= layer0_outputs(5014);
    outputs(4849) <= (layer0_outputs(3791)) and (layer0_outputs(1226));
    outputs(4850) <= (layer0_outputs(1346)) and (layer0_outputs(3872));
    outputs(4851) <= layer0_outputs(975);
    outputs(4852) <= layer0_outputs(2439);
    outputs(4853) <= not((layer0_outputs(336)) or (layer0_outputs(3784)));
    outputs(4854) <= (layer0_outputs(3629)) and (layer0_outputs(1626));
    outputs(4855) <= layer0_outputs(627);
    outputs(4856) <= (layer0_outputs(4998)) and not (layer0_outputs(3848));
    outputs(4857) <= not(layer0_outputs(2021)) or (layer0_outputs(2231));
    outputs(4858) <= (layer0_outputs(4564)) and (layer0_outputs(1111));
    outputs(4859) <= (layer0_outputs(772)) and not (layer0_outputs(2708));
    outputs(4860) <= not(layer0_outputs(1797));
    outputs(4861) <= (layer0_outputs(3421)) xor (layer0_outputs(4455));
    outputs(4862) <= (layer0_outputs(9)) and not (layer0_outputs(2555));
    outputs(4863) <= not(layer0_outputs(4945));
    outputs(4864) <= not(layer0_outputs(4031));
    outputs(4865) <= (layer0_outputs(4450)) and not (layer0_outputs(924));
    outputs(4866) <= (layer0_outputs(4496)) and not (layer0_outputs(770));
    outputs(4867) <= layer0_outputs(1931);
    outputs(4868) <= (layer0_outputs(3872)) and not (layer0_outputs(2473));
    outputs(4869) <= not(layer0_outputs(184));
    outputs(4870) <= layer0_outputs(1823);
    outputs(4871) <= layer0_outputs(3812);
    outputs(4872) <= not((layer0_outputs(4121)) or (layer0_outputs(2284)));
    outputs(4873) <= (layer0_outputs(2229)) and not (layer0_outputs(3172));
    outputs(4874) <= layer0_outputs(3568);
    outputs(4875) <= (layer0_outputs(753)) and not (layer0_outputs(1657));
    outputs(4876) <= not(layer0_outputs(2203)) or (layer0_outputs(4680));
    outputs(4877) <= layer0_outputs(948);
    outputs(4878) <= (layer0_outputs(3080)) and not (layer0_outputs(2369));
    outputs(4879) <= not(layer0_outputs(2448));
    outputs(4880) <= layer0_outputs(3309);
    outputs(4881) <= not(layer0_outputs(1557));
    outputs(4882) <= (layer0_outputs(510)) and (layer0_outputs(4679));
    outputs(4883) <= not((layer0_outputs(3514)) xor (layer0_outputs(941)));
    outputs(4884) <= layer0_outputs(1007);
    outputs(4885) <= (layer0_outputs(431)) and (layer0_outputs(71));
    outputs(4886) <= not(layer0_outputs(3799));
    outputs(4887) <= not((layer0_outputs(125)) or (layer0_outputs(3542)));
    outputs(4888) <= (layer0_outputs(2180)) and (layer0_outputs(534));
    outputs(4889) <= layer0_outputs(2446);
    outputs(4890) <= not((layer0_outputs(2837)) or (layer0_outputs(639)));
    outputs(4891) <= layer0_outputs(401);
    outputs(4892) <= not(layer0_outputs(1258));
    outputs(4893) <= not(layer0_outputs(270));
    outputs(4894) <= (layer0_outputs(3789)) and not (layer0_outputs(507));
    outputs(4895) <= not((layer0_outputs(2822)) or (layer0_outputs(4074)));
    outputs(4896) <= not(layer0_outputs(3539));
    outputs(4897) <= (layer0_outputs(1791)) and (layer0_outputs(2268));
    outputs(4898) <= layer0_outputs(117);
    outputs(4899) <= (layer0_outputs(218)) and not (layer0_outputs(2537));
    outputs(4900) <= not(layer0_outputs(4893));
    outputs(4901) <= layer0_outputs(4962);
    outputs(4902) <= not(layer0_outputs(2810));
    outputs(4903) <= layer0_outputs(3904);
    outputs(4904) <= not(layer0_outputs(2291));
    outputs(4905) <= layer0_outputs(5087);
    outputs(4906) <= not(layer0_outputs(1003));
    outputs(4907) <= (layer0_outputs(898)) and not (layer0_outputs(2526));
    outputs(4908) <= layer0_outputs(2765);
    outputs(4909) <= layer0_outputs(4978);
    outputs(4910) <= layer0_outputs(5050);
    outputs(4911) <= (layer0_outputs(2582)) and not (layer0_outputs(1188));
    outputs(4912) <= layer0_outputs(2562);
    outputs(4913) <= not(layer0_outputs(687)) or (layer0_outputs(4811));
    outputs(4914) <= not((layer0_outputs(2769)) xor (layer0_outputs(1480)));
    outputs(4915) <= layer0_outputs(4390);
    outputs(4916) <= layer0_outputs(3067);
    outputs(4917) <= (layer0_outputs(2180)) and (layer0_outputs(1839));
    outputs(4918) <= not(layer0_outputs(1679));
    outputs(4919) <= (layer0_outputs(3831)) and (layer0_outputs(2055));
    outputs(4920) <= not((layer0_outputs(2739)) or (layer0_outputs(2904)));
    outputs(4921) <= layer0_outputs(3902);
    outputs(4922) <= not((layer0_outputs(1090)) and (layer0_outputs(2746)));
    outputs(4923) <= not((layer0_outputs(1126)) xor (layer0_outputs(4646)));
    outputs(4924) <= (layer0_outputs(1230)) and (layer0_outputs(4275));
    outputs(4925) <= layer0_outputs(565);
    outputs(4926) <= not(layer0_outputs(3886));
    outputs(4927) <= (layer0_outputs(2418)) and not (layer0_outputs(1557));
    outputs(4928) <= (layer0_outputs(2634)) and not (layer0_outputs(107));
    outputs(4929) <= not(layer0_outputs(2281));
    outputs(4930) <= not(layer0_outputs(2146));
    outputs(4931) <= not((layer0_outputs(4609)) or (layer0_outputs(3231)));
    outputs(4932) <= layer0_outputs(783);
    outputs(4933) <= not((layer0_outputs(4829)) or (layer0_outputs(591)));
    outputs(4934) <= layer0_outputs(1133);
    outputs(4935) <= layer0_outputs(3975);
    outputs(4936) <= (layer0_outputs(4288)) and not (layer0_outputs(2682));
    outputs(4937) <= not(layer0_outputs(2531)) or (layer0_outputs(96));
    outputs(4938) <= not(layer0_outputs(3480));
    outputs(4939) <= layer0_outputs(1978);
    outputs(4940) <= not(layer0_outputs(3577));
    outputs(4941) <= (layer0_outputs(2686)) and (layer0_outputs(3360));
    outputs(4942) <= not((layer0_outputs(2351)) or (layer0_outputs(112)));
    outputs(4943) <= not((layer0_outputs(3964)) or (layer0_outputs(2397)));
    outputs(4944) <= (layer0_outputs(3612)) and not (layer0_outputs(2782));
    outputs(4945) <= (layer0_outputs(177)) and (layer0_outputs(4312));
    outputs(4946) <= (layer0_outputs(489)) or (layer0_outputs(208));
    outputs(4947) <= not(layer0_outputs(3199)) or (layer0_outputs(3185));
    outputs(4948) <= (layer0_outputs(1533)) and not (layer0_outputs(4773));
    outputs(4949) <= not(layer0_outputs(1864));
    outputs(4950) <= (layer0_outputs(461)) and not (layer0_outputs(4927));
    outputs(4951) <= (layer0_outputs(896)) xor (layer0_outputs(2043));
    outputs(4952) <= (layer0_outputs(3012)) xor (layer0_outputs(3929));
    outputs(4953) <= (layer0_outputs(1315)) and not (layer0_outputs(3970));
    outputs(4954) <= not((layer0_outputs(207)) or (layer0_outputs(1059)));
    outputs(4955) <= layer0_outputs(2018);
    outputs(4956) <= layer0_outputs(2609);
    outputs(4957) <= layer0_outputs(1628);
    outputs(4958) <= (layer0_outputs(2505)) and (layer0_outputs(2938));
    outputs(4959) <= (layer0_outputs(3363)) and not (layer0_outputs(809));
    outputs(4960) <= layer0_outputs(4368);
    outputs(4961) <= not(layer0_outputs(3751)) or (layer0_outputs(1978));
    outputs(4962) <= not(layer0_outputs(3743));
    outputs(4963) <= not(layer0_outputs(675));
    outputs(4964) <= not(layer0_outputs(3952));
    outputs(4965) <= layer0_outputs(3222);
    outputs(4966) <= layer0_outputs(1881);
    outputs(4967) <= not(layer0_outputs(4394));
    outputs(4968) <= layer0_outputs(2646);
    outputs(4969) <= (layer0_outputs(2069)) or (layer0_outputs(1492));
    outputs(4970) <= not((layer0_outputs(537)) xor (layer0_outputs(4996)));
    outputs(4971) <= not(layer0_outputs(1598));
    outputs(4972) <= not((layer0_outputs(509)) or (layer0_outputs(3747)));
    outputs(4973) <= (layer0_outputs(2336)) and not (layer0_outputs(4489));
    outputs(4974) <= (layer0_outputs(2879)) and not (layer0_outputs(937));
    outputs(4975) <= (layer0_outputs(4545)) and not (layer0_outputs(2472));
    outputs(4976) <= not(layer0_outputs(2607));
    outputs(4977) <= (layer0_outputs(296)) and not (layer0_outputs(3447));
    outputs(4978) <= not((layer0_outputs(2437)) and (layer0_outputs(541)));
    outputs(4979) <= not((layer0_outputs(4860)) or (layer0_outputs(3826)));
    outputs(4980) <= (layer0_outputs(893)) and (layer0_outputs(4904));
    outputs(4981) <= not((layer0_outputs(1984)) or (layer0_outputs(856)));
    outputs(4982) <= layer0_outputs(1381);
    outputs(4983) <= (layer0_outputs(3975)) and not (layer0_outputs(4130));
    outputs(4984) <= layer0_outputs(2806);
    outputs(4985) <= (layer0_outputs(2225)) and not (layer0_outputs(1352));
    outputs(4986) <= (layer0_outputs(3835)) and not (layer0_outputs(3054));
    outputs(4987) <= not(layer0_outputs(2477)) or (layer0_outputs(2444));
    outputs(4988) <= not(layer0_outputs(3596)) or (layer0_outputs(5087));
    outputs(4989) <= (layer0_outputs(2206)) and not (layer0_outputs(247));
    outputs(4990) <= layer0_outputs(3518);
    outputs(4991) <= (layer0_outputs(473)) and not (layer0_outputs(1198));
    outputs(4992) <= not((layer0_outputs(2598)) xor (layer0_outputs(594)));
    outputs(4993) <= layer0_outputs(1084);
    outputs(4994) <= not(layer0_outputs(4501));
    outputs(4995) <= not(layer0_outputs(910));
    outputs(4996) <= (layer0_outputs(3556)) and not (layer0_outputs(2275));
    outputs(4997) <= not(layer0_outputs(2933)) or (layer0_outputs(1708));
    outputs(4998) <= (layer0_outputs(725)) and not (layer0_outputs(3199));
    outputs(4999) <= (layer0_outputs(664)) and (layer0_outputs(3058));
    outputs(5000) <= (layer0_outputs(2972)) and (layer0_outputs(3670));
    outputs(5001) <= layer0_outputs(4263);
    outputs(5002) <= not(layer0_outputs(3023));
    outputs(5003) <= not(layer0_outputs(76));
    outputs(5004) <= (layer0_outputs(36)) and (layer0_outputs(4348));
    outputs(5005) <= not(layer0_outputs(367));
    outputs(5006) <= layer0_outputs(1910);
    outputs(5007) <= not(layer0_outputs(4808));
    outputs(5008) <= layer0_outputs(2380);
    outputs(5009) <= (layer0_outputs(4153)) and not (layer0_outputs(4053));
    outputs(5010) <= not((layer0_outputs(4175)) xor (layer0_outputs(216)));
    outputs(5011) <= not((layer0_outputs(1697)) or (layer0_outputs(4597)));
    outputs(5012) <= (layer0_outputs(485)) and not (layer0_outputs(1774));
    outputs(5013) <= not(layer0_outputs(1010));
    outputs(5014) <= (layer0_outputs(3234)) and not (layer0_outputs(3874));
    outputs(5015) <= not(layer0_outputs(5));
    outputs(5016) <= layer0_outputs(3538);
    outputs(5017) <= not(layer0_outputs(4785)) or (layer0_outputs(2095));
    outputs(5018) <= not(layer0_outputs(3435));
    outputs(5019) <= not((layer0_outputs(2368)) xor (layer0_outputs(1842)));
    outputs(5020) <= not(layer0_outputs(1754));
    outputs(5021) <= not((layer0_outputs(3417)) and (layer0_outputs(2832)));
    outputs(5022) <= (layer0_outputs(2317)) and (layer0_outputs(1654));
    outputs(5023) <= not((layer0_outputs(1553)) or (layer0_outputs(3539)));
    outputs(5024) <= layer0_outputs(4599);
    outputs(5025) <= not(layer0_outputs(1551)) or (layer0_outputs(4003));
    outputs(5026) <= layer0_outputs(2208);
    outputs(5027) <= layer0_outputs(984);
    outputs(5028) <= (layer0_outputs(3791)) and not (layer0_outputs(1920));
    outputs(5029) <= (layer0_outputs(1018)) and not (layer0_outputs(3315));
    outputs(5030) <= (layer0_outputs(1675)) and (layer0_outputs(3410));
    outputs(5031) <= (layer0_outputs(3720)) or (layer0_outputs(3664));
    outputs(5032) <= (layer0_outputs(3234)) and not (layer0_outputs(1691));
    outputs(5033) <= (layer0_outputs(626)) and not (layer0_outputs(487));
    outputs(5034) <= not(layer0_outputs(61));
    outputs(5035) <= not(layer0_outputs(1622));
    outputs(5036) <= not(layer0_outputs(1648));
    outputs(5037) <= not(layer0_outputs(3342)) or (layer0_outputs(1712));
    outputs(5038) <= not(layer0_outputs(4511));
    outputs(5039) <= not((layer0_outputs(2875)) or (layer0_outputs(2158)));
    outputs(5040) <= not(layer0_outputs(2126));
    outputs(5041) <= (layer0_outputs(3364)) and (layer0_outputs(2046));
    outputs(5042) <= not((layer0_outputs(4989)) xor (layer0_outputs(4331)));
    outputs(5043) <= layer0_outputs(503);
    outputs(5044) <= not((layer0_outputs(4711)) xor (layer0_outputs(2269)));
    outputs(5045) <= not((layer0_outputs(2256)) xor (layer0_outputs(1160)));
    outputs(5046) <= (layer0_outputs(4755)) and not (layer0_outputs(4055));
    outputs(5047) <= (layer0_outputs(2697)) or (layer0_outputs(2871));
    outputs(5048) <= layer0_outputs(3614);
    outputs(5049) <= (layer0_outputs(797)) and not (layer0_outputs(2391));
    outputs(5050) <= (layer0_outputs(48)) and not (layer0_outputs(2391));
    outputs(5051) <= not((layer0_outputs(3179)) and (layer0_outputs(4676)));
    outputs(5052) <= layer0_outputs(2317);
    outputs(5053) <= layer0_outputs(3795);
    outputs(5054) <= layer0_outputs(2313);
    outputs(5055) <= layer0_outputs(4873);
    outputs(5056) <= layer0_outputs(1671);
    outputs(5057) <= layer0_outputs(3411);
    outputs(5058) <= not(layer0_outputs(2753));
    outputs(5059) <= (layer0_outputs(5114)) and (layer0_outputs(2092));
    outputs(5060) <= (layer0_outputs(2072)) and not (layer0_outputs(3298));
    outputs(5061) <= not(layer0_outputs(1735));
    outputs(5062) <= (layer0_outputs(1361)) and not (layer0_outputs(3712));
    outputs(5063) <= (layer0_outputs(680)) and not (layer0_outputs(4283));
    outputs(5064) <= not((layer0_outputs(4903)) or (layer0_outputs(331)));
    outputs(5065) <= layer0_outputs(4658);
    outputs(5066) <= layer0_outputs(4642);
    outputs(5067) <= (layer0_outputs(3707)) and (layer0_outputs(222));
    outputs(5068) <= not(layer0_outputs(2585));
    outputs(5069) <= layer0_outputs(2034);
    outputs(5070) <= not(layer0_outputs(625));
    outputs(5071) <= (layer0_outputs(5031)) and (layer0_outputs(3891));
    outputs(5072) <= not((layer0_outputs(3408)) or (layer0_outputs(3148)));
    outputs(5073) <= (layer0_outputs(2781)) and not (layer0_outputs(2673));
    outputs(5074) <= not((layer0_outputs(1289)) xor (layer0_outputs(992)));
    outputs(5075) <= not(layer0_outputs(2021));
    outputs(5076) <= not((layer0_outputs(3940)) xor (layer0_outputs(23)));
    outputs(5077) <= not((layer0_outputs(4205)) or (layer0_outputs(1877)));
    outputs(5078) <= (layer0_outputs(328)) and (layer0_outputs(4919));
    outputs(5079) <= layer0_outputs(3520);
    outputs(5080) <= not(layer0_outputs(2832)) or (layer0_outputs(3898));
    outputs(5081) <= (layer0_outputs(4697)) and (layer0_outputs(4643));
    outputs(5082) <= layer0_outputs(2570);
    outputs(5083) <= not(layer0_outputs(3254));
    outputs(5084) <= layer0_outputs(824);
    outputs(5085) <= not((layer0_outputs(3406)) xor (layer0_outputs(2501)));
    outputs(5086) <= layer0_outputs(1868);
    outputs(5087) <= (layer0_outputs(2130)) and (layer0_outputs(464));
    outputs(5088) <= not((layer0_outputs(2961)) or (layer0_outputs(3734)));
    outputs(5089) <= (layer0_outputs(1075)) and not (layer0_outputs(1221));
    outputs(5090) <= (layer0_outputs(4106)) and not (layer0_outputs(190));
    outputs(5091) <= (layer0_outputs(3291)) xor (layer0_outputs(742));
    outputs(5092) <= not(layer0_outputs(3132));
    outputs(5093) <= not(layer0_outputs(3745));
    outputs(5094) <= not(layer0_outputs(2663)) or (layer0_outputs(2680));
    outputs(5095) <= not((layer0_outputs(3248)) or (layer0_outputs(4714)));
    outputs(5096) <= (layer0_outputs(845)) and (layer0_outputs(2859));
    outputs(5097) <= (layer0_outputs(1644)) and not (layer0_outputs(533));
    outputs(5098) <= layer0_outputs(364);
    outputs(5099) <= (layer0_outputs(3942)) and (layer0_outputs(295));
    outputs(5100) <= layer0_outputs(678);
    outputs(5101) <= not((layer0_outputs(4063)) or (layer0_outputs(2249)));
    outputs(5102) <= not(layer0_outputs(1290));
    outputs(5103) <= layer0_outputs(4554);
    outputs(5104) <= layer0_outputs(2187);
    outputs(5105) <= (layer0_outputs(3982)) xor (layer0_outputs(2105));
    outputs(5106) <= not((layer0_outputs(603)) or (layer0_outputs(2556)));
    outputs(5107) <= (layer0_outputs(147)) xor (layer0_outputs(1773));
    outputs(5108) <= (layer0_outputs(127)) xor (layer0_outputs(3002));
    outputs(5109) <= not(layer0_outputs(441));
    outputs(5110) <= (layer0_outputs(1182)) and not (layer0_outputs(269));
    outputs(5111) <= (layer0_outputs(1292)) and not (layer0_outputs(1249));
    outputs(5112) <= not(layer0_outputs(2752));
    outputs(5113) <= (layer0_outputs(942)) and not (layer0_outputs(2774));
    outputs(5114) <= (layer0_outputs(1434)) and not (layer0_outputs(1336));
    outputs(5115) <= (layer0_outputs(1349)) or (layer0_outputs(4161));
    outputs(5116) <= (layer0_outputs(365)) and not (layer0_outputs(4887));
    outputs(5117) <= (layer0_outputs(2903)) and (layer0_outputs(3950));
    outputs(5118) <= not((layer0_outputs(2600)) or (layer0_outputs(4455)));
    outputs(5119) <= not(layer0_outputs(4007)) or (layer0_outputs(3441));

end Behavioral;
