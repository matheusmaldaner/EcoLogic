library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs: in std_logic_vector(1023 downto 0);
        outputs: out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs: std_logic_vector(10239 downto 0);
    signal layer1_outputs: std_logic_vector(10239 downto 0);
    signal layer2_outputs: std_logic_vector(10239 downto 0);

begin
    layer0_outputs(0) <= a or b;
    layer0_outputs(1) <= b;
    layer0_outputs(2) <= not b;
    layer0_outputs(3) <= a or b;
    layer0_outputs(4) <= not b;
    layer0_outputs(5) <= not (a or b);
    layer0_outputs(6) <= not a or b;
    layer0_outputs(7) <= a or b;
    layer0_outputs(8) <= not a;
    layer0_outputs(9) <= a and not b;
    layer0_outputs(10) <= not (a and b);
    layer0_outputs(11) <= not a;
    layer0_outputs(12) <= a and b;
    layer0_outputs(13) <= b;
    layer0_outputs(14) <= a or b;
    layer0_outputs(15) <= not a;
    layer0_outputs(16) <= a and not b;
    layer0_outputs(17) <= b and not a;
    layer0_outputs(18) <= '1';
    layer0_outputs(19) <= not (a or b);
    layer0_outputs(20) <= not a or b;
    layer0_outputs(21) <= a and not b;
    layer0_outputs(22) <= not (a xor b);
    layer0_outputs(23) <= b;
    layer0_outputs(24) <= not (a and b);
    layer0_outputs(25) <= a or b;
    layer0_outputs(26) <= not (a or b);
    layer0_outputs(27) <= not (a or b);
    layer0_outputs(28) <= a;
    layer0_outputs(29) <= a or b;
    layer0_outputs(30) <= a and not b;
    layer0_outputs(31) <= '0';
    layer0_outputs(32) <= b;
    layer0_outputs(33) <= a or b;
    layer0_outputs(34) <= not b or a;
    layer0_outputs(35) <= not b;
    layer0_outputs(36) <= not (a xor b);
    layer0_outputs(37) <= a or b;
    layer0_outputs(38) <= not b or a;
    layer0_outputs(39) <= not (a or b);
    layer0_outputs(40) <= not b;
    layer0_outputs(41) <= a or b;
    layer0_outputs(42) <= b and not a;
    layer0_outputs(43) <= '0';
    layer0_outputs(44) <= not (a or b);
    layer0_outputs(45) <= not b;
    layer0_outputs(46) <= not (a xor b);
    layer0_outputs(47) <= not (a xor b);
    layer0_outputs(48) <= '0';
    layer0_outputs(49) <= a xor b;
    layer0_outputs(50) <= a or b;
    layer0_outputs(51) <= not b;
    layer0_outputs(52) <= a xor b;
    layer0_outputs(53) <= b and not a;
    layer0_outputs(54) <= b and not a;
    layer0_outputs(55) <= not (a or b);
    layer0_outputs(56) <= a;
    layer0_outputs(57) <= '1';
    layer0_outputs(58) <= b and not a;
    layer0_outputs(59) <= a;
    layer0_outputs(60) <= not b or a;
    layer0_outputs(61) <= not (a or b);
    layer0_outputs(62) <= a;
    layer0_outputs(63) <= a or b;
    layer0_outputs(64) <= a;
    layer0_outputs(65) <= not (a and b);
    layer0_outputs(66) <= a or b;
    layer0_outputs(67) <= a or b;
    layer0_outputs(68) <= a;
    layer0_outputs(69) <= b and not a;
    layer0_outputs(70) <= a and b;
    layer0_outputs(71) <= a xor b;
    layer0_outputs(72) <= not a;
    layer0_outputs(73) <= b and not a;
    layer0_outputs(74) <= a and not b;
    layer0_outputs(75) <= b and not a;
    layer0_outputs(76) <= a xor b;
    layer0_outputs(77) <= a and not b;
    layer0_outputs(78) <= a or b;
    layer0_outputs(79) <= a or b;
    layer0_outputs(80) <= b and not a;
    layer0_outputs(81) <= a or b;
    layer0_outputs(82) <= a and b;
    layer0_outputs(83) <= not (a xor b);
    layer0_outputs(84) <= not (a xor b);
    layer0_outputs(85) <= not (a xor b);
    layer0_outputs(86) <= a or b;
    layer0_outputs(87) <= b;
    layer0_outputs(88) <= a;
    layer0_outputs(89) <= not (a xor b);
    layer0_outputs(90) <= not a;
    layer0_outputs(91) <= a xor b;
    layer0_outputs(92) <= not a;
    layer0_outputs(93) <= not a or b;
    layer0_outputs(94) <= b;
    layer0_outputs(95) <= a and not b;
    layer0_outputs(96) <= not a;
    layer0_outputs(97) <= not (a and b);
    layer0_outputs(98) <= a and not b;
    layer0_outputs(99) <= not (a xor b);
    layer0_outputs(100) <= not (a xor b);
    layer0_outputs(101) <= a xor b;
    layer0_outputs(102) <= a or b;
    layer0_outputs(103) <= b and not a;
    layer0_outputs(104) <= not (a and b);
    layer0_outputs(105) <= b;
    layer0_outputs(106) <= not a;
    layer0_outputs(107) <= a and not b;
    layer0_outputs(108) <= not b or a;
    layer0_outputs(109) <= not (a or b);
    layer0_outputs(110) <= a xor b;
    layer0_outputs(111) <= b;
    layer0_outputs(112) <= not b or a;
    layer0_outputs(113) <= not b or a;
    layer0_outputs(114) <= a xor b;
    layer0_outputs(115) <= not b;
    layer0_outputs(116) <= a or b;
    layer0_outputs(117) <= a;
    layer0_outputs(118) <= b and not a;
    layer0_outputs(119) <= a and not b;
    layer0_outputs(120) <= not a;
    layer0_outputs(121) <= not b or a;
    layer0_outputs(122) <= '0';
    layer0_outputs(123) <= '1';
    layer0_outputs(124) <= '0';
    layer0_outputs(125) <= not (a or b);
    layer0_outputs(126) <= a or b;
    layer0_outputs(127) <= not b;
    layer0_outputs(128) <= a or b;
    layer0_outputs(129) <= a;
    layer0_outputs(130) <= not b or a;
    layer0_outputs(131) <= not (a or b);
    layer0_outputs(132) <= a and not b;
    layer0_outputs(133) <= not (a or b);
    layer0_outputs(134) <= a or b;
    layer0_outputs(135) <= not (a or b);
    layer0_outputs(136) <= '1';
    layer0_outputs(137) <= a or b;
    layer0_outputs(138) <= '1';
    layer0_outputs(139) <= a xor b;
    layer0_outputs(140) <= a;
    layer0_outputs(141) <= not b or a;
    layer0_outputs(142) <= b and not a;
    layer0_outputs(143) <= '1';
    layer0_outputs(144) <= not (a or b);
    layer0_outputs(145) <= not a;
    layer0_outputs(146) <= a and not b;
    layer0_outputs(147) <= not (a and b);
    layer0_outputs(148) <= not b or a;
    layer0_outputs(149) <= not b;
    layer0_outputs(150) <= not (a or b);
    layer0_outputs(151) <= b and not a;
    layer0_outputs(152) <= not a;
    layer0_outputs(153) <= not a or b;
    layer0_outputs(154) <= not (a or b);
    layer0_outputs(155) <= a xor b;
    layer0_outputs(156) <= a or b;
    layer0_outputs(157) <= not a or b;
    layer0_outputs(158) <= a xor b;
    layer0_outputs(159) <= b;
    layer0_outputs(160) <= not b or a;
    layer0_outputs(161) <= not a or b;
    layer0_outputs(162) <= a and not b;
    layer0_outputs(163) <= not (a xor b);
    layer0_outputs(164) <= not a or b;
    layer0_outputs(165) <= not b;
    layer0_outputs(166) <= a and b;
    layer0_outputs(167) <= b and not a;
    layer0_outputs(168) <= not b;
    layer0_outputs(169) <= not (a xor b);
    layer0_outputs(170) <= '1';
    layer0_outputs(171) <= a xor b;
    layer0_outputs(172) <= b and not a;
    layer0_outputs(173) <= not (a xor b);
    layer0_outputs(174) <= a xor b;
    layer0_outputs(175) <= a and not b;
    layer0_outputs(176) <= not b;
    layer0_outputs(177) <= a xor b;
    layer0_outputs(178) <= not a;
    layer0_outputs(179) <= b;
    layer0_outputs(180) <= not a;
    layer0_outputs(181) <= not (a xor b);
    layer0_outputs(182) <= not a;
    layer0_outputs(183) <= a;
    layer0_outputs(184) <= '1';
    layer0_outputs(185) <= not a or b;
    layer0_outputs(186) <= not (a xor b);
    layer0_outputs(187) <= a;
    layer0_outputs(188) <= a or b;
    layer0_outputs(189) <= not b;
    layer0_outputs(190) <= a or b;
    layer0_outputs(191) <= a and b;
    layer0_outputs(192) <= a xor b;
    layer0_outputs(193) <= b;
    layer0_outputs(194) <= b;
    layer0_outputs(195) <= not a or b;
    layer0_outputs(196) <= b;
    layer0_outputs(197) <= a;
    layer0_outputs(198) <= a or b;
    layer0_outputs(199) <= a and not b;
    layer0_outputs(200) <= a xor b;
    layer0_outputs(201) <= a;
    layer0_outputs(202) <= b;
    layer0_outputs(203) <= a and not b;
    layer0_outputs(204) <= not (a or b);
    layer0_outputs(205) <= b;
    layer0_outputs(206) <= not (a xor b);
    layer0_outputs(207) <= a or b;
    layer0_outputs(208) <= not (a or b);
    layer0_outputs(209) <= a or b;
    layer0_outputs(210) <= a or b;
    layer0_outputs(211) <= not b or a;
    layer0_outputs(212) <= a xor b;
    layer0_outputs(213) <= b;
    layer0_outputs(214) <= not b;
    layer0_outputs(215) <= not b;
    layer0_outputs(216) <= not (a or b);
    layer0_outputs(217) <= not (a or b);
    layer0_outputs(218) <= not (a xor b);
    layer0_outputs(219) <= a and not b;
    layer0_outputs(220) <= a;
    layer0_outputs(221) <= not a;
    layer0_outputs(222) <= not b or a;
    layer0_outputs(223) <= not a or b;
    layer0_outputs(224) <= '1';
    layer0_outputs(225) <= a xor b;
    layer0_outputs(226) <= not (a xor b);
    layer0_outputs(227) <= not a;
    layer0_outputs(228) <= b;
    layer0_outputs(229) <= a xor b;
    layer0_outputs(230) <= a and b;
    layer0_outputs(231) <= a and b;
    layer0_outputs(232) <= b and not a;
    layer0_outputs(233) <= a;
    layer0_outputs(234) <= a and not b;
    layer0_outputs(235) <= not (a xor b);
    layer0_outputs(236) <= not b or a;
    layer0_outputs(237) <= a;
    layer0_outputs(238) <= not b or a;
    layer0_outputs(239) <= not (a or b);
    layer0_outputs(240) <= '1';
    layer0_outputs(241) <= not (a xor b);
    layer0_outputs(242) <= not a;
    layer0_outputs(243) <= not b;
    layer0_outputs(244) <= not (a and b);
    layer0_outputs(245) <= not a;
    layer0_outputs(246) <= '1';
    layer0_outputs(247) <= not (a or b);
    layer0_outputs(248) <= '0';
    layer0_outputs(249) <= not (a xor b);
    layer0_outputs(250) <= not a;
    layer0_outputs(251) <= not a;
    layer0_outputs(252) <= not (a or b);
    layer0_outputs(253) <= not (a or b);
    layer0_outputs(254) <= not (a or b);
    layer0_outputs(255) <= not a or b;
    layer0_outputs(256) <= a;
    layer0_outputs(257) <= not a;
    layer0_outputs(258) <= not (a or b);
    layer0_outputs(259) <= not a;
    layer0_outputs(260) <= b;
    layer0_outputs(261) <= not (a or b);
    layer0_outputs(262) <= not (a and b);
    layer0_outputs(263) <= a or b;
    layer0_outputs(264) <= not (a or b);
    layer0_outputs(265) <= a;
    layer0_outputs(266) <= b;
    layer0_outputs(267) <= a xor b;
    layer0_outputs(268) <= a xor b;
    layer0_outputs(269) <= a xor b;
    layer0_outputs(270) <= not b;
    layer0_outputs(271) <= a;
    layer0_outputs(272) <= not a or b;
    layer0_outputs(273) <= not a;
    layer0_outputs(274) <= not a;
    layer0_outputs(275) <= not b;
    layer0_outputs(276) <= not (a xor b);
    layer0_outputs(277) <= not a;
    layer0_outputs(278) <= a or b;
    layer0_outputs(279) <= not b or a;
    layer0_outputs(280) <= a or b;
    layer0_outputs(281) <= a and not b;
    layer0_outputs(282) <= not (a or b);
    layer0_outputs(283) <= b;
    layer0_outputs(284) <= not a;
    layer0_outputs(285) <= not (a xor b);
    layer0_outputs(286) <= b and not a;
    layer0_outputs(287) <= not (a or b);
    layer0_outputs(288) <= not a;
    layer0_outputs(289) <= b;
    layer0_outputs(290) <= not a or b;
    layer0_outputs(291) <= not b or a;
    layer0_outputs(292) <= not b or a;
    layer0_outputs(293) <= b;
    layer0_outputs(294) <= not (a or b);
    layer0_outputs(295) <= '0';
    layer0_outputs(296) <= '1';
    layer0_outputs(297) <= a;
    layer0_outputs(298) <= not (a or b);
    layer0_outputs(299) <= not a;
    layer0_outputs(300) <= b;
    layer0_outputs(301) <= a or b;
    layer0_outputs(302) <= not (a xor b);
    layer0_outputs(303) <= a or b;
    layer0_outputs(304) <= b and not a;
    layer0_outputs(305) <= a or b;
    layer0_outputs(306) <= a and not b;
    layer0_outputs(307) <= not a;
    layer0_outputs(308) <= b and not a;
    layer0_outputs(309) <= not (a or b);
    layer0_outputs(310) <= not (a or b);
    layer0_outputs(311) <= not a or b;
    layer0_outputs(312) <= not a or b;
    layer0_outputs(313) <= a xor b;
    layer0_outputs(314) <= not a;
    layer0_outputs(315) <= a xor b;
    layer0_outputs(316) <= not (a xor b);
    layer0_outputs(317) <= a or b;
    layer0_outputs(318) <= '1';
    layer0_outputs(319) <= a;
    layer0_outputs(320) <= '1';
    layer0_outputs(321) <= not (a xor b);
    layer0_outputs(322) <= not (a or b);
    layer0_outputs(323) <= a and not b;
    layer0_outputs(324) <= not b;
    layer0_outputs(325) <= a or b;
    layer0_outputs(326) <= not (a or b);
    layer0_outputs(327) <= a and not b;
    layer0_outputs(328) <= not (a or b);
    layer0_outputs(329) <= not a or b;
    layer0_outputs(330) <= not a;
    layer0_outputs(331) <= a and not b;
    layer0_outputs(332) <= a or b;
    layer0_outputs(333) <= a xor b;
    layer0_outputs(334) <= a xor b;
    layer0_outputs(335) <= a and not b;
    layer0_outputs(336) <= not b;
    layer0_outputs(337) <= not (a xor b);
    layer0_outputs(338) <= a or b;
    layer0_outputs(339) <= a;
    layer0_outputs(340) <= a or b;
    layer0_outputs(341) <= '0';
    layer0_outputs(342) <= not (a xor b);
    layer0_outputs(343) <= a xor b;
    layer0_outputs(344) <= not (a and b);
    layer0_outputs(345) <= not a or b;
    layer0_outputs(346) <= a or b;
    layer0_outputs(347) <= not (a xor b);
    layer0_outputs(348) <= not (a or b);
    layer0_outputs(349) <= b;
    layer0_outputs(350) <= not (a and b);
    layer0_outputs(351) <= a xor b;
    layer0_outputs(352) <= a or b;
    layer0_outputs(353) <= b;
    layer0_outputs(354) <= not b or a;
    layer0_outputs(355) <= not (a or b);
    layer0_outputs(356) <= b and not a;
    layer0_outputs(357) <= b;
    layer0_outputs(358) <= not b or a;
    layer0_outputs(359) <= not (a xor b);
    layer0_outputs(360) <= a or b;
    layer0_outputs(361) <= not (a or b);
    layer0_outputs(362) <= not a;
    layer0_outputs(363) <= '1';
    layer0_outputs(364) <= a xor b;
    layer0_outputs(365) <= not (a or b);
    layer0_outputs(366) <= not (a or b);
    layer0_outputs(367) <= not b or a;
    layer0_outputs(368) <= not (a or b);
    layer0_outputs(369) <= not (a xor b);
    layer0_outputs(370) <= a;
    layer0_outputs(371) <= not (a and b);
    layer0_outputs(372) <= not (a or b);
    layer0_outputs(373) <= not (a xor b);
    layer0_outputs(374) <= not a;
    layer0_outputs(375) <= not a;
    layer0_outputs(376) <= not (a or b);
    layer0_outputs(377) <= a or b;
    layer0_outputs(378) <= not (a or b);
    layer0_outputs(379) <= not (a or b);
    layer0_outputs(380) <= not b;
    layer0_outputs(381) <= not (a xor b);
    layer0_outputs(382) <= a and not b;
    layer0_outputs(383) <= a;
    layer0_outputs(384) <= not (a xor b);
    layer0_outputs(385) <= a xor b;
    layer0_outputs(386) <= not b;
    layer0_outputs(387) <= a or b;
    layer0_outputs(388) <= a or b;
    layer0_outputs(389) <= not a;
    layer0_outputs(390) <= not b or a;
    layer0_outputs(391) <= not (a xor b);
    layer0_outputs(392) <= a;
    layer0_outputs(393) <= not b;
    layer0_outputs(394) <= not b or a;
    layer0_outputs(395) <= not (a and b);
    layer0_outputs(396) <= b;
    layer0_outputs(397) <= not (a or b);
    layer0_outputs(398) <= a;
    layer0_outputs(399) <= a;
    layer0_outputs(400) <= a xor b;
    layer0_outputs(401) <= not (a and b);
    layer0_outputs(402) <= b;
    layer0_outputs(403) <= not (a xor b);
    layer0_outputs(404) <= not (a xor b);
    layer0_outputs(405) <= not a or b;
    layer0_outputs(406) <= a and not b;
    layer0_outputs(407) <= not a or b;
    layer0_outputs(408) <= b;
    layer0_outputs(409) <= a and not b;
    layer0_outputs(410) <= a and not b;
    layer0_outputs(411) <= a;
    layer0_outputs(412) <= '0';
    layer0_outputs(413) <= not (a xor b);
    layer0_outputs(414) <= not (a or b);
    layer0_outputs(415) <= a and not b;
    layer0_outputs(416) <= a xor b;
    layer0_outputs(417) <= '1';
    layer0_outputs(418) <= a or b;
    layer0_outputs(419) <= not b;
    layer0_outputs(420) <= not a or b;
    layer0_outputs(421) <= not b or a;
    layer0_outputs(422) <= a or b;
    layer0_outputs(423) <= not (a xor b);
    layer0_outputs(424) <= not a or b;
    layer0_outputs(425) <= not b or a;
    layer0_outputs(426) <= not (a xor b);
    layer0_outputs(427) <= not (a xor b);
    layer0_outputs(428) <= a;
    layer0_outputs(429) <= b and not a;
    layer0_outputs(430) <= a and not b;
    layer0_outputs(431) <= not (a or b);
    layer0_outputs(432) <= a xor b;
    layer0_outputs(433) <= a and b;
    layer0_outputs(434) <= not b or a;
    layer0_outputs(435) <= a or b;
    layer0_outputs(436) <= a;
    layer0_outputs(437) <= a;
    layer0_outputs(438) <= a and not b;
    layer0_outputs(439) <= not b;
    layer0_outputs(440) <= '1';
    layer0_outputs(441) <= a;
    layer0_outputs(442) <= b;
    layer0_outputs(443) <= a and not b;
    layer0_outputs(444) <= a or b;
    layer0_outputs(445) <= a and not b;
    layer0_outputs(446) <= not b;
    layer0_outputs(447) <= b and not a;
    layer0_outputs(448) <= a xor b;
    layer0_outputs(449) <= not (a or b);
    layer0_outputs(450) <= b and not a;
    layer0_outputs(451) <= not b;
    layer0_outputs(452) <= b;
    layer0_outputs(453) <= not a or b;
    layer0_outputs(454) <= b and not a;
    layer0_outputs(455) <= b and not a;
    layer0_outputs(456) <= not (a or b);
    layer0_outputs(457) <= a or b;
    layer0_outputs(458) <= a;
    layer0_outputs(459) <= not b;
    layer0_outputs(460) <= '0';
    layer0_outputs(461) <= not (a or b);
    layer0_outputs(462) <= b;
    layer0_outputs(463) <= a xor b;
    layer0_outputs(464) <= a or b;
    layer0_outputs(465) <= not a or b;
    layer0_outputs(466) <= b;
    layer0_outputs(467) <= not (a and b);
    layer0_outputs(468) <= b;
    layer0_outputs(469) <= not (a or b);
    layer0_outputs(470) <= not (a or b);
    layer0_outputs(471) <= b and not a;
    layer0_outputs(472) <= a;
    layer0_outputs(473) <= not a;
    layer0_outputs(474) <= not (a and b);
    layer0_outputs(475) <= a and not b;
    layer0_outputs(476) <= a and not b;
    layer0_outputs(477) <= b and not a;
    layer0_outputs(478) <= a xor b;
    layer0_outputs(479) <= not b or a;
    layer0_outputs(480) <= a and not b;
    layer0_outputs(481) <= not (a or b);
    layer0_outputs(482) <= not (a xor b);
    layer0_outputs(483) <= a or b;
    layer0_outputs(484) <= a and not b;
    layer0_outputs(485) <= a xor b;
    layer0_outputs(486) <= b;
    layer0_outputs(487) <= a or b;
    layer0_outputs(488) <= not (a and b);
    layer0_outputs(489) <= a and not b;
    layer0_outputs(490) <= a xor b;
    layer0_outputs(491) <= a or b;
    layer0_outputs(492) <= not (a xor b);
    layer0_outputs(493) <= not (a xor b);
    layer0_outputs(494) <= '1';
    layer0_outputs(495) <= '1';
    layer0_outputs(496) <= a xor b;
    layer0_outputs(497) <= not (a or b);
    layer0_outputs(498) <= not a or b;
    layer0_outputs(499) <= a;
    layer0_outputs(500) <= not b;
    layer0_outputs(501) <= not b;
    layer0_outputs(502) <= a or b;
    layer0_outputs(503) <= '0';
    layer0_outputs(504) <= not b;
    layer0_outputs(505) <= a xor b;
    layer0_outputs(506) <= not (a or b);
    layer0_outputs(507) <= b;
    layer0_outputs(508) <= a;
    layer0_outputs(509) <= a;
    layer0_outputs(510) <= not b or a;
    layer0_outputs(511) <= a and not b;
    layer0_outputs(512) <= not b or a;
    layer0_outputs(513) <= b and not a;
    layer0_outputs(514) <= not a;
    layer0_outputs(515) <= a or b;
    layer0_outputs(516) <= b;
    layer0_outputs(517) <= a;
    layer0_outputs(518) <= b;
    layer0_outputs(519) <= not (a xor b);
    layer0_outputs(520) <= a xor b;
    layer0_outputs(521) <= a and not b;
    layer0_outputs(522) <= not a;
    layer0_outputs(523) <= a;
    layer0_outputs(524) <= a and not b;
    layer0_outputs(525) <= not b or a;
    layer0_outputs(526) <= not a or b;
    layer0_outputs(527) <= not (a or b);
    layer0_outputs(528) <= not b;
    layer0_outputs(529) <= not (a or b);
    layer0_outputs(530) <= a or b;
    layer0_outputs(531) <= b;
    layer0_outputs(532) <= not (a or b);
    layer0_outputs(533) <= not a or b;
    layer0_outputs(534) <= b and not a;
    layer0_outputs(535) <= '1';
    layer0_outputs(536) <= not a;
    layer0_outputs(537) <= not a or b;
    layer0_outputs(538) <= b;
    layer0_outputs(539) <= b and not a;
    layer0_outputs(540) <= not b or a;
    layer0_outputs(541) <= not (a and b);
    layer0_outputs(542) <= not a;
    layer0_outputs(543) <= a or b;
    layer0_outputs(544) <= not b or a;
    layer0_outputs(545) <= a xor b;
    layer0_outputs(546) <= b and not a;
    layer0_outputs(547) <= a or b;
    layer0_outputs(548) <= a or b;
    layer0_outputs(549) <= a and not b;
    layer0_outputs(550) <= a and b;
    layer0_outputs(551) <= a xor b;
    layer0_outputs(552) <= '0';
    layer0_outputs(553) <= not a or b;
    layer0_outputs(554) <= a xor b;
    layer0_outputs(555) <= b;
    layer0_outputs(556) <= not a;
    layer0_outputs(557) <= not (a or b);
    layer0_outputs(558) <= not (a and b);
    layer0_outputs(559) <= '0';
    layer0_outputs(560) <= b;
    layer0_outputs(561) <= a or b;
    layer0_outputs(562) <= not b;
    layer0_outputs(563) <= b and not a;
    layer0_outputs(564) <= a or b;
    layer0_outputs(565) <= a xor b;
    layer0_outputs(566) <= b;
    layer0_outputs(567) <= not (a or b);
    layer0_outputs(568) <= not (a or b);
    layer0_outputs(569) <= not a or b;
    layer0_outputs(570) <= b;
    layer0_outputs(571) <= b and not a;
    layer0_outputs(572) <= a;
    layer0_outputs(573) <= not (a or b);
    layer0_outputs(574) <= not a or b;
    layer0_outputs(575) <= not b;
    layer0_outputs(576) <= a and not b;
    layer0_outputs(577) <= '0';
    layer0_outputs(578) <= not a;
    layer0_outputs(579) <= b;
    layer0_outputs(580) <= not (a xor b);
    layer0_outputs(581) <= not (a xor b);
    layer0_outputs(582) <= not (a or b);
    layer0_outputs(583) <= not (a or b);
    layer0_outputs(584) <= not a or b;
    layer0_outputs(585) <= '0';
    layer0_outputs(586) <= a and not b;
    layer0_outputs(587) <= a or b;
    layer0_outputs(588) <= not (a or b);
    layer0_outputs(589) <= not (a or b);
    layer0_outputs(590) <= a;
    layer0_outputs(591) <= not (a or b);
    layer0_outputs(592) <= a or b;
    layer0_outputs(593) <= not a;
    layer0_outputs(594) <= not (a xor b);
    layer0_outputs(595) <= not (a xor b);
    layer0_outputs(596) <= b and not a;
    layer0_outputs(597) <= not (a xor b);
    layer0_outputs(598) <= not a or b;
    layer0_outputs(599) <= not (a and b);
    layer0_outputs(600) <= '0';
    layer0_outputs(601) <= not (a and b);
    layer0_outputs(602) <= not (a or b);
    layer0_outputs(603) <= not (a or b);
    layer0_outputs(604) <= a or b;
    layer0_outputs(605) <= a or b;
    layer0_outputs(606) <= a or b;
    layer0_outputs(607) <= b;
    layer0_outputs(608) <= a xor b;
    layer0_outputs(609) <= a and b;
    layer0_outputs(610) <= '0';
    layer0_outputs(611) <= a;
    layer0_outputs(612) <= '1';
    layer0_outputs(613) <= not a or b;
    layer0_outputs(614) <= not (a xor b);
    layer0_outputs(615) <= not (a xor b);
    layer0_outputs(616) <= a or b;
    layer0_outputs(617) <= not (a or b);
    layer0_outputs(618) <= a or b;
    layer0_outputs(619) <= not (a xor b);
    layer0_outputs(620) <= a and b;
    layer0_outputs(621) <= a and not b;
    layer0_outputs(622) <= not b;
    layer0_outputs(623) <= not a;
    layer0_outputs(624) <= a and not b;
    layer0_outputs(625) <= a and not b;
    layer0_outputs(626) <= b and not a;
    layer0_outputs(627) <= not (a or b);
    layer0_outputs(628) <= not (a or b);
    layer0_outputs(629) <= a and b;
    layer0_outputs(630) <= not (a or b);
    layer0_outputs(631) <= not a;
    layer0_outputs(632) <= a;
    layer0_outputs(633) <= a xor b;
    layer0_outputs(634) <= b;
    layer0_outputs(635) <= not (a or b);
    layer0_outputs(636) <= not (a or b);
    layer0_outputs(637) <= a and not b;
    layer0_outputs(638) <= a and not b;
    layer0_outputs(639) <= a xor b;
    layer0_outputs(640) <= not (a or b);
    layer0_outputs(641) <= not b;
    layer0_outputs(642) <= a or b;
    layer0_outputs(643) <= a and b;
    layer0_outputs(644) <= a and not b;
    layer0_outputs(645) <= b and not a;
    layer0_outputs(646) <= b;
    layer0_outputs(647) <= not b or a;
    layer0_outputs(648) <= a or b;
    layer0_outputs(649) <= b and not a;
    layer0_outputs(650) <= not a or b;
    layer0_outputs(651) <= a xor b;
    layer0_outputs(652) <= not (a or b);
    layer0_outputs(653) <= not (a or b);
    layer0_outputs(654) <= not a or b;
    layer0_outputs(655) <= a xor b;
    layer0_outputs(656) <= not (a xor b);
    layer0_outputs(657) <= a;
    layer0_outputs(658) <= a;
    layer0_outputs(659) <= not a or b;
    layer0_outputs(660) <= b;
    layer0_outputs(661) <= b and not a;
    layer0_outputs(662) <= a or b;
    layer0_outputs(663) <= not a;
    layer0_outputs(664) <= not b or a;
    layer0_outputs(665) <= not (a xor b);
    layer0_outputs(666) <= a or b;
    layer0_outputs(667) <= not b;
    layer0_outputs(668) <= not a or b;
    layer0_outputs(669) <= not (a or b);
    layer0_outputs(670) <= b;
    layer0_outputs(671) <= not a;
    layer0_outputs(672) <= not b;
    layer0_outputs(673) <= not a;
    layer0_outputs(674) <= a or b;
    layer0_outputs(675) <= not b or a;
    layer0_outputs(676) <= not b;
    layer0_outputs(677) <= not (a or b);
    layer0_outputs(678) <= not a or b;
    layer0_outputs(679) <= a and not b;
    layer0_outputs(680) <= b;
    layer0_outputs(681) <= not (a or b);
    layer0_outputs(682) <= a xor b;
    layer0_outputs(683) <= a or b;
    layer0_outputs(684) <= not b;
    layer0_outputs(685) <= a and not b;
    layer0_outputs(686) <= not a;
    layer0_outputs(687) <= not (a xor b);
    layer0_outputs(688) <= b;
    layer0_outputs(689) <= not (a or b);
    layer0_outputs(690) <= a xor b;
    layer0_outputs(691) <= not (a xor b);
    layer0_outputs(692) <= a;
    layer0_outputs(693) <= a xor b;
    layer0_outputs(694) <= not (a or b);
    layer0_outputs(695) <= not b;
    layer0_outputs(696) <= not (a xor b);
    layer0_outputs(697) <= a xor b;
    layer0_outputs(698) <= not (a xor b);
    layer0_outputs(699) <= not (a or b);
    layer0_outputs(700) <= b and not a;
    layer0_outputs(701) <= a and b;
    layer0_outputs(702) <= not b;
    layer0_outputs(703) <= not a or b;
    layer0_outputs(704) <= not b or a;
    layer0_outputs(705) <= not (a xor b);
    layer0_outputs(706) <= a and not b;
    layer0_outputs(707) <= a or b;
    layer0_outputs(708) <= a xor b;
    layer0_outputs(709) <= not a or b;
    layer0_outputs(710) <= b;
    layer0_outputs(711) <= not (a xor b);
    layer0_outputs(712) <= not b or a;
    layer0_outputs(713) <= not a;
    layer0_outputs(714) <= a xor b;
    layer0_outputs(715) <= not a;
    layer0_outputs(716) <= '1';
    layer0_outputs(717) <= '1';
    layer0_outputs(718) <= b;
    layer0_outputs(719) <= a and not b;
    layer0_outputs(720) <= '1';
    layer0_outputs(721) <= '1';
    layer0_outputs(722) <= a xor b;
    layer0_outputs(723) <= '0';
    layer0_outputs(724) <= not (a xor b);
    layer0_outputs(725) <= not a;
    layer0_outputs(726) <= not (a or b);
    layer0_outputs(727) <= not b or a;
    layer0_outputs(728) <= b and not a;
    layer0_outputs(729) <= not a;
    layer0_outputs(730) <= not (a xor b);
    layer0_outputs(731) <= a xor b;
    layer0_outputs(732) <= a xor b;
    layer0_outputs(733) <= a or b;
    layer0_outputs(734) <= '1';
    layer0_outputs(735) <= a and b;
    layer0_outputs(736) <= not b;
    layer0_outputs(737) <= b and not a;
    layer0_outputs(738) <= '1';
    layer0_outputs(739) <= b;
    layer0_outputs(740) <= a xor b;
    layer0_outputs(741) <= not b;
    layer0_outputs(742) <= b and not a;
    layer0_outputs(743) <= a or b;
    layer0_outputs(744) <= not (a or b);
    layer0_outputs(745) <= a;
    layer0_outputs(746) <= not (a or b);
    layer0_outputs(747) <= not b;
    layer0_outputs(748) <= not b;
    layer0_outputs(749) <= '0';
    layer0_outputs(750) <= a or b;
    layer0_outputs(751) <= b;
    layer0_outputs(752) <= not (a or b);
    layer0_outputs(753) <= a;
    layer0_outputs(754) <= '0';
    layer0_outputs(755) <= a or b;
    layer0_outputs(756) <= a and not b;
    layer0_outputs(757) <= not (a xor b);
    layer0_outputs(758) <= not a;
    layer0_outputs(759) <= not b;
    layer0_outputs(760) <= '0';
    layer0_outputs(761) <= a;
    layer0_outputs(762) <= not (a xor b);
    layer0_outputs(763) <= a;
    layer0_outputs(764) <= a xor b;
    layer0_outputs(765) <= not (a xor b);
    layer0_outputs(766) <= a or b;
    layer0_outputs(767) <= a or b;
    layer0_outputs(768) <= not (a and b);
    layer0_outputs(769) <= not (a or b);
    layer0_outputs(770) <= a xor b;
    layer0_outputs(771) <= b and not a;
    layer0_outputs(772) <= a or b;
    layer0_outputs(773) <= b and not a;
    layer0_outputs(774) <= a or b;
    layer0_outputs(775) <= b;
    layer0_outputs(776) <= not b;
    layer0_outputs(777) <= a or b;
    layer0_outputs(778) <= not b;
    layer0_outputs(779) <= not a or b;
    layer0_outputs(780) <= a or b;
    layer0_outputs(781) <= not a;
    layer0_outputs(782) <= a and b;
    layer0_outputs(783) <= a xor b;
    layer0_outputs(784) <= not (a or b);
    layer0_outputs(785) <= a or b;
    layer0_outputs(786) <= b and not a;
    layer0_outputs(787) <= not (a or b);
    layer0_outputs(788) <= not a or b;
    layer0_outputs(789) <= a xor b;
    layer0_outputs(790) <= not (a xor b);
    layer0_outputs(791) <= b and not a;
    layer0_outputs(792) <= a and not b;
    layer0_outputs(793) <= '0';
    layer0_outputs(794) <= not b;
    layer0_outputs(795) <= not (a or b);
    layer0_outputs(796) <= a and b;
    layer0_outputs(797) <= a xor b;
    layer0_outputs(798) <= not (a or b);
    layer0_outputs(799) <= a and not b;
    layer0_outputs(800) <= b;
    layer0_outputs(801) <= a or b;
    layer0_outputs(802) <= not a or b;
    layer0_outputs(803) <= not b;
    layer0_outputs(804) <= a;
    layer0_outputs(805) <= a xor b;
    layer0_outputs(806) <= not b;
    layer0_outputs(807) <= a xor b;
    layer0_outputs(808) <= not b;
    layer0_outputs(809) <= a;
    layer0_outputs(810) <= b;
    layer0_outputs(811) <= not b or a;
    layer0_outputs(812) <= a xor b;
    layer0_outputs(813) <= not b or a;
    layer0_outputs(814) <= not (a or b);
    layer0_outputs(815) <= not (a xor b);
    layer0_outputs(816) <= a or b;
    layer0_outputs(817) <= a or b;
    layer0_outputs(818) <= not b or a;
    layer0_outputs(819) <= '0';
    layer0_outputs(820) <= a and not b;
    layer0_outputs(821) <= not a or b;
    layer0_outputs(822) <= a;
    layer0_outputs(823) <= not (a or b);
    layer0_outputs(824) <= a or b;
    layer0_outputs(825) <= b;
    layer0_outputs(826) <= b and not a;
    layer0_outputs(827) <= not b;
    layer0_outputs(828) <= not (a or b);
    layer0_outputs(829) <= a and not b;
    layer0_outputs(830) <= '1';
    layer0_outputs(831) <= '1';
    layer0_outputs(832) <= b;
    layer0_outputs(833) <= '1';
    layer0_outputs(834) <= a or b;
    layer0_outputs(835) <= not b or a;
    layer0_outputs(836) <= not (a or b);
    layer0_outputs(837) <= a and not b;
    layer0_outputs(838) <= b;
    layer0_outputs(839) <= a and not b;
    layer0_outputs(840) <= not a;
    layer0_outputs(841) <= not (a xor b);
    layer0_outputs(842) <= b;
    layer0_outputs(843) <= a and b;
    layer0_outputs(844) <= not b;
    layer0_outputs(845) <= a and not b;
    layer0_outputs(846) <= not b;
    layer0_outputs(847) <= not b or a;
    layer0_outputs(848) <= '0';
    layer0_outputs(849) <= not (a or b);
    layer0_outputs(850) <= not a or b;
    layer0_outputs(851) <= not (a xor b);
    layer0_outputs(852) <= a or b;
    layer0_outputs(853) <= a or b;
    layer0_outputs(854) <= not a or b;
    layer0_outputs(855) <= b;
    layer0_outputs(856) <= not (a or b);
    layer0_outputs(857) <= not (a and b);
    layer0_outputs(858) <= not b;
    layer0_outputs(859) <= not b;
    layer0_outputs(860) <= b and not a;
    layer0_outputs(861) <= not (a or b);
    layer0_outputs(862) <= a;
    layer0_outputs(863) <= not a;
    layer0_outputs(864) <= not b or a;
    layer0_outputs(865) <= not (a xor b);
    layer0_outputs(866) <= b and not a;
    layer0_outputs(867) <= not a or b;
    layer0_outputs(868) <= not (a or b);
    layer0_outputs(869) <= a xor b;
    layer0_outputs(870) <= a or b;
    layer0_outputs(871) <= not (a or b);
    layer0_outputs(872) <= not a or b;
    layer0_outputs(873) <= not b;
    layer0_outputs(874) <= not b;
    layer0_outputs(875) <= not (a or b);
    layer0_outputs(876) <= a;
    layer0_outputs(877) <= not (a or b);
    layer0_outputs(878) <= a xor b;
    layer0_outputs(879) <= a or b;
    layer0_outputs(880) <= b;
    layer0_outputs(881) <= not a or b;
    layer0_outputs(882) <= not (a xor b);
    layer0_outputs(883) <= not b;
    layer0_outputs(884) <= a or b;
    layer0_outputs(885) <= a and not b;
    layer0_outputs(886) <= not (a xor b);
    layer0_outputs(887) <= not (a or b);
    layer0_outputs(888) <= not (a xor b);
    layer0_outputs(889) <= not a;
    layer0_outputs(890) <= b;
    layer0_outputs(891) <= b and not a;
    layer0_outputs(892) <= a xor b;
    layer0_outputs(893) <= b and not a;
    layer0_outputs(894) <= a or b;
    layer0_outputs(895) <= a;
    layer0_outputs(896) <= b;
    layer0_outputs(897) <= not a or b;
    layer0_outputs(898) <= a;
    layer0_outputs(899) <= not b;
    layer0_outputs(900) <= not a or b;
    layer0_outputs(901) <= not (a or b);
    layer0_outputs(902) <= not a;
    layer0_outputs(903) <= '1';
    layer0_outputs(904) <= b and not a;
    layer0_outputs(905) <= not a or b;
    layer0_outputs(906) <= a and not b;
    layer0_outputs(907) <= a and b;
    layer0_outputs(908) <= b;
    layer0_outputs(909) <= a xor b;
    layer0_outputs(910) <= b;
    layer0_outputs(911) <= a;
    layer0_outputs(912) <= not (a xor b);
    layer0_outputs(913) <= a or b;
    layer0_outputs(914) <= b;
    layer0_outputs(915) <= not (a xor b);
    layer0_outputs(916) <= not (a or b);
    layer0_outputs(917) <= a and not b;
    layer0_outputs(918) <= not (a or b);
    layer0_outputs(919) <= a or b;
    layer0_outputs(920) <= a or b;
    layer0_outputs(921) <= a or b;
    layer0_outputs(922) <= not (a xor b);
    layer0_outputs(923) <= b;
    layer0_outputs(924) <= not b;
    layer0_outputs(925) <= a;
    layer0_outputs(926) <= not (a or b);
    layer0_outputs(927) <= a xor b;
    layer0_outputs(928) <= a;
    layer0_outputs(929) <= not (a xor b);
    layer0_outputs(930) <= not (a or b);
    layer0_outputs(931) <= a;
    layer0_outputs(932) <= a or b;
    layer0_outputs(933) <= not a or b;
    layer0_outputs(934) <= a;
    layer0_outputs(935) <= not a or b;
    layer0_outputs(936) <= a xor b;
    layer0_outputs(937) <= not (a or b);
    layer0_outputs(938) <= not b or a;
    layer0_outputs(939) <= a or b;
    layer0_outputs(940) <= not (a xor b);
    layer0_outputs(941) <= a xor b;
    layer0_outputs(942) <= a xor b;
    layer0_outputs(943) <= a xor b;
    layer0_outputs(944) <= b and not a;
    layer0_outputs(945) <= not a;
    layer0_outputs(946) <= a and not b;
    layer0_outputs(947) <= b;
    layer0_outputs(948) <= not b;
    layer0_outputs(949) <= not (a or b);
    layer0_outputs(950) <= a and not b;
    layer0_outputs(951) <= b;
    layer0_outputs(952) <= not (a and b);
    layer0_outputs(953) <= a or b;
    layer0_outputs(954) <= a or b;
    layer0_outputs(955) <= not (a xor b);
    layer0_outputs(956) <= not a or b;
    layer0_outputs(957) <= b;
    layer0_outputs(958) <= not (a xor b);
    layer0_outputs(959) <= not b;
    layer0_outputs(960) <= a or b;
    layer0_outputs(961) <= a or b;
    layer0_outputs(962) <= not b;
    layer0_outputs(963) <= b;
    layer0_outputs(964) <= a or b;
    layer0_outputs(965) <= not a;
    layer0_outputs(966) <= a xor b;
    layer0_outputs(967) <= b and not a;
    layer0_outputs(968) <= not (a or b);
    layer0_outputs(969) <= not a or b;
    layer0_outputs(970) <= not a;
    layer0_outputs(971) <= not a or b;
    layer0_outputs(972) <= not a;
    layer0_outputs(973) <= b;
    layer0_outputs(974) <= not (a or b);
    layer0_outputs(975) <= a or b;
    layer0_outputs(976) <= a and not b;
    layer0_outputs(977) <= a and not b;
    layer0_outputs(978) <= a xor b;
    layer0_outputs(979) <= not (a xor b);
    layer0_outputs(980) <= a and not b;
    layer0_outputs(981) <= not b;
    layer0_outputs(982) <= a and not b;
    layer0_outputs(983) <= '1';
    layer0_outputs(984) <= not (a or b);
    layer0_outputs(985) <= not (a or b);
    layer0_outputs(986) <= not a;
    layer0_outputs(987) <= a xor b;
    layer0_outputs(988) <= a or b;
    layer0_outputs(989) <= not a;
    layer0_outputs(990) <= not (a or b);
    layer0_outputs(991) <= '0';
    layer0_outputs(992) <= not (a or b);
    layer0_outputs(993) <= a or b;
    layer0_outputs(994) <= not a or b;
    layer0_outputs(995) <= '0';
    layer0_outputs(996) <= not (a or b);
    layer0_outputs(997) <= not (a or b);
    layer0_outputs(998) <= b;
    layer0_outputs(999) <= not b or a;
    layer0_outputs(1000) <= b and not a;
    layer0_outputs(1001) <= b and not a;
    layer0_outputs(1002) <= not a or b;
    layer0_outputs(1003) <= a xor b;
    layer0_outputs(1004) <= not (a and b);
    layer0_outputs(1005) <= b and not a;
    layer0_outputs(1006) <= a or b;
    layer0_outputs(1007) <= not (a xor b);
    layer0_outputs(1008) <= '1';
    layer0_outputs(1009) <= not (a xor b);
    layer0_outputs(1010) <= not (a xor b);
    layer0_outputs(1011) <= a xor b;
    layer0_outputs(1012) <= a;
    layer0_outputs(1013) <= not (a xor b);
    layer0_outputs(1014) <= not b or a;
    layer0_outputs(1015) <= not a or b;
    layer0_outputs(1016) <= not (a xor b);
    layer0_outputs(1017) <= b;
    layer0_outputs(1018) <= a or b;
    layer0_outputs(1019) <= not (a xor b);
    layer0_outputs(1020) <= a xor b;
    layer0_outputs(1021) <= b;
    layer0_outputs(1022) <= a and not b;
    layer0_outputs(1023) <= not (a xor b);
    layer0_outputs(1024) <= not (a xor b);
    layer0_outputs(1025) <= '0';
    layer0_outputs(1026) <= a;
    layer0_outputs(1027) <= a or b;
    layer0_outputs(1028) <= '0';
    layer0_outputs(1029) <= not b;
    layer0_outputs(1030) <= '1';
    layer0_outputs(1031) <= b and not a;
    layer0_outputs(1032) <= not b;
    layer0_outputs(1033) <= a or b;
    layer0_outputs(1034) <= a xor b;
    layer0_outputs(1035) <= not a;
    layer0_outputs(1036) <= not a;
    layer0_outputs(1037) <= b;
    layer0_outputs(1038) <= not b or a;
    layer0_outputs(1039) <= not a;
    layer0_outputs(1040) <= a xor b;
    layer0_outputs(1041) <= '0';
    layer0_outputs(1042) <= a or b;
    layer0_outputs(1043) <= b and not a;
    layer0_outputs(1044) <= not b;
    layer0_outputs(1045) <= not a or b;
    layer0_outputs(1046) <= not b;
    layer0_outputs(1047) <= not a;
    layer0_outputs(1048) <= a;
    layer0_outputs(1049) <= b;
    layer0_outputs(1050) <= not (a xor b);
    layer0_outputs(1051) <= not a or b;
    layer0_outputs(1052) <= not b or a;
    layer0_outputs(1053) <= not b;
    layer0_outputs(1054) <= a or b;
    layer0_outputs(1055) <= b;
    layer0_outputs(1056) <= not b;
    layer0_outputs(1057) <= not (a or b);
    layer0_outputs(1058) <= not a or b;
    layer0_outputs(1059) <= not (a xor b);
    layer0_outputs(1060) <= not a or b;
    layer0_outputs(1061) <= not b or a;
    layer0_outputs(1062) <= a;
    layer0_outputs(1063) <= b;
    layer0_outputs(1064) <= not a or b;
    layer0_outputs(1065) <= not (a xor b);
    layer0_outputs(1066) <= b;
    layer0_outputs(1067) <= not b or a;
    layer0_outputs(1068) <= not b;
    layer0_outputs(1069) <= not (a xor b);
    layer0_outputs(1070) <= a or b;
    layer0_outputs(1071) <= a;
    layer0_outputs(1072) <= not (a and b);
    layer0_outputs(1073) <= not b or a;
    layer0_outputs(1074) <= b;
    layer0_outputs(1075) <= a;
    layer0_outputs(1076) <= not b or a;
    layer0_outputs(1077) <= b;
    layer0_outputs(1078) <= not a or b;
    layer0_outputs(1079) <= not a;
    layer0_outputs(1080) <= a;
    layer0_outputs(1081) <= not (a or b);
    layer0_outputs(1082) <= a and b;
    layer0_outputs(1083) <= '0';
    layer0_outputs(1084) <= a or b;
    layer0_outputs(1085) <= not (a or b);
    layer0_outputs(1086) <= not b or a;
    layer0_outputs(1087) <= not (a xor b);
    layer0_outputs(1088) <= '0';
    layer0_outputs(1089) <= not (a xor b);
    layer0_outputs(1090) <= a and not b;
    layer0_outputs(1091) <= not a;
    layer0_outputs(1092) <= not b;
    layer0_outputs(1093) <= not b or a;
    layer0_outputs(1094) <= not a or b;
    layer0_outputs(1095) <= not a;
    layer0_outputs(1096) <= a and b;
    layer0_outputs(1097) <= '1';
    layer0_outputs(1098) <= not (a and b);
    layer0_outputs(1099) <= a xor b;
    layer0_outputs(1100) <= not b or a;
    layer0_outputs(1101) <= b;
    layer0_outputs(1102) <= b;
    layer0_outputs(1103) <= not (a or b);
    layer0_outputs(1104) <= not a;
    layer0_outputs(1105) <= not a;
    layer0_outputs(1106) <= a;
    layer0_outputs(1107) <= b and not a;
    layer0_outputs(1108) <= '1';
    layer0_outputs(1109) <= not (a or b);
    layer0_outputs(1110) <= not a or b;
    layer0_outputs(1111) <= not (a or b);
    layer0_outputs(1112) <= not (a or b);
    layer0_outputs(1113) <= a or b;
    layer0_outputs(1114) <= not b;
    layer0_outputs(1115) <= not (a and b);
    layer0_outputs(1116) <= a xor b;
    layer0_outputs(1117) <= a or b;
    layer0_outputs(1118) <= a xor b;
    layer0_outputs(1119) <= not (a xor b);
    layer0_outputs(1120) <= not (a or b);
    layer0_outputs(1121) <= a;
    layer0_outputs(1122) <= a or b;
    layer0_outputs(1123) <= not (a and b);
    layer0_outputs(1124) <= not (a and b);
    layer0_outputs(1125) <= not (a or b);
    layer0_outputs(1126) <= a xor b;
    layer0_outputs(1127) <= not (a or b);
    layer0_outputs(1128) <= not a;
    layer0_outputs(1129) <= not b;
    layer0_outputs(1130) <= not a;
    layer0_outputs(1131) <= a or b;
    layer0_outputs(1132) <= b;
    layer0_outputs(1133) <= a;
    layer0_outputs(1134) <= not a or b;
    layer0_outputs(1135) <= not a;
    layer0_outputs(1136) <= not (a xor b);
    layer0_outputs(1137) <= not (a and b);
    layer0_outputs(1138) <= a and not b;
    layer0_outputs(1139) <= not b;
    layer0_outputs(1140) <= not a;
    layer0_outputs(1141) <= not a or b;
    layer0_outputs(1142) <= not a;
    layer0_outputs(1143) <= not (a xor b);
    layer0_outputs(1144) <= not (a and b);
    layer0_outputs(1145) <= a or b;
    layer0_outputs(1146) <= a and not b;
    layer0_outputs(1147) <= a and b;
    layer0_outputs(1148) <= b;
    layer0_outputs(1149) <= not a;
    layer0_outputs(1150) <= b and not a;
    layer0_outputs(1151) <= not a;
    layer0_outputs(1152) <= not (a or b);
    layer0_outputs(1153) <= not (a or b);
    layer0_outputs(1154) <= not a;
    layer0_outputs(1155) <= a;
    layer0_outputs(1156) <= b;
    layer0_outputs(1157) <= a xor b;
    layer0_outputs(1158) <= a;
    layer0_outputs(1159) <= a;
    layer0_outputs(1160) <= not (a or b);
    layer0_outputs(1161) <= not a or b;
    layer0_outputs(1162) <= b;
    layer0_outputs(1163) <= not (a or b);
    layer0_outputs(1164) <= '1';
    layer0_outputs(1165) <= a and not b;
    layer0_outputs(1166) <= not (a xor b);
    layer0_outputs(1167) <= a;
    layer0_outputs(1168) <= a or b;
    layer0_outputs(1169) <= not b;
    layer0_outputs(1170) <= a;
    layer0_outputs(1171) <= not a or b;
    layer0_outputs(1172) <= not b or a;
    layer0_outputs(1173) <= a or b;
    layer0_outputs(1174) <= not (a xor b);
    layer0_outputs(1175) <= not (a or b);
    layer0_outputs(1176) <= '1';
    layer0_outputs(1177) <= a and not b;
    layer0_outputs(1178) <= a and not b;
    layer0_outputs(1179) <= '1';
    layer0_outputs(1180) <= not a;
    layer0_outputs(1181) <= not b or a;
    layer0_outputs(1182) <= not (a or b);
    layer0_outputs(1183) <= b and not a;
    layer0_outputs(1184) <= b;
    layer0_outputs(1185) <= not a;
    layer0_outputs(1186) <= a and not b;
    layer0_outputs(1187) <= not (a or b);
    layer0_outputs(1188) <= '0';
    layer0_outputs(1189) <= a and b;
    layer0_outputs(1190) <= not a or b;
    layer0_outputs(1191) <= a and b;
    layer0_outputs(1192) <= b;
    layer0_outputs(1193) <= not (a or b);
    layer0_outputs(1194) <= a or b;
    layer0_outputs(1195) <= a xor b;
    layer0_outputs(1196) <= not (a or b);
    layer0_outputs(1197) <= not (a xor b);
    layer0_outputs(1198) <= a or b;
    layer0_outputs(1199) <= not (a or b);
    layer0_outputs(1200) <= a;
    layer0_outputs(1201) <= not (a xor b);
    layer0_outputs(1202) <= not a or b;
    layer0_outputs(1203) <= not a;
    layer0_outputs(1204) <= not b;
    layer0_outputs(1205) <= b;
    layer0_outputs(1206) <= a or b;
    layer0_outputs(1207) <= b;
    layer0_outputs(1208) <= a;
    layer0_outputs(1209) <= '1';
    layer0_outputs(1210) <= not b or a;
    layer0_outputs(1211) <= a;
    layer0_outputs(1212) <= '1';
    layer0_outputs(1213) <= a;
    layer0_outputs(1214) <= not a;
    layer0_outputs(1215) <= not (a or b);
    layer0_outputs(1216) <= b and not a;
    layer0_outputs(1217) <= a and not b;
    layer0_outputs(1218) <= not a or b;
    layer0_outputs(1219) <= a xor b;
    layer0_outputs(1220) <= not a;
    layer0_outputs(1221) <= a and not b;
    layer0_outputs(1222) <= b and not a;
    layer0_outputs(1223) <= not b;
    layer0_outputs(1224) <= a xor b;
    layer0_outputs(1225) <= a;
    layer0_outputs(1226) <= not a;
    layer0_outputs(1227) <= not b;
    layer0_outputs(1228) <= a xor b;
    layer0_outputs(1229) <= not a;
    layer0_outputs(1230) <= a and not b;
    layer0_outputs(1231) <= not (a or b);
    layer0_outputs(1232) <= a or b;
    layer0_outputs(1233) <= not (a or b);
    layer0_outputs(1234) <= not (a or b);
    layer0_outputs(1235) <= not (a xor b);
    layer0_outputs(1236) <= a;
    layer0_outputs(1237) <= a xor b;
    layer0_outputs(1238) <= a xor b;
    layer0_outputs(1239) <= not (a xor b);
    layer0_outputs(1240) <= a;
    layer0_outputs(1241) <= a or b;
    layer0_outputs(1242) <= not (a or b);
    layer0_outputs(1243) <= not a or b;
    layer0_outputs(1244) <= not (a xor b);
    layer0_outputs(1245) <= not b;
    layer0_outputs(1246) <= not (a xor b);
    layer0_outputs(1247) <= not a or b;
    layer0_outputs(1248) <= not (a xor b);
    layer0_outputs(1249) <= a xor b;
    layer0_outputs(1250) <= a or b;
    layer0_outputs(1251) <= not (a or b);
    layer0_outputs(1252) <= '0';
    layer0_outputs(1253) <= b;
    layer0_outputs(1254) <= a xor b;
    layer0_outputs(1255) <= not (a or b);
    layer0_outputs(1256) <= a and b;
    layer0_outputs(1257) <= a and not b;
    layer0_outputs(1258) <= a;
    layer0_outputs(1259) <= b and not a;
    layer0_outputs(1260) <= not b;
    layer0_outputs(1261) <= '1';
    layer0_outputs(1262) <= a or b;
    layer0_outputs(1263) <= not a;
    layer0_outputs(1264) <= a or b;
    layer0_outputs(1265) <= not (a or b);
    layer0_outputs(1266) <= b and not a;
    layer0_outputs(1267) <= a and not b;
    layer0_outputs(1268) <= a and b;
    layer0_outputs(1269) <= a or b;
    layer0_outputs(1270) <= '0';
    layer0_outputs(1271) <= '1';
    layer0_outputs(1272) <= not (a or b);
    layer0_outputs(1273) <= a or b;
    layer0_outputs(1274) <= not (a xor b);
    layer0_outputs(1275) <= b and not a;
    layer0_outputs(1276) <= not (a or b);
    layer0_outputs(1277) <= not a;
    layer0_outputs(1278) <= a or b;
    layer0_outputs(1279) <= '0';
    layer0_outputs(1280) <= not (a xor b);
    layer0_outputs(1281) <= not b or a;
    layer0_outputs(1282) <= a and not b;
    layer0_outputs(1283) <= '1';
    layer0_outputs(1284) <= not (a or b);
    layer0_outputs(1285) <= not (a or b);
    layer0_outputs(1286) <= a and b;
    layer0_outputs(1287) <= b;
    layer0_outputs(1288) <= a xor b;
    layer0_outputs(1289) <= not (a and b);
    layer0_outputs(1290) <= a;
    layer0_outputs(1291) <= not b or a;
    layer0_outputs(1292) <= a xor b;
    layer0_outputs(1293) <= not (a and b);
    layer0_outputs(1294) <= '0';
    layer0_outputs(1295) <= a or b;
    layer0_outputs(1296) <= a xor b;
    layer0_outputs(1297) <= a xor b;
    layer0_outputs(1298) <= '0';
    layer0_outputs(1299) <= a and not b;
    layer0_outputs(1300) <= not a;
    layer0_outputs(1301) <= a xor b;
    layer0_outputs(1302) <= not b;
    layer0_outputs(1303) <= b;
    layer0_outputs(1304) <= a;
    layer0_outputs(1305) <= not a;
    layer0_outputs(1306) <= b;
    layer0_outputs(1307) <= not (a xor b);
    layer0_outputs(1308) <= a xor b;
    layer0_outputs(1309) <= not (a and b);
    layer0_outputs(1310) <= not b or a;
    layer0_outputs(1311) <= a and not b;
    layer0_outputs(1312) <= not a;
    layer0_outputs(1313) <= not (a xor b);
    layer0_outputs(1314) <= '0';
    layer0_outputs(1315) <= a xor b;
    layer0_outputs(1316) <= not (a or b);
    layer0_outputs(1317) <= not (a and b);
    layer0_outputs(1318) <= a and not b;
    layer0_outputs(1319) <= a xor b;
    layer0_outputs(1320) <= a and not b;
    layer0_outputs(1321) <= not b or a;
    layer0_outputs(1322) <= '1';
    layer0_outputs(1323) <= not (a or b);
    layer0_outputs(1324) <= a or b;
    layer0_outputs(1325) <= a or b;
    layer0_outputs(1326) <= a and not b;
    layer0_outputs(1327) <= '0';
    layer0_outputs(1328) <= b;
    layer0_outputs(1329) <= not a or b;
    layer0_outputs(1330) <= a xor b;
    layer0_outputs(1331) <= a;
    layer0_outputs(1332) <= not a or b;
    layer0_outputs(1333) <= not a or b;
    layer0_outputs(1334) <= not (a and b);
    layer0_outputs(1335) <= '0';
    layer0_outputs(1336) <= not (a xor b);
    layer0_outputs(1337) <= a or b;
    layer0_outputs(1338) <= a or b;
    layer0_outputs(1339) <= b;
    layer0_outputs(1340) <= not b;
    layer0_outputs(1341) <= b;
    layer0_outputs(1342) <= a xor b;
    layer0_outputs(1343) <= not (a or b);
    layer0_outputs(1344) <= a or b;
    layer0_outputs(1345) <= not a;
    layer0_outputs(1346) <= not (a or b);
    layer0_outputs(1347) <= a xor b;
    layer0_outputs(1348) <= not a or b;
    layer0_outputs(1349) <= a xor b;
    layer0_outputs(1350) <= not a or b;
    layer0_outputs(1351) <= not (a or b);
    layer0_outputs(1352) <= not a;
    layer0_outputs(1353) <= not (a or b);
    layer0_outputs(1354) <= not (a or b);
    layer0_outputs(1355) <= a;
    layer0_outputs(1356) <= a and not b;
    layer0_outputs(1357) <= '1';
    layer0_outputs(1358) <= not b;
    layer0_outputs(1359) <= not (a and b);
    layer0_outputs(1360) <= not b;
    layer0_outputs(1361) <= a xor b;
    layer0_outputs(1362) <= a and not b;
    layer0_outputs(1363) <= a or b;
    layer0_outputs(1364) <= a or b;
    layer0_outputs(1365) <= not b;
    layer0_outputs(1366) <= not (a or b);
    layer0_outputs(1367) <= b and not a;
    layer0_outputs(1368) <= a xor b;
    layer0_outputs(1369) <= '1';
    layer0_outputs(1370) <= not (a xor b);
    layer0_outputs(1371) <= a or b;
    layer0_outputs(1372) <= not (a or b);
    layer0_outputs(1373) <= b;
    layer0_outputs(1374) <= a xor b;
    layer0_outputs(1375) <= not a;
    layer0_outputs(1376) <= not b or a;
    layer0_outputs(1377) <= a xor b;
    layer0_outputs(1378) <= a or b;
    layer0_outputs(1379) <= not (a xor b);
    layer0_outputs(1380) <= not b or a;
    layer0_outputs(1381) <= not a or b;
    layer0_outputs(1382) <= b and not a;
    layer0_outputs(1383) <= a;
    layer0_outputs(1384) <= a or b;
    layer0_outputs(1385) <= a xor b;
    layer0_outputs(1386) <= not a;
    layer0_outputs(1387) <= a and not b;
    layer0_outputs(1388) <= a and not b;
    layer0_outputs(1389) <= a xor b;
    layer0_outputs(1390) <= not (a and b);
    layer0_outputs(1391) <= '1';
    layer0_outputs(1392) <= not a or b;
    layer0_outputs(1393) <= b and not a;
    layer0_outputs(1394) <= not b or a;
    layer0_outputs(1395) <= not (a or b);
    layer0_outputs(1396) <= a xor b;
    layer0_outputs(1397) <= not (a xor b);
    layer0_outputs(1398) <= not (a xor b);
    layer0_outputs(1399) <= a and not b;
    layer0_outputs(1400) <= a and not b;
    layer0_outputs(1401) <= b;
    layer0_outputs(1402) <= not b or a;
    layer0_outputs(1403) <= b and not a;
    layer0_outputs(1404) <= a or b;
    layer0_outputs(1405) <= not (a xor b);
    layer0_outputs(1406) <= b and not a;
    layer0_outputs(1407) <= b and not a;
    layer0_outputs(1408) <= not (a xor b);
    layer0_outputs(1409) <= '1';
    layer0_outputs(1410) <= b and not a;
    layer0_outputs(1411) <= a or b;
    layer0_outputs(1412) <= a xor b;
    layer0_outputs(1413) <= not a;
    layer0_outputs(1414) <= b and not a;
    layer0_outputs(1415) <= not a or b;
    layer0_outputs(1416) <= a and not b;
    layer0_outputs(1417) <= not (a and b);
    layer0_outputs(1418) <= not b or a;
    layer0_outputs(1419) <= a or b;
    layer0_outputs(1420) <= a xor b;
    layer0_outputs(1421) <= b and not a;
    layer0_outputs(1422) <= not (a or b);
    layer0_outputs(1423) <= not (a or b);
    layer0_outputs(1424) <= a and not b;
    layer0_outputs(1425) <= not b or a;
    layer0_outputs(1426) <= a or b;
    layer0_outputs(1427) <= b;
    layer0_outputs(1428) <= a;
    layer0_outputs(1429) <= b;
    layer0_outputs(1430) <= not b;
    layer0_outputs(1431) <= not b;
    layer0_outputs(1432) <= not (a or b);
    layer0_outputs(1433) <= a xor b;
    layer0_outputs(1434) <= not b or a;
    layer0_outputs(1435) <= '1';
    layer0_outputs(1436) <= not b or a;
    layer0_outputs(1437) <= not a or b;
    layer0_outputs(1438) <= b;
    layer0_outputs(1439) <= a and not b;
    layer0_outputs(1440) <= not a;
    layer0_outputs(1441) <= a;
    layer0_outputs(1442) <= a;
    layer0_outputs(1443) <= not (a or b);
    layer0_outputs(1444) <= not b;
    layer0_outputs(1445) <= a;
    layer0_outputs(1446) <= a and not b;
    layer0_outputs(1447) <= not (a or b);
    layer0_outputs(1448) <= not a or b;
    layer0_outputs(1449) <= not a or b;
    layer0_outputs(1450) <= b;
    layer0_outputs(1451) <= not a or b;
    layer0_outputs(1452) <= a and not b;
    layer0_outputs(1453) <= b and not a;
    layer0_outputs(1454) <= not a or b;
    layer0_outputs(1455) <= not b;
    layer0_outputs(1456) <= a xor b;
    layer0_outputs(1457) <= '0';
    layer0_outputs(1458) <= '1';
    layer0_outputs(1459) <= a and b;
    layer0_outputs(1460) <= not (a or b);
    layer0_outputs(1461) <= a and b;
    layer0_outputs(1462) <= not b;
    layer0_outputs(1463) <= not (a or b);
    layer0_outputs(1464) <= not (a xor b);
    layer0_outputs(1465) <= a or b;
    layer0_outputs(1466) <= a;
    layer0_outputs(1467) <= not a or b;
    layer0_outputs(1468) <= a;
    layer0_outputs(1469) <= not (a and b);
    layer0_outputs(1470) <= b and not a;
    layer0_outputs(1471) <= a or b;
    layer0_outputs(1472) <= a;
    layer0_outputs(1473) <= not (a or b);
    layer0_outputs(1474) <= not b;
    layer0_outputs(1475) <= '1';
    layer0_outputs(1476) <= not b or a;
    layer0_outputs(1477) <= a xor b;
    layer0_outputs(1478) <= a or b;
    layer0_outputs(1479) <= not a;
    layer0_outputs(1480) <= b and not a;
    layer0_outputs(1481) <= '0';
    layer0_outputs(1482) <= a and not b;
    layer0_outputs(1483) <= b and not a;
    layer0_outputs(1484) <= not (a or b);
    layer0_outputs(1485) <= not (a xor b);
    layer0_outputs(1486) <= not a or b;
    layer0_outputs(1487) <= a;
    layer0_outputs(1488) <= not (a or b);
    layer0_outputs(1489) <= b and not a;
    layer0_outputs(1490) <= a;
    layer0_outputs(1491) <= not (a xor b);
    layer0_outputs(1492) <= not (a xor b);
    layer0_outputs(1493) <= a xor b;
    layer0_outputs(1494) <= a xor b;
    layer0_outputs(1495) <= a and b;
    layer0_outputs(1496) <= not a;
    layer0_outputs(1497) <= a xor b;
    layer0_outputs(1498) <= a and not b;
    layer0_outputs(1499) <= a and not b;
    layer0_outputs(1500) <= not (a and b);
    layer0_outputs(1501) <= b;
    layer0_outputs(1502) <= not (a or b);
    layer0_outputs(1503) <= not a or b;
    layer0_outputs(1504) <= not (a or b);
    layer0_outputs(1505) <= a and not b;
    layer0_outputs(1506) <= not (a or b);
    layer0_outputs(1507) <= not b;
    layer0_outputs(1508) <= a xor b;
    layer0_outputs(1509) <= not (a xor b);
    layer0_outputs(1510) <= a or b;
    layer0_outputs(1511) <= not b;
    layer0_outputs(1512) <= b;
    layer0_outputs(1513) <= not (a or b);
    layer0_outputs(1514) <= b;
    layer0_outputs(1515) <= not (a or b);
    layer0_outputs(1516) <= not (a or b);
    layer0_outputs(1517) <= a or b;
    layer0_outputs(1518) <= '1';
    layer0_outputs(1519) <= not a;
    layer0_outputs(1520) <= a or b;
    layer0_outputs(1521) <= not b or a;
    layer0_outputs(1522) <= not a or b;
    layer0_outputs(1523) <= b;
    layer0_outputs(1524) <= b and not a;
    layer0_outputs(1525) <= '0';
    layer0_outputs(1526) <= a;
    layer0_outputs(1527) <= b;
    layer0_outputs(1528) <= b and not a;
    layer0_outputs(1529) <= a and not b;
    layer0_outputs(1530) <= b and not a;
    layer0_outputs(1531) <= not a;
    layer0_outputs(1532) <= a xor b;
    layer0_outputs(1533) <= b;
    layer0_outputs(1534) <= b and not a;
    layer0_outputs(1535) <= not (a xor b);
    layer0_outputs(1536) <= a;
    layer0_outputs(1537) <= not b;
    layer0_outputs(1538) <= not a or b;
    layer0_outputs(1539) <= not (a and b);
    layer0_outputs(1540) <= a and not b;
    layer0_outputs(1541) <= b and not a;
    layer0_outputs(1542) <= '0';
    layer0_outputs(1543) <= not a;
    layer0_outputs(1544) <= not a or b;
    layer0_outputs(1545) <= not b or a;
    layer0_outputs(1546) <= '1';
    layer0_outputs(1547) <= not (a or b);
    layer0_outputs(1548) <= a or b;
    layer0_outputs(1549) <= b and not a;
    layer0_outputs(1550) <= a;
    layer0_outputs(1551) <= not (a or b);
    layer0_outputs(1552) <= not (a and b);
    layer0_outputs(1553) <= not (a xor b);
    layer0_outputs(1554) <= not b;
    layer0_outputs(1555) <= b;
    layer0_outputs(1556) <= b;
    layer0_outputs(1557) <= not (a xor b);
    layer0_outputs(1558) <= not b or a;
    layer0_outputs(1559) <= a xor b;
    layer0_outputs(1560) <= a xor b;
    layer0_outputs(1561) <= a;
    layer0_outputs(1562) <= not (a xor b);
    layer0_outputs(1563) <= not a;
    layer0_outputs(1564) <= not a;
    layer0_outputs(1565) <= a xor b;
    layer0_outputs(1566) <= not a;
    layer0_outputs(1567) <= a xor b;
    layer0_outputs(1568) <= a xor b;
    layer0_outputs(1569) <= b and not a;
    layer0_outputs(1570) <= not a;
    layer0_outputs(1571) <= not b;
    layer0_outputs(1572) <= not a;
    layer0_outputs(1573) <= b;
    layer0_outputs(1574) <= b;
    layer0_outputs(1575) <= not (a or b);
    layer0_outputs(1576) <= a or b;
    layer0_outputs(1577) <= not b;
    layer0_outputs(1578) <= a;
    layer0_outputs(1579) <= not (a xor b);
    layer0_outputs(1580) <= a;
    layer0_outputs(1581) <= a or b;
    layer0_outputs(1582) <= not a or b;
    layer0_outputs(1583) <= not b;
    layer0_outputs(1584) <= a or b;
    layer0_outputs(1585) <= '1';
    layer0_outputs(1586) <= not b;
    layer0_outputs(1587) <= a and not b;
    layer0_outputs(1588) <= b and not a;
    layer0_outputs(1589) <= b and not a;
    layer0_outputs(1590) <= not (a or b);
    layer0_outputs(1591) <= b and not a;
    layer0_outputs(1592) <= b;
    layer0_outputs(1593) <= not (a and b);
    layer0_outputs(1594) <= not (a xor b);
    layer0_outputs(1595) <= '1';
    layer0_outputs(1596) <= not (a or b);
    layer0_outputs(1597) <= b and not a;
    layer0_outputs(1598) <= not b or a;
    layer0_outputs(1599) <= a;
    layer0_outputs(1600) <= not (a and b);
    layer0_outputs(1601) <= not b;
    layer0_outputs(1602) <= a;
    layer0_outputs(1603) <= '0';
    layer0_outputs(1604) <= not (a or b);
    layer0_outputs(1605) <= b and not a;
    layer0_outputs(1606) <= not a;
    layer0_outputs(1607) <= b;
    layer0_outputs(1608) <= a or b;
    layer0_outputs(1609) <= not (a or b);
    layer0_outputs(1610) <= b;
    layer0_outputs(1611) <= not a;
    layer0_outputs(1612) <= not b;
    layer0_outputs(1613) <= not (a or b);
    layer0_outputs(1614) <= not b or a;
    layer0_outputs(1615) <= a xor b;
    layer0_outputs(1616) <= not (a xor b);
    layer0_outputs(1617) <= '1';
    layer0_outputs(1618) <= a and not b;
    layer0_outputs(1619) <= a or b;
    layer0_outputs(1620) <= not (a and b);
    layer0_outputs(1621) <= not (a or b);
    layer0_outputs(1622) <= a xor b;
    layer0_outputs(1623) <= not (a or b);
    layer0_outputs(1624) <= b and not a;
    layer0_outputs(1625) <= not a or b;
    layer0_outputs(1626) <= a xor b;
    layer0_outputs(1627) <= not (a or b);
    layer0_outputs(1628) <= not a or b;
    layer0_outputs(1629) <= not a or b;
    layer0_outputs(1630) <= a xor b;
    layer0_outputs(1631) <= not (a or b);
    layer0_outputs(1632) <= not b;
    layer0_outputs(1633) <= not b or a;
    layer0_outputs(1634) <= not b;
    layer0_outputs(1635) <= '0';
    layer0_outputs(1636) <= b and not a;
    layer0_outputs(1637) <= a or b;
    layer0_outputs(1638) <= a and not b;
    layer0_outputs(1639) <= b and not a;
    layer0_outputs(1640) <= not a or b;
    layer0_outputs(1641) <= not b or a;
    layer0_outputs(1642) <= a or b;
    layer0_outputs(1643) <= a or b;
    layer0_outputs(1644) <= a xor b;
    layer0_outputs(1645) <= b and not a;
    layer0_outputs(1646) <= a and not b;
    layer0_outputs(1647) <= not (a xor b);
    layer0_outputs(1648) <= b and not a;
    layer0_outputs(1649) <= a and not b;
    layer0_outputs(1650) <= not b or a;
    layer0_outputs(1651) <= a or b;
    layer0_outputs(1652) <= b and not a;
    layer0_outputs(1653) <= not b;
    layer0_outputs(1654) <= '0';
    layer0_outputs(1655) <= not a or b;
    layer0_outputs(1656) <= not b or a;
    layer0_outputs(1657) <= b and not a;
    layer0_outputs(1658) <= not b;
    layer0_outputs(1659) <= not (a or b);
    layer0_outputs(1660) <= not (a or b);
    layer0_outputs(1661) <= a;
    layer0_outputs(1662) <= b;
    layer0_outputs(1663) <= a or b;
    layer0_outputs(1664) <= b;
    layer0_outputs(1665) <= not (a xor b);
    layer0_outputs(1666) <= not a;
    layer0_outputs(1667) <= not a or b;
    layer0_outputs(1668) <= a;
    layer0_outputs(1669) <= a;
    layer0_outputs(1670) <= not (a xor b);
    layer0_outputs(1671) <= not (a or b);
    layer0_outputs(1672) <= not b;
    layer0_outputs(1673) <= a;
    layer0_outputs(1674) <= not (a xor b);
    layer0_outputs(1675) <= b and not a;
    layer0_outputs(1676) <= a or b;
    layer0_outputs(1677) <= not (a or b);
    layer0_outputs(1678) <= a or b;
    layer0_outputs(1679) <= a or b;
    layer0_outputs(1680) <= a;
    layer0_outputs(1681) <= a xor b;
    layer0_outputs(1682) <= not (a and b);
    layer0_outputs(1683) <= a or b;
    layer0_outputs(1684) <= a and not b;
    layer0_outputs(1685) <= not b;
    layer0_outputs(1686) <= not a;
    layer0_outputs(1687) <= b;
    layer0_outputs(1688) <= not (a xor b);
    layer0_outputs(1689) <= not (a or b);
    layer0_outputs(1690) <= not (a and b);
    layer0_outputs(1691) <= not (a or b);
    layer0_outputs(1692) <= a xor b;
    layer0_outputs(1693) <= a and not b;
    layer0_outputs(1694) <= a or b;
    layer0_outputs(1695) <= not a;
    layer0_outputs(1696) <= not a or b;
    layer0_outputs(1697) <= a or b;
    layer0_outputs(1698) <= a;
    layer0_outputs(1699) <= not (a and b);
    layer0_outputs(1700) <= '1';
    layer0_outputs(1701) <= a or b;
    layer0_outputs(1702) <= not (a and b);
    layer0_outputs(1703) <= not a;
    layer0_outputs(1704) <= not a or b;
    layer0_outputs(1705) <= a and b;
    layer0_outputs(1706) <= not b;
    layer0_outputs(1707) <= not (a or b);
    layer0_outputs(1708) <= a;
    layer0_outputs(1709) <= not (a and b);
    layer0_outputs(1710) <= a;
    layer0_outputs(1711) <= b;
    layer0_outputs(1712) <= a xor b;
    layer0_outputs(1713) <= not a;
    layer0_outputs(1714) <= not b;
    layer0_outputs(1715) <= b and not a;
    layer0_outputs(1716) <= b;
    layer0_outputs(1717) <= b;
    layer0_outputs(1718) <= not b;
    layer0_outputs(1719) <= a xor b;
    layer0_outputs(1720) <= not (a or b);
    layer0_outputs(1721) <= a xor b;
    layer0_outputs(1722) <= not a or b;
    layer0_outputs(1723) <= not a;
    layer0_outputs(1724) <= not (a and b);
    layer0_outputs(1725) <= not b;
    layer0_outputs(1726) <= b and not a;
    layer0_outputs(1727) <= b and not a;
    layer0_outputs(1728) <= not b;
    layer0_outputs(1729) <= a xor b;
    layer0_outputs(1730) <= b;
    layer0_outputs(1731) <= not a;
    layer0_outputs(1732) <= a or b;
    layer0_outputs(1733) <= '0';
    layer0_outputs(1734) <= not (a or b);
    layer0_outputs(1735) <= a or b;
    layer0_outputs(1736) <= not (a or b);
    layer0_outputs(1737) <= not (a or b);
    layer0_outputs(1738) <= a and not b;
    layer0_outputs(1739) <= a xor b;
    layer0_outputs(1740) <= a;
    layer0_outputs(1741) <= a or b;
    layer0_outputs(1742) <= not b;
    layer0_outputs(1743) <= b and not a;
    layer0_outputs(1744) <= not (a or b);
    layer0_outputs(1745) <= a or b;
    layer0_outputs(1746) <= '1';
    layer0_outputs(1747) <= a;
    layer0_outputs(1748) <= a or b;
    layer0_outputs(1749) <= not (a or b);
    layer0_outputs(1750) <= a and not b;
    layer0_outputs(1751) <= not (a or b);
    layer0_outputs(1752) <= not a or b;
    layer0_outputs(1753) <= a and b;
    layer0_outputs(1754) <= not (a or b);
    layer0_outputs(1755) <= a xor b;
    layer0_outputs(1756) <= not a;
    layer0_outputs(1757) <= not b;
    layer0_outputs(1758) <= not a;
    layer0_outputs(1759) <= not (a and b);
    layer0_outputs(1760) <= a xor b;
    layer0_outputs(1761) <= not b;
    layer0_outputs(1762) <= not (a or b);
    layer0_outputs(1763) <= not a;
    layer0_outputs(1764) <= a;
    layer0_outputs(1765) <= not (a xor b);
    layer0_outputs(1766) <= a and not b;
    layer0_outputs(1767) <= a;
    layer0_outputs(1768) <= b;
    layer0_outputs(1769) <= a;
    layer0_outputs(1770) <= not a or b;
    layer0_outputs(1771) <= a;
    layer0_outputs(1772) <= not (a and b);
    layer0_outputs(1773) <= not b or a;
    layer0_outputs(1774) <= not a or b;
    layer0_outputs(1775) <= a or b;
    layer0_outputs(1776) <= a;
    layer0_outputs(1777) <= '0';
    layer0_outputs(1778) <= not a or b;
    layer0_outputs(1779) <= not a;
    layer0_outputs(1780) <= not a;
    layer0_outputs(1781) <= not b;
    layer0_outputs(1782) <= b;
    layer0_outputs(1783) <= b;
    layer0_outputs(1784) <= a xor b;
    layer0_outputs(1785) <= not b;
    layer0_outputs(1786) <= a or b;
    layer0_outputs(1787) <= not (a or b);
    layer0_outputs(1788) <= a;
    layer0_outputs(1789) <= a;
    layer0_outputs(1790) <= '0';
    layer0_outputs(1791) <= a and not b;
    layer0_outputs(1792) <= not b or a;
    layer0_outputs(1793) <= '1';
    layer0_outputs(1794) <= not (a xor b);
    layer0_outputs(1795) <= a or b;
    layer0_outputs(1796) <= a or b;
    layer0_outputs(1797) <= a xor b;
    layer0_outputs(1798) <= a and not b;
    layer0_outputs(1799) <= not (a and b);
    layer0_outputs(1800) <= not a;
    layer0_outputs(1801) <= not b;
    layer0_outputs(1802) <= not (a xor b);
    layer0_outputs(1803) <= not (a or b);
    layer0_outputs(1804) <= not (a or b);
    layer0_outputs(1805) <= a and not b;
    layer0_outputs(1806) <= a and not b;
    layer0_outputs(1807) <= b and not a;
    layer0_outputs(1808) <= a or b;
    layer0_outputs(1809) <= a or b;
    layer0_outputs(1810) <= not (a or b);
    layer0_outputs(1811) <= a xor b;
    layer0_outputs(1812) <= b;
    layer0_outputs(1813) <= b;
    layer0_outputs(1814) <= not a;
    layer0_outputs(1815) <= not a;
    layer0_outputs(1816) <= not (a or b);
    layer0_outputs(1817) <= b;
    layer0_outputs(1818) <= not b;
    layer0_outputs(1819) <= not b or a;
    layer0_outputs(1820) <= a and not b;
    layer0_outputs(1821) <= a;
    layer0_outputs(1822) <= a;
    layer0_outputs(1823) <= a or b;
    layer0_outputs(1824) <= not a;
    layer0_outputs(1825) <= a and b;
    layer0_outputs(1826) <= a xor b;
    layer0_outputs(1827) <= not b or a;
    layer0_outputs(1828) <= not b or a;
    layer0_outputs(1829) <= not (a xor b);
    layer0_outputs(1830) <= not (a or b);
    layer0_outputs(1831) <= a xor b;
    layer0_outputs(1832) <= not (a or b);
    layer0_outputs(1833) <= not (a and b);
    layer0_outputs(1834) <= not b or a;
    layer0_outputs(1835) <= b;
    layer0_outputs(1836) <= not (a xor b);
    layer0_outputs(1837) <= not (a or b);
    layer0_outputs(1838) <= not b or a;
    layer0_outputs(1839) <= '1';
    layer0_outputs(1840) <= not (a xor b);
    layer0_outputs(1841) <= a and not b;
    layer0_outputs(1842) <= not b;
    layer0_outputs(1843) <= a xor b;
    layer0_outputs(1844) <= '1';
    layer0_outputs(1845) <= a and not b;
    layer0_outputs(1846) <= not b;
    layer0_outputs(1847) <= not a or b;
    layer0_outputs(1848) <= b and not a;
    layer0_outputs(1849) <= a xor b;
    layer0_outputs(1850) <= a or b;
    layer0_outputs(1851) <= a xor b;
    layer0_outputs(1852) <= not a or b;
    layer0_outputs(1853) <= not a;
    layer0_outputs(1854) <= not b or a;
    layer0_outputs(1855) <= not (a or b);
    layer0_outputs(1856) <= not a or b;
    layer0_outputs(1857) <= b and not a;
    layer0_outputs(1858) <= a xor b;
    layer0_outputs(1859) <= a;
    layer0_outputs(1860) <= '1';
    layer0_outputs(1861) <= not (a xor b);
    layer0_outputs(1862) <= a;
    layer0_outputs(1863) <= not a or b;
    layer0_outputs(1864) <= b and not a;
    layer0_outputs(1865) <= b and not a;
    layer0_outputs(1866) <= a xor b;
    layer0_outputs(1867) <= b and not a;
    layer0_outputs(1868) <= a xor b;
    layer0_outputs(1869) <= a xor b;
    layer0_outputs(1870) <= not (a or b);
    layer0_outputs(1871) <= not a or b;
    layer0_outputs(1872) <= not a;
    layer0_outputs(1873) <= not a;
    layer0_outputs(1874) <= not a;
    layer0_outputs(1875) <= a xor b;
    layer0_outputs(1876) <= not (a xor b);
    layer0_outputs(1877) <= a or b;
    layer0_outputs(1878) <= a or b;
    layer0_outputs(1879) <= not b;
    layer0_outputs(1880) <= not a or b;
    layer0_outputs(1881) <= not b;
    layer0_outputs(1882) <= not a or b;
    layer0_outputs(1883) <= not a;
    layer0_outputs(1884) <= b;
    layer0_outputs(1885) <= not (a or b);
    layer0_outputs(1886) <= a xor b;
    layer0_outputs(1887) <= not a;
    layer0_outputs(1888) <= not b or a;
    layer0_outputs(1889) <= a or b;
    layer0_outputs(1890) <= not b or a;
    layer0_outputs(1891) <= not b;
    layer0_outputs(1892) <= a;
    layer0_outputs(1893) <= b and not a;
    layer0_outputs(1894) <= not a or b;
    layer0_outputs(1895) <= not b;
    layer0_outputs(1896) <= b and not a;
    layer0_outputs(1897) <= a and not b;
    layer0_outputs(1898) <= not (a xor b);
    layer0_outputs(1899) <= b;
    layer0_outputs(1900) <= a or b;
    layer0_outputs(1901) <= not b;
    layer0_outputs(1902) <= not (a or b);
    layer0_outputs(1903) <= not a or b;
    layer0_outputs(1904) <= a or b;
    layer0_outputs(1905) <= a or b;
    layer0_outputs(1906) <= a or b;
    layer0_outputs(1907) <= a or b;
    layer0_outputs(1908) <= not (a xor b);
    layer0_outputs(1909) <= not (a or b);
    layer0_outputs(1910) <= a or b;
    layer0_outputs(1911) <= not (a or b);
    layer0_outputs(1912) <= not (a and b);
    layer0_outputs(1913) <= a or b;
    layer0_outputs(1914) <= '1';
    layer0_outputs(1915) <= not a;
    layer0_outputs(1916) <= '1';
    layer0_outputs(1917) <= a and not b;
    layer0_outputs(1918) <= not (a or b);
    layer0_outputs(1919) <= b;
    layer0_outputs(1920) <= a and not b;
    layer0_outputs(1921) <= not b;
    layer0_outputs(1922) <= not b or a;
    layer0_outputs(1923) <= not (a xor b);
    layer0_outputs(1924) <= a or b;
    layer0_outputs(1925) <= a and not b;
    layer0_outputs(1926) <= a or b;
    layer0_outputs(1927) <= b;
    layer0_outputs(1928) <= a and not b;
    layer0_outputs(1929) <= not a;
    layer0_outputs(1930) <= a;
    layer0_outputs(1931) <= not (a or b);
    layer0_outputs(1932) <= not b or a;
    layer0_outputs(1933) <= a xor b;
    layer0_outputs(1934) <= a or b;
    layer0_outputs(1935) <= a and b;
    layer0_outputs(1936) <= not a;
    layer0_outputs(1937) <= not a or b;
    layer0_outputs(1938) <= not (a xor b);
    layer0_outputs(1939) <= b;
    layer0_outputs(1940) <= b and not a;
    layer0_outputs(1941) <= a;
    layer0_outputs(1942) <= not b;
    layer0_outputs(1943) <= not b;
    layer0_outputs(1944) <= not a or b;
    layer0_outputs(1945) <= not a or b;
    layer0_outputs(1946) <= b;
    layer0_outputs(1947) <= a;
    layer0_outputs(1948) <= not a;
    layer0_outputs(1949) <= not (a xor b);
    layer0_outputs(1950) <= b;
    layer0_outputs(1951) <= a xor b;
    layer0_outputs(1952) <= not b;
    layer0_outputs(1953) <= a and not b;
    layer0_outputs(1954) <= a and not b;
    layer0_outputs(1955) <= not (a xor b);
    layer0_outputs(1956) <= not a or b;
    layer0_outputs(1957) <= not (a xor b);
    layer0_outputs(1958) <= a or b;
    layer0_outputs(1959) <= not b or a;
    layer0_outputs(1960) <= not (a or b);
    layer0_outputs(1961) <= not b;
    layer0_outputs(1962) <= a xor b;
    layer0_outputs(1963) <= not b;
    layer0_outputs(1964) <= not (a or b);
    layer0_outputs(1965) <= a;
    layer0_outputs(1966) <= not a or b;
    layer0_outputs(1967) <= a or b;
    layer0_outputs(1968) <= a or b;
    layer0_outputs(1969) <= a;
    layer0_outputs(1970) <= a or b;
    layer0_outputs(1971) <= not (a or b);
    layer0_outputs(1972) <= b;
    layer0_outputs(1973) <= not b;
    layer0_outputs(1974) <= not (a xor b);
    layer0_outputs(1975) <= '1';
    layer0_outputs(1976) <= not b or a;
    layer0_outputs(1977) <= not a or b;
    layer0_outputs(1978) <= not (a xor b);
    layer0_outputs(1979) <= not a or b;
    layer0_outputs(1980) <= not (a or b);
    layer0_outputs(1981) <= not a or b;
    layer0_outputs(1982) <= a or b;
    layer0_outputs(1983) <= not (a xor b);
    layer0_outputs(1984) <= not a;
    layer0_outputs(1985) <= b;
    layer0_outputs(1986) <= not (a or b);
    layer0_outputs(1987) <= a or b;
    layer0_outputs(1988) <= not a or b;
    layer0_outputs(1989) <= a or b;
    layer0_outputs(1990) <= not (a xor b);
    layer0_outputs(1991) <= not (a or b);
    layer0_outputs(1992) <= not b;
    layer0_outputs(1993) <= not (a or b);
    layer0_outputs(1994) <= not b;
    layer0_outputs(1995) <= not a or b;
    layer0_outputs(1996) <= a and not b;
    layer0_outputs(1997) <= '1';
    layer0_outputs(1998) <= a;
    layer0_outputs(1999) <= not b or a;
    layer0_outputs(2000) <= not (a and b);
    layer0_outputs(2001) <= not b or a;
    layer0_outputs(2002) <= not (a or b);
    layer0_outputs(2003) <= a and not b;
    layer0_outputs(2004) <= not a;
    layer0_outputs(2005) <= b and not a;
    layer0_outputs(2006) <= a or b;
    layer0_outputs(2007) <= a and b;
    layer0_outputs(2008) <= not a;
    layer0_outputs(2009) <= a;
    layer0_outputs(2010) <= a and b;
    layer0_outputs(2011) <= a xor b;
    layer0_outputs(2012) <= not (a xor b);
    layer0_outputs(2013) <= a or b;
    layer0_outputs(2014) <= not (a and b);
    layer0_outputs(2015) <= a and b;
    layer0_outputs(2016) <= not b or a;
    layer0_outputs(2017) <= not (a or b);
    layer0_outputs(2018) <= not (a xor b);
    layer0_outputs(2019) <= a or b;
    layer0_outputs(2020) <= b;
    layer0_outputs(2021) <= a;
    layer0_outputs(2022) <= a and not b;
    layer0_outputs(2023) <= b;
    layer0_outputs(2024) <= b;
    layer0_outputs(2025) <= a xor b;
    layer0_outputs(2026) <= a xor b;
    layer0_outputs(2027) <= not a or b;
    layer0_outputs(2028) <= not a or b;
    layer0_outputs(2029) <= a or b;
    layer0_outputs(2030) <= a xor b;
    layer0_outputs(2031) <= not b;
    layer0_outputs(2032) <= a and not b;
    layer0_outputs(2033) <= not (a xor b);
    layer0_outputs(2034) <= b;
    layer0_outputs(2035) <= a;
    layer0_outputs(2036) <= a or b;
    layer0_outputs(2037) <= not b or a;
    layer0_outputs(2038) <= a or b;
    layer0_outputs(2039) <= not (a or b);
    layer0_outputs(2040) <= not (a xor b);
    layer0_outputs(2041) <= not b or a;
    layer0_outputs(2042) <= a or b;
    layer0_outputs(2043) <= a xor b;
    layer0_outputs(2044) <= a;
    layer0_outputs(2045) <= not (a or b);
    layer0_outputs(2046) <= not (a or b);
    layer0_outputs(2047) <= b and not a;
    layer0_outputs(2048) <= b and not a;
    layer0_outputs(2049) <= not (a xor b);
    layer0_outputs(2050) <= a or b;
    layer0_outputs(2051) <= not (a xor b);
    layer0_outputs(2052) <= a and not b;
    layer0_outputs(2053) <= b;
    layer0_outputs(2054) <= not (a xor b);
    layer0_outputs(2055) <= not (a or b);
    layer0_outputs(2056) <= b and not a;
    layer0_outputs(2057) <= a or b;
    layer0_outputs(2058) <= not (a and b);
    layer0_outputs(2059) <= not (a and b);
    layer0_outputs(2060) <= not a;
    layer0_outputs(2061) <= a or b;
    layer0_outputs(2062) <= not (a xor b);
    layer0_outputs(2063) <= not a;
    layer0_outputs(2064) <= a or b;
    layer0_outputs(2065) <= not (a xor b);
    layer0_outputs(2066) <= not (a or b);
    layer0_outputs(2067) <= a and not b;
    layer0_outputs(2068) <= not a or b;
    layer0_outputs(2069) <= not b;
    layer0_outputs(2070) <= not (a xor b);
    layer0_outputs(2071) <= a or b;
    layer0_outputs(2072) <= not b;
    layer0_outputs(2073) <= a;
    layer0_outputs(2074) <= a;
    layer0_outputs(2075) <= a;
    layer0_outputs(2076) <= not a;
    layer0_outputs(2077) <= b and not a;
    layer0_outputs(2078) <= b;
    layer0_outputs(2079) <= not (a or b);
    layer0_outputs(2080) <= not (a xor b);
    layer0_outputs(2081) <= a or b;
    layer0_outputs(2082) <= not (a xor b);
    layer0_outputs(2083) <= not a;
    layer0_outputs(2084) <= a;
    layer0_outputs(2085) <= b;
    layer0_outputs(2086) <= a xor b;
    layer0_outputs(2087) <= b;
    layer0_outputs(2088) <= not a or b;
    layer0_outputs(2089) <= a or b;
    layer0_outputs(2090) <= not (a and b);
    layer0_outputs(2091) <= not (a xor b);
    layer0_outputs(2092) <= a or b;
    layer0_outputs(2093) <= not a;
    layer0_outputs(2094) <= a xor b;
    layer0_outputs(2095) <= a;
    layer0_outputs(2096) <= not (a or b);
    layer0_outputs(2097) <= not (a or b);
    layer0_outputs(2098) <= a xor b;
    layer0_outputs(2099) <= not a;
    layer0_outputs(2100) <= not b;
    layer0_outputs(2101) <= not a or b;
    layer0_outputs(2102) <= not (a or b);
    layer0_outputs(2103) <= not b;
    layer0_outputs(2104) <= not b or a;
    layer0_outputs(2105) <= a or b;
    layer0_outputs(2106) <= not b;
    layer0_outputs(2107) <= a and not b;
    layer0_outputs(2108) <= a and not b;
    layer0_outputs(2109) <= a xor b;
    layer0_outputs(2110) <= not (a xor b);
    layer0_outputs(2111) <= not (a xor b);
    layer0_outputs(2112) <= b;
    layer0_outputs(2113) <= a and b;
    layer0_outputs(2114) <= not b;
    layer0_outputs(2115) <= not (a or b);
    layer0_outputs(2116) <= a;
    layer0_outputs(2117) <= not b;
    layer0_outputs(2118) <= not (a or b);
    layer0_outputs(2119) <= a;
    layer0_outputs(2120) <= not (a or b);
    layer0_outputs(2121) <= not (a or b);
    layer0_outputs(2122) <= not (a xor b);
    layer0_outputs(2123) <= not b or a;
    layer0_outputs(2124) <= a or b;
    layer0_outputs(2125) <= not (a or b);
    layer0_outputs(2126) <= a xor b;
    layer0_outputs(2127) <= not a or b;
    layer0_outputs(2128) <= b;
    layer0_outputs(2129) <= a or b;
    layer0_outputs(2130) <= a or b;
    layer0_outputs(2131) <= not b or a;
    layer0_outputs(2132) <= not b;
    layer0_outputs(2133) <= not b or a;
    layer0_outputs(2134) <= a and not b;
    layer0_outputs(2135) <= not (a xor b);
    layer0_outputs(2136) <= not (a xor b);
    layer0_outputs(2137) <= not a;
    layer0_outputs(2138) <= not b or a;
    layer0_outputs(2139) <= not (a xor b);
    layer0_outputs(2140) <= a;
    layer0_outputs(2141) <= a xor b;
    layer0_outputs(2142) <= a or b;
    layer0_outputs(2143) <= a and not b;
    layer0_outputs(2144) <= a;
    layer0_outputs(2145) <= not b or a;
    layer0_outputs(2146) <= not b;
    layer0_outputs(2147) <= not a;
    layer0_outputs(2148) <= not a or b;
    layer0_outputs(2149) <= a xor b;
    layer0_outputs(2150) <= not a;
    layer0_outputs(2151) <= not b;
    layer0_outputs(2152) <= a and not b;
    layer0_outputs(2153) <= not (a xor b);
    layer0_outputs(2154) <= a;
    layer0_outputs(2155) <= not a or b;
    layer0_outputs(2156) <= not b;
    layer0_outputs(2157) <= not a;
    layer0_outputs(2158) <= not a;
    layer0_outputs(2159) <= b and not a;
    layer0_outputs(2160) <= a xor b;
    layer0_outputs(2161) <= not b or a;
    layer0_outputs(2162) <= '0';
    layer0_outputs(2163) <= not a or b;
    layer0_outputs(2164) <= not a;
    layer0_outputs(2165) <= not a or b;
    layer0_outputs(2166) <= not (a xor b);
    layer0_outputs(2167) <= a and not b;
    layer0_outputs(2168) <= a;
    layer0_outputs(2169) <= a;
    layer0_outputs(2170) <= a;
    layer0_outputs(2171) <= b and not a;
    layer0_outputs(2172) <= a;
    layer0_outputs(2173) <= not (a xor b);
    layer0_outputs(2174) <= b;
    layer0_outputs(2175) <= a and not b;
    layer0_outputs(2176) <= not (a and b);
    layer0_outputs(2177) <= b and not a;
    layer0_outputs(2178) <= a and not b;
    layer0_outputs(2179) <= '1';
    layer0_outputs(2180) <= a and b;
    layer0_outputs(2181) <= a xor b;
    layer0_outputs(2182) <= b;
    layer0_outputs(2183) <= not a or b;
    layer0_outputs(2184) <= b;
    layer0_outputs(2185) <= not a;
    layer0_outputs(2186) <= a xor b;
    layer0_outputs(2187) <= not (a or b);
    layer0_outputs(2188) <= not (a xor b);
    layer0_outputs(2189) <= not (a xor b);
    layer0_outputs(2190) <= a;
    layer0_outputs(2191) <= a or b;
    layer0_outputs(2192) <= not (a or b);
    layer0_outputs(2193) <= a or b;
    layer0_outputs(2194) <= a or b;
    layer0_outputs(2195) <= a and not b;
    layer0_outputs(2196) <= not a;
    layer0_outputs(2197) <= a xor b;
    layer0_outputs(2198) <= not a or b;
    layer0_outputs(2199) <= not (a or b);
    layer0_outputs(2200) <= not (a xor b);
    layer0_outputs(2201) <= a xor b;
    layer0_outputs(2202) <= not (a or b);
    layer0_outputs(2203) <= a and b;
    layer0_outputs(2204) <= a or b;
    layer0_outputs(2205) <= not b;
    layer0_outputs(2206) <= not (a xor b);
    layer0_outputs(2207) <= not (a xor b);
    layer0_outputs(2208) <= not a;
    layer0_outputs(2209) <= not (a xor b);
    layer0_outputs(2210) <= a and not b;
    layer0_outputs(2211) <= b;
    layer0_outputs(2212) <= a or b;
    layer0_outputs(2213) <= not b or a;
    layer0_outputs(2214) <= a or b;
    layer0_outputs(2215) <= not a;
    layer0_outputs(2216) <= b;
    layer0_outputs(2217) <= a and not b;
    layer0_outputs(2218) <= not a or b;
    layer0_outputs(2219) <= a xor b;
    layer0_outputs(2220) <= a;
    layer0_outputs(2221) <= not a or b;
    layer0_outputs(2222) <= a xor b;
    layer0_outputs(2223) <= not (a xor b);
    layer0_outputs(2224) <= not a;
    layer0_outputs(2225) <= a;
    layer0_outputs(2226) <= not a or b;
    layer0_outputs(2227) <= not a or b;
    layer0_outputs(2228) <= a and not b;
    layer0_outputs(2229) <= '1';
    layer0_outputs(2230) <= b;
    layer0_outputs(2231) <= not a;
    layer0_outputs(2232) <= b and not a;
    layer0_outputs(2233) <= not a or b;
    layer0_outputs(2234) <= a and not b;
    layer0_outputs(2235) <= b and not a;
    layer0_outputs(2236) <= not (a and b);
    layer0_outputs(2237) <= b and not a;
    layer0_outputs(2238) <= not (a or b);
    layer0_outputs(2239) <= a or b;
    layer0_outputs(2240) <= b and not a;
    layer0_outputs(2241) <= a;
    layer0_outputs(2242) <= b;
    layer0_outputs(2243) <= not (a xor b);
    layer0_outputs(2244) <= b;
    layer0_outputs(2245) <= a;
    layer0_outputs(2246) <= a or b;
    layer0_outputs(2247) <= a and not b;
    layer0_outputs(2248) <= not (a xor b);
    layer0_outputs(2249) <= not a or b;
    layer0_outputs(2250) <= a and not b;
    layer0_outputs(2251) <= not (a and b);
    layer0_outputs(2252) <= not (a and b);
    layer0_outputs(2253) <= b;
    layer0_outputs(2254) <= not (a and b);
    layer0_outputs(2255) <= not b or a;
    layer0_outputs(2256) <= not (a or b);
    layer0_outputs(2257) <= not a or b;
    layer0_outputs(2258) <= not (a or b);
    layer0_outputs(2259) <= a and not b;
    layer0_outputs(2260) <= not a;
    layer0_outputs(2261) <= not (a or b);
    layer0_outputs(2262) <= not (a or b);
    layer0_outputs(2263) <= not (a xor b);
    layer0_outputs(2264) <= a or b;
    layer0_outputs(2265) <= not (a xor b);
    layer0_outputs(2266) <= b;
    layer0_outputs(2267) <= not (a xor b);
    layer0_outputs(2268) <= not (a or b);
    layer0_outputs(2269) <= not a or b;
    layer0_outputs(2270) <= not b;
    layer0_outputs(2271) <= not b or a;
    layer0_outputs(2272) <= a or b;
    layer0_outputs(2273) <= a or b;
    layer0_outputs(2274) <= not a;
    layer0_outputs(2275) <= a and not b;
    layer0_outputs(2276) <= not b or a;
    layer0_outputs(2277) <= a xor b;
    layer0_outputs(2278) <= not (a or b);
    layer0_outputs(2279) <= a and not b;
    layer0_outputs(2280) <= b and not a;
    layer0_outputs(2281) <= not (a and b);
    layer0_outputs(2282) <= a;
    layer0_outputs(2283) <= not (a xor b);
    layer0_outputs(2284) <= b;
    layer0_outputs(2285) <= a or b;
    layer0_outputs(2286) <= a or b;
    layer0_outputs(2287) <= b;
    layer0_outputs(2288) <= a and not b;
    layer0_outputs(2289) <= a or b;
    layer0_outputs(2290) <= not a or b;
    layer0_outputs(2291) <= not (a xor b);
    layer0_outputs(2292) <= a or b;
    layer0_outputs(2293) <= not b or a;
    layer0_outputs(2294) <= a xor b;
    layer0_outputs(2295) <= a and not b;
    layer0_outputs(2296) <= a and not b;
    layer0_outputs(2297) <= b and not a;
    layer0_outputs(2298) <= a and not b;
    layer0_outputs(2299) <= not (a xor b);
    layer0_outputs(2300) <= a xor b;
    layer0_outputs(2301) <= a and not b;
    layer0_outputs(2302) <= b and not a;
    layer0_outputs(2303) <= not (a xor b);
    layer0_outputs(2304) <= b;
    layer0_outputs(2305) <= not (a or b);
    layer0_outputs(2306) <= a and not b;
    layer0_outputs(2307) <= a and b;
    layer0_outputs(2308) <= not b;
    layer0_outputs(2309) <= b;
    layer0_outputs(2310) <= not (a xor b);
    layer0_outputs(2311) <= not (a or b);
    layer0_outputs(2312) <= not (a xor b);
    layer0_outputs(2313) <= a xor b;
    layer0_outputs(2314) <= '0';
    layer0_outputs(2315) <= not (a or b);
    layer0_outputs(2316) <= b and not a;
    layer0_outputs(2317) <= not b;
    layer0_outputs(2318) <= not b or a;
    layer0_outputs(2319) <= a or b;
    layer0_outputs(2320) <= not b or a;
    layer0_outputs(2321) <= a and not b;
    layer0_outputs(2322) <= b;
    layer0_outputs(2323) <= '0';
    layer0_outputs(2324) <= a;
    layer0_outputs(2325) <= not (a xor b);
    layer0_outputs(2326) <= not b;
    layer0_outputs(2327) <= a xor b;
    layer0_outputs(2328) <= not b;
    layer0_outputs(2329) <= not (a xor b);
    layer0_outputs(2330) <= b and not a;
    layer0_outputs(2331) <= a and not b;
    layer0_outputs(2332) <= not b;
    layer0_outputs(2333) <= a or b;
    layer0_outputs(2334) <= b;
    layer0_outputs(2335) <= a and b;
    layer0_outputs(2336) <= b;
    layer0_outputs(2337) <= a and not b;
    layer0_outputs(2338) <= a xor b;
    layer0_outputs(2339) <= a and not b;
    layer0_outputs(2340) <= a and not b;
    layer0_outputs(2341) <= a or b;
    layer0_outputs(2342) <= a;
    layer0_outputs(2343) <= not (a or b);
    layer0_outputs(2344) <= a xor b;
    layer0_outputs(2345) <= not (a or b);
    layer0_outputs(2346) <= not (a or b);
    layer0_outputs(2347) <= a;
    layer0_outputs(2348) <= a or b;
    layer0_outputs(2349) <= a and not b;
    layer0_outputs(2350) <= a xor b;
    layer0_outputs(2351) <= not b;
    layer0_outputs(2352) <= not a;
    layer0_outputs(2353) <= not a;
    layer0_outputs(2354) <= not b;
    layer0_outputs(2355) <= a or b;
    layer0_outputs(2356) <= not b;
    layer0_outputs(2357) <= not (a xor b);
    layer0_outputs(2358) <= a;
    layer0_outputs(2359) <= b and not a;
    layer0_outputs(2360) <= not a;
    layer0_outputs(2361) <= not a;
    layer0_outputs(2362) <= a xor b;
    layer0_outputs(2363) <= not (a or b);
    layer0_outputs(2364) <= not (a or b);
    layer0_outputs(2365) <= not (a or b);
    layer0_outputs(2366) <= not a or b;
    layer0_outputs(2367) <= '0';
    layer0_outputs(2368) <= a xor b;
    layer0_outputs(2369) <= '0';
    layer0_outputs(2370) <= '1';
    layer0_outputs(2371) <= a and b;
    layer0_outputs(2372) <= not (a or b);
    layer0_outputs(2373) <= a xor b;
    layer0_outputs(2374) <= b and not a;
    layer0_outputs(2375) <= not a;
    layer0_outputs(2376) <= not a;
    layer0_outputs(2377) <= not a or b;
    layer0_outputs(2378) <= a xor b;
    layer0_outputs(2379) <= not a;
    layer0_outputs(2380) <= a or b;
    layer0_outputs(2381) <= a xor b;
    layer0_outputs(2382) <= b;
    layer0_outputs(2383) <= not a or b;
    layer0_outputs(2384) <= a or b;
    layer0_outputs(2385) <= not (a or b);
    layer0_outputs(2386) <= not (a or b);
    layer0_outputs(2387) <= not (a or b);
    layer0_outputs(2388) <= not b or a;
    layer0_outputs(2389) <= not b;
    layer0_outputs(2390) <= not b or a;
    layer0_outputs(2391) <= not a;
    layer0_outputs(2392) <= not (a xor b);
    layer0_outputs(2393) <= a xor b;
    layer0_outputs(2394) <= not b or a;
    layer0_outputs(2395) <= a and b;
    layer0_outputs(2396) <= a and b;
    layer0_outputs(2397) <= b and not a;
    layer0_outputs(2398) <= not (a or b);
    layer0_outputs(2399) <= b;
    layer0_outputs(2400) <= a and not b;
    layer0_outputs(2401) <= a or b;
    layer0_outputs(2402) <= '0';
    layer0_outputs(2403) <= not a;
    layer0_outputs(2404) <= b;
    layer0_outputs(2405) <= '0';
    layer0_outputs(2406) <= not (a or b);
    layer0_outputs(2407) <= not (a or b);
    layer0_outputs(2408) <= a or b;
    layer0_outputs(2409) <= b;
    layer0_outputs(2410) <= not (a or b);
    layer0_outputs(2411) <= not b;
    layer0_outputs(2412) <= not a;
    layer0_outputs(2413) <= not a or b;
    layer0_outputs(2414) <= not b or a;
    layer0_outputs(2415) <= not (a and b);
    layer0_outputs(2416) <= b and not a;
    layer0_outputs(2417) <= a or b;
    layer0_outputs(2418) <= not (a xor b);
    layer0_outputs(2419) <= a xor b;
    layer0_outputs(2420) <= not b or a;
    layer0_outputs(2421) <= not b or a;
    layer0_outputs(2422) <= a or b;
    layer0_outputs(2423) <= not (a xor b);
    layer0_outputs(2424) <= not (a or b);
    layer0_outputs(2425) <= not a;
    layer0_outputs(2426) <= not a;
    layer0_outputs(2427) <= b and not a;
    layer0_outputs(2428) <= a;
    layer0_outputs(2429) <= not (a or b);
    layer0_outputs(2430) <= a;
    layer0_outputs(2431) <= '1';
    layer0_outputs(2432) <= a and b;
    layer0_outputs(2433) <= b and not a;
    layer0_outputs(2434) <= not a or b;
    layer0_outputs(2435) <= not a;
    layer0_outputs(2436) <= a;
    layer0_outputs(2437) <= not (a or b);
    layer0_outputs(2438) <= '0';
    layer0_outputs(2439) <= not b or a;
    layer0_outputs(2440) <= a xor b;
    layer0_outputs(2441) <= a or b;
    layer0_outputs(2442) <= a and not b;
    layer0_outputs(2443) <= not b or a;
    layer0_outputs(2444) <= not a or b;
    layer0_outputs(2445) <= not (a xor b);
    layer0_outputs(2446) <= b;
    layer0_outputs(2447) <= b;
    layer0_outputs(2448) <= a and b;
    layer0_outputs(2449) <= a and not b;
    layer0_outputs(2450) <= not a or b;
    layer0_outputs(2451) <= a and not b;
    layer0_outputs(2452) <= a or b;
    layer0_outputs(2453) <= not a;
    layer0_outputs(2454) <= a xor b;
    layer0_outputs(2455) <= a xor b;
    layer0_outputs(2456) <= a;
    layer0_outputs(2457) <= not (a or b);
    layer0_outputs(2458) <= a or b;
    layer0_outputs(2459) <= a;
    layer0_outputs(2460) <= a or b;
    layer0_outputs(2461) <= not (a xor b);
    layer0_outputs(2462) <= '1';
    layer0_outputs(2463) <= b and not a;
    layer0_outputs(2464) <= a or b;
    layer0_outputs(2465) <= a;
    layer0_outputs(2466) <= a xor b;
    layer0_outputs(2467) <= a;
    layer0_outputs(2468) <= not b or a;
    layer0_outputs(2469) <= a;
    layer0_outputs(2470) <= a;
    layer0_outputs(2471) <= not b;
    layer0_outputs(2472) <= not a or b;
    layer0_outputs(2473) <= b and not a;
    layer0_outputs(2474) <= not a;
    layer0_outputs(2475) <= a and b;
    layer0_outputs(2476) <= not (a xor b);
    layer0_outputs(2477) <= not b or a;
    layer0_outputs(2478) <= a xor b;
    layer0_outputs(2479) <= a xor b;
    layer0_outputs(2480) <= not a;
    layer0_outputs(2481) <= b;
    layer0_outputs(2482) <= not b;
    layer0_outputs(2483) <= b and not a;
    layer0_outputs(2484) <= not b;
    layer0_outputs(2485) <= b;
    layer0_outputs(2486) <= not (a or b);
    layer0_outputs(2487) <= not a;
    layer0_outputs(2488) <= not a or b;
    layer0_outputs(2489) <= not b;
    layer0_outputs(2490) <= a xor b;
    layer0_outputs(2491) <= not a;
    layer0_outputs(2492) <= not b;
    layer0_outputs(2493) <= a xor b;
    layer0_outputs(2494) <= a;
    layer0_outputs(2495) <= not (a or b);
    layer0_outputs(2496) <= b;
    layer0_outputs(2497) <= b and not a;
    layer0_outputs(2498) <= b;
    layer0_outputs(2499) <= not a or b;
    layer0_outputs(2500) <= not (a xor b);
    layer0_outputs(2501) <= b and not a;
    layer0_outputs(2502) <= a xor b;
    layer0_outputs(2503) <= not (a or b);
    layer0_outputs(2504) <= a or b;
    layer0_outputs(2505) <= a;
    layer0_outputs(2506) <= a and not b;
    layer0_outputs(2507) <= b and not a;
    layer0_outputs(2508) <= a xor b;
    layer0_outputs(2509) <= not (a or b);
    layer0_outputs(2510) <= not b;
    layer0_outputs(2511) <= not (a or b);
    layer0_outputs(2512) <= not b or a;
    layer0_outputs(2513) <= not (a or b);
    layer0_outputs(2514) <= a or b;
    layer0_outputs(2515) <= '0';
    layer0_outputs(2516) <= not (a xor b);
    layer0_outputs(2517) <= b;
    layer0_outputs(2518) <= b and not a;
    layer0_outputs(2519) <= not (a xor b);
    layer0_outputs(2520) <= a or b;
    layer0_outputs(2521) <= not (a xor b);
    layer0_outputs(2522) <= b;
    layer0_outputs(2523) <= a;
    layer0_outputs(2524) <= not (a or b);
    layer0_outputs(2525) <= a or b;
    layer0_outputs(2526) <= not (a xor b);
    layer0_outputs(2527) <= not (a or b);
    layer0_outputs(2528) <= a xor b;
    layer0_outputs(2529) <= not b;
    layer0_outputs(2530) <= not (a xor b);
    layer0_outputs(2531) <= a xor b;
    layer0_outputs(2532) <= not b;
    layer0_outputs(2533) <= b;
    layer0_outputs(2534) <= a or b;
    layer0_outputs(2535) <= a and not b;
    layer0_outputs(2536) <= not (a or b);
    layer0_outputs(2537) <= b and not a;
    layer0_outputs(2538) <= a;
    layer0_outputs(2539) <= not a;
    layer0_outputs(2540) <= a;
    layer0_outputs(2541) <= not a;
    layer0_outputs(2542) <= not a;
    layer0_outputs(2543) <= not (a xor b);
    layer0_outputs(2544) <= not b or a;
    layer0_outputs(2545) <= not (a xor b);
    layer0_outputs(2546) <= a and not b;
    layer0_outputs(2547) <= a or b;
    layer0_outputs(2548) <= a and b;
    layer0_outputs(2549) <= not b or a;
    layer0_outputs(2550) <= not (a or b);
    layer0_outputs(2551) <= a or b;
    layer0_outputs(2552) <= not (a xor b);
    layer0_outputs(2553) <= a xor b;
    layer0_outputs(2554) <= not (a or b);
    layer0_outputs(2555) <= a;
    layer0_outputs(2556) <= a and b;
    layer0_outputs(2557) <= not b or a;
    layer0_outputs(2558) <= not (a xor b);
    layer0_outputs(2559) <= b and not a;
    layer0_outputs(2560) <= a or b;
    layer0_outputs(2561) <= a;
    layer0_outputs(2562) <= a or b;
    layer0_outputs(2563) <= not b;
    layer0_outputs(2564) <= not a or b;
    layer0_outputs(2565) <= a and b;
    layer0_outputs(2566) <= a;
    layer0_outputs(2567) <= not a;
    layer0_outputs(2568) <= b and not a;
    layer0_outputs(2569) <= a and not b;
    layer0_outputs(2570) <= a or b;
    layer0_outputs(2571) <= not a or b;
    layer0_outputs(2572) <= not (a or b);
    layer0_outputs(2573) <= a or b;
    layer0_outputs(2574) <= not a;
    layer0_outputs(2575) <= not b or a;
    layer0_outputs(2576) <= '0';
    layer0_outputs(2577) <= not a;
    layer0_outputs(2578) <= not b or a;
    layer0_outputs(2579) <= a;
    layer0_outputs(2580) <= a and not b;
    layer0_outputs(2581) <= a and not b;
    layer0_outputs(2582) <= not (a and b);
    layer0_outputs(2583) <= not a or b;
    layer0_outputs(2584) <= a and b;
    layer0_outputs(2585) <= a and b;
    layer0_outputs(2586) <= a or b;
    layer0_outputs(2587) <= a or b;
    layer0_outputs(2588) <= a;
    layer0_outputs(2589) <= not b;
    layer0_outputs(2590) <= not (a xor b);
    layer0_outputs(2591) <= a;
    layer0_outputs(2592) <= not (a or b);
    layer0_outputs(2593) <= a or b;
    layer0_outputs(2594) <= a and not b;
    layer0_outputs(2595) <= b and not a;
    layer0_outputs(2596) <= not a or b;
    layer0_outputs(2597) <= a or b;
    layer0_outputs(2598) <= not a or b;
    layer0_outputs(2599) <= not (a and b);
    layer0_outputs(2600) <= a;
    layer0_outputs(2601) <= not (a and b);
    layer0_outputs(2602) <= b;
    layer0_outputs(2603) <= b and not a;
    layer0_outputs(2604) <= not a;
    layer0_outputs(2605) <= not b or a;
    layer0_outputs(2606) <= not (a or b);
    layer0_outputs(2607) <= '0';
    layer0_outputs(2608) <= not (a xor b);
    layer0_outputs(2609) <= a or b;
    layer0_outputs(2610) <= not b;
    layer0_outputs(2611) <= not (a or b);
    layer0_outputs(2612) <= '0';
    layer0_outputs(2613) <= not (a xor b);
    layer0_outputs(2614) <= a xor b;
    layer0_outputs(2615) <= not b;
    layer0_outputs(2616) <= not (a and b);
    layer0_outputs(2617) <= not (a or b);
    layer0_outputs(2618) <= not (a xor b);
    layer0_outputs(2619) <= a or b;
    layer0_outputs(2620) <= not (a xor b);
    layer0_outputs(2621) <= b and not a;
    layer0_outputs(2622) <= a xor b;
    layer0_outputs(2623) <= not b or a;
    layer0_outputs(2624) <= not b or a;
    layer0_outputs(2625) <= not (a or b);
    layer0_outputs(2626) <= a or b;
    layer0_outputs(2627) <= '0';
    layer0_outputs(2628) <= not a or b;
    layer0_outputs(2629) <= a xor b;
    layer0_outputs(2630) <= a;
    layer0_outputs(2631) <= not (a or b);
    layer0_outputs(2632) <= a or b;
    layer0_outputs(2633) <= a;
    layer0_outputs(2634) <= not b;
    layer0_outputs(2635) <= not b;
    layer0_outputs(2636) <= b;
    layer0_outputs(2637) <= b;
    layer0_outputs(2638) <= not (a and b);
    layer0_outputs(2639) <= not b;
    layer0_outputs(2640) <= '1';
    layer0_outputs(2641) <= not a;
    layer0_outputs(2642) <= b and not a;
    layer0_outputs(2643) <= not b;
    layer0_outputs(2644) <= a or b;
    layer0_outputs(2645) <= a or b;
    layer0_outputs(2646) <= a xor b;
    layer0_outputs(2647) <= a and b;
    layer0_outputs(2648) <= a and b;
    layer0_outputs(2649) <= a and b;
    layer0_outputs(2650) <= a xor b;
    layer0_outputs(2651) <= a and b;
    layer0_outputs(2652) <= not a;
    layer0_outputs(2653) <= a xor b;
    layer0_outputs(2654) <= a;
    layer0_outputs(2655) <= not (a or b);
    layer0_outputs(2656) <= not b or a;
    layer0_outputs(2657) <= not (a or b);
    layer0_outputs(2658) <= not a or b;
    layer0_outputs(2659) <= not a or b;
    layer0_outputs(2660) <= a and not b;
    layer0_outputs(2661) <= not a;
    layer0_outputs(2662) <= b and not a;
    layer0_outputs(2663) <= b and not a;
    layer0_outputs(2664) <= a or b;
    layer0_outputs(2665) <= a;
    layer0_outputs(2666) <= '0';
    layer0_outputs(2667) <= not a or b;
    layer0_outputs(2668) <= a and not b;
    layer0_outputs(2669) <= not a or b;
    layer0_outputs(2670) <= not (a or b);
    layer0_outputs(2671) <= a xor b;
    layer0_outputs(2672) <= not (a and b);
    layer0_outputs(2673) <= not a;
    layer0_outputs(2674) <= not b;
    layer0_outputs(2675) <= a xor b;
    layer0_outputs(2676) <= not a;
    layer0_outputs(2677) <= not b or a;
    layer0_outputs(2678) <= not (a or b);
    layer0_outputs(2679) <= not b or a;
    layer0_outputs(2680) <= not b or a;
    layer0_outputs(2681) <= not (a xor b);
    layer0_outputs(2682) <= not (a and b);
    layer0_outputs(2683) <= not a;
    layer0_outputs(2684) <= '1';
    layer0_outputs(2685) <= not a or b;
    layer0_outputs(2686) <= not b or a;
    layer0_outputs(2687) <= b and not a;
    layer0_outputs(2688) <= a;
    layer0_outputs(2689) <= '1';
    layer0_outputs(2690) <= not (a or b);
    layer0_outputs(2691) <= not (a and b);
    layer0_outputs(2692) <= a and not b;
    layer0_outputs(2693) <= a xor b;
    layer0_outputs(2694) <= a or b;
    layer0_outputs(2695) <= b and not a;
    layer0_outputs(2696) <= not a or b;
    layer0_outputs(2697) <= '0';
    layer0_outputs(2698) <= a or b;
    layer0_outputs(2699) <= not a or b;
    layer0_outputs(2700) <= not b;
    layer0_outputs(2701) <= '0';
    layer0_outputs(2702) <= not a;
    layer0_outputs(2703) <= a xor b;
    layer0_outputs(2704) <= a or b;
    layer0_outputs(2705) <= a or b;
    layer0_outputs(2706) <= a or b;
    layer0_outputs(2707) <= not (a and b);
    layer0_outputs(2708) <= not (a or b);
    layer0_outputs(2709) <= a xor b;
    layer0_outputs(2710) <= not (a or b);
    layer0_outputs(2711) <= a or b;
    layer0_outputs(2712) <= not (a xor b);
    layer0_outputs(2713) <= not b or a;
    layer0_outputs(2714) <= not (a xor b);
    layer0_outputs(2715) <= b and not a;
    layer0_outputs(2716) <= not a;
    layer0_outputs(2717) <= not (a xor b);
    layer0_outputs(2718) <= not b or a;
    layer0_outputs(2719) <= a or b;
    layer0_outputs(2720) <= not a;
    layer0_outputs(2721) <= a or b;
    layer0_outputs(2722) <= a or b;
    layer0_outputs(2723) <= b and not a;
    layer0_outputs(2724) <= a;
    layer0_outputs(2725) <= a or b;
    layer0_outputs(2726) <= a and not b;
    layer0_outputs(2727) <= not (a xor b);
    layer0_outputs(2728) <= not a or b;
    layer0_outputs(2729) <= not a;
    layer0_outputs(2730) <= a xor b;
    layer0_outputs(2731) <= not b or a;
    layer0_outputs(2732) <= not b or a;
    layer0_outputs(2733) <= not a;
    layer0_outputs(2734) <= a or b;
    layer0_outputs(2735) <= a or b;
    layer0_outputs(2736) <= not (a or b);
    layer0_outputs(2737) <= a;
    layer0_outputs(2738) <= a or b;
    layer0_outputs(2739) <= a;
    layer0_outputs(2740) <= a or b;
    layer0_outputs(2741) <= a or b;
    layer0_outputs(2742) <= not a or b;
    layer0_outputs(2743) <= not (a or b);
    layer0_outputs(2744) <= not a;
    layer0_outputs(2745) <= b;
    layer0_outputs(2746) <= a or b;
    layer0_outputs(2747) <= a or b;
    layer0_outputs(2748) <= a xor b;
    layer0_outputs(2749) <= '0';
    layer0_outputs(2750) <= a xor b;
    layer0_outputs(2751) <= not b;
    layer0_outputs(2752) <= not b or a;
    layer0_outputs(2753) <= a and not b;
    layer0_outputs(2754) <= not (a xor b);
    layer0_outputs(2755) <= a or b;
    layer0_outputs(2756) <= a xor b;
    layer0_outputs(2757) <= b;
    layer0_outputs(2758) <= not a or b;
    layer0_outputs(2759) <= not (a or b);
    layer0_outputs(2760) <= a xor b;
    layer0_outputs(2761) <= not (a xor b);
    layer0_outputs(2762) <= not a or b;
    layer0_outputs(2763) <= not a or b;
    layer0_outputs(2764) <= a xor b;
    layer0_outputs(2765) <= a xor b;
    layer0_outputs(2766) <= not (a or b);
    layer0_outputs(2767) <= a or b;
    layer0_outputs(2768) <= a or b;
    layer0_outputs(2769) <= not (a xor b);
    layer0_outputs(2770) <= not (a or b);
    layer0_outputs(2771) <= not a or b;
    layer0_outputs(2772) <= not a or b;
    layer0_outputs(2773) <= not a;
    layer0_outputs(2774) <= a xor b;
    layer0_outputs(2775) <= not b;
    layer0_outputs(2776) <= '0';
    layer0_outputs(2777) <= a xor b;
    layer0_outputs(2778) <= not b;
    layer0_outputs(2779) <= not a;
    layer0_outputs(2780) <= not (a xor b);
    layer0_outputs(2781) <= a and not b;
    layer0_outputs(2782) <= a and b;
    layer0_outputs(2783) <= not a or b;
    layer0_outputs(2784) <= b and not a;
    layer0_outputs(2785) <= '1';
    layer0_outputs(2786) <= b and not a;
    layer0_outputs(2787) <= '1';
    layer0_outputs(2788) <= not a;
    layer0_outputs(2789) <= a or b;
    layer0_outputs(2790) <= a;
    layer0_outputs(2791) <= a;
    layer0_outputs(2792) <= a and not b;
    layer0_outputs(2793) <= not a;
    layer0_outputs(2794) <= a or b;
    layer0_outputs(2795) <= b;
    layer0_outputs(2796) <= not b or a;
    layer0_outputs(2797) <= not b or a;
    layer0_outputs(2798) <= not (a or b);
    layer0_outputs(2799) <= b;
    layer0_outputs(2800) <= not a;
    layer0_outputs(2801) <= not a;
    layer0_outputs(2802) <= a;
    layer0_outputs(2803) <= a or b;
    layer0_outputs(2804) <= '1';
    layer0_outputs(2805) <= not b or a;
    layer0_outputs(2806) <= a or b;
    layer0_outputs(2807) <= not (a and b);
    layer0_outputs(2808) <= a;
    layer0_outputs(2809) <= a;
    layer0_outputs(2810) <= a and not b;
    layer0_outputs(2811) <= not b;
    layer0_outputs(2812) <= a;
    layer0_outputs(2813) <= a and not b;
    layer0_outputs(2814) <= '1';
    layer0_outputs(2815) <= not (a or b);
    layer0_outputs(2816) <= not (a xor b);
    layer0_outputs(2817) <= a xor b;
    layer0_outputs(2818) <= a or b;
    layer0_outputs(2819) <= not b;
    layer0_outputs(2820) <= b;
    layer0_outputs(2821) <= not (a and b);
    layer0_outputs(2822) <= b and not a;
    layer0_outputs(2823) <= not b or a;
    layer0_outputs(2824) <= b;
    layer0_outputs(2825) <= a and not b;
    layer0_outputs(2826) <= not (a or b);
    layer0_outputs(2827) <= a;
    layer0_outputs(2828) <= a;
    layer0_outputs(2829) <= a;
    layer0_outputs(2830) <= not (a xor b);
    layer0_outputs(2831) <= a xor b;
    layer0_outputs(2832) <= not (a and b);
    layer0_outputs(2833) <= not b or a;
    layer0_outputs(2834) <= b and not a;
    layer0_outputs(2835) <= b;
    layer0_outputs(2836) <= not b;
    layer0_outputs(2837) <= a xor b;
    layer0_outputs(2838) <= b;
    layer0_outputs(2839) <= not (a or b);
    layer0_outputs(2840) <= not (a or b);
    layer0_outputs(2841) <= a and b;
    layer0_outputs(2842) <= a;
    layer0_outputs(2843) <= a xor b;
    layer0_outputs(2844) <= b;
    layer0_outputs(2845) <= a or b;
    layer0_outputs(2846) <= b and not a;
    layer0_outputs(2847) <= '1';
    layer0_outputs(2848) <= not (a or b);
    layer0_outputs(2849) <= '1';
    layer0_outputs(2850) <= a xor b;
    layer0_outputs(2851) <= not (a or b);
    layer0_outputs(2852) <= b;
    layer0_outputs(2853) <= not (a or b);
    layer0_outputs(2854) <= a xor b;
    layer0_outputs(2855) <= not b or a;
    layer0_outputs(2856) <= '0';
    layer0_outputs(2857) <= a or b;
    layer0_outputs(2858) <= not b;
    layer0_outputs(2859) <= b;
    layer0_outputs(2860) <= not a;
    layer0_outputs(2861) <= not a or b;
    layer0_outputs(2862) <= a and b;
    layer0_outputs(2863) <= a xor b;
    layer0_outputs(2864) <= a xor b;
    layer0_outputs(2865) <= a;
    layer0_outputs(2866) <= a;
    layer0_outputs(2867) <= '1';
    layer0_outputs(2868) <= not (a or b);
    layer0_outputs(2869) <= b;
    layer0_outputs(2870) <= not (a xor b);
    layer0_outputs(2871) <= not b or a;
    layer0_outputs(2872) <= not b;
    layer0_outputs(2873) <= not a;
    layer0_outputs(2874) <= not b or a;
    layer0_outputs(2875) <= b;
    layer0_outputs(2876) <= not a or b;
    layer0_outputs(2877) <= a and b;
    layer0_outputs(2878) <= not b;
    layer0_outputs(2879) <= not (a xor b);
    layer0_outputs(2880) <= a xor b;
    layer0_outputs(2881) <= a xor b;
    layer0_outputs(2882) <= b;
    layer0_outputs(2883) <= not a;
    layer0_outputs(2884) <= not b;
    layer0_outputs(2885) <= not (a xor b);
    layer0_outputs(2886) <= not a;
    layer0_outputs(2887) <= a xor b;
    layer0_outputs(2888) <= '0';
    layer0_outputs(2889) <= not (a xor b);
    layer0_outputs(2890) <= a or b;
    layer0_outputs(2891) <= a or b;
    layer0_outputs(2892) <= not (a or b);
    layer0_outputs(2893) <= not a;
    layer0_outputs(2894) <= a or b;
    layer0_outputs(2895) <= a;
    layer0_outputs(2896) <= not (a xor b);
    layer0_outputs(2897) <= a or b;
    layer0_outputs(2898) <= not b;
    layer0_outputs(2899) <= b and not a;
    layer0_outputs(2900) <= b;
    layer0_outputs(2901) <= a xor b;
    layer0_outputs(2902) <= a xor b;
    layer0_outputs(2903) <= not (a or b);
    layer0_outputs(2904) <= b;
    layer0_outputs(2905) <= b and not a;
    layer0_outputs(2906) <= '1';
    layer0_outputs(2907) <= b;
    layer0_outputs(2908) <= a or b;
    layer0_outputs(2909) <= b and not a;
    layer0_outputs(2910) <= a;
    layer0_outputs(2911) <= not (a xor b);
    layer0_outputs(2912) <= not (a or b);
    layer0_outputs(2913) <= not (a xor b);
    layer0_outputs(2914) <= not b or a;
    layer0_outputs(2915) <= not (a and b);
    layer0_outputs(2916) <= b;
    layer0_outputs(2917) <= a xor b;
    layer0_outputs(2918) <= not (a xor b);
    layer0_outputs(2919) <= a and b;
    layer0_outputs(2920) <= b and not a;
    layer0_outputs(2921) <= not a or b;
    layer0_outputs(2922) <= a xor b;
    layer0_outputs(2923) <= a and not b;
    layer0_outputs(2924) <= a xor b;
    layer0_outputs(2925) <= a or b;
    layer0_outputs(2926) <= a and b;
    layer0_outputs(2927) <= a;
    layer0_outputs(2928) <= b;
    layer0_outputs(2929) <= not a;
    layer0_outputs(2930) <= not (a or b);
    layer0_outputs(2931) <= not a or b;
    layer0_outputs(2932) <= a and b;
    layer0_outputs(2933) <= not b or a;
    layer0_outputs(2934) <= not (a or b);
    layer0_outputs(2935) <= not (a xor b);
    layer0_outputs(2936) <= a or b;
    layer0_outputs(2937) <= not (a xor b);
    layer0_outputs(2938) <= not a or b;
    layer0_outputs(2939) <= not (a xor b);
    layer0_outputs(2940) <= a or b;
    layer0_outputs(2941) <= a xor b;
    layer0_outputs(2942) <= a and not b;
    layer0_outputs(2943) <= a or b;
    layer0_outputs(2944) <= not a;
    layer0_outputs(2945) <= a xor b;
    layer0_outputs(2946) <= not a;
    layer0_outputs(2947) <= not (a and b);
    layer0_outputs(2948) <= b and not a;
    layer0_outputs(2949) <= not a;
    layer0_outputs(2950) <= a;
    layer0_outputs(2951) <= not a;
    layer0_outputs(2952) <= a;
    layer0_outputs(2953) <= not b or a;
    layer0_outputs(2954) <= a or b;
    layer0_outputs(2955) <= not a;
    layer0_outputs(2956) <= not b;
    layer0_outputs(2957) <= not (a and b);
    layer0_outputs(2958) <= not (a or b);
    layer0_outputs(2959) <= b and not a;
    layer0_outputs(2960) <= a;
    layer0_outputs(2961) <= a;
    layer0_outputs(2962) <= b;
    layer0_outputs(2963) <= not (a xor b);
    layer0_outputs(2964) <= '0';
    layer0_outputs(2965) <= not (a or b);
    layer0_outputs(2966) <= not (a or b);
    layer0_outputs(2967) <= not (a xor b);
    layer0_outputs(2968) <= not (a or b);
    layer0_outputs(2969) <= b;
    layer0_outputs(2970) <= not (a xor b);
    layer0_outputs(2971) <= b;
    layer0_outputs(2972) <= not a or b;
    layer0_outputs(2973) <= not b or a;
    layer0_outputs(2974) <= not b;
    layer0_outputs(2975) <= a and b;
    layer0_outputs(2976) <= not a;
    layer0_outputs(2977) <= a or b;
    layer0_outputs(2978) <= a;
    layer0_outputs(2979) <= b and not a;
    layer0_outputs(2980) <= not a or b;
    layer0_outputs(2981) <= '0';
    layer0_outputs(2982) <= not b;
    layer0_outputs(2983) <= a xor b;
    layer0_outputs(2984) <= a or b;
    layer0_outputs(2985) <= '1';
    layer0_outputs(2986) <= b and not a;
    layer0_outputs(2987) <= a xor b;
    layer0_outputs(2988) <= not (a or b);
    layer0_outputs(2989) <= a xor b;
    layer0_outputs(2990) <= a xor b;
    layer0_outputs(2991) <= '0';
    layer0_outputs(2992) <= b and not a;
    layer0_outputs(2993) <= not (a or b);
    layer0_outputs(2994) <= not (a and b);
    layer0_outputs(2995) <= not b or a;
    layer0_outputs(2996) <= a xor b;
    layer0_outputs(2997) <= b;
    layer0_outputs(2998) <= a or b;
    layer0_outputs(2999) <= not b or a;
    layer0_outputs(3000) <= not b;
    layer0_outputs(3001) <= not (a or b);
    layer0_outputs(3002) <= '1';
    layer0_outputs(3003) <= a or b;
    layer0_outputs(3004) <= a or b;
    layer0_outputs(3005) <= a;
    layer0_outputs(3006) <= not (a or b);
    layer0_outputs(3007) <= not b or a;
    layer0_outputs(3008) <= not b or a;
    layer0_outputs(3009) <= a and not b;
    layer0_outputs(3010) <= not (a or b);
    layer0_outputs(3011) <= a xor b;
    layer0_outputs(3012) <= a or b;
    layer0_outputs(3013) <= a and not b;
    layer0_outputs(3014) <= a xor b;
    layer0_outputs(3015) <= a or b;
    layer0_outputs(3016) <= not (a or b);
    layer0_outputs(3017) <= b;
    layer0_outputs(3018) <= not (a or b);
    layer0_outputs(3019) <= not a;
    layer0_outputs(3020) <= not b or a;
    layer0_outputs(3021) <= not b or a;
    layer0_outputs(3022) <= not a or b;
    layer0_outputs(3023) <= a;
    layer0_outputs(3024) <= a or b;
    layer0_outputs(3025) <= not b;
    layer0_outputs(3026) <= not b;
    layer0_outputs(3027) <= b;
    layer0_outputs(3028) <= a xor b;
    layer0_outputs(3029) <= not b or a;
    layer0_outputs(3030) <= not b or a;
    layer0_outputs(3031) <= not b;
    layer0_outputs(3032) <= b;
    layer0_outputs(3033) <= not (a xor b);
    layer0_outputs(3034) <= a;
    layer0_outputs(3035) <= not (a or b);
    layer0_outputs(3036) <= not b;
    layer0_outputs(3037) <= not a;
    layer0_outputs(3038) <= a;
    layer0_outputs(3039) <= b and not a;
    layer0_outputs(3040) <= a xor b;
    layer0_outputs(3041) <= b and not a;
    layer0_outputs(3042) <= a and not b;
    layer0_outputs(3043) <= not b or a;
    layer0_outputs(3044) <= '0';
    layer0_outputs(3045) <= not (a xor b);
    layer0_outputs(3046) <= not a or b;
    layer0_outputs(3047) <= not a;
    layer0_outputs(3048) <= not a;
    layer0_outputs(3049) <= a xor b;
    layer0_outputs(3050) <= not (a or b);
    layer0_outputs(3051) <= not (a xor b);
    layer0_outputs(3052) <= not (a xor b);
    layer0_outputs(3053) <= not a or b;
    layer0_outputs(3054) <= b;
    layer0_outputs(3055) <= not b;
    layer0_outputs(3056) <= not b or a;
    layer0_outputs(3057) <= b;
    layer0_outputs(3058) <= not b or a;
    layer0_outputs(3059) <= a and not b;
    layer0_outputs(3060) <= a xor b;
    layer0_outputs(3061) <= not (a or b);
    layer0_outputs(3062) <= b;
    layer0_outputs(3063) <= '1';
    layer0_outputs(3064) <= a and not b;
    layer0_outputs(3065) <= b and not a;
    layer0_outputs(3066) <= a;
    layer0_outputs(3067) <= a or b;
    layer0_outputs(3068) <= not (a or b);
    layer0_outputs(3069) <= b;
    layer0_outputs(3070) <= a or b;
    layer0_outputs(3071) <= b;
    layer0_outputs(3072) <= not (a or b);
    layer0_outputs(3073) <= b and not a;
    layer0_outputs(3074) <= not (a or b);
    layer0_outputs(3075) <= a;
    layer0_outputs(3076) <= b;
    layer0_outputs(3077) <= b and not a;
    layer0_outputs(3078) <= not b;
    layer0_outputs(3079) <= not b;
    layer0_outputs(3080) <= not a;
    layer0_outputs(3081) <= a and not b;
    layer0_outputs(3082) <= a or b;
    layer0_outputs(3083) <= b and not a;
    layer0_outputs(3084) <= not a or b;
    layer0_outputs(3085) <= '1';
    layer0_outputs(3086) <= not b or a;
    layer0_outputs(3087) <= a xor b;
    layer0_outputs(3088) <= b and not a;
    layer0_outputs(3089) <= not (a xor b);
    layer0_outputs(3090) <= b;
    layer0_outputs(3091) <= '1';
    layer0_outputs(3092) <= not (a or b);
    layer0_outputs(3093) <= a and b;
    layer0_outputs(3094) <= not (a or b);
    layer0_outputs(3095) <= not a;
    layer0_outputs(3096) <= b and not a;
    layer0_outputs(3097) <= not b;
    layer0_outputs(3098) <= b and not a;
    layer0_outputs(3099) <= '0';
    layer0_outputs(3100) <= not (a or b);
    layer0_outputs(3101) <= a xor b;
    layer0_outputs(3102) <= a and not b;
    layer0_outputs(3103) <= not (a or b);
    layer0_outputs(3104) <= a xor b;
    layer0_outputs(3105) <= a xor b;
    layer0_outputs(3106) <= a xor b;
    layer0_outputs(3107) <= not a;
    layer0_outputs(3108) <= a and not b;
    layer0_outputs(3109) <= not (a xor b);
    layer0_outputs(3110) <= not (a or b);
    layer0_outputs(3111) <= not (a or b);
    layer0_outputs(3112) <= a and b;
    layer0_outputs(3113) <= a or b;
    layer0_outputs(3114) <= not a or b;
    layer0_outputs(3115) <= not (a xor b);
    layer0_outputs(3116) <= a and not b;
    layer0_outputs(3117) <= not (a xor b);
    layer0_outputs(3118) <= a and b;
    layer0_outputs(3119) <= not a or b;
    layer0_outputs(3120) <= a or b;
    layer0_outputs(3121) <= b and not a;
    layer0_outputs(3122) <= a or b;
    layer0_outputs(3123) <= '0';
    layer0_outputs(3124) <= a xor b;
    layer0_outputs(3125) <= a or b;
    layer0_outputs(3126) <= a xor b;
    layer0_outputs(3127) <= a xor b;
    layer0_outputs(3128) <= not (a or b);
    layer0_outputs(3129) <= not (a or b);
    layer0_outputs(3130) <= a xor b;
    layer0_outputs(3131) <= not a;
    layer0_outputs(3132) <= not (a or b);
    layer0_outputs(3133) <= not (a xor b);
    layer0_outputs(3134) <= not (a or b);
    layer0_outputs(3135) <= not (a xor b);
    layer0_outputs(3136) <= not a or b;
    layer0_outputs(3137) <= not a;
    layer0_outputs(3138) <= not a;
    layer0_outputs(3139) <= '0';
    layer0_outputs(3140) <= a xor b;
    layer0_outputs(3141) <= not b;
    layer0_outputs(3142) <= not (a xor b);
    layer0_outputs(3143) <= a and not b;
    layer0_outputs(3144) <= not (a xor b);
    layer0_outputs(3145) <= a xor b;
    layer0_outputs(3146) <= a xor b;
    layer0_outputs(3147) <= not b;
    layer0_outputs(3148) <= a and b;
    layer0_outputs(3149) <= not a;
    layer0_outputs(3150) <= a and not b;
    layer0_outputs(3151) <= not (a or b);
    layer0_outputs(3152) <= not a or b;
    layer0_outputs(3153) <= a and not b;
    layer0_outputs(3154) <= not (a or b);
    layer0_outputs(3155) <= a xor b;
    layer0_outputs(3156) <= not a or b;
    layer0_outputs(3157) <= a and not b;
    layer0_outputs(3158) <= not (a or b);
    layer0_outputs(3159) <= not (a or b);
    layer0_outputs(3160) <= b;
    layer0_outputs(3161) <= a;
    layer0_outputs(3162) <= a or b;
    layer0_outputs(3163) <= b and not a;
    layer0_outputs(3164) <= not (a or b);
    layer0_outputs(3165) <= not a;
    layer0_outputs(3166) <= not (a xor b);
    layer0_outputs(3167) <= a xor b;
    layer0_outputs(3168) <= not (a xor b);
    layer0_outputs(3169) <= '0';
    layer0_outputs(3170) <= not b;
    layer0_outputs(3171) <= b;
    layer0_outputs(3172) <= not b or a;
    layer0_outputs(3173) <= a or b;
    layer0_outputs(3174) <= not (a or b);
    layer0_outputs(3175) <= not b or a;
    layer0_outputs(3176) <= not a;
    layer0_outputs(3177) <= not b or a;
    layer0_outputs(3178) <= a xor b;
    layer0_outputs(3179) <= a and not b;
    layer0_outputs(3180) <= not b;
    layer0_outputs(3181) <= a and b;
    layer0_outputs(3182) <= b;
    layer0_outputs(3183) <= a or b;
    layer0_outputs(3184) <= not (a and b);
    layer0_outputs(3185) <= b;
    layer0_outputs(3186) <= not (a or b);
    layer0_outputs(3187) <= not (a xor b);
    layer0_outputs(3188) <= a xor b;
    layer0_outputs(3189) <= a xor b;
    layer0_outputs(3190) <= not b or a;
    layer0_outputs(3191) <= not b;
    layer0_outputs(3192) <= a or b;
    layer0_outputs(3193) <= a xor b;
    layer0_outputs(3194) <= a and not b;
    layer0_outputs(3195) <= not b or a;
    layer0_outputs(3196) <= b;
    layer0_outputs(3197) <= not (a and b);
    layer0_outputs(3198) <= not a;
    layer0_outputs(3199) <= a and not b;
    layer0_outputs(3200) <= not b;
    layer0_outputs(3201) <= b and not a;
    layer0_outputs(3202) <= b and not a;
    layer0_outputs(3203) <= not (a xor b);
    layer0_outputs(3204) <= not (a or b);
    layer0_outputs(3205) <= a xor b;
    layer0_outputs(3206) <= a or b;
    layer0_outputs(3207) <= not a;
    layer0_outputs(3208) <= a or b;
    layer0_outputs(3209) <= not a;
    layer0_outputs(3210) <= a;
    layer0_outputs(3211) <= b and not a;
    layer0_outputs(3212) <= b and not a;
    layer0_outputs(3213) <= a and not b;
    layer0_outputs(3214) <= not (a and b);
    layer0_outputs(3215) <= not (a or b);
    layer0_outputs(3216) <= not a;
    layer0_outputs(3217) <= not a;
    layer0_outputs(3218) <= b;
    layer0_outputs(3219) <= a and not b;
    layer0_outputs(3220) <= not (a and b);
    layer0_outputs(3221) <= b and not a;
    layer0_outputs(3222) <= b;
    layer0_outputs(3223) <= a;
    layer0_outputs(3224) <= not (a or b);
    layer0_outputs(3225) <= not a;
    layer0_outputs(3226) <= not (a or b);
    layer0_outputs(3227) <= not a or b;
    layer0_outputs(3228) <= not b;
    layer0_outputs(3229) <= not (a or b);
    layer0_outputs(3230) <= not b;
    layer0_outputs(3231) <= not (a or b);
    layer0_outputs(3232) <= not b or a;
    layer0_outputs(3233) <= not a;
    layer0_outputs(3234) <= not b;
    layer0_outputs(3235) <= '1';
    layer0_outputs(3236) <= not (a or b);
    layer0_outputs(3237) <= a and b;
    layer0_outputs(3238) <= a or b;
    layer0_outputs(3239) <= a or b;
    layer0_outputs(3240) <= not a;
    layer0_outputs(3241) <= not a;
    layer0_outputs(3242) <= not a;
    layer0_outputs(3243) <= b and not a;
    layer0_outputs(3244) <= not (a or b);
    layer0_outputs(3245) <= '0';
    layer0_outputs(3246) <= a or b;
    layer0_outputs(3247) <= a;
    layer0_outputs(3248) <= b;
    layer0_outputs(3249) <= b;
    layer0_outputs(3250) <= '0';
    layer0_outputs(3251) <= not (a or b);
    layer0_outputs(3252) <= not b or a;
    layer0_outputs(3253) <= not b;
    layer0_outputs(3254) <= b and not a;
    layer0_outputs(3255) <= a;
    layer0_outputs(3256) <= '1';
    layer0_outputs(3257) <= a xor b;
    layer0_outputs(3258) <= b and not a;
    layer0_outputs(3259) <= not b;
    layer0_outputs(3260) <= a xor b;
    layer0_outputs(3261) <= not (a or b);
    layer0_outputs(3262) <= not (a xor b);
    layer0_outputs(3263) <= a or b;
    layer0_outputs(3264) <= not (a xor b);
    layer0_outputs(3265) <= not a;
    layer0_outputs(3266) <= not (a xor b);
    layer0_outputs(3267) <= a or b;
    layer0_outputs(3268) <= a or b;
    layer0_outputs(3269) <= not (a or b);
    layer0_outputs(3270) <= b;
    layer0_outputs(3271) <= a and b;
    layer0_outputs(3272) <= not (a xor b);
    layer0_outputs(3273) <= a xor b;
    layer0_outputs(3274) <= b;
    layer0_outputs(3275) <= a or b;
    layer0_outputs(3276) <= a xor b;
    layer0_outputs(3277) <= a xor b;
    layer0_outputs(3278) <= a;
    layer0_outputs(3279) <= '1';
    layer0_outputs(3280) <= not a;
    layer0_outputs(3281) <= not a;
    layer0_outputs(3282) <= not (a xor b);
    layer0_outputs(3283) <= not b;
    layer0_outputs(3284) <= a;
    layer0_outputs(3285) <= not b or a;
    layer0_outputs(3286) <= not (a or b);
    layer0_outputs(3287) <= a;
    layer0_outputs(3288) <= not (a and b);
    layer0_outputs(3289) <= b;
    layer0_outputs(3290) <= not a or b;
    layer0_outputs(3291) <= a or b;
    layer0_outputs(3292) <= b and not a;
    layer0_outputs(3293) <= a xor b;
    layer0_outputs(3294) <= a and not b;
    layer0_outputs(3295) <= not a or b;
    layer0_outputs(3296) <= b and not a;
    layer0_outputs(3297) <= not (a xor b);
    layer0_outputs(3298) <= not b or a;
    layer0_outputs(3299) <= a and not b;
    layer0_outputs(3300) <= a and not b;
    layer0_outputs(3301) <= not (a or b);
    layer0_outputs(3302) <= a;
    layer0_outputs(3303) <= not a or b;
    layer0_outputs(3304) <= a or b;
    layer0_outputs(3305) <= b;
    layer0_outputs(3306) <= not a;
    layer0_outputs(3307) <= a or b;
    layer0_outputs(3308) <= a xor b;
    layer0_outputs(3309) <= not (a or b);
    layer0_outputs(3310) <= a xor b;
    layer0_outputs(3311) <= a xor b;
    layer0_outputs(3312) <= a and not b;
    layer0_outputs(3313) <= not (a or b);
    layer0_outputs(3314) <= a xor b;
    layer0_outputs(3315) <= not b or a;
    layer0_outputs(3316) <= a xor b;
    layer0_outputs(3317) <= not b or a;
    layer0_outputs(3318) <= not (a or b);
    layer0_outputs(3319) <= '1';
    layer0_outputs(3320) <= a or b;
    layer0_outputs(3321) <= a or b;
    layer0_outputs(3322) <= a and not b;
    layer0_outputs(3323) <= not a or b;
    layer0_outputs(3324) <= b and not a;
    layer0_outputs(3325) <= a or b;
    layer0_outputs(3326) <= a xor b;
    layer0_outputs(3327) <= '0';
    layer0_outputs(3328) <= not a;
    layer0_outputs(3329) <= not (a xor b);
    layer0_outputs(3330) <= '1';
    layer0_outputs(3331) <= a or b;
    layer0_outputs(3332) <= not a or b;
    layer0_outputs(3333) <= b;
    layer0_outputs(3334) <= not (a or b);
    layer0_outputs(3335) <= not b;
    layer0_outputs(3336) <= not a;
    layer0_outputs(3337) <= not a;
    layer0_outputs(3338) <= not b or a;
    layer0_outputs(3339) <= b and not a;
    layer0_outputs(3340) <= a;
    layer0_outputs(3341) <= not a or b;
    layer0_outputs(3342) <= not b or a;
    layer0_outputs(3343) <= a xor b;
    layer0_outputs(3344) <= a;
    layer0_outputs(3345) <= not (a xor b);
    layer0_outputs(3346) <= not (a or b);
    layer0_outputs(3347) <= a or b;
    layer0_outputs(3348) <= a xor b;
    layer0_outputs(3349) <= b and not a;
    layer0_outputs(3350) <= a;
    layer0_outputs(3351) <= a and b;
    layer0_outputs(3352) <= b and not a;
    layer0_outputs(3353) <= a xor b;
    layer0_outputs(3354) <= a;
    layer0_outputs(3355) <= not (a or b);
    layer0_outputs(3356) <= not (a xor b);
    layer0_outputs(3357) <= b and not a;
    layer0_outputs(3358) <= not b or a;
    layer0_outputs(3359) <= b;
    layer0_outputs(3360) <= not b or a;
    layer0_outputs(3361) <= not b or a;
    layer0_outputs(3362) <= a or b;
    layer0_outputs(3363) <= a or b;
    layer0_outputs(3364) <= a or b;
    layer0_outputs(3365) <= not (a or b);
    layer0_outputs(3366) <= not a or b;
    layer0_outputs(3367) <= not b or a;
    layer0_outputs(3368) <= a;
    layer0_outputs(3369) <= a;
    layer0_outputs(3370) <= a or b;
    layer0_outputs(3371) <= not a;
    layer0_outputs(3372) <= not (a or b);
    layer0_outputs(3373) <= not (a xor b);
    layer0_outputs(3374) <= '0';
    layer0_outputs(3375) <= a or b;
    layer0_outputs(3376) <= not (a or b);
    layer0_outputs(3377) <= a and not b;
    layer0_outputs(3378) <= a xor b;
    layer0_outputs(3379) <= not a;
    layer0_outputs(3380) <= b and not a;
    layer0_outputs(3381) <= a or b;
    layer0_outputs(3382) <= b;
    layer0_outputs(3383) <= not (a or b);
    layer0_outputs(3384) <= not (a or b);
    layer0_outputs(3385) <= not b or a;
    layer0_outputs(3386) <= '1';
    layer0_outputs(3387) <= not (a and b);
    layer0_outputs(3388) <= not (a or b);
    layer0_outputs(3389) <= a or b;
    layer0_outputs(3390) <= '0';
    layer0_outputs(3391) <= b and not a;
    layer0_outputs(3392) <= not b;
    layer0_outputs(3393) <= a;
    layer0_outputs(3394) <= not b or a;
    layer0_outputs(3395) <= a and not b;
    layer0_outputs(3396) <= a or b;
    layer0_outputs(3397) <= a xor b;
    layer0_outputs(3398) <= a or b;
    layer0_outputs(3399) <= not a;
    layer0_outputs(3400) <= not b;
    layer0_outputs(3401) <= not a;
    layer0_outputs(3402) <= not b or a;
    layer0_outputs(3403) <= not b;
    layer0_outputs(3404) <= not a or b;
    layer0_outputs(3405) <= a or b;
    layer0_outputs(3406) <= a;
    layer0_outputs(3407) <= not (a and b);
    layer0_outputs(3408) <= '0';
    layer0_outputs(3409) <= not (a or b);
    layer0_outputs(3410) <= not a;
    layer0_outputs(3411) <= a or b;
    layer0_outputs(3412) <= not a;
    layer0_outputs(3413) <= a or b;
    layer0_outputs(3414) <= not (a or b);
    layer0_outputs(3415) <= not a or b;
    layer0_outputs(3416) <= not (a xor b);
    layer0_outputs(3417) <= a;
    layer0_outputs(3418) <= not (a or b);
    layer0_outputs(3419) <= a;
    layer0_outputs(3420) <= b;
    layer0_outputs(3421) <= a;
    layer0_outputs(3422) <= not a or b;
    layer0_outputs(3423) <= a or b;
    layer0_outputs(3424) <= a or b;
    layer0_outputs(3425) <= not (a or b);
    layer0_outputs(3426) <= b and not a;
    layer0_outputs(3427) <= '0';
    layer0_outputs(3428) <= not a or b;
    layer0_outputs(3429) <= a xor b;
    layer0_outputs(3430) <= not (a or b);
    layer0_outputs(3431) <= not a;
    layer0_outputs(3432) <= b;
    layer0_outputs(3433) <= a and not b;
    layer0_outputs(3434) <= a or b;
    layer0_outputs(3435) <= a and not b;
    layer0_outputs(3436) <= a xor b;
    layer0_outputs(3437) <= not a;
    layer0_outputs(3438) <= not (a xor b);
    layer0_outputs(3439) <= b;
    layer0_outputs(3440) <= not a or b;
    layer0_outputs(3441) <= a and b;
    layer0_outputs(3442) <= not (a xor b);
    layer0_outputs(3443) <= not a or b;
    layer0_outputs(3444) <= not (a or b);
    layer0_outputs(3445) <= b;
    layer0_outputs(3446) <= a and not b;
    layer0_outputs(3447) <= a and b;
    layer0_outputs(3448) <= not a or b;
    layer0_outputs(3449) <= not (a or b);
    layer0_outputs(3450) <= not (a and b);
    layer0_outputs(3451) <= not (a xor b);
    layer0_outputs(3452) <= a and b;
    layer0_outputs(3453) <= not (a xor b);
    layer0_outputs(3454) <= a and not b;
    layer0_outputs(3455) <= not b;
    layer0_outputs(3456) <= not (a or b);
    layer0_outputs(3457) <= b and not a;
    layer0_outputs(3458) <= a or b;
    layer0_outputs(3459) <= not a or b;
    layer0_outputs(3460) <= not a or b;
    layer0_outputs(3461) <= not (a or b);
    layer0_outputs(3462) <= a or b;
    layer0_outputs(3463) <= not (a and b);
    layer0_outputs(3464) <= not b;
    layer0_outputs(3465) <= not a or b;
    layer0_outputs(3466) <= b and not a;
    layer0_outputs(3467) <= not a or b;
    layer0_outputs(3468) <= b and not a;
    layer0_outputs(3469) <= '0';
    layer0_outputs(3470) <= b and not a;
    layer0_outputs(3471) <= not b;
    layer0_outputs(3472) <= '1';
    layer0_outputs(3473) <= '1';
    layer0_outputs(3474) <= a xor b;
    layer0_outputs(3475) <= '0';
    layer0_outputs(3476) <= not b;
    layer0_outputs(3477) <= '0';
    layer0_outputs(3478) <= not b;
    layer0_outputs(3479) <= not b;
    layer0_outputs(3480) <= not a;
    layer0_outputs(3481) <= not (a xor b);
    layer0_outputs(3482) <= not (a and b);
    layer0_outputs(3483) <= not a;
    layer0_outputs(3484) <= a or b;
    layer0_outputs(3485) <= not a;
    layer0_outputs(3486) <= not b;
    layer0_outputs(3487) <= a or b;
    layer0_outputs(3488) <= a and b;
    layer0_outputs(3489) <= b and not a;
    layer0_outputs(3490) <= a or b;
    layer0_outputs(3491) <= not a or b;
    layer0_outputs(3492) <= a or b;
    layer0_outputs(3493) <= not (a xor b);
    layer0_outputs(3494) <= b and not a;
    layer0_outputs(3495) <= not (a xor b);
    layer0_outputs(3496) <= not (a or b);
    layer0_outputs(3497) <= not (a or b);
    layer0_outputs(3498) <= not (a xor b);
    layer0_outputs(3499) <= a or b;
    layer0_outputs(3500) <= a or b;
    layer0_outputs(3501) <= not a;
    layer0_outputs(3502) <= b and not a;
    layer0_outputs(3503) <= a or b;
    layer0_outputs(3504) <= a or b;
    layer0_outputs(3505) <= not b;
    layer0_outputs(3506) <= not (a xor b);
    layer0_outputs(3507) <= '1';
    layer0_outputs(3508) <= not a;
    layer0_outputs(3509) <= a or b;
    layer0_outputs(3510) <= a xor b;
    layer0_outputs(3511) <= a and not b;
    layer0_outputs(3512) <= a or b;
    layer0_outputs(3513) <= a;
    layer0_outputs(3514) <= not (a xor b);
    layer0_outputs(3515) <= a;
    layer0_outputs(3516) <= a and b;
    layer0_outputs(3517) <= not a;
    layer0_outputs(3518) <= not a;
    layer0_outputs(3519) <= not a or b;
    layer0_outputs(3520) <= not b;
    layer0_outputs(3521) <= not a;
    layer0_outputs(3522) <= not a;
    layer0_outputs(3523) <= b and not a;
    layer0_outputs(3524) <= a or b;
    layer0_outputs(3525) <= a or b;
    layer0_outputs(3526) <= b and not a;
    layer0_outputs(3527) <= not (a or b);
    layer0_outputs(3528) <= a or b;
    layer0_outputs(3529) <= a xor b;
    layer0_outputs(3530) <= not b;
    layer0_outputs(3531) <= '0';
    layer0_outputs(3532) <= a or b;
    layer0_outputs(3533) <= not (a xor b);
    layer0_outputs(3534) <= a;
    layer0_outputs(3535) <= b and not a;
    layer0_outputs(3536) <= a or b;
    layer0_outputs(3537) <= not (a or b);
    layer0_outputs(3538) <= not (a or b);
    layer0_outputs(3539) <= a and not b;
    layer0_outputs(3540) <= '0';
    layer0_outputs(3541) <= not a or b;
    layer0_outputs(3542) <= a;
    layer0_outputs(3543) <= not b;
    layer0_outputs(3544) <= not b or a;
    layer0_outputs(3545) <= b and not a;
    layer0_outputs(3546) <= not a;
    layer0_outputs(3547) <= not (a xor b);
    layer0_outputs(3548) <= a;
    layer0_outputs(3549) <= not b or a;
    layer0_outputs(3550) <= a;
    layer0_outputs(3551) <= a and not b;
    layer0_outputs(3552) <= not a or b;
    layer0_outputs(3553) <= not (a and b);
    layer0_outputs(3554) <= not (a xor b);
    layer0_outputs(3555) <= a xor b;
    layer0_outputs(3556) <= b and not a;
    layer0_outputs(3557) <= a xor b;
    layer0_outputs(3558) <= a;
    layer0_outputs(3559) <= a or b;
    layer0_outputs(3560) <= not (a xor b);
    layer0_outputs(3561) <= not (a or b);
    layer0_outputs(3562) <= a xor b;
    layer0_outputs(3563) <= a and not b;
    layer0_outputs(3564) <= a or b;
    layer0_outputs(3565) <= b and not a;
    layer0_outputs(3566) <= '0';
    layer0_outputs(3567) <= not b;
    layer0_outputs(3568) <= not b;
    layer0_outputs(3569) <= a;
    layer0_outputs(3570) <= a and not b;
    layer0_outputs(3571) <= not (a and b);
    layer0_outputs(3572) <= a and not b;
    layer0_outputs(3573) <= a xor b;
    layer0_outputs(3574) <= a and not b;
    layer0_outputs(3575) <= not a;
    layer0_outputs(3576) <= not a or b;
    layer0_outputs(3577) <= a or b;
    layer0_outputs(3578) <= not (a xor b);
    layer0_outputs(3579) <= a xor b;
    layer0_outputs(3580) <= not b or a;
    layer0_outputs(3581) <= a;
    layer0_outputs(3582) <= b;
    layer0_outputs(3583) <= not a;
    layer0_outputs(3584) <= b;
    layer0_outputs(3585) <= not (a or b);
    layer0_outputs(3586) <= not (a and b);
    layer0_outputs(3587) <= a or b;
    layer0_outputs(3588) <= a;
    layer0_outputs(3589) <= a xor b;
    layer0_outputs(3590) <= not a;
    layer0_outputs(3591) <= not (a xor b);
    layer0_outputs(3592) <= b;
    layer0_outputs(3593) <= '0';
    layer0_outputs(3594) <= not b or a;
    layer0_outputs(3595) <= b;
    layer0_outputs(3596) <= a or b;
    layer0_outputs(3597) <= a or b;
    layer0_outputs(3598) <= not a or b;
    layer0_outputs(3599) <= a xor b;
    layer0_outputs(3600) <= b;
    layer0_outputs(3601) <= not (a xor b);
    layer0_outputs(3602) <= a or b;
    layer0_outputs(3603) <= not a or b;
    layer0_outputs(3604) <= not b or a;
    layer0_outputs(3605) <= a or b;
    layer0_outputs(3606) <= b;
    layer0_outputs(3607) <= a;
    layer0_outputs(3608) <= a;
    layer0_outputs(3609) <= b;
    layer0_outputs(3610) <= a;
    layer0_outputs(3611) <= a or b;
    layer0_outputs(3612) <= a or b;
    layer0_outputs(3613) <= b;
    layer0_outputs(3614) <= a or b;
    layer0_outputs(3615) <= not (a xor b);
    layer0_outputs(3616) <= b and not a;
    layer0_outputs(3617) <= not b or a;
    layer0_outputs(3618) <= b;
    layer0_outputs(3619) <= not (a and b);
    layer0_outputs(3620) <= not (a or b);
    layer0_outputs(3621) <= not a or b;
    layer0_outputs(3622) <= not (a xor b);
    layer0_outputs(3623) <= not a;
    layer0_outputs(3624) <= a;
    layer0_outputs(3625) <= b and not a;
    layer0_outputs(3626) <= not (a xor b);
    layer0_outputs(3627) <= a or b;
    layer0_outputs(3628) <= b and not a;
    layer0_outputs(3629) <= a xor b;
    layer0_outputs(3630) <= not b or a;
    layer0_outputs(3631) <= a and not b;
    layer0_outputs(3632) <= b and not a;
    layer0_outputs(3633) <= not b or a;
    layer0_outputs(3634) <= not b or a;
    layer0_outputs(3635) <= b;
    layer0_outputs(3636) <= b;
    layer0_outputs(3637) <= not a or b;
    layer0_outputs(3638) <= not (a or b);
    layer0_outputs(3639) <= a xor b;
    layer0_outputs(3640) <= a;
    layer0_outputs(3641) <= a;
    layer0_outputs(3642) <= a;
    layer0_outputs(3643) <= not (a xor b);
    layer0_outputs(3644) <= '0';
    layer0_outputs(3645) <= a or b;
    layer0_outputs(3646) <= not a;
    layer0_outputs(3647) <= not a;
    layer0_outputs(3648) <= not (a xor b);
    layer0_outputs(3649) <= not a or b;
    layer0_outputs(3650) <= not b;
    layer0_outputs(3651) <= '0';
    layer0_outputs(3652) <= a and b;
    layer0_outputs(3653) <= not (a or b);
    layer0_outputs(3654) <= a xor b;
    layer0_outputs(3655) <= a xor b;
    layer0_outputs(3656) <= a;
    layer0_outputs(3657) <= not (a xor b);
    layer0_outputs(3658) <= not b or a;
    layer0_outputs(3659) <= '0';
    layer0_outputs(3660) <= b;
    layer0_outputs(3661) <= not (a or b);
    layer0_outputs(3662) <= a or b;
    layer0_outputs(3663) <= '0';
    layer0_outputs(3664) <= a;
    layer0_outputs(3665) <= a;
    layer0_outputs(3666) <= not b;
    layer0_outputs(3667) <= not a;
    layer0_outputs(3668) <= b and not a;
    layer0_outputs(3669) <= not a or b;
    layer0_outputs(3670) <= a xor b;
    layer0_outputs(3671) <= not a;
    layer0_outputs(3672) <= not (a xor b);
    layer0_outputs(3673) <= not a;
    layer0_outputs(3674) <= b;
    layer0_outputs(3675) <= a xor b;
    layer0_outputs(3676) <= a and b;
    layer0_outputs(3677) <= not a or b;
    layer0_outputs(3678) <= '0';
    layer0_outputs(3679) <= a xor b;
    layer0_outputs(3680) <= not (a and b);
    layer0_outputs(3681) <= b and not a;
    layer0_outputs(3682) <= not b;
    layer0_outputs(3683) <= not b;
    layer0_outputs(3684) <= a xor b;
    layer0_outputs(3685) <= not a;
    layer0_outputs(3686) <= b and not a;
    layer0_outputs(3687) <= not a;
    layer0_outputs(3688) <= a or b;
    layer0_outputs(3689) <= not (a or b);
    layer0_outputs(3690) <= a and not b;
    layer0_outputs(3691) <= a xor b;
    layer0_outputs(3692) <= a;
    layer0_outputs(3693) <= not a or b;
    layer0_outputs(3694) <= a xor b;
    layer0_outputs(3695) <= not a or b;
    layer0_outputs(3696) <= a;
    layer0_outputs(3697) <= '1';
    layer0_outputs(3698) <= a xor b;
    layer0_outputs(3699) <= a and b;
    layer0_outputs(3700) <= b and not a;
    layer0_outputs(3701) <= not (a or b);
    layer0_outputs(3702) <= not b;
    layer0_outputs(3703) <= not b or a;
    layer0_outputs(3704) <= not (a or b);
    layer0_outputs(3705) <= a or b;
    layer0_outputs(3706) <= not a;
    layer0_outputs(3707) <= b and not a;
    layer0_outputs(3708) <= not a;
    layer0_outputs(3709) <= b;
    layer0_outputs(3710) <= not (a or b);
    layer0_outputs(3711) <= not a;
    layer0_outputs(3712) <= not a or b;
    layer0_outputs(3713) <= a or b;
    layer0_outputs(3714) <= a;
    layer0_outputs(3715) <= b;
    layer0_outputs(3716) <= b;
    layer0_outputs(3717) <= b and not a;
    layer0_outputs(3718) <= a or b;
    layer0_outputs(3719) <= not b or a;
    layer0_outputs(3720) <= not (a xor b);
    layer0_outputs(3721) <= not a or b;
    layer0_outputs(3722) <= a and not b;
    layer0_outputs(3723) <= not a;
    layer0_outputs(3724) <= not a or b;
    layer0_outputs(3725) <= a or b;
    layer0_outputs(3726) <= not a or b;
    layer0_outputs(3727) <= a;
    layer0_outputs(3728) <= not a;
    layer0_outputs(3729) <= b and not a;
    layer0_outputs(3730) <= not (a or b);
    layer0_outputs(3731) <= not (a or b);
    layer0_outputs(3732) <= not (a and b);
    layer0_outputs(3733) <= '0';
    layer0_outputs(3734) <= not a;
    layer0_outputs(3735) <= not (a or b);
    layer0_outputs(3736) <= b and not a;
    layer0_outputs(3737) <= b;
    layer0_outputs(3738) <= a and b;
    layer0_outputs(3739) <= not a or b;
    layer0_outputs(3740) <= a and not b;
    layer0_outputs(3741) <= not (a xor b);
    layer0_outputs(3742) <= b;
    layer0_outputs(3743) <= not a or b;
    layer0_outputs(3744) <= b and not a;
    layer0_outputs(3745) <= a and not b;
    layer0_outputs(3746) <= b;
    layer0_outputs(3747) <= a;
    layer0_outputs(3748) <= not a or b;
    layer0_outputs(3749) <= not a;
    layer0_outputs(3750) <= a;
    layer0_outputs(3751) <= not (a or b);
    layer0_outputs(3752) <= a;
    layer0_outputs(3753) <= not (a or b);
    layer0_outputs(3754) <= a;
    layer0_outputs(3755) <= not b;
    layer0_outputs(3756) <= not a or b;
    layer0_outputs(3757) <= not (a xor b);
    layer0_outputs(3758) <= not a;
    layer0_outputs(3759) <= '1';
    layer0_outputs(3760) <= not (a xor b);
    layer0_outputs(3761) <= b;
    layer0_outputs(3762) <= not (a or b);
    layer0_outputs(3763) <= a and not b;
    layer0_outputs(3764) <= not (a xor b);
    layer0_outputs(3765) <= not (a xor b);
    layer0_outputs(3766) <= a or b;
    layer0_outputs(3767) <= '0';
    layer0_outputs(3768) <= not (a xor b);
    layer0_outputs(3769) <= not a;
    layer0_outputs(3770) <= a or b;
    layer0_outputs(3771) <= not (a or b);
    layer0_outputs(3772) <= b;
    layer0_outputs(3773) <= not b;
    layer0_outputs(3774) <= a or b;
    layer0_outputs(3775) <= not (a xor b);
    layer0_outputs(3776) <= not (a xor b);
    layer0_outputs(3777) <= not (a or b);
    layer0_outputs(3778) <= a and b;
    layer0_outputs(3779) <= a and not b;
    layer0_outputs(3780) <= not a;
    layer0_outputs(3781) <= a xor b;
    layer0_outputs(3782) <= not (a xor b);
    layer0_outputs(3783) <= not (a or b);
    layer0_outputs(3784) <= a;
    layer0_outputs(3785) <= not (a and b);
    layer0_outputs(3786) <= a and b;
    layer0_outputs(3787) <= b and not a;
    layer0_outputs(3788) <= a xor b;
    layer0_outputs(3789) <= not a or b;
    layer0_outputs(3790) <= a or b;
    layer0_outputs(3791) <= b and not a;
    layer0_outputs(3792) <= not (a xor b);
    layer0_outputs(3793) <= not a;
    layer0_outputs(3794) <= a xor b;
    layer0_outputs(3795) <= not b;
    layer0_outputs(3796) <= not b or a;
    layer0_outputs(3797) <= not (a xor b);
    layer0_outputs(3798) <= a;
    layer0_outputs(3799) <= a xor b;
    layer0_outputs(3800) <= a xor b;
    layer0_outputs(3801) <= a or b;
    layer0_outputs(3802) <= a or b;
    layer0_outputs(3803) <= a and not b;
    layer0_outputs(3804) <= not b or a;
    layer0_outputs(3805) <= b;
    layer0_outputs(3806) <= a and b;
    layer0_outputs(3807) <= a;
    layer0_outputs(3808) <= not b;
    layer0_outputs(3809) <= a or b;
    layer0_outputs(3810) <= not a;
    layer0_outputs(3811) <= not (a xor b);
    layer0_outputs(3812) <= a and not b;
    layer0_outputs(3813) <= '0';
    layer0_outputs(3814) <= not (a xor b);
    layer0_outputs(3815) <= a or b;
    layer0_outputs(3816) <= a xor b;
    layer0_outputs(3817) <= not b;
    layer0_outputs(3818) <= a;
    layer0_outputs(3819) <= a and b;
    layer0_outputs(3820) <= a and b;
    layer0_outputs(3821) <= not b or a;
    layer0_outputs(3822) <= a or b;
    layer0_outputs(3823) <= not (a xor b);
    layer0_outputs(3824) <= a or b;
    layer0_outputs(3825) <= not (a or b);
    layer0_outputs(3826) <= not a;
    layer0_outputs(3827) <= not a or b;
    layer0_outputs(3828) <= not a or b;
    layer0_outputs(3829) <= not b;
    layer0_outputs(3830) <= b;
    layer0_outputs(3831) <= '0';
    layer0_outputs(3832) <= a and not b;
    layer0_outputs(3833) <= a xor b;
    layer0_outputs(3834) <= a xor b;
    layer0_outputs(3835) <= a and not b;
    layer0_outputs(3836) <= not b or a;
    layer0_outputs(3837) <= a or b;
    layer0_outputs(3838) <= a xor b;
    layer0_outputs(3839) <= not a;
    layer0_outputs(3840) <= not (a or b);
    layer0_outputs(3841) <= a xor b;
    layer0_outputs(3842) <= b;
    layer0_outputs(3843) <= a;
    layer0_outputs(3844) <= a;
    layer0_outputs(3845) <= not (a xor b);
    layer0_outputs(3846) <= a and b;
    layer0_outputs(3847) <= b;
    layer0_outputs(3848) <= not (a or b);
    layer0_outputs(3849) <= a and not b;
    layer0_outputs(3850) <= not b or a;
    layer0_outputs(3851) <= a or b;
    layer0_outputs(3852) <= not b;
    layer0_outputs(3853) <= a or b;
    layer0_outputs(3854) <= not (a or b);
    layer0_outputs(3855) <= a xor b;
    layer0_outputs(3856) <= a or b;
    layer0_outputs(3857) <= a or b;
    layer0_outputs(3858) <= b;
    layer0_outputs(3859) <= not b;
    layer0_outputs(3860) <= b and not a;
    layer0_outputs(3861) <= a or b;
    layer0_outputs(3862) <= '1';
    layer0_outputs(3863) <= a and not b;
    layer0_outputs(3864) <= not a or b;
    layer0_outputs(3865) <= a or b;
    layer0_outputs(3866) <= not a or b;
    layer0_outputs(3867) <= not a or b;
    layer0_outputs(3868) <= not (a or b);
    layer0_outputs(3869) <= not (a and b);
    layer0_outputs(3870) <= not a or b;
    layer0_outputs(3871) <= b and not a;
    layer0_outputs(3872) <= a xor b;
    layer0_outputs(3873) <= not a;
    layer0_outputs(3874) <= b;
    layer0_outputs(3875) <= not (a or b);
    layer0_outputs(3876) <= not b or a;
    layer0_outputs(3877) <= '0';
    layer0_outputs(3878) <= a and not b;
    layer0_outputs(3879) <= a and not b;
    layer0_outputs(3880) <= not (a and b);
    layer0_outputs(3881) <= not (a or b);
    layer0_outputs(3882) <= not (a or b);
    layer0_outputs(3883) <= a;
    layer0_outputs(3884) <= not b or a;
    layer0_outputs(3885) <= not (a or b);
    layer0_outputs(3886) <= '0';
    layer0_outputs(3887) <= a or b;
    layer0_outputs(3888) <= a;
    layer0_outputs(3889) <= not b or a;
    layer0_outputs(3890) <= not a;
    layer0_outputs(3891) <= not b or a;
    layer0_outputs(3892) <= not (a xor b);
    layer0_outputs(3893) <= a;
    layer0_outputs(3894) <= a and not b;
    layer0_outputs(3895) <= a or b;
    layer0_outputs(3896) <= not (a xor b);
    layer0_outputs(3897) <= not a or b;
    layer0_outputs(3898) <= not b or a;
    layer0_outputs(3899) <= b and not a;
    layer0_outputs(3900) <= a and not b;
    layer0_outputs(3901) <= a or b;
    layer0_outputs(3902) <= a and not b;
    layer0_outputs(3903) <= not (a or b);
    layer0_outputs(3904) <= not (a or b);
    layer0_outputs(3905) <= a;
    layer0_outputs(3906) <= b and not a;
    layer0_outputs(3907) <= a xor b;
    layer0_outputs(3908) <= a and not b;
    layer0_outputs(3909) <= a xor b;
    layer0_outputs(3910) <= a or b;
    layer0_outputs(3911) <= a xor b;
    layer0_outputs(3912) <= not (a or b);
    layer0_outputs(3913) <= not a or b;
    layer0_outputs(3914) <= a xor b;
    layer0_outputs(3915) <= b and not a;
    layer0_outputs(3916) <= b and not a;
    layer0_outputs(3917) <= not (a or b);
    layer0_outputs(3918) <= a;
    layer0_outputs(3919) <= not a or b;
    layer0_outputs(3920) <= a or b;
    layer0_outputs(3921) <= a and not b;
    layer0_outputs(3922) <= a;
    layer0_outputs(3923) <= b and not a;
    layer0_outputs(3924) <= a or b;
    layer0_outputs(3925) <= a xor b;
    layer0_outputs(3926) <= not (a or b);
    layer0_outputs(3927) <= b;
    layer0_outputs(3928) <= not (a and b);
    layer0_outputs(3929) <= a or b;
    layer0_outputs(3930) <= a or b;
    layer0_outputs(3931) <= not (a and b);
    layer0_outputs(3932) <= a and not b;
    layer0_outputs(3933) <= a or b;
    layer0_outputs(3934) <= b;
    layer0_outputs(3935) <= a xor b;
    layer0_outputs(3936) <= a;
    layer0_outputs(3937) <= not a or b;
    layer0_outputs(3938) <= not a;
    layer0_outputs(3939) <= b;
    layer0_outputs(3940) <= not b;
    layer0_outputs(3941) <= not a;
    layer0_outputs(3942) <= not b;
    layer0_outputs(3943) <= b and not a;
    layer0_outputs(3944) <= a or b;
    layer0_outputs(3945) <= a and not b;
    layer0_outputs(3946) <= a xor b;
    layer0_outputs(3947) <= not b or a;
    layer0_outputs(3948) <= a xor b;
    layer0_outputs(3949) <= a;
    layer0_outputs(3950) <= not b or a;
    layer0_outputs(3951) <= not (a or b);
    layer0_outputs(3952) <= not (a xor b);
    layer0_outputs(3953) <= not (a or b);
    layer0_outputs(3954) <= not b or a;
    layer0_outputs(3955) <= b;
    layer0_outputs(3956) <= b and not a;
    layer0_outputs(3957) <= not (a xor b);
    layer0_outputs(3958) <= '0';
    layer0_outputs(3959) <= not (a or b);
    layer0_outputs(3960) <= a;
    layer0_outputs(3961) <= not b;
    layer0_outputs(3962) <= not (a or b);
    layer0_outputs(3963) <= b and not a;
    layer0_outputs(3964) <= a and b;
    layer0_outputs(3965) <= a xor b;
    layer0_outputs(3966) <= not (a or b);
    layer0_outputs(3967) <= a or b;
    layer0_outputs(3968) <= b and not a;
    layer0_outputs(3969) <= not (a or b);
    layer0_outputs(3970) <= a or b;
    layer0_outputs(3971) <= b;
    layer0_outputs(3972) <= not a or b;
    layer0_outputs(3973) <= not a or b;
    layer0_outputs(3974) <= not (a or b);
    layer0_outputs(3975) <= a xor b;
    layer0_outputs(3976) <= not b or a;
    layer0_outputs(3977) <= not a;
    layer0_outputs(3978) <= b and not a;
    layer0_outputs(3979) <= not a or b;
    layer0_outputs(3980) <= not (a or b);
    layer0_outputs(3981) <= b and not a;
    layer0_outputs(3982) <= a xor b;
    layer0_outputs(3983) <= not a or b;
    layer0_outputs(3984) <= b and not a;
    layer0_outputs(3985) <= a and not b;
    layer0_outputs(3986) <= not a;
    layer0_outputs(3987) <= a;
    layer0_outputs(3988) <= a;
    layer0_outputs(3989) <= '0';
    layer0_outputs(3990) <= not (a or b);
    layer0_outputs(3991) <= not (a xor b);
    layer0_outputs(3992) <= a or b;
    layer0_outputs(3993) <= not a or b;
    layer0_outputs(3994) <= a and b;
    layer0_outputs(3995) <= a and b;
    layer0_outputs(3996) <= a and not b;
    layer0_outputs(3997) <= b and not a;
    layer0_outputs(3998) <= '0';
    layer0_outputs(3999) <= not a;
    layer0_outputs(4000) <= not (a xor b);
    layer0_outputs(4001) <= not a;
    layer0_outputs(4002) <= b and not a;
    layer0_outputs(4003) <= not b or a;
    layer0_outputs(4004) <= not (a or b);
    layer0_outputs(4005) <= not (a xor b);
    layer0_outputs(4006) <= '0';
    layer0_outputs(4007) <= a and not b;
    layer0_outputs(4008) <= not (a or b);
    layer0_outputs(4009) <= a xor b;
    layer0_outputs(4010) <= b and not a;
    layer0_outputs(4011) <= not a;
    layer0_outputs(4012) <= not b or a;
    layer0_outputs(4013) <= a xor b;
    layer0_outputs(4014) <= not b or a;
    layer0_outputs(4015) <= not (a and b);
    layer0_outputs(4016) <= a and b;
    layer0_outputs(4017) <= not (a xor b);
    layer0_outputs(4018) <= a xor b;
    layer0_outputs(4019) <= '1';
    layer0_outputs(4020) <= '0';
    layer0_outputs(4021) <= a or b;
    layer0_outputs(4022) <= not (a xor b);
    layer0_outputs(4023) <= not a;
    layer0_outputs(4024) <= a xor b;
    layer0_outputs(4025) <= not b;
    layer0_outputs(4026) <= not (a xor b);
    layer0_outputs(4027) <= b;
    layer0_outputs(4028) <= b;
    layer0_outputs(4029) <= not a;
    layer0_outputs(4030) <= not (a xor b);
    layer0_outputs(4031) <= a or b;
    layer0_outputs(4032) <= not a;
    layer0_outputs(4033) <= not b or a;
    layer0_outputs(4034) <= a or b;
    layer0_outputs(4035) <= a and not b;
    layer0_outputs(4036) <= a or b;
    layer0_outputs(4037) <= a or b;
    layer0_outputs(4038) <= not b;
    layer0_outputs(4039) <= not b or a;
    layer0_outputs(4040) <= not (a and b);
    layer0_outputs(4041) <= not b or a;
    layer0_outputs(4042) <= not b or a;
    layer0_outputs(4043) <= b;
    layer0_outputs(4044) <= a and b;
    layer0_outputs(4045) <= not a;
    layer0_outputs(4046) <= a or b;
    layer0_outputs(4047) <= a xor b;
    layer0_outputs(4048) <= not (a or b);
    layer0_outputs(4049) <= not (a or b);
    layer0_outputs(4050) <= not (a xor b);
    layer0_outputs(4051) <= b and not a;
    layer0_outputs(4052) <= not (a or b);
    layer0_outputs(4053) <= b and not a;
    layer0_outputs(4054) <= not (a xor b);
    layer0_outputs(4055) <= a or b;
    layer0_outputs(4056) <= not b or a;
    layer0_outputs(4057) <= b and not a;
    layer0_outputs(4058) <= not (a xor b);
    layer0_outputs(4059) <= not (a or b);
    layer0_outputs(4060) <= a or b;
    layer0_outputs(4061) <= not a or b;
    layer0_outputs(4062) <= b;
    layer0_outputs(4063) <= not b;
    layer0_outputs(4064) <= b;
    layer0_outputs(4065) <= not a;
    layer0_outputs(4066) <= not a;
    layer0_outputs(4067) <= b;
    layer0_outputs(4068) <= a xor b;
    layer0_outputs(4069) <= a;
    layer0_outputs(4070) <= not b or a;
    layer0_outputs(4071) <= a;
    layer0_outputs(4072) <= a xor b;
    layer0_outputs(4073) <= not (a xor b);
    layer0_outputs(4074) <= not (a xor b);
    layer0_outputs(4075) <= not b;
    layer0_outputs(4076) <= a and not b;
    layer0_outputs(4077) <= not (a or b);
    layer0_outputs(4078) <= a;
    layer0_outputs(4079) <= not (a or b);
    layer0_outputs(4080) <= not b or a;
    layer0_outputs(4081) <= not (a or b);
    layer0_outputs(4082) <= b;
    layer0_outputs(4083) <= not a;
    layer0_outputs(4084) <= not a;
    layer0_outputs(4085) <= not a or b;
    layer0_outputs(4086) <= a and b;
    layer0_outputs(4087) <= not (a xor b);
    layer0_outputs(4088) <= a xor b;
    layer0_outputs(4089) <= a or b;
    layer0_outputs(4090) <= '0';
    layer0_outputs(4091) <= b;
    layer0_outputs(4092) <= not a or b;
    layer0_outputs(4093) <= '0';
    layer0_outputs(4094) <= not b;
    layer0_outputs(4095) <= a and b;
    layer0_outputs(4096) <= not (a or b);
    layer0_outputs(4097) <= a xor b;
    layer0_outputs(4098) <= not (a or b);
    layer0_outputs(4099) <= b and not a;
    layer0_outputs(4100) <= not b or a;
    layer0_outputs(4101) <= a or b;
    layer0_outputs(4102) <= a or b;
    layer0_outputs(4103) <= a;
    layer0_outputs(4104) <= not (a xor b);
    layer0_outputs(4105) <= not (a or b);
    layer0_outputs(4106) <= not (a or b);
    layer0_outputs(4107) <= a xor b;
    layer0_outputs(4108) <= not (a and b);
    layer0_outputs(4109) <= not (a xor b);
    layer0_outputs(4110) <= not (a or b);
    layer0_outputs(4111) <= b;
    layer0_outputs(4112) <= not a;
    layer0_outputs(4113) <= not (a and b);
    layer0_outputs(4114) <= a;
    layer0_outputs(4115) <= '0';
    layer0_outputs(4116) <= not a or b;
    layer0_outputs(4117) <= a or b;
    layer0_outputs(4118) <= not a or b;
    layer0_outputs(4119) <= not (a or b);
    layer0_outputs(4120) <= a xor b;
    layer0_outputs(4121) <= '1';
    layer0_outputs(4122) <= a xor b;
    layer0_outputs(4123) <= a xor b;
    layer0_outputs(4124) <= b;
    layer0_outputs(4125) <= not (a or b);
    layer0_outputs(4126) <= not (a xor b);
    layer0_outputs(4127) <= not b;
    layer0_outputs(4128) <= not (a or b);
    layer0_outputs(4129) <= not (a xor b);
    layer0_outputs(4130) <= '1';
    layer0_outputs(4131) <= a;
    layer0_outputs(4132) <= a and not b;
    layer0_outputs(4133) <= not (a xor b);
    layer0_outputs(4134) <= not a or b;
    layer0_outputs(4135) <= a or b;
    layer0_outputs(4136) <= a xor b;
    layer0_outputs(4137) <= not b;
    layer0_outputs(4138) <= not a or b;
    layer0_outputs(4139) <= '1';
    layer0_outputs(4140) <= '1';
    layer0_outputs(4141) <= not b;
    layer0_outputs(4142) <= not a;
    layer0_outputs(4143) <= a or b;
    layer0_outputs(4144) <= not (a xor b);
    layer0_outputs(4145) <= a or b;
    layer0_outputs(4146) <= b and not a;
    layer0_outputs(4147) <= not (a and b);
    layer0_outputs(4148) <= not b;
    layer0_outputs(4149) <= not a;
    layer0_outputs(4150) <= b;
    layer0_outputs(4151) <= a;
    layer0_outputs(4152) <= not a or b;
    layer0_outputs(4153) <= not a;
    layer0_outputs(4154) <= not a;
    layer0_outputs(4155) <= a xor b;
    layer0_outputs(4156) <= a;
    layer0_outputs(4157) <= '1';
    layer0_outputs(4158) <= not b;
    layer0_outputs(4159) <= not a;
    layer0_outputs(4160) <= not (a or b);
    layer0_outputs(4161) <= b;
    layer0_outputs(4162) <= not a or b;
    layer0_outputs(4163) <= '0';
    layer0_outputs(4164) <= not a;
    layer0_outputs(4165) <= not (a xor b);
    layer0_outputs(4166) <= not (a or b);
    layer0_outputs(4167) <= not a;
    layer0_outputs(4168) <= a;
    layer0_outputs(4169) <= not (a or b);
    layer0_outputs(4170) <= a;
    layer0_outputs(4171) <= not b or a;
    layer0_outputs(4172) <= not (a and b);
    layer0_outputs(4173) <= '1';
    layer0_outputs(4174) <= a;
    layer0_outputs(4175) <= not b;
    layer0_outputs(4176) <= not a or b;
    layer0_outputs(4177) <= a or b;
    layer0_outputs(4178) <= a xor b;
    layer0_outputs(4179) <= not (a or b);
    layer0_outputs(4180) <= b;
    layer0_outputs(4181) <= not (a or b);
    layer0_outputs(4182) <= '0';
    layer0_outputs(4183) <= not b or a;
    layer0_outputs(4184) <= not (a xor b);
    layer0_outputs(4185) <= not a;
    layer0_outputs(4186) <= a or b;
    layer0_outputs(4187) <= a xor b;
    layer0_outputs(4188) <= not (a or b);
    layer0_outputs(4189) <= a or b;
    layer0_outputs(4190) <= not (a xor b);
    layer0_outputs(4191) <= not (a or b);
    layer0_outputs(4192) <= b and not a;
    layer0_outputs(4193) <= a or b;
    layer0_outputs(4194) <= not (a and b);
    layer0_outputs(4195) <= not a;
    layer0_outputs(4196) <= not b;
    layer0_outputs(4197) <= b and not a;
    layer0_outputs(4198) <= b;
    layer0_outputs(4199) <= not (a xor b);
    layer0_outputs(4200) <= a and b;
    layer0_outputs(4201) <= not (a or b);
    layer0_outputs(4202) <= a or b;
    layer0_outputs(4203) <= not a or b;
    layer0_outputs(4204) <= b and not a;
    layer0_outputs(4205) <= a and b;
    layer0_outputs(4206) <= a and not b;
    layer0_outputs(4207) <= not (a xor b);
    layer0_outputs(4208) <= not (a or b);
    layer0_outputs(4209) <= not (a or b);
    layer0_outputs(4210) <= b;
    layer0_outputs(4211) <= not (a xor b);
    layer0_outputs(4212) <= a;
    layer0_outputs(4213) <= b;
    layer0_outputs(4214) <= a or b;
    layer0_outputs(4215) <= a and not b;
    layer0_outputs(4216) <= not (a xor b);
    layer0_outputs(4217) <= b;
    layer0_outputs(4218) <= not (a or b);
    layer0_outputs(4219) <= a;
    layer0_outputs(4220) <= a or b;
    layer0_outputs(4221) <= not b or a;
    layer0_outputs(4222) <= not a or b;
    layer0_outputs(4223) <= a or b;
    layer0_outputs(4224) <= not b;
    layer0_outputs(4225) <= not b;
    layer0_outputs(4226) <= a;
    layer0_outputs(4227) <= a or b;
    layer0_outputs(4228) <= a xor b;
    layer0_outputs(4229) <= not b or a;
    layer0_outputs(4230) <= not (a or b);
    layer0_outputs(4231) <= not a;
    layer0_outputs(4232) <= '1';
    layer0_outputs(4233) <= a or b;
    layer0_outputs(4234) <= not b or a;
    layer0_outputs(4235) <= not a;
    layer0_outputs(4236) <= not a;
    layer0_outputs(4237) <= not b;
    layer0_outputs(4238) <= a or b;
    layer0_outputs(4239) <= a xor b;
    layer0_outputs(4240) <= a xor b;
    layer0_outputs(4241) <= not b;
    layer0_outputs(4242) <= not b;
    layer0_outputs(4243) <= b;
    layer0_outputs(4244) <= not (a xor b);
    layer0_outputs(4245) <= not b;
    layer0_outputs(4246) <= not a;
    layer0_outputs(4247) <= not (a or b);
    layer0_outputs(4248) <= a xor b;
    layer0_outputs(4249) <= not (a xor b);
    layer0_outputs(4250) <= a xor b;
    layer0_outputs(4251) <= b and not a;
    layer0_outputs(4252) <= not a or b;
    layer0_outputs(4253) <= a;
    layer0_outputs(4254) <= a or b;
    layer0_outputs(4255) <= not (a xor b);
    layer0_outputs(4256) <= a;
    layer0_outputs(4257) <= not a or b;
    layer0_outputs(4258) <= b;
    layer0_outputs(4259) <= not (a xor b);
    layer0_outputs(4260) <= b;
    layer0_outputs(4261) <= not a;
    layer0_outputs(4262) <= a or b;
    layer0_outputs(4263) <= not b or a;
    layer0_outputs(4264) <= a;
    layer0_outputs(4265) <= not a or b;
    layer0_outputs(4266) <= a xor b;
    layer0_outputs(4267) <= a;
    layer0_outputs(4268) <= not b;
    layer0_outputs(4269) <= b and not a;
    layer0_outputs(4270) <= not a;
    layer0_outputs(4271) <= not a;
    layer0_outputs(4272) <= b;
    layer0_outputs(4273) <= b;
    layer0_outputs(4274) <= a or b;
    layer0_outputs(4275) <= a;
    layer0_outputs(4276) <= a xor b;
    layer0_outputs(4277) <= not b or a;
    layer0_outputs(4278) <= not (a or b);
    layer0_outputs(4279) <= a or b;
    layer0_outputs(4280) <= not a;
    layer0_outputs(4281) <= not (a or b);
    layer0_outputs(4282) <= not (a xor b);
    layer0_outputs(4283) <= a or b;
    layer0_outputs(4284) <= a xor b;
    layer0_outputs(4285) <= not (a or b);
    layer0_outputs(4286) <= '0';
    layer0_outputs(4287) <= '1';
    layer0_outputs(4288) <= a xor b;
    layer0_outputs(4289) <= not b;
    layer0_outputs(4290) <= not (a xor b);
    layer0_outputs(4291) <= a;
    layer0_outputs(4292) <= not b or a;
    layer0_outputs(4293) <= a or b;
    layer0_outputs(4294) <= not b;
    layer0_outputs(4295) <= a and not b;
    layer0_outputs(4296) <= '1';
    layer0_outputs(4297) <= not (a or b);
    layer0_outputs(4298) <= a and not b;
    layer0_outputs(4299) <= a and not b;
    layer0_outputs(4300) <= a xor b;
    layer0_outputs(4301) <= not (a or b);
    layer0_outputs(4302) <= not (a xor b);
    layer0_outputs(4303) <= b and not a;
    layer0_outputs(4304) <= not a or b;
    layer0_outputs(4305) <= a or b;
    layer0_outputs(4306) <= not (a xor b);
    layer0_outputs(4307) <= not b;
    layer0_outputs(4308) <= a xor b;
    layer0_outputs(4309) <= a;
    layer0_outputs(4310) <= not a;
    layer0_outputs(4311) <= not b or a;
    layer0_outputs(4312) <= b and not a;
    layer0_outputs(4313) <= a xor b;
    layer0_outputs(4314) <= b and not a;
    layer0_outputs(4315) <= not (a or b);
    layer0_outputs(4316) <= not b or a;
    layer0_outputs(4317) <= '1';
    layer0_outputs(4318) <= b and not a;
    layer0_outputs(4319) <= not (a xor b);
    layer0_outputs(4320) <= not a;
    layer0_outputs(4321) <= not a or b;
    layer0_outputs(4322) <= b;
    layer0_outputs(4323) <= not (a or b);
    layer0_outputs(4324) <= a;
    layer0_outputs(4325) <= not a;
    layer0_outputs(4326) <= not (a or b);
    layer0_outputs(4327) <= not (a xor b);
    layer0_outputs(4328) <= a;
    layer0_outputs(4329) <= not b or a;
    layer0_outputs(4330) <= a;
    layer0_outputs(4331) <= '0';
    layer0_outputs(4332) <= a and not b;
    layer0_outputs(4333) <= b and not a;
    layer0_outputs(4334) <= a xor b;
    layer0_outputs(4335) <= not b;
    layer0_outputs(4336) <= a and not b;
    layer0_outputs(4337) <= not a;
    layer0_outputs(4338) <= not b or a;
    layer0_outputs(4339) <= not (a or b);
    layer0_outputs(4340) <= not a or b;
    layer0_outputs(4341) <= b and not a;
    layer0_outputs(4342) <= a and not b;
    layer0_outputs(4343) <= b and not a;
    layer0_outputs(4344) <= b;
    layer0_outputs(4345) <= a and not b;
    layer0_outputs(4346) <= a or b;
    layer0_outputs(4347) <= a xor b;
    layer0_outputs(4348) <= a or b;
    layer0_outputs(4349) <= a xor b;
    layer0_outputs(4350) <= not a or b;
    layer0_outputs(4351) <= b and not a;
    layer0_outputs(4352) <= a and b;
    layer0_outputs(4353) <= not a;
    layer0_outputs(4354) <= not (a xor b);
    layer0_outputs(4355) <= '0';
    layer0_outputs(4356) <= a xor b;
    layer0_outputs(4357) <= not (a or b);
    layer0_outputs(4358) <= b;
    layer0_outputs(4359) <= a;
    layer0_outputs(4360) <= not (a or b);
    layer0_outputs(4361) <= a;
    layer0_outputs(4362) <= not a or b;
    layer0_outputs(4363) <= a and not b;
    layer0_outputs(4364) <= a and not b;
    layer0_outputs(4365) <= not (a or b);
    layer0_outputs(4366) <= not b;
    layer0_outputs(4367) <= not a;
    layer0_outputs(4368) <= not (a or b);
    layer0_outputs(4369) <= '1';
    layer0_outputs(4370) <= not a;
    layer0_outputs(4371) <= '0';
    layer0_outputs(4372) <= not (a or b);
    layer0_outputs(4373) <= a or b;
    layer0_outputs(4374) <= not (a and b);
    layer0_outputs(4375) <= a and not b;
    layer0_outputs(4376) <= not a or b;
    layer0_outputs(4377) <= not b;
    layer0_outputs(4378) <= not a or b;
    layer0_outputs(4379) <= '1';
    layer0_outputs(4380) <= a or b;
    layer0_outputs(4381) <= not (a xor b);
    layer0_outputs(4382) <= a and b;
    layer0_outputs(4383) <= not b or a;
    layer0_outputs(4384) <= a xor b;
    layer0_outputs(4385) <= not b;
    layer0_outputs(4386) <= a xor b;
    layer0_outputs(4387) <= not a;
    layer0_outputs(4388) <= not b or a;
    layer0_outputs(4389) <= a and not b;
    layer0_outputs(4390) <= not (a or b);
    layer0_outputs(4391) <= '1';
    layer0_outputs(4392) <= a and not b;
    layer0_outputs(4393) <= b and not a;
    layer0_outputs(4394) <= b;
    layer0_outputs(4395) <= not (a and b);
    layer0_outputs(4396) <= a or b;
    layer0_outputs(4397) <= not (a xor b);
    layer0_outputs(4398) <= b and not a;
    layer0_outputs(4399) <= a and b;
    layer0_outputs(4400) <= b and not a;
    layer0_outputs(4401) <= '0';
    layer0_outputs(4402) <= a or b;
    layer0_outputs(4403) <= not a;
    layer0_outputs(4404) <= a or b;
    layer0_outputs(4405) <= not (a or b);
    layer0_outputs(4406) <= a or b;
    layer0_outputs(4407) <= not (a xor b);
    layer0_outputs(4408) <= b and not a;
    layer0_outputs(4409) <= a or b;
    layer0_outputs(4410) <= not (a xor b);
    layer0_outputs(4411) <= not (a or b);
    layer0_outputs(4412) <= not a;
    layer0_outputs(4413) <= not b;
    layer0_outputs(4414) <= not (a or b);
    layer0_outputs(4415) <= a;
    layer0_outputs(4416) <= a xor b;
    layer0_outputs(4417) <= not (a or b);
    layer0_outputs(4418) <= not (a or b);
    layer0_outputs(4419) <= not a;
    layer0_outputs(4420) <= not b;
    layer0_outputs(4421) <= a and not b;
    layer0_outputs(4422) <= a and not b;
    layer0_outputs(4423) <= not a;
    layer0_outputs(4424) <= not a or b;
    layer0_outputs(4425) <= not a;
    layer0_outputs(4426) <= a or b;
    layer0_outputs(4427) <= a and b;
    layer0_outputs(4428) <= not (a xor b);
    layer0_outputs(4429) <= not a;
    layer0_outputs(4430) <= b;
    layer0_outputs(4431) <= a and not b;
    layer0_outputs(4432) <= a;
    layer0_outputs(4433) <= a and not b;
    layer0_outputs(4434) <= not (a or b);
    layer0_outputs(4435) <= not (a and b);
    layer0_outputs(4436) <= not a;
    layer0_outputs(4437) <= not b;
    layer0_outputs(4438) <= a xor b;
    layer0_outputs(4439) <= not b;
    layer0_outputs(4440) <= not a;
    layer0_outputs(4441) <= a;
    layer0_outputs(4442) <= a and b;
    layer0_outputs(4443) <= not a or b;
    layer0_outputs(4444) <= a or b;
    layer0_outputs(4445) <= a and b;
    layer0_outputs(4446) <= a or b;
    layer0_outputs(4447) <= b and not a;
    layer0_outputs(4448) <= not b or a;
    layer0_outputs(4449) <= not (a or b);
    layer0_outputs(4450) <= not (a xor b);
    layer0_outputs(4451) <= not a or b;
    layer0_outputs(4452) <= not (a and b);
    layer0_outputs(4453) <= b and not a;
    layer0_outputs(4454) <= a or b;
    layer0_outputs(4455) <= not (a xor b);
    layer0_outputs(4456) <= a or b;
    layer0_outputs(4457) <= not b or a;
    layer0_outputs(4458) <= not b;
    layer0_outputs(4459) <= not (a xor b);
    layer0_outputs(4460) <= b;
    layer0_outputs(4461) <= not a;
    layer0_outputs(4462) <= a or b;
    layer0_outputs(4463) <= a or b;
    layer0_outputs(4464) <= a;
    layer0_outputs(4465) <= '1';
    layer0_outputs(4466) <= a xor b;
    layer0_outputs(4467) <= not a or b;
    layer0_outputs(4468) <= a or b;
    layer0_outputs(4469) <= a or b;
    layer0_outputs(4470) <= not b;
    layer0_outputs(4471) <= '0';
    layer0_outputs(4472) <= a xor b;
    layer0_outputs(4473) <= '1';
    layer0_outputs(4474) <= not (a xor b);
    layer0_outputs(4475) <= not b;
    layer0_outputs(4476) <= a;
    layer0_outputs(4477) <= a xor b;
    layer0_outputs(4478) <= not b;
    layer0_outputs(4479) <= a xor b;
    layer0_outputs(4480) <= not a or b;
    layer0_outputs(4481) <= a and b;
    layer0_outputs(4482) <= not (a and b);
    layer0_outputs(4483) <= not b or a;
    layer0_outputs(4484) <= a and not b;
    layer0_outputs(4485) <= a xor b;
    layer0_outputs(4486) <= not a;
    layer0_outputs(4487) <= a;
    layer0_outputs(4488) <= not b or a;
    layer0_outputs(4489) <= not (a or b);
    layer0_outputs(4490) <= b and not a;
    layer0_outputs(4491) <= not (a and b);
    layer0_outputs(4492) <= b;
    layer0_outputs(4493) <= not a;
    layer0_outputs(4494) <= b;
    layer0_outputs(4495) <= not b or a;
    layer0_outputs(4496) <= a xor b;
    layer0_outputs(4497) <= not a or b;
    layer0_outputs(4498) <= a or b;
    layer0_outputs(4499) <= not (a or b);
    layer0_outputs(4500) <= not a;
    layer0_outputs(4501) <= b;
    layer0_outputs(4502) <= not (a xor b);
    layer0_outputs(4503) <= a or b;
    layer0_outputs(4504) <= b;
    layer0_outputs(4505) <= a and not b;
    layer0_outputs(4506) <= not a or b;
    layer0_outputs(4507) <= a xor b;
    layer0_outputs(4508) <= '0';
    layer0_outputs(4509) <= a xor b;
    layer0_outputs(4510) <= not a or b;
    layer0_outputs(4511) <= a and not b;
    layer0_outputs(4512) <= a or b;
    layer0_outputs(4513) <= b;
    layer0_outputs(4514) <= not a;
    layer0_outputs(4515) <= a and not b;
    layer0_outputs(4516) <= '1';
    layer0_outputs(4517) <= a or b;
    layer0_outputs(4518) <= not a or b;
    layer0_outputs(4519) <= not a;
    layer0_outputs(4520) <= b and not a;
    layer0_outputs(4521) <= b and not a;
    layer0_outputs(4522) <= b and not a;
    layer0_outputs(4523) <= b and not a;
    layer0_outputs(4524) <= b;
    layer0_outputs(4525) <= not (a xor b);
    layer0_outputs(4526) <= not (a and b);
    layer0_outputs(4527) <= a or b;
    layer0_outputs(4528) <= a or b;
    layer0_outputs(4529) <= a or b;
    layer0_outputs(4530) <= not (a xor b);
    layer0_outputs(4531) <= a xor b;
    layer0_outputs(4532) <= a or b;
    layer0_outputs(4533) <= not (a or b);
    layer0_outputs(4534) <= '0';
    layer0_outputs(4535) <= a xor b;
    layer0_outputs(4536) <= not a or b;
    layer0_outputs(4537) <= not b;
    layer0_outputs(4538) <= a and not b;
    layer0_outputs(4539) <= a xor b;
    layer0_outputs(4540) <= a or b;
    layer0_outputs(4541) <= a or b;
    layer0_outputs(4542) <= not (a xor b);
    layer0_outputs(4543) <= not (a xor b);
    layer0_outputs(4544) <= a;
    layer0_outputs(4545) <= a xor b;
    layer0_outputs(4546) <= not (a xor b);
    layer0_outputs(4547) <= not (a xor b);
    layer0_outputs(4548) <= not (a or b);
    layer0_outputs(4549) <= a xor b;
    layer0_outputs(4550) <= not (a xor b);
    layer0_outputs(4551) <= a xor b;
    layer0_outputs(4552) <= a and not b;
    layer0_outputs(4553) <= a or b;
    layer0_outputs(4554) <= not b or a;
    layer0_outputs(4555) <= not (a xor b);
    layer0_outputs(4556) <= not (a xor b);
    layer0_outputs(4557) <= not (a and b);
    layer0_outputs(4558) <= b;
    layer0_outputs(4559) <= a and not b;
    layer0_outputs(4560) <= not a;
    layer0_outputs(4561) <= not (a xor b);
    layer0_outputs(4562) <= a xor b;
    layer0_outputs(4563) <= a;
    layer0_outputs(4564) <= a;
    layer0_outputs(4565) <= not a;
    layer0_outputs(4566) <= '1';
    layer0_outputs(4567) <= b and not a;
    layer0_outputs(4568) <= not a or b;
    layer0_outputs(4569) <= not (a or b);
    layer0_outputs(4570) <= a xor b;
    layer0_outputs(4571) <= not (a or b);
    layer0_outputs(4572) <= a and b;
    layer0_outputs(4573) <= a and b;
    layer0_outputs(4574) <= not b;
    layer0_outputs(4575) <= a xor b;
    layer0_outputs(4576) <= a or b;
    layer0_outputs(4577) <= a and b;
    layer0_outputs(4578) <= not (a and b);
    layer0_outputs(4579) <= a;
    layer0_outputs(4580) <= not (a and b);
    layer0_outputs(4581) <= not b;
    layer0_outputs(4582) <= b;
    layer0_outputs(4583) <= '1';
    layer0_outputs(4584) <= not (a or b);
    layer0_outputs(4585) <= '1';
    layer0_outputs(4586) <= b and not a;
    layer0_outputs(4587) <= a and not b;
    layer0_outputs(4588) <= b;
    layer0_outputs(4589) <= not (a xor b);
    layer0_outputs(4590) <= not (a or b);
    layer0_outputs(4591) <= a xor b;
    layer0_outputs(4592) <= not (a or b);
    layer0_outputs(4593) <= not b;
    layer0_outputs(4594) <= not a;
    layer0_outputs(4595) <= a or b;
    layer0_outputs(4596) <= a xor b;
    layer0_outputs(4597) <= not (a and b);
    layer0_outputs(4598) <= a or b;
    layer0_outputs(4599) <= '1';
    layer0_outputs(4600) <= a;
    layer0_outputs(4601) <= a or b;
    layer0_outputs(4602) <= not a or b;
    layer0_outputs(4603) <= not (a xor b);
    layer0_outputs(4604) <= a xor b;
    layer0_outputs(4605) <= not (a xor b);
    layer0_outputs(4606) <= b;
    layer0_outputs(4607) <= not a;
    layer0_outputs(4608) <= a and b;
    layer0_outputs(4609) <= not b;
    layer0_outputs(4610) <= b;
    layer0_outputs(4611) <= a;
    layer0_outputs(4612) <= not b or a;
    layer0_outputs(4613) <= not b;
    layer0_outputs(4614) <= b;
    layer0_outputs(4615) <= b and not a;
    layer0_outputs(4616) <= not (a and b);
    layer0_outputs(4617) <= b;
    layer0_outputs(4618) <= not (a or b);
    layer0_outputs(4619) <= not (a xor b);
    layer0_outputs(4620) <= not a;
    layer0_outputs(4621) <= not (a or b);
    layer0_outputs(4622) <= not b;
    layer0_outputs(4623) <= not (a and b);
    layer0_outputs(4624) <= b;
    layer0_outputs(4625) <= a and not b;
    layer0_outputs(4626) <= not a or b;
    layer0_outputs(4627) <= b and not a;
    layer0_outputs(4628) <= a or b;
    layer0_outputs(4629) <= not b or a;
    layer0_outputs(4630) <= not a or b;
    layer0_outputs(4631) <= a or b;
    layer0_outputs(4632) <= a or b;
    layer0_outputs(4633) <= a xor b;
    layer0_outputs(4634) <= not a or b;
    layer0_outputs(4635) <= not (a or b);
    layer0_outputs(4636) <= a or b;
    layer0_outputs(4637) <= a or b;
    layer0_outputs(4638) <= b and not a;
    layer0_outputs(4639) <= not b;
    layer0_outputs(4640) <= not a;
    layer0_outputs(4641) <= not b;
    layer0_outputs(4642) <= not (a or b);
    layer0_outputs(4643) <= not b or a;
    layer0_outputs(4644) <= not a;
    layer0_outputs(4645) <= not b or a;
    layer0_outputs(4646) <= a or b;
    layer0_outputs(4647) <= '1';
    layer0_outputs(4648) <= not a;
    layer0_outputs(4649) <= b;
    layer0_outputs(4650) <= b;
    layer0_outputs(4651) <= a xor b;
    layer0_outputs(4652) <= not (a or b);
    layer0_outputs(4653) <= not b;
    layer0_outputs(4654) <= not (a or b);
    layer0_outputs(4655) <= b and not a;
    layer0_outputs(4656) <= not (a or b);
    layer0_outputs(4657) <= a xor b;
    layer0_outputs(4658) <= b and not a;
    layer0_outputs(4659) <= a and b;
    layer0_outputs(4660) <= b and not a;
    layer0_outputs(4661) <= b;
    layer0_outputs(4662) <= not (a or b);
    layer0_outputs(4663) <= not (a xor b);
    layer0_outputs(4664) <= a and not b;
    layer0_outputs(4665) <= a xor b;
    layer0_outputs(4666) <= a or b;
    layer0_outputs(4667) <= not b or a;
    layer0_outputs(4668) <= not (a or b);
    layer0_outputs(4669) <= not (a or b);
    layer0_outputs(4670) <= not b or a;
    layer0_outputs(4671) <= not b or a;
    layer0_outputs(4672) <= not (a and b);
    layer0_outputs(4673) <= not (a or b);
    layer0_outputs(4674) <= not b or a;
    layer0_outputs(4675) <= a or b;
    layer0_outputs(4676) <= not (a xor b);
    layer0_outputs(4677) <= not b;
    layer0_outputs(4678) <= not a;
    layer0_outputs(4679) <= a xor b;
    layer0_outputs(4680) <= a and not b;
    layer0_outputs(4681) <= a;
    layer0_outputs(4682) <= a;
    layer0_outputs(4683) <= a;
    layer0_outputs(4684) <= not b or a;
    layer0_outputs(4685) <= not (a xor b);
    layer0_outputs(4686) <= not b or a;
    layer0_outputs(4687) <= a;
    layer0_outputs(4688) <= not b or a;
    layer0_outputs(4689) <= not b;
    layer0_outputs(4690) <= not (a or b);
    layer0_outputs(4691) <= not b;
    layer0_outputs(4692) <= not (a xor b);
    layer0_outputs(4693) <= not a or b;
    layer0_outputs(4694) <= a or b;
    layer0_outputs(4695) <= a or b;
    layer0_outputs(4696) <= b;
    layer0_outputs(4697) <= a xor b;
    layer0_outputs(4698) <= not a;
    layer0_outputs(4699) <= a xor b;
    layer0_outputs(4700) <= b;
    layer0_outputs(4701) <= a or b;
    layer0_outputs(4702) <= a;
    layer0_outputs(4703) <= not b;
    layer0_outputs(4704) <= a;
    layer0_outputs(4705) <= not (a or b);
    layer0_outputs(4706) <= b;
    layer0_outputs(4707) <= not a;
    layer0_outputs(4708) <= b and not a;
    layer0_outputs(4709) <= b and not a;
    layer0_outputs(4710) <= not a;
    layer0_outputs(4711) <= a xor b;
    layer0_outputs(4712) <= a and not b;
    layer0_outputs(4713) <= a or b;
    layer0_outputs(4714) <= a and not b;
    layer0_outputs(4715) <= not (a and b);
    layer0_outputs(4716) <= b;
    layer0_outputs(4717) <= not a or b;
    layer0_outputs(4718) <= not a;
    layer0_outputs(4719) <= not (a xor b);
    layer0_outputs(4720) <= not a or b;
    layer0_outputs(4721) <= not (a or b);
    layer0_outputs(4722) <= not b or a;
    layer0_outputs(4723) <= a;
    layer0_outputs(4724) <= '0';
    layer0_outputs(4725) <= a or b;
    layer0_outputs(4726) <= not (a xor b);
    layer0_outputs(4727) <= a and not b;
    layer0_outputs(4728) <= '0';
    layer0_outputs(4729) <= not (a or b);
    layer0_outputs(4730) <= b;
    layer0_outputs(4731) <= a or b;
    layer0_outputs(4732) <= not a or b;
    layer0_outputs(4733) <= not (a or b);
    layer0_outputs(4734) <= a or b;
    layer0_outputs(4735) <= b;
    layer0_outputs(4736) <= not (a xor b);
    layer0_outputs(4737) <= a;
    layer0_outputs(4738) <= not (a xor b);
    layer0_outputs(4739) <= not b;
    layer0_outputs(4740) <= '1';
    layer0_outputs(4741) <= not (a or b);
    layer0_outputs(4742) <= not a;
    layer0_outputs(4743) <= a or b;
    layer0_outputs(4744) <= not a or b;
    layer0_outputs(4745) <= b and not a;
    layer0_outputs(4746) <= not (a xor b);
    layer0_outputs(4747) <= not (a xor b);
    layer0_outputs(4748) <= not a or b;
    layer0_outputs(4749) <= not (a xor b);
    layer0_outputs(4750) <= a and b;
    layer0_outputs(4751) <= not a or b;
    layer0_outputs(4752) <= b;
    layer0_outputs(4753) <= not b or a;
    layer0_outputs(4754) <= a and not b;
    layer0_outputs(4755) <= b;
    layer0_outputs(4756) <= a;
    layer0_outputs(4757) <= not a or b;
    layer0_outputs(4758) <= not (a xor b);
    layer0_outputs(4759) <= not (a xor b);
    layer0_outputs(4760) <= a or b;
    layer0_outputs(4761) <= not b;
    layer0_outputs(4762) <= not (a and b);
    layer0_outputs(4763) <= not a;
    layer0_outputs(4764) <= not a or b;
    layer0_outputs(4765) <= a and not b;
    layer0_outputs(4766) <= a or b;
    layer0_outputs(4767) <= a xor b;
    layer0_outputs(4768) <= a;
    layer0_outputs(4769) <= not b or a;
    layer0_outputs(4770) <= a or b;
    layer0_outputs(4771) <= '0';
    layer0_outputs(4772) <= a and b;
    layer0_outputs(4773) <= a;
    layer0_outputs(4774) <= not b;
    layer0_outputs(4775) <= not (a or b);
    layer0_outputs(4776) <= a or b;
    layer0_outputs(4777) <= not a or b;
    layer0_outputs(4778) <= not b;
    layer0_outputs(4779) <= a and not b;
    layer0_outputs(4780) <= not (a or b);
    layer0_outputs(4781) <= not (a or b);
    layer0_outputs(4782) <= a xor b;
    layer0_outputs(4783) <= a and not b;
    layer0_outputs(4784) <= a and not b;
    layer0_outputs(4785) <= not b;
    layer0_outputs(4786) <= a or b;
    layer0_outputs(4787) <= not a or b;
    layer0_outputs(4788) <= not a or b;
    layer0_outputs(4789) <= a and b;
    layer0_outputs(4790) <= not (a or b);
    layer0_outputs(4791) <= a or b;
    layer0_outputs(4792) <= not (a xor b);
    layer0_outputs(4793) <= not a or b;
    layer0_outputs(4794) <= not (a and b);
    layer0_outputs(4795) <= '0';
    layer0_outputs(4796) <= a or b;
    layer0_outputs(4797) <= not a or b;
    layer0_outputs(4798) <= not (a xor b);
    layer0_outputs(4799) <= not (a or b);
    layer0_outputs(4800) <= a and not b;
    layer0_outputs(4801) <= a or b;
    layer0_outputs(4802) <= not a;
    layer0_outputs(4803) <= a or b;
    layer0_outputs(4804) <= a xor b;
    layer0_outputs(4805) <= not (a xor b);
    layer0_outputs(4806) <= not a or b;
    layer0_outputs(4807) <= b and not a;
    layer0_outputs(4808) <= a;
    layer0_outputs(4809) <= not b;
    layer0_outputs(4810) <= a;
    layer0_outputs(4811) <= b and not a;
    layer0_outputs(4812) <= not b;
    layer0_outputs(4813) <= '1';
    layer0_outputs(4814) <= a or b;
    layer0_outputs(4815) <= not b or a;
    layer0_outputs(4816) <= not (a xor b);
    layer0_outputs(4817) <= a xor b;
    layer0_outputs(4818) <= a or b;
    layer0_outputs(4819) <= not a or b;
    layer0_outputs(4820) <= a xor b;
    layer0_outputs(4821) <= a and b;
    layer0_outputs(4822) <= not (a or b);
    layer0_outputs(4823) <= not (a and b);
    layer0_outputs(4824) <= a xor b;
    layer0_outputs(4825) <= not a;
    layer0_outputs(4826) <= a and b;
    layer0_outputs(4827) <= a xor b;
    layer0_outputs(4828) <= not b;
    layer0_outputs(4829) <= b;
    layer0_outputs(4830) <= a or b;
    layer0_outputs(4831) <= '0';
    layer0_outputs(4832) <= b and not a;
    layer0_outputs(4833) <= not (a xor b);
    layer0_outputs(4834) <= a xor b;
    layer0_outputs(4835) <= not (a or b);
    layer0_outputs(4836) <= a or b;
    layer0_outputs(4837) <= a xor b;
    layer0_outputs(4838) <= not a or b;
    layer0_outputs(4839) <= b;
    layer0_outputs(4840) <= not b or a;
    layer0_outputs(4841) <= b and not a;
    layer0_outputs(4842) <= not (a xor b);
    layer0_outputs(4843) <= a and not b;
    layer0_outputs(4844) <= a or b;
    layer0_outputs(4845) <= a;
    layer0_outputs(4846) <= a;
    layer0_outputs(4847) <= not b or a;
    layer0_outputs(4848) <= a and not b;
    layer0_outputs(4849) <= a and not b;
    layer0_outputs(4850) <= not b or a;
    layer0_outputs(4851) <= b and not a;
    layer0_outputs(4852) <= not b or a;
    layer0_outputs(4853) <= a or b;
    layer0_outputs(4854) <= a xor b;
    layer0_outputs(4855) <= b;
    layer0_outputs(4856) <= not (a or b);
    layer0_outputs(4857) <= '0';
    layer0_outputs(4858) <= not (a or b);
    layer0_outputs(4859) <= not b;
    layer0_outputs(4860) <= a;
    layer0_outputs(4861) <= a xor b;
    layer0_outputs(4862) <= not a or b;
    layer0_outputs(4863) <= a;
    layer0_outputs(4864) <= b and not a;
    layer0_outputs(4865) <= not (a or b);
    layer0_outputs(4866) <= not (a or b);
    layer0_outputs(4867) <= not (a or b);
    layer0_outputs(4868) <= a xor b;
    layer0_outputs(4869) <= a;
    layer0_outputs(4870) <= not (a xor b);
    layer0_outputs(4871) <= not (a xor b);
    layer0_outputs(4872) <= not (a xor b);
    layer0_outputs(4873) <= a or b;
    layer0_outputs(4874) <= not (a or b);
    layer0_outputs(4875) <= not b or a;
    layer0_outputs(4876) <= a or b;
    layer0_outputs(4877) <= b and not a;
    layer0_outputs(4878) <= a and b;
    layer0_outputs(4879) <= not b;
    layer0_outputs(4880) <= a;
    layer0_outputs(4881) <= not a or b;
    layer0_outputs(4882) <= b and not a;
    layer0_outputs(4883) <= a xor b;
    layer0_outputs(4884) <= not a or b;
    layer0_outputs(4885) <= a;
    layer0_outputs(4886) <= not (a xor b);
    layer0_outputs(4887) <= not (a xor b);
    layer0_outputs(4888) <= a and b;
    layer0_outputs(4889) <= not (a or b);
    layer0_outputs(4890) <= a xor b;
    layer0_outputs(4891) <= b and not a;
    layer0_outputs(4892) <= '1';
    layer0_outputs(4893) <= a xor b;
    layer0_outputs(4894) <= a xor b;
    layer0_outputs(4895) <= not (a xor b);
    layer0_outputs(4896) <= not (a or b);
    layer0_outputs(4897) <= not a or b;
    layer0_outputs(4898) <= b and not a;
    layer0_outputs(4899) <= b and not a;
    layer0_outputs(4900) <= not (a and b);
    layer0_outputs(4901) <= a and b;
    layer0_outputs(4902) <= not b;
    layer0_outputs(4903) <= not b or a;
    layer0_outputs(4904) <= '1';
    layer0_outputs(4905) <= a;
    layer0_outputs(4906) <= a and not b;
    layer0_outputs(4907) <= not (a and b);
    layer0_outputs(4908) <= a;
    layer0_outputs(4909) <= a and not b;
    layer0_outputs(4910) <= not (a or b);
    layer0_outputs(4911) <= b;
    layer0_outputs(4912) <= not (a xor b);
    layer0_outputs(4913) <= not (a or b);
    layer0_outputs(4914) <= not a;
    layer0_outputs(4915) <= b and not a;
    layer0_outputs(4916) <= a xor b;
    layer0_outputs(4917) <= a;
    layer0_outputs(4918) <= a xor b;
    layer0_outputs(4919) <= a;
    layer0_outputs(4920) <= a or b;
    layer0_outputs(4921) <= not (a or b);
    layer0_outputs(4922) <= a and not b;
    layer0_outputs(4923) <= not (a or b);
    layer0_outputs(4924) <= '0';
    layer0_outputs(4925) <= not (a or b);
    layer0_outputs(4926) <= a and not b;
    layer0_outputs(4927) <= not (a or b);
    layer0_outputs(4928) <= not a or b;
    layer0_outputs(4929) <= not (a xor b);
    layer0_outputs(4930) <= b;
    layer0_outputs(4931) <= '0';
    layer0_outputs(4932) <= a or b;
    layer0_outputs(4933) <= b and not a;
    layer0_outputs(4934) <= a xor b;
    layer0_outputs(4935) <= a xor b;
    layer0_outputs(4936) <= not a or b;
    layer0_outputs(4937) <= not (a or b);
    layer0_outputs(4938) <= a xor b;
    layer0_outputs(4939) <= not (a and b);
    layer0_outputs(4940) <= '0';
    layer0_outputs(4941) <= b;
    layer0_outputs(4942) <= a or b;
    layer0_outputs(4943) <= a and b;
    layer0_outputs(4944) <= not (a xor b);
    layer0_outputs(4945) <= not a;
    layer0_outputs(4946) <= not (a xor b);
    layer0_outputs(4947) <= a;
    layer0_outputs(4948) <= a xor b;
    layer0_outputs(4949) <= '1';
    layer0_outputs(4950) <= not (a or b);
    layer0_outputs(4951) <= a or b;
    layer0_outputs(4952) <= b;
    layer0_outputs(4953) <= a or b;
    layer0_outputs(4954) <= b;
    layer0_outputs(4955) <= '1';
    layer0_outputs(4956) <= not (a xor b);
    layer0_outputs(4957) <= '0';
    layer0_outputs(4958) <= not (a or b);
    layer0_outputs(4959) <= a and not b;
    layer0_outputs(4960) <= a and not b;
    layer0_outputs(4961) <= a and not b;
    layer0_outputs(4962) <= not a or b;
    layer0_outputs(4963) <= not (a or b);
    layer0_outputs(4964) <= '0';
    layer0_outputs(4965) <= not a or b;
    layer0_outputs(4966) <= not b;
    layer0_outputs(4967) <= not a or b;
    layer0_outputs(4968) <= '0';
    layer0_outputs(4969) <= not (a xor b);
    layer0_outputs(4970) <= not (a xor b);
    layer0_outputs(4971) <= not a;
    layer0_outputs(4972) <= not b or a;
    layer0_outputs(4973) <= not (a or b);
    layer0_outputs(4974) <= a xor b;
    layer0_outputs(4975) <= b and not a;
    layer0_outputs(4976) <= a or b;
    layer0_outputs(4977) <= not (a xor b);
    layer0_outputs(4978) <= a;
    layer0_outputs(4979) <= a or b;
    layer0_outputs(4980) <= not b or a;
    layer0_outputs(4981) <= not (a and b);
    layer0_outputs(4982) <= not (a or b);
    layer0_outputs(4983) <= a;
    layer0_outputs(4984) <= not (a xor b);
    layer0_outputs(4985) <= a;
    layer0_outputs(4986) <= a;
    layer0_outputs(4987) <= '0';
    layer0_outputs(4988) <= a;
    layer0_outputs(4989) <= a;
    layer0_outputs(4990) <= '1';
    layer0_outputs(4991) <= not (a xor b);
    layer0_outputs(4992) <= not (a and b);
    layer0_outputs(4993) <= b;
    layer0_outputs(4994) <= not b;
    layer0_outputs(4995) <= a or b;
    layer0_outputs(4996) <= not a;
    layer0_outputs(4997) <= not a or b;
    layer0_outputs(4998) <= not (a xor b);
    layer0_outputs(4999) <= a;
    layer0_outputs(5000) <= not (a xor b);
    layer0_outputs(5001) <= not (a or b);
    layer0_outputs(5002) <= a and b;
    layer0_outputs(5003) <= a and not b;
    layer0_outputs(5004) <= b and not a;
    layer0_outputs(5005) <= not (a or b);
    layer0_outputs(5006) <= not (a xor b);
    layer0_outputs(5007) <= a or b;
    layer0_outputs(5008) <= a and not b;
    layer0_outputs(5009) <= b and not a;
    layer0_outputs(5010) <= b and not a;
    layer0_outputs(5011) <= '1';
    layer0_outputs(5012) <= not (a or b);
    layer0_outputs(5013) <= a;
    layer0_outputs(5014) <= b and not a;
    layer0_outputs(5015) <= not (a or b);
    layer0_outputs(5016) <= a or b;
    layer0_outputs(5017) <= not (a xor b);
    layer0_outputs(5018) <= a;
    layer0_outputs(5019) <= a or b;
    layer0_outputs(5020) <= a xor b;
    layer0_outputs(5021) <= not (a or b);
    layer0_outputs(5022) <= a xor b;
    layer0_outputs(5023) <= not a;
    layer0_outputs(5024) <= not a;
    layer0_outputs(5025) <= a;
    layer0_outputs(5026) <= b and not a;
    layer0_outputs(5027) <= a xor b;
    layer0_outputs(5028) <= not a or b;
    layer0_outputs(5029) <= not a;
    layer0_outputs(5030) <= not a or b;
    layer0_outputs(5031) <= not (a or b);
    layer0_outputs(5032) <= b and not a;
    layer0_outputs(5033) <= not b;
    layer0_outputs(5034) <= not b;
    layer0_outputs(5035) <= not (a xor b);
    layer0_outputs(5036) <= not (a or b);
    layer0_outputs(5037) <= b and not a;
    layer0_outputs(5038) <= not (a and b);
    layer0_outputs(5039) <= a and b;
    layer0_outputs(5040) <= not (a xor b);
    layer0_outputs(5041) <= not a or b;
    layer0_outputs(5042) <= not b or a;
    layer0_outputs(5043) <= b and not a;
    layer0_outputs(5044) <= '0';
    layer0_outputs(5045) <= a;
    layer0_outputs(5046) <= not a;
    layer0_outputs(5047) <= not a or b;
    layer0_outputs(5048) <= a and b;
    layer0_outputs(5049) <= a and not b;
    layer0_outputs(5050) <= not (a xor b);
    layer0_outputs(5051) <= a and not b;
    layer0_outputs(5052) <= not b or a;
    layer0_outputs(5053) <= '1';
    layer0_outputs(5054) <= not b;
    layer0_outputs(5055) <= not a;
    layer0_outputs(5056) <= not (a xor b);
    layer0_outputs(5057) <= not (a xor b);
    layer0_outputs(5058) <= not a or b;
    layer0_outputs(5059) <= not (a or b);
    layer0_outputs(5060) <= a and b;
    layer0_outputs(5061) <= not b;
    layer0_outputs(5062) <= not b;
    layer0_outputs(5063) <= not b;
    layer0_outputs(5064) <= a or b;
    layer0_outputs(5065) <= a or b;
    layer0_outputs(5066) <= a xor b;
    layer0_outputs(5067) <= b and not a;
    layer0_outputs(5068) <= a;
    layer0_outputs(5069) <= a or b;
    layer0_outputs(5070) <= not (a or b);
    layer0_outputs(5071) <= a;
    layer0_outputs(5072) <= a and b;
    layer0_outputs(5073) <= '0';
    layer0_outputs(5074) <= a xor b;
    layer0_outputs(5075) <= not (a or b);
    layer0_outputs(5076) <= not a or b;
    layer0_outputs(5077) <= not (a xor b);
    layer0_outputs(5078) <= a xor b;
    layer0_outputs(5079) <= not (a or b);
    layer0_outputs(5080) <= not b or a;
    layer0_outputs(5081) <= not (a or b);
    layer0_outputs(5082) <= '1';
    layer0_outputs(5083) <= a xor b;
    layer0_outputs(5084) <= a xor b;
    layer0_outputs(5085) <= not (a xor b);
    layer0_outputs(5086) <= not a or b;
    layer0_outputs(5087) <= not (a xor b);
    layer0_outputs(5088) <= b and not a;
    layer0_outputs(5089) <= b;
    layer0_outputs(5090) <= not a;
    layer0_outputs(5091) <= b;
    layer0_outputs(5092) <= a and not b;
    layer0_outputs(5093) <= a or b;
    layer0_outputs(5094) <= b;
    layer0_outputs(5095) <= not b;
    layer0_outputs(5096) <= not a or b;
    layer0_outputs(5097) <= not (a and b);
    layer0_outputs(5098) <= a and not b;
    layer0_outputs(5099) <= a or b;
    layer0_outputs(5100) <= b and not a;
    layer0_outputs(5101) <= not a or b;
    layer0_outputs(5102) <= a or b;
    layer0_outputs(5103) <= '0';
    layer0_outputs(5104) <= not b or a;
    layer0_outputs(5105) <= not a or b;
    layer0_outputs(5106) <= a or b;
    layer0_outputs(5107) <= not (a xor b);
    layer0_outputs(5108) <= not a or b;
    layer0_outputs(5109) <= not (a xor b);
    layer0_outputs(5110) <= not (a or b);
    layer0_outputs(5111) <= not a or b;
    layer0_outputs(5112) <= a and not b;
    layer0_outputs(5113) <= b;
    layer0_outputs(5114) <= b;
    layer0_outputs(5115) <= not a or b;
    layer0_outputs(5116) <= a xor b;
    layer0_outputs(5117) <= a xor b;
    layer0_outputs(5118) <= not b or a;
    layer0_outputs(5119) <= a or b;
    layer0_outputs(5120) <= not b or a;
    layer0_outputs(5121) <= a xor b;
    layer0_outputs(5122) <= a;
    layer0_outputs(5123) <= not a or b;
    layer0_outputs(5124) <= not (a xor b);
    layer0_outputs(5125) <= not a or b;
    layer0_outputs(5126) <= a or b;
    layer0_outputs(5127) <= not b;
    layer0_outputs(5128) <= a xor b;
    layer0_outputs(5129) <= a and b;
    layer0_outputs(5130) <= a;
    layer0_outputs(5131) <= not b or a;
    layer0_outputs(5132) <= a and not b;
    layer0_outputs(5133) <= not a;
    layer0_outputs(5134) <= not a or b;
    layer0_outputs(5135) <= not (a or b);
    layer0_outputs(5136) <= not (a or b);
    layer0_outputs(5137) <= not (a or b);
    layer0_outputs(5138) <= a xor b;
    layer0_outputs(5139) <= a or b;
    layer0_outputs(5140) <= not (a xor b);
    layer0_outputs(5141) <= not b or a;
    layer0_outputs(5142) <= a xor b;
    layer0_outputs(5143) <= not (a xor b);
    layer0_outputs(5144) <= not (a or b);
    layer0_outputs(5145) <= a or b;
    layer0_outputs(5146) <= not a or b;
    layer0_outputs(5147) <= '0';
    layer0_outputs(5148) <= not a or b;
    layer0_outputs(5149) <= not b;
    layer0_outputs(5150) <= a and b;
    layer0_outputs(5151) <= not b or a;
    layer0_outputs(5152) <= b;
    layer0_outputs(5153) <= a or b;
    layer0_outputs(5154) <= not (a and b);
    layer0_outputs(5155) <= not b;
    layer0_outputs(5156) <= b;
    layer0_outputs(5157) <= a and b;
    layer0_outputs(5158) <= a and not b;
    layer0_outputs(5159) <= a xor b;
    layer0_outputs(5160) <= not b;
    layer0_outputs(5161) <= not a or b;
    layer0_outputs(5162) <= not b or a;
    layer0_outputs(5163) <= b;
    layer0_outputs(5164) <= not (a or b);
    layer0_outputs(5165) <= not (a or b);
    layer0_outputs(5166) <= a;
    layer0_outputs(5167) <= not (a and b);
    layer0_outputs(5168) <= a or b;
    layer0_outputs(5169) <= a xor b;
    layer0_outputs(5170) <= b and not a;
    layer0_outputs(5171) <= not (a and b);
    layer0_outputs(5172) <= not a;
    layer0_outputs(5173) <= a;
    layer0_outputs(5174) <= a xor b;
    layer0_outputs(5175) <= not (a and b);
    layer0_outputs(5176) <= not b or a;
    layer0_outputs(5177) <= a or b;
    layer0_outputs(5178) <= not (a xor b);
    layer0_outputs(5179) <= a xor b;
    layer0_outputs(5180) <= not (a xor b);
    layer0_outputs(5181) <= not (a xor b);
    layer0_outputs(5182) <= not (a xor b);
    layer0_outputs(5183) <= a or b;
    layer0_outputs(5184) <= '1';
    layer0_outputs(5185) <= not a or b;
    layer0_outputs(5186) <= '0';
    layer0_outputs(5187) <= a xor b;
    layer0_outputs(5188) <= a or b;
    layer0_outputs(5189) <= a xor b;
    layer0_outputs(5190) <= not (a or b);
    layer0_outputs(5191) <= not b or a;
    layer0_outputs(5192) <= not b;
    layer0_outputs(5193) <= not b;
    layer0_outputs(5194) <= b and not a;
    layer0_outputs(5195) <= not (a or b);
    layer0_outputs(5196) <= a xor b;
    layer0_outputs(5197) <= not (a or b);
    layer0_outputs(5198) <= not (a or b);
    layer0_outputs(5199) <= a xor b;
    layer0_outputs(5200) <= a and not b;
    layer0_outputs(5201) <= not (a xor b);
    layer0_outputs(5202) <= a xor b;
    layer0_outputs(5203) <= b;
    layer0_outputs(5204) <= a and not b;
    layer0_outputs(5205) <= b and not a;
    layer0_outputs(5206) <= '0';
    layer0_outputs(5207) <= not b;
    layer0_outputs(5208) <= a and not b;
    layer0_outputs(5209) <= not b;
    layer0_outputs(5210) <= a or b;
    layer0_outputs(5211) <= a and not b;
    layer0_outputs(5212) <= a;
    layer0_outputs(5213) <= a and not b;
    layer0_outputs(5214) <= not b;
    layer0_outputs(5215) <= not b;
    layer0_outputs(5216) <= not (a or b);
    layer0_outputs(5217) <= a;
    layer0_outputs(5218) <= not (a xor b);
    layer0_outputs(5219) <= not a;
    layer0_outputs(5220) <= a;
    layer0_outputs(5221) <= not a or b;
    layer0_outputs(5222) <= not b or a;
    layer0_outputs(5223) <= not b or a;
    layer0_outputs(5224) <= a and b;
    layer0_outputs(5225) <= not b or a;
    layer0_outputs(5226) <= not (a xor b);
    layer0_outputs(5227) <= a or b;
    layer0_outputs(5228) <= a and not b;
    layer0_outputs(5229) <= not b or a;
    layer0_outputs(5230) <= b;
    layer0_outputs(5231) <= not (a and b);
    layer0_outputs(5232) <= not b or a;
    layer0_outputs(5233) <= b;
    layer0_outputs(5234) <= b and not a;
    layer0_outputs(5235) <= not (a xor b);
    layer0_outputs(5236) <= a;
    layer0_outputs(5237) <= not b or a;
    layer0_outputs(5238) <= not (a or b);
    layer0_outputs(5239) <= '0';
    layer0_outputs(5240) <= '1';
    layer0_outputs(5241) <= not a or b;
    layer0_outputs(5242) <= a;
    layer0_outputs(5243) <= not b;
    layer0_outputs(5244) <= a xor b;
    layer0_outputs(5245) <= a and not b;
    layer0_outputs(5246) <= not (a or b);
    layer0_outputs(5247) <= a or b;
    layer0_outputs(5248) <= a or b;
    layer0_outputs(5249) <= not b;
    layer0_outputs(5250) <= '1';
    layer0_outputs(5251) <= a xor b;
    layer0_outputs(5252) <= not (a or b);
    layer0_outputs(5253) <= a or b;
    layer0_outputs(5254) <= a;
    layer0_outputs(5255) <= not a;
    layer0_outputs(5256) <= a xor b;
    layer0_outputs(5257) <= not (a or b);
    layer0_outputs(5258) <= b;
    layer0_outputs(5259) <= '1';
    layer0_outputs(5260) <= a or b;
    layer0_outputs(5261) <= a;
    layer0_outputs(5262) <= a and b;
    layer0_outputs(5263) <= b;
    layer0_outputs(5264) <= not (a or b);
    layer0_outputs(5265) <= not b;
    layer0_outputs(5266) <= not b or a;
    layer0_outputs(5267) <= not b or a;
    layer0_outputs(5268) <= a xor b;
    layer0_outputs(5269) <= a and b;
    layer0_outputs(5270) <= not a or b;
    layer0_outputs(5271) <= not a;
    layer0_outputs(5272) <= not b;
    layer0_outputs(5273) <= a and not b;
    layer0_outputs(5274) <= not b;
    layer0_outputs(5275) <= a and not b;
    layer0_outputs(5276) <= a and b;
    layer0_outputs(5277) <= b;
    layer0_outputs(5278) <= not a;
    layer0_outputs(5279) <= not a;
    layer0_outputs(5280) <= not a or b;
    layer0_outputs(5281) <= not b or a;
    layer0_outputs(5282) <= not b or a;
    layer0_outputs(5283) <= not (a xor b);
    layer0_outputs(5284) <= a;
    layer0_outputs(5285) <= not b;
    layer0_outputs(5286) <= a and not b;
    layer0_outputs(5287) <= a xor b;
    layer0_outputs(5288) <= b;
    layer0_outputs(5289) <= a xor b;
    layer0_outputs(5290) <= a xor b;
    layer0_outputs(5291) <= not a;
    layer0_outputs(5292) <= not a or b;
    layer0_outputs(5293) <= a and not b;
    layer0_outputs(5294) <= not a or b;
    layer0_outputs(5295) <= not (a and b);
    layer0_outputs(5296) <= a or b;
    layer0_outputs(5297) <= not (a or b);
    layer0_outputs(5298) <= a or b;
    layer0_outputs(5299) <= a and b;
    layer0_outputs(5300) <= a;
    layer0_outputs(5301) <= a and not b;
    layer0_outputs(5302) <= not (a or b);
    layer0_outputs(5303) <= a or b;
    layer0_outputs(5304) <= not (a and b);
    layer0_outputs(5305) <= not b or a;
    layer0_outputs(5306) <= not a or b;
    layer0_outputs(5307) <= not (a xor b);
    layer0_outputs(5308) <= a or b;
    layer0_outputs(5309) <= not (a xor b);
    layer0_outputs(5310) <= b;
    layer0_outputs(5311) <= b and not a;
    layer0_outputs(5312) <= a and not b;
    layer0_outputs(5313) <= b;
    layer0_outputs(5314) <= not a or b;
    layer0_outputs(5315) <= not (a xor b);
    layer0_outputs(5316) <= not (a or b);
    layer0_outputs(5317) <= a and not b;
    layer0_outputs(5318) <= b;
    layer0_outputs(5319) <= not a;
    layer0_outputs(5320) <= a and b;
    layer0_outputs(5321) <= not b;
    layer0_outputs(5322) <= a or b;
    layer0_outputs(5323) <= not b or a;
    layer0_outputs(5324) <= a or b;
    layer0_outputs(5325) <= not (a or b);
    layer0_outputs(5326) <= a xor b;
    layer0_outputs(5327) <= not b or a;
    layer0_outputs(5328) <= b and not a;
    layer0_outputs(5329) <= a;
    layer0_outputs(5330) <= a;
    layer0_outputs(5331) <= not (a or b);
    layer0_outputs(5332) <= not a or b;
    layer0_outputs(5333) <= not a;
    layer0_outputs(5334) <= a or b;
    layer0_outputs(5335) <= not (a xor b);
    layer0_outputs(5336) <= a xor b;
    layer0_outputs(5337) <= not (a xor b);
    layer0_outputs(5338) <= not a or b;
    layer0_outputs(5339) <= a or b;
    layer0_outputs(5340) <= not a or b;
    layer0_outputs(5341) <= not (a or b);
    layer0_outputs(5342) <= a or b;
    layer0_outputs(5343) <= b and not a;
    layer0_outputs(5344) <= '0';
    layer0_outputs(5345) <= b and not a;
    layer0_outputs(5346) <= b;
    layer0_outputs(5347) <= a and not b;
    layer0_outputs(5348) <= not (a or b);
    layer0_outputs(5349) <= a or b;
    layer0_outputs(5350) <= a or b;
    layer0_outputs(5351) <= a xor b;
    layer0_outputs(5352) <= not b;
    layer0_outputs(5353) <= b;
    layer0_outputs(5354) <= a;
    layer0_outputs(5355) <= not (a xor b);
    layer0_outputs(5356) <= a xor b;
    layer0_outputs(5357) <= not a or b;
    layer0_outputs(5358) <= not b or a;
    layer0_outputs(5359) <= '0';
    layer0_outputs(5360) <= b and not a;
    layer0_outputs(5361) <= a;
    layer0_outputs(5362) <= a xor b;
    layer0_outputs(5363) <= b and not a;
    layer0_outputs(5364) <= a xor b;
    layer0_outputs(5365) <= not b or a;
    layer0_outputs(5366) <= b and not a;
    layer0_outputs(5367) <= b;
    layer0_outputs(5368) <= not (a or b);
    layer0_outputs(5369) <= a xor b;
    layer0_outputs(5370) <= b;
    layer0_outputs(5371) <= not (a xor b);
    layer0_outputs(5372) <= not b or a;
    layer0_outputs(5373) <= not (a or b);
    layer0_outputs(5374) <= not (a xor b);
    layer0_outputs(5375) <= '1';
    layer0_outputs(5376) <= a and not b;
    layer0_outputs(5377) <= a or b;
    layer0_outputs(5378) <= not b or a;
    layer0_outputs(5379) <= '1';
    layer0_outputs(5380) <= a;
    layer0_outputs(5381) <= not a or b;
    layer0_outputs(5382) <= a xor b;
    layer0_outputs(5383) <= a and not b;
    layer0_outputs(5384) <= b;
    layer0_outputs(5385) <= not (a xor b);
    layer0_outputs(5386) <= a;
    layer0_outputs(5387) <= not (a or b);
    layer0_outputs(5388) <= a and not b;
    layer0_outputs(5389) <= not a;
    layer0_outputs(5390) <= not b or a;
    layer0_outputs(5391) <= b and not a;
    layer0_outputs(5392) <= not a or b;
    layer0_outputs(5393) <= not (a or b);
    layer0_outputs(5394) <= a or b;
    layer0_outputs(5395) <= a xor b;
    layer0_outputs(5396) <= not a;
    layer0_outputs(5397) <= not (a or b);
    layer0_outputs(5398) <= not a or b;
    layer0_outputs(5399) <= not (a and b);
    layer0_outputs(5400) <= not b or a;
    layer0_outputs(5401) <= a or b;
    layer0_outputs(5402) <= not (a or b);
    layer0_outputs(5403) <= a or b;
    layer0_outputs(5404) <= a xor b;
    layer0_outputs(5405) <= a or b;
    layer0_outputs(5406) <= not b;
    layer0_outputs(5407) <= not a;
    layer0_outputs(5408) <= b and not a;
    layer0_outputs(5409) <= a xor b;
    layer0_outputs(5410) <= a or b;
    layer0_outputs(5411) <= not (a xor b);
    layer0_outputs(5412) <= a xor b;
    layer0_outputs(5413) <= not a;
    layer0_outputs(5414) <= not a;
    layer0_outputs(5415) <= a or b;
    layer0_outputs(5416) <= a xor b;
    layer0_outputs(5417) <= a xor b;
    layer0_outputs(5418) <= '0';
    layer0_outputs(5419) <= a and not b;
    layer0_outputs(5420) <= not (a xor b);
    layer0_outputs(5421) <= a or b;
    layer0_outputs(5422) <= a or b;
    layer0_outputs(5423) <= a or b;
    layer0_outputs(5424) <= '1';
    layer0_outputs(5425) <= not (a or b);
    layer0_outputs(5426) <= not (a xor b);
    layer0_outputs(5427) <= a and not b;
    layer0_outputs(5428) <= a;
    layer0_outputs(5429) <= not b or a;
    layer0_outputs(5430) <= not b or a;
    layer0_outputs(5431) <= a;
    layer0_outputs(5432) <= a or b;
    layer0_outputs(5433) <= not (a and b);
    layer0_outputs(5434) <= '0';
    layer0_outputs(5435) <= a or b;
    layer0_outputs(5436) <= '1';
    layer0_outputs(5437) <= not (a xor b);
    layer0_outputs(5438) <= not (a or b);
    layer0_outputs(5439) <= not a or b;
    layer0_outputs(5440) <= not (a or b);
    layer0_outputs(5441) <= not a or b;
    layer0_outputs(5442) <= not a or b;
    layer0_outputs(5443) <= a and not b;
    layer0_outputs(5444) <= a or b;
    layer0_outputs(5445) <= not (a xor b);
    layer0_outputs(5446) <= a and not b;
    layer0_outputs(5447) <= '0';
    layer0_outputs(5448) <= b;
    layer0_outputs(5449) <= a xor b;
    layer0_outputs(5450) <= not b;
    layer0_outputs(5451) <= not a or b;
    layer0_outputs(5452) <= not a;
    layer0_outputs(5453) <= not a;
    layer0_outputs(5454) <= '0';
    layer0_outputs(5455) <= not a or b;
    layer0_outputs(5456) <= b;
    layer0_outputs(5457) <= '0';
    layer0_outputs(5458) <= a and b;
    layer0_outputs(5459) <= a xor b;
    layer0_outputs(5460) <= a and b;
    layer0_outputs(5461) <= not a;
    layer0_outputs(5462) <= not a;
    layer0_outputs(5463) <= not (a xor b);
    layer0_outputs(5464) <= '0';
    layer0_outputs(5465) <= not b;
    layer0_outputs(5466) <= a and b;
    layer0_outputs(5467) <= a;
    layer0_outputs(5468) <= not a or b;
    layer0_outputs(5469) <= b and not a;
    layer0_outputs(5470) <= not b or a;
    layer0_outputs(5471) <= not b or a;
    layer0_outputs(5472) <= a and not b;
    layer0_outputs(5473) <= not a or b;
    layer0_outputs(5474) <= a;
    layer0_outputs(5475) <= not (a and b);
    layer0_outputs(5476) <= a;
    layer0_outputs(5477) <= not (a xor b);
    layer0_outputs(5478) <= not a or b;
    layer0_outputs(5479) <= a and not b;
    layer0_outputs(5480) <= a xor b;
    layer0_outputs(5481) <= a;
    layer0_outputs(5482) <= b and not a;
    layer0_outputs(5483) <= a or b;
    layer0_outputs(5484) <= '1';
    layer0_outputs(5485) <= '1';
    layer0_outputs(5486) <= b;
    layer0_outputs(5487) <= a or b;
    layer0_outputs(5488) <= a or b;
    layer0_outputs(5489) <= not b or a;
    layer0_outputs(5490) <= a or b;
    layer0_outputs(5491) <= '0';
    layer0_outputs(5492) <= not (a or b);
    layer0_outputs(5493) <= not b;
    layer0_outputs(5494) <= a or b;
    layer0_outputs(5495) <= not (a and b);
    layer0_outputs(5496) <= not (a or b);
    layer0_outputs(5497) <= a xor b;
    layer0_outputs(5498) <= b;
    layer0_outputs(5499) <= a and b;
    layer0_outputs(5500) <= a or b;
    layer0_outputs(5501) <= a or b;
    layer0_outputs(5502) <= b and not a;
    layer0_outputs(5503) <= not (a and b);
    layer0_outputs(5504) <= not b or a;
    layer0_outputs(5505) <= a or b;
    layer0_outputs(5506) <= not a;
    layer0_outputs(5507) <= not a;
    layer0_outputs(5508) <= not (a or b);
    layer0_outputs(5509) <= not b or a;
    layer0_outputs(5510) <= a;
    layer0_outputs(5511) <= a xor b;
    layer0_outputs(5512) <= not (a and b);
    layer0_outputs(5513) <= b and not a;
    layer0_outputs(5514) <= a xor b;
    layer0_outputs(5515) <= not b;
    layer0_outputs(5516) <= b;
    layer0_outputs(5517) <= not a;
    layer0_outputs(5518) <= not a;
    layer0_outputs(5519) <= not a or b;
    layer0_outputs(5520) <= a;
    layer0_outputs(5521) <= b and not a;
    layer0_outputs(5522) <= not (a xor b);
    layer0_outputs(5523) <= a or b;
    layer0_outputs(5524) <= b;
    layer0_outputs(5525) <= not a or b;
    layer0_outputs(5526) <= a xor b;
    layer0_outputs(5527) <= a xor b;
    layer0_outputs(5528) <= not (a xor b);
    layer0_outputs(5529) <= not b;
    layer0_outputs(5530) <= not a;
    layer0_outputs(5531) <= not (a or b);
    layer0_outputs(5532) <= a or b;
    layer0_outputs(5533) <= not a or b;
    layer0_outputs(5534) <= not (a xor b);
    layer0_outputs(5535) <= a or b;
    layer0_outputs(5536) <= not (a xor b);
    layer0_outputs(5537) <= not (a or b);
    layer0_outputs(5538) <= not a or b;
    layer0_outputs(5539) <= not b;
    layer0_outputs(5540) <= not a;
    layer0_outputs(5541) <= not b or a;
    layer0_outputs(5542) <= a and not b;
    layer0_outputs(5543) <= not (a or b);
    layer0_outputs(5544) <= not b;
    layer0_outputs(5545) <= not b;
    layer0_outputs(5546) <= not a or b;
    layer0_outputs(5547) <= a;
    layer0_outputs(5548) <= not (a or b);
    layer0_outputs(5549) <= '1';
    layer0_outputs(5550) <= not b;
    layer0_outputs(5551) <= not (a or b);
    layer0_outputs(5552) <= not (a or b);
    layer0_outputs(5553) <= not a or b;
    layer0_outputs(5554) <= b and not a;
    layer0_outputs(5555) <= a or b;
    layer0_outputs(5556) <= a xor b;
    layer0_outputs(5557) <= not a;
    layer0_outputs(5558) <= b and not a;
    layer0_outputs(5559) <= a or b;
    layer0_outputs(5560) <= not a;
    layer0_outputs(5561) <= a and not b;
    layer0_outputs(5562) <= not (a xor b);
    layer0_outputs(5563) <= b;
    layer0_outputs(5564) <= not (a xor b);
    layer0_outputs(5565) <= a and b;
    layer0_outputs(5566) <= not b;
    layer0_outputs(5567) <= '0';
    layer0_outputs(5568) <= b;
    layer0_outputs(5569) <= '1';
    layer0_outputs(5570) <= '0';
    layer0_outputs(5571) <= not a;
    layer0_outputs(5572) <= a or b;
    layer0_outputs(5573) <= not a or b;
    layer0_outputs(5574) <= not b;
    layer0_outputs(5575) <= not (a or b);
    layer0_outputs(5576) <= '0';
    layer0_outputs(5577) <= '0';
    layer0_outputs(5578) <= b and not a;
    layer0_outputs(5579) <= not (a or b);
    layer0_outputs(5580) <= a or b;
    layer0_outputs(5581) <= b;
    layer0_outputs(5582) <= a and not b;
    layer0_outputs(5583) <= not a;
    layer0_outputs(5584) <= not a;
    layer0_outputs(5585) <= a and not b;
    layer0_outputs(5586) <= not (a or b);
    layer0_outputs(5587) <= b;
    layer0_outputs(5588) <= b and not a;
    layer0_outputs(5589) <= not a or b;
    layer0_outputs(5590) <= not (a and b);
    layer0_outputs(5591) <= '0';
    layer0_outputs(5592) <= b and not a;
    layer0_outputs(5593) <= not a;
    layer0_outputs(5594) <= b;
    layer0_outputs(5595) <= not (a xor b);
    layer0_outputs(5596) <= a xor b;
    layer0_outputs(5597) <= a xor b;
    layer0_outputs(5598) <= not (a xor b);
    layer0_outputs(5599) <= not (a or b);
    layer0_outputs(5600) <= not a;
    layer0_outputs(5601) <= b and not a;
    layer0_outputs(5602) <= a xor b;
    layer0_outputs(5603) <= '0';
    layer0_outputs(5604) <= not (a xor b);
    layer0_outputs(5605) <= a or b;
    layer0_outputs(5606) <= not b;
    layer0_outputs(5607) <= not (a xor b);
    layer0_outputs(5608) <= not (a xor b);
    layer0_outputs(5609) <= not (a or b);
    layer0_outputs(5610) <= a and not b;
    layer0_outputs(5611) <= not a or b;
    layer0_outputs(5612) <= a and not b;
    layer0_outputs(5613) <= '1';
    layer0_outputs(5614) <= not b;
    layer0_outputs(5615) <= a xor b;
    layer0_outputs(5616) <= a and not b;
    layer0_outputs(5617) <= b;
    layer0_outputs(5618) <= b;
    layer0_outputs(5619) <= a;
    layer0_outputs(5620) <= not (a xor b);
    layer0_outputs(5621) <= a xor b;
    layer0_outputs(5622) <= not a;
    layer0_outputs(5623) <= not a;
    layer0_outputs(5624) <= not (a or b);
    layer0_outputs(5625) <= a xor b;
    layer0_outputs(5626) <= a xor b;
    layer0_outputs(5627) <= not (a xor b);
    layer0_outputs(5628) <= a xor b;
    layer0_outputs(5629) <= not (a xor b);
    layer0_outputs(5630) <= a and not b;
    layer0_outputs(5631) <= not (a or b);
    layer0_outputs(5632) <= a;
    layer0_outputs(5633) <= not a or b;
    layer0_outputs(5634) <= '1';
    layer0_outputs(5635) <= a;
    layer0_outputs(5636) <= a;
    layer0_outputs(5637) <= '1';
    layer0_outputs(5638) <= not b;
    layer0_outputs(5639) <= a or b;
    layer0_outputs(5640) <= a and not b;
    layer0_outputs(5641) <= a and b;
    layer0_outputs(5642) <= not (a xor b);
    layer0_outputs(5643) <= not a or b;
    layer0_outputs(5644) <= b and not a;
    layer0_outputs(5645) <= not (a or b);
    layer0_outputs(5646) <= not (a or b);
    layer0_outputs(5647) <= '1';
    layer0_outputs(5648) <= a and not b;
    layer0_outputs(5649) <= not (a or b);
    layer0_outputs(5650) <= a xor b;
    layer0_outputs(5651) <= not (a xor b);
    layer0_outputs(5652) <= not b;
    layer0_outputs(5653) <= not (a and b);
    layer0_outputs(5654) <= not (a xor b);
    layer0_outputs(5655) <= not b;
    layer0_outputs(5656) <= not (a or b);
    layer0_outputs(5657) <= not (a xor b);
    layer0_outputs(5658) <= a or b;
    layer0_outputs(5659) <= a;
    layer0_outputs(5660) <= b;
    layer0_outputs(5661) <= not (a xor b);
    layer0_outputs(5662) <= '1';
    layer0_outputs(5663) <= not a or b;
    layer0_outputs(5664) <= not (a or b);
    layer0_outputs(5665) <= not (a or b);
    layer0_outputs(5666) <= b and not a;
    layer0_outputs(5667) <= not (a and b);
    layer0_outputs(5668) <= b;
    layer0_outputs(5669) <= not (a or b);
    layer0_outputs(5670) <= a and not b;
    layer0_outputs(5671) <= a and not b;
    layer0_outputs(5672) <= a xor b;
    layer0_outputs(5673) <= not (a xor b);
    layer0_outputs(5674) <= '1';
    layer0_outputs(5675) <= not a;
    layer0_outputs(5676) <= b and not a;
    layer0_outputs(5677) <= not (a or b);
    layer0_outputs(5678) <= a or b;
    layer0_outputs(5679) <= not (a xor b);
    layer0_outputs(5680) <= not a;
    layer0_outputs(5681) <= not a or b;
    layer0_outputs(5682) <= not b;
    layer0_outputs(5683) <= '1';
    layer0_outputs(5684) <= a or b;
    layer0_outputs(5685) <= b;
    layer0_outputs(5686) <= not b or a;
    layer0_outputs(5687) <= not a or b;
    layer0_outputs(5688) <= b;
    layer0_outputs(5689) <= not b;
    layer0_outputs(5690) <= a or b;
    layer0_outputs(5691) <= not b or a;
    layer0_outputs(5692) <= not (a xor b);
    layer0_outputs(5693) <= a or b;
    layer0_outputs(5694) <= b and not a;
    layer0_outputs(5695) <= not a;
    layer0_outputs(5696) <= not (a xor b);
    layer0_outputs(5697) <= '0';
    layer0_outputs(5698) <= a or b;
    layer0_outputs(5699) <= not b or a;
    layer0_outputs(5700) <= not b;
    layer0_outputs(5701) <= a and not b;
    layer0_outputs(5702) <= not a;
    layer0_outputs(5703) <= not (a or b);
    layer0_outputs(5704) <= not b or a;
    layer0_outputs(5705) <= '1';
    layer0_outputs(5706) <= a or b;
    layer0_outputs(5707) <= a or b;
    layer0_outputs(5708) <= not b;
    layer0_outputs(5709) <= b;
    layer0_outputs(5710) <= not b or a;
    layer0_outputs(5711) <= not b or a;
    layer0_outputs(5712) <= a and b;
    layer0_outputs(5713) <= not a;
    layer0_outputs(5714) <= '1';
    layer0_outputs(5715) <= a and not b;
    layer0_outputs(5716) <= b;
    layer0_outputs(5717) <= not a;
    layer0_outputs(5718) <= not (a or b);
    layer0_outputs(5719) <= not (a or b);
    layer0_outputs(5720) <= not (a and b);
    layer0_outputs(5721) <= b and not a;
    layer0_outputs(5722) <= not a or b;
    layer0_outputs(5723) <= a and b;
    layer0_outputs(5724) <= not (a xor b);
    layer0_outputs(5725) <= not b;
    layer0_outputs(5726) <= a or b;
    layer0_outputs(5727) <= a and not b;
    layer0_outputs(5728) <= a or b;
    layer0_outputs(5729) <= b and not a;
    layer0_outputs(5730) <= a xor b;
    layer0_outputs(5731) <= '0';
    layer0_outputs(5732) <= not (a or b);
    layer0_outputs(5733) <= not (a xor b);
    layer0_outputs(5734) <= a xor b;
    layer0_outputs(5735) <= not b;
    layer0_outputs(5736) <= a or b;
    layer0_outputs(5737) <= not (a xor b);
    layer0_outputs(5738) <= b and not a;
    layer0_outputs(5739) <= a;
    layer0_outputs(5740) <= b;
    layer0_outputs(5741) <= '1';
    layer0_outputs(5742) <= not b;
    layer0_outputs(5743) <= a or b;
    layer0_outputs(5744) <= not (a and b);
    layer0_outputs(5745) <= a or b;
    layer0_outputs(5746) <= a xor b;
    layer0_outputs(5747) <= b;
    layer0_outputs(5748) <= not (a xor b);
    layer0_outputs(5749) <= not (a xor b);
    layer0_outputs(5750) <= not (a xor b);
    layer0_outputs(5751) <= a and b;
    layer0_outputs(5752) <= not (a or b);
    layer0_outputs(5753) <= not a;
    layer0_outputs(5754) <= a or b;
    layer0_outputs(5755) <= a or b;
    layer0_outputs(5756) <= not a;
    layer0_outputs(5757) <= a xor b;
    layer0_outputs(5758) <= not (a or b);
    layer0_outputs(5759) <= not b or a;
    layer0_outputs(5760) <= not b;
    layer0_outputs(5761) <= b and not a;
    layer0_outputs(5762) <= a or b;
    layer0_outputs(5763) <= b;
    layer0_outputs(5764) <= a xor b;
    layer0_outputs(5765) <= not a;
    layer0_outputs(5766) <= b;
    layer0_outputs(5767) <= not (a or b);
    layer0_outputs(5768) <= not (a or b);
    layer0_outputs(5769) <= a and not b;
    layer0_outputs(5770) <= '0';
    layer0_outputs(5771) <= a or b;
    layer0_outputs(5772) <= a or b;
    layer0_outputs(5773) <= b;
    layer0_outputs(5774) <= a;
    layer0_outputs(5775) <= b and not a;
    layer0_outputs(5776) <= not a or b;
    layer0_outputs(5777) <= b;
    layer0_outputs(5778) <= not b or a;
    layer0_outputs(5779) <= not (a or b);
    layer0_outputs(5780) <= a or b;
    layer0_outputs(5781) <= a or b;
    layer0_outputs(5782) <= a xor b;
    layer0_outputs(5783) <= not (a xor b);
    layer0_outputs(5784) <= not a or b;
    layer0_outputs(5785) <= not a or b;
    layer0_outputs(5786) <= a and not b;
    layer0_outputs(5787) <= not a;
    layer0_outputs(5788) <= a or b;
    layer0_outputs(5789) <= a and b;
    layer0_outputs(5790) <= not (a or b);
    layer0_outputs(5791) <= a or b;
    layer0_outputs(5792) <= not a;
    layer0_outputs(5793) <= not a or b;
    layer0_outputs(5794) <= not (a or b);
    layer0_outputs(5795) <= not b or a;
    layer0_outputs(5796) <= not (a xor b);
    layer0_outputs(5797) <= not a;
    layer0_outputs(5798) <= a or b;
    layer0_outputs(5799) <= a;
    layer0_outputs(5800) <= not b;
    layer0_outputs(5801) <= not (a xor b);
    layer0_outputs(5802) <= b;
    layer0_outputs(5803) <= a and not b;
    layer0_outputs(5804) <= not (a xor b);
    layer0_outputs(5805) <= '0';
    layer0_outputs(5806) <= not b;
    layer0_outputs(5807) <= b and not a;
    layer0_outputs(5808) <= b and not a;
    layer0_outputs(5809) <= not a;
    layer0_outputs(5810) <= '1';
    layer0_outputs(5811) <= not (a or b);
    layer0_outputs(5812) <= b and not a;
    layer0_outputs(5813) <= b;
    layer0_outputs(5814) <= not a;
    layer0_outputs(5815) <= not a or b;
    layer0_outputs(5816) <= b and not a;
    layer0_outputs(5817) <= not b or a;
    layer0_outputs(5818) <= b and not a;
    layer0_outputs(5819) <= not a or b;
    layer0_outputs(5820) <= not b;
    layer0_outputs(5821) <= b;
    layer0_outputs(5822) <= a or b;
    layer0_outputs(5823) <= not b or a;
    layer0_outputs(5824) <= not (a xor b);
    layer0_outputs(5825) <= a and b;
    layer0_outputs(5826) <= not (a or b);
    layer0_outputs(5827) <= not (a or b);
    layer0_outputs(5828) <= not a;
    layer0_outputs(5829) <= b and not a;
    layer0_outputs(5830) <= b and not a;
    layer0_outputs(5831) <= not a;
    layer0_outputs(5832) <= not (a and b);
    layer0_outputs(5833) <= not (a xor b);
    layer0_outputs(5834) <= b;
    layer0_outputs(5835) <= b;
    layer0_outputs(5836) <= not (a or b);
    layer0_outputs(5837) <= not a or b;
    layer0_outputs(5838) <= a xor b;
    layer0_outputs(5839) <= b and not a;
    layer0_outputs(5840) <= a and not b;
    layer0_outputs(5841) <= not b or a;
    layer0_outputs(5842) <= a or b;
    layer0_outputs(5843) <= not (a and b);
    layer0_outputs(5844) <= b;
    layer0_outputs(5845) <= not a;
    layer0_outputs(5846) <= a and b;
    layer0_outputs(5847) <= a and not b;
    layer0_outputs(5848) <= not (a or b);
    layer0_outputs(5849) <= not (a xor b);
    layer0_outputs(5850) <= a and b;
    layer0_outputs(5851) <= not b;
    layer0_outputs(5852) <= a;
    layer0_outputs(5853) <= not (a xor b);
    layer0_outputs(5854) <= not b;
    layer0_outputs(5855) <= b;
    layer0_outputs(5856) <= a;
    layer0_outputs(5857) <= not a;
    layer0_outputs(5858) <= b and not a;
    layer0_outputs(5859) <= not (a or b);
    layer0_outputs(5860) <= not (a or b);
    layer0_outputs(5861) <= '0';
    layer0_outputs(5862) <= b;
    layer0_outputs(5863) <= '1';
    layer0_outputs(5864) <= a and not b;
    layer0_outputs(5865) <= not (a xor b);
    layer0_outputs(5866) <= not b;
    layer0_outputs(5867) <= not b or a;
    layer0_outputs(5868) <= not (a xor b);
    layer0_outputs(5869) <= not (a xor b);
    layer0_outputs(5870) <= not a or b;
    layer0_outputs(5871) <= b and not a;
    layer0_outputs(5872) <= not (a xor b);
    layer0_outputs(5873) <= a and not b;
    layer0_outputs(5874) <= a;
    layer0_outputs(5875) <= a xor b;
    layer0_outputs(5876) <= not b or a;
    layer0_outputs(5877) <= a or b;
    layer0_outputs(5878) <= not (a or b);
    layer0_outputs(5879) <= not a;
    layer0_outputs(5880) <= not b;
    layer0_outputs(5881) <= not b;
    layer0_outputs(5882) <= not a;
    layer0_outputs(5883) <= b and not a;
    layer0_outputs(5884) <= b;
    layer0_outputs(5885) <= a or b;
    layer0_outputs(5886) <= b;
    layer0_outputs(5887) <= not a;
    layer0_outputs(5888) <= not (a or b);
    layer0_outputs(5889) <= not b or a;
    layer0_outputs(5890) <= not a or b;
    layer0_outputs(5891) <= not (a xor b);
    layer0_outputs(5892) <= b and not a;
    layer0_outputs(5893) <= not (a or b);
    layer0_outputs(5894) <= not (a and b);
    layer0_outputs(5895) <= not (a xor b);
    layer0_outputs(5896) <= '0';
    layer0_outputs(5897) <= not b or a;
    layer0_outputs(5898) <= a or b;
    layer0_outputs(5899) <= a or b;
    layer0_outputs(5900) <= b and not a;
    layer0_outputs(5901) <= a xor b;
    layer0_outputs(5902) <= '1';
    layer0_outputs(5903) <= not b or a;
    layer0_outputs(5904) <= not b;
    layer0_outputs(5905) <= a and not b;
    layer0_outputs(5906) <= not a;
    layer0_outputs(5907) <= a or b;
    layer0_outputs(5908) <= not a or b;
    layer0_outputs(5909) <= not a;
    layer0_outputs(5910) <= b;
    layer0_outputs(5911) <= not a or b;
    layer0_outputs(5912) <= not (a or b);
    layer0_outputs(5913) <= a xor b;
    layer0_outputs(5914) <= a;
    layer0_outputs(5915) <= a;
    layer0_outputs(5916) <= not b or a;
    layer0_outputs(5917) <= a or b;
    layer0_outputs(5918) <= a xor b;
    layer0_outputs(5919) <= a or b;
    layer0_outputs(5920) <= not a or b;
    layer0_outputs(5921) <= a;
    layer0_outputs(5922) <= a xor b;
    layer0_outputs(5923) <= a and b;
    layer0_outputs(5924) <= a;
    layer0_outputs(5925) <= b and not a;
    layer0_outputs(5926) <= not a;
    layer0_outputs(5927) <= b;
    layer0_outputs(5928) <= not (a xor b);
    layer0_outputs(5929) <= not (a or b);
    layer0_outputs(5930) <= b;
    layer0_outputs(5931) <= a or b;
    layer0_outputs(5932) <= b;
    layer0_outputs(5933) <= b and not a;
    layer0_outputs(5934) <= a xor b;
    layer0_outputs(5935) <= b and not a;
    layer0_outputs(5936) <= not a;
    layer0_outputs(5937) <= not (a xor b);
    layer0_outputs(5938) <= a xor b;
    layer0_outputs(5939) <= not a;
    layer0_outputs(5940) <= not (a or b);
    layer0_outputs(5941) <= not (a or b);
    layer0_outputs(5942) <= not b;
    layer0_outputs(5943) <= not (a xor b);
    layer0_outputs(5944) <= not a or b;
    layer0_outputs(5945) <= a or b;
    layer0_outputs(5946) <= '1';
    layer0_outputs(5947) <= not (a or b);
    layer0_outputs(5948) <= a xor b;
    layer0_outputs(5949) <= not b;
    layer0_outputs(5950) <= a or b;
    layer0_outputs(5951) <= a xor b;
    layer0_outputs(5952) <= not a;
    layer0_outputs(5953) <= a and b;
    layer0_outputs(5954) <= a or b;
    layer0_outputs(5955) <= a or b;
    layer0_outputs(5956) <= not a or b;
    layer0_outputs(5957) <= a or b;
    layer0_outputs(5958) <= b;
    layer0_outputs(5959) <= a or b;
    layer0_outputs(5960) <= not b;
    layer0_outputs(5961) <= not a;
    layer0_outputs(5962) <= a xor b;
    layer0_outputs(5963) <= not (a xor b);
    layer0_outputs(5964) <= not (a or b);
    layer0_outputs(5965) <= not (a or b);
    layer0_outputs(5966) <= not (a and b);
    layer0_outputs(5967) <= a or b;
    layer0_outputs(5968) <= not (a xor b);
    layer0_outputs(5969) <= a;
    layer0_outputs(5970) <= not b;
    layer0_outputs(5971) <= not a;
    layer0_outputs(5972) <= b;
    layer0_outputs(5973) <= a and not b;
    layer0_outputs(5974) <= not (a or b);
    layer0_outputs(5975) <= b and not a;
    layer0_outputs(5976) <= a or b;
    layer0_outputs(5977) <= a;
    layer0_outputs(5978) <= a xor b;
    layer0_outputs(5979) <= a or b;
    layer0_outputs(5980) <= not b;
    layer0_outputs(5981) <= not a;
    layer0_outputs(5982) <= b;
    layer0_outputs(5983) <= a xor b;
    layer0_outputs(5984) <= a xor b;
    layer0_outputs(5985) <= not a or b;
    layer0_outputs(5986) <= a or b;
    layer0_outputs(5987) <= not b or a;
    layer0_outputs(5988) <= not (a and b);
    layer0_outputs(5989) <= b;
    layer0_outputs(5990) <= not (a xor b);
    layer0_outputs(5991) <= not b;
    layer0_outputs(5992) <= not (a xor b);
    layer0_outputs(5993) <= a or b;
    layer0_outputs(5994) <= not a or b;
    layer0_outputs(5995) <= a;
    layer0_outputs(5996) <= b;
    layer0_outputs(5997) <= not a;
    layer0_outputs(5998) <= b and not a;
    layer0_outputs(5999) <= not a;
    layer0_outputs(6000) <= not (a or b);
    layer0_outputs(6001) <= not a;
    layer0_outputs(6002) <= not b or a;
    layer0_outputs(6003) <= a or b;
    layer0_outputs(6004) <= not (a and b);
    layer0_outputs(6005) <= b;
    layer0_outputs(6006) <= not b;
    layer0_outputs(6007) <= not (a or b);
    layer0_outputs(6008) <= a and b;
    layer0_outputs(6009) <= not b or a;
    layer0_outputs(6010) <= a xor b;
    layer0_outputs(6011) <= not a;
    layer0_outputs(6012) <= b and not a;
    layer0_outputs(6013) <= not b;
    layer0_outputs(6014) <= a;
    layer0_outputs(6015) <= not (a and b);
    layer0_outputs(6016) <= not a or b;
    layer0_outputs(6017) <= a;
    layer0_outputs(6018) <= a and not b;
    layer0_outputs(6019) <= b and not a;
    layer0_outputs(6020) <= not a or b;
    layer0_outputs(6021) <= b;
    layer0_outputs(6022) <= a and b;
    layer0_outputs(6023) <= not (a xor b);
    layer0_outputs(6024) <= not b or a;
    layer0_outputs(6025) <= a or b;
    layer0_outputs(6026) <= not a or b;
    layer0_outputs(6027) <= not b or a;
    layer0_outputs(6028) <= a;
    layer0_outputs(6029) <= not a or b;
    layer0_outputs(6030) <= a and not b;
    layer0_outputs(6031) <= not b;
    layer0_outputs(6032) <= not b or a;
    layer0_outputs(6033) <= a;
    layer0_outputs(6034) <= a;
    layer0_outputs(6035) <= b;
    layer0_outputs(6036) <= a;
    layer0_outputs(6037) <= a and b;
    layer0_outputs(6038) <= a or b;
    layer0_outputs(6039) <= not a;
    layer0_outputs(6040) <= not b or a;
    layer0_outputs(6041) <= not b or a;
    layer0_outputs(6042) <= a xor b;
    layer0_outputs(6043) <= a;
    layer0_outputs(6044) <= not (a xor b);
    layer0_outputs(6045) <= a;
    layer0_outputs(6046) <= not b or a;
    layer0_outputs(6047) <= a and not b;
    layer0_outputs(6048) <= not (a or b);
    layer0_outputs(6049) <= a or b;
    layer0_outputs(6050) <= a and not b;
    layer0_outputs(6051) <= a xor b;
    layer0_outputs(6052) <= not b or a;
    layer0_outputs(6053) <= not (a and b);
    layer0_outputs(6054) <= not a or b;
    layer0_outputs(6055) <= not a;
    layer0_outputs(6056) <= a xor b;
    layer0_outputs(6057) <= a and b;
    layer0_outputs(6058) <= a and not b;
    layer0_outputs(6059) <= not b or a;
    layer0_outputs(6060) <= not (a or b);
    layer0_outputs(6061) <= not a;
    layer0_outputs(6062) <= a and b;
    layer0_outputs(6063) <= not a;
    layer0_outputs(6064) <= not (a and b);
    layer0_outputs(6065) <= a or b;
    layer0_outputs(6066) <= not a;
    layer0_outputs(6067) <= not a;
    layer0_outputs(6068) <= not (a or b);
    layer0_outputs(6069) <= not b or a;
    layer0_outputs(6070) <= a and not b;
    layer0_outputs(6071) <= b;
    layer0_outputs(6072) <= not a or b;
    layer0_outputs(6073) <= a;
    layer0_outputs(6074) <= not b;
    layer0_outputs(6075) <= not a;
    layer0_outputs(6076) <= a;
    layer0_outputs(6077) <= not a or b;
    layer0_outputs(6078) <= not b or a;
    layer0_outputs(6079) <= a;
    layer0_outputs(6080) <= a xor b;
    layer0_outputs(6081) <= a and not b;
    layer0_outputs(6082) <= b;
    layer0_outputs(6083) <= a or b;
    layer0_outputs(6084) <= not (a xor b);
    layer0_outputs(6085) <= b;
    layer0_outputs(6086) <= a;
    layer0_outputs(6087) <= not (a or b);
    layer0_outputs(6088) <= a or b;
    layer0_outputs(6089) <= b and not a;
    layer0_outputs(6090) <= a;
    layer0_outputs(6091) <= b;
    layer0_outputs(6092) <= not b;
    layer0_outputs(6093) <= a or b;
    layer0_outputs(6094) <= not a or b;
    layer0_outputs(6095) <= not (a and b);
    layer0_outputs(6096) <= '1';
    layer0_outputs(6097) <= a or b;
    layer0_outputs(6098) <= not b;
    layer0_outputs(6099) <= a and b;
    layer0_outputs(6100) <= b;
    layer0_outputs(6101) <= not a;
    layer0_outputs(6102) <= a xor b;
    layer0_outputs(6103) <= not a;
    layer0_outputs(6104) <= not a;
    layer0_outputs(6105) <= a;
    layer0_outputs(6106) <= not b or a;
    layer0_outputs(6107) <= not (a or b);
    layer0_outputs(6108) <= not b or a;
    layer0_outputs(6109) <= b;
    layer0_outputs(6110) <= a;
    layer0_outputs(6111) <= not (a or b);
    layer0_outputs(6112) <= not a;
    layer0_outputs(6113) <= not (a and b);
    layer0_outputs(6114) <= not b;
    layer0_outputs(6115) <= '0';
    layer0_outputs(6116) <= a or b;
    layer0_outputs(6117) <= not (a and b);
    layer0_outputs(6118) <= not (a or b);
    layer0_outputs(6119) <= '0';
    layer0_outputs(6120) <= b and not a;
    layer0_outputs(6121) <= not (a and b);
    layer0_outputs(6122) <= a xor b;
    layer0_outputs(6123) <= a;
    layer0_outputs(6124) <= a or b;
    layer0_outputs(6125) <= not (a xor b);
    layer0_outputs(6126) <= a and not b;
    layer0_outputs(6127) <= a xor b;
    layer0_outputs(6128) <= a or b;
    layer0_outputs(6129) <= b;
    layer0_outputs(6130) <= not (a xor b);
    layer0_outputs(6131) <= not (a or b);
    layer0_outputs(6132) <= '0';
    layer0_outputs(6133) <= not (a or b);
    layer0_outputs(6134) <= a;
    layer0_outputs(6135) <= not (a xor b);
    layer0_outputs(6136) <= b and not a;
    layer0_outputs(6137) <= a or b;
    layer0_outputs(6138) <= not (a or b);
    layer0_outputs(6139) <= '0';
    layer0_outputs(6140) <= not a;
    layer0_outputs(6141) <= a;
    layer0_outputs(6142) <= not b;
    layer0_outputs(6143) <= not a;
    layer0_outputs(6144) <= not b;
    layer0_outputs(6145) <= a xor b;
    layer0_outputs(6146) <= not a;
    layer0_outputs(6147) <= a;
    layer0_outputs(6148) <= not (a or b);
    layer0_outputs(6149) <= a xor b;
    layer0_outputs(6150) <= not (a xor b);
    layer0_outputs(6151) <= b;
    layer0_outputs(6152) <= not (a or b);
    layer0_outputs(6153) <= not a or b;
    layer0_outputs(6154) <= not (a or b);
    layer0_outputs(6155) <= not b or a;
    layer0_outputs(6156) <= not a;
    layer0_outputs(6157) <= a and b;
    layer0_outputs(6158) <= a or b;
    layer0_outputs(6159) <= b;
    layer0_outputs(6160) <= '1';
    layer0_outputs(6161) <= not a;
    layer0_outputs(6162) <= not a or b;
    layer0_outputs(6163) <= a or b;
    layer0_outputs(6164) <= b;
    layer0_outputs(6165) <= a and not b;
    layer0_outputs(6166) <= not b or a;
    layer0_outputs(6167) <= a and b;
    layer0_outputs(6168) <= not b or a;
    layer0_outputs(6169) <= a xor b;
    layer0_outputs(6170) <= a or b;
    layer0_outputs(6171) <= b and not a;
    layer0_outputs(6172) <= not (a and b);
    layer0_outputs(6173) <= not a;
    layer0_outputs(6174) <= a xor b;
    layer0_outputs(6175) <= not b or a;
    layer0_outputs(6176) <= '1';
    layer0_outputs(6177) <= not b;
    layer0_outputs(6178) <= a and b;
    layer0_outputs(6179) <= not a or b;
    layer0_outputs(6180) <= a and not b;
    layer0_outputs(6181) <= not (a xor b);
    layer0_outputs(6182) <= not (a or b);
    layer0_outputs(6183) <= a xor b;
    layer0_outputs(6184) <= not (a or b);
    layer0_outputs(6185) <= not b or a;
    layer0_outputs(6186) <= not b;
    layer0_outputs(6187) <= a;
    layer0_outputs(6188) <= not a or b;
    layer0_outputs(6189) <= not a;
    layer0_outputs(6190) <= not b;
    layer0_outputs(6191) <= not b or a;
    layer0_outputs(6192) <= not a;
    layer0_outputs(6193) <= not (a xor b);
    layer0_outputs(6194) <= b;
    layer0_outputs(6195) <= '0';
    layer0_outputs(6196) <= a xor b;
    layer0_outputs(6197) <= not a;
    layer0_outputs(6198) <= a;
    layer0_outputs(6199) <= a or b;
    layer0_outputs(6200) <= not (a xor b);
    layer0_outputs(6201) <= not (a or b);
    layer0_outputs(6202) <= a;
    layer0_outputs(6203) <= a or b;
    layer0_outputs(6204) <= not (a or b);
    layer0_outputs(6205) <= b and not a;
    layer0_outputs(6206) <= a and not b;
    layer0_outputs(6207) <= a and b;
    layer0_outputs(6208) <= b and not a;
    layer0_outputs(6209) <= a or b;
    layer0_outputs(6210) <= not (a or b);
    layer0_outputs(6211) <= a xor b;
    layer0_outputs(6212) <= b;
    layer0_outputs(6213) <= b and not a;
    layer0_outputs(6214) <= a;
    layer0_outputs(6215) <= not b or a;
    layer0_outputs(6216) <= b;
    layer0_outputs(6217) <= not (a or b);
    layer0_outputs(6218) <= not (a or b);
    layer0_outputs(6219) <= not b or a;
    layer0_outputs(6220) <= a or b;
    layer0_outputs(6221) <= not a;
    layer0_outputs(6222) <= '0';
    layer0_outputs(6223) <= not b;
    layer0_outputs(6224) <= b and not a;
    layer0_outputs(6225) <= a;
    layer0_outputs(6226) <= a and not b;
    layer0_outputs(6227) <= a and b;
    layer0_outputs(6228) <= not (a or b);
    layer0_outputs(6229) <= not b;
    layer0_outputs(6230) <= not a or b;
    layer0_outputs(6231) <= b;
    layer0_outputs(6232) <= a or b;
    layer0_outputs(6233) <= not b;
    layer0_outputs(6234) <= a or b;
    layer0_outputs(6235) <= a;
    layer0_outputs(6236) <= not a;
    layer0_outputs(6237) <= not b or a;
    layer0_outputs(6238) <= a or b;
    layer0_outputs(6239) <= b and not a;
    layer0_outputs(6240) <= b and not a;
    layer0_outputs(6241) <= not a or b;
    layer0_outputs(6242) <= not b;
    layer0_outputs(6243) <= a or b;
    layer0_outputs(6244) <= a and not b;
    layer0_outputs(6245) <= not a;
    layer0_outputs(6246) <= not b;
    layer0_outputs(6247) <= not b or a;
    layer0_outputs(6248) <= not (a xor b);
    layer0_outputs(6249) <= b;
    layer0_outputs(6250) <= not (a or b);
    layer0_outputs(6251) <= a or b;
    layer0_outputs(6252) <= b and not a;
    layer0_outputs(6253) <= a or b;
    layer0_outputs(6254) <= a or b;
    layer0_outputs(6255) <= not (a and b);
    layer0_outputs(6256) <= a or b;
    layer0_outputs(6257) <= not (a or b);
    layer0_outputs(6258) <= not a or b;
    layer0_outputs(6259) <= a or b;
    layer0_outputs(6260) <= a or b;
    layer0_outputs(6261) <= not (a xor b);
    layer0_outputs(6262) <= not (a and b);
    layer0_outputs(6263) <= b;
    layer0_outputs(6264) <= not b or a;
    layer0_outputs(6265) <= b and not a;
    layer0_outputs(6266) <= a or b;
    layer0_outputs(6267) <= not b;
    layer0_outputs(6268) <= '0';
    layer0_outputs(6269) <= b and not a;
    layer0_outputs(6270) <= a;
    layer0_outputs(6271) <= a xor b;
    layer0_outputs(6272) <= b;
    layer0_outputs(6273) <= a;
    layer0_outputs(6274) <= a xor b;
    layer0_outputs(6275) <= a or b;
    layer0_outputs(6276) <= not a;
    layer0_outputs(6277) <= not b or a;
    layer0_outputs(6278) <= not b;
    layer0_outputs(6279) <= a and not b;
    layer0_outputs(6280) <= b and not a;
    layer0_outputs(6281) <= not a or b;
    layer0_outputs(6282) <= not b;
    layer0_outputs(6283) <= b;
    layer0_outputs(6284) <= not (a and b);
    layer0_outputs(6285) <= not (a and b);
    layer0_outputs(6286) <= a or b;
    layer0_outputs(6287) <= a xor b;
    layer0_outputs(6288) <= not (a xor b);
    layer0_outputs(6289) <= not (a or b);
    layer0_outputs(6290) <= a or b;
    layer0_outputs(6291) <= b;
    layer0_outputs(6292) <= a or b;
    layer0_outputs(6293) <= a and not b;
    layer0_outputs(6294) <= a and b;
    layer0_outputs(6295) <= not (a or b);
    layer0_outputs(6296) <= not (a and b);
    layer0_outputs(6297) <= not (a and b);
    layer0_outputs(6298) <= a;
    layer0_outputs(6299) <= a or b;
    layer0_outputs(6300) <= '0';
    layer0_outputs(6301) <= a;
    layer0_outputs(6302) <= a or b;
    layer0_outputs(6303) <= a;
    layer0_outputs(6304) <= a xor b;
    layer0_outputs(6305) <= a and not b;
    layer0_outputs(6306) <= a or b;
    layer0_outputs(6307) <= not (a and b);
    layer0_outputs(6308) <= not a or b;
    layer0_outputs(6309) <= not a or b;
    layer0_outputs(6310) <= not (a or b);
    layer0_outputs(6311) <= b;
    layer0_outputs(6312) <= not (a xor b);
    layer0_outputs(6313) <= not (a or b);
    layer0_outputs(6314) <= not a;
    layer0_outputs(6315) <= a;
    layer0_outputs(6316) <= b and not a;
    layer0_outputs(6317) <= not (a or b);
    layer0_outputs(6318) <= not b or a;
    layer0_outputs(6319) <= b;
    layer0_outputs(6320) <= not b;
    layer0_outputs(6321) <= not a or b;
    layer0_outputs(6322) <= not b;
    layer0_outputs(6323) <= not b;
    layer0_outputs(6324) <= b;
    layer0_outputs(6325) <= b and not a;
    layer0_outputs(6326) <= not (a or b);
    layer0_outputs(6327) <= a;
    layer0_outputs(6328) <= not a;
    layer0_outputs(6329) <= b;
    layer0_outputs(6330) <= a xor b;
    layer0_outputs(6331) <= '1';
    layer0_outputs(6332) <= not (a and b);
    layer0_outputs(6333) <= not a;
    layer0_outputs(6334) <= not a;
    layer0_outputs(6335) <= b and not a;
    layer0_outputs(6336) <= a or b;
    layer0_outputs(6337) <= a xor b;
    layer0_outputs(6338) <= not a or b;
    layer0_outputs(6339) <= not b;
    layer0_outputs(6340) <= a;
    layer0_outputs(6341) <= a or b;
    layer0_outputs(6342) <= not b;
    layer0_outputs(6343) <= a xor b;
    layer0_outputs(6344) <= not (a or b);
    layer0_outputs(6345) <= b;
    layer0_outputs(6346) <= b;
    layer0_outputs(6347) <= a xor b;
    layer0_outputs(6348) <= a or b;
    layer0_outputs(6349) <= not (a or b);
    layer0_outputs(6350) <= a and b;
    layer0_outputs(6351) <= not (a xor b);
    layer0_outputs(6352) <= not (a or b);
    layer0_outputs(6353) <= a and not b;
    layer0_outputs(6354) <= a and b;
    layer0_outputs(6355) <= a or b;
    layer0_outputs(6356) <= a and not b;
    layer0_outputs(6357) <= a or b;
    layer0_outputs(6358) <= a or b;
    layer0_outputs(6359) <= not (a or b);
    layer0_outputs(6360) <= a;
    layer0_outputs(6361) <= a or b;
    layer0_outputs(6362) <= b and not a;
    layer0_outputs(6363) <= not (a or b);
    layer0_outputs(6364) <= not (a xor b);
    layer0_outputs(6365) <= a xor b;
    layer0_outputs(6366) <= b;
    layer0_outputs(6367) <= b and not a;
    layer0_outputs(6368) <= b and not a;
    layer0_outputs(6369) <= not (a or b);
    layer0_outputs(6370) <= a or b;
    layer0_outputs(6371) <= a and b;
    layer0_outputs(6372) <= b;
    layer0_outputs(6373) <= not a or b;
    layer0_outputs(6374) <= a;
    layer0_outputs(6375) <= a or b;
    layer0_outputs(6376) <= b;
    layer0_outputs(6377) <= '1';
    layer0_outputs(6378) <= not b or a;
    layer0_outputs(6379) <= not b;
    layer0_outputs(6380) <= b and not a;
    layer0_outputs(6381) <= a xor b;
    layer0_outputs(6382) <= not b;
    layer0_outputs(6383) <= b and not a;
    layer0_outputs(6384) <= not (a or b);
    layer0_outputs(6385) <= b and not a;
    layer0_outputs(6386) <= not b;
    layer0_outputs(6387) <= a or b;
    layer0_outputs(6388) <= a xor b;
    layer0_outputs(6389) <= b;
    layer0_outputs(6390) <= a or b;
    layer0_outputs(6391) <= a or b;
    layer0_outputs(6392) <= not (a or b);
    layer0_outputs(6393) <= not (a and b);
    layer0_outputs(6394) <= not (a or b);
    layer0_outputs(6395) <= '1';
    layer0_outputs(6396) <= a xor b;
    layer0_outputs(6397) <= not a;
    layer0_outputs(6398) <= a xor b;
    layer0_outputs(6399) <= not (a or b);
    layer0_outputs(6400) <= a and b;
    layer0_outputs(6401) <= b and not a;
    layer0_outputs(6402) <= b and not a;
    layer0_outputs(6403) <= not (a xor b);
    layer0_outputs(6404) <= a and not b;
    layer0_outputs(6405) <= b and not a;
    layer0_outputs(6406) <= not b;
    layer0_outputs(6407) <= not (a and b);
    layer0_outputs(6408) <= not (a or b);
    layer0_outputs(6409) <= b;
    layer0_outputs(6410) <= a and not b;
    layer0_outputs(6411) <= not a;
    layer0_outputs(6412) <= not (a and b);
    layer0_outputs(6413) <= a and not b;
    layer0_outputs(6414) <= a;
    layer0_outputs(6415) <= not (a or b);
    layer0_outputs(6416) <= a and not b;
    layer0_outputs(6417) <= not b or a;
    layer0_outputs(6418) <= a xor b;
    layer0_outputs(6419) <= not (a or b);
    layer0_outputs(6420) <= not b or a;
    layer0_outputs(6421) <= not a or b;
    layer0_outputs(6422) <= not (a or b);
    layer0_outputs(6423) <= a xor b;
    layer0_outputs(6424) <= not b;
    layer0_outputs(6425) <= '0';
    layer0_outputs(6426) <= not (a and b);
    layer0_outputs(6427) <= not (a xor b);
    layer0_outputs(6428) <= b;
    layer0_outputs(6429) <= a and b;
    layer0_outputs(6430) <= a xor b;
    layer0_outputs(6431) <= not (a or b);
    layer0_outputs(6432) <= a or b;
    layer0_outputs(6433) <= not b;
    layer0_outputs(6434) <= not b;
    layer0_outputs(6435) <= not a or b;
    layer0_outputs(6436) <= a and not b;
    layer0_outputs(6437) <= b and not a;
    layer0_outputs(6438) <= not (a xor b);
    layer0_outputs(6439) <= b and not a;
    layer0_outputs(6440) <= not b or a;
    layer0_outputs(6441) <= '1';
    layer0_outputs(6442) <= not (a or b);
    layer0_outputs(6443) <= a and b;
    layer0_outputs(6444) <= not a;
    layer0_outputs(6445) <= not a or b;
    layer0_outputs(6446) <= not b;
    layer0_outputs(6447) <= not a;
    layer0_outputs(6448) <= a and not b;
    layer0_outputs(6449) <= a;
    layer0_outputs(6450) <= b and not a;
    layer0_outputs(6451) <= not a;
    layer0_outputs(6452) <= a or b;
    layer0_outputs(6453) <= b and not a;
    layer0_outputs(6454) <= not (a or b);
    layer0_outputs(6455) <= a or b;
    layer0_outputs(6456) <= not b;
    layer0_outputs(6457) <= '1';
    layer0_outputs(6458) <= not b or a;
    layer0_outputs(6459) <= a xor b;
    layer0_outputs(6460) <= a or b;
    layer0_outputs(6461) <= a and b;
    layer0_outputs(6462) <= not (a and b);
    layer0_outputs(6463) <= '0';
    layer0_outputs(6464) <= not b or a;
    layer0_outputs(6465) <= not a;
    layer0_outputs(6466) <= not (a or b);
    layer0_outputs(6467) <= '0';
    layer0_outputs(6468) <= a xor b;
    layer0_outputs(6469) <= '1';
    layer0_outputs(6470) <= a xor b;
    layer0_outputs(6471) <= a;
    layer0_outputs(6472) <= not b;
    layer0_outputs(6473) <= not a or b;
    layer0_outputs(6474) <= a and b;
    layer0_outputs(6475) <= not (a or b);
    layer0_outputs(6476) <= not (a or b);
    layer0_outputs(6477) <= not a or b;
    layer0_outputs(6478) <= a xor b;
    layer0_outputs(6479) <= b;
    layer0_outputs(6480) <= not b;
    layer0_outputs(6481) <= '1';
    layer0_outputs(6482) <= not (a or b);
    layer0_outputs(6483) <= a xor b;
    layer0_outputs(6484) <= not (a and b);
    layer0_outputs(6485) <= not a or b;
    layer0_outputs(6486) <= not (a or b);
    layer0_outputs(6487) <= a;
    layer0_outputs(6488) <= not a;
    layer0_outputs(6489) <= a and not b;
    layer0_outputs(6490) <= a;
    layer0_outputs(6491) <= not (a or b);
    layer0_outputs(6492) <= a;
    layer0_outputs(6493) <= not (a or b);
    layer0_outputs(6494) <= a and not b;
    layer0_outputs(6495) <= not a or b;
    layer0_outputs(6496) <= not a or b;
    layer0_outputs(6497) <= not (a xor b);
    layer0_outputs(6498) <= a or b;
    layer0_outputs(6499) <= not (a or b);
    layer0_outputs(6500) <= b;
    layer0_outputs(6501) <= a or b;
    layer0_outputs(6502) <= not (a or b);
    layer0_outputs(6503) <= not a or b;
    layer0_outputs(6504) <= not (a or b);
    layer0_outputs(6505) <= not b or a;
    layer0_outputs(6506) <= not a or b;
    layer0_outputs(6507) <= a;
    layer0_outputs(6508) <= not a or b;
    layer0_outputs(6509) <= not b or a;
    layer0_outputs(6510) <= not (a and b);
    layer0_outputs(6511) <= not b or a;
    layer0_outputs(6512) <= a and b;
    layer0_outputs(6513) <= not a;
    layer0_outputs(6514) <= a or b;
    layer0_outputs(6515) <= not a;
    layer0_outputs(6516) <= a xor b;
    layer0_outputs(6517) <= a and not b;
    layer0_outputs(6518) <= not (a or b);
    layer0_outputs(6519) <= '0';
    layer0_outputs(6520) <= not (a or b);
    layer0_outputs(6521) <= a and not b;
    layer0_outputs(6522) <= a;
    layer0_outputs(6523) <= not b;
    layer0_outputs(6524) <= a and not b;
    layer0_outputs(6525) <= a and b;
    layer0_outputs(6526) <= a and b;
    layer0_outputs(6527) <= not (a or b);
    layer0_outputs(6528) <= not a or b;
    layer0_outputs(6529) <= not (a or b);
    layer0_outputs(6530) <= a;
    layer0_outputs(6531) <= a;
    layer0_outputs(6532) <= a or b;
    layer0_outputs(6533) <= not (a or b);
    layer0_outputs(6534) <= not a or b;
    layer0_outputs(6535) <= not (a and b);
    layer0_outputs(6536) <= not (a xor b);
    layer0_outputs(6537) <= not (a xor b);
    layer0_outputs(6538) <= b and not a;
    layer0_outputs(6539) <= a xor b;
    layer0_outputs(6540) <= a xor b;
    layer0_outputs(6541) <= not (a or b);
    layer0_outputs(6542) <= not a;
    layer0_outputs(6543) <= not a or b;
    layer0_outputs(6544) <= b and not a;
    layer0_outputs(6545) <= a or b;
    layer0_outputs(6546) <= not (a xor b);
    layer0_outputs(6547) <= not (a xor b);
    layer0_outputs(6548) <= a or b;
    layer0_outputs(6549) <= '1';
    layer0_outputs(6550) <= not a or b;
    layer0_outputs(6551) <= not b or a;
    layer0_outputs(6552) <= a xor b;
    layer0_outputs(6553) <= not a;
    layer0_outputs(6554) <= '1';
    layer0_outputs(6555) <= not b or a;
    layer0_outputs(6556) <= a;
    layer0_outputs(6557) <= not a;
    layer0_outputs(6558) <= b;
    layer0_outputs(6559) <= '1';
    layer0_outputs(6560) <= '1';
    layer0_outputs(6561) <= not (a or b);
    layer0_outputs(6562) <= not (a and b);
    layer0_outputs(6563) <= not b;
    layer0_outputs(6564) <= b;
    layer0_outputs(6565) <= not (a xor b);
    layer0_outputs(6566) <= a xor b;
    layer0_outputs(6567) <= not a;
    layer0_outputs(6568) <= not b;
    layer0_outputs(6569) <= not b or a;
    layer0_outputs(6570) <= a and not b;
    layer0_outputs(6571) <= a xor b;
    layer0_outputs(6572) <= not b or a;
    layer0_outputs(6573) <= a or b;
    layer0_outputs(6574) <= b;
    layer0_outputs(6575) <= b and not a;
    layer0_outputs(6576) <= a xor b;
    layer0_outputs(6577) <= a or b;
    layer0_outputs(6578) <= not b;
    layer0_outputs(6579) <= not (a xor b);
    layer0_outputs(6580) <= b and not a;
    layer0_outputs(6581) <= not a or b;
    layer0_outputs(6582) <= not (a and b);
    layer0_outputs(6583) <= not b or a;
    layer0_outputs(6584) <= not (a or b);
    layer0_outputs(6585) <= not a or b;
    layer0_outputs(6586) <= a xor b;
    layer0_outputs(6587) <= a xor b;
    layer0_outputs(6588) <= b;
    layer0_outputs(6589) <= a xor b;
    layer0_outputs(6590) <= a xor b;
    layer0_outputs(6591) <= a or b;
    layer0_outputs(6592) <= not (a xor b);
    layer0_outputs(6593) <= a and not b;
    layer0_outputs(6594) <= a xor b;
    layer0_outputs(6595) <= b and not a;
    layer0_outputs(6596) <= a xor b;
    layer0_outputs(6597) <= not b;
    layer0_outputs(6598) <= not (a or b);
    layer0_outputs(6599) <= not (a or b);
    layer0_outputs(6600) <= not b;
    layer0_outputs(6601) <= b;
    layer0_outputs(6602) <= not (a or b);
    layer0_outputs(6603) <= b;
    layer0_outputs(6604) <= not a;
    layer0_outputs(6605) <= not (a or b);
    layer0_outputs(6606) <= a xor b;
    layer0_outputs(6607) <= not a;
    layer0_outputs(6608) <= a;
    layer0_outputs(6609) <= a or b;
    layer0_outputs(6610) <= not (a or b);
    layer0_outputs(6611) <= a;
    layer0_outputs(6612) <= a;
    layer0_outputs(6613) <= b;
    layer0_outputs(6614) <= a and b;
    layer0_outputs(6615) <= a or b;
    layer0_outputs(6616) <= not b or a;
    layer0_outputs(6617) <= a;
    layer0_outputs(6618) <= not b;
    layer0_outputs(6619) <= not (a or b);
    layer0_outputs(6620) <= a and b;
    layer0_outputs(6621) <= a or b;
    layer0_outputs(6622) <= not a or b;
    layer0_outputs(6623) <= not (a xor b);
    layer0_outputs(6624) <= a or b;
    layer0_outputs(6625) <= b and not a;
    layer0_outputs(6626) <= a;
    layer0_outputs(6627) <= not (a xor b);
    layer0_outputs(6628) <= a;
    layer0_outputs(6629) <= b and not a;
    layer0_outputs(6630) <= b;
    layer0_outputs(6631) <= a xor b;
    layer0_outputs(6632) <= a and b;
    layer0_outputs(6633) <= not (a or b);
    layer0_outputs(6634) <= not a;
    layer0_outputs(6635) <= a and b;
    layer0_outputs(6636) <= not a or b;
    layer0_outputs(6637) <= not a or b;
    layer0_outputs(6638) <= '1';
    layer0_outputs(6639) <= b and not a;
    layer0_outputs(6640) <= b;
    layer0_outputs(6641) <= a xor b;
    layer0_outputs(6642) <= not a;
    layer0_outputs(6643) <= a or b;
    layer0_outputs(6644) <= not (a or b);
    layer0_outputs(6645) <= a and b;
    layer0_outputs(6646) <= a and not b;
    layer0_outputs(6647) <= not b;
    layer0_outputs(6648) <= not (a or b);
    layer0_outputs(6649) <= not b;
    layer0_outputs(6650) <= a or b;
    layer0_outputs(6651) <= '1';
    layer0_outputs(6652) <= not (a xor b);
    layer0_outputs(6653) <= not a or b;
    layer0_outputs(6654) <= not a;
    layer0_outputs(6655) <= not b or a;
    layer0_outputs(6656) <= a;
    layer0_outputs(6657) <= a or b;
    layer0_outputs(6658) <= not b;
    layer0_outputs(6659) <= b;
    layer0_outputs(6660) <= '1';
    layer0_outputs(6661) <= a or b;
    layer0_outputs(6662) <= a or b;
    layer0_outputs(6663) <= not (a xor b);
    layer0_outputs(6664) <= b;
    layer0_outputs(6665) <= b;
    layer0_outputs(6666) <= a xor b;
    layer0_outputs(6667) <= a;
    layer0_outputs(6668) <= not (a or b);
    layer0_outputs(6669) <= not (a xor b);
    layer0_outputs(6670) <= not (a and b);
    layer0_outputs(6671) <= not a or b;
    layer0_outputs(6672) <= a xor b;
    layer0_outputs(6673) <= not b or a;
    layer0_outputs(6674) <= not b;
    layer0_outputs(6675) <= a and not b;
    layer0_outputs(6676) <= not (a xor b);
    layer0_outputs(6677) <= a or b;
    layer0_outputs(6678) <= not a or b;
    layer0_outputs(6679) <= not (a xor b);
    layer0_outputs(6680) <= '0';
    layer0_outputs(6681) <= not (a or b);
    layer0_outputs(6682) <= a;
    layer0_outputs(6683) <= not (a or b);
    layer0_outputs(6684) <= a or b;
    layer0_outputs(6685) <= a xor b;
    layer0_outputs(6686) <= a and not b;
    layer0_outputs(6687) <= not (a xor b);
    layer0_outputs(6688) <= not a;
    layer0_outputs(6689) <= b;
    layer0_outputs(6690) <= not (a and b);
    layer0_outputs(6691) <= not b or a;
    layer0_outputs(6692) <= not b or a;
    layer0_outputs(6693) <= not (a or b);
    layer0_outputs(6694) <= not a;
    layer0_outputs(6695) <= a xor b;
    layer0_outputs(6696) <= not b;
    layer0_outputs(6697) <= not (a xor b);
    layer0_outputs(6698) <= not a;
    layer0_outputs(6699) <= a xor b;
    layer0_outputs(6700) <= not b or a;
    layer0_outputs(6701) <= a and b;
    layer0_outputs(6702) <= a;
    layer0_outputs(6703) <= not (a xor b);
    layer0_outputs(6704) <= not (a xor b);
    layer0_outputs(6705) <= '1';
    layer0_outputs(6706) <= not (a or b);
    layer0_outputs(6707) <= a and b;
    layer0_outputs(6708) <= not (a or b);
    layer0_outputs(6709) <= a xor b;
    layer0_outputs(6710) <= not a or b;
    layer0_outputs(6711) <= '1';
    layer0_outputs(6712) <= a or b;
    layer0_outputs(6713) <= not (a xor b);
    layer0_outputs(6714) <= b;
    layer0_outputs(6715) <= a and not b;
    layer0_outputs(6716) <= b;
    layer0_outputs(6717) <= not (a xor b);
    layer0_outputs(6718) <= a xor b;
    layer0_outputs(6719) <= a or b;
    layer0_outputs(6720) <= '0';
    layer0_outputs(6721) <= '0';
    layer0_outputs(6722) <= a and not b;
    layer0_outputs(6723) <= a or b;
    layer0_outputs(6724) <= a and b;
    layer0_outputs(6725) <= '0';
    layer0_outputs(6726) <= not a;
    layer0_outputs(6727) <= not a or b;
    layer0_outputs(6728) <= a;
    layer0_outputs(6729) <= not b or a;
    layer0_outputs(6730) <= not (a xor b);
    layer0_outputs(6731) <= not (a xor b);
    layer0_outputs(6732) <= a and not b;
    layer0_outputs(6733) <= a or b;
    layer0_outputs(6734) <= not (a xor b);
    layer0_outputs(6735) <= a or b;
    layer0_outputs(6736) <= a and not b;
    layer0_outputs(6737) <= b and not a;
    layer0_outputs(6738) <= a;
    layer0_outputs(6739) <= not b;
    layer0_outputs(6740) <= '1';
    layer0_outputs(6741) <= a;
    layer0_outputs(6742) <= not (a or b);
    layer0_outputs(6743) <= a and b;
    layer0_outputs(6744) <= not (a or b);
    layer0_outputs(6745) <= a;
    layer0_outputs(6746) <= a or b;
    layer0_outputs(6747) <= not b;
    layer0_outputs(6748) <= not (a or b);
    layer0_outputs(6749) <= not b or a;
    layer0_outputs(6750) <= not a;
    layer0_outputs(6751) <= b and not a;
    layer0_outputs(6752) <= not b or a;
    layer0_outputs(6753) <= a;
    layer0_outputs(6754) <= a xor b;
    layer0_outputs(6755) <= a and not b;
    layer0_outputs(6756) <= a and not b;
    layer0_outputs(6757) <= a;
    layer0_outputs(6758) <= not (a or b);
    layer0_outputs(6759) <= not (a xor b);
    layer0_outputs(6760) <= b;
    layer0_outputs(6761) <= a or b;
    layer0_outputs(6762) <= not (a xor b);
    layer0_outputs(6763) <= not (a or b);
    layer0_outputs(6764) <= not a;
    layer0_outputs(6765) <= a or b;
    layer0_outputs(6766) <= b;
    layer0_outputs(6767) <= not a;
    layer0_outputs(6768) <= not (a or b);
    layer0_outputs(6769) <= not (a and b);
    layer0_outputs(6770) <= a or b;
    layer0_outputs(6771) <= not (a or b);
    layer0_outputs(6772) <= not b or a;
    layer0_outputs(6773) <= not b;
    layer0_outputs(6774) <= b and not a;
    layer0_outputs(6775) <= '1';
    layer0_outputs(6776) <= a or b;
    layer0_outputs(6777) <= not (a xor b);
    layer0_outputs(6778) <= not b or a;
    layer0_outputs(6779) <= a xor b;
    layer0_outputs(6780) <= not (a or b);
    layer0_outputs(6781) <= not a;
    layer0_outputs(6782) <= a or b;
    layer0_outputs(6783) <= a or b;
    layer0_outputs(6784) <= a or b;
    layer0_outputs(6785) <= not (a or b);
    layer0_outputs(6786) <= not (a or b);
    layer0_outputs(6787) <= not (a xor b);
    layer0_outputs(6788) <= not b or a;
    layer0_outputs(6789) <= not (a xor b);
    layer0_outputs(6790) <= a;
    layer0_outputs(6791) <= a xor b;
    layer0_outputs(6792) <= not (a or b);
    layer0_outputs(6793) <= not b or a;
    layer0_outputs(6794) <= a xor b;
    layer0_outputs(6795) <= a or b;
    layer0_outputs(6796) <= not a or b;
    layer0_outputs(6797) <= a or b;
    layer0_outputs(6798) <= not a;
    layer0_outputs(6799) <= b and not a;
    layer0_outputs(6800) <= not (a and b);
    layer0_outputs(6801) <= b and not a;
    layer0_outputs(6802) <= a;
    layer0_outputs(6803) <= not (a xor b);
    layer0_outputs(6804) <= b and not a;
    layer0_outputs(6805) <= a and not b;
    layer0_outputs(6806) <= a and b;
    layer0_outputs(6807) <= a and not b;
    layer0_outputs(6808) <= b and not a;
    layer0_outputs(6809) <= not (a xor b);
    layer0_outputs(6810) <= a;
    layer0_outputs(6811) <= a or b;
    layer0_outputs(6812) <= not (a or b);
    layer0_outputs(6813) <= b;
    layer0_outputs(6814) <= not (a or b);
    layer0_outputs(6815) <= not b;
    layer0_outputs(6816) <= a or b;
    layer0_outputs(6817) <= a;
    layer0_outputs(6818) <= not a or b;
    layer0_outputs(6819) <= a and b;
    layer0_outputs(6820) <= a or b;
    layer0_outputs(6821) <= b;
    layer0_outputs(6822) <= a;
    layer0_outputs(6823) <= a and not b;
    layer0_outputs(6824) <= a and not b;
    layer0_outputs(6825) <= not (a or b);
    layer0_outputs(6826) <= not b or a;
    layer0_outputs(6827) <= '0';
    layer0_outputs(6828) <= '0';
    layer0_outputs(6829) <= not (a or b);
    layer0_outputs(6830) <= not a;
    layer0_outputs(6831) <= b and not a;
    layer0_outputs(6832) <= not a;
    layer0_outputs(6833) <= not b;
    layer0_outputs(6834) <= b and not a;
    layer0_outputs(6835) <= not (a xor b);
    layer0_outputs(6836) <= b;
    layer0_outputs(6837) <= a or b;
    layer0_outputs(6838) <= not (a xor b);
    layer0_outputs(6839) <= a;
    layer0_outputs(6840) <= not a or b;
    layer0_outputs(6841) <= a and not b;
    layer0_outputs(6842) <= a or b;
    layer0_outputs(6843) <= a or b;
    layer0_outputs(6844) <= '0';
    layer0_outputs(6845) <= not (a and b);
    layer0_outputs(6846) <= not b;
    layer0_outputs(6847) <= a and not b;
    layer0_outputs(6848) <= not a or b;
    layer0_outputs(6849) <= not (a xor b);
    layer0_outputs(6850) <= not (a xor b);
    layer0_outputs(6851) <= a xor b;
    layer0_outputs(6852) <= '1';
    layer0_outputs(6853) <= a xor b;
    layer0_outputs(6854) <= a or b;
    layer0_outputs(6855) <= not b;
    layer0_outputs(6856) <= '1';
    layer0_outputs(6857) <= not b or a;
    layer0_outputs(6858) <= not b or a;
    layer0_outputs(6859) <= a or b;
    layer0_outputs(6860) <= not a;
    layer0_outputs(6861) <= not (a or b);
    layer0_outputs(6862) <= not a;
    layer0_outputs(6863) <= a and not b;
    layer0_outputs(6864) <= not (a xor b);
    layer0_outputs(6865) <= a or b;
    layer0_outputs(6866) <= a and not b;
    layer0_outputs(6867) <= a;
    layer0_outputs(6868) <= a;
    layer0_outputs(6869) <= a and not b;
    layer0_outputs(6870) <= not (a and b);
    layer0_outputs(6871) <= '1';
    layer0_outputs(6872) <= b and not a;
    layer0_outputs(6873) <= not b;
    layer0_outputs(6874) <= not b or a;
    layer0_outputs(6875) <= a and not b;
    layer0_outputs(6876) <= a and not b;
    layer0_outputs(6877) <= not a or b;
    layer0_outputs(6878) <= a and b;
    layer0_outputs(6879) <= not b or a;
    layer0_outputs(6880) <= not b or a;
    layer0_outputs(6881) <= a xor b;
    layer0_outputs(6882) <= a xor b;
    layer0_outputs(6883) <= not (a or b);
    layer0_outputs(6884) <= a xor b;
    layer0_outputs(6885) <= not (a xor b);
    layer0_outputs(6886) <= not b or a;
    layer0_outputs(6887) <= not (a or b);
    layer0_outputs(6888) <= a xor b;
    layer0_outputs(6889) <= not (a or b);
    layer0_outputs(6890) <= a xor b;
    layer0_outputs(6891) <= b;
    layer0_outputs(6892) <= b;
    layer0_outputs(6893) <= a and not b;
    layer0_outputs(6894) <= a xor b;
    layer0_outputs(6895) <= not a;
    layer0_outputs(6896) <= not (a and b);
    layer0_outputs(6897) <= not b or a;
    layer0_outputs(6898) <= a xor b;
    layer0_outputs(6899) <= not b;
    layer0_outputs(6900) <= not b or a;
    layer0_outputs(6901) <= b and not a;
    layer0_outputs(6902) <= a xor b;
    layer0_outputs(6903) <= b;
    layer0_outputs(6904) <= a or b;
    layer0_outputs(6905) <= not (a and b);
    layer0_outputs(6906) <= not a;
    layer0_outputs(6907) <= a xor b;
    layer0_outputs(6908) <= a and not b;
    layer0_outputs(6909) <= not (a or b);
    layer0_outputs(6910) <= not b;
    layer0_outputs(6911) <= not (a and b);
    layer0_outputs(6912) <= not a;
    layer0_outputs(6913) <= not (a or b);
    layer0_outputs(6914) <= not a;
    layer0_outputs(6915) <= a;
    layer0_outputs(6916) <= not b or a;
    layer0_outputs(6917) <= not (a or b);
    layer0_outputs(6918) <= not a;
    layer0_outputs(6919) <= b and not a;
    layer0_outputs(6920) <= a or b;
    layer0_outputs(6921) <= not (a or b);
    layer0_outputs(6922) <= not a or b;
    layer0_outputs(6923) <= a xor b;
    layer0_outputs(6924) <= not (a or b);
    layer0_outputs(6925) <= '1';
    layer0_outputs(6926) <= not a or b;
    layer0_outputs(6927) <= not a;
    layer0_outputs(6928) <= not b;
    layer0_outputs(6929) <= a and b;
    layer0_outputs(6930) <= not (a or b);
    layer0_outputs(6931) <= not (a or b);
    layer0_outputs(6932) <= b;
    layer0_outputs(6933) <= not a;
    layer0_outputs(6934) <= '0';
    layer0_outputs(6935) <= not (a or b);
    layer0_outputs(6936) <= a;
    layer0_outputs(6937) <= '1';
    layer0_outputs(6938) <= a or b;
    layer0_outputs(6939) <= not (a xor b);
    layer0_outputs(6940) <= not b or a;
    layer0_outputs(6941) <= not (a or b);
    layer0_outputs(6942) <= not (a or b);
    layer0_outputs(6943) <= a xor b;
    layer0_outputs(6944) <= b;
    layer0_outputs(6945) <= a xor b;
    layer0_outputs(6946) <= b and not a;
    layer0_outputs(6947) <= not (a or b);
    layer0_outputs(6948) <= not b;
    layer0_outputs(6949) <= not b;
    layer0_outputs(6950) <= not (a or b);
    layer0_outputs(6951) <= not a;
    layer0_outputs(6952) <= not (a and b);
    layer0_outputs(6953) <= not (a xor b);
    layer0_outputs(6954) <= not (a or b);
    layer0_outputs(6955) <= not a;
    layer0_outputs(6956) <= '0';
    layer0_outputs(6957) <= b;
    layer0_outputs(6958) <= not b or a;
    layer0_outputs(6959) <= not b or a;
    layer0_outputs(6960) <= a xor b;
    layer0_outputs(6961) <= not b or a;
    layer0_outputs(6962) <= a and not b;
    layer0_outputs(6963) <= a xor b;
    layer0_outputs(6964) <= a xor b;
    layer0_outputs(6965) <= a;
    layer0_outputs(6966) <= not (a or b);
    layer0_outputs(6967) <= not a or b;
    layer0_outputs(6968) <= not (a and b);
    layer0_outputs(6969) <= a and not b;
    layer0_outputs(6970) <= not a or b;
    layer0_outputs(6971) <= a;
    layer0_outputs(6972) <= not a or b;
    layer0_outputs(6973) <= b;
    layer0_outputs(6974) <= not (a or b);
    layer0_outputs(6975) <= b;
    layer0_outputs(6976) <= '0';
    layer0_outputs(6977) <= not (a or b);
    layer0_outputs(6978) <= not a;
    layer0_outputs(6979) <= '1';
    layer0_outputs(6980) <= a xor b;
    layer0_outputs(6981) <= b and not a;
    layer0_outputs(6982) <= a and b;
    layer0_outputs(6983) <= not b;
    layer0_outputs(6984) <= a xor b;
    layer0_outputs(6985) <= not (a or b);
    layer0_outputs(6986) <= '1';
    layer0_outputs(6987) <= a and not b;
    layer0_outputs(6988) <= not (a or b);
    layer0_outputs(6989) <= a and not b;
    layer0_outputs(6990) <= b and not a;
    layer0_outputs(6991) <= b and not a;
    layer0_outputs(6992) <= not b or a;
    layer0_outputs(6993) <= '0';
    layer0_outputs(6994) <= not a;
    layer0_outputs(6995) <= a xor b;
    layer0_outputs(6996) <= not b or a;
    layer0_outputs(6997) <= a xor b;
    layer0_outputs(6998) <= b and not a;
    layer0_outputs(6999) <= not b;
    layer0_outputs(7000) <= a and not b;
    layer0_outputs(7001) <= a or b;
    layer0_outputs(7002) <= not a or b;
    layer0_outputs(7003) <= not a;
    layer0_outputs(7004) <= b;
    layer0_outputs(7005) <= a;
    layer0_outputs(7006) <= not (a or b);
    layer0_outputs(7007) <= not (a xor b);
    layer0_outputs(7008) <= a;
    layer0_outputs(7009) <= not (a xor b);
    layer0_outputs(7010) <= b and not a;
    layer0_outputs(7011) <= not a;
    layer0_outputs(7012) <= a and b;
    layer0_outputs(7013) <= a;
    layer0_outputs(7014) <= not a;
    layer0_outputs(7015) <= a and not b;
    layer0_outputs(7016) <= not b or a;
    layer0_outputs(7017) <= not (a xor b);
    layer0_outputs(7018) <= a xor b;
    layer0_outputs(7019) <= a xor b;
    layer0_outputs(7020) <= b and not a;
    layer0_outputs(7021) <= not a;
    layer0_outputs(7022) <= not a;
    layer0_outputs(7023) <= not a or b;
    layer0_outputs(7024) <= not (a xor b);
    layer0_outputs(7025) <= a xor b;
    layer0_outputs(7026) <= not b or a;
    layer0_outputs(7027) <= a xor b;
    layer0_outputs(7028) <= a or b;
    layer0_outputs(7029) <= not (a xor b);
    layer0_outputs(7030) <= a;
    layer0_outputs(7031) <= a or b;
    layer0_outputs(7032) <= not (a xor b);
    layer0_outputs(7033) <= not (a or b);
    layer0_outputs(7034) <= not b or a;
    layer0_outputs(7035) <= not (a or b);
    layer0_outputs(7036) <= b and not a;
    layer0_outputs(7037) <= not (a or b);
    layer0_outputs(7038) <= not b or a;
    layer0_outputs(7039) <= a or b;
    layer0_outputs(7040) <= not b or a;
    layer0_outputs(7041) <= '1';
    layer0_outputs(7042) <= not (a or b);
    layer0_outputs(7043) <= a and b;
    layer0_outputs(7044) <= not (a and b);
    layer0_outputs(7045) <= not a;
    layer0_outputs(7046) <= b;
    layer0_outputs(7047) <= not a or b;
    layer0_outputs(7048) <= not (a xor b);
    layer0_outputs(7049) <= '1';
    layer0_outputs(7050) <= not (a and b);
    layer0_outputs(7051) <= a and not b;
    layer0_outputs(7052) <= not (a and b);
    layer0_outputs(7053) <= a xor b;
    layer0_outputs(7054) <= not (a or b);
    layer0_outputs(7055) <= '1';
    layer0_outputs(7056) <= not b or a;
    layer0_outputs(7057) <= not a;
    layer0_outputs(7058) <= a xor b;
    layer0_outputs(7059) <= not b or a;
    layer0_outputs(7060) <= not (a or b);
    layer0_outputs(7061) <= not (a or b);
    layer0_outputs(7062) <= a xor b;
    layer0_outputs(7063) <= b;
    layer0_outputs(7064) <= a and not b;
    layer0_outputs(7065) <= a or b;
    layer0_outputs(7066) <= not (a xor b);
    layer0_outputs(7067) <= a and not b;
    layer0_outputs(7068) <= '0';
    layer0_outputs(7069) <= a and not b;
    layer0_outputs(7070) <= a or b;
    layer0_outputs(7071) <= a;
    layer0_outputs(7072) <= not a or b;
    layer0_outputs(7073) <= not (a or b);
    layer0_outputs(7074) <= a;
    layer0_outputs(7075) <= a;
    layer0_outputs(7076) <= a or b;
    layer0_outputs(7077) <= '1';
    layer0_outputs(7078) <= a xor b;
    layer0_outputs(7079) <= a;
    layer0_outputs(7080) <= not (a xor b);
    layer0_outputs(7081) <= a;
    layer0_outputs(7082) <= a or b;
    layer0_outputs(7083) <= not (a xor b);
    layer0_outputs(7084) <= not (a or b);
    layer0_outputs(7085) <= b and not a;
    layer0_outputs(7086) <= not (a or b);
    layer0_outputs(7087) <= a or b;
    layer0_outputs(7088) <= not a or b;
    layer0_outputs(7089) <= b and not a;
    layer0_outputs(7090) <= '0';
    layer0_outputs(7091) <= a or b;
    layer0_outputs(7092) <= a;
    layer0_outputs(7093) <= not b;
    layer0_outputs(7094) <= a;
    layer0_outputs(7095) <= not (a xor b);
    layer0_outputs(7096) <= a;
    layer0_outputs(7097) <= not (a xor b);
    layer0_outputs(7098) <= not (a xor b);
    layer0_outputs(7099) <= not b;
    layer0_outputs(7100) <= '0';
    layer0_outputs(7101) <= a and b;
    layer0_outputs(7102) <= b and not a;
    layer0_outputs(7103) <= a;
    layer0_outputs(7104) <= a and b;
    layer0_outputs(7105) <= not (a or b);
    layer0_outputs(7106) <= a and not b;
    layer0_outputs(7107) <= a or b;
    layer0_outputs(7108) <= '1';
    layer0_outputs(7109) <= not a;
    layer0_outputs(7110) <= a;
    layer0_outputs(7111) <= not (a and b);
    layer0_outputs(7112) <= not (a or b);
    layer0_outputs(7113) <= b;
    layer0_outputs(7114) <= not (a or b);
    layer0_outputs(7115) <= b and not a;
    layer0_outputs(7116) <= not (a xor b);
    layer0_outputs(7117) <= not (a xor b);
    layer0_outputs(7118) <= b;
    layer0_outputs(7119) <= a;
    layer0_outputs(7120) <= not (a xor b);
    layer0_outputs(7121) <= a xor b;
    layer0_outputs(7122) <= a or b;
    layer0_outputs(7123) <= not a or b;
    layer0_outputs(7124) <= a or b;
    layer0_outputs(7125) <= not b or a;
    layer0_outputs(7126) <= b and not a;
    layer0_outputs(7127) <= not (a or b);
    layer0_outputs(7128) <= not (a xor b);
    layer0_outputs(7129) <= not (a xor b);
    layer0_outputs(7130) <= not (a or b);
    layer0_outputs(7131) <= a and not b;
    layer0_outputs(7132) <= not (a or b);
    layer0_outputs(7133) <= b and not a;
    layer0_outputs(7134) <= a or b;
    layer0_outputs(7135) <= b and not a;
    layer0_outputs(7136) <= a or b;
    layer0_outputs(7137) <= not a or b;
    layer0_outputs(7138) <= a;
    layer0_outputs(7139) <= not b or a;
    layer0_outputs(7140) <= a xor b;
    layer0_outputs(7141) <= '0';
    layer0_outputs(7142) <= a and not b;
    layer0_outputs(7143) <= not (a xor b);
    layer0_outputs(7144) <= not b or a;
    layer0_outputs(7145) <= not (a or b);
    layer0_outputs(7146) <= a;
    layer0_outputs(7147) <= not (a xor b);
    layer0_outputs(7148) <= a and not b;
    layer0_outputs(7149) <= not a;
    layer0_outputs(7150) <= a and not b;
    layer0_outputs(7151) <= a;
    layer0_outputs(7152) <= a or b;
    layer0_outputs(7153) <= not b;
    layer0_outputs(7154) <= not (a or b);
    layer0_outputs(7155) <= not (a xor b);
    layer0_outputs(7156) <= a xor b;
    layer0_outputs(7157) <= a xor b;
    layer0_outputs(7158) <= not (a or b);
    layer0_outputs(7159) <= a;
    layer0_outputs(7160) <= not b;
    layer0_outputs(7161) <= '0';
    layer0_outputs(7162) <= not (a xor b);
    layer0_outputs(7163) <= a;
    layer0_outputs(7164) <= not b;
    layer0_outputs(7165) <= b and not a;
    layer0_outputs(7166) <= not (a and b);
    layer0_outputs(7167) <= b;
    layer0_outputs(7168) <= not (a and b);
    layer0_outputs(7169) <= a or b;
    layer0_outputs(7170) <= '0';
    layer0_outputs(7171) <= b and not a;
    layer0_outputs(7172) <= not (a or b);
    layer0_outputs(7173) <= not (a xor b);
    layer0_outputs(7174) <= not (a or b);
    layer0_outputs(7175) <= a or b;
    layer0_outputs(7176) <= not a or b;
    layer0_outputs(7177) <= not a;
    layer0_outputs(7178) <= a and not b;
    layer0_outputs(7179) <= not (a or b);
    layer0_outputs(7180) <= not (a xor b);
    layer0_outputs(7181) <= not (a or b);
    layer0_outputs(7182) <= a and not b;
    layer0_outputs(7183) <= b;
    layer0_outputs(7184) <= not b or a;
    layer0_outputs(7185) <= '0';
    layer0_outputs(7186) <= not (a or b);
    layer0_outputs(7187) <= not a;
    layer0_outputs(7188) <= b;
    layer0_outputs(7189) <= a and not b;
    layer0_outputs(7190) <= b and not a;
    layer0_outputs(7191) <= a;
    layer0_outputs(7192) <= '1';
    layer0_outputs(7193) <= '0';
    layer0_outputs(7194) <= not a or b;
    layer0_outputs(7195) <= a and b;
    layer0_outputs(7196) <= not (a xor b);
    layer0_outputs(7197) <= not (a xor b);
    layer0_outputs(7198) <= '0';
    layer0_outputs(7199) <= not (a or b);
    layer0_outputs(7200) <= a;
    layer0_outputs(7201) <= not (a xor b);
    layer0_outputs(7202) <= not b or a;
    layer0_outputs(7203) <= not (a xor b);
    layer0_outputs(7204) <= not (a xor b);
    layer0_outputs(7205) <= not a or b;
    layer0_outputs(7206) <= a or b;
    layer0_outputs(7207) <= b and not a;
    layer0_outputs(7208) <= not a;
    layer0_outputs(7209) <= not (a and b);
    layer0_outputs(7210) <= b;
    layer0_outputs(7211) <= not (a or b);
    layer0_outputs(7212) <= not (a xor b);
    layer0_outputs(7213) <= not (a and b);
    layer0_outputs(7214) <= not (a or b);
    layer0_outputs(7215) <= '0';
    layer0_outputs(7216) <= a xor b;
    layer0_outputs(7217) <= a;
    layer0_outputs(7218) <= b;
    layer0_outputs(7219) <= not (a or b);
    layer0_outputs(7220) <= b and not a;
    layer0_outputs(7221) <= a;
    layer0_outputs(7222) <= b and not a;
    layer0_outputs(7223) <= not a or b;
    layer0_outputs(7224) <= b and not a;
    layer0_outputs(7225) <= not (a or b);
    layer0_outputs(7226) <= b and not a;
    layer0_outputs(7227) <= not (a or b);
    layer0_outputs(7228) <= not b;
    layer0_outputs(7229) <= not a;
    layer0_outputs(7230) <= a xor b;
    layer0_outputs(7231) <= a and b;
    layer0_outputs(7232) <= a or b;
    layer0_outputs(7233) <= b;
    layer0_outputs(7234) <= a;
    layer0_outputs(7235) <= a xor b;
    layer0_outputs(7236) <= not (a xor b);
    layer0_outputs(7237) <= b;
    layer0_outputs(7238) <= b;
    layer0_outputs(7239) <= b and not a;
    layer0_outputs(7240) <= not (a or b);
    layer0_outputs(7241) <= a xor b;
    layer0_outputs(7242) <= not a or b;
    layer0_outputs(7243) <= a xor b;
    layer0_outputs(7244) <= not (a xor b);
    layer0_outputs(7245) <= not a;
    layer0_outputs(7246) <= not (a or b);
    layer0_outputs(7247) <= b;
    layer0_outputs(7248) <= a or b;
    layer0_outputs(7249) <= a or b;
    layer0_outputs(7250) <= b;
    layer0_outputs(7251) <= not a;
    layer0_outputs(7252) <= not a or b;
    layer0_outputs(7253) <= b;
    layer0_outputs(7254) <= a;
    layer0_outputs(7255) <= a and not b;
    layer0_outputs(7256) <= not (a xor b);
    layer0_outputs(7257) <= b and not a;
    layer0_outputs(7258) <= not b;
    layer0_outputs(7259) <= not (a xor b);
    layer0_outputs(7260) <= a or b;
    layer0_outputs(7261) <= a or b;
    layer0_outputs(7262) <= a;
    layer0_outputs(7263) <= not a;
    layer0_outputs(7264) <= a xor b;
    layer0_outputs(7265) <= not (a xor b);
    layer0_outputs(7266) <= not a or b;
    layer0_outputs(7267) <= a;
    layer0_outputs(7268) <= a or b;
    layer0_outputs(7269) <= a and not b;
    layer0_outputs(7270) <= a or b;
    layer0_outputs(7271) <= a and b;
    layer0_outputs(7272) <= a or b;
    layer0_outputs(7273) <= not (a or b);
    layer0_outputs(7274) <= not b or a;
    layer0_outputs(7275) <= '0';
    layer0_outputs(7276) <= a xor b;
    layer0_outputs(7277) <= '1';
    layer0_outputs(7278) <= not (a xor b);
    layer0_outputs(7279) <= a;
    layer0_outputs(7280) <= a and b;
    layer0_outputs(7281) <= a or b;
    layer0_outputs(7282) <= not (a or b);
    layer0_outputs(7283) <= not (a and b);
    layer0_outputs(7284) <= a;
    layer0_outputs(7285) <= not (a or b);
    layer0_outputs(7286) <= not b or a;
    layer0_outputs(7287) <= a;
    layer0_outputs(7288) <= a or b;
    layer0_outputs(7289) <= not (a xor b);
    layer0_outputs(7290) <= not a;
    layer0_outputs(7291) <= not a or b;
    layer0_outputs(7292) <= a or b;
    layer0_outputs(7293) <= a;
    layer0_outputs(7294) <= a or b;
    layer0_outputs(7295) <= not a or b;
    layer0_outputs(7296) <= b and not a;
    layer0_outputs(7297) <= not (a and b);
    layer0_outputs(7298) <= not (a xor b);
    layer0_outputs(7299) <= b;
    layer0_outputs(7300) <= not (a xor b);
    layer0_outputs(7301) <= not b;
    layer0_outputs(7302) <= not (a and b);
    layer0_outputs(7303) <= '0';
    layer0_outputs(7304) <= a xor b;
    layer0_outputs(7305) <= a or b;
    layer0_outputs(7306) <= b;
    layer0_outputs(7307) <= not a;
    layer0_outputs(7308) <= a and b;
    layer0_outputs(7309) <= a and not b;
    layer0_outputs(7310) <= b and not a;
    layer0_outputs(7311) <= '1';
    layer0_outputs(7312) <= a or b;
    layer0_outputs(7313) <= not (a and b);
    layer0_outputs(7314) <= a xor b;
    layer0_outputs(7315) <= not a;
    layer0_outputs(7316) <= b;
    layer0_outputs(7317) <= not b or a;
    layer0_outputs(7318) <= b and not a;
    layer0_outputs(7319) <= not a or b;
    layer0_outputs(7320) <= a;
    layer0_outputs(7321) <= a and not b;
    layer0_outputs(7322) <= a;
    layer0_outputs(7323) <= not a or b;
    layer0_outputs(7324) <= a xor b;
    layer0_outputs(7325) <= a or b;
    layer0_outputs(7326) <= a xor b;
    layer0_outputs(7327) <= a and not b;
    layer0_outputs(7328) <= not (a and b);
    layer0_outputs(7329) <= a or b;
    layer0_outputs(7330) <= not a;
    layer0_outputs(7331) <= a xor b;
    layer0_outputs(7332) <= a or b;
    layer0_outputs(7333) <= a or b;
    layer0_outputs(7334) <= a and b;
    layer0_outputs(7335) <= not b or a;
    layer0_outputs(7336) <= not a or b;
    layer0_outputs(7337) <= a and b;
    layer0_outputs(7338) <= b;
    layer0_outputs(7339) <= b;
    layer0_outputs(7340) <= not a or b;
    layer0_outputs(7341) <= not (a xor b);
    layer0_outputs(7342) <= not (a or b);
    layer0_outputs(7343) <= not (a and b);
    layer0_outputs(7344) <= a and not b;
    layer0_outputs(7345) <= not a;
    layer0_outputs(7346) <= not a or b;
    layer0_outputs(7347) <= b;
    layer0_outputs(7348) <= not b;
    layer0_outputs(7349) <= not b;
    layer0_outputs(7350) <= not b;
    layer0_outputs(7351) <= not a or b;
    layer0_outputs(7352) <= not a or b;
    layer0_outputs(7353) <= a and b;
    layer0_outputs(7354) <= not (a xor b);
    layer0_outputs(7355) <= not b;
    layer0_outputs(7356) <= not (a xor b);
    layer0_outputs(7357) <= a;
    layer0_outputs(7358) <= not (a xor b);
    layer0_outputs(7359) <= not (a or b);
    layer0_outputs(7360) <= a and not b;
    layer0_outputs(7361) <= a xor b;
    layer0_outputs(7362) <= a or b;
    layer0_outputs(7363) <= b and not a;
    layer0_outputs(7364) <= a xor b;
    layer0_outputs(7365) <= b and not a;
    layer0_outputs(7366) <= a or b;
    layer0_outputs(7367) <= b;
    layer0_outputs(7368) <= a;
    layer0_outputs(7369) <= not a;
    layer0_outputs(7370) <= not b;
    layer0_outputs(7371) <= not (a or b);
    layer0_outputs(7372) <= not a;
    layer0_outputs(7373) <= not (a xor b);
    layer0_outputs(7374) <= a and b;
    layer0_outputs(7375) <= not a;
    layer0_outputs(7376) <= not a or b;
    layer0_outputs(7377) <= '1';
    layer0_outputs(7378) <= not b;
    layer0_outputs(7379) <= '1';
    layer0_outputs(7380) <= not b;
    layer0_outputs(7381) <= a and not b;
    layer0_outputs(7382) <= not (a xor b);
    layer0_outputs(7383) <= a xor b;
    layer0_outputs(7384) <= '0';
    layer0_outputs(7385) <= a and not b;
    layer0_outputs(7386) <= not a;
    layer0_outputs(7387) <= b and not a;
    layer0_outputs(7388) <= '1';
    layer0_outputs(7389) <= not (a xor b);
    layer0_outputs(7390) <= '1';
    layer0_outputs(7391) <= a xor b;
    layer0_outputs(7392) <= not b or a;
    layer0_outputs(7393) <= not b;
    layer0_outputs(7394) <= not (a or b);
    layer0_outputs(7395) <= a or b;
    layer0_outputs(7396) <= not a or b;
    layer0_outputs(7397) <= b;
    layer0_outputs(7398) <= not b;
    layer0_outputs(7399) <= b and not a;
    layer0_outputs(7400) <= not (a or b);
    layer0_outputs(7401) <= not (a xor b);
    layer0_outputs(7402) <= not (a and b);
    layer0_outputs(7403) <= not (a or b);
    layer0_outputs(7404) <= not a or b;
    layer0_outputs(7405) <= not (a and b);
    layer0_outputs(7406) <= not (a xor b);
    layer0_outputs(7407) <= a xor b;
    layer0_outputs(7408) <= not a;
    layer0_outputs(7409) <= '0';
    layer0_outputs(7410) <= not b or a;
    layer0_outputs(7411) <= a and not b;
    layer0_outputs(7412) <= a or b;
    layer0_outputs(7413) <= a;
    layer0_outputs(7414) <= not a;
    layer0_outputs(7415) <= a or b;
    layer0_outputs(7416) <= b;
    layer0_outputs(7417) <= a or b;
    layer0_outputs(7418) <= a xor b;
    layer0_outputs(7419) <= not a;
    layer0_outputs(7420) <= not a or b;
    layer0_outputs(7421) <= not a or b;
    layer0_outputs(7422) <= a;
    layer0_outputs(7423) <= a or b;
    layer0_outputs(7424) <= a;
    layer0_outputs(7425) <= a and not b;
    layer0_outputs(7426) <= b and not a;
    layer0_outputs(7427) <= b;
    layer0_outputs(7428) <= not (a xor b);
    layer0_outputs(7429) <= not (a and b);
    layer0_outputs(7430) <= a or b;
    layer0_outputs(7431) <= not b or a;
    layer0_outputs(7432) <= a;
    layer0_outputs(7433) <= not (a or b);
    layer0_outputs(7434) <= not b;
    layer0_outputs(7435) <= not (a and b);
    layer0_outputs(7436) <= b;
    layer0_outputs(7437) <= b and not a;
    layer0_outputs(7438) <= not b;
    layer0_outputs(7439) <= a and not b;
    layer0_outputs(7440) <= a;
    layer0_outputs(7441) <= a and not b;
    layer0_outputs(7442) <= a xor b;
    layer0_outputs(7443) <= not b or a;
    layer0_outputs(7444) <= b;
    layer0_outputs(7445) <= not (a or b);
    layer0_outputs(7446) <= a and not b;
    layer0_outputs(7447) <= not b;
    layer0_outputs(7448) <= a;
    layer0_outputs(7449) <= not b;
    layer0_outputs(7450) <= a or b;
    layer0_outputs(7451) <= b;
    layer0_outputs(7452) <= not a or b;
    layer0_outputs(7453) <= a or b;
    layer0_outputs(7454) <= a;
    layer0_outputs(7455) <= a or b;
    layer0_outputs(7456) <= not b;
    layer0_outputs(7457) <= a or b;
    layer0_outputs(7458) <= not a;
    layer0_outputs(7459) <= b;
    layer0_outputs(7460) <= b;
    layer0_outputs(7461) <= a;
    layer0_outputs(7462) <= not a or b;
    layer0_outputs(7463) <= a xor b;
    layer0_outputs(7464) <= not (a or b);
    layer0_outputs(7465) <= a xor b;
    layer0_outputs(7466) <= not a or b;
    layer0_outputs(7467) <= not (a or b);
    layer0_outputs(7468) <= a or b;
    layer0_outputs(7469) <= not b or a;
    layer0_outputs(7470) <= a and b;
    layer0_outputs(7471) <= not a or b;
    layer0_outputs(7472) <= not b;
    layer0_outputs(7473) <= b and not a;
    layer0_outputs(7474) <= a xor b;
    layer0_outputs(7475) <= a xor b;
    layer0_outputs(7476) <= a xor b;
    layer0_outputs(7477) <= b;
    layer0_outputs(7478) <= not (a and b);
    layer0_outputs(7479) <= a;
    layer0_outputs(7480) <= not (a and b);
    layer0_outputs(7481) <= a and b;
    layer0_outputs(7482) <= a or b;
    layer0_outputs(7483) <= a or b;
    layer0_outputs(7484) <= b and not a;
    layer0_outputs(7485) <= not (a xor b);
    layer0_outputs(7486) <= not (a xor b);
    layer0_outputs(7487) <= b and not a;
    layer0_outputs(7488) <= a or b;
    layer0_outputs(7489) <= a or b;
    layer0_outputs(7490) <= not (a or b);
    layer0_outputs(7491) <= a xor b;
    layer0_outputs(7492) <= not (a or b);
    layer0_outputs(7493) <= b and not a;
    layer0_outputs(7494) <= b and not a;
    layer0_outputs(7495) <= not (a or b);
    layer0_outputs(7496) <= not b;
    layer0_outputs(7497) <= b and not a;
    layer0_outputs(7498) <= b and not a;
    layer0_outputs(7499) <= not a;
    layer0_outputs(7500) <= not a or b;
    layer0_outputs(7501) <= b;
    layer0_outputs(7502) <= a;
    layer0_outputs(7503) <= not (a or b);
    layer0_outputs(7504) <= not (a or b);
    layer0_outputs(7505) <= not (a and b);
    layer0_outputs(7506) <= a or b;
    layer0_outputs(7507) <= not b;
    layer0_outputs(7508) <= a xor b;
    layer0_outputs(7509) <= not (a or b);
    layer0_outputs(7510) <= a or b;
    layer0_outputs(7511) <= not b;
    layer0_outputs(7512) <= a or b;
    layer0_outputs(7513) <= a or b;
    layer0_outputs(7514) <= not (a xor b);
    layer0_outputs(7515) <= not (a or b);
    layer0_outputs(7516) <= b and not a;
    layer0_outputs(7517) <= not (a or b);
    layer0_outputs(7518) <= a and not b;
    layer0_outputs(7519) <= not (a and b);
    layer0_outputs(7520) <= a and not b;
    layer0_outputs(7521) <= '1';
    layer0_outputs(7522) <= a or b;
    layer0_outputs(7523) <= not b or a;
    layer0_outputs(7524) <= a xor b;
    layer0_outputs(7525) <= a or b;
    layer0_outputs(7526) <= b;
    layer0_outputs(7527) <= not (a or b);
    layer0_outputs(7528) <= not a or b;
    layer0_outputs(7529) <= not (a or b);
    layer0_outputs(7530) <= a xor b;
    layer0_outputs(7531) <= not a or b;
    layer0_outputs(7532) <= a or b;
    layer0_outputs(7533) <= '0';
    layer0_outputs(7534) <= not a or b;
    layer0_outputs(7535) <= a or b;
    layer0_outputs(7536) <= not a;
    layer0_outputs(7537) <= b;
    layer0_outputs(7538) <= not b;
    layer0_outputs(7539) <= not b;
    layer0_outputs(7540) <= not (a and b);
    layer0_outputs(7541) <= not (a xor b);
    layer0_outputs(7542) <= not a or b;
    layer0_outputs(7543) <= b and not a;
    layer0_outputs(7544) <= a and not b;
    layer0_outputs(7545) <= not a;
    layer0_outputs(7546) <= not (a xor b);
    layer0_outputs(7547) <= b;
    layer0_outputs(7548) <= not (a xor b);
    layer0_outputs(7549) <= b and not a;
    layer0_outputs(7550) <= a;
    layer0_outputs(7551) <= '0';
    layer0_outputs(7552) <= not b or a;
    layer0_outputs(7553) <= not b or a;
    layer0_outputs(7554) <= not a;
    layer0_outputs(7555) <= a;
    layer0_outputs(7556) <= not (a xor b);
    layer0_outputs(7557) <= not a;
    layer0_outputs(7558) <= '0';
    layer0_outputs(7559) <= a xor b;
    layer0_outputs(7560) <= '1';
    layer0_outputs(7561) <= not (a or b);
    layer0_outputs(7562) <= a or b;
    layer0_outputs(7563) <= '0';
    layer0_outputs(7564) <= a and b;
    layer0_outputs(7565) <= a or b;
    layer0_outputs(7566) <= not b or a;
    layer0_outputs(7567) <= a xor b;
    layer0_outputs(7568) <= a xor b;
    layer0_outputs(7569) <= not b;
    layer0_outputs(7570) <= a and not b;
    layer0_outputs(7571) <= not (a or b);
    layer0_outputs(7572) <= a;
    layer0_outputs(7573) <= not (a or b);
    layer0_outputs(7574) <= a xor b;
    layer0_outputs(7575) <= '0';
    layer0_outputs(7576) <= not a;
    layer0_outputs(7577) <= a or b;
    layer0_outputs(7578) <= a and not b;
    layer0_outputs(7579) <= a;
    layer0_outputs(7580) <= a or b;
    layer0_outputs(7581) <= not (a and b);
    layer0_outputs(7582) <= b;
    layer0_outputs(7583) <= not (a xor b);
    layer0_outputs(7584) <= b;
    layer0_outputs(7585) <= b;
    layer0_outputs(7586) <= b;
    layer0_outputs(7587) <= b;
    layer0_outputs(7588) <= a or b;
    layer0_outputs(7589) <= not a or b;
    layer0_outputs(7590) <= not (a or b);
    layer0_outputs(7591) <= not (a xor b);
    layer0_outputs(7592) <= a xor b;
    layer0_outputs(7593) <= b;
    layer0_outputs(7594) <= not (a or b);
    layer0_outputs(7595) <= a or b;
    layer0_outputs(7596) <= a xor b;
    layer0_outputs(7597) <= not (a or b);
    layer0_outputs(7598) <= not a;
    layer0_outputs(7599) <= not (a or b);
    layer0_outputs(7600) <= '0';
    layer0_outputs(7601) <= a or b;
    layer0_outputs(7602) <= a and not b;
    layer0_outputs(7603) <= '1';
    layer0_outputs(7604) <= not (a or b);
    layer0_outputs(7605) <= not (a and b);
    layer0_outputs(7606) <= not b or a;
    layer0_outputs(7607) <= not (a or b);
    layer0_outputs(7608) <= a and b;
    layer0_outputs(7609) <= b;
    layer0_outputs(7610) <= not (a xor b);
    layer0_outputs(7611) <= b and not a;
    layer0_outputs(7612) <= not a;
    layer0_outputs(7613) <= not a or b;
    layer0_outputs(7614) <= b;
    layer0_outputs(7615) <= not a;
    layer0_outputs(7616) <= not (a or b);
    layer0_outputs(7617) <= a or b;
    layer0_outputs(7618) <= a and not b;
    layer0_outputs(7619) <= not a or b;
    layer0_outputs(7620) <= not a;
    layer0_outputs(7621) <= not a;
    layer0_outputs(7622) <= b and not a;
    layer0_outputs(7623) <= not (a xor b);
    layer0_outputs(7624) <= a;
    layer0_outputs(7625) <= not a;
    layer0_outputs(7626) <= a xor b;
    layer0_outputs(7627) <= not b or a;
    layer0_outputs(7628) <= not b or a;
    layer0_outputs(7629) <= '0';
    layer0_outputs(7630) <= b;
    layer0_outputs(7631) <= a or b;
    layer0_outputs(7632) <= not b;
    layer0_outputs(7633) <= a xor b;
    layer0_outputs(7634) <= not b;
    layer0_outputs(7635) <= not a or b;
    layer0_outputs(7636) <= not (a or b);
    layer0_outputs(7637) <= b and not a;
    layer0_outputs(7638) <= a or b;
    layer0_outputs(7639) <= a and not b;
    layer0_outputs(7640) <= not (a or b);
    layer0_outputs(7641) <= not (a xor b);
    layer0_outputs(7642) <= not (a or b);
    layer0_outputs(7643) <= b;
    layer0_outputs(7644) <= a and not b;
    layer0_outputs(7645) <= a or b;
    layer0_outputs(7646) <= a or b;
    layer0_outputs(7647) <= a;
    layer0_outputs(7648) <= not a or b;
    layer0_outputs(7649) <= not a or b;
    layer0_outputs(7650) <= b and not a;
    layer0_outputs(7651) <= a;
    layer0_outputs(7652) <= a xor b;
    layer0_outputs(7653) <= a xor b;
    layer0_outputs(7654) <= not (a or b);
    layer0_outputs(7655) <= a or b;
    layer0_outputs(7656) <= not b or a;
    layer0_outputs(7657) <= a xor b;
    layer0_outputs(7658) <= '0';
    layer0_outputs(7659) <= a;
    layer0_outputs(7660) <= a or b;
    layer0_outputs(7661) <= a or b;
    layer0_outputs(7662) <= not (a or b);
    layer0_outputs(7663) <= not b;
    layer0_outputs(7664) <= not a;
    layer0_outputs(7665) <= not b or a;
    layer0_outputs(7666) <= not (a and b);
    layer0_outputs(7667) <= not a;
    layer0_outputs(7668) <= not (a or b);
    layer0_outputs(7669) <= not b;
    layer0_outputs(7670) <= not b;
    layer0_outputs(7671) <= a and not b;
    layer0_outputs(7672) <= a or b;
    layer0_outputs(7673) <= a xor b;
    layer0_outputs(7674) <= b and not a;
    layer0_outputs(7675) <= not a;
    layer0_outputs(7676) <= a xor b;
    layer0_outputs(7677) <= a or b;
    layer0_outputs(7678) <= b and not a;
    layer0_outputs(7679) <= a and b;
    layer0_outputs(7680) <= not a;
    layer0_outputs(7681) <= b;
    layer0_outputs(7682) <= not b;
    layer0_outputs(7683) <= b;
    layer0_outputs(7684) <= not (a xor b);
    layer0_outputs(7685) <= not b;
    layer0_outputs(7686) <= not b;
    layer0_outputs(7687) <= not a or b;
    layer0_outputs(7688) <= not (a or b);
    layer0_outputs(7689) <= a or b;
    layer0_outputs(7690) <= a and not b;
    layer0_outputs(7691) <= not (a or b);
    layer0_outputs(7692) <= '1';
    layer0_outputs(7693) <= not a;
    layer0_outputs(7694) <= not (a xor b);
    layer0_outputs(7695) <= a xor b;
    layer0_outputs(7696) <= not (a or b);
    layer0_outputs(7697) <= not (a or b);
    layer0_outputs(7698) <= a or b;
    layer0_outputs(7699) <= not (a xor b);
    layer0_outputs(7700) <= b and not a;
    layer0_outputs(7701) <= b;
    layer0_outputs(7702) <= '1';
    layer0_outputs(7703) <= not b or a;
    layer0_outputs(7704) <= not (a or b);
    layer0_outputs(7705) <= not a;
    layer0_outputs(7706) <= a and not b;
    layer0_outputs(7707) <= not (a xor b);
    layer0_outputs(7708) <= not (a or b);
    layer0_outputs(7709) <= a xor b;
    layer0_outputs(7710) <= a xor b;
    layer0_outputs(7711) <= not b;
    layer0_outputs(7712) <= not a or b;
    layer0_outputs(7713) <= '0';
    layer0_outputs(7714) <= b and not a;
    layer0_outputs(7715) <= a xor b;
    layer0_outputs(7716) <= not (a or b);
    layer0_outputs(7717) <= not (a xor b);
    layer0_outputs(7718) <= a xor b;
    layer0_outputs(7719) <= not b or a;
    layer0_outputs(7720) <= a or b;
    layer0_outputs(7721) <= a and not b;
    layer0_outputs(7722) <= a or b;
    layer0_outputs(7723) <= a and not b;
    layer0_outputs(7724) <= a or b;
    layer0_outputs(7725) <= not a;
    layer0_outputs(7726) <= a;
    layer0_outputs(7727) <= a;
    layer0_outputs(7728) <= not (a xor b);
    layer0_outputs(7729) <= not (a and b);
    layer0_outputs(7730) <= not (a or b);
    layer0_outputs(7731) <= not (a xor b);
    layer0_outputs(7732) <= a xor b;
    layer0_outputs(7733) <= a or b;
    layer0_outputs(7734) <= not b or a;
    layer0_outputs(7735) <= not (a xor b);
    layer0_outputs(7736) <= a;
    layer0_outputs(7737) <= not a or b;
    layer0_outputs(7738) <= not b or a;
    layer0_outputs(7739) <= a xor b;
    layer0_outputs(7740) <= not (a xor b);
    layer0_outputs(7741) <= a or b;
    layer0_outputs(7742) <= '1';
    layer0_outputs(7743) <= not (a xor b);
    layer0_outputs(7744) <= not b or a;
    layer0_outputs(7745) <= b and not a;
    layer0_outputs(7746) <= not a or b;
    layer0_outputs(7747) <= not b;
    layer0_outputs(7748) <= a xor b;
    layer0_outputs(7749) <= not b or a;
    layer0_outputs(7750) <= a or b;
    layer0_outputs(7751) <= '1';
    layer0_outputs(7752) <= a;
    layer0_outputs(7753) <= a xor b;
    layer0_outputs(7754) <= a xor b;
    layer0_outputs(7755) <= not (a and b);
    layer0_outputs(7756) <= a and b;
    layer0_outputs(7757) <= not (a or b);
    layer0_outputs(7758) <= not (a or b);
    layer0_outputs(7759) <= b;
    layer0_outputs(7760) <= not (a xor b);
    layer0_outputs(7761) <= not b;
    layer0_outputs(7762) <= not (a or b);
    layer0_outputs(7763) <= b and not a;
    layer0_outputs(7764) <= b;
    layer0_outputs(7765) <= '0';
    layer0_outputs(7766) <= b and not a;
    layer0_outputs(7767) <= not (a xor b);
    layer0_outputs(7768) <= not b;
    layer0_outputs(7769) <= b;
    layer0_outputs(7770) <= a or b;
    layer0_outputs(7771) <= not a;
    layer0_outputs(7772) <= '1';
    layer0_outputs(7773) <= a or b;
    layer0_outputs(7774) <= not b;
    layer0_outputs(7775) <= '0';
    layer0_outputs(7776) <= not (a or b);
    layer0_outputs(7777) <= a and not b;
    layer0_outputs(7778) <= not a or b;
    layer0_outputs(7779) <= a or b;
    layer0_outputs(7780) <= not a;
    layer0_outputs(7781) <= '0';
    layer0_outputs(7782) <= not b or a;
    layer0_outputs(7783) <= not (a xor b);
    layer0_outputs(7784) <= a or b;
    layer0_outputs(7785) <= a or b;
    layer0_outputs(7786) <= b and not a;
    layer0_outputs(7787) <= a or b;
    layer0_outputs(7788) <= not (a xor b);
    layer0_outputs(7789) <= not (a xor b);
    layer0_outputs(7790) <= not (a xor b);
    layer0_outputs(7791) <= a;
    layer0_outputs(7792) <= a;
    layer0_outputs(7793) <= not b or a;
    layer0_outputs(7794) <= not b or a;
    layer0_outputs(7795) <= not b or a;
    layer0_outputs(7796) <= b and not a;
    layer0_outputs(7797) <= b and not a;
    layer0_outputs(7798) <= not (a or b);
    layer0_outputs(7799) <= a;
    layer0_outputs(7800) <= not a or b;
    layer0_outputs(7801) <= not (a xor b);
    layer0_outputs(7802) <= not (a xor b);
    layer0_outputs(7803) <= not (a xor b);
    layer0_outputs(7804) <= '1';
    layer0_outputs(7805) <= a and b;
    layer0_outputs(7806) <= a or b;
    layer0_outputs(7807) <= a or b;
    layer0_outputs(7808) <= not (a xor b);
    layer0_outputs(7809) <= a;
    layer0_outputs(7810) <= a or b;
    layer0_outputs(7811) <= a xor b;
    layer0_outputs(7812) <= b and not a;
    layer0_outputs(7813) <= not b or a;
    layer0_outputs(7814) <= not (a xor b);
    layer0_outputs(7815) <= not (a and b);
    layer0_outputs(7816) <= not a;
    layer0_outputs(7817) <= a or b;
    layer0_outputs(7818) <= a or b;
    layer0_outputs(7819) <= a;
    layer0_outputs(7820) <= a or b;
    layer0_outputs(7821) <= '1';
    layer0_outputs(7822) <= not (a or b);
    layer0_outputs(7823) <= b and not a;
    layer0_outputs(7824) <= b and not a;
    layer0_outputs(7825) <= a or b;
    layer0_outputs(7826) <= a or b;
    layer0_outputs(7827) <= not b;
    layer0_outputs(7828) <= a;
    layer0_outputs(7829) <= not b or a;
    layer0_outputs(7830) <= not a;
    layer0_outputs(7831) <= not (a or b);
    layer0_outputs(7832) <= a or b;
    layer0_outputs(7833) <= b and not a;
    layer0_outputs(7834) <= b;
    layer0_outputs(7835) <= not a or b;
    layer0_outputs(7836) <= a xor b;
    layer0_outputs(7837) <= not b or a;
    layer0_outputs(7838) <= not b;
    layer0_outputs(7839) <= not (a or b);
    layer0_outputs(7840) <= b;
    layer0_outputs(7841) <= not b;
    layer0_outputs(7842) <= a or b;
    layer0_outputs(7843) <= not b;
    layer0_outputs(7844) <= not (a xor b);
    layer0_outputs(7845) <= a xor b;
    layer0_outputs(7846) <= not b;
    layer0_outputs(7847) <= not b or a;
    layer0_outputs(7848) <= not a or b;
    layer0_outputs(7849) <= not (a or b);
    layer0_outputs(7850) <= a or b;
    layer0_outputs(7851) <= a or b;
    layer0_outputs(7852) <= b and not a;
    layer0_outputs(7853) <= a or b;
    layer0_outputs(7854) <= not b or a;
    layer0_outputs(7855) <= a;
    layer0_outputs(7856) <= not b or a;
    layer0_outputs(7857) <= not (a or b);
    layer0_outputs(7858) <= a and b;
    layer0_outputs(7859) <= a;
    layer0_outputs(7860) <= not (a and b);
    layer0_outputs(7861) <= a and b;
    layer0_outputs(7862) <= not (a xor b);
    layer0_outputs(7863) <= not a;
    layer0_outputs(7864) <= not (a xor b);
    layer0_outputs(7865) <= a or b;
    layer0_outputs(7866) <= a and not b;
    layer0_outputs(7867) <= not a;
    layer0_outputs(7868) <= b and not a;
    layer0_outputs(7869) <= not (a xor b);
    layer0_outputs(7870) <= a or b;
    layer0_outputs(7871) <= b;
    layer0_outputs(7872) <= not (a xor b);
    layer0_outputs(7873) <= not (a xor b);
    layer0_outputs(7874) <= a xor b;
    layer0_outputs(7875) <= a and not b;
    layer0_outputs(7876) <= a or b;
    layer0_outputs(7877) <= a;
    layer0_outputs(7878) <= a and b;
    layer0_outputs(7879) <= b and not a;
    layer0_outputs(7880) <= not (a or b);
    layer0_outputs(7881) <= not b;
    layer0_outputs(7882) <= a;
    layer0_outputs(7883) <= a;
    layer0_outputs(7884) <= b;
    layer0_outputs(7885) <= a xor b;
    layer0_outputs(7886) <= not a;
    layer0_outputs(7887) <= a or b;
    layer0_outputs(7888) <= b;
    layer0_outputs(7889) <= b and not a;
    layer0_outputs(7890) <= a xor b;
    layer0_outputs(7891) <= not a or b;
    layer0_outputs(7892) <= not b;
    layer0_outputs(7893) <= not (a or b);
    layer0_outputs(7894) <= not (a or b);
    layer0_outputs(7895) <= not a;
    layer0_outputs(7896) <= not b;
    layer0_outputs(7897) <= a;
    layer0_outputs(7898) <= a;
    layer0_outputs(7899) <= a or b;
    layer0_outputs(7900) <= '0';
    layer0_outputs(7901) <= a or b;
    layer0_outputs(7902) <= a xor b;
    layer0_outputs(7903) <= a xor b;
    layer0_outputs(7904) <= a or b;
    layer0_outputs(7905) <= not (a and b);
    layer0_outputs(7906) <= '1';
    layer0_outputs(7907) <= not (a xor b);
    layer0_outputs(7908) <= a and not b;
    layer0_outputs(7909) <= a;
    layer0_outputs(7910) <= a or b;
    layer0_outputs(7911) <= not (a and b);
    layer0_outputs(7912) <= a or b;
    layer0_outputs(7913) <= a and not b;
    layer0_outputs(7914) <= b;
    layer0_outputs(7915) <= not (a xor b);
    layer0_outputs(7916) <= a and not b;
    layer0_outputs(7917) <= a or b;
    layer0_outputs(7918) <= not (a xor b);
    layer0_outputs(7919) <= not a or b;
    layer0_outputs(7920) <= not a or b;
    layer0_outputs(7921) <= not (a and b);
    layer0_outputs(7922) <= a xor b;
    layer0_outputs(7923) <= not (a and b);
    layer0_outputs(7924) <= not b;
    layer0_outputs(7925) <= not (a and b);
    layer0_outputs(7926) <= not b or a;
    layer0_outputs(7927) <= not a or b;
    layer0_outputs(7928) <= not b;
    layer0_outputs(7929) <= a and not b;
    layer0_outputs(7930) <= not b;
    layer0_outputs(7931) <= b;
    layer0_outputs(7932) <= a xor b;
    layer0_outputs(7933) <= a;
    layer0_outputs(7934) <= not b or a;
    layer0_outputs(7935) <= not b or a;
    layer0_outputs(7936) <= not a or b;
    layer0_outputs(7937) <= not b or a;
    layer0_outputs(7938) <= not (a xor b);
    layer0_outputs(7939) <= a or b;
    layer0_outputs(7940) <= not a or b;
    layer0_outputs(7941) <= not (a xor b);
    layer0_outputs(7942) <= not b;
    layer0_outputs(7943) <= a and not b;
    layer0_outputs(7944) <= a;
    layer0_outputs(7945) <= not (a or b);
    layer0_outputs(7946) <= a xor b;
    layer0_outputs(7947) <= a or b;
    layer0_outputs(7948) <= not b;
    layer0_outputs(7949) <= b and not a;
    layer0_outputs(7950) <= not a or b;
    layer0_outputs(7951) <= not b or a;
    layer0_outputs(7952) <= not b;
    layer0_outputs(7953) <= not a or b;
    layer0_outputs(7954) <= not a;
    layer0_outputs(7955) <= a or b;
    layer0_outputs(7956) <= not (a or b);
    layer0_outputs(7957) <= not (a or b);
    layer0_outputs(7958) <= a xor b;
    layer0_outputs(7959) <= not (a or b);
    layer0_outputs(7960) <= not (a or b);
    layer0_outputs(7961) <= b;
    layer0_outputs(7962) <= a or b;
    layer0_outputs(7963) <= '1';
    layer0_outputs(7964) <= a xor b;
    layer0_outputs(7965) <= b and not a;
    layer0_outputs(7966) <= not a or b;
    layer0_outputs(7967) <= '0';
    layer0_outputs(7968) <= not (a or b);
    layer0_outputs(7969) <= a and not b;
    layer0_outputs(7970) <= a or b;
    layer0_outputs(7971) <= a and not b;
    layer0_outputs(7972) <= not (a xor b);
    layer0_outputs(7973) <= a xor b;
    layer0_outputs(7974) <= not b or a;
    layer0_outputs(7975) <= not b or a;
    layer0_outputs(7976) <= '1';
    layer0_outputs(7977) <= a;
    layer0_outputs(7978) <= not a;
    layer0_outputs(7979) <= a and b;
    layer0_outputs(7980) <= a and not b;
    layer0_outputs(7981) <= not (a xor b);
    layer0_outputs(7982) <= a;
    layer0_outputs(7983) <= not b;
    layer0_outputs(7984) <= b;
    layer0_outputs(7985) <= not a;
    layer0_outputs(7986) <= not (a or b);
    layer0_outputs(7987) <= b;
    layer0_outputs(7988) <= not (a xor b);
    layer0_outputs(7989) <= not (a or b);
    layer0_outputs(7990) <= b and not a;
    layer0_outputs(7991) <= a xor b;
    layer0_outputs(7992) <= a and not b;
    layer0_outputs(7993) <= not (a or b);
    layer0_outputs(7994) <= not (a or b);
    layer0_outputs(7995) <= not (a xor b);
    layer0_outputs(7996) <= a;
    layer0_outputs(7997) <= a or b;
    layer0_outputs(7998) <= not a;
    layer0_outputs(7999) <= a xor b;
    layer0_outputs(8000) <= not (a and b);
    layer0_outputs(8001) <= a or b;
    layer0_outputs(8002) <= a xor b;
    layer0_outputs(8003) <= '1';
    layer0_outputs(8004) <= a or b;
    layer0_outputs(8005) <= not a;
    layer0_outputs(8006) <= a;
    layer0_outputs(8007) <= a and b;
    layer0_outputs(8008) <= not (a xor b);
    layer0_outputs(8009) <= b;
    layer0_outputs(8010) <= '1';
    layer0_outputs(8011) <= a xor b;
    layer0_outputs(8012) <= a or b;
    layer0_outputs(8013) <= not (a or b);
    layer0_outputs(8014) <= not a;
    layer0_outputs(8015) <= a or b;
    layer0_outputs(8016) <= a xor b;
    layer0_outputs(8017) <= a or b;
    layer0_outputs(8018) <= not a;
    layer0_outputs(8019) <= not a;
    layer0_outputs(8020) <= not (a or b);
    layer0_outputs(8021) <= not a;
    layer0_outputs(8022) <= not (a or b);
    layer0_outputs(8023) <= '0';
    layer0_outputs(8024) <= not a;
    layer0_outputs(8025) <= a and not b;
    layer0_outputs(8026) <= a xor b;
    layer0_outputs(8027) <= a and not b;
    layer0_outputs(8028) <= not a or b;
    layer0_outputs(8029) <= a or b;
    layer0_outputs(8030) <= not a;
    layer0_outputs(8031) <= not a;
    layer0_outputs(8032) <= not (a and b);
    layer0_outputs(8033) <= not (a or b);
    layer0_outputs(8034) <= not b;
    layer0_outputs(8035) <= not (a xor b);
    layer0_outputs(8036) <= not (a or b);
    layer0_outputs(8037) <= a and not b;
    layer0_outputs(8038) <= not (a or b);
    layer0_outputs(8039) <= not (a xor b);
    layer0_outputs(8040) <= a or b;
    layer0_outputs(8041) <= a and b;
    layer0_outputs(8042) <= not b or a;
    layer0_outputs(8043) <= not (a or b);
    layer0_outputs(8044) <= not a or b;
    layer0_outputs(8045) <= not b or a;
    layer0_outputs(8046) <= not (a xor b);
    layer0_outputs(8047) <= not (a or b);
    layer0_outputs(8048) <= a or b;
    layer0_outputs(8049) <= a or b;
    layer0_outputs(8050) <= a or b;
    layer0_outputs(8051) <= a;
    layer0_outputs(8052) <= not b or a;
    layer0_outputs(8053) <= a or b;
    layer0_outputs(8054) <= not (a xor b);
    layer0_outputs(8055) <= not b;
    layer0_outputs(8056) <= a xor b;
    layer0_outputs(8057) <= '0';
    layer0_outputs(8058) <= not a or b;
    layer0_outputs(8059) <= not a;
    layer0_outputs(8060) <= not (a and b);
    layer0_outputs(8061) <= not (a xor b);
    layer0_outputs(8062) <= not (a xor b);
    layer0_outputs(8063) <= a and b;
    layer0_outputs(8064) <= not b;
    layer0_outputs(8065) <= b and not a;
    layer0_outputs(8066) <= b;
    layer0_outputs(8067) <= a and not b;
    layer0_outputs(8068) <= '0';
    layer0_outputs(8069) <= not b or a;
    layer0_outputs(8070) <= b;
    layer0_outputs(8071) <= a and not b;
    layer0_outputs(8072) <= b and not a;
    layer0_outputs(8073) <= a and not b;
    layer0_outputs(8074) <= b;
    layer0_outputs(8075) <= a and not b;
    layer0_outputs(8076) <= not a;
    layer0_outputs(8077) <= not b;
    layer0_outputs(8078) <= b and not a;
    layer0_outputs(8079) <= a and not b;
    layer0_outputs(8080) <= not a or b;
    layer0_outputs(8081) <= not (a or b);
    layer0_outputs(8082) <= not a or b;
    layer0_outputs(8083) <= '1';
    layer0_outputs(8084) <= a or b;
    layer0_outputs(8085) <= not b or a;
    layer0_outputs(8086) <= not (a xor b);
    layer0_outputs(8087) <= not (a or b);
    layer0_outputs(8088) <= not (a or b);
    layer0_outputs(8089) <= not (a xor b);
    layer0_outputs(8090) <= b;
    layer0_outputs(8091) <= a xor b;
    layer0_outputs(8092) <= a xor b;
    layer0_outputs(8093) <= not (a xor b);
    layer0_outputs(8094) <= not (a or b);
    layer0_outputs(8095) <= not a;
    layer0_outputs(8096) <= b and not a;
    layer0_outputs(8097) <= not a or b;
    layer0_outputs(8098) <= a and not b;
    layer0_outputs(8099) <= b and not a;
    layer0_outputs(8100) <= not (a xor b);
    layer0_outputs(8101) <= a and not b;
    layer0_outputs(8102) <= a;
    layer0_outputs(8103) <= not a;
    layer0_outputs(8104) <= not a;
    layer0_outputs(8105) <= a or b;
    layer0_outputs(8106) <= not (a or b);
    layer0_outputs(8107) <= b;
    layer0_outputs(8108) <= not (a or b);
    layer0_outputs(8109) <= b;
    layer0_outputs(8110) <= '0';
    layer0_outputs(8111) <= b;
    layer0_outputs(8112) <= a xor b;
    layer0_outputs(8113) <= not a or b;
    layer0_outputs(8114) <= not a or b;
    layer0_outputs(8115) <= not (a or b);
    layer0_outputs(8116) <= a and not b;
    layer0_outputs(8117) <= b;
    layer0_outputs(8118) <= a or b;
    layer0_outputs(8119) <= '0';
    layer0_outputs(8120) <= a xor b;
    layer0_outputs(8121) <= b;
    layer0_outputs(8122) <= not b;
    layer0_outputs(8123) <= not b or a;
    layer0_outputs(8124) <= not (a or b);
    layer0_outputs(8125) <= a xor b;
    layer0_outputs(8126) <= a or b;
    layer0_outputs(8127) <= not a or b;
    layer0_outputs(8128) <= not (a or b);
    layer0_outputs(8129) <= not b;
    layer0_outputs(8130) <= a or b;
    layer0_outputs(8131) <= b and not a;
    layer0_outputs(8132) <= a xor b;
    layer0_outputs(8133) <= not b;
    layer0_outputs(8134) <= b;
    layer0_outputs(8135) <= not b;
    layer0_outputs(8136) <= a and not b;
    layer0_outputs(8137) <= not (a or b);
    layer0_outputs(8138) <= b;
    layer0_outputs(8139) <= a xor b;
    layer0_outputs(8140) <= not a or b;
    layer0_outputs(8141) <= not (a or b);
    layer0_outputs(8142) <= a and b;
    layer0_outputs(8143) <= not (a or b);
    layer0_outputs(8144) <= a and not b;
    layer0_outputs(8145) <= not a or b;
    layer0_outputs(8146) <= b and not a;
    layer0_outputs(8147) <= not (a xor b);
    layer0_outputs(8148) <= b and not a;
    layer0_outputs(8149) <= a;
    layer0_outputs(8150) <= not b;
    layer0_outputs(8151) <= a;
    layer0_outputs(8152) <= not (a or b);
    layer0_outputs(8153) <= b;
    layer0_outputs(8154) <= not a;
    layer0_outputs(8155) <= not (a or b);
    layer0_outputs(8156) <= a;
    layer0_outputs(8157) <= not (a xor b);
    layer0_outputs(8158) <= not a or b;
    layer0_outputs(8159) <= not a;
    layer0_outputs(8160) <= a xor b;
    layer0_outputs(8161) <= a or b;
    layer0_outputs(8162) <= a or b;
    layer0_outputs(8163) <= a or b;
    layer0_outputs(8164) <= '1';
    layer0_outputs(8165) <= not a;
    layer0_outputs(8166) <= not b;
    layer0_outputs(8167) <= not b or a;
    layer0_outputs(8168) <= a and not b;
    layer0_outputs(8169) <= a;
    layer0_outputs(8170) <= not (a or b);
    layer0_outputs(8171) <= not (a or b);
    layer0_outputs(8172) <= a or b;
    layer0_outputs(8173) <= not (a or b);
    layer0_outputs(8174) <= a;
    layer0_outputs(8175) <= not (a xor b);
    layer0_outputs(8176) <= a or b;
    layer0_outputs(8177) <= not (a and b);
    layer0_outputs(8178) <= a and not b;
    layer0_outputs(8179) <= a xor b;
    layer0_outputs(8180) <= a;
    layer0_outputs(8181) <= a and not b;
    layer0_outputs(8182) <= a or b;
    layer0_outputs(8183) <= b;
    layer0_outputs(8184) <= not (a and b);
    layer0_outputs(8185) <= not a;
    layer0_outputs(8186) <= '1';
    layer0_outputs(8187) <= b and not a;
    layer0_outputs(8188) <= not a;
    layer0_outputs(8189) <= a xor b;
    layer0_outputs(8190) <= a xor b;
    layer0_outputs(8191) <= a and not b;
    layer0_outputs(8192) <= a xor b;
    layer0_outputs(8193) <= a;
    layer0_outputs(8194) <= a or b;
    layer0_outputs(8195) <= not (a and b);
    layer0_outputs(8196) <= b and not a;
    layer0_outputs(8197) <= not (a and b);
    layer0_outputs(8198) <= a or b;
    layer0_outputs(8199) <= b and not a;
    layer0_outputs(8200) <= b;
    layer0_outputs(8201) <= a;
    layer0_outputs(8202) <= not (a or b);
    layer0_outputs(8203) <= a xor b;
    layer0_outputs(8204) <= not a or b;
    layer0_outputs(8205) <= not a;
    layer0_outputs(8206) <= not b or a;
    layer0_outputs(8207) <= a or b;
    layer0_outputs(8208) <= not a;
    layer0_outputs(8209) <= not (a or b);
    layer0_outputs(8210) <= a or b;
    layer0_outputs(8211) <= not b;
    layer0_outputs(8212) <= b and not a;
    layer0_outputs(8213) <= a or b;
    layer0_outputs(8214) <= not (a or b);
    layer0_outputs(8215) <= not b or a;
    layer0_outputs(8216) <= b and not a;
    layer0_outputs(8217) <= not b or a;
    layer0_outputs(8218) <= not a or b;
    layer0_outputs(8219) <= '1';
    layer0_outputs(8220) <= b;
    layer0_outputs(8221) <= a or b;
    layer0_outputs(8222) <= a;
    layer0_outputs(8223) <= a and not b;
    layer0_outputs(8224) <= b;
    layer0_outputs(8225) <= a;
    layer0_outputs(8226) <= a xor b;
    layer0_outputs(8227) <= not (a xor b);
    layer0_outputs(8228) <= not a;
    layer0_outputs(8229) <= b and not a;
    layer0_outputs(8230) <= '1';
    layer0_outputs(8231) <= a xor b;
    layer0_outputs(8232) <= a xor b;
    layer0_outputs(8233) <= not (a or b);
    layer0_outputs(8234) <= '1';
    layer0_outputs(8235) <= not a;
    layer0_outputs(8236) <= a or b;
    layer0_outputs(8237) <= not b;
    layer0_outputs(8238) <= a or b;
    layer0_outputs(8239) <= not (a or b);
    layer0_outputs(8240) <= a xor b;
    layer0_outputs(8241) <= not b or a;
    layer0_outputs(8242) <= a;
    layer0_outputs(8243) <= a xor b;
    layer0_outputs(8244) <= not b or a;
    layer0_outputs(8245) <= b and not a;
    layer0_outputs(8246) <= a xor b;
    layer0_outputs(8247) <= not b;
    layer0_outputs(8248) <= a or b;
    layer0_outputs(8249) <= not (a or b);
    layer0_outputs(8250) <= not b or a;
    layer0_outputs(8251) <= not a or b;
    layer0_outputs(8252) <= a xor b;
    layer0_outputs(8253) <= a or b;
    layer0_outputs(8254) <= a;
    layer0_outputs(8255) <= not (a or b);
    layer0_outputs(8256) <= a and b;
    layer0_outputs(8257) <= a or b;
    layer0_outputs(8258) <= a or b;
    layer0_outputs(8259) <= not (a or b);
    layer0_outputs(8260) <= not a;
    layer0_outputs(8261) <= not a or b;
    layer0_outputs(8262) <= a or b;
    layer0_outputs(8263) <= b;
    layer0_outputs(8264) <= '1';
    layer0_outputs(8265) <= a;
    layer0_outputs(8266) <= b and not a;
    layer0_outputs(8267) <= not (a or b);
    layer0_outputs(8268) <= not a;
    layer0_outputs(8269) <= not (a or b);
    layer0_outputs(8270) <= a or b;
    layer0_outputs(8271) <= a or b;
    layer0_outputs(8272) <= a or b;
    layer0_outputs(8273) <= a xor b;
    layer0_outputs(8274) <= not (a and b);
    layer0_outputs(8275) <= b and not a;
    layer0_outputs(8276) <= b and not a;
    layer0_outputs(8277) <= a or b;
    layer0_outputs(8278) <= not b;
    layer0_outputs(8279) <= not b or a;
    layer0_outputs(8280) <= not a or b;
    layer0_outputs(8281) <= not (a or b);
    layer0_outputs(8282) <= not b;
    layer0_outputs(8283) <= not (a xor b);
    layer0_outputs(8284) <= not (a and b);
    layer0_outputs(8285) <= not a or b;
    layer0_outputs(8286) <= a xor b;
    layer0_outputs(8287) <= not b;
    layer0_outputs(8288) <= not b;
    layer0_outputs(8289) <= a;
    layer0_outputs(8290) <= a and b;
    layer0_outputs(8291) <= not (a or b);
    layer0_outputs(8292) <= a and not b;
    layer0_outputs(8293) <= not (a or b);
    layer0_outputs(8294) <= a or b;
    layer0_outputs(8295) <= b and not a;
    layer0_outputs(8296) <= a xor b;
    layer0_outputs(8297) <= a;
    layer0_outputs(8298) <= not (a and b);
    layer0_outputs(8299) <= not a or b;
    layer0_outputs(8300) <= not (a or b);
    layer0_outputs(8301) <= not a;
    layer0_outputs(8302) <= not (a xor b);
    layer0_outputs(8303) <= not (a or b);
    layer0_outputs(8304) <= not a;
    layer0_outputs(8305) <= a or b;
    layer0_outputs(8306) <= not (a or b);
    layer0_outputs(8307) <= a;
    layer0_outputs(8308) <= a or b;
    layer0_outputs(8309) <= a xor b;
    layer0_outputs(8310) <= not (a xor b);
    layer0_outputs(8311) <= not (a xor b);
    layer0_outputs(8312) <= '1';
    layer0_outputs(8313) <= not (a xor b);
    layer0_outputs(8314) <= not b or a;
    layer0_outputs(8315) <= a and not b;
    layer0_outputs(8316) <= not a;
    layer0_outputs(8317) <= not a or b;
    layer0_outputs(8318) <= not b;
    layer0_outputs(8319) <= not (a xor b);
    layer0_outputs(8320) <= not b;
    layer0_outputs(8321) <= not (a or b);
    layer0_outputs(8322) <= not (a or b);
    layer0_outputs(8323) <= not (a or b);
    layer0_outputs(8324) <= not a;
    layer0_outputs(8325) <= a and not b;
    layer0_outputs(8326) <= a xor b;
    layer0_outputs(8327) <= a and b;
    layer0_outputs(8328) <= not a or b;
    layer0_outputs(8329) <= not b or a;
    layer0_outputs(8330) <= b;
    layer0_outputs(8331) <= not (a xor b);
    layer0_outputs(8332) <= not (a or b);
    layer0_outputs(8333) <= not (a and b);
    layer0_outputs(8334) <= not (a xor b);
    layer0_outputs(8335) <= a or b;
    layer0_outputs(8336) <= not b;
    layer0_outputs(8337) <= a xor b;
    layer0_outputs(8338) <= not (a or b);
    layer0_outputs(8339) <= not (a or b);
    layer0_outputs(8340) <= a or b;
    layer0_outputs(8341) <= a;
    layer0_outputs(8342) <= a or b;
    layer0_outputs(8343) <= b and not a;
    layer0_outputs(8344) <= not a;
    layer0_outputs(8345) <= a xor b;
    layer0_outputs(8346) <= a;
    layer0_outputs(8347) <= not b;
    layer0_outputs(8348) <= not b;
    layer0_outputs(8349) <= not b or a;
    layer0_outputs(8350) <= b and not a;
    layer0_outputs(8351) <= not b;
    layer0_outputs(8352) <= a and b;
    layer0_outputs(8353) <= a xor b;
    layer0_outputs(8354) <= not b;
    layer0_outputs(8355) <= not b;
    layer0_outputs(8356) <= not (a or b);
    layer0_outputs(8357) <= b;
    layer0_outputs(8358) <= not (a or b);
    layer0_outputs(8359) <= not b or a;
    layer0_outputs(8360) <= a xor b;
    layer0_outputs(8361) <= not b;
    layer0_outputs(8362) <= not b;
    layer0_outputs(8363) <= a or b;
    layer0_outputs(8364) <= '1';
    layer0_outputs(8365) <= b and not a;
    layer0_outputs(8366) <= a or b;
    layer0_outputs(8367) <= not (a xor b);
    layer0_outputs(8368) <= a or b;
    layer0_outputs(8369) <= a or b;
    layer0_outputs(8370) <= not b;
    layer0_outputs(8371) <= a and b;
    layer0_outputs(8372) <= not b;
    layer0_outputs(8373) <= not (a or b);
    layer0_outputs(8374) <= not (a and b);
    layer0_outputs(8375) <= not a or b;
    layer0_outputs(8376) <= not (a xor b);
    layer0_outputs(8377) <= not (a xor b);
    layer0_outputs(8378) <= not a or b;
    layer0_outputs(8379) <= not a;
    layer0_outputs(8380) <= not (a xor b);
    layer0_outputs(8381) <= not (a xor b);
    layer0_outputs(8382) <= not (a and b);
    layer0_outputs(8383) <= b;
    layer0_outputs(8384) <= not a;
    layer0_outputs(8385) <= not (a and b);
    layer0_outputs(8386) <= a or b;
    layer0_outputs(8387) <= a and not b;
    layer0_outputs(8388) <= not (a xor b);
    layer0_outputs(8389) <= a xor b;
    layer0_outputs(8390) <= a and not b;
    layer0_outputs(8391) <= '1';
    layer0_outputs(8392) <= '0';
    layer0_outputs(8393) <= a or b;
    layer0_outputs(8394) <= not a or b;
    layer0_outputs(8395) <= not (a xor b);
    layer0_outputs(8396) <= a xor b;
    layer0_outputs(8397) <= not a;
    layer0_outputs(8398) <= not b;
    layer0_outputs(8399) <= a;
    layer0_outputs(8400) <= not a or b;
    layer0_outputs(8401) <= a xor b;
    layer0_outputs(8402) <= a;
    layer0_outputs(8403) <= a;
    layer0_outputs(8404) <= not b or a;
    layer0_outputs(8405) <= not a;
    layer0_outputs(8406) <= not (a xor b);
    layer0_outputs(8407) <= a or b;
    layer0_outputs(8408) <= not a or b;
    layer0_outputs(8409) <= a;
    layer0_outputs(8410) <= not (a and b);
    layer0_outputs(8411) <= not (a or b);
    layer0_outputs(8412) <= not b or a;
    layer0_outputs(8413) <= b and not a;
    layer0_outputs(8414) <= b;
    layer0_outputs(8415) <= a or b;
    layer0_outputs(8416) <= b;
    layer0_outputs(8417) <= b and not a;
    layer0_outputs(8418) <= a and b;
    layer0_outputs(8419) <= not b or a;
    layer0_outputs(8420) <= not (a or b);
    layer0_outputs(8421) <= a and b;
    layer0_outputs(8422) <= not b;
    layer0_outputs(8423) <= a or b;
    layer0_outputs(8424) <= not b;
    layer0_outputs(8425) <= a or b;
    layer0_outputs(8426) <= not (a xor b);
    layer0_outputs(8427) <= a and b;
    layer0_outputs(8428) <= b and not a;
    layer0_outputs(8429) <= not a or b;
    layer0_outputs(8430) <= a and not b;
    layer0_outputs(8431) <= a and not b;
    layer0_outputs(8432) <= a;
    layer0_outputs(8433) <= not a;
    layer0_outputs(8434) <= a or b;
    layer0_outputs(8435) <= not (a and b);
    layer0_outputs(8436) <= '0';
    layer0_outputs(8437) <= a or b;
    layer0_outputs(8438) <= b;
    layer0_outputs(8439) <= b and not a;
    layer0_outputs(8440) <= not b;
    layer0_outputs(8441) <= b;
    layer0_outputs(8442) <= a or b;
    layer0_outputs(8443) <= a xor b;
    layer0_outputs(8444) <= a;
    layer0_outputs(8445) <= not a;
    layer0_outputs(8446) <= not b;
    layer0_outputs(8447) <= a or b;
    layer0_outputs(8448) <= not (a xor b);
    layer0_outputs(8449) <= not a or b;
    layer0_outputs(8450) <= a xor b;
    layer0_outputs(8451) <= not b or a;
    layer0_outputs(8452) <= not (a xor b);
    layer0_outputs(8453) <= not b;
    layer0_outputs(8454) <= b and not a;
    layer0_outputs(8455) <= b and not a;
    layer0_outputs(8456) <= not (a xor b);
    layer0_outputs(8457) <= a and b;
    layer0_outputs(8458) <= a and b;
    layer0_outputs(8459) <= a;
    layer0_outputs(8460) <= a or b;
    layer0_outputs(8461) <= a and not b;
    layer0_outputs(8462) <= a xor b;
    layer0_outputs(8463) <= not (a or b);
    layer0_outputs(8464) <= b;
    layer0_outputs(8465) <= b;
    layer0_outputs(8466) <= b and not a;
    layer0_outputs(8467) <= a xor b;
    layer0_outputs(8468) <= not a or b;
    layer0_outputs(8469) <= not (a and b);
    layer0_outputs(8470) <= a;
    layer0_outputs(8471) <= a and not b;
    layer0_outputs(8472) <= b;
    layer0_outputs(8473) <= not b or a;
    layer0_outputs(8474) <= '0';
    layer0_outputs(8475) <= b;
    layer0_outputs(8476) <= not (a and b);
    layer0_outputs(8477) <= not a or b;
    layer0_outputs(8478) <= not (a xor b);
    layer0_outputs(8479) <= not (a xor b);
    layer0_outputs(8480) <= not a;
    layer0_outputs(8481) <= a or b;
    layer0_outputs(8482) <= not (a or b);
    layer0_outputs(8483) <= not a;
    layer0_outputs(8484) <= a or b;
    layer0_outputs(8485) <= not (a and b);
    layer0_outputs(8486) <= a;
    layer0_outputs(8487) <= not (a or b);
    layer0_outputs(8488) <= a or b;
    layer0_outputs(8489) <= '1';
    layer0_outputs(8490) <= a xor b;
    layer0_outputs(8491) <= a or b;
    layer0_outputs(8492) <= not (a or b);
    layer0_outputs(8493) <= a xor b;
    layer0_outputs(8494) <= a xor b;
    layer0_outputs(8495) <= not (a and b);
    layer0_outputs(8496) <= a or b;
    layer0_outputs(8497) <= b and not a;
    layer0_outputs(8498) <= a xor b;
    layer0_outputs(8499) <= a or b;
    layer0_outputs(8500) <= not b or a;
    layer0_outputs(8501) <= a or b;
    layer0_outputs(8502) <= not a;
    layer0_outputs(8503) <= b;
    layer0_outputs(8504) <= not (a xor b);
    layer0_outputs(8505) <= not (a xor b);
    layer0_outputs(8506) <= not a;
    layer0_outputs(8507) <= b and not a;
    layer0_outputs(8508) <= not a or b;
    layer0_outputs(8509) <= not a;
    layer0_outputs(8510) <= a;
    layer0_outputs(8511) <= not (a xor b);
    layer0_outputs(8512) <= b and not a;
    layer0_outputs(8513) <= b;
    layer0_outputs(8514) <= b and not a;
    layer0_outputs(8515) <= not a or b;
    layer0_outputs(8516) <= a or b;
    layer0_outputs(8517) <= a and b;
    layer0_outputs(8518) <= not (a xor b);
    layer0_outputs(8519) <= not (a or b);
    layer0_outputs(8520) <= not a or b;
    layer0_outputs(8521) <= not (a or b);
    layer0_outputs(8522) <= b and not a;
    layer0_outputs(8523) <= not (a or b);
    layer0_outputs(8524) <= not a or b;
    layer0_outputs(8525) <= b;
    layer0_outputs(8526) <= not a or b;
    layer0_outputs(8527) <= not a;
    layer0_outputs(8528) <= b;
    layer0_outputs(8529) <= not b;
    layer0_outputs(8530) <= not (a or b);
    layer0_outputs(8531) <= a xor b;
    layer0_outputs(8532) <= not (a xor b);
    layer0_outputs(8533) <= not (a or b);
    layer0_outputs(8534) <= a xor b;
    layer0_outputs(8535) <= a or b;
    layer0_outputs(8536) <= not (a or b);
    layer0_outputs(8537) <= b;
    layer0_outputs(8538) <= not (a or b);
    layer0_outputs(8539) <= not (a and b);
    layer0_outputs(8540) <= b and not a;
    layer0_outputs(8541) <= not b;
    layer0_outputs(8542) <= a xor b;
    layer0_outputs(8543) <= a or b;
    layer0_outputs(8544) <= not b or a;
    layer0_outputs(8545) <= a or b;
    layer0_outputs(8546) <= not (a and b);
    layer0_outputs(8547) <= a or b;
    layer0_outputs(8548) <= not b or a;
    layer0_outputs(8549) <= b and not a;
    layer0_outputs(8550) <= a or b;
    layer0_outputs(8551) <= not (a or b);
    layer0_outputs(8552) <= not a;
    layer0_outputs(8553) <= '0';
    layer0_outputs(8554) <= not a;
    layer0_outputs(8555) <= not a or b;
    layer0_outputs(8556) <= '0';
    layer0_outputs(8557) <= not b;
    layer0_outputs(8558) <= a and not b;
    layer0_outputs(8559) <= not b or a;
    layer0_outputs(8560) <= not a or b;
    layer0_outputs(8561) <= not (a or b);
    layer0_outputs(8562) <= '1';
    layer0_outputs(8563) <= not b or a;
    layer0_outputs(8564) <= not a or b;
    layer0_outputs(8565) <= not (a xor b);
    layer0_outputs(8566) <= '1';
    layer0_outputs(8567) <= not (a or b);
    layer0_outputs(8568) <= not (a xor b);
    layer0_outputs(8569) <= not (a or b);
    layer0_outputs(8570) <= not (a or b);
    layer0_outputs(8571) <= '1';
    layer0_outputs(8572) <= a or b;
    layer0_outputs(8573) <= not b or a;
    layer0_outputs(8574) <= b and not a;
    layer0_outputs(8575) <= a or b;
    layer0_outputs(8576) <= a or b;
    layer0_outputs(8577) <= a and not b;
    layer0_outputs(8578) <= a or b;
    layer0_outputs(8579) <= a or b;
    layer0_outputs(8580) <= not b or a;
    layer0_outputs(8581) <= not (a xor b);
    layer0_outputs(8582) <= not a;
    layer0_outputs(8583) <= a or b;
    layer0_outputs(8584) <= not (a or b);
    layer0_outputs(8585) <= a or b;
    layer0_outputs(8586) <= not b;
    layer0_outputs(8587) <= '1';
    layer0_outputs(8588) <= a and not b;
    layer0_outputs(8589) <= not a;
    layer0_outputs(8590) <= a and not b;
    layer0_outputs(8591) <= b and not a;
    layer0_outputs(8592) <= a xor b;
    layer0_outputs(8593) <= not b or a;
    layer0_outputs(8594) <= '1';
    layer0_outputs(8595) <= a and b;
    layer0_outputs(8596) <= not (a or b);
    layer0_outputs(8597) <= not b or a;
    layer0_outputs(8598) <= b;
    layer0_outputs(8599) <= not a or b;
    layer0_outputs(8600) <= a or b;
    layer0_outputs(8601) <= '0';
    layer0_outputs(8602) <= not b or a;
    layer0_outputs(8603) <= not (a or b);
    layer0_outputs(8604) <= a;
    layer0_outputs(8605) <= not a or b;
    layer0_outputs(8606) <= not a or b;
    layer0_outputs(8607) <= b;
    layer0_outputs(8608) <= not b;
    layer0_outputs(8609) <= a and not b;
    layer0_outputs(8610) <= not (a or b);
    layer0_outputs(8611) <= b and not a;
    layer0_outputs(8612) <= not b or a;
    layer0_outputs(8613) <= a and not b;
    layer0_outputs(8614) <= a xor b;
    layer0_outputs(8615) <= a xor b;
    layer0_outputs(8616) <= not a;
    layer0_outputs(8617) <= a xor b;
    layer0_outputs(8618) <= not b;
    layer0_outputs(8619) <= a xor b;
    layer0_outputs(8620) <= not b;
    layer0_outputs(8621) <= a xor b;
    layer0_outputs(8622) <= a xor b;
    layer0_outputs(8623) <= not a;
    layer0_outputs(8624) <= not a;
    layer0_outputs(8625) <= a or b;
    layer0_outputs(8626) <= not (a or b);
    layer0_outputs(8627) <= '0';
    layer0_outputs(8628) <= a or b;
    layer0_outputs(8629) <= not (a xor b);
    layer0_outputs(8630) <= not b;
    layer0_outputs(8631) <= a xor b;
    layer0_outputs(8632) <= b;
    layer0_outputs(8633) <= a or b;
    layer0_outputs(8634) <= not b;
    layer0_outputs(8635) <= not (a or b);
    layer0_outputs(8636) <= a xor b;
    layer0_outputs(8637) <= a or b;
    layer0_outputs(8638) <= not (a or b);
    layer0_outputs(8639) <= a or b;
    layer0_outputs(8640) <= not b;
    layer0_outputs(8641) <= b;
    layer0_outputs(8642) <= b;
    layer0_outputs(8643) <= not (a xor b);
    layer0_outputs(8644) <= not (a or b);
    layer0_outputs(8645) <= not (a xor b);
    layer0_outputs(8646) <= not a or b;
    layer0_outputs(8647) <= not b or a;
    layer0_outputs(8648) <= not (a or b);
    layer0_outputs(8649) <= not b or a;
    layer0_outputs(8650) <= not (a or b);
    layer0_outputs(8651) <= not (a or b);
    layer0_outputs(8652) <= b;
    layer0_outputs(8653) <= not (a and b);
    layer0_outputs(8654) <= a;
    layer0_outputs(8655) <= not a;
    layer0_outputs(8656) <= not a;
    layer0_outputs(8657) <= '0';
    layer0_outputs(8658) <= a and not b;
    layer0_outputs(8659) <= not (a or b);
    layer0_outputs(8660) <= not (a or b);
    layer0_outputs(8661) <= not (a xor b);
    layer0_outputs(8662) <= not (a or b);
    layer0_outputs(8663) <= not (a or b);
    layer0_outputs(8664) <= a or b;
    layer0_outputs(8665) <= b and not a;
    layer0_outputs(8666) <= not b or a;
    layer0_outputs(8667) <= not b or a;
    layer0_outputs(8668) <= not a or b;
    layer0_outputs(8669) <= a or b;
    layer0_outputs(8670) <= a xor b;
    layer0_outputs(8671) <= a and b;
    layer0_outputs(8672) <= not b;
    layer0_outputs(8673) <= a;
    layer0_outputs(8674) <= a or b;
    layer0_outputs(8675) <= a or b;
    layer0_outputs(8676) <= '0';
    layer0_outputs(8677) <= a and not b;
    layer0_outputs(8678) <= a xor b;
    layer0_outputs(8679) <= a;
    layer0_outputs(8680) <= a xor b;
    layer0_outputs(8681) <= not a;
    layer0_outputs(8682) <= a or b;
    layer0_outputs(8683) <= a or b;
    layer0_outputs(8684) <= a xor b;
    layer0_outputs(8685) <= b;
    layer0_outputs(8686) <= a and not b;
    layer0_outputs(8687) <= b and not a;
    layer0_outputs(8688) <= not a or b;
    layer0_outputs(8689) <= b;
    layer0_outputs(8690) <= b;
    layer0_outputs(8691) <= b and not a;
    layer0_outputs(8692) <= not (a and b);
    layer0_outputs(8693) <= not (a xor b);
    layer0_outputs(8694) <= b;
    layer0_outputs(8695) <= a xor b;
    layer0_outputs(8696) <= not a;
    layer0_outputs(8697) <= a xor b;
    layer0_outputs(8698) <= a xor b;
    layer0_outputs(8699) <= a xor b;
    layer0_outputs(8700) <= not (a or b);
    layer0_outputs(8701) <= not (a or b);
    layer0_outputs(8702) <= b and not a;
    layer0_outputs(8703) <= not (a or b);
    layer0_outputs(8704) <= a or b;
    layer0_outputs(8705) <= not a or b;
    layer0_outputs(8706) <= not a;
    layer0_outputs(8707) <= '0';
    layer0_outputs(8708) <= a or b;
    layer0_outputs(8709) <= a or b;
    layer0_outputs(8710) <= not a;
    layer0_outputs(8711) <= a and not b;
    layer0_outputs(8712) <= a or b;
    layer0_outputs(8713) <= a;
    layer0_outputs(8714) <= a or b;
    layer0_outputs(8715) <= a xor b;
    layer0_outputs(8716) <= not (a or b);
    layer0_outputs(8717) <= a xor b;
    layer0_outputs(8718) <= not a;
    layer0_outputs(8719) <= a or b;
    layer0_outputs(8720) <= b;
    layer0_outputs(8721) <= a;
    layer0_outputs(8722) <= not a or b;
    layer0_outputs(8723) <= not b;
    layer0_outputs(8724) <= a or b;
    layer0_outputs(8725) <= b;
    layer0_outputs(8726) <= b and not a;
    layer0_outputs(8727) <= not a;
    layer0_outputs(8728) <= b and not a;
    layer0_outputs(8729) <= '1';
    layer0_outputs(8730) <= not a or b;
    layer0_outputs(8731) <= a and not b;
    layer0_outputs(8732) <= not a;
    layer0_outputs(8733) <= a or b;
    layer0_outputs(8734) <= a;
    layer0_outputs(8735) <= a and b;
    layer0_outputs(8736) <= a xor b;
    layer0_outputs(8737) <= '0';
    layer0_outputs(8738) <= not a;
    layer0_outputs(8739) <= '1';
    layer0_outputs(8740) <= a;
    layer0_outputs(8741) <= not (a or b);
    layer0_outputs(8742) <= b;
    layer0_outputs(8743) <= a;
    layer0_outputs(8744) <= not b;
    layer0_outputs(8745) <= not b or a;
    layer0_outputs(8746) <= b;
    layer0_outputs(8747) <= not (a xor b);
    layer0_outputs(8748) <= not a or b;
    layer0_outputs(8749) <= not a;
    layer0_outputs(8750) <= b;
    layer0_outputs(8751) <= not (a and b);
    layer0_outputs(8752) <= a and not b;
    layer0_outputs(8753) <= not (a or b);
    layer0_outputs(8754) <= b and not a;
    layer0_outputs(8755) <= not (a or b);
    layer0_outputs(8756) <= b and not a;
    layer0_outputs(8757) <= not (a or b);
    layer0_outputs(8758) <= not (a xor b);
    layer0_outputs(8759) <= a and b;
    layer0_outputs(8760) <= a and not b;
    layer0_outputs(8761) <= not (a xor b);
    layer0_outputs(8762) <= not (a and b);
    layer0_outputs(8763) <= not b;
    layer0_outputs(8764) <= not a;
    layer0_outputs(8765) <= not b;
    layer0_outputs(8766) <= not b;
    layer0_outputs(8767) <= not a or b;
    layer0_outputs(8768) <= not (a xor b);
    layer0_outputs(8769) <= a xor b;
    layer0_outputs(8770) <= a;
    layer0_outputs(8771) <= b and not a;
    layer0_outputs(8772) <= a or b;
    layer0_outputs(8773) <= b;
    layer0_outputs(8774) <= not a;
    layer0_outputs(8775) <= '1';
    layer0_outputs(8776) <= b;
    layer0_outputs(8777) <= a xor b;
    layer0_outputs(8778) <= not a;
    layer0_outputs(8779) <= a xor b;
    layer0_outputs(8780) <= not b;
    layer0_outputs(8781) <= a;
    layer0_outputs(8782) <= a;
    layer0_outputs(8783) <= not (a and b);
    layer0_outputs(8784) <= a;
    layer0_outputs(8785) <= not (a or b);
    layer0_outputs(8786) <= a or b;
    layer0_outputs(8787) <= b and not a;
    layer0_outputs(8788) <= b;
    layer0_outputs(8789) <= a;
    layer0_outputs(8790) <= not (a or b);
    layer0_outputs(8791) <= b and not a;
    layer0_outputs(8792) <= a or b;
    layer0_outputs(8793) <= not (a or b);
    layer0_outputs(8794) <= not b;
    layer0_outputs(8795) <= b;
    layer0_outputs(8796) <= not a;
    layer0_outputs(8797) <= b and not a;
    layer0_outputs(8798) <= not a or b;
    layer0_outputs(8799) <= not (a or b);
    layer0_outputs(8800) <= b and not a;
    layer0_outputs(8801) <= not b;
    layer0_outputs(8802) <= a or b;
    layer0_outputs(8803) <= a and not b;
    layer0_outputs(8804) <= a xor b;
    layer0_outputs(8805) <= a or b;
    layer0_outputs(8806) <= a and b;
    layer0_outputs(8807) <= not (a xor b);
    layer0_outputs(8808) <= not b or a;
    layer0_outputs(8809) <= not b;
    layer0_outputs(8810) <= not a or b;
    layer0_outputs(8811) <= a or b;
    layer0_outputs(8812) <= '1';
    layer0_outputs(8813) <= a;
    layer0_outputs(8814) <= b and not a;
    layer0_outputs(8815) <= not a or b;
    layer0_outputs(8816) <= '0';
    layer0_outputs(8817) <= a or b;
    layer0_outputs(8818) <= a xor b;
    layer0_outputs(8819) <= a and b;
    layer0_outputs(8820) <= not b;
    layer0_outputs(8821) <= '1';
    layer0_outputs(8822) <= not (a or b);
    layer0_outputs(8823) <= a;
    layer0_outputs(8824) <= not (a or b);
    layer0_outputs(8825) <= a and not b;
    layer0_outputs(8826) <= a or b;
    layer0_outputs(8827) <= a or b;
    layer0_outputs(8828) <= not (a xor b);
    layer0_outputs(8829) <= a;
    layer0_outputs(8830) <= '0';
    layer0_outputs(8831) <= a;
    layer0_outputs(8832) <= a;
    layer0_outputs(8833) <= a xor b;
    layer0_outputs(8834) <= not (a xor b);
    layer0_outputs(8835) <= a xor b;
    layer0_outputs(8836) <= not (a or b);
    layer0_outputs(8837) <= not a;
    layer0_outputs(8838) <= not (a and b);
    layer0_outputs(8839) <= a xor b;
    layer0_outputs(8840) <= a xor b;
    layer0_outputs(8841) <= b;
    layer0_outputs(8842) <= a;
    layer0_outputs(8843) <= not (a or b);
    layer0_outputs(8844) <= b and not a;
    layer0_outputs(8845) <= '1';
    layer0_outputs(8846) <= not (a xor b);
    layer0_outputs(8847) <= a or b;
    layer0_outputs(8848) <= not b or a;
    layer0_outputs(8849) <= a;
    layer0_outputs(8850) <= not (a or b);
    layer0_outputs(8851) <= not (a or b);
    layer0_outputs(8852) <= b and not a;
    layer0_outputs(8853) <= not b;
    layer0_outputs(8854) <= not (a xor b);
    layer0_outputs(8855) <= not a or b;
    layer0_outputs(8856) <= not (a or b);
    layer0_outputs(8857) <= not (a or b);
    layer0_outputs(8858) <= not (a or b);
    layer0_outputs(8859) <= not (a or b);
    layer0_outputs(8860) <= a;
    layer0_outputs(8861) <= not (a xor b);
    layer0_outputs(8862) <= a or b;
    layer0_outputs(8863) <= a or b;
    layer0_outputs(8864) <= a xor b;
    layer0_outputs(8865) <= a xor b;
    layer0_outputs(8866) <= not b or a;
    layer0_outputs(8867) <= a and not b;
    layer0_outputs(8868) <= a;
    layer0_outputs(8869) <= a;
    layer0_outputs(8870) <= a and not b;
    layer0_outputs(8871) <= a or b;
    layer0_outputs(8872) <= not (a or b);
    layer0_outputs(8873) <= a xor b;
    layer0_outputs(8874) <= not (a xor b);
    layer0_outputs(8875) <= not a;
    layer0_outputs(8876) <= not (a or b);
    layer0_outputs(8877) <= not a;
    layer0_outputs(8878) <= not b or a;
    layer0_outputs(8879) <= not b;
    layer0_outputs(8880) <= not b or a;
    layer0_outputs(8881) <= not b;
    layer0_outputs(8882) <= a xor b;
    layer0_outputs(8883) <= a xor b;
    layer0_outputs(8884) <= not b or a;
    layer0_outputs(8885) <= not b or a;
    layer0_outputs(8886) <= not (a and b);
    layer0_outputs(8887) <= a xor b;
    layer0_outputs(8888) <= not (a or b);
    layer0_outputs(8889) <= not (a xor b);
    layer0_outputs(8890) <= not b or a;
    layer0_outputs(8891) <= a or b;
    layer0_outputs(8892) <= not a or b;
    layer0_outputs(8893) <= a or b;
    layer0_outputs(8894) <= a and not b;
    layer0_outputs(8895) <= not (a or b);
    layer0_outputs(8896) <= not (a and b);
    layer0_outputs(8897) <= not (a and b);
    layer0_outputs(8898) <= not a;
    layer0_outputs(8899) <= b and not a;
    layer0_outputs(8900) <= not a or b;
    layer0_outputs(8901) <= not (a or b);
    layer0_outputs(8902) <= not (a xor b);
    layer0_outputs(8903) <= not (a xor b);
    layer0_outputs(8904) <= a and not b;
    layer0_outputs(8905) <= not b;
    layer0_outputs(8906) <= not (a or b);
    layer0_outputs(8907) <= b;
    layer0_outputs(8908) <= not (a xor b);
    layer0_outputs(8909) <= not b or a;
    layer0_outputs(8910) <= a and b;
    layer0_outputs(8911) <= not (a or b);
    layer0_outputs(8912) <= not (a xor b);
    layer0_outputs(8913) <= b and not a;
    layer0_outputs(8914) <= not (a or b);
    layer0_outputs(8915) <= not a;
    layer0_outputs(8916) <= not b or a;
    layer0_outputs(8917) <= not a or b;
    layer0_outputs(8918) <= not (a xor b);
    layer0_outputs(8919) <= not (a or b);
    layer0_outputs(8920) <= not b;
    layer0_outputs(8921) <= b and not a;
    layer0_outputs(8922) <= a or b;
    layer0_outputs(8923) <= '1';
    layer0_outputs(8924) <= a xor b;
    layer0_outputs(8925) <= not (a xor b);
    layer0_outputs(8926) <= not (a or b);
    layer0_outputs(8927) <= not b;
    layer0_outputs(8928) <= not a;
    layer0_outputs(8929) <= a xor b;
    layer0_outputs(8930) <= a xor b;
    layer0_outputs(8931) <= b;
    layer0_outputs(8932) <= a or b;
    layer0_outputs(8933) <= not b or a;
    layer0_outputs(8934) <= not (a xor b);
    layer0_outputs(8935) <= a xor b;
    layer0_outputs(8936) <= '1';
    layer0_outputs(8937) <= not (a and b);
    layer0_outputs(8938) <= not (a and b);
    layer0_outputs(8939) <= not a;
    layer0_outputs(8940) <= not a;
    layer0_outputs(8941) <= b;
    layer0_outputs(8942) <= a;
    layer0_outputs(8943) <= not b;
    layer0_outputs(8944) <= a or b;
    layer0_outputs(8945) <= not b or a;
    layer0_outputs(8946) <= not b;
    layer0_outputs(8947) <= a or b;
    layer0_outputs(8948) <= not a or b;
    layer0_outputs(8949) <= not a;
    layer0_outputs(8950) <= not a;
    layer0_outputs(8951) <= a;
    layer0_outputs(8952) <= not a or b;
    layer0_outputs(8953) <= not b;
    layer0_outputs(8954) <= a or b;
    layer0_outputs(8955) <= not (a or b);
    layer0_outputs(8956) <= a and not b;
    layer0_outputs(8957) <= b and not a;
    layer0_outputs(8958) <= not b;
    layer0_outputs(8959) <= not b;
    layer0_outputs(8960) <= not (a or b);
    layer0_outputs(8961) <= not (a or b);
    layer0_outputs(8962) <= not (a or b);
    layer0_outputs(8963) <= not (a or b);
    layer0_outputs(8964) <= a and not b;
    layer0_outputs(8965) <= a or b;
    layer0_outputs(8966) <= b;
    layer0_outputs(8967) <= not (a xor b);
    layer0_outputs(8968) <= a xor b;
    layer0_outputs(8969) <= a and b;
    layer0_outputs(8970) <= not b or a;
    layer0_outputs(8971) <= a and not b;
    layer0_outputs(8972) <= a or b;
    layer0_outputs(8973) <= not (a xor b);
    layer0_outputs(8974) <= not (a or b);
    layer0_outputs(8975) <= not a;
    layer0_outputs(8976) <= a and not b;
    layer0_outputs(8977) <= '1';
    layer0_outputs(8978) <= not (a xor b);
    layer0_outputs(8979) <= not b or a;
    layer0_outputs(8980) <= not (a and b);
    layer0_outputs(8981) <= not (a or b);
    layer0_outputs(8982) <= not (a xor b);
    layer0_outputs(8983) <= a and b;
    layer0_outputs(8984) <= b and not a;
    layer0_outputs(8985) <= a or b;
    layer0_outputs(8986) <= b;
    layer0_outputs(8987) <= not (a xor b);
    layer0_outputs(8988) <= '1';
    layer0_outputs(8989) <= b and not a;
    layer0_outputs(8990) <= a and b;
    layer0_outputs(8991) <= not a or b;
    layer0_outputs(8992) <= not (a or b);
    layer0_outputs(8993) <= not b or a;
    layer0_outputs(8994) <= not a;
    layer0_outputs(8995) <= not (a and b);
    layer0_outputs(8996) <= a;
    layer0_outputs(8997) <= b;
    layer0_outputs(8998) <= not b or a;
    layer0_outputs(8999) <= a;
    layer0_outputs(9000) <= b;
    layer0_outputs(9001) <= b;
    layer0_outputs(9002) <= '1';
    layer0_outputs(9003) <= not b or a;
    layer0_outputs(9004) <= not a;
    layer0_outputs(9005) <= not (a or b);
    layer0_outputs(9006) <= b;
    layer0_outputs(9007) <= a or b;
    layer0_outputs(9008) <= not b;
    layer0_outputs(9009) <= not a or b;
    layer0_outputs(9010) <= not (a or b);
    layer0_outputs(9011) <= not a or b;
    layer0_outputs(9012) <= b and not a;
    layer0_outputs(9013) <= a;
    layer0_outputs(9014) <= a or b;
    layer0_outputs(9015) <= not (a xor b);
    layer0_outputs(9016) <= a xor b;
    layer0_outputs(9017) <= a xor b;
    layer0_outputs(9018) <= a or b;
    layer0_outputs(9019) <= not (a or b);
    layer0_outputs(9020) <= a xor b;
    layer0_outputs(9021) <= a and not b;
    layer0_outputs(9022) <= not (a or b);
    layer0_outputs(9023) <= a or b;
    layer0_outputs(9024) <= '0';
    layer0_outputs(9025) <= a;
    layer0_outputs(9026) <= b and not a;
    layer0_outputs(9027) <= a;
    layer0_outputs(9028) <= not (a or b);
    layer0_outputs(9029) <= not (a or b);
    layer0_outputs(9030) <= not (a and b);
    layer0_outputs(9031) <= '0';
    layer0_outputs(9032) <= not b;
    layer0_outputs(9033) <= not b or a;
    layer0_outputs(9034) <= a and not b;
    layer0_outputs(9035) <= not (a or b);
    layer0_outputs(9036) <= a;
    layer0_outputs(9037) <= not (a or b);
    layer0_outputs(9038) <= a and not b;
    layer0_outputs(9039) <= not b;
    layer0_outputs(9040) <= a and not b;
    layer0_outputs(9041) <= not a or b;
    layer0_outputs(9042) <= '1';
    layer0_outputs(9043) <= not b;
    layer0_outputs(9044) <= '0';
    layer0_outputs(9045) <= not b or a;
    layer0_outputs(9046) <= a or b;
    layer0_outputs(9047) <= '0';
    layer0_outputs(9048) <= not a or b;
    layer0_outputs(9049) <= a and not b;
    layer0_outputs(9050) <= not (a xor b);
    layer0_outputs(9051) <= not (a xor b);
    layer0_outputs(9052) <= a and b;
    layer0_outputs(9053) <= a or b;
    layer0_outputs(9054) <= not b;
    layer0_outputs(9055) <= b and not a;
    layer0_outputs(9056) <= a xor b;
    layer0_outputs(9057) <= not (a or b);
    layer0_outputs(9058) <= a;
    layer0_outputs(9059) <= not (a or b);
    layer0_outputs(9060) <= a or b;
    layer0_outputs(9061) <= a xor b;
    layer0_outputs(9062) <= b;
    layer0_outputs(9063) <= b;
    layer0_outputs(9064) <= not (a and b);
    layer0_outputs(9065) <= not (a or b);
    layer0_outputs(9066) <= not (a xor b);
    layer0_outputs(9067) <= not b;
    layer0_outputs(9068) <= not (a xor b);
    layer0_outputs(9069) <= not b or a;
    layer0_outputs(9070) <= b;
    layer0_outputs(9071) <= b;
    layer0_outputs(9072) <= not b;
    layer0_outputs(9073) <= a or b;
    layer0_outputs(9074) <= a and not b;
    layer0_outputs(9075) <= not a or b;
    layer0_outputs(9076) <= a and not b;
    layer0_outputs(9077) <= a or b;
    layer0_outputs(9078) <= a;
    layer0_outputs(9079) <= '0';
    layer0_outputs(9080) <= '0';
    layer0_outputs(9081) <= a xor b;
    layer0_outputs(9082) <= not a or b;
    layer0_outputs(9083) <= not (a or b);
    layer0_outputs(9084) <= not a;
    layer0_outputs(9085) <= b;
    layer0_outputs(9086) <= '0';
    layer0_outputs(9087) <= a or b;
    layer0_outputs(9088) <= a and b;
    layer0_outputs(9089) <= '0';
    layer0_outputs(9090) <= a or b;
    layer0_outputs(9091) <= not (a or b);
    layer0_outputs(9092) <= not (a and b);
    layer0_outputs(9093) <= not b;
    layer0_outputs(9094) <= a and not b;
    layer0_outputs(9095) <= not b;
    layer0_outputs(9096) <= a or b;
    layer0_outputs(9097) <= b;
    layer0_outputs(9098) <= a or b;
    layer0_outputs(9099) <= not (a xor b);
    layer0_outputs(9100) <= a and b;
    layer0_outputs(9101) <= not b;
    layer0_outputs(9102) <= a xor b;
    layer0_outputs(9103) <= not b or a;
    layer0_outputs(9104) <= b;
    layer0_outputs(9105) <= b and not a;
    layer0_outputs(9106) <= '0';
    layer0_outputs(9107) <= a and not b;
    layer0_outputs(9108) <= not a;
    layer0_outputs(9109) <= a xor b;
    layer0_outputs(9110) <= a;
    layer0_outputs(9111) <= a or b;
    layer0_outputs(9112) <= not (a or b);
    layer0_outputs(9113) <= not (a or b);
    layer0_outputs(9114) <= a or b;
    layer0_outputs(9115) <= not b;
    layer0_outputs(9116) <= not (a xor b);
    layer0_outputs(9117) <= b and not a;
    layer0_outputs(9118) <= a;
    layer0_outputs(9119) <= not (a or b);
    layer0_outputs(9120) <= a or b;
    layer0_outputs(9121) <= not (a xor b);
    layer0_outputs(9122) <= not (a or b);
    layer0_outputs(9123) <= a or b;
    layer0_outputs(9124) <= b;
    layer0_outputs(9125) <= '0';
    layer0_outputs(9126) <= b;
    layer0_outputs(9127) <= not (a or b);
    layer0_outputs(9128) <= a and not b;
    layer0_outputs(9129) <= a or b;
    layer0_outputs(9130) <= '1';
    layer0_outputs(9131) <= not (a or b);
    layer0_outputs(9132) <= a and b;
    layer0_outputs(9133) <= b;
    layer0_outputs(9134) <= a xor b;
    layer0_outputs(9135) <= not a or b;
    layer0_outputs(9136) <= not (a and b);
    layer0_outputs(9137) <= b and not a;
    layer0_outputs(9138) <= b and not a;
    layer0_outputs(9139) <= not b;
    layer0_outputs(9140) <= a or b;
    layer0_outputs(9141) <= a and not b;
    layer0_outputs(9142) <= a and b;
    layer0_outputs(9143) <= b;
    layer0_outputs(9144) <= b and not a;
    layer0_outputs(9145) <= not (a or b);
    layer0_outputs(9146) <= not a or b;
    layer0_outputs(9147) <= not (a or b);
    layer0_outputs(9148) <= a or b;
    layer0_outputs(9149) <= a xor b;
    layer0_outputs(9150) <= not (a xor b);
    layer0_outputs(9151) <= b;
    layer0_outputs(9152) <= not a or b;
    layer0_outputs(9153) <= a or b;
    layer0_outputs(9154) <= not (a xor b);
    layer0_outputs(9155) <= '0';
    layer0_outputs(9156) <= b and not a;
    layer0_outputs(9157) <= not b;
    layer0_outputs(9158) <= a;
    layer0_outputs(9159) <= a;
    layer0_outputs(9160) <= a or b;
    layer0_outputs(9161) <= not b or a;
    layer0_outputs(9162) <= a and not b;
    layer0_outputs(9163) <= '0';
    layer0_outputs(9164) <= a xor b;
    layer0_outputs(9165) <= not a or b;
    layer0_outputs(9166) <= b and not a;
    layer0_outputs(9167) <= '1';
    layer0_outputs(9168) <= b and not a;
    layer0_outputs(9169) <= not b;
    layer0_outputs(9170) <= not (a xor b);
    layer0_outputs(9171) <= a;
    layer0_outputs(9172) <= b and not a;
    layer0_outputs(9173) <= a xor b;
    layer0_outputs(9174) <= '1';
    layer0_outputs(9175) <= not b;
    layer0_outputs(9176) <= not (a or b);
    layer0_outputs(9177) <= not b;
    layer0_outputs(9178) <= not b;
    layer0_outputs(9179) <= '1';
    layer0_outputs(9180) <= not a;
    layer0_outputs(9181) <= b and not a;
    layer0_outputs(9182) <= a or b;
    layer0_outputs(9183) <= a or b;
    layer0_outputs(9184) <= not a;
    layer0_outputs(9185) <= a or b;
    layer0_outputs(9186) <= a and b;
    layer0_outputs(9187) <= not (a or b);
    layer0_outputs(9188) <= '0';
    layer0_outputs(9189) <= not b or a;
    layer0_outputs(9190) <= not b;
    layer0_outputs(9191) <= not b;
    layer0_outputs(9192) <= a or b;
    layer0_outputs(9193) <= a or b;
    layer0_outputs(9194) <= a or b;
    layer0_outputs(9195) <= not (a and b);
    layer0_outputs(9196) <= b;
    layer0_outputs(9197) <= not (a or b);
    layer0_outputs(9198) <= not b or a;
    layer0_outputs(9199) <= a;
    layer0_outputs(9200) <= a or b;
    layer0_outputs(9201) <= b and not a;
    layer0_outputs(9202) <= not a;
    layer0_outputs(9203) <= not b or a;
    layer0_outputs(9204) <= not b;
    layer0_outputs(9205) <= not (a or b);
    layer0_outputs(9206) <= a or b;
    layer0_outputs(9207) <= a xor b;
    layer0_outputs(9208) <= not b;
    layer0_outputs(9209) <= b;
    layer0_outputs(9210) <= not (a xor b);
    layer0_outputs(9211) <= not (a or b);
    layer0_outputs(9212) <= a xor b;
    layer0_outputs(9213) <= not b;
    layer0_outputs(9214) <= not b or a;
    layer0_outputs(9215) <= b;
    layer0_outputs(9216) <= not a;
    layer0_outputs(9217) <= a or b;
    layer0_outputs(9218) <= not b or a;
    layer0_outputs(9219) <= a;
    layer0_outputs(9220) <= b;
    layer0_outputs(9221) <= not b;
    layer0_outputs(9222) <= b and not a;
    layer0_outputs(9223) <= a or b;
    layer0_outputs(9224) <= not (a or b);
    layer0_outputs(9225) <= b;
    layer0_outputs(9226) <= not a;
    layer0_outputs(9227) <= a and not b;
    layer0_outputs(9228) <= not (a xor b);
    layer0_outputs(9229) <= a and not b;
    layer0_outputs(9230) <= not (a or b);
    layer0_outputs(9231) <= not a;
    layer0_outputs(9232) <= '1';
    layer0_outputs(9233) <= a xor b;
    layer0_outputs(9234) <= not (a or b);
    layer0_outputs(9235) <= '1';
    layer0_outputs(9236) <= b and not a;
    layer0_outputs(9237) <= b and not a;
    layer0_outputs(9238) <= a or b;
    layer0_outputs(9239) <= not b or a;
    layer0_outputs(9240) <= a and not b;
    layer0_outputs(9241) <= not (a xor b);
    layer0_outputs(9242) <= b;
    layer0_outputs(9243) <= not a or b;
    layer0_outputs(9244) <= not b;
    layer0_outputs(9245) <= not (a or b);
    layer0_outputs(9246) <= not b;
    layer0_outputs(9247) <= not a or b;
    layer0_outputs(9248) <= a xor b;
    layer0_outputs(9249) <= b;
    layer0_outputs(9250) <= not b;
    layer0_outputs(9251) <= not (a xor b);
    layer0_outputs(9252) <= b and not a;
    layer0_outputs(9253) <= a and b;
    layer0_outputs(9254) <= b and not a;
    layer0_outputs(9255) <= not b or a;
    layer0_outputs(9256) <= not (a or b);
    layer0_outputs(9257) <= a;
    layer0_outputs(9258) <= a and not b;
    layer0_outputs(9259) <= a or b;
    layer0_outputs(9260) <= not b or a;
    layer0_outputs(9261) <= not (a or b);
    layer0_outputs(9262) <= '1';
    layer0_outputs(9263) <= not b or a;
    layer0_outputs(9264) <= a or b;
    layer0_outputs(9265) <= not a;
    layer0_outputs(9266) <= not (a or b);
    layer0_outputs(9267) <= a and not b;
    layer0_outputs(9268) <= a or b;
    layer0_outputs(9269) <= not (a xor b);
    layer0_outputs(9270) <= not (a or b);
    layer0_outputs(9271) <= a and not b;
    layer0_outputs(9272) <= b and not a;
    layer0_outputs(9273) <= not b;
    layer0_outputs(9274) <= a or b;
    layer0_outputs(9275) <= a or b;
    layer0_outputs(9276) <= b;
    layer0_outputs(9277) <= a xor b;
    layer0_outputs(9278) <= a;
    layer0_outputs(9279) <= not b or a;
    layer0_outputs(9280) <= not b;
    layer0_outputs(9281) <= a or b;
    layer0_outputs(9282) <= a;
    layer0_outputs(9283) <= not b or a;
    layer0_outputs(9284) <= b and not a;
    layer0_outputs(9285) <= not a or b;
    layer0_outputs(9286) <= not (a or b);
    layer0_outputs(9287) <= '1';
    layer0_outputs(9288) <= not (a or b);
    layer0_outputs(9289) <= b;
    layer0_outputs(9290) <= not b or a;
    layer0_outputs(9291) <= not (a and b);
    layer0_outputs(9292) <= a or b;
    layer0_outputs(9293) <= a or b;
    layer0_outputs(9294) <= not a or b;
    layer0_outputs(9295) <= b;
    layer0_outputs(9296) <= not b or a;
    layer0_outputs(9297) <= a or b;
    layer0_outputs(9298) <= b and not a;
    layer0_outputs(9299) <= not b;
    layer0_outputs(9300) <= not b or a;
    layer0_outputs(9301) <= a xor b;
    layer0_outputs(9302) <= a or b;
    layer0_outputs(9303) <= not b;
    layer0_outputs(9304) <= not b or a;
    layer0_outputs(9305) <= a or b;
    layer0_outputs(9306) <= not a or b;
    layer0_outputs(9307) <= '0';
    layer0_outputs(9308) <= not a or b;
    layer0_outputs(9309) <= a;
    layer0_outputs(9310) <= not a;
    layer0_outputs(9311) <= not (a xor b);
    layer0_outputs(9312) <= a;
    layer0_outputs(9313) <= a xor b;
    layer0_outputs(9314) <= a xor b;
    layer0_outputs(9315) <= a;
    layer0_outputs(9316) <= a xor b;
    layer0_outputs(9317) <= a xor b;
    layer0_outputs(9318) <= a and not b;
    layer0_outputs(9319) <= not b;
    layer0_outputs(9320) <= not (a xor b);
    layer0_outputs(9321) <= b;
    layer0_outputs(9322) <= not b or a;
    layer0_outputs(9323) <= a;
    layer0_outputs(9324) <= b and not a;
    layer0_outputs(9325) <= not (a or b);
    layer0_outputs(9326) <= '1';
    layer0_outputs(9327) <= a and b;
    layer0_outputs(9328) <= not a or b;
    layer0_outputs(9329) <= '1';
    layer0_outputs(9330) <= b;
    layer0_outputs(9331) <= not (a or b);
    layer0_outputs(9332) <= a and b;
    layer0_outputs(9333) <= a or b;
    layer0_outputs(9334) <= not a;
    layer0_outputs(9335) <= a or b;
    layer0_outputs(9336) <= '1';
    layer0_outputs(9337) <= not (a xor b);
    layer0_outputs(9338) <= not a or b;
    layer0_outputs(9339) <= not b or a;
    layer0_outputs(9340) <= a xor b;
    layer0_outputs(9341) <= a;
    layer0_outputs(9342) <= not b;
    layer0_outputs(9343) <= not b;
    layer0_outputs(9344) <= not b;
    layer0_outputs(9345) <= a xor b;
    layer0_outputs(9346) <= not b or a;
    layer0_outputs(9347) <= a;
    layer0_outputs(9348) <= not (a xor b);
    layer0_outputs(9349) <= not a or b;
    layer0_outputs(9350) <= a and not b;
    layer0_outputs(9351) <= not (a xor b);
    layer0_outputs(9352) <= not b or a;
    layer0_outputs(9353) <= a and b;
    layer0_outputs(9354) <= not (a or b);
    layer0_outputs(9355) <= a xor b;
    layer0_outputs(9356) <= b and not a;
    layer0_outputs(9357) <= not (a xor b);
    layer0_outputs(9358) <= not (a xor b);
    layer0_outputs(9359) <= not b;
    layer0_outputs(9360) <= not a;
    layer0_outputs(9361) <= not b;
    layer0_outputs(9362) <= a;
    layer0_outputs(9363) <= not (a xor b);
    layer0_outputs(9364) <= not (a or b);
    layer0_outputs(9365) <= not b;
    layer0_outputs(9366) <= a and not b;
    layer0_outputs(9367) <= not b;
    layer0_outputs(9368) <= not (a or b);
    layer0_outputs(9369) <= not a;
    layer0_outputs(9370) <= a;
    layer0_outputs(9371) <= not a;
    layer0_outputs(9372) <= not b or a;
    layer0_outputs(9373) <= a or b;
    layer0_outputs(9374) <= a and b;
    layer0_outputs(9375) <= not (a and b);
    layer0_outputs(9376) <= not a or b;
    layer0_outputs(9377) <= a;
    layer0_outputs(9378) <= a and b;
    layer0_outputs(9379) <= not (a or b);
    layer0_outputs(9380) <= a or b;
    layer0_outputs(9381) <= '1';
    layer0_outputs(9382) <= not b;
    layer0_outputs(9383) <= a and not b;
    layer0_outputs(9384) <= a and b;
    layer0_outputs(9385) <= a xor b;
    layer0_outputs(9386) <= b;
    layer0_outputs(9387) <= b and not a;
    layer0_outputs(9388) <= b;
    layer0_outputs(9389) <= a and b;
    layer0_outputs(9390) <= not a or b;
    layer0_outputs(9391) <= not a or b;
    layer0_outputs(9392) <= '0';
    layer0_outputs(9393) <= a xor b;
    layer0_outputs(9394) <= a and not b;
    layer0_outputs(9395) <= not (a or b);
    layer0_outputs(9396) <= not b;
    layer0_outputs(9397) <= a;
    layer0_outputs(9398) <= a xor b;
    layer0_outputs(9399) <= a or b;
    layer0_outputs(9400) <= not b;
    layer0_outputs(9401) <= not (a or b);
    layer0_outputs(9402) <= not (a xor b);
    layer0_outputs(9403) <= not a;
    layer0_outputs(9404) <= a;
    layer0_outputs(9405) <= a;
    layer0_outputs(9406) <= a or b;
    layer0_outputs(9407) <= '1';
    layer0_outputs(9408) <= a or b;
    layer0_outputs(9409) <= not a;
    layer0_outputs(9410) <= b;
    layer0_outputs(9411) <= not a or b;
    layer0_outputs(9412) <= not a;
    layer0_outputs(9413) <= not (a or b);
    layer0_outputs(9414) <= a xor b;
    layer0_outputs(9415) <= not (a or b);
    layer0_outputs(9416) <= b;
    layer0_outputs(9417) <= not b or a;
    layer0_outputs(9418) <= a;
    layer0_outputs(9419) <= a xor b;
    layer0_outputs(9420) <= b and not a;
    layer0_outputs(9421) <= not a or b;
    layer0_outputs(9422) <= b;
    layer0_outputs(9423) <= b;
    layer0_outputs(9424) <= not b or a;
    layer0_outputs(9425) <= not (a or b);
    layer0_outputs(9426) <= not a or b;
    layer0_outputs(9427) <= b;
    layer0_outputs(9428) <= '0';
    layer0_outputs(9429) <= not (a and b);
    layer0_outputs(9430) <= b;
    layer0_outputs(9431) <= a or b;
    layer0_outputs(9432) <= a or b;
    layer0_outputs(9433) <= not (a or b);
    layer0_outputs(9434) <= a and b;
    layer0_outputs(9435) <= not (a or b);
    layer0_outputs(9436) <= not (a or b);
    layer0_outputs(9437) <= not a;
    layer0_outputs(9438) <= not (a or b);
    layer0_outputs(9439) <= not b or a;
    layer0_outputs(9440) <= b and not a;
    layer0_outputs(9441) <= a or b;
    layer0_outputs(9442) <= a;
    layer0_outputs(9443) <= not b;
    layer0_outputs(9444) <= b and not a;
    layer0_outputs(9445) <= a or b;
    layer0_outputs(9446) <= not (a or b);
    layer0_outputs(9447) <= not (a xor b);
    layer0_outputs(9448) <= not b or a;
    layer0_outputs(9449) <= not a;
    layer0_outputs(9450) <= a;
    layer0_outputs(9451) <= a and not b;
    layer0_outputs(9452) <= not (a xor b);
    layer0_outputs(9453) <= a and not b;
    layer0_outputs(9454) <= not b;
    layer0_outputs(9455) <= not b or a;
    layer0_outputs(9456) <= not (a and b);
    layer0_outputs(9457) <= not b;
    layer0_outputs(9458) <= '1';
    layer0_outputs(9459) <= a and b;
    layer0_outputs(9460) <= not (a xor b);
    layer0_outputs(9461) <= a and not b;
    layer0_outputs(9462) <= '0';
    layer0_outputs(9463) <= a and not b;
    layer0_outputs(9464) <= not b;
    layer0_outputs(9465) <= not a;
    layer0_outputs(9466) <= a xor b;
    layer0_outputs(9467) <= not b;
    layer0_outputs(9468) <= not b;
    layer0_outputs(9469) <= b;
    layer0_outputs(9470) <= a and not b;
    layer0_outputs(9471) <= a or b;
    layer0_outputs(9472) <= b and not a;
    layer0_outputs(9473) <= not (a xor b);
    layer0_outputs(9474) <= a xor b;
    layer0_outputs(9475) <= b and not a;
    layer0_outputs(9476) <= not b;
    layer0_outputs(9477) <= b;
    layer0_outputs(9478) <= not b;
    layer0_outputs(9479) <= b and not a;
    layer0_outputs(9480) <= b;
    layer0_outputs(9481) <= not (a xor b);
    layer0_outputs(9482) <= not a or b;
    layer0_outputs(9483) <= not (a xor b);
    layer0_outputs(9484) <= b and not a;
    layer0_outputs(9485) <= not b or a;
    layer0_outputs(9486) <= not (a or b);
    layer0_outputs(9487) <= a or b;
    layer0_outputs(9488) <= not (a or b);
    layer0_outputs(9489) <= not b;
    layer0_outputs(9490) <= a or b;
    layer0_outputs(9491) <= a or b;
    layer0_outputs(9492) <= not b or a;
    layer0_outputs(9493) <= b;
    layer0_outputs(9494) <= '0';
    layer0_outputs(9495) <= not a or b;
    layer0_outputs(9496) <= b;
    layer0_outputs(9497) <= not b or a;
    layer0_outputs(9498) <= not a or b;
    layer0_outputs(9499) <= not a or b;
    layer0_outputs(9500) <= not a or b;
    layer0_outputs(9501) <= b;
    layer0_outputs(9502) <= b;
    layer0_outputs(9503) <= not (a xor b);
    layer0_outputs(9504) <= a xor b;
    layer0_outputs(9505) <= not (a xor b);
    layer0_outputs(9506) <= not (a or b);
    layer0_outputs(9507) <= a xor b;
    layer0_outputs(9508) <= not (a or b);
    layer0_outputs(9509) <= not (a or b);
    layer0_outputs(9510) <= a and not b;
    layer0_outputs(9511) <= not a or b;
    layer0_outputs(9512) <= not (a xor b);
    layer0_outputs(9513) <= not a or b;
    layer0_outputs(9514) <= a xor b;
    layer0_outputs(9515) <= a or b;
    layer0_outputs(9516) <= not (a xor b);
    layer0_outputs(9517) <= not (a and b);
    layer0_outputs(9518) <= a and b;
    layer0_outputs(9519) <= a;
    layer0_outputs(9520) <= '1';
    layer0_outputs(9521) <= not b;
    layer0_outputs(9522) <= a and b;
    layer0_outputs(9523) <= not b or a;
    layer0_outputs(9524) <= b and not a;
    layer0_outputs(9525) <= b and not a;
    layer0_outputs(9526) <= '0';
    layer0_outputs(9527) <= a xor b;
    layer0_outputs(9528) <= a and not b;
    layer0_outputs(9529) <= b;
    layer0_outputs(9530) <= not a;
    layer0_outputs(9531) <= not (a xor b);
    layer0_outputs(9532) <= a and not b;
    layer0_outputs(9533) <= not a or b;
    layer0_outputs(9534) <= not b;
    layer0_outputs(9535) <= not b;
    layer0_outputs(9536) <= a or b;
    layer0_outputs(9537) <= a or b;
    layer0_outputs(9538) <= a and not b;
    layer0_outputs(9539) <= a or b;
    layer0_outputs(9540) <= not b;
    layer0_outputs(9541) <= not a;
    layer0_outputs(9542) <= b and not a;
    layer0_outputs(9543) <= a and b;
    layer0_outputs(9544) <= b;
    layer0_outputs(9545) <= not b;
    layer0_outputs(9546) <= not a or b;
    layer0_outputs(9547) <= not a;
    layer0_outputs(9548) <= not (a or b);
    layer0_outputs(9549) <= '1';
    layer0_outputs(9550) <= not (a or b);
    layer0_outputs(9551) <= a xor b;
    layer0_outputs(9552) <= not (a xor b);
    layer0_outputs(9553) <= a or b;
    layer0_outputs(9554) <= a or b;
    layer0_outputs(9555) <= a or b;
    layer0_outputs(9556) <= b and not a;
    layer0_outputs(9557) <= b and not a;
    layer0_outputs(9558) <= not (a or b);
    layer0_outputs(9559) <= not a;
    layer0_outputs(9560) <= not (a xor b);
    layer0_outputs(9561) <= not (a and b);
    layer0_outputs(9562) <= a;
    layer0_outputs(9563) <= not b;
    layer0_outputs(9564) <= not (a xor b);
    layer0_outputs(9565) <= not (a or b);
    layer0_outputs(9566) <= a or b;
    layer0_outputs(9567) <= not a or b;
    layer0_outputs(9568) <= b and not a;
    layer0_outputs(9569) <= b and not a;
    layer0_outputs(9570) <= not b;
    layer0_outputs(9571) <= not (a xor b);
    layer0_outputs(9572) <= not (a or b);
    layer0_outputs(9573) <= a xor b;
    layer0_outputs(9574) <= a and not b;
    layer0_outputs(9575) <= '0';
    layer0_outputs(9576) <= a xor b;
    layer0_outputs(9577) <= not b or a;
    layer0_outputs(9578) <= '1';
    layer0_outputs(9579) <= a;
    layer0_outputs(9580) <= a;
    layer0_outputs(9581) <= not (a or b);
    layer0_outputs(9582) <= not (a or b);
    layer0_outputs(9583) <= b;
    layer0_outputs(9584) <= a or b;
    layer0_outputs(9585) <= a xor b;
    layer0_outputs(9586) <= '0';
    layer0_outputs(9587) <= a;
    layer0_outputs(9588) <= not (a or b);
    layer0_outputs(9589) <= a and not b;
    layer0_outputs(9590) <= a and not b;
    layer0_outputs(9591) <= not (a and b);
    layer0_outputs(9592) <= not (a and b);
    layer0_outputs(9593) <= not (a or b);
    layer0_outputs(9594) <= not (a or b);
    layer0_outputs(9595) <= b;
    layer0_outputs(9596) <= not a;
    layer0_outputs(9597) <= not b or a;
    layer0_outputs(9598) <= a or b;
    layer0_outputs(9599) <= not b;
    layer0_outputs(9600) <= a xor b;
    layer0_outputs(9601) <= a and not b;
    layer0_outputs(9602) <= not (a xor b);
    layer0_outputs(9603) <= b;
    layer0_outputs(9604) <= not b or a;
    layer0_outputs(9605) <= a and not b;
    layer0_outputs(9606) <= a;
    layer0_outputs(9607) <= not a or b;
    layer0_outputs(9608) <= not b;
    layer0_outputs(9609) <= not b or a;
    layer0_outputs(9610) <= not b or a;
    layer0_outputs(9611) <= a or b;
    layer0_outputs(9612) <= not a;
    layer0_outputs(9613) <= a;
    layer0_outputs(9614) <= not (a or b);
    layer0_outputs(9615) <= a or b;
    layer0_outputs(9616) <= not (a or b);
    layer0_outputs(9617) <= a or b;
    layer0_outputs(9618) <= not (a xor b);
    layer0_outputs(9619) <= not a;
    layer0_outputs(9620) <= not a or b;
    layer0_outputs(9621) <= b;
    layer0_outputs(9622) <= not a or b;
    layer0_outputs(9623) <= a or b;
    layer0_outputs(9624) <= not b or a;
    layer0_outputs(9625) <= not (a xor b);
    layer0_outputs(9626) <= a and not b;
    layer0_outputs(9627) <= a xor b;
    layer0_outputs(9628) <= a and not b;
    layer0_outputs(9629) <= not (a xor b);
    layer0_outputs(9630) <= a and not b;
    layer0_outputs(9631) <= b;
    layer0_outputs(9632) <= a and not b;
    layer0_outputs(9633) <= not (a or b);
    layer0_outputs(9634) <= not a or b;
    layer0_outputs(9635) <= '1';
    layer0_outputs(9636) <= not (a or b);
    layer0_outputs(9637) <= not b;
    layer0_outputs(9638) <= not b;
    layer0_outputs(9639) <= a or b;
    layer0_outputs(9640) <= a;
    layer0_outputs(9641) <= not a;
    layer0_outputs(9642) <= a or b;
    layer0_outputs(9643) <= not (a xor b);
    layer0_outputs(9644) <= not a or b;
    layer0_outputs(9645) <= a;
    layer0_outputs(9646) <= a or b;
    layer0_outputs(9647) <= a xor b;
    layer0_outputs(9648) <= a;
    layer0_outputs(9649) <= a and b;
    layer0_outputs(9650) <= a or b;
    layer0_outputs(9651) <= '1';
    layer0_outputs(9652) <= not a or b;
    layer0_outputs(9653) <= not (a or b);
    layer0_outputs(9654) <= a;
    layer0_outputs(9655) <= b;
    layer0_outputs(9656) <= not a or b;
    layer0_outputs(9657) <= not b or a;
    layer0_outputs(9658) <= not (a or b);
    layer0_outputs(9659) <= b and not a;
    layer0_outputs(9660) <= a and not b;
    layer0_outputs(9661) <= a or b;
    layer0_outputs(9662) <= a xor b;
    layer0_outputs(9663) <= not (a or b);
    layer0_outputs(9664) <= a or b;
    layer0_outputs(9665) <= not a or b;
    layer0_outputs(9666) <= a or b;
    layer0_outputs(9667) <= a xor b;
    layer0_outputs(9668) <= a and not b;
    layer0_outputs(9669) <= '1';
    layer0_outputs(9670) <= a or b;
    layer0_outputs(9671) <= '1';
    layer0_outputs(9672) <= a and not b;
    layer0_outputs(9673) <= a xor b;
    layer0_outputs(9674) <= b;
    layer0_outputs(9675) <= a or b;
    layer0_outputs(9676) <= not a or b;
    layer0_outputs(9677) <= b and not a;
    layer0_outputs(9678) <= b;
    layer0_outputs(9679) <= a and not b;
    layer0_outputs(9680) <= a or b;
    layer0_outputs(9681) <= not (a or b);
    layer0_outputs(9682) <= not b or a;
    layer0_outputs(9683) <= a xor b;
    layer0_outputs(9684) <= a or b;
    layer0_outputs(9685) <= a xor b;
    layer0_outputs(9686) <= not (a or b);
    layer0_outputs(9687) <= '1';
    layer0_outputs(9688) <= a xor b;
    layer0_outputs(9689) <= not (a or b);
    layer0_outputs(9690) <= not b;
    layer0_outputs(9691) <= a and not b;
    layer0_outputs(9692) <= not (a xor b);
    layer0_outputs(9693) <= not (a or b);
    layer0_outputs(9694) <= not b or a;
    layer0_outputs(9695) <= not b;
    layer0_outputs(9696) <= b;
    layer0_outputs(9697) <= a and not b;
    layer0_outputs(9698) <= not b or a;
    layer0_outputs(9699) <= b;
    layer0_outputs(9700) <= not a;
    layer0_outputs(9701) <= not a or b;
    layer0_outputs(9702) <= not (a or b);
    layer0_outputs(9703) <= b;
    layer0_outputs(9704) <= a and not b;
    layer0_outputs(9705) <= b and not a;
    layer0_outputs(9706) <= a;
    layer0_outputs(9707) <= a xor b;
    layer0_outputs(9708) <= not (a and b);
    layer0_outputs(9709) <= a and not b;
    layer0_outputs(9710) <= a xor b;
    layer0_outputs(9711) <= not (a or b);
    layer0_outputs(9712) <= a xor b;
    layer0_outputs(9713) <= not (a or b);
    layer0_outputs(9714) <= b;
    layer0_outputs(9715) <= not (a xor b);
    layer0_outputs(9716) <= a xor b;
    layer0_outputs(9717) <= a xor b;
    layer0_outputs(9718) <= not (a or b);
    layer0_outputs(9719) <= not (a or b);
    layer0_outputs(9720) <= a xor b;
    layer0_outputs(9721) <= a;
    layer0_outputs(9722) <= b and not a;
    layer0_outputs(9723) <= not a;
    layer0_outputs(9724) <= not b;
    layer0_outputs(9725) <= a and not b;
    layer0_outputs(9726) <= not b;
    layer0_outputs(9727) <= a;
    layer0_outputs(9728) <= not (a xor b);
    layer0_outputs(9729) <= not (a xor b);
    layer0_outputs(9730) <= b;
    layer0_outputs(9731) <= not (a xor b);
    layer0_outputs(9732) <= not (a and b);
    layer0_outputs(9733) <= b;
    layer0_outputs(9734) <= a or b;
    layer0_outputs(9735) <= b;
    layer0_outputs(9736) <= not (a or b);
    layer0_outputs(9737) <= not (a or b);
    layer0_outputs(9738) <= not a;
    layer0_outputs(9739) <= '1';
    layer0_outputs(9740) <= not (a xor b);
    layer0_outputs(9741) <= not a;
    layer0_outputs(9742) <= a;
    layer0_outputs(9743) <= a and b;
    layer0_outputs(9744) <= not b;
    layer0_outputs(9745) <= a or b;
    layer0_outputs(9746) <= not (a xor b);
    layer0_outputs(9747) <= a;
    layer0_outputs(9748) <= b and not a;
    layer0_outputs(9749) <= a;
    layer0_outputs(9750) <= a or b;
    layer0_outputs(9751) <= a or b;
    layer0_outputs(9752) <= a;
    layer0_outputs(9753) <= a;
    layer0_outputs(9754) <= not b or a;
    layer0_outputs(9755) <= not b;
    layer0_outputs(9756) <= a or b;
    layer0_outputs(9757) <= a or b;
    layer0_outputs(9758) <= not (a xor b);
    layer0_outputs(9759) <= not a or b;
    layer0_outputs(9760) <= a or b;
    layer0_outputs(9761) <= a or b;
    layer0_outputs(9762) <= not a or b;
    layer0_outputs(9763) <= a and b;
    layer0_outputs(9764) <= not (a or b);
    layer0_outputs(9765) <= b;
    layer0_outputs(9766) <= b and not a;
    layer0_outputs(9767) <= b;
    layer0_outputs(9768) <= a or b;
    layer0_outputs(9769) <= not b or a;
    layer0_outputs(9770) <= a;
    layer0_outputs(9771) <= not b or a;
    layer0_outputs(9772) <= '0';
    layer0_outputs(9773) <= b and not a;
    layer0_outputs(9774) <= a or b;
    layer0_outputs(9775) <= not b or a;
    layer0_outputs(9776) <= a or b;
    layer0_outputs(9777) <= a xor b;
    layer0_outputs(9778) <= a xor b;
    layer0_outputs(9779) <= a and not b;
    layer0_outputs(9780) <= not (a or b);
    layer0_outputs(9781) <= not b or a;
    layer0_outputs(9782) <= not (a or b);
    layer0_outputs(9783) <= not a;
    layer0_outputs(9784) <= a;
    layer0_outputs(9785) <= not (a or b);
    layer0_outputs(9786) <= a or b;
    layer0_outputs(9787) <= a;
    layer0_outputs(9788) <= a;
    layer0_outputs(9789) <= a or b;
    layer0_outputs(9790) <= a or b;
    layer0_outputs(9791) <= b;
    layer0_outputs(9792) <= not (a or b);
    layer0_outputs(9793) <= a or b;
    layer0_outputs(9794) <= not (a or b);
    layer0_outputs(9795) <= not a or b;
    layer0_outputs(9796) <= a;
    layer0_outputs(9797) <= a or b;
    layer0_outputs(9798) <= a and b;
    layer0_outputs(9799) <= a xor b;
    layer0_outputs(9800) <= not b or a;
    layer0_outputs(9801) <= not b;
    layer0_outputs(9802) <= not b or a;
    layer0_outputs(9803) <= a and not b;
    layer0_outputs(9804) <= a;
    layer0_outputs(9805) <= not a or b;
    layer0_outputs(9806) <= not (a xor b);
    layer0_outputs(9807) <= a or b;
    layer0_outputs(9808) <= a or b;
    layer0_outputs(9809) <= not (a xor b);
    layer0_outputs(9810) <= not a or b;
    layer0_outputs(9811) <= not a;
    layer0_outputs(9812) <= '1';
    layer0_outputs(9813) <= not (a or b);
    layer0_outputs(9814) <= a or b;
    layer0_outputs(9815) <= not b;
    layer0_outputs(9816) <= a or b;
    layer0_outputs(9817) <= not a;
    layer0_outputs(9818) <= not a or b;
    layer0_outputs(9819) <= not (a or b);
    layer0_outputs(9820) <= a or b;
    layer0_outputs(9821) <= a or b;
    layer0_outputs(9822) <= not b;
    layer0_outputs(9823) <= not b or a;
    layer0_outputs(9824) <= a xor b;
    layer0_outputs(9825) <= not b or a;
    layer0_outputs(9826) <= a or b;
    layer0_outputs(9827) <= '0';
    layer0_outputs(9828) <= not a or b;
    layer0_outputs(9829) <= a or b;
    layer0_outputs(9830) <= a and not b;
    layer0_outputs(9831) <= not b or a;
    layer0_outputs(9832) <= not a;
    layer0_outputs(9833) <= a xor b;
    layer0_outputs(9834) <= not b or a;
    layer0_outputs(9835) <= not (a and b);
    layer0_outputs(9836) <= b and not a;
    layer0_outputs(9837) <= not (a or b);
    layer0_outputs(9838) <= a or b;
    layer0_outputs(9839) <= a or b;
    layer0_outputs(9840) <= a or b;
    layer0_outputs(9841) <= not (a xor b);
    layer0_outputs(9842) <= a and not b;
    layer0_outputs(9843) <= not (a or b);
    layer0_outputs(9844) <= not (a or b);
    layer0_outputs(9845) <= not (a or b);
    layer0_outputs(9846) <= b and not a;
    layer0_outputs(9847) <= not (a or b);
    layer0_outputs(9848) <= not b;
    layer0_outputs(9849) <= '1';
    layer0_outputs(9850) <= not (a or b);
    layer0_outputs(9851) <= a or b;
    layer0_outputs(9852) <= not a;
    layer0_outputs(9853) <= not (a xor b);
    layer0_outputs(9854) <= a or b;
    layer0_outputs(9855) <= a xor b;
    layer0_outputs(9856) <= '0';
    layer0_outputs(9857) <= a;
    layer0_outputs(9858) <= a xor b;
    layer0_outputs(9859) <= a and b;
    layer0_outputs(9860) <= not b;
    layer0_outputs(9861) <= b and not a;
    layer0_outputs(9862) <= not (a or b);
    layer0_outputs(9863) <= b;
    layer0_outputs(9864) <= not b or a;
    layer0_outputs(9865) <= '0';
    layer0_outputs(9866) <= b and not a;
    layer0_outputs(9867) <= not (a or b);
    layer0_outputs(9868) <= a;
    layer0_outputs(9869) <= b;
    layer0_outputs(9870) <= not a;
    layer0_outputs(9871) <= a and not b;
    layer0_outputs(9872) <= a and b;
    layer0_outputs(9873) <= '1';
    layer0_outputs(9874) <= not (a xor b);
    layer0_outputs(9875) <= a or b;
    layer0_outputs(9876) <= a;
    layer0_outputs(9877) <= b and not a;
    layer0_outputs(9878) <= b and not a;
    layer0_outputs(9879) <= not a;
    layer0_outputs(9880) <= b;
    layer0_outputs(9881) <= a and b;
    layer0_outputs(9882) <= a and not b;
    layer0_outputs(9883) <= '1';
    layer0_outputs(9884) <= not a;
    layer0_outputs(9885) <= not (a xor b);
    layer0_outputs(9886) <= a or b;
    layer0_outputs(9887) <= not a or b;
    layer0_outputs(9888) <= b;
    layer0_outputs(9889) <= a or b;
    layer0_outputs(9890) <= not b;
    layer0_outputs(9891) <= a and not b;
    layer0_outputs(9892) <= a and b;
    layer0_outputs(9893) <= a xor b;
    layer0_outputs(9894) <= a or b;
    layer0_outputs(9895) <= not a;
    layer0_outputs(9896) <= not a;
    layer0_outputs(9897) <= a or b;
    layer0_outputs(9898) <= not b;
    layer0_outputs(9899) <= not (a xor b);
    layer0_outputs(9900) <= not (a or b);
    layer0_outputs(9901) <= not (a xor b);
    layer0_outputs(9902) <= a;
    layer0_outputs(9903) <= a;
    layer0_outputs(9904) <= a or b;
    layer0_outputs(9905) <= not (a or b);
    layer0_outputs(9906) <= a;
    layer0_outputs(9907) <= a and not b;
    layer0_outputs(9908) <= not a;
    layer0_outputs(9909) <= a;
    layer0_outputs(9910) <= not (a xor b);
    layer0_outputs(9911) <= a and not b;
    layer0_outputs(9912) <= not a;
    layer0_outputs(9913) <= a xor b;
    layer0_outputs(9914) <= a or b;
    layer0_outputs(9915) <= a xor b;
    layer0_outputs(9916) <= not (a or b);
    layer0_outputs(9917) <= b;
    layer0_outputs(9918) <= not a or b;
    layer0_outputs(9919) <= not b;
    layer0_outputs(9920) <= a;
    layer0_outputs(9921) <= not a or b;
    layer0_outputs(9922) <= a xor b;
    layer0_outputs(9923) <= not (a xor b);
    layer0_outputs(9924) <= a and b;
    layer0_outputs(9925) <= a or b;
    layer0_outputs(9926) <= not (a and b);
    layer0_outputs(9927) <= not a or b;
    layer0_outputs(9928) <= not (a or b);
    layer0_outputs(9929) <= a or b;
    layer0_outputs(9930) <= a;
    layer0_outputs(9931) <= not a or b;
    layer0_outputs(9932) <= a xor b;
    layer0_outputs(9933) <= not (a or b);
    layer0_outputs(9934) <= not b;
    layer0_outputs(9935) <= not (a xor b);
    layer0_outputs(9936) <= not a;
    layer0_outputs(9937) <= not b;
    layer0_outputs(9938) <= not b;
    layer0_outputs(9939) <= a;
    layer0_outputs(9940) <= not a;
    layer0_outputs(9941) <= not b or a;
    layer0_outputs(9942) <= not a or b;
    layer0_outputs(9943) <= a;
    layer0_outputs(9944) <= a;
    layer0_outputs(9945) <= a or b;
    layer0_outputs(9946) <= not a or b;
    layer0_outputs(9947) <= a or b;
    layer0_outputs(9948) <= a xor b;
    layer0_outputs(9949) <= not (a xor b);
    layer0_outputs(9950) <= not (a or b);
    layer0_outputs(9951) <= b;
    layer0_outputs(9952) <= not (a xor b);
    layer0_outputs(9953) <= not b or a;
    layer0_outputs(9954) <= b;
    layer0_outputs(9955) <= a;
    layer0_outputs(9956) <= a or b;
    layer0_outputs(9957) <= not (a and b);
    layer0_outputs(9958) <= a and b;
    layer0_outputs(9959) <= not b;
    layer0_outputs(9960) <= not (a xor b);
    layer0_outputs(9961) <= not (a xor b);
    layer0_outputs(9962) <= a and b;
    layer0_outputs(9963) <= a xor b;
    layer0_outputs(9964) <= a or b;
    layer0_outputs(9965) <= a or b;
    layer0_outputs(9966) <= not b or a;
    layer0_outputs(9967) <= not (a or b);
    layer0_outputs(9968) <= a;
    layer0_outputs(9969) <= a xor b;
    layer0_outputs(9970) <= not b or a;
    layer0_outputs(9971) <= not a or b;
    layer0_outputs(9972) <= not (a or b);
    layer0_outputs(9973) <= not (a or b);
    layer0_outputs(9974) <= a or b;
    layer0_outputs(9975) <= b;
    layer0_outputs(9976) <= not b or a;
    layer0_outputs(9977) <= not (a or b);
    layer0_outputs(9978) <= not (a xor b);
    layer0_outputs(9979) <= not (a or b);
    layer0_outputs(9980) <= b;
    layer0_outputs(9981) <= not a;
    layer0_outputs(9982) <= not a or b;
    layer0_outputs(9983) <= a xor b;
    layer0_outputs(9984) <= b and not a;
    layer0_outputs(9985) <= not a;
    layer0_outputs(9986) <= not a;
    layer0_outputs(9987) <= not a or b;
    layer0_outputs(9988) <= b;
    layer0_outputs(9989) <= not a or b;
    layer0_outputs(9990) <= not (a xor b);
    layer0_outputs(9991) <= a and b;
    layer0_outputs(9992) <= not a or b;
    layer0_outputs(9993) <= not b or a;
    layer0_outputs(9994) <= a;
    layer0_outputs(9995) <= b;
    layer0_outputs(9996) <= not (a xor b);
    layer0_outputs(9997) <= b and not a;
    layer0_outputs(9998) <= a;
    layer0_outputs(9999) <= a and not b;
    layer0_outputs(10000) <= not (a and b);
    layer0_outputs(10001) <= a or b;
    layer0_outputs(10002) <= '0';
    layer0_outputs(10003) <= '1';
    layer0_outputs(10004) <= not a;
    layer0_outputs(10005) <= not b;
    layer0_outputs(10006) <= not a;
    layer0_outputs(10007) <= b;
    layer0_outputs(10008) <= not (a xor b);
    layer0_outputs(10009) <= a;
    layer0_outputs(10010) <= a or b;
    layer0_outputs(10011) <= not a or b;
    layer0_outputs(10012) <= a and b;
    layer0_outputs(10013) <= b and not a;
    layer0_outputs(10014) <= a xor b;
    layer0_outputs(10015) <= not (a or b);
    layer0_outputs(10016) <= not (a xor b);
    layer0_outputs(10017) <= not b or a;
    layer0_outputs(10018) <= not a;
    layer0_outputs(10019) <= b;
    layer0_outputs(10020) <= a;
    layer0_outputs(10021) <= not (a or b);
    layer0_outputs(10022) <= a or b;
    layer0_outputs(10023) <= a xor b;
    layer0_outputs(10024) <= a and not b;
    layer0_outputs(10025) <= a or b;
    layer0_outputs(10026) <= not (a xor b);
    layer0_outputs(10027) <= not (a or b);
    layer0_outputs(10028) <= a or b;
    layer0_outputs(10029) <= b;
    layer0_outputs(10030) <= not a or b;
    layer0_outputs(10031) <= not (a and b);
    layer0_outputs(10032) <= a xor b;
    layer0_outputs(10033) <= not (a xor b);
    layer0_outputs(10034) <= not a;
    layer0_outputs(10035) <= a and b;
    layer0_outputs(10036) <= not b or a;
    layer0_outputs(10037) <= not a;
    layer0_outputs(10038) <= a and not b;
    layer0_outputs(10039) <= not b or a;
    layer0_outputs(10040) <= a;
    layer0_outputs(10041) <= a and b;
    layer0_outputs(10042) <= '0';
    layer0_outputs(10043) <= not a or b;
    layer0_outputs(10044) <= not (a or b);
    layer0_outputs(10045) <= a xor b;
    layer0_outputs(10046) <= b;
    layer0_outputs(10047) <= b;
    layer0_outputs(10048) <= '1';
    layer0_outputs(10049) <= a;
    layer0_outputs(10050) <= not a;
    layer0_outputs(10051) <= not (a xor b);
    layer0_outputs(10052) <= a xor b;
    layer0_outputs(10053) <= a xor b;
    layer0_outputs(10054) <= not b or a;
    layer0_outputs(10055) <= not b;
    layer0_outputs(10056) <= a xor b;
    layer0_outputs(10057) <= a or b;
    layer0_outputs(10058) <= not (a or b);
    layer0_outputs(10059) <= a or b;
    layer0_outputs(10060) <= a;
    layer0_outputs(10061) <= not b;
    layer0_outputs(10062) <= not (a or b);
    layer0_outputs(10063) <= a;
    layer0_outputs(10064) <= '1';
    layer0_outputs(10065) <= a or b;
    layer0_outputs(10066) <= not (a xor b);
    layer0_outputs(10067) <= not (a or b);
    layer0_outputs(10068) <= a or b;
    layer0_outputs(10069) <= a;
    layer0_outputs(10070) <= b and not a;
    layer0_outputs(10071) <= not (a xor b);
    layer0_outputs(10072) <= a or b;
    layer0_outputs(10073) <= a and not b;
    layer0_outputs(10074) <= a or b;
    layer0_outputs(10075) <= '0';
    layer0_outputs(10076) <= not a or b;
    layer0_outputs(10077) <= not b or a;
    layer0_outputs(10078) <= a;
    layer0_outputs(10079) <= not (a and b);
    layer0_outputs(10080) <= a and not b;
    layer0_outputs(10081) <= not (a or b);
    layer0_outputs(10082) <= not b;
    layer0_outputs(10083) <= not b;
    layer0_outputs(10084) <= not (a xor b);
    layer0_outputs(10085) <= b;
    layer0_outputs(10086) <= a xor b;
    layer0_outputs(10087) <= not b or a;
    layer0_outputs(10088) <= not b;
    layer0_outputs(10089) <= not (a and b);
    layer0_outputs(10090) <= not a;
    layer0_outputs(10091) <= not (a or b);
    layer0_outputs(10092) <= not (a xor b);
    layer0_outputs(10093) <= a or b;
    layer0_outputs(10094) <= a;
    layer0_outputs(10095) <= a;
    layer0_outputs(10096) <= not a or b;
    layer0_outputs(10097) <= a;
    layer0_outputs(10098) <= b and not a;
    layer0_outputs(10099) <= not (a or b);
    layer0_outputs(10100) <= b;
    layer0_outputs(10101) <= b and not a;
    layer0_outputs(10102) <= not b;
    layer0_outputs(10103) <= a and not b;
    layer0_outputs(10104) <= b and not a;
    layer0_outputs(10105) <= a;
    layer0_outputs(10106) <= b;
    layer0_outputs(10107) <= '1';
    layer0_outputs(10108) <= not a;
    layer0_outputs(10109) <= not b;
    layer0_outputs(10110) <= a and b;
    layer0_outputs(10111) <= a or b;
    layer0_outputs(10112) <= a or b;
    layer0_outputs(10113) <= not b;
    layer0_outputs(10114) <= a or b;
    layer0_outputs(10115) <= a and not b;
    layer0_outputs(10116) <= not (a and b);
    layer0_outputs(10117) <= not b;
    layer0_outputs(10118) <= a and not b;
    layer0_outputs(10119) <= a;
    layer0_outputs(10120) <= a and not b;
    layer0_outputs(10121) <= a and not b;
    layer0_outputs(10122) <= '0';
    layer0_outputs(10123) <= a;
    layer0_outputs(10124) <= a or b;
    layer0_outputs(10125) <= b and not a;
    layer0_outputs(10126) <= b;
    layer0_outputs(10127) <= a xor b;
    layer0_outputs(10128) <= '1';
    layer0_outputs(10129) <= not a;
    layer0_outputs(10130) <= a or b;
    layer0_outputs(10131) <= a or b;
    layer0_outputs(10132) <= a;
    layer0_outputs(10133) <= '0';
    layer0_outputs(10134) <= a and not b;
    layer0_outputs(10135) <= not b or a;
    layer0_outputs(10136) <= not (a or b);
    layer0_outputs(10137) <= a and not b;
    layer0_outputs(10138) <= not b or a;
    layer0_outputs(10139) <= not (a xor b);
    layer0_outputs(10140) <= b;
    layer0_outputs(10141) <= not (a xor b);
    layer0_outputs(10142) <= a or b;
    layer0_outputs(10143) <= a and not b;
    layer0_outputs(10144) <= a or b;
    layer0_outputs(10145) <= not (a or b);
    layer0_outputs(10146) <= not (a xor b);
    layer0_outputs(10147) <= a and not b;
    layer0_outputs(10148) <= not (a or b);
    layer0_outputs(10149) <= a xor b;
    layer0_outputs(10150) <= a;
    layer0_outputs(10151) <= not (a or b);
    layer0_outputs(10152) <= b;
    layer0_outputs(10153) <= b;
    layer0_outputs(10154) <= b;
    layer0_outputs(10155) <= not a;
    layer0_outputs(10156) <= a;
    layer0_outputs(10157) <= not a;
    layer0_outputs(10158) <= a xor b;
    layer0_outputs(10159) <= not (a or b);
    layer0_outputs(10160) <= not a;
    layer0_outputs(10161) <= '0';
    layer0_outputs(10162) <= not (a xor b);
    layer0_outputs(10163) <= a and not b;
    layer0_outputs(10164) <= a or b;
    layer0_outputs(10165) <= not (a or b);
    layer0_outputs(10166) <= not a;
    layer0_outputs(10167) <= a;
    layer0_outputs(10168) <= a xor b;
    layer0_outputs(10169) <= not (a xor b);
    layer0_outputs(10170) <= not b or a;
    layer0_outputs(10171) <= not (a xor b);
    layer0_outputs(10172) <= not (a or b);
    layer0_outputs(10173) <= b;
    layer0_outputs(10174) <= a or b;
    layer0_outputs(10175) <= not (a xor b);
    layer0_outputs(10176) <= not a or b;
    layer0_outputs(10177) <= b;
    layer0_outputs(10178) <= not a;
    layer0_outputs(10179) <= a and not b;
    layer0_outputs(10180) <= not a;
    layer0_outputs(10181) <= a xor b;
    layer0_outputs(10182) <= not (a or b);
    layer0_outputs(10183) <= b and not a;
    layer0_outputs(10184) <= a and not b;
    layer0_outputs(10185) <= a;
    layer0_outputs(10186) <= not b;
    layer0_outputs(10187) <= not (a or b);
    layer0_outputs(10188) <= a and not b;
    layer0_outputs(10189) <= '0';
    layer0_outputs(10190) <= a or b;
    layer0_outputs(10191) <= a xor b;
    layer0_outputs(10192) <= b and not a;
    layer0_outputs(10193) <= b and not a;
    layer0_outputs(10194) <= not a or b;
    layer0_outputs(10195) <= not (a or b);
    layer0_outputs(10196) <= not a;
    layer0_outputs(10197) <= b;
    layer0_outputs(10198) <= a and b;
    layer0_outputs(10199) <= a and b;
    layer0_outputs(10200) <= not (a xor b);
    layer0_outputs(10201) <= '0';
    layer0_outputs(10202) <= not (a or b);
    layer0_outputs(10203) <= not b;
    layer0_outputs(10204) <= not (a or b);
    layer0_outputs(10205) <= b and not a;
    layer0_outputs(10206) <= not b or a;
    layer0_outputs(10207) <= not a or b;
    layer0_outputs(10208) <= not b;
    layer0_outputs(10209) <= a and not b;
    layer0_outputs(10210) <= a and not b;
    layer0_outputs(10211) <= not b;
    layer0_outputs(10212) <= not (a or b);
    layer0_outputs(10213) <= not a;
    layer0_outputs(10214) <= not (a xor b);
    layer0_outputs(10215) <= b;
    layer0_outputs(10216) <= not b;
    layer0_outputs(10217) <= not (a or b);
    layer0_outputs(10218) <= a;
    layer0_outputs(10219) <= a and b;
    layer0_outputs(10220) <= b and not a;
    layer0_outputs(10221) <= a xor b;
    layer0_outputs(10222) <= not b;
    layer0_outputs(10223) <= a or b;
    layer0_outputs(10224) <= not a;
    layer0_outputs(10225) <= not (a xor b);
    layer0_outputs(10226) <= a;
    layer0_outputs(10227) <= a and not b;
    layer0_outputs(10228) <= a or b;
    layer0_outputs(10229) <= not (a or b);
    layer0_outputs(10230) <= a xor b;
    layer0_outputs(10231) <= a;
    layer0_outputs(10232) <= not (a or b);
    layer0_outputs(10233) <= not a or b;
    layer0_outputs(10234) <= not a;
    layer0_outputs(10235) <= b;
    layer0_outputs(10236) <= not (a or b);
    layer0_outputs(10237) <= not (a and b);
    layer0_outputs(10238) <= a or b;
    layer0_outputs(10239) <= not b;
    layer1_outputs(0) <= not (a or b);
    layer1_outputs(1) <= not (a or b);
    layer1_outputs(2) <= a and b;
    layer1_outputs(3) <= not b;
    layer1_outputs(4) <= b;
    layer1_outputs(5) <= not b;
    layer1_outputs(6) <= not a or b;
    layer1_outputs(7) <= a xor b;
    layer1_outputs(8) <= a or b;
    layer1_outputs(9) <= not (a or b);
    layer1_outputs(10) <= not b;
    layer1_outputs(11) <= b;
    layer1_outputs(12) <= not (a or b);
    layer1_outputs(13) <= not b;
    layer1_outputs(14) <= a;
    layer1_outputs(15) <= a and not b;
    layer1_outputs(16) <= not (a or b);
    layer1_outputs(17) <= a and not b;
    layer1_outputs(18) <= a;
    layer1_outputs(19) <= a xor b;
    layer1_outputs(20) <= a or b;
    layer1_outputs(21) <= not (a xor b);
    layer1_outputs(22) <= not b;
    layer1_outputs(23) <= a or b;
    layer1_outputs(24) <= not b;
    layer1_outputs(25) <= not b;
    layer1_outputs(26) <= not (a xor b);
    layer1_outputs(27) <= b;
    layer1_outputs(28) <= b;
    layer1_outputs(29) <= not b or a;
    layer1_outputs(30) <= a xor b;
    layer1_outputs(31) <= b;
    layer1_outputs(32) <= a xor b;
    layer1_outputs(33) <= b and not a;
    layer1_outputs(34) <= b and not a;
    layer1_outputs(35) <= a xor b;
    layer1_outputs(36) <= a and b;
    layer1_outputs(37) <= not a;
    layer1_outputs(38) <= not b;
    layer1_outputs(39) <= a;
    layer1_outputs(40) <= not b;
    layer1_outputs(41) <= b;
    layer1_outputs(42) <= not b;
    layer1_outputs(43) <= a and not b;
    layer1_outputs(44) <= a xor b;
    layer1_outputs(45) <= not (a xor b);
    layer1_outputs(46) <= not a;
    layer1_outputs(47) <= not (a xor b);
    layer1_outputs(48) <= not (a xor b);
    layer1_outputs(49) <= not (a xor b);
    layer1_outputs(50) <= a;
    layer1_outputs(51) <= not (a xor b);
    layer1_outputs(52) <= a;
    layer1_outputs(53) <= not b;
    layer1_outputs(54) <= not b;
    layer1_outputs(55) <= not (a and b);
    layer1_outputs(56) <= not a or b;
    layer1_outputs(57) <= not b;
    layer1_outputs(58) <= a or b;
    layer1_outputs(59) <= a and not b;
    layer1_outputs(60) <= not a;
    layer1_outputs(61) <= not a;
    layer1_outputs(62) <= a or b;
    layer1_outputs(63) <= not b;
    layer1_outputs(64) <= a and b;
    layer1_outputs(65) <= b;
    layer1_outputs(66) <= a xor b;
    layer1_outputs(67) <= a;
    layer1_outputs(68) <= not (a or b);
    layer1_outputs(69) <= a;
    layer1_outputs(70) <= not b or a;
    layer1_outputs(71) <= a xor b;
    layer1_outputs(72) <= not (a xor b);
    layer1_outputs(73) <= b and not a;
    layer1_outputs(74) <= a and b;
    layer1_outputs(75) <= b;
    layer1_outputs(76) <= b and not a;
    layer1_outputs(77) <= not (a xor b);
    layer1_outputs(78) <= not a;
    layer1_outputs(79) <= b;
    layer1_outputs(80) <= a or b;
    layer1_outputs(81) <= not a;
    layer1_outputs(82) <= b;
    layer1_outputs(83) <= not b;
    layer1_outputs(84) <= a and b;
    layer1_outputs(85) <= not b;
    layer1_outputs(86) <= a xor b;
    layer1_outputs(87) <= not b;
    layer1_outputs(88) <= a and not b;
    layer1_outputs(89) <= a xor b;
    layer1_outputs(90) <= not a or b;
    layer1_outputs(91) <= a and not b;
    layer1_outputs(92) <= not (a xor b);
    layer1_outputs(93) <= b;
    layer1_outputs(94) <= not a or b;
    layer1_outputs(95) <= b;
    layer1_outputs(96) <= not (a or b);
    layer1_outputs(97) <= a;
    layer1_outputs(98) <= a xor b;
    layer1_outputs(99) <= not b or a;
    layer1_outputs(100) <= not (a xor b);
    layer1_outputs(101) <= not a;
    layer1_outputs(102) <= not (a or b);
    layer1_outputs(103) <= not (a xor b);
    layer1_outputs(104) <= a and not b;
    layer1_outputs(105) <= not a;
    layer1_outputs(106) <= a xor b;
    layer1_outputs(107) <= not a or b;
    layer1_outputs(108) <= a and not b;
    layer1_outputs(109) <= not (a xor b);
    layer1_outputs(110) <= not b;
    layer1_outputs(111) <= not b or a;
    layer1_outputs(112) <= b;
    layer1_outputs(113) <= b and not a;
    layer1_outputs(114) <= a and b;
    layer1_outputs(115) <= a;
    layer1_outputs(116) <= not a;
    layer1_outputs(117) <= not (a or b);
    layer1_outputs(118) <= b and not a;
    layer1_outputs(119) <= not (a xor b);
    layer1_outputs(120) <= not a;
    layer1_outputs(121) <= a xor b;
    layer1_outputs(122) <= a or b;
    layer1_outputs(123) <= not (a xor b);
    layer1_outputs(124) <= not a;
    layer1_outputs(125) <= a xor b;
    layer1_outputs(126) <= not b or a;
    layer1_outputs(127) <= not (a or b);
    layer1_outputs(128) <= not a or b;
    layer1_outputs(129) <= not a or b;
    layer1_outputs(130) <= a xor b;
    layer1_outputs(131) <= a and b;
    layer1_outputs(132) <= a;
    layer1_outputs(133) <= a or b;
    layer1_outputs(134) <= b and not a;
    layer1_outputs(135) <= b and not a;
    layer1_outputs(136) <= a;
    layer1_outputs(137) <= a and b;
    layer1_outputs(138) <= b and not a;
    layer1_outputs(139) <= not a or b;
    layer1_outputs(140) <= not b or a;
    layer1_outputs(141) <= a and b;
    layer1_outputs(142) <= not b or a;
    layer1_outputs(143) <= a;
    layer1_outputs(144) <= a and b;
    layer1_outputs(145) <= a xor b;
    layer1_outputs(146) <= a and not b;
    layer1_outputs(147) <= not a;
    layer1_outputs(148) <= not b;
    layer1_outputs(149) <= a and not b;
    layer1_outputs(150) <= not (a xor b);
    layer1_outputs(151) <= not (a and b);
    layer1_outputs(152) <= a or b;
    layer1_outputs(153) <= not b or a;
    layer1_outputs(154) <= a xor b;
    layer1_outputs(155) <= not (a xor b);
    layer1_outputs(156) <= a;
    layer1_outputs(157) <= a xor b;
    layer1_outputs(158) <= a and not b;
    layer1_outputs(159) <= not b or a;
    layer1_outputs(160) <= not (a or b);
    layer1_outputs(161) <= not b;
    layer1_outputs(162) <= not b or a;
    layer1_outputs(163) <= a;
    layer1_outputs(164) <= not (a or b);
    layer1_outputs(165) <= not (a and b);
    layer1_outputs(166) <= not a or b;
    layer1_outputs(167) <= a;
    layer1_outputs(168) <= not (a xor b);
    layer1_outputs(169) <= not (a xor b);
    layer1_outputs(170) <= not a;
    layer1_outputs(171) <= not (a xor b);
    layer1_outputs(172) <= a xor b;
    layer1_outputs(173) <= not (a xor b);
    layer1_outputs(174) <= b;
    layer1_outputs(175) <= a;
    layer1_outputs(176) <= a xor b;
    layer1_outputs(177) <= not (a or b);
    layer1_outputs(178) <= b and not a;
    layer1_outputs(179) <= not b or a;
    layer1_outputs(180) <= a;
    layer1_outputs(181) <= a and b;
    layer1_outputs(182) <= a or b;
    layer1_outputs(183) <= not (a xor b);
    layer1_outputs(184) <= not (a or b);
    layer1_outputs(185) <= b;
    layer1_outputs(186) <= not (a and b);
    layer1_outputs(187) <= a or b;
    layer1_outputs(188) <= not (a xor b);
    layer1_outputs(189) <= a xor b;
    layer1_outputs(190) <= a and b;
    layer1_outputs(191) <= a;
    layer1_outputs(192) <= a or b;
    layer1_outputs(193) <= b;
    layer1_outputs(194) <= not b;
    layer1_outputs(195) <= not a or b;
    layer1_outputs(196) <= not a;
    layer1_outputs(197) <= not a or b;
    layer1_outputs(198) <= not (a or b);
    layer1_outputs(199) <= a and not b;
    layer1_outputs(200) <= not (a or b);
    layer1_outputs(201) <= a or b;
    layer1_outputs(202) <= not a;
    layer1_outputs(203) <= not b or a;
    layer1_outputs(204) <= a;
    layer1_outputs(205) <= not a;
    layer1_outputs(206) <= a xor b;
    layer1_outputs(207) <= a xor b;
    layer1_outputs(208) <= '0';
    layer1_outputs(209) <= a and not b;
    layer1_outputs(210) <= a or b;
    layer1_outputs(211) <= a and b;
    layer1_outputs(212) <= not a or b;
    layer1_outputs(213) <= b;
    layer1_outputs(214) <= not (a xor b);
    layer1_outputs(215) <= a or b;
    layer1_outputs(216) <= not a;
    layer1_outputs(217) <= a or b;
    layer1_outputs(218) <= a xor b;
    layer1_outputs(219) <= a and b;
    layer1_outputs(220) <= a and b;
    layer1_outputs(221) <= a and not b;
    layer1_outputs(222) <= not a or b;
    layer1_outputs(223) <= not b;
    layer1_outputs(224) <= not b;
    layer1_outputs(225) <= a and b;
    layer1_outputs(226) <= not a or b;
    layer1_outputs(227) <= not b or a;
    layer1_outputs(228) <= not a;
    layer1_outputs(229) <= a and not b;
    layer1_outputs(230) <= not (a xor b);
    layer1_outputs(231) <= not (a or b);
    layer1_outputs(232) <= b and not a;
    layer1_outputs(233) <= b;
    layer1_outputs(234) <= a xor b;
    layer1_outputs(235) <= a and b;
    layer1_outputs(236) <= a and not b;
    layer1_outputs(237) <= a xor b;
    layer1_outputs(238) <= b;
    layer1_outputs(239) <= not a or b;
    layer1_outputs(240) <= b;
    layer1_outputs(241) <= not a or b;
    layer1_outputs(242) <= b and not a;
    layer1_outputs(243) <= not (a and b);
    layer1_outputs(244) <= a or b;
    layer1_outputs(245) <= not (a xor b);
    layer1_outputs(246) <= a;
    layer1_outputs(247) <= not a or b;
    layer1_outputs(248) <= not (a xor b);
    layer1_outputs(249) <= a;
    layer1_outputs(250) <= a and not b;
    layer1_outputs(251) <= b and not a;
    layer1_outputs(252) <= not (a xor b);
    layer1_outputs(253) <= b;
    layer1_outputs(254) <= a or b;
    layer1_outputs(255) <= not (a and b);
    layer1_outputs(256) <= b and not a;
    layer1_outputs(257) <= not (a xor b);
    layer1_outputs(258) <= a or b;
    layer1_outputs(259) <= not a or b;
    layer1_outputs(260) <= not (a xor b);
    layer1_outputs(261) <= a xor b;
    layer1_outputs(262) <= not b;
    layer1_outputs(263) <= not b or a;
    layer1_outputs(264) <= a;
    layer1_outputs(265) <= not b or a;
    layer1_outputs(266) <= not a;
    layer1_outputs(267) <= not b;
    layer1_outputs(268) <= a or b;
    layer1_outputs(269) <= not b;
    layer1_outputs(270) <= '0';
    layer1_outputs(271) <= not (a and b);
    layer1_outputs(272) <= not a or b;
    layer1_outputs(273) <= a or b;
    layer1_outputs(274) <= b and not a;
    layer1_outputs(275) <= b;
    layer1_outputs(276) <= not a;
    layer1_outputs(277) <= not (a and b);
    layer1_outputs(278) <= b;
    layer1_outputs(279) <= not b or a;
    layer1_outputs(280) <= not (a xor b);
    layer1_outputs(281) <= not (a xor b);
    layer1_outputs(282) <= not a or b;
    layer1_outputs(283) <= a and b;
    layer1_outputs(284) <= b and not a;
    layer1_outputs(285) <= not b or a;
    layer1_outputs(286) <= b;
    layer1_outputs(287) <= a and b;
    layer1_outputs(288) <= not a or b;
    layer1_outputs(289) <= a or b;
    layer1_outputs(290) <= not (a xor b);
    layer1_outputs(291) <= not a or b;
    layer1_outputs(292) <= not (a or b);
    layer1_outputs(293) <= a and not b;
    layer1_outputs(294) <= not (a or b);
    layer1_outputs(295) <= not (a xor b);
    layer1_outputs(296) <= b;
    layer1_outputs(297) <= not (a and b);
    layer1_outputs(298) <= '0';
    layer1_outputs(299) <= a;
    layer1_outputs(300) <= not b;
    layer1_outputs(301) <= a and b;
    layer1_outputs(302) <= a and not b;
    layer1_outputs(303) <= a and b;
    layer1_outputs(304) <= not a or b;
    layer1_outputs(305) <= a;
    layer1_outputs(306) <= a;
    layer1_outputs(307) <= '1';
    layer1_outputs(308) <= b and not a;
    layer1_outputs(309) <= a or b;
    layer1_outputs(310) <= b;
    layer1_outputs(311) <= not (a or b);
    layer1_outputs(312) <= not b;
    layer1_outputs(313) <= a or b;
    layer1_outputs(314) <= b;
    layer1_outputs(315) <= not a;
    layer1_outputs(316) <= not b;
    layer1_outputs(317) <= a or b;
    layer1_outputs(318) <= not b;
    layer1_outputs(319) <= a and not b;
    layer1_outputs(320) <= a;
    layer1_outputs(321) <= not (a or b);
    layer1_outputs(322) <= b and not a;
    layer1_outputs(323) <= not (a xor b);
    layer1_outputs(324) <= b;
    layer1_outputs(325) <= not (a or b);
    layer1_outputs(326) <= not (a or b);
    layer1_outputs(327) <= a or b;
    layer1_outputs(328) <= not a or b;
    layer1_outputs(329) <= a xor b;
    layer1_outputs(330) <= not a or b;
    layer1_outputs(331) <= not (a and b);
    layer1_outputs(332) <= a and not b;
    layer1_outputs(333) <= b;
    layer1_outputs(334) <= not (a xor b);
    layer1_outputs(335) <= b and not a;
    layer1_outputs(336) <= b;
    layer1_outputs(337) <= a and b;
    layer1_outputs(338) <= b and not a;
    layer1_outputs(339) <= a and b;
    layer1_outputs(340) <= not (a or b);
    layer1_outputs(341) <= a and not b;
    layer1_outputs(342) <= not a or b;
    layer1_outputs(343) <= not (a and b);
    layer1_outputs(344) <= not a;
    layer1_outputs(345) <= a;
    layer1_outputs(346) <= not b;
    layer1_outputs(347) <= not (a or b);
    layer1_outputs(348) <= not a or b;
    layer1_outputs(349) <= not b;
    layer1_outputs(350) <= b;
    layer1_outputs(351) <= not (a or b);
    layer1_outputs(352) <= b and not a;
    layer1_outputs(353) <= b and not a;
    layer1_outputs(354) <= '1';
    layer1_outputs(355) <= b;
    layer1_outputs(356) <= not (a or b);
    layer1_outputs(357) <= a xor b;
    layer1_outputs(358) <= not (a xor b);
    layer1_outputs(359) <= not a;
    layer1_outputs(360) <= b;
    layer1_outputs(361) <= '1';
    layer1_outputs(362) <= a and not b;
    layer1_outputs(363) <= b;
    layer1_outputs(364) <= a;
    layer1_outputs(365) <= not (a or b);
    layer1_outputs(366) <= a;
    layer1_outputs(367) <= a;
    layer1_outputs(368) <= not (a xor b);
    layer1_outputs(369) <= a;
    layer1_outputs(370) <= not (a xor b);
    layer1_outputs(371) <= not b;
    layer1_outputs(372) <= not b or a;
    layer1_outputs(373) <= not (a and b);
    layer1_outputs(374) <= not a;
    layer1_outputs(375) <= a and b;
    layer1_outputs(376) <= a and not b;
    layer1_outputs(377) <= b;
    layer1_outputs(378) <= not a or b;
    layer1_outputs(379) <= a xor b;
    layer1_outputs(380) <= a;
    layer1_outputs(381) <= not a or b;
    layer1_outputs(382) <= not (a and b);
    layer1_outputs(383) <= not (a and b);
    layer1_outputs(384) <= a;
    layer1_outputs(385) <= not a;
    layer1_outputs(386) <= not (a and b);
    layer1_outputs(387) <= a and not b;
    layer1_outputs(388) <= b and not a;
    layer1_outputs(389) <= a;
    layer1_outputs(390) <= b;
    layer1_outputs(391) <= a and not b;
    layer1_outputs(392) <= not b or a;
    layer1_outputs(393) <= not a;
    layer1_outputs(394) <= not (a xor b);
    layer1_outputs(395) <= not (a and b);
    layer1_outputs(396) <= not a;
    layer1_outputs(397) <= a;
    layer1_outputs(398) <= b and not a;
    layer1_outputs(399) <= a or b;
    layer1_outputs(400) <= a;
    layer1_outputs(401) <= not (a or b);
    layer1_outputs(402) <= a;
    layer1_outputs(403) <= not (a and b);
    layer1_outputs(404) <= a xor b;
    layer1_outputs(405) <= a or b;
    layer1_outputs(406) <= b and not a;
    layer1_outputs(407) <= not (a xor b);
    layer1_outputs(408) <= a and not b;
    layer1_outputs(409) <= b;
    layer1_outputs(410) <= not b;
    layer1_outputs(411) <= a xor b;
    layer1_outputs(412) <= not (a or b);
    layer1_outputs(413) <= a and not b;
    layer1_outputs(414) <= a and not b;
    layer1_outputs(415) <= not b;
    layer1_outputs(416) <= not a;
    layer1_outputs(417) <= not b;
    layer1_outputs(418) <= a;
    layer1_outputs(419) <= not a or b;
    layer1_outputs(420) <= b;
    layer1_outputs(421) <= a xor b;
    layer1_outputs(422) <= not (a and b);
    layer1_outputs(423) <= a or b;
    layer1_outputs(424) <= b;
    layer1_outputs(425) <= not (a xor b);
    layer1_outputs(426) <= not a;
    layer1_outputs(427) <= not a;
    layer1_outputs(428) <= a and not b;
    layer1_outputs(429) <= not a;
    layer1_outputs(430) <= not a;
    layer1_outputs(431) <= b;
    layer1_outputs(432) <= b and not a;
    layer1_outputs(433) <= b;
    layer1_outputs(434) <= not b;
    layer1_outputs(435) <= not b or a;
    layer1_outputs(436) <= not a;
    layer1_outputs(437) <= a xor b;
    layer1_outputs(438) <= not (a or b);
    layer1_outputs(439) <= a xor b;
    layer1_outputs(440) <= not (a or b);
    layer1_outputs(441) <= not (a and b);
    layer1_outputs(442) <= not b;
    layer1_outputs(443) <= a and not b;
    layer1_outputs(444) <= not (a xor b);
    layer1_outputs(445) <= a or b;
    layer1_outputs(446) <= not (a or b);
    layer1_outputs(447) <= not (a and b);
    layer1_outputs(448) <= not (a xor b);
    layer1_outputs(449) <= a or b;
    layer1_outputs(450) <= not b or a;
    layer1_outputs(451) <= b;
    layer1_outputs(452) <= not b or a;
    layer1_outputs(453) <= a and not b;
    layer1_outputs(454) <= a and b;
    layer1_outputs(455) <= not (a or b);
    layer1_outputs(456) <= not (a and b);
    layer1_outputs(457) <= a and not b;
    layer1_outputs(458) <= not (a xor b);
    layer1_outputs(459) <= not (a and b);
    layer1_outputs(460) <= a and b;
    layer1_outputs(461) <= a or b;
    layer1_outputs(462) <= b;
    layer1_outputs(463) <= not b or a;
    layer1_outputs(464) <= b and not a;
    layer1_outputs(465) <= a or b;
    layer1_outputs(466) <= '1';
    layer1_outputs(467) <= a;
    layer1_outputs(468) <= a and not b;
    layer1_outputs(469) <= a and b;
    layer1_outputs(470) <= a or b;
    layer1_outputs(471) <= a;
    layer1_outputs(472) <= a or b;
    layer1_outputs(473) <= not a or b;
    layer1_outputs(474) <= not (a or b);
    layer1_outputs(475) <= not b;
    layer1_outputs(476) <= not b;
    layer1_outputs(477) <= not b;
    layer1_outputs(478) <= not (a and b);
    layer1_outputs(479) <= a or b;
    layer1_outputs(480) <= a xor b;
    layer1_outputs(481) <= not a;
    layer1_outputs(482) <= b;
    layer1_outputs(483) <= not (a xor b);
    layer1_outputs(484) <= a;
    layer1_outputs(485) <= b;
    layer1_outputs(486) <= not (a xor b);
    layer1_outputs(487) <= not (a xor b);
    layer1_outputs(488) <= a or b;
    layer1_outputs(489) <= b;
    layer1_outputs(490) <= b;
    layer1_outputs(491) <= a and not b;
    layer1_outputs(492) <= not a;
    layer1_outputs(493) <= not b;
    layer1_outputs(494) <= not a or b;
    layer1_outputs(495) <= not (a and b);
    layer1_outputs(496) <= not a;
    layer1_outputs(497) <= a;
    layer1_outputs(498) <= not (a xor b);
    layer1_outputs(499) <= a and b;
    layer1_outputs(500) <= b and not a;
    layer1_outputs(501) <= not b or a;
    layer1_outputs(502) <= a or b;
    layer1_outputs(503) <= not a;
    layer1_outputs(504) <= a and b;
    layer1_outputs(505) <= not (a xor b);
    layer1_outputs(506) <= a and not b;
    layer1_outputs(507) <= b;
    layer1_outputs(508) <= not a;
    layer1_outputs(509) <= a xor b;
    layer1_outputs(510) <= a and b;
    layer1_outputs(511) <= not (a or b);
    layer1_outputs(512) <= a xor b;
    layer1_outputs(513) <= not a;
    layer1_outputs(514) <= a and not b;
    layer1_outputs(515) <= a and b;
    layer1_outputs(516) <= not a;
    layer1_outputs(517) <= a xor b;
    layer1_outputs(518) <= not (a or b);
    layer1_outputs(519) <= not a;
    layer1_outputs(520) <= a and not b;
    layer1_outputs(521) <= not (a xor b);
    layer1_outputs(522) <= b and not a;
    layer1_outputs(523) <= a;
    layer1_outputs(524) <= b and not a;
    layer1_outputs(525) <= a or b;
    layer1_outputs(526) <= '0';
    layer1_outputs(527) <= not (a and b);
    layer1_outputs(528) <= b and not a;
    layer1_outputs(529) <= not (a and b);
    layer1_outputs(530) <= not b or a;
    layer1_outputs(531) <= not a;
    layer1_outputs(532) <= not (a xor b);
    layer1_outputs(533) <= a xor b;
    layer1_outputs(534) <= not a;
    layer1_outputs(535) <= not b;
    layer1_outputs(536) <= not (a and b);
    layer1_outputs(537) <= a xor b;
    layer1_outputs(538) <= not (a xor b);
    layer1_outputs(539) <= b;
    layer1_outputs(540) <= not b;
    layer1_outputs(541) <= not (a xor b);
    layer1_outputs(542) <= a or b;
    layer1_outputs(543) <= not (a and b);
    layer1_outputs(544) <= '0';
    layer1_outputs(545) <= not a;
    layer1_outputs(546) <= b and not a;
    layer1_outputs(547) <= b and not a;
    layer1_outputs(548) <= a or b;
    layer1_outputs(549) <= a xor b;
    layer1_outputs(550) <= a and not b;
    layer1_outputs(551) <= not b;
    layer1_outputs(552) <= a xor b;
    layer1_outputs(553) <= a;
    layer1_outputs(554) <= a and b;
    layer1_outputs(555) <= b;
    layer1_outputs(556) <= not b or a;
    layer1_outputs(557) <= not (a or b);
    layer1_outputs(558) <= not a or b;
    layer1_outputs(559) <= not (a xor b);
    layer1_outputs(560) <= a or b;
    layer1_outputs(561) <= b and not a;
    layer1_outputs(562) <= b;
    layer1_outputs(563) <= a;
    layer1_outputs(564) <= not a;
    layer1_outputs(565) <= not b;
    layer1_outputs(566) <= a;
    layer1_outputs(567) <= a and not b;
    layer1_outputs(568) <= a xor b;
    layer1_outputs(569) <= b;
    layer1_outputs(570) <= a xor b;
    layer1_outputs(571) <= not b;
    layer1_outputs(572) <= not b;
    layer1_outputs(573) <= a xor b;
    layer1_outputs(574) <= b and not a;
    layer1_outputs(575) <= b;
    layer1_outputs(576) <= a or b;
    layer1_outputs(577) <= '0';
    layer1_outputs(578) <= a and not b;
    layer1_outputs(579) <= not b;
    layer1_outputs(580) <= b and not a;
    layer1_outputs(581) <= b;
    layer1_outputs(582) <= not b or a;
    layer1_outputs(583) <= not (a and b);
    layer1_outputs(584) <= not (a and b);
    layer1_outputs(585) <= not b or a;
    layer1_outputs(586) <= not b;
    layer1_outputs(587) <= not (a xor b);
    layer1_outputs(588) <= not a or b;
    layer1_outputs(589) <= not b;
    layer1_outputs(590) <= a and not b;
    layer1_outputs(591) <= b and not a;
    layer1_outputs(592) <= a and b;
    layer1_outputs(593) <= not (a or b);
    layer1_outputs(594) <= not (a xor b);
    layer1_outputs(595) <= a;
    layer1_outputs(596) <= not (a and b);
    layer1_outputs(597) <= a and not b;
    layer1_outputs(598) <= not a or b;
    layer1_outputs(599) <= a xor b;
    layer1_outputs(600) <= not b or a;
    layer1_outputs(601) <= b;
    layer1_outputs(602) <= a;
    layer1_outputs(603) <= not b;
    layer1_outputs(604) <= a or b;
    layer1_outputs(605) <= b;
    layer1_outputs(606) <= b and not a;
    layer1_outputs(607) <= not (a or b);
    layer1_outputs(608) <= a and b;
    layer1_outputs(609) <= not a or b;
    layer1_outputs(610) <= a or b;
    layer1_outputs(611) <= not (a and b);
    layer1_outputs(612) <= not (a and b);
    layer1_outputs(613) <= b and not a;
    layer1_outputs(614) <= not b;
    layer1_outputs(615) <= not (a and b);
    layer1_outputs(616) <= b;
    layer1_outputs(617) <= a xor b;
    layer1_outputs(618) <= not a;
    layer1_outputs(619) <= not a or b;
    layer1_outputs(620) <= not (a and b);
    layer1_outputs(621) <= not a;
    layer1_outputs(622) <= not a;
    layer1_outputs(623) <= not b;
    layer1_outputs(624) <= not b;
    layer1_outputs(625) <= b;
    layer1_outputs(626) <= not (a or b);
    layer1_outputs(627) <= a and b;
    layer1_outputs(628) <= a and b;
    layer1_outputs(629) <= not (a or b);
    layer1_outputs(630) <= a xor b;
    layer1_outputs(631) <= b and not a;
    layer1_outputs(632) <= b;
    layer1_outputs(633) <= b and not a;
    layer1_outputs(634) <= a;
    layer1_outputs(635) <= not (a or b);
    layer1_outputs(636) <= b and not a;
    layer1_outputs(637) <= a xor b;
    layer1_outputs(638) <= not (a xor b);
    layer1_outputs(639) <= a;
    layer1_outputs(640) <= a xor b;
    layer1_outputs(641) <= '0';
    layer1_outputs(642) <= not (a or b);
    layer1_outputs(643) <= '1';
    layer1_outputs(644) <= not b;
    layer1_outputs(645) <= not b;
    layer1_outputs(646) <= b and not a;
    layer1_outputs(647) <= b;
    layer1_outputs(648) <= a xor b;
    layer1_outputs(649) <= a or b;
    layer1_outputs(650) <= not a or b;
    layer1_outputs(651) <= a and not b;
    layer1_outputs(652) <= b;
    layer1_outputs(653) <= b and not a;
    layer1_outputs(654) <= not a or b;
    layer1_outputs(655) <= a and b;
    layer1_outputs(656) <= '0';
    layer1_outputs(657) <= b;
    layer1_outputs(658) <= a xor b;
    layer1_outputs(659) <= not (a or b);
    layer1_outputs(660) <= not a or b;
    layer1_outputs(661) <= a xor b;
    layer1_outputs(662) <= a and not b;
    layer1_outputs(663) <= not (a xor b);
    layer1_outputs(664) <= not (a xor b);
    layer1_outputs(665) <= a or b;
    layer1_outputs(666) <= a xor b;
    layer1_outputs(667) <= not b;
    layer1_outputs(668) <= a;
    layer1_outputs(669) <= not (a xor b);
    layer1_outputs(670) <= b and not a;
    layer1_outputs(671) <= not a;
    layer1_outputs(672) <= not (a xor b);
    layer1_outputs(673) <= not (a xor b);
    layer1_outputs(674) <= not b or a;
    layer1_outputs(675) <= a xor b;
    layer1_outputs(676) <= b;
    layer1_outputs(677) <= not a or b;
    layer1_outputs(678) <= a xor b;
    layer1_outputs(679) <= a or b;
    layer1_outputs(680) <= not b or a;
    layer1_outputs(681) <= a and b;
    layer1_outputs(682) <= '1';
    layer1_outputs(683) <= a;
    layer1_outputs(684) <= not (a xor b);
    layer1_outputs(685) <= not b or a;
    layer1_outputs(686) <= b and not a;
    layer1_outputs(687) <= b;
    layer1_outputs(688) <= not a or b;
    layer1_outputs(689) <= a;
    layer1_outputs(690) <= a;
    layer1_outputs(691) <= a;
    layer1_outputs(692) <= a and not b;
    layer1_outputs(693) <= a and not b;
    layer1_outputs(694) <= not a;
    layer1_outputs(695) <= a or b;
    layer1_outputs(696) <= a xor b;
    layer1_outputs(697) <= not (a xor b);
    layer1_outputs(698) <= a xor b;
    layer1_outputs(699) <= not (a or b);
    layer1_outputs(700) <= not (a or b);
    layer1_outputs(701) <= not (a xor b);
    layer1_outputs(702) <= a;
    layer1_outputs(703) <= not b or a;
    layer1_outputs(704) <= not (a and b);
    layer1_outputs(705) <= a and b;
    layer1_outputs(706) <= b and not a;
    layer1_outputs(707) <= not (a or b);
    layer1_outputs(708) <= a xor b;
    layer1_outputs(709) <= not (a xor b);
    layer1_outputs(710) <= not a;
    layer1_outputs(711) <= a;
    layer1_outputs(712) <= not a;
    layer1_outputs(713) <= a and b;
    layer1_outputs(714) <= not (a and b);
    layer1_outputs(715) <= b;
    layer1_outputs(716) <= b and not a;
    layer1_outputs(717) <= a;
    layer1_outputs(718) <= not b;
    layer1_outputs(719) <= not a;
    layer1_outputs(720) <= a and b;
    layer1_outputs(721) <= a xor b;
    layer1_outputs(722) <= a or b;
    layer1_outputs(723) <= a;
    layer1_outputs(724) <= a xor b;
    layer1_outputs(725) <= not b;
    layer1_outputs(726) <= a xor b;
    layer1_outputs(727) <= a xor b;
    layer1_outputs(728) <= a or b;
    layer1_outputs(729) <= not b or a;
    layer1_outputs(730) <= not b;
    layer1_outputs(731) <= a and b;
    layer1_outputs(732) <= a or b;
    layer1_outputs(733) <= not a or b;
    layer1_outputs(734) <= a or b;
    layer1_outputs(735) <= not b;
    layer1_outputs(736) <= a and b;
    layer1_outputs(737) <= b and not a;
    layer1_outputs(738) <= a xor b;
    layer1_outputs(739) <= not (a and b);
    layer1_outputs(740) <= not b;
    layer1_outputs(741) <= b;
    layer1_outputs(742) <= a and not b;
    layer1_outputs(743) <= not a;
    layer1_outputs(744) <= not a or b;
    layer1_outputs(745) <= a xor b;
    layer1_outputs(746) <= not a or b;
    layer1_outputs(747) <= a;
    layer1_outputs(748) <= a;
    layer1_outputs(749) <= not b or a;
    layer1_outputs(750) <= a;
    layer1_outputs(751) <= not (a xor b);
    layer1_outputs(752) <= not b;
    layer1_outputs(753) <= not (a xor b);
    layer1_outputs(754) <= b and not a;
    layer1_outputs(755) <= b and not a;
    layer1_outputs(756) <= not (a and b);
    layer1_outputs(757) <= a and b;
    layer1_outputs(758) <= not a;
    layer1_outputs(759) <= not b or a;
    layer1_outputs(760) <= a and b;
    layer1_outputs(761) <= b and not a;
    layer1_outputs(762) <= a xor b;
    layer1_outputs(763) <= not (a or b);
    layer1_outputs(764) <= a xor b;
    layer1_outputs(765) <= not b;
    layer1_outputs(766) <= b;
    layer1_outputs(767) <= not (a or b);
    layer1_outputs(768) <= a and b;
    layer1_outputs(769) <= a xor b;
    layer1_outputs(770) <= not a or b;
    layer1_outputs(771) <= not a;
    layer1_outputs(772) <= not a;
    layer1_outputs(773) <= a or b;
    layer1_outputs(774) <= not (a xor b);
    layer1_outputs(775) <= a xor b;
    layer1_outputs(776) <= not b;
    layer1_outputs(777) <= not (a or b);
    layer1_outputs(778) <= a and not b;
    layer1_outputs(779) <= not (a xor b);
    layer1_outputs(780) <= not a;
    layer1_outputs(781) <= not (a and b);
    layer1_outputs(782) <= b;
    layer1_outputs(783) <= not a or b;
    layer1_outputs(784) <= a and b;
    layer1_outputs(785) <= not b;
    layer1_outputs(786) <= not b or a;
    layer1_outputs(787) <= not (a or b);
    layer1_outputs(788) <= not b;
    layer1_outputs(789) <= not a or b;
    layer1_outputs(790) <= a or b;
    layer1_outputs(791) <= not b;
    layer1_outputs(792) <= not a or b;
    layer1_outputs(793) <= a and b;
    layer1_outputs(794) <= a xor b;
    layer1_outputs(795) <= a;
    layer1_outputs(796) <= a or b;
    layer1_outputs(797) <= not a;
    layer1_outputs(798) <= a and b;
    layer1_outputs(799) <= a or b;
    layer1_outputs(800) <= a;
    layer1_outputs(801) <= a and not b;
    layer1_outputs(802) <= b;
    layer1_outputs(803) <= a and not b;
    layer1_outputs(804) <= not (a or b);
    layer1_outputs(805) <= not b;
    layer1_outputs(806) <= not a or b;
    layer1_outputs(807) <= not b or a;
    layer1_outputs(808) <= a xor b;
    layer1_outputs(809) <= a and b;
    layer1_outputs(810) <= not (a or b);
    layer1_outputs(811) <= b and not a;
    layer1_outputs(812) <= b;
    layer1_outputs(813) <= a and not b;
    layer1_outputs(814) <= not (a and b);
    layer1_outputs(815) <= not a or b;
    layer1_outputs(816) <= '0';
    layer1_outputs(817) <= not (a and b);
    layer1_outputs(818) <= not a;
    layer1_outputs(819) <= a;
    layer1_outputs(820) <= b;
    layer1_outputs(821) <= not a;
    layer1_outputs(822) <= not b;
    layer1_outputs(823) <= not (a and b);
    layer1_outputs(824) <= a or b;
    layer1_outputs(825) <= not b;
    layer1_outputs(826) <= not a or b;
    layer1_outputs(827) <= a and not b;
    layer1_outputs(828) <= a;
    layer1_outputs(829) <= a and not b;
    layer1_outputs(830) <= not a;
    layer1_outputs(831) <= not b;
    layer1_outputs(832) <= not a;
    layer1_outputs(833) <= not (a and b);
    layer1_outputs(834) <= a or b;
    layer1_outputs(835) <= a xor b;
    layer1_outputs(836) <= a or b;
    layer1_outputs(837) <= b and not a;
    layer1_outputs(838) <= not a;
    layer1_outputs(839) <= not b or a;
    layer1_outputs(840) <= not b;
    layer1_outputs(841) <= not b or a;
    layer1_outputs(842) <= a and b;
    layer1_outputs(843) <= a or b;
    layer1_outputs(844) <= a xor b;
    layer1_outputs(845) <= not b;
    layer1_outputs(846) <= b;
    layer1_outputs(847) <= a;
    layer1_outputs(848) <= b;
    layer1_outputs(849) <= not b;
    layer1_outputs(850) <= not a;
    layer1_outputs(851) <= a and b;
    layer1_outputs(852) <= a and b;
    layer1_outputs(853) <= not (a or b);
    layer1_outputs(854) <= not b or a;
    layer1_outputs(855) <= not b or a;
    layer1_outputs(856) <= not a;
    layer1_outputs(857) <= a;
    layer1_outputs(858) <= not (a xor b);
    layer1_outputs(859) <= a and b;
    layer1_outputs(860) <= not (a xor b);
    layer1_outputs(861) <= not (a and b);
    layer1_outputs(862) <= a and b;
    layer1_outputs(863) <= not b;
    layer1_outputs(864) <= a or b;
    layer1_outputs(865) <= not a or b;
    layer1_outputs(866) <= a xor b;
    layer1_outputs(867) <= not a;
    layer1_outputs(868) <= not (a and b);
    layer1_outputs(869) <= a xor b;
    layer1_outputs(870) <= a or b;
    layer1_outputs(871) <= a and b;
    layer1_outputs(872) <= b and not a;
    layer1_outputs(873) <= a;
    layer1_outputs(874) <= not a;
    layer1_outputs(875) <= a and not b;
    layer1_outputs(876) <= a xor b;
    layer1_outputs(877) <= not a or b;
    layer1_outputs(878) <= not (a or b);
    layer1_outputs(879) <= not a;
    layer1_outputs(880) <= b and not a;
    layer1_outputs(881) <= not b or a;
    layer1_outputs(882) <= a xor b;
    layer1_outputs(883) <= not a or b;
    layer1_outputs(884) <= a and b;
    layer1_outputs(885) <= not a;
    layer1_outputs(886) <= a and not b;
    layer1_outputs(887) <= not (a xor b);
    layer1_outputs(888) <= not b or a;
    layer1_outputs(889) <= '1';
    layer1_outputs(890) <= not (a or b);
    layer1_outputs(891) <= b and not a;
    layer1_outputs(892) <= a;
    layer1_outputs(893) <= not (a xor b);
    layer1_outputs(894) <= not a;
    layer1_outputs(895) <= a or b;
    layer1_outputs(896) <= a;
    layer1_outputs(897) <= a xor b;
    layer1_outputs(898) <= a;
    layer1_outputs(899) <= a and b;
    layer1_outputs(900) <= '0';
    layer1_outputs(901) <= a;
    layer1_outputs(902) <= a or b;
    layer1_outputs(903) <= not (a or b);
    layer1_outputs(904) <= not (a or b);
    layer1_outputs(905) <= not a;
    layer1_outputs(906) <= not b or a;
    layer1_outputs(907) <= not (a or b);
    layer1_outputs(908) <= not b;
    layer1_outputs(909) <= b and not a;
    layer1_outputs(910) <= not a or b;
    layer1_outputs(911) <= not b or a;
    layer1_outputs(912) <= b;
    layer1_outputs(913) <= a;
    layer1_outputs(914) <= '1';
    layer1_outputs(915) <= not (a and b);
    layer1_outputs(916) <= b and not a;
    layer1_outputs(917) <= not b;
    layer1_outputs(918) <= b and not a;
    layer1_outputs(919) <= not (a or b);
    layer1_outputs(920) <= b and not a;
    layer1_outputs(921) <= not (a or b);
    layer1_outputs(922) <= b and not a;
    layer1_outputs(923) <= not a or b;
    layer1_outputs(924) <= b and not a;
    layer1_outputs(925) <= not b or a;
    layer1_outputs(926) <= not b;
    layer1_outputs(927) <= not (a xor b);
    layer1_outputs(928) <= not a;
    layer1_outputs(929) <= not (a xor b);
    layer1_outputs(930) <= b and not a;
    layer1_outputs(931) <= a xor b;
    layer1_outputs(932) <= b and not a;
    layer1_outputs(933) <= not b;
    layer1_outputs(934) <= b;
    layer1_outputs(935) <= a;
    layer1_outputs(936) <= not a or b;
    layer1_outputs(937) <= not (a or b);
    layer1_outputs(938) <= not b;
    layer1_outputs(939) <= not a;
    layer1_outputs(940) <= b and not a;
    layer1_outputs(941) <= a;
    layer1_outputs(942) <= b;
    layer1_outputs(943) <= not (a xor b);
    layer1_outputs(944) <= a;
    layer1_outputs(945) <= a and not b;
    layer1_outputs(946) <= not (a and b);
    layer1_outputs(947) <= not (a xor b);
    layer1_outputs(948) <= '0';
    layer1_outputs(949) <= a;
    layer1_outputs(950) <= not b or a;
    layer1_outputs(951) <= not a;
    layer1_outputs(952) <= not (a xor b);
    layer1_outputs(953) <= a xor b;
    layer1_outputs(954) <= b;
    layer1_outputs(955) <= a and not b;
    layer1_outputs(956) <= b;
    layer1_outputs(957) <= not b or a;
    layer1_outputs(958) <= '0';
    layer1_outputs(959) <= not a;
    layer1_outputs(960) <= not a;
    layer1_outputs(961) <= not b;
    layer1_outputs(962) <= not b;
    layer1_outputs(963) <= not b;
    layer1_outputs(964) <= not a or b;
    layer1_outputs(965) <= not (a or b);
    layer1_outputs(966) <= not (a xor b);
    layer1_outputs(967) <= a xor b;
    layer1_outputs(968) <= not a;
    layer1_outputs(969) <= a and b;
    layer1_outputs(970) <= a;
    layer1_outputs(971) <= '0';
    layer1_outputs(972) <= not b;
    layer1_outputs(973) <= a xor b;
    layer1_outputs(974) <= a xor b;
    layer1_outputs(975) <= b;
    layer1_outputs(976) <= a;
    layer1_outputs(977) <= b and not a;
    layer1_outputs(978) <= b;
    layer1_outputs(979) <= not (a and b);
    layer1_outputs(980) <= a or b;
    layer1_outputs(981) <= b and not a;
    layer1_outputs(982) <= not (a or b);
    layer1_outputs(983) <= not a;
    layer1_outputs(984) <= a xor b;
    layer1_outputs(985) <= a xor b;
    layer1_outputs(986) <= a xor b;
    layer1_outputs(987) <= not a;
    layer1_outputs(988) <= not b;
    layer1_outputs(989) <= a and not b;
    layer1_outputs(990) <= not b;
    layer1_outputs(991) <= not b;
    layer1_outputs(992) <= not b;
    layer1_outputs(993) <= not (a xor b);
    layer1_outputs(994) <= not b or a;
    layer1_outputs(995) <= not (a or b);
    layer1_outputs(996) <= not (a and b);
    layer1_outputs(997) <= b;
    layer1_outputs(998) <= not (a xor b);
    layer1_outputs(999) <= not a;
    layer1_outputs(1000) <= not (a xor b);
    layer1_outputs(1001) <= not a or b;
    layer1_outputs(1002) <= not b or a;
    layer1_outputs(1003) <= a or b;
    layer1_outputs(1004) <= a;
    layer1_outputs(1005) <= not b;
    layer1_outputs(1006) <= not (a and b);
    layer1_outputs(1007) <= a and not b;
    layer1_outputs(1008) <= not a;
    layer1_outputs(1009) <= a and not b;
    layer1_outputs(1010) <= not (a and b);
    layer1_outputs(1011) <= a and b;
    layer1_outputs(1012) <= b and not a;
    layer1_outputs(1013) <= not b or a;
    layer1_outputs(1014) <= a and b;
    layer1_outputs(1015) <= a;
    layer1_outputs(1016) <= b and not a;
    layer1_outputs(1017) <= not (a xor b);
    layer1_outputs(1018) <= b;
    layer1_outputs(1019) <= a or b;
    layer1_outputs(1020) <= not (a and b);
    layer1_outputs(1021) <= not a;
    layer1_outputs(1022) <= b and not a;
    layer1_outputs(1023) <= not a or b;
    layer1_outputs(1024) <= '0';
    layer1_outputs(1025) <= not (a xor b);
    layer1_outputs(1026) <= not b;
    layer1_outputs(1027) <= not b;
    layer1_outputs(1028) <= not b or a;
    layer1_outputs(1029) <= a xor b;
    layer1_outputs(1030) <= b;
    layer1_outputs(1031) <= a and b;
    layer1_outputs(1032) <= not (a and b);
    layer1_outputs(1033) <= a xor b;
    layer1_outputs(1034) <= a and not b;
    layer1_outputs(1035) <= a and not b;
    layer1_outputs(1036) <= not b;
    layer1_outputs(1037) <= '1';
    layer1_outputs(1038) <= not (a xor b);
    layer1_outputs(1039) <= not (a xor b);
    layer1_outputs(1040) <= a or b;
    layer1_outputs(1041) <= not a;
    layer1_outputs(1042) <= a;
    layer1_outputs(1043) <= a and not b;
    layer1_outputs(1044) <= not a or b;
    layer1_outputs(1045) <= '1';
    layer1_outputs(1046) <= not (a and b);
    layer1_outputs(1047) <= not a;
    layer1_outputs(1048) <= not b;
    layer1_outputs(1049) <= a and not b;
    layer1_outputs(1050) <= not (a and b);
    layer1_outputs(1051) <= a and b;
    layer1_outputs(1052) <= not b;
    layer1_outputs(1053) <= a xor b;
    layer1_outputs(1054) <= not b or a;
    layer1_outputs(1055) <= not b or a;
    layer1_outputs(1056) <= a xor b;
    layer1_outputs(1057) <= a;
    layer1_outputs(1058) <= a xor b;
    layer1_outputs(1059) <= not (a or b);
    layer1_outputs(1060) <= a and b;
    layer1_outputs(1061) <= not a or b;
    layer1_outputs(1062) <= b;
    layer1_outputs(1063) <= not b or a;
    layer1_outputs(1064) <= a xor b;
    layer1_outputs(1065) <= not (a xor b);
    layer1_outputs(1066) <= a;
    layer1_outputs(1067) <= a and not b;
    layer1_outputs(1068) <= not a or b;
    layer1_outputs(1069) <= not a;
    layer1_outputs(1070) <= a and not b;
    layer1_outputs(1071) <= '0';
    layer1_outputs(1072) <= not b;
    layer1_outputs(1073) <= not a;
    layer1_outputs(1074) <= a and b;
    layer1_outputs(1075) <= not a or b;
    layer1_outputs(1076) <= a or b;
    layer1_outputs(1077) <= not (a and b);
    layer1_outputs(1078) <= a and b;
    layer1_outputs(1079) <= not b or a;
    layer1_outputs(1080) <= not b;
    layer1_outputs(1081) <= a or b;
    layer1_outputs(1082) <= not (a xor b);
    layer1_outputs(1083) <= not (a or b);
    layer1_outputs(1084) <= b;
    layer1_outputs(1085) <= b and not a;
    layer1_outputs(1086) <= b;
    layer1_outputs(1087) <= not b;
    layer1_outputs(1088) <= b and not a;
    layer1_outputs(1089) <= not a;
    layer1_outputs(1090) <= b;
    layer1_outputs(1091) <= not b;
    layer1_outputs(1092) <= a xor b;
    layer1_outputs(1093) <= not (a xor b);
    layer1_outputs(1094) <= not (a or b);
    layer1_outputs(1095) <= a and not b;
    layer1_outputs(1096) <= not (a and b);
    layer1_outputs(1097) <= not (a and b);
    layer1_outputs(1098) <= not (a xor b);
    layer1_outputs(1099) <= not a;
    layer1_outputs(1100) <= a;
    layer1_outputs(1101) <= not a or b;
    layer1_outputs(1102) <= a and not b;
    layer1_outputs(1103) <= not a;
    layer1_outputs(1104) <= a;
    layer1_outputs(1105) <= not b or a;
    layer1_outputs(1106) <= a xor b;
    layer1_outputs(1107) <= a;
    layer1_outputs(1108) <= b;
    layer1_outputs(1109) <= not b or a;
    layer1_outputs(1110) <= a;
    layer1_outputs(1111) <= a;
    layer1_outputs(1112) <= b;
    layer1_outputs(1113) <= not b;
    layer1_outputs(1114) <= a xor b;
    layer1_outputs(1115) <= b;
    layer1_outputs(1116) <= not b;
    layer1_outputs(1117) <= not (a xor b);
    layer1_outputs(1118) <= b and not a;
    layer1_outputs(1119) <= a;
    layer1_outputs(1120) <= b;
    layer1_outputs(1121) <= b;
    layer1_outputs(1122) <= not a;
    layer1_outputs(1123) <= b;
    layer1_outputs(1124) <= not b;
    layer1_outputs(1125) <= a;
    layer1_outputs(1126) <= a and not b;
    layer1_outputs(1127) <= not (a or b);
    layer1_outputs(1128) <= not b;
    layer1_outputs(1129) <= a or b;
    layer1_outputs(1130) <= not b or a;
    layer1_outputs(1131) <= a;
    layer1_outputs(1132) <= b and not a;
    layer1_outputs(1133) <= b;
    layer1_outputs(1134) <= b;
    layer1_outputs(1135) <= not (a xor b);
    layer1_outputs(1136) <= b and not a;
    layer1_outputs(1137) <= not (a or b);
    layer1_outputs(1138) <= a or b;
    layer1_outputs(1139) <= b;
    layer1_outputs(1140) <= not a;
    layer1_outputs(1141) <= a or b;
    layer1_outputs(1142) <= a or b;
    layer1_outputs(1143) <= a and b;
    layer1_outputs(1144) <= b;
    layer1_outputs(1145) <= b;
    layer1_outputs(1146) <= not b or a;
    layer1_outputs(1147) <= not b;
    layer1_outputs(1148) <= b;
    layer1_outputs(1149) <= a;
    layer1_outputs(1150) <= a and b;
    layer1_outputs(1151) <= a;
    layer1_outputs(1152) <= a;
    layer1_outputs(1153) <= not (a or b);
    layer1_outputs(1154) <= b;
    layer1_outputs(1155) <= a xor b;
    layer1_outputs(1156) <= b and not a;
    layer1_outputs(1157) <= not b;
    layer1_outputs(1158) <= '0';
    layer1_outputs(1159) <= not (a xor b);
    layer1_outputs(1160) <= '1';
    layer1_outputs(1161) <= a and not b;
    layer1_outputs(1162) <= not b;
    layer1_outputs(1163) <= not a;
    layer1_outputs(1164) <= b and not a;
    layer1_outputs(1165) <= b and not a;
    layer1_outputs(1166) <= not (a xor b);
    layer1_outputs(1167) <= not (a or b);
    layer1_outputs(1168) <= not b;
    layer1_outputs(1169) <= not (a and b);
    layer1_outputs(1170) <= a;
    layer1_outputs(1171) <= a and not b;
    layer1_outputs(1172) <= not (a and b);
    layer1_outputs(1173) <= a;
    layer1_outputs(1174) <= a xor b;
    layer1_outputs(1175) <= not b;
    layer1_outputs(1176) <= b;
    layer1_outputs(1177) <= a and b;
    layer1_outputs(1178) <= b and not a;
    layer1_outputs(1179) <= b;
    layer1_outputs(1180) <= a xor b;
    layer1_outputs(1181) <= a;
    layer1_outputs(1182) <= not (a xor b);
    layer1_outputs(1183) <= a and b;
    layer1_outputs(1184) <= a or b;
    layer1_outputs(1185) <= not b;
    layer1_outputs(1186) <= not a;
    layer1_outputs(1187) <= not b or a;
    layer1_outputs(1188) <= not b;
    layer1_outputs(1189) <= not (a and b);
    layer1_outputs(1190) <= not a;
    layer1_outputs(1191) <= not a or b;
    layer1_outputs(1192) <= not (a xor b);
    layer1_outputs(1193) <= a and not b;
    layer1_outputs(1194) <= b;
    layer1_outputs(1195) <= a xor b;
    layer1_outputs(1196) <= not b;
    layer1_outputs(1197) <= a;
    layer1_outputs(1198) <= not b;
    layer1_outputs(1199) <= a and b;
    layer1_outputs(1200) <= b and not a;
    layer1_outputs(1201) <= not (a xor b);
    layer1_outputs(1202) <= a;
    layer1_outputs(1203) <= not b;
    layer1_outputs(1204) <= a and b;
    layer1_outputs(1205) <= a or b;
    layer1_outputs(1206) <= b;
    layer1_outputs(1207) <= a xor b;
    layer1_outputs(1208) <= a and b;
    layer1_outputs(1209) <= not a;
    layer1_outputs(1210) <= b;
    layer1_outputs(1211) <= not (a or b);
    layer1_outputs(1212) <= not (a and b);
    layer1_outputs(1213) <= a;
    layer1_outputs(1214) <= a;
    layer1_outputs(1215) <= not b or a;
    layer1_outputs(1216) <= not (a xor b);
    layer1_outputs(1217) <= a and not b;
    layer1_outputs(1218) <= not a or b;
    layer1_outputs(1219) <= not (a and b);
    layer1_outputs(1220) <= not a;
    layer1_outputs(1221) <= not a or b;
    layer1_outputs(1222) <= a;
    layer1_outputs(1223) <= b;
    layer1_outputs(1224) <= b and not a;
    layer1_outputs(1225) <= not b or a;
    layer1_outputs(1226) <= not a;
    layer1_outputs(1227) <= a xor b;
    layer1_outputs(1228) <= b;
    layer1_outputs(1229) <= not b;
    layer1_outputs(1230) <= not a;
    layer1_outputs(1231) <= b;
    layer1_outputs(1232) <= not a or b;
    layer1_outputs(1233) <= not a;
    layer1_outputs(1234) <= a and not b;
    layer1_outputs(1235) <= not b;
    layer1_outputs(1236) <= a and b;
    layer1_outputs(1237) <= not b or a;
    layer1_outputs(1238) <= not (a or b);
    layer1_outputs(1239) <= a xor b;
    layer1_outputs(1240) <= a or b;
    layer1_outputs(1241) <= b and not a;
    layer1_outputs(1242) <= not a;
    layer1_outputs(1243) <= not b;
    layer1_outputs(1244) <= b and not a;
    layer1_outputs(1245) <= not (a or b);
    layer1_outputs(1246) <= b;
    layer1_outputs(1247) <= b and not a;
    layer1_outputs(1248) <= not b;
    layer1_outputs(1249) <= a and b;
    layer1_outputs(1250) <= a xor b;
    layer1_outputs(1251) <= b;
    layer1_outputs(1252) <= not a or b;
    layer1_outputs(1253) <= not b;
    layer1_outputs(1254) <= not a;
    layer1_outputs(1255) <= a and b;
    layer1_outputs(1256) <= b;
    layer1_outputs(1257) <= not (a and b);
    layer1_outputs(1258) <= not a or b;
    layer1_outputs(1259) <= not a;
    layer1_outputs(1260) <= a;
    layer1_outputs(1261) <= not a or b;
    layer1_outputs(1262) <= a;
    layer1_outputs(1263) <= not (a and b);
    layer1_outputs(1264) <= not b;
    layer1_outputs(1265) <= not a;
    layer1_outputs(1266) <= b;
    layer1_outputs(1267) <= not a or b;
    layer1_outputs(1268) <= not b;
    layer1_outputs(1269) <= not a or b;
    layer1_outputs(1270) <= not (a or b);
    layer1_outputs(1271) <= not (a and b);
    layer1_outputs(1272) <= not (a xor b);
    layer1_outputs(1273) <= not a;
    layer1_outputs(1274) <= not b;
    layer1_outputs(1275) <= a xor b;
    layer1_outputs(1276) <= a and not b;
    layer1_outputs(1277) <= a and b;
    layer1_outputs(1278) <= b;
    layer1_outputs(1279) <= b and not a;
    layer1_outputs(1280) <= not a;
    layer1_outputs(1281) <= not (a xor b);
    layer1_outputs(1282) <= not b or a;
    layer1_outputs(1283) <= a;
    layer1_outputs(1284) <= not b;
    layer1_outputs(1285) <= a and b;
    layer1_outputs(1286) <= not (a xor b);
    layer1_outputs(1287) <= not b;
    layer1_outputs(1288) <= not (a xor b);
    layer1_outputs(1289) <= b;
    layer1_outputs(1290) <= a and b;
    layer1_outputs(1291) <= a or b;
    layer1_outputs(1292) <= b;
    layer1_outputs(1293) <= not b or a;
    layer1_outputs(1294) <= not (a or b);
    layer1_outputs(1295) <= a or b;
    layer1_outputs(1296) <= b and not a;
    layer1_outputs(1297) <= a;
    layer1_outputs(1298) <= b and not a;
    layer1_outputs(1299) <= not (a and b);
    layer1_outputs(1300) <= not b;
    layer1_outputs(1301) <= not a or b;
    layer1_outputs(1302) <= a;
    layer1_outputs(1303) <= not b;
    layer1_outputs(1304) <= not a or b;
    layer1_outputs(1305) <= not b;
    layer1_outputs(1306) <= a xor b;
    layer1_outputs(1307) <= not a or b;
    layer1_outputs(1308) <= b and not a;
    layer1_outputs(1309) <= not b or a;
    layer1_outputs(1310) <= not (a xor b);
    layer1_outputs(1311) <= '1';
    layer1_outputs(1312) <= a and b;
    layer1_outputs(1313) <= '0';
    layer1_outputs(1314) <= '1';
    layer1_outputs(1315) <= a or b;
    layer1_outputs(1316) <= a and not b;
    layer1_outputs(1317) <= a xor b;
    layer1_outputs(1318) <= not a or b;
    layer1_outputs(1319) <= b;
    layer1_outputs(1320) <= not a or b;
    layer1_outputs(1321) <= a or b;
    layer1_outputs(1322) <= a xor b;
    layer1_outputs(1323) <= not a;
    layer1_outputs(1324) <= not (a or b);
    layer1_outputs(1325) <= a and b;
    layer1_outputs(1326) <= not a;
    layer1_outputs(1327) <= not b;
    layer1_outputs(1328) <= not b or a;
    layer1_outputs(1329) <= a;
    layer1_outputs(1330) <= not (a or b);
    layer1_outputs(1331) <= a or b;
    layer1_outputs(1332) <= b and not a;
    layer1_outputs(1333) <= a and b;
    layer1_outputs(1334) <= not (a or b);
    layer1_outputs(1335) <= not b or a;
    layer1_outputs(1336) <= a or b;
    layer1_outputs(1337) <= not b;
    layer1_outputs(1338) <= a xor b;
    layer1_outputs(1339) <= '0';
    layer1_outputs(1340) <= not b;
    layer1_outputs(1341) <= b;
    layer1_outputs(1342) <= b;
    layer1_outputs(1343) <= not a;
    layer1_outputs(1344) <= a xor b;
    layer1_outputs(1345) <= not (a and b);
    layer1_outputs(1346) <= a and b;
    layer1_outputs(1347) <= not (a xor b);
    layer1_outputs(1348) <= not a;
    layer1_outputs(1349) <= b and not a;
    layer1_outputs(1350) <= a and not b;
    layer1_outputs(1351) <= a or b;
    layer1_outputs(1352) <= not (a and b);
    layer1_outputs(1353) <= b and not a;
    layer1_outputs(1354) <= a;
    layer1_outputs(1355) <= a or b;
    layer1_outputs(1356) <= not (a xor b);
    layer1_outputs(1357) <= a and not b;
    layer1_outputs(1358) <= not b or a;
    layer1_outputs(1359) <= not b;
    layer1_outputs(1360) <= not (a xor b);
    layer1_outputs(1361) <= a and not b;
    layer1_outputs(1362) <= a;
    layer1_outputs(1363) <= not b or a;
    layer1_outputs(1364) <= not b;
    layer1_outputs(1365) <= not a;
    layer1_outputs(1366) <= a and not b;
    layer1_outputs(1367) <= not b;
    layer1_outputs(1368) <= not (a or b);
    layer1_outputs(1369) <= not (a xor b);
    layer1_outputs(1370) <= a xor b;
    layer1_outputs(1371) <= not b or a;
    layer1_outputs(1372) <= not (a xor b);
    layer1_outputs(1373) <= a xor b;
    layer1_outputs(1374) <= not a or b;
    layer1_outputs(1375) <= not b;
    layer1_outputs(1376) <= b;
    layer1_outputs(1377) <= a;
    layer1_outputs(1378) <= '0';
    layer1_outputs(1379) <= not b or a;
    layer1_outputs(1380) <= not a;
    layer1_outputs(1381) <= not b;
    layer1_outputs(1382) <= b and not a;
    layer1_outputs(1383) <= a and not b;
    layer1_outputs(1384) <= not (a or b);
    layer1_outputs(1385) <= a and b;
    layer1_outputs(1386) <= b;
    layer1_outputs(1387) <= not (a or b);
    layer1_outputs(1388) <= a and b;
    layer1_outputs(1389) <= a and b;
    layer1_outputs(1390) <= a;
    layer1_outputs(1391) <= not (a xor b);
    layer1_outputs(1392) <= not b;
    layer1_outputs(1393) <= b;
    layer1_outputs(1394) <= b;
    layer1_outputs(1395) <= a or b;
    layer1_outputs(1396) <= not a;
    layer1_outputs(1397) <= not a;
    layer1_outputs(1398) <= a and b;
    layer1_outputs(1399) <= not b;
    layer1_outputs(1400) <= b and not a;
    layer1_outputs(1401) <= a or b;
    layer1_outputs(1402) <= a and b;
    layer1_outputs(1403) <= not b or a;
    layer1_outputs(1404) <= not a or b;
    layer1_outputs(1405) <= b;
    layer1_outputs(1406) <= a;
    layer1_outputs(1407) <= a and b;
    layer1_outputs(1408) <= b;
    layer1_outputs(1409) <= not a or b;
    layer1_outputs(1410) <= a and b;
    layer1_outputs(1411) <= not a or b;
    layer1_outputs(1412) <= not b or a;
    layer1_outputs(1413) <= a and not b;
    layer1_outputs(1414) <= not b or a;
    layer1_outputs(1415) <= a and not b;
    layer1_outputs(1416) <= a;
    layer1_outputs(1417) <= a xor b;
    layer1_outputs(1418) <= not (a or b);
    layer1_outputs(1419) <= a or b;
    layer1_outputs(1420) <= a or b;
    layer1_outputs(1421) <= a;
    layer1_outputs(1422) <= not b;
    layer1_outputs(1423) <= not b;
    layer1_outputs(1424) <= not a;
    layer1_outputs(1425) <= not a or b;
    layer1_outputs(1426) <= not b or a;
    layer1_outputs(1427) <= a xor b;
    layer1_outputs(1428) <= not (a and b);
    layer1_outputs(1429) <= a;
    layer1_outputs(1430) <= not b or a;
    layer1_outputs(1431) <= not b;
    layer1_outputs(1432) <= a or b;
    layer1_outputs(1433) <= not (a xor b);
    layer1_outputs(1434) <= a or b;
    layer1_outputs(1435) <= a or b;
    layer1_outputs(1436) <= not b or a;
    layer1_outputs(1437) <= a xor b;
    layer1_outputs(1438) <= b;
    layer1_outputs(1439) <= not (a or b);
    layer1_outputs(1440) <= not a;
    layer1_outputs(1441) <= not a;
    layer1_outputs(1442) <= not (a and b);
    layer1_outputs(1443) <= a xor b;
    layer1_outputs(1444) <= a and not b;
    layer1_outputs(1445) <= not (a or b);
    layer1_outputs(1446) <= a and b;
    layer1_outputs(1447) <= not (a and b);
    layer1_outputs(1448) <= a or b;
    layer1_outputs(1449) <= a;
    layer1_outputs(1450) <= a xor b;
    layer1_outputs(1451) <= not b;
    layer1_outputs(1452) <= b and not a;
    layer1_outputs(1453) <= b and not a;
    layer1_outputs(1454) <= not b;
    layer1_outputs(1455) <= a;
    layer1_outputs(1456) <= b;
    layer1_outputs(1457) <= b;
    layer1_outputs(1458) <= b;
    layer1_outputs(1459) <= not b;
    layer1_outputs(1460) <= a;
    layer1_outputs(1461) <= a;
    layer1_outputs(1462) <= a and b;
    layer1_outputs(1463) <= not a or b;
    layer1_outputs(1464) <= a;
    layer1_outputs(1465) <= a or b;
    layer1_outputs(1466) <= not b;
    layer1_outputs(1467) <= a and not b;
    layer1_outputs(1468) <= not a;
    layer1_outputs(1469) <= not b;
    layer1_outputs(1470) <= not a or b;
    layer1_outputs(1471) <= b;
    layer1_outputs(1472) <= not (a or b);
    layer1_outputs(1473) <= not (a or b);
    layer1_outputs(1474) <= not a;
    layer1_outputs(1475) <= not a;
    layer1_outputs(1476) <= not (a and b);
    layer1_outputs(1477) <= not b;
    layer1_outputs(1478) <= a xor b;
    layer1_outputs(1479) <= a and not b;
    layer1_outputs(1480) <= b and not a;
    layer1_outputs(1481) <= a and not b;
    layer1_outputs(1482) <= not (a and b);
    layer1_outputs(1483) <= not a;
    layer1_outputs(1484) <= not (a xor b);
    layer1_outputs(1485) <= not (a or b);
    layer1_outputs(1486) <= not b or a;
    layer1_outputs(1487) <= not (a or b);
    layer1_outputs(1488) <= a or b;
    layer1_outputs(1489) <= a and b;
    layer1_outputs(1490) <= not a;
    layer1_outputs(1491) <= b;
    layer1_outputs(1492) <= a and not b;
    layer1_outputs(1493) <= b;
    layer1_outputs(1494) <= a xor b;
    layer1_outputs(1495) <= not (a or b);
    layer1_outputs(1496) <= not a or b;
    layer1_outputs(1497) <= not b;
    layer1_outputs(1498) <= not b or a;
    layer1_outputs(1499) <= b;
    layer1_outputs(1500) <= a xor b;
    layer1_outputs(1501) <= a;
    layer1_outputs(1502) <= a;
    layer1_outputs(1503) <= not (a xor b);
    layer1_outputs(1504) <= not (a or b);
    layer1_outputs(1505) <= not (a or b);
    layer1_outputs(1506) <= not (a xor b);
    layer1_outputs(1507) <= not a;
    layer1_outputs(1508) <= a and b;
    layer1_outputs(1509) <= b;
    layer1_outputs(1510) <= b;
    layer1_outputs(1511) <= not (a xor b);
    layer1_outputs(1512) <= b;
    layer1_outputs(1513) <= b and not a;
    layer1_outputs(1514) <= not a;
    layer1_outputs(1515) <= not b;
    layer1_outputs(1516) <= not (a and b);
    layer1_outputs(1517) <= not a or b;
    layer1_outputs(1518) <= not a or b;
    layer1_outputs(1519) <= not (a or b);
    layer1_outputs(1520) <= b;
    layer1_outputs(1521) <= a and not b;
    layer1_outputs(1522) <= not (a xor b);
    layer1_outputs(1523) <= not (a xor b);
    layer1_outputs(1524) <= a and b;
    layer1_outputs(1525) <= not a;
    layer1_outputs(1526) <= not (a xor b);
    layer1_outputs(1527) <= not a;
    layer1_outputs(1528) <= not a;
    layer1_outputs(1529) <= not b or a;
    layer1_outputs(1530) <= not (a and b);
    layer1_outputs(1531) <= not (a xor b);
    layer1_outputs(1532) <= '1';
    layer1_outputs(1533) <= a or b;
    layer1_outputs(1534) <= a;
    layer1_outputs(1535) <= a or b;
    layer1_outputs(1536) <= a or b;
    layer1_outputs(1537) <= not b or a;
    layer1_outputs(1538) <= not b;
    layer1_outputs(1539) <= not a;
    layer1_outputs(1540) <= not b;
    layer1_outputs(1541) <= a and not b;
    layer1_outputs(1542) <= '0';
    layer1_outputs(1543) <= not b;
    layer1_outputs(1544) <= a or b;
    layer1_outputs(1545) <= not b;
    layer1_outputs(1546) <= not (a and b);
    layer1_outputs(1547) <= not (a and b);
    layer1_outputs(1548) <= a xor b;
    layer1_outputs(1549) <= not (a and b);
    layer1_outputs(1550) <= b;
    layer1_outputs(1551) <= b;
    layer1_outputs(1552) <= not (a xor b);
    layer1_outputs(1553) <= a xor b;
    layer1_outputs(1554) <= '0';
    layer1_outputs(1555) <= b;
    layer1_outputs(1556) <= not b or a;
    layer1_outputs(1557) <= a xor b;
    layer1_outputs(1558) <= a or b;
    layer1_outputs(1559) <= a;
    layer1_outputs(1560) <= not (a xor b);
    layer1_outputs(1561) <= not b;
    layer1_outputs(1562) <= b and not a;
    layer1_outputs(1563) <= not b;
    layer1_outputs(1564) <= a;
    layer1_outputs(1565) <= not a;
    layer1_outputs(1566) <= a or b;
    layer1_outputs(1567) <= not a or b;
    layer1_outputs(1568) <= not (a or b);
    layer1_outputs(1569) <= a;
    layer1_outputs(1570) <= a xor b;
    layer1_outputs(1571) <= a;
    layer1_outputs(1572) <= b;
    layer1_outputs(1573) <= b;
    layer1_outputs(1574) <= not a or b;
    layer1_outputs(1575) <= a or b;
    layer1_outputs(1576) <= not b or a;
    layer1_outputs(1577) <= b;
    layer1_outputs(1578) <= not (a xor b);
    layer1_outputs(1579) <= not b;
    layer1_outputs(1580) <= a xor b;
    layer1_outputs(1581) <= a and not b;
    layer1_outputs(1582) <= not a or b;
    layer1_outputs(1583) <= '1';
    layer1_outputs(1584) <= b;
    layer1_outputs(1585) <= a and not b;
    layer1_outputs(1586) <= not a or b;
    layer1_outputs(1587) <= '1';
    layer1_outputs(1588) <= not b;
    layer1_outputs(1589) <= b and not a;
    layer1_outputs(1590) <= not (a or b);
    layer1_outputs(1591) <= not (a and b);
    layer1_outputs(1592) <= not a or b;
    layer1_outputs(1593) <= a and not b;
    layer1_outputs(1594) <= not b;
    layer1_outputs(1595) <= not a or b;
    layer1_outputs(1596) <= a and not b;
    layer1_outputs(1597) <= b;
    layer1_outputs(1598) <= not (a xor b);
    layer1_outputs(1599) <= a and not b;
    layer1_outputs(1600) <= a xor b;
    layer1_outputs(1601) <= not (a or b);
    layer1_outputs(1602) <= b;
    layer1_outputs(1603) <= not (a xor b);
    layer1_outputs(1604) <= a and b;
    layer1_outputs(1605) <= not a or b;
    layer1_outputs(1606) <= not b;
    layer1_outputs(1607) <= not a;
    layer1_outputs(1608) <= a xor b;
    layer1_outputs(1609) <= a and b;
    layer1_outputs(1610) <= not (a or b);
    layer1_outputs(1611) <= a;
    layer1_outputs(1612) <= a xor b;
    layer1_outputs(1613) <= a or b;
    layer1_outputs(1614) <= b;
    layer1_outputs(1615) <= not a or b;
    layer1_outputs(1616) <= b;
    layer1_outputs(1617) <= not b;
    layer1_outputs(1618) <= not a;
    layer1_outputs(1619) <= a and b;
    layer1_outputs(1620) <= a or b;
    layer1_outputs(1621) <= not b;
    layer1_outputs(1622) <= not a;
    layer1_outputs(1623) <= not (a or b);
    layer1_outputs(1624) <= not b;
    layer1_outputs(1625) <= a and not b;
    layer1_outputs(1626) <= a and not b;
    layer1_outputs(1627) <= not (a and b);
    layer1_outputs(1628) <= a;
    layer1_outputs(1629) <= not a or b;
    layer1_outputs(1630) <= a;
    layer1_outputs(1631) <= not b or a;
    layer1_outputs(1632) <= b;
    layer1_outputs(1633) <= b and not a;
    layer1_outputs(1634) <= a and b;
    layer1_outputs(1635) <= not a or b;
    layer1_outputs(1636) <= not (a xor b);
    layer1_outputs(1637) <= a and not b;
    layer1_outputs(1638) <= b and not a;
    layer1_outputs(1639) <= not a;
    layer1_outputs(1640) <= not (a and b);
    layer1_outputs(1641) <= not (a xor b);
    layer1_outputs(1642) <= a or b;
    layer1_outputs(1643) <= not a;
    layer1_outputs(1644) <= not (a or b);
    layer1_outputs(1645) <= a and not b;
    layer1_outputs(1646) <= not b;
    layer1_outputs(1647) <= b;
    layer1_outputs(1648) <= not b;
    layer1_outputs(1649) <= not (a xor b);
    layer1_outputs(1650) <= not (a or b);
    layer1_outputs(1651) <= '1';
    layer1_outputs(1652) <= not b or a;
    layer1_outputs(1653) <= a and b;
    layer1_outputs(1654) <= not a;
    layer1_outputs(1655) <= not a;
    layer1_outputs(1656) <= a xor b;
    layer1_outputs(1657) <= b and not a;
    layer1_outputs(1658) <= b and not a;
    layer1_outputs(1659) <= b;
    layer1_outputs(1660) <= not (a and b);
    layer1_outputs(1661) <= not b;
    layer1_outputs(1662) <= not a or b;
    layer1_outputs(1663) <= not b or a;
    layer1_outputs(1664) <= not a or b;
    layer1_outputs(1665) <= a xor b;
    layer1_outputs(1666) <= a or b;
    layer1_outputs(1667) <= b and not a;
    layer1_outputs(1668) <= a and b;
    layer1_outputs(1669) <= not b;
    layer1_outputs(1670) <= a or b;
    layer1_outputs(1671) <= a or b;
    layer1_outputs(1672) <= a xor b;
    layer1_outputs(1673) <= a or b;
    layer1_outputs(1674) <= not b or a;
    layer1_outputs(1675) <= b;
    layer1_outputs(1676) <= not b;
    layer1_outputs(1677) <= b;
    layer1_outputs(1678) <= not b;
    layer1_outputs(1679) <= b;
    layer1_outputs(1680) <= b;
    layer1_outputs(1681) <= a and not b;
    layer1_outputs(1682) <= a and not b;
    layer1_outputs(1683) <= not a;
    layer1_outputs(1684) <= not (a xor b);
    layer1_outputs(1685) <= not b;
    layer1_outputs(1686) <= b;
    layer1_outputs(1687) <= a and b;
    layer1_outputs(1688) <= not b or a;
    layer1_outputs(1689) <= not (a and b);
    layer1_outputs(1690) <= not a or b;
    layer1_outputs(1691) <= not (a and b);
    layer1_outputs(1692) <= not (a and b);
    layer1_outputs(1693) <= a;
    layer1_outputs(1694) <= not (a xor b);
    layer1_outputs(1695) <= not b or a;
    layer1_outputs(1696) <= not b;
    layer1_outputs(1697) <= a and b;
    layer1_outputs(1698) <= not b;
    layer1_outputs(1699) <= a xor b;
    layer1_outputs(1700) <= a and not b;
    layer1_outputs(1701) <= not b;
    layer1_outputs(1702) <= b;
    layer1_outputs(1703) <= b;
    layer1_outputs(1704) <= not (a xor b);
    layer1_outputs(1705) <= not a or b;
    layer1_outputs(1706) <= not a or b;
    layer1_outputs(1707) <= not b;
    layer1_outputs(1708) <= a and not b;
    layer1_outputs(1709) <= b and not a;
    layer1_outputs(1710) <= b;
    layer1_outputs(1711) <= not a;
    layer1_outputs(1712) <= not b;
    layer1_outputs(1713) <= a xor b;
    layer1_outputs(1714) <= not b;
    layer1_outputs(1715) <= not (a and b);
    layer1_outputs(1716) <= a and b;
    layer1_outputs(1717) <= a or b;
    layer1_outputs(1718) <= not (a and b);
    layer1_outputs(1719) <= '0';
    layer1_outputs(1720) <= b and not a;
    layer1_outputs(1721) <= not (a and b);
    layer1_outputs(1722) <= a;
    layer1_outputs(1723) <= not (a xor b);
    layer1_outputs(1724) <= not b;
    layer1_outputs(1725) <= not b or a;
    layer1_outputs(1726) <= not b;
    layer1_outputs(1727) <= a;
    layer1_outputs(1728) <= a xor b;
    layer1_outputs(1729) <= a or b;
    layer1_outputs(1730) <= not a;
    layer1_outputs(1731) <= a xor b;
    layer1_outputs(1732) <= not (a or b);
    layer1_outputs(1733) <= a and b;
    layer1_outputs(1734) <= '0';
    layer1_outputs(1735) <= not a or b;
    layer1_outputs(1736) <= a and not b;
    layer1_outputs(1737) <= a xor b;
    layer1_outputs(1738) <= not b or a;
    layer1_outputs(1739) <= not (a or b);
    layer1_outputs(1740) <= b;
    layer1_outputs(1741) <= b;
    layer1_outputs(1742) <= b;
    layer1_outputs(1743) <= a xor b;
    layer1_outputs(1744) <= b and not a;
    layer1_outputs(1745) <= b and not a;
    layer1_outputs(1746) <= not a;
    layer1_outputs(1747) <= not b;
    layer1_outputs(1748) <= b;
    layer1_outputs(1749) <= b;
    layer1_outputs(1750) <= b and not a;
    layer1_outputs(1751) <= a and b;
    layer1_outputs(1752) <= a or b;
    layer1_outputs(1753) <= not (a or b);
    layer1_outputs(1754) <= a xor b;
    layer1_outputs(1755) <= a xor b;
    layer1_outputs(1756) <= a and not b;
    layer1_outputs(1757) <= '0';
    layer1_outputs(1758) <= not b;
    layer1_outputs(1759) <= not (a xor b);
    layer1_outputs(1760) <= not a or b;
    layer1_outputs(1761) <= a or b;
    layer1_outputs(1762) <= a xor b;
    layer1_outputs(1763) <= a;
    layer1_outputs(1764) <= not (a and b);
    layer1_outputs(1765) <= a and b;
    layer1_outputs(1766) <= not b;
    layer1_outputs(1767) <= not (a or b);
    layer1_outputs(1768) <= '0';
    layer1_outputs(1769) <= a;
    layer1_outputs(1770) <= b;
    layer1_outputs(1771) <= a xor b;
    layer1_outputs(1772) <= b and not a;
    layer1_outputs(1773) <= a;
    layer1_outputs(1774) <= not a;
    layer1_outputs(1775) <= not (a or b);
    layer1_outputs(1776) <= not a or b;
    layer1_outputs(1777) <= b;
    layer1_outputs(1778) <= not b;
    layer1_outputs(1779) <= not (a and b);
    layer1_outputs(1780) <= a or b;
    layer1_outputs(1781) <= a xor b;
    layer1_outputs(1782) <= a or b;
    layer1_outputs(1783) <= b and not a;
    layer1_outputs(1784) <= a and b;
    layer1_outputs(1785) <= a;
    layer1_outputs(1786) <= a xor b;
    layer1_outputs(1787) <= not a;
    layer1_outputs(1788) <= a;
    layer1_outputs(1789) <= a;
    layer1_outputs(1790) <= b;
    layer1_outputs(1791) <= not (a or b);
    layer1_outputs(1792) <= a and b;
    layer1_outputs(1793) <= a and not b;
    layer1_outputs(1794) <= '1';
    layer1_outputs(1795) <= a xor b;
    layer1_outputs(1796) <= not a;
    layer1_outputs(1797) <= a and b;
    layer1_outputs(1798) <= not b or a;
    layer1_outputs(1799) <= not (a xor b);
    layer1_outputs(1800) <= a;
    layer1_outputs(1801) <= b and not a;
    layer1_outputs(1802) <= not a or b;
    layer1_outputs(1803) <= a xor b;
    layer1_outputs(1804) <= a;
    layer1_outputs(1805) <= a;
    layer1_outputs(1806) <= a and b;
    layer1_outputs(1807) <= not (a and b);
    layer1_outputs(1808) <= not b or a;
    layer1_outputs(1809) <= b and not a;
    layer1_outputs(1810) <= not (a or b);
    layer1_outputs(1811) <= a or b;
    layer1_outputs(1812) <= not (a and b);
    layer1_outputs(1813) <= not b;
    layer1_outputs(1814) <= a;
    layer1_outputs(1815) <= a and not b;
    layer1_outputs(1816) <= a or b;
    layer1_outputs(1817) <= b;
    layer1_outputs(1818) <= a and b;
    layer1_outputs(1819) <= b;
    layer1_outputs(1820) <= not a;
    layer1_outputs(1821) <= a;
    layer1_outputs(1822) <= not b or a;
    layer1_outputs(1823) <= a and not b;
    layer1_outputs(1824) <= not a;
    layer1_outputs(1825) <= a xor b;
    layer1_outputs(1826) <= a xor b;
    layer1_outputs(1827) <= not a;
    layer1_outputs(1828) <= not (a or b);
    layer1_outputs(1829) <= not b or a;
    layer1_outputs(1830) <= a or b;
    layer1_outputs(1831) <= b;
    layer1_outputs(1832) <= a and b;
    layer1_outputs(1833) <= a and b;
    layer1_outputs(1834) <= not b or a;
    layer1_outputs(1835) <= a or b;
    layer1_outputs(1836) <= not (a and b);
    layer1_outputs(1837) <= '0';
    layer1_outputs(1838) <= a;
    layer1_outputs(1839) <= a;
    layer1_outputs(1840) <= a and b;
    layer1_outputs(1841) <= not a;
    layer1_outputs(1842) <= b and not a;
    layer1_outputs(1843) <= not (a or b);
    layer1_outputs(1844) <= not b;
    layer1_outputs(1845) <= a or b;
    layer1_outputs(1846) <= a xor b;
    layer1_outputs(1847) <= a and not b;
    layer1_outputs(1848) <= not a;
    layer1_outputs(1849) <= not (a xor b);
    layer1_outputs(1850) <= not (a xor b);
    layer1_outputs(1851) <= not a or b;
    layer1_outputs(1852) <= not a or b;
    layer1_outputs(1853) <= '1';
    layer1_outputs(1854) <= a;
    layer1_outputs(1855) <= not (a xor b);
    layer1_outputs(1856) <= a or b;
    layer1_outputs(1857) <= a;
    layer1_outputs(1858) <= a and not b;
    layer1_outputs(1859) <= a or b;
    layer1_outputs(1860) <= not b;
    layer1_outputs(1861) <= not (a xor b);
    layer1_outputs(1862) <= a;
    layer1_outputs(1863) <= b and not a;
    layer1_outputs(1864) <= a and not b;
    layer1_outputs(1865) <= '1';
    layer1_outputs(1866) <= a or b;
    layer1_outputs(1867) <= a xor b;
    layer1_outputs(1868) <= not a;
    layer1_outputs(1869) <= not (a and b);
    layer1_outputs(1870) <= a;
    layer1_outputs(1871) <= not b;
    layer1_outputs(1872) <= not a;
    layer1_outputs(1873) <= a xor b;
    layer1_outputs(1874) <= not (a xor b);
    layer1_outputs(1875) <= b;
    layer1_outputs(1876) <= a xor b;
    layer1_outputs(1877) <= not a;
    layer1_outputs(1878) <= a or b;
    layer1_outputs(1879) <= not (a and b);
    layer1_outputs(1880) <= not b or a;
    layer1_outputs(1881) <= a and b;
    layer1_outputs(1882) <= not b or a;
    layer1_outputs(1883) <= not (a or b);
    layer1_outputs(1884) <= not (a xor b);
    layer1_outputs(1885) <= not b or a;
    layer1_outputs(1886) <= b;
    layer1_outputs(1887) <= b and not a;
    layer1_outputs(1888) <= a or b;
    layer1_outputs(1889) <= a xor b;
    layer1_outputs(1890) <= a and b;
    layer1_outputs(1891) <= a;
    layer1_outputs(1892) <= a xor b;
    layer1_outputs(1893) <= not (a xor b);
    layer1_outputs(1894) <= not (a and b);
    layer1_outputs(1895) <= a;
    layer1_outputs(1896) <= '0';
    layer1_outputs(1897) <= b and not a;
    layer1_outputs(1898) <= not (a and b);
    layer1_outputs(1899) <= not b;
    layer1_outputs(1900) <= b;
    layer1_outputs(1901) <= not b or a;
    layer1_outputs(1902) <= not (a or b);
    layer1_outputs(1903) <= not (a and b);
    layer1_outputs(1904) <= b;
    layer1_outputs(1905) <= a;
    layer1_outputs(1906) <= not (a and b);
    layer1_outputs(1907) <= not a or b;
    layer1_outputs(1908) <= a;
    layer1_outputs(1909) <= b;
    layer1_outputs(1910) <= not (a and b);
    layer1_outputs(1911) <= a xor b;
    layer1_outputs(1912) <= not b;
    layer1_outputs(1913) <= b;
    layer1_outputs(1914) <= not (a and b);
    layer1_outputs(1915) <= b;
    layer1_outputs(1916) <= a;
    layer1_outputs(1917) <= a;
    layer1_outputs(1918) <= not a or b;
    layer1_outputs(1919) <= a or b;
    layer1_outputs(1920) <= not b;
    layer1_outputs(1921) <= a or b;
    layer1_outputs(1922) <= a or b;
    layer1_outputs(1923) <= a xor b;
    layer1_outputs(1924) <= not a or b;
    layer1_outputs(1925) <= not (a xor b);
    layer1_outputs(1926) <= not a;
    layer1_outputs(1927) <= not b;
    layer1_outputs(1928) <= a or b;
    layer1_outputs(1929) <= not a;
    layer1_outputs(1930) <= not (a xor b);
    layer1_outputs(1931) <= not (a and b);
    layer1_outputs(1932) <= not b;
    layer1_outputs(1933) <= not (a xor b);
    layer1_outputs(1934) <= a and not b;
    layer1_outputs(1935) <= a and b;
    layer1_outputs(1936) <= b;
    layer1_outputs(1937) <= not b;
    layer1_outputs(1938) <= not b or a;
    layer1_outputs(1939) <= a and b;
    layer1_outputs(1940) <= b;
    layer1_outputs(1941) <= a xor b;
    layer1_outputs(1942) <= not a or b;
    layer1_outputs(1943) <= not (a or b);
    layer1_outputs(1944) <= not b;
    layer1_outputs(1945) <= b;
    layer1_outputs(1946) <= not b;
    layer1_outputs(1947) <= a;
    layer1_outputs(1948) <= a;
    layer1_outputs(1949) <= b and not a;
    layer1_outputs(1950) <= b and not a;
    layer1_outputs(1951) <= a and b;
    layer1_outputs(1952) <= not (a and b);
    layer1_outputs(1953) <= not b;
    layer1_outputs(1954) <= a;
    layer1_outputs(1955) <= not (a or b);
    layer1_outputs(1956) <= b;
    layer1_outputs(1957) <= b;
    layer1_outputs(1958) <= a;
    layer1_outputs(1959) <= not a;
    layer1_outputs(1960) <= not a;
    layer1_outputs(1961) <= a or b;
    layer1_outputs(1962) <= a and b;
    layer1_outputs(1963) <= not b;
    layer1_outputs(1964) <= a and not b;
    layer1_outputs(1965) <= a or b;
    layer1_outputs(1966) <= not (a xor b);
    layer1_outputs(1967) <= b and not a;
    layer1_outputs(1968) <= not (a and b);
    layer1_outputs(1969) <= b and not a;
    layer1_outputs(1970) <= not b or a;
    layer1_outputs(1971) <= not (a xor b);
    layer1_outputs(1972) <= b;
    layer1_outputs(1973) <= b and not a;
    layer1_outputs(1974) <= not (a and b);
    layer1_outputs(1975) <= not (a xor b);
    layer1_outputs(1976) <= a or b;
    layer1_outputs(1977) <= not b;
    layer1_outputs(1978) <= '0';
    layer1_outputs(1979) <= not (a and b);
    layer1_outputs(1980) <= not (a or b);
    layer1_outputs(1981) <= not b;
    layer1_outputs(1982) <= not (a xor b);
    layer1_outputs(1983) <= not (a or b);
    layer1_outputs(1984) <= a;
    layer1_outputs(1985) <= b and not a;
    layer1_outputs(1986) <= a;
    layer1_outputs(1987) <= not b;
    layer1_outputs(1988) <= a and b;
    layer1_outputs(1989) <= a xor b;
    layer1_outputs(1990) <= a and b;
    layer1_outputs(1991) <= a xor b;
    layer1_outputs(1992) <= not b or a;
    layer1_outputs(1993) <= not b or a;
    layer1_outputs(1994) <= not b;
    layer1_outputs(1995) <= b;
    layer1_outputs(1996) <= not (a and b);
    layer1_outputs(1997) <= a or b;
    layer1_outputs(1998) <= b;
    layer1_outputs(1999) <= b;
    layer1_outputs(2000) <= not b or a;
    layer1_outputs(2001) <= b and not a;
    layer1_outputs(2002) <= not a;
    layer1_outputs(2003) <= not (a and b);
    layer1_outputs(2004) <= a or b;
    layer1_outputs(2005) <= a and b;
    layer1_outputs(2006) <= a;
    layer1_outputs(2007) <= not (a xor b);
    layer1_outputs(2008) <= not b or a;
    layer1_outputs(2009) <= not b;
    layer1_outputs(2010) <= not b or a;
    layer1_outputs(2011) <= not (a and b);
    layer1_outputs(2012) <= a;
    layer1_outputs(2013) <= a or b;
    layer1_outputs(2014) <= b and not a;
    layer1_outputs(2015) <= not (a or b);
    layer1_outputs(2016) <= a;
    layer1_outputs(2017) <= not b;
    layer1_outputs(2018) <= a or b;
    layer1_outputs(2019) <= a;
    layer1_outputs(2020) <= not b;
    layer1_outputs(2021) <= not b or a;
    layer1_outputs(2022) <= not a;
    layer1_outputs(2023) <= not (a xor b);
    layer1_outputs(2024) <= not (a or b);
    layer1_outputs(2025) <= b;
    layer1_outputs(2026) <= not b;
    layer1_outputs(2027) <= a or b;
    layer1_outputs(2028) <= not a;
    layer1_outputs(2029) <= a;
    layer1_outputs(2030) <= not a;
    layer1_outputs(2031) <= a;
    layer1_outputs(2032) <= not (a or b);
    layer1_outputs(2033) <= a and b;
    layer1_outputs(2034) <= b;
    layer1_outputs(2035) <= b;
    layer1_outputs(2036) <= not a or b;
    layer1_outputs(2037) <= a or b;
    layer1_outputs(2038) <= not (a or b);
    layer1_outputs(2039) <= a xor b;
    layer1_outputs(2040) <= not (a xor b);
    layer1_outputs(2041) <= not (a and b);
    layer1_outputs(2042) <= b and not a;
    layer1_outputs(2043) <= a or b;
    layer1_outputs(2044) <= not a or b;
    layer1_outputs(2045) <= a and b;
    layer1_outputs(2046) <= not (a xor b);
    layer1_outputs(2047) <= a and not b;
    layer1_outputs(2048) <= not (a and b);
    layer1_outputs(2049) <= a xor b;
    layer1_outputs(2050) <= a and not b;
    layer1_outputs(2051) <= not a;
    layer1_outputs(2052) <= not (a and b);
    layer1_outputs(2053) <= a;
    layer1_outputs(2054) <= a or b;
    layer1_outputs(2055) <= a;
    layer1_outputs(2056) <= not a or b;
    layer1_outputs(2057) <= not b;
    layer1_outputs(2058) <= not b or a;
    layer1_outputs(2059) <= a and not b;
    layer1_outputs(2060) <= not a;
    layer1_outputs(2061) <= a and not b;
    layer1_outputs(2062) <= a or b;
    layer1_outputs(2063) <= not (a xor b);
    layer1_outputs(2064) <= not a;
    layer1_outputs(2065) <= a xor b;
    layer1_outputs(2066) <= not (a or b);
    layer1_outputs(2067) <= a and not b;
    layer1_outputs(2068) <= not a or b;
    layer1_outputs(2069) <= a and b;
    layer1_outputs(2070) <= not a or b;
    layer1_outputs(2071) <= not a or b;
    layer1_outputs(2072) <= not (a xor b);
    layer1_outputs(2073) <= a;
    layer1_outputs(2074) <= not a or b;
    layer1_outputs(2075) <= not (a or b);
    layer1_outputs(2076) <= '1';
    layer1_outputs(2077) <= not (a and b);
    layer1_outputs(2078) <= a and b;
    layer1_outputs(2079) <= b;
    layer1_outputs(2080) <= a;
    layer1_outputs(2081) <= a or b;
    layer1_outputs(2082) <= b and not a;
    layer1_outputs(2083) <= b and not a;
    layer1_outputs(2084) <= a or b;
    layer1_outputs(2085) <= not a or b;
    layer1_outputs(2086) <= b;
    layer1_outputs(2087) <= a xor b;
    layer1_outputs(2088) <= not (a xor b);
    layer1_outputs(2089) <= a;
    layer1_outputs(2090) <= a and b;
    layer1_outputs(2091) <= a;
    layer1_outputs(2092) <= not a;
    layer1_outputs(2093) <= not (a or b);
    layer1_outputs(2094) <= not (a or b);
    layer1_outputs(2095) <= b and not a;
    layer1_outputs(2096) <= a and not b;
    layer1_outputs(2097) <= a;
    layer1_outputs(2098) <= not (a and b);
    layer1_outputs(2099) <= a and b;
    layer1_outputs(2100) <= not (a xor b);
    layer1_outputs(2101) <= b;
    layer1_outputs(2102) <= a and b;
    layer1_outputs(2103) <= not (a xor b);
    layer1_outputs(2104) <= not a;
    layer1_outputs(2105) <= not (a xor b);
    layer1_outputs(2106) <= not a;
    layer1_outputs(2107) <= a xor b;
    layer1_outputs(2108) <= not (a and b);
    layer1_outputs(2109) <= a;
    layer1_outputs(2110) <= not a;
    layer1_outputs(2111) <= a;
    layer1_outputs(2112) <= a and b;
    layer1_outputs(2113) <= not b or a;
    layer1_outputs(2114) <= not (a and b);
    layer1_outputs(2115) <= not a;
    layer1_outputs(2116) <= not a;
    layer1_outputs(2117) <= not a or b;
    layer1_outputs(2118) <= not b;
    layer1_outputs(2119) <= not a;
    layer1_outputs(2120) <= b;
    layer1_outputs(2121) <= not (a and b);
    layer1_outputs(2122) <= not (a or b);
    layer1_outputs(2123) <= not (a and b);
    layer1_outputs(2124) <= not b or a;
    layer1_outputs(2125) <= not a;
    layer1_outputs(2126) <= not a;
    layer1_outputs(2127) <= b;
    layer1_outputs(2128) <= a;
    layer1_outputs(2129) <= b;
    layer1_outputs(2130) <= not a or b;
    layer1_outputs(2131) <= a;
    layer1_outputs(2132) <= not a or b;
    layer1_outputs(2133) <= not (a or b);
    layer1_outputs(2134) <= not (a xor b);
    layer1_outputs(2135) <= a and not b;
    layer1_outputs(2136) <= a and b;
    layer1_outputs(2137) <= not (a xor b);
    layer1_outputs(2138) <= a;
    layer1_outputs(2139) <= not b or a;
    layer1_outputs(2140) <= a xor b;
    layer1_outputs(2141) <= not (a and b);
    layer1_outputs(2142) <= a;
    layer1_outputs(2143) <= b;
    layer1_outputs(2144) <= not a or b;
    layer1_outputs(2145) <= a or b;
    layer1_outputs(2146) <= not (a xor b);
    layer1_outputs(2147) <= not (a or b);
    layer1_outputs(2148) <= a and b;
    layer1_outputs(2149) <= not b;
    layer1_outputs(2150) <= not b;
    layer1_outputs(2151) <= a and b;
    layer1_outputs(2152) <= a and b;
    layer1_outputs(2153) <= a or b;
    layer1_outputs(2154) <= a xor b;
    layer1_outputs(2155) <= a;
    layer1_outputs(2156) <= not (a or b);
    layer1_outputs(2157) <= not b or a;
    layer1_outputs(2158) <= b;
    layer1_outputs(2159) <= a;
    layer1_outputs(2160) <= a or b;
    layer1_outputs(2161) <= not a;
    layer1_outputs(2162) <= not (a xor b);
    layer1_outputs(2163) <= not b;
    layer1_outputs(2164) <= not b;
    layer1_outputs(2165) <= not (a and b);
    layer1_outputs(2166) <= not a;
    layer1_outputs(2167) <= not a or b;
    layer1_outputs(2168) <= a and b;
    layer1_outputs(2169) <= not (a xor b);
    layer1_outputs(2170) <= a;
    layer1_outputs(2171) <= a or b;
    layer1_outputs(2172) <= a;
    layer1_outputs(2173) <= a xor b;
    layer1_outputs(2174) <= a;
    layer1_outputs(2175) <= not (a or b);
    layer1_outputs(2176) <= not a;
    layer1_outputs(2177) <= a and b;
    layer1_outputs(2178) <= not (a xor b);
    layer1_outputs(2179) <= b;
    layer1_outputs(2180) <= a xor b;
    layer1_outputs(2181) <= not a or b;
    layer1_outputs(2182) <= b;
    layer1_outputs(2183) <= not a or b;
    layer1_outputs(2184) <= a and b;
    layer1_outputs(2185) <= not a or b;
    layer1_outputs(2186) <= not a;
    layer1_outputs(2187) <= not (a xor b);
    layer1_outputs(2188) <= not b or a;
    layer1_outputs(2189) <= a xor b;
    layer1_outputs(2190) <= not b or a;
    layer1_outputs(2191) <= not b or a;
    layer1_outputs(2192) <= not b;
    layer1_outputs(2193) <= a and b;
    layer1_outputs(2194) <= a and b;
    layer1_outputs(2195) <= not b;
    layer1_outputs(2196) <= b;
    layer1_outputs(2197) <= a;
    layer1_outputs(2198) <= not (a or b);
    layer1_outputs(2199) <= not b or a;
    layer1_outputs(2200) <= not b;
    layer1_outputs(2201) <= b;
    layer1_outputs(2202) <= b and not a;
    layer1_outputs(2203) <= a;
    layer1_outputs(2204) <= not b or a;
    layer1_outputs(2205) <= a;
    layer1_outputs(2206) <= a xor b;
    layer1_outputs(2207) <= a and not b;
    layer1_outputs(2208) <= not (a xor b);
    layer1_outputs(2209) <= a;
    layer1_outputs(2210) <= not (a or b);
    layer1_outputs(2211) <= a;
    layer1_outputs(2212) <= not b or a;
    layer1_outputs(2213) <= not a;
    layer1_outputs(2214) <= a and not b;
    layer1_outputs(2215) <= a;
    layer1_outputs(2216) <= b;
    layer1_outputs(2217) <= b and not a;
    layer1_outputs(2218) <= a;
    layer1_outputs(2219) <= a xor b;
    layer1_outputs(2220) <= not (a or b);
    layer1_outputs(2221) <= not (a and b);
    layer1_outputs(2222) <= not a;
    layer1_outputs(2223) <= not a;
    layer1_outputs(2224) <= not a;
    layer1_outputs(2225) <= not b or a;
    layer1_outputs(2226) <= not (a and b);
    layer1_outputs(2227) <= b;
    layer1_outputs(2228) <= a xor b;
    layer1_outputs(2229) <= a;
    layer1_outputs(2230) <= not a;
    layer1_outputs(2231) <= not (a or b);
    layer1_outputs(2232) <= not b;
    layer1_outputs(2233) <= b;
    layer1_outputs(2234) <= not b;
    layer1_outputs(2235) <= not a or b;
    layer1_outputs(2236) <= not (a or b);
    layer1_outputs(2237) <= a and b;
    layer1_outputs(2238) <= a or b;
    layer1_outputs(2239) <= not (a or b);
    layer1_outputs(2240) <= not (a xor b);
    layer1_outputs(2241) <= not (a or b);
    layer1_outputs(2242) <= a;
    layer1_outputs(2243) <= not (a and b);
    layer1_outputs(2244) <= not a;
    layer1_outputs(2245) <= a xor b;
    layer1_outputs(2246) <= not (a or b);
    layer1_outputs(2247) <= a or b;
    layer1_outputs(2248) <= b and not a;
    layer1_outputs(2249) <= not (a or b);
    layer1_outputs(2250) <= not (a xor b);
    layer1_outputs(2251) <= not (a xor b);
    layer1_outputs(2252) <= a xor b;
    layer1_outputs(2253) <= not (a and b);
    layer1_outputs(2254) <= a and not b;
    layer1_outputs(2255) <= not b;
    layer1_outputs(2256) <= a;
    layer1_outputs(2257) <= b and not a;
    layer1_outputs(2258) <= not b;
    layer1_outputs(2259) <= b and not a;
    layer1_outputs(2260) <= not a;
    layer1_outputs(2261) <= not b or a;
    layer1_outputs(2262) <= not b or a;
    layer1_outputs(2263) <= not a or b;
    layer1_outputs(2264) <= a xor b;
    layer1_outputs(2265) <= not (a xor b);
    layer1_outputs(2266) <= not (a or b);
    layer1_outputs(2267) <= a;
    layer1_outputs(2268) <= a and not b;
    layer1_outputs(2269) <= not a;
    layer1_outputs(2270) <= b;
    layer1_outputs(2271) <= not b;
    layer1_outputs(2272) <= b;
    layer1_outputs(2273) <= b;
    layer1_outputs(2274) <= a and b;
    layer1_outputs(2275) <= a;
    layer1_outputs(2276) <= not (a xor b);
    layer1_outputs(2277) <= '1';
    layer1_outputs(2278) <= not b;
    layer1_outputs(2279) <= a;
    layer1_outputs(2280) <= a;
    layer1_outputs(2281) <= not (a xor b);
    layer1_outputs(2282) <= a and b;
    layer1_outputs(2283) <= a xor b;
    layer1_outputs(2284) <= a or b;
    layer1_outputs(2285) <= not b;
    layer1_outputs(2286) <= a or b;
    layer1_outputs(2287) <= b and not a;
    layer1_outputs(2288) <= '1';
    layer1_outputs(2289) <= not b;
    layer1_outputs(2290) <= not (a or b);
    layer1_outputs(2291) <= a and b;
    layer1_outputs(2292) <= not (a or b);
    layer1_outputs(2293) <= not (a xor b);
    layer1_outputs(2294) <= a;
    layer1_outputs(2295) <= not b;
    layer1_outputs(2296) <= not (a xor b);
    layer1_outputs(2297) <= b;
    layer1_outputs(2298) <= b and not a;
    layer1_outputs(2299) <= a;
    layer1_outputs(2300) <= not (a xor b);
    layer1_outputs(2301) <= b and not a;
    layer1_outputs(2302) <= b and not a;
    layer1_outputs(2303) <= not (a or b);
    layer1_outputs(2304) <= a and not b;
    layer1_outputs(2305) <= not a;
    layer1_outputs(2306) <= not (a and b);
    layer1_outputs(2307) <= not b;
    layer1_outputs(2308) <= a xor b;
    layer1_outputs(2309) <= a or b;
    layer1_outputs(2310) <= not a or b;
    layer1_outputs(2311) <= b and not a;
    layer1_outputs(2312) <= not a;
    layer1_outputs(2313) <= a xor b;
    layer1_outputs(2314) <= a and not b;
    layer1_outputs(2315) <= a xor b;
    layer1_outputs(2316) <= not (a or b);
    layer1_outputs(2317) <= a;
    layer1_outputs(2318) <= a or b;
    layer1_outputs(2319) <= not (a and b);
    layer1_outputs(2320) <= a and not b;
    layer1_outputs(2321) <= not a or b;
    layer1_outputs(2322) <= not a or b;
    layer1_outputs(2323) <= not b or a;
    layer1_outputs(2324) <= not a or b;
    layer1_outputs(2325) <= b;
    layer1_outputs(2326) <= a or b;
    layer1_outputs(2327) <= a xor b;
    layer1_outputs(2328) <= b;
    layer1_outputs(2329) <= b;
    layer1_outputs(2330) <= b;
    layer1_outputs(2331) <= not (a or b);
    layer1_outputs(2332) <= a and not b;
    layer1_outputs(2333) <= '1';
    layer1_outputs(2334) <= not a;
    layer1_outputs(2335) <= not b;
    layer1_outputs(2336) <= not a;
    layer1_outputs(2337) <= a or b;
    layer1_outputs(2338) <= a xor b;
    layer1_outputs(2339) <= not (a or b);
    layer1_outputs(2340) <= not b;
    layer1_outputs(2341) <= not a;
    layer1_outputs(2342) <= not a;
    layer1_outputs(2343) <= '1';
    layer1_outputs(2344) <= a and not b;
    layer1_outputs(2345) <= not b;
    layer1_outputs(2346) <= b and not a;
    layer1_outputs(2347) <= a or b;
    layer1_outputs(2348) <= a;
    layer1_outputs(2349) <= a xor b;
    layer1_outputs(2350) <= not b or a;
    layer1_outputs(2351) <= a and b;
    layer1_outputs(2352) <= not (a or b);
    layer1_outputs(2353) <= a;
    layer1_outputs(2354) <= a and b;
    layer1_outputs(2355) <= not b or a;
    layer1_outputs(2356) <= a and not b;
    layer1_outputs(2357) <= not (a or b);
    layer1_outputs(2358) <= not (a xor b);
    layer1_outputs(2359) <= not a;
    layer1_outputs(2360) <= not a;
    layer1_outputs(2361) <= not b;
    layer1_outputs(2362) <= not a;
    layer1_outputs(2363) <= a and b;
    layer1_outputs(2364) <= '0';
    layer1_outputs(2365) <= not a;
    layer1_outputs(2366) <= b and not a;
    layer1_outputs(2367) <= not (a or b);
    layer1_outputs(2368) <= not (a or b);
    layer1_outputs(2369) <= a and b;
    layer1_outputs(2370) <= not b;
    layer1_outputs(2371) <= a and not b;
    layer1_outputs(2372) <= not (a or b);
    layer1_outputs(2373) <= not (a and b);
    layer1_outputs(2374) <= a xor b;
    layer1_outputs(2375) <= not a;
    layer1_outputs(2376) <= not (a and b);
    layer1_outputs(2377) <= not (a or b);
    layer1_outputs(2378) <= a and b;
    layer1_outputs(2379) <= '0';
    layer1_outputs(2380) <= a and b;
    layer1_outputs(2381) <= a and b;
    layer1_outputs(2382) <= '1';
    layer1_outputs(2383) <= not (a or b);
    layer1_outputs(2384) <= a;
    layer1_outputs(2385) <= b;
    layer1_outputs(2386) <= a and b;
    layer1_outputs(2387) <= a;
    layer1_outputs(2388) <= a and not b;
    layer1_outputs(2389) <= not a;
    layer1_outputs(2390) <= a and not b;
    layer1_outputs(2391) <= not (a xor b);
    layer1_outputs(2392) <= not b;
    layer1_outputs(2393) <= a and not b;
    layer1_outputs(2394) <= a xor b;
    layer1_outputs(2395) <= a and b;
    layer1_outputs(2396) <= a and not b;
    layer1_outputs(2397) <= a xor b;
    layer1_outputs(2398) <= a and not b;
    layer1_outputs(2399) <= a and not b;
    layer1_outputs(2400) <= b and not a;
    layer1_outputs(2401) <= not (a and b);
    layer1_outputs(2402) <= not (a or b);
    layer1_outputs(2403) <= not (a or b);
    layer1_outputs(2404) <= b and not a;
    layer1_outputs(2405) <= not a;
    layer1_outputs(2406) <= a and not b;
    layer1_outputs(2407) <= not (a xor b);
    layer1_outputs(2408) <= b;
    layer1_outputs(2409) <= b and not a;
    layer1_outputs(2410) <= b;
    layer1_outputs(2411) <= a or b;
    layer1_outputs(2412) <= not a;
    layer1_outputs(2413) <= not (a xor b);
    layer1_outputs(2414) <= not b or a;
    layer1_outputs(2415) <= not a or b;
    layer1_outputs(2416) <= a;
    layer1_outputs(2417) <= not a;
    layer1_outputs(2418) <= not b;
    layer1_outputs(2419) <= b and not a;
    layer1_outputs(2420) <= '0';
    layer1_outputs(2421) <= b;
    layer1_outputs(2422) <= a and not b;
    layer1_outputs(2423) <= b;
    layer1_outputs(2424) <= a xor b;
    layer1_outputs(2425) <= not a;
    layer1_outputs(2426) <= a and not b;
    layer1_outputs(2427) <= a;
    layer1_outputs(2428) <= not b or a;
    layer1_outputs(2429) <= not (a xor b);
    layer1_outputs(2430) <= a xor b;
    layer1_outputs(2431) <= not (a or b);
    layer1_outputs(2432) <= b;
    layer1_outputs(2433) <= a xor b;
    layer1_outputs(2434) <= not b;
    layer1_outputs(2435) <= b;
    layer1_outputs(2436) <= a xor b;
    layer1_outputs(2437) <= a or b;
    layer1_outputs(2438) <= not b;
    layer1_outputs(2439) <= a and not b;
    layer1_outputs(2440) <= a and not b;
    layer1_outputs(2441) <= a or b;
    layer1_outputs(2442) <= b;
    layer1_outputs(2443) <= not b or a;
    layer1_outputs(2444) <= not (a and b);
    layer1_outputs(2445) <= b;
    layer1_outputs(2446) <= a and b;
    layer1_outputs(2447) <= a or b;
    layer1_outputs(2448) <= a and b;
    layer1_outputs(2449) <= b;
    layer1_outputs(2450) <= b and not a;
    layer1_outputs(2451) <= not (a or b);
    layer1_outputs(2452) <= '0';
    layer1_outputs(2453) <= a and not b;
    layer1_outputs(2454) <= a;
    layer1_outputs(2455) <= not a or b;
    layer1_outputs(2456) <= not b;
    layer1_outputs(2457) <= b;
    layer1_outputs(2458) <= a or b;
    layer1_outputs(2459) <= not (a or b);
    layer1_outputs(2460) <= not (a or b);
    layer1_outputs(2461) <= not b;
    layer1_outputs(2462) <= not (a xor b);
    layer1_outputs(2463) <= a;
    layer1_outputs(2464) <= not (a or b);
    layer1_outputs(2465) <= a;
    layer1_outputs(2466) <= a and b;
    layer1_outputs(2467) <= a xor b;
    layer1_outputs(2468) <= not b or a;
    layer1_outputs(2469) <= not (a xor b);
    layer1_outputs(2470) <= not b;
    layer1_outputs(2471) <= a;
    layer1_outputs(2472) <= not b or a;
    layer1_outputs(2473) <= not b or a;
    layer1_outputs(2474) <= not (a and b);
    layer1_outputs(2475) <= a and b;
    layer1_outputs(2476) <= a xor b;
    layer1_outputs(2477) <= b;
    layer1_outputs(2478) <= a xor b;
    layer1_outputs(2479) <= not b or a;
    layer1_outputs(2480) <= not (a or b);
    layer1_outputs(2481) <= b and not a;
    layer1_outputs(2482) <= a xor b;
    layer1_outputs(2483) <= not a or b;
    layer1_outputs(2484) <= not a or b;
    layer1_outputs(2485) <= a and b;
    layer1_outputs(2486) <= a and not b;
    layer1_outputs(2487) <= a xor b;
    layer1_outputs(2488) <= a;
    layer1_outputs(2489) <= not b;
    layer1_outputs(2490) <= not (a and b);
    layer1_outputs(2491) <= a and b;
    layer1_outputs(2492) <= not a;
    layer1_outputs(2493) <= a or b;
    layer1_outputs(2494) <= a and not b;
    layer1_outputs(2495) <= not b;
    layer1_outputs(2496) <= a;
    layer1_outputs(2497) <= not a;
    layer1_outputs(2498) <= a;
    layer1_outputs(2499) <= not b;
    layer1_outputs(2500) <= not a;
    layer1_outputs(2501) <= a xor b;
    layer1_outputs(2502) <= a;
    layer1_outputs(2503) <= b and not a;
    layer1_outputs(2504) <= not b or a;
    layer1_outputs(2505) <= not a;
    layer1_outputs(2506) <= not a;
    layer1_outputs(2507) <= a;
    layer1_outputs(2508) <= not b;
    layer1_outputs(2509) <= b;
    layer1_outputs(2510) <= a;
    layer1_outputs(2511) <= not (a and b);
    layer1_outputs(2512) <= not a or b;
    layer1_outputs(2513) <= a or b;
    layer1_outputs(2514) <= not (a xor b);
    layer1_outputs(2515) <= '1';
    layer1_outputs(2516) <= b and not a;
    layer1_outputs(2517) <= b and not a;
    layer1_outputs(2518) <= not (a xor b);
    layer1_outputs(2519) <= a or b;
    layer1_outputs(2520) <= not b;
    layer1_outputs(2521) <= not (a and b);
    layer1_outputs(2522) <= a and b;
    layer1_outputs(2523) <= b;
    layer1_outputs(2524) <= a;
    layer1_outputs(2525) <= b and not a;
    layer1_outputs(2526) <= a and b;
    layer1_outputs(2527) <= not a;
    layer1_outputs(2528) <= a and b;
    layer1_outputs(2529) <= not b;
    layer1_outputs(2530) <= a or b;
    layer1_outputs(2531) <= a and not b;
    layer1_outputs(2532) <= not (a and b);
    layer1_outputs(2533) <= a or b;
    layer1_outputs(2534) <= not (a and b);
    layer1_outputs(2535) <= not a;
    layer1_outputs(2536) <= a or b;
    layer1_outputs(2537) <= '0';
    layer1_outputs(2538) <= a and b;
    layer1_outputs(2539) <= not b;
    layer1_outputs(2540) <= not a;
    layer1_outputs(2541) <= a;
    layer1_outputs(2542) <= b and not a;
    layer1_outputs(2543) <= not b;
    layer1_outputs(2544) <= not b;
    layer1_outputs(2545) <= a xor b;
    layer1_outputs(2546) <= not b or a;
    layer1_outputs(2547) <= a and not b;
    layer1_outputs(2548) <= not b;
    layer1_outputs(2549) <= a or b;
    layer1_outputs(2550) <= b and not a;
    layer1_outputs(2551) <= b and not a;
    layer1_outputs(2552) <= a;
    layer1_outputs(2553) <= b;
    layer1_outputs(2554) <= not a or b;
    layer1_outputs(2555) <= b;
    layer1_outputs(2556) <= not (a and b);
    layer1_outputs(2557) <= not (a and b);
    layer1_outputs(2558) <= not (a or b);
    layer1_outputs(2559) <= not a or b;
    layer1_outputs(2560) <= not b;
    layer1_outputs(2561) <= a;
    layer1_outputs(2562) <= a xor b;
    layer1_outputs(2563) <= a xor b;
    layer1_outputs(2564) <= not (a or b);
    layer1_outputs(2565) <= a and b;
    layer1_outputs(2566) <= a and not b;
    layer1_outputs(2567) <= a and not b;
    layer1_outputs(2568) <= not a;
    layer1_outputs(2569) <= not (a and b);
    layer1_outputs(2570) <= not a;
    layer1_outputs(2571) <= a and not b;
    layer1_outputs(2572) <= not a;
    layer1_outputs(2573) <= a or b;
    layer1_outputs(2574) <= not b;
    layer1_outputs(2575) <= b and not a;
    layer1_outputs(2576) <= not b;
    layer1_outputs(2577) <= not (a and b);
    layer1_outputs(2578) <= not b;
    layer1_outputs(2579) <= not a;
    layer1_outputs(2580) <= not (a or b);
    layer1_outputs(2581) <= not b;
    layer1_outputs(2582) <= a;
    layer1_outputs(2583) <= not (a or b);
    layer1_outputs(2584) <= not a;
    layer1_outputs(2585) <= b and not a;
    layer1_outputs(2586) <= b;
    layer1_outputs(2587) <= not a;
    layer1_outputs(2588) <= b and not a;
    layer1_outputs(2589) <= a;
    layer1_outputs(2590) <= a or b;
    layer1_outputs(2591) <= not b;
    layer1_outputs(2592) <= not b;
    layer1_outputs(2593) <= not (a xor b);
    layer1_outputs(2594) <= not a or b;
    layer1_outputs(2595) <= b and not a;
    layer1_outputs(2596) <= a or b;
    layer1_outputs(2597) <= not b;
    layer1_outputs(2598) <= not (a xor b);
    layer1_outputs(2599) <= a or b;
    layer1_outputs(2600) <= not (a xor b);
    layer1_outputs(2601) <= '0';
    layer1_outputs(2602) <= not (a and b);
    layer1_outputs(2603) <= b and not a;
    layer1_outputs(2604) <= a and not b;
    layer1_outputs(2605) <= not b or a;
    layer1_outputs(2606) <= a;
    layer1_outputs(2607) <= not a or b;
    layer1_outputs(2608) <= a xor b;
    layer1_outputs(2609) <= not (a xor b);
    layer1_outputs(2610) <= a xor b;
    layer1_outputs(2611) <= not (a xor b);
    layer1_outputs(2612) <= a and b;
    layer1_outputs(2613) <= not a;
    layer1_outputs(2614) <= '0';
    layer1_outputs(2615) <= a xor b;
    layer1_outputs(2616) <= not b or a;
    layer1_outputs(2617) <= not (a xor b);
    layer1_outputs(2618) <= not a;
    layer1_outputs(2619) <= not (a or b);
    layer1_outputs(2620) <= b;
    layer1_outputs(2621) <= a or b;
    layer1_outputs(2622) <= a xor b;
    layer1_outputs(2623) <= not a;
    layer1_outputs(2624) <= a;
    layer1_outputs(2625) <= not b;
    layer1_outputs(2626) <= not b;
    layer1_outputs(2627) <= a or b;
    layer1_outputs(2628) <= a xor b;
    layer1_outputs(2629) <= not a or b;
    layer1_outputs(2630) <= not b;
    layer1_outputs(2631) <= a and b;
    layer1_outputs(2632) <= not b or a;
    layer1_outputs(2633) <= a and b;
    layer1_outputs(2634) <= a xor b;
    layer1_outputs(2635) <= not b or a;
    layer1_outputs(2636) <= a;
    layer1_outputs(2637) <= a;
    layer1_outputs(2638) <= not (a xor b);
    layer1_outputs(2639) <= not b or a;
    layer1_outputs(2640) <= a and not b;
    layer1_outputs(2641) <= a;
    layer1_outputs(2642) <= not a;
    layer1_outputs(2643) <= a xor b;
    layer1_outputs(2644) <= a xor b;
    layer1_outputs(2645) <= not a or b;
    layer1_outputs(2646) <= b and not a;
    layer1_outputs(2647) <= not (a and b);
    layer1_outputs(2648) <= a or b;
    layer1_outputs(2649) <= not a or b;
    layer1_outputs(2650) <= not a;
    layer1_outputs(2651) <= b;
    layer1_outputs(2652) <= not b;
    layer1_outputs(2653) <= not b or a;
    layer1_outputs(2654) <= not (a or b);
    layer1_outputs(2655) <= not a;
    layer1_outputs(2656) <= b;
    layer1_outputs(2657) <= b;
    layer1_outputs(2658) <= a xor b;
    layer1_outputs(2659) <= not (a xor b);
    layer1_outputs(2660) <= not (a or b);
    layer1_outputs(2661) <= a and not b;
    layer1_outputs(2662) <= a or b;
    layer1_outputs(2663) <= a and b;
    layer1_outputs(2664) <= not a or b;
    layer1_outputs(2665) <= not (a and b);
    layer1_outputs(2666) <= not b;
    layer1_outputs(2667) <= not a or b;
    layer1_outputs(2668) <= a and not b;
    layer1_outputs(2669) <= not b or a;
    layer1_outputs(2670) <= a or b;
    layer1_outputs(2671) <= not b or a;
    layer1_outputs(2672) <= not b;
    layer1_outputs(2673) <= a and b;
    layer1_outputs(2674) <= b and not a;
    layer1_outputs(2675) <= a and b;
    layer1_outputs(2676) <= not (a or b);
    layer1_outputs(2677) <= not (a and b);
    layer1_outputs(2678) <= not b;
    layer1_outputs(2679) <= not b;
    layer1_outputs(2680) <= a;
    layer1_outputs(2681) <= not (a and b);
    layer1_outputs(2682) <= b;
    layer1_outputs(2683) <= not b or a;
    layer1_outputs(2684) <= not (a and b);
    layer1_outputs(2685) <= not b;
    layer1_outputs(2686) <= b;
    layer1_outputs(2687) <= '1';
    layer1_outputs(2688) <= a xor b;
    layer1_outputs(2689) <= a or b;
    layer1_outputs(2690) <= not b;
    layer1_outputs(2691) <= b and not a;
    layer1_outputs(2692) <= not (a xor b);
    layer1_outputs(2693) <= not b;
    layer1_outputs(2694) <= a or b;
    layer1_outputs(2695) <= a;
    layer1_outputs(2696) <= b;
    layer1_outputs(2697) <= a and b;
    layer1_outputs(2698) <= a xor b;
    layer1_outputs(2699) <= b and not a;
    layer1_outputs(2700) <= not a;
    layer1_outputs(2701) <= a and b;
    layer1_outputs(2702) <= not (a xor b);
    layer1_outputs(2703) <= not (a or b);
    layer1_outputs(2704) <= a and b;
    layer1_outputs(2705) <= not b;
    layer1_outputs(2706) <= a;
    layer1_outputs(2707) <= b and not a;
    layer1_outputs(2708) <= not b;
    layer1_outputs(2709) <= b and not a;
    layer1_outputs(2710) <= not (a xor b);
    layer1_outputs(2711) <= not a or b;
    layer1_outputs(2712) <= not b;
    layer1_outputs(2713) <= a;
    layer1_outputs(2714) <= b;
    layer1_outputs(2715) <= a;
    layer1_outputs(2716) <= b;
    layer1_outputs(2717) <= not b or a;
    layer1_outputs(2718) <= not (a or b);
    layer1_outputs(2719) <= not b;
    layer1_outputs(2720) <= a xor b;
    layer1_outputs(2721) <= a and not b;
    layer1_outputs(2722) <= not (a or b);
    layer1_outputs(2723) <= not b;
    layer1_outputs(2724) <= not a;
    layer1_outputs(2725) <= not (a xor b);
    layer1_outputs(2726) <= not (a xor b);
    layer1_outputs(2727) <= not (a xor b);
    layer1_outputs(2728) <= not a or b;
    layer1_outputs(2729) <= not (a xor b);
    layer1_outputs(2730) <= not a;
    layer1_outputs(2731) <= a xor b;
    layer1_outputs(2732) <= a;
    layer1_outputs(2733) <= b and not a;
    layer1_outputs(2734) <= not b or a;
    layer1_outputs(2735) <= not b or a;
    layer1_outputs(2736) <= a or b;
    layer1_outputs(2737) <= not (a xor b);
    layer1_outputs(2738) <= '1';
    layer1_outputs(2739) <= not a or b;
    layer1_outputs(2740) <= b;
    layer1_outputs(2741) <= not b;
    layer1_outputs(2742) <= not a;
    layer1_outputs(2743) <= not (a xor b);
    layer1_outputs(2744) <= not b;
    layer1_outputs(2745) <= not (a xor b);
    layer1_outputs(2746) <= not (a or b);
    layer1_outputs(2747) <= not a;
    layer1_outputs(2748) <= not b;
    layer1_outputs(2749) <= a;
    layer1_outputs(2750) <= b and not a;
    layer1_outputs(2751) <= not b;
    layer1_outputs(2752) <= a;
    layer1_outputs(2753) <= not a;
    layer1_outputs(2754) <= not (a and b);
    layer1_outputs(2755) <= a;
    layer1_outputs(2756) <= a xor b;
    layer1_outputs(2757) <= '1';
    layer1_outputs(2758) <= a or b;
    layer1_outputs(2759) <= a and b;
    layer1_outputs(2760) <= not a or b;
    layer1_outputs(2761) <= not b or a;
    layer1_outputs(2762) <= not b or a;
    layer1_outputs(2763) <= a;
    layer1_outputs(2764) <= not a or b;
    layer1_outputs(2765) <= a or b;
    layer1_outputs(2766) <= a xor b;
    layer1_outputs(2767) <= not a;
    layer1_outputs(2768) <= a;
    layer1_outputs(2769) <= a and not b;
    layer1_outputs(2770) <= not (a or b);
    layer1_outputs(2771) <= a;
    layer1_outputs(2772) <= not (a or b);
    layer1_outputs(2773) <= not (a and b);
    layer1_outputs(2774) <= not a;
    layer1_outputs(2775) <= '0';
    layer1_outputs(2776) <= not (a or b);
    layer1_outputs(2777) <= a and not b;
    layer1_outputs(2778) <= not b;
    layer1_outputs(2779) <= not (a xor b);
    layer1_outputs(2780) <= not a;
    layer1_outputs(2781) <= a and b;
    layer1_outputs(2782) <= b;
    layer1_outputs(2783) <= b;
    layer1_outputs(2784) <= b;
    layer1_outputs(2785) <= a or b;
    layer1_outputs(2786) <= not (a xor b);
    layer1_outputs(2787) <= not (a and b);
    layer1_outputs(2788) <= not a or b;
    layer1_outputs(2789) <= b;
    layer1_outputs(2790) <= a or b;
    layer1_outputs(2791) <= not a;
    layer1_outputs(2792) <= not a;
    layer1_outputs(2793) <= not b;
    layer1_outputs(2794) <= not (a xor b);
    layer1_outputs(2795) <= not a;
    layer1_outputs(2796) <= not (a and b);
    layer1_outputs(2797) <= not (a xor b);
    layer1_outputs(2798) <= not (a xor b);
    layer1_outputs(2799) <= not b or a;
    layer1_outputs(2800) <= not (a xor b);
    layer1_outputs(2801) <= b;
    layer1_outputs(2802) <= b and not a;
    layer1_outputs(2803) <= b;
    layer1_outputs(2804) <= not (a xor b);
    layer1_outputs(2805) <= not b or a;
    layer1_outputs(2806) <= b and not a;
    layer1_outputs(2807) <= not (a xor b);
    layer1_outputs(2808) <= b;
    layer1_outputs(2809) <= a and not b;
    layer1_outputs(2810) <= a xor b;
    layer1_outputs(2811) <= b;
    layer1_outputs(2812) <= b and not a;
    layer1_outputs(2813) <= not (a or b);
    layer1_outputs(2814) <= b and not a;
    layer1_outputs(2815) <= b;
    layer1_outputs(2816) <= not a or b;
    layer1_outputs(2817) <= not b or a;
    layer1_outputs(2818) <= not (a xor b);
    layer1_outputs(2819) <= b and not a;
    layer1_outputs(2820) <= b;
    layer1_outputs(2821) <= a and b;
    layer1_outputs(2822) <= a;
    layer1_outputs(2823) <= not a;
    layer1_outputs(2824) <= b;
    layer1_outputs(2825) <= '1';
    layer1_outputs(2826) <= not b;
    layer1_outputs(2827) <= a;
    layer1_outputs(2828) <= not (a xor b);
    layer1_outputs(2829) <= b;
    layer1_outputs(2830) <= not a;
    layer1_outputs(2831) <= b;
    layer1_outputs(2832) <= b;
    layer1_outputs(2833) <= not b or a;
    layer1_outputs(2834) <= a and not b;
    layer1_outputs(2835) <= a or b;
    layer1_outputs(2836) <= not b;
    layer1_outputs(2837) <= not (a and b);
    layer1_outputs(2838) <= b;
    layer1_outputs(2839) <= not b;
    layer1_outputs(2840) <= not (a xor b);
    layer1_outputs(2841) <= not a or b;
    layer1_outputs(2842) <= a and b;
    layer1_outputs(2843) <= a;
    layer1_outputs(2844) <= a and not b;
    layer1_outputs(2845) <= '1';
    layer1_outputs(2846) <= a or b;
    layer1_outputs(2847) <= not b;
    layer1_outputs(2848) <= not a;
    layer1_outputs(2849) <= not b;
    layer1_outputs(2850) <= not (a and b);
    layer1_outputs(2851) <= not b;
    layer1_outputs(2852) <= a xor b;
    layer1_outputs(2853) <= '0';
    layer1_outputs(2854) <= b and not a;
    layer1_outputs(2855) <= a xor b;
    layer1_outputs(2856) <= a;
    layer1_outputs(2857) <= not (a and b);
    layer1_outputs(2858) <= '0';
    layer1_outputs(2859) <= a;
    layer1_outputs(2860) <= a;
    layer1_outputs(2861) <= not b or a;
    layer1_outputs(2862) <= not a;
    layer1_outputs(2863) <= not b or a;
    layer1_outputs(2864) <= not b or a;
    layer1_outputs(2865) <= a and not b;
    layer1_outputs(2866) <= not b;
    layer1_outputs(2867) <= b and not a;
    layer1_outputs(2868) <= a;
    layer1_outputs(2869) <= b and not a;
    layer1_outputs(2870) <= a and b;
    layer1_outputs(2871) <= a and b;
    layer1_outputs(2872) <= a or b;
    layer1_outputs(2873) <= not a or b;
    layer1_outputs(2874) <= a xor b;
    layer1_outputs(2875) <= not a or b;
    layer1_outputs(2876) <= b;
    layer1_outputs(2877) <= not (a or b);
    layer1_outputs(2878) <= not a;
    layer1_outputs(2879) <= not (a and b);
    layer1_outputs(2880) <= not a or b;
    layer1_outputs(2881) <= not b or a;
    layer1_outputs(2882) <= a and not b;
    layer1_outputs(2883) <= not b;
    layer1_outputs(2884) <= not (a or b);
    layer1_outputs(2885) <= a xor b;
    layer1_outputs(2886) <= not (a xor b);
    layer1_outputs(2887) <= b;
    layer1_outputs(2888) <= not b;
    layer1_outputs(2889) <= not a;
    layer1_outputs(2890) <= b;
    layer1_outputs(2891) <= not (a xor b);
    layer1_outputs(2892) <= a xor b;
    layer1_outputs(2893) <= not b or a;
    layer1_outputs(2894) <= not b;
    layer1_outputs(2895) <= a and not b;
    layer1_outputs(2896) <= not a or b;
    layer1_outputs(2897) <= a xor b;
    layer1_outputs(2898) <= a;
    layer1_outputs(2899) <= a;
    layer1_outputs(2900) <= not (a or b);
    layer1_outputs(2901) <= a;
    layer1_outputs(2902) <= not b;
    layer1_outputs(2903) <= '1';
    layer1_outputs(2904) <= not b or a;
    layer1_outputs(2905) <= not (a xor b);
    layer1_outputs(2906) <= not b or a;
    layer1_outputs(2907) <= not (a and b);
    layer1_outputs(2908) <= b;
    layer1_outputs(2909) <= not b;
    layer1_outputs(2910) <= not a;
    layer1_outputs(2911) <= a xor b;
    layer1_outputs(2912) <= a xor b;
    layer1_outputs(2913) <= b;
    layer1_outputs(2914) <= a;
    layer1_outputs(2915) <= a and b;
    layer1_outputs(2916) <= b and not a;
    layer1_outputs(2917) <= not a or b;
    layer1_outputs(2918) <= a;
    layer1_outputs(2919) <= not (a and b);
    layer1_outputs(2920) <= not a;
    layer1_outputs(2921) <= a and not b;
    layer1_outputs(2922) <= a xor b;
    layer1_outputs(2923) <= not (a xor b);
    layer1_outputs(2924) <= a and not b;
    layer1_outputs(2925) <= a xor b;
    layer1_outputs(2926) <= a and b;
    layer1_outputs(2927) <= not a or b;
    layer1_outputs(2928) <= b and not a;
    layer1_outputs(2929) <= a;
    layer1_outputs(2930) <= not (a xor b);
    layer1_outputs(2931) <= b;
    layer1_outputs(2932) <= a or b;
    layer1_outputs(2933) <= '1';
    layer1_outputs(2934) <= b and not a;
    layer1_outputs(2935) <= not a;
    layer1_outputs(2936) <= b;
    layer1_outputs(2937) <= a;
    layer1_outputs(2938) <= a or b;
    layer1_outputs(2939) <= a;
    layer1_outputs(2940) <= not (a xor b);
    layer1_outputs(2941) <= not a or b;
    layer1_outputs(2942) <= not (a xor b);
    layer1_outputs(2943) <= a and b;
    layer1_outputs(2944) <= not a or b;
    layer1_outputs(2945) <= not a;
    layer1_outputs(2946) <= a and b;
    layer1_outputs(2947) <= b and not a;
    layer1_outputs(2948) <= not b;
    layer1_outputs(2949) <= not b or a;
    layer1_outputs(2950) <= a or b;
    layer1_outputs(2951) <= a and b;
    layer1_outputs(2952) <= a or b;
    layer1_outputs(2953) <= a;
    layer1_outputs(2954) <= a or b;
    layer1_outputs(2955) <= not (a or b);
    layer1_outputs(2956) <= a xor b;
    layer1_outputs(2957) <= a;
    layer1_outputs(2958) <= a;
    layer1_outputs(2959) <= b;
    layer1_outputs(2960) <= not (a and b);
    layer1_outputs(2961) <= a and not b;
    layer1_outputs(2962) <= not (a xor b);
    layer1_outputs(2963) <= a xor b;
    layer1_outputs(2964) <= not (a or b);
    layer1_outputs(2965) <= a xor b;
    layer1_outputs(2966) <= b and not a;
    layer1_outputs(2967) <= not (a and b);
    layer1_outputs(2968) <= a and b;
    layer1_outputs(2969) <= a and b;
    layer1_outputs(2970) <= b;
    layer1_outputs(2971) <= not a or b;
    layer1_outputs(2972) <= not b;
    layer1_outputs(2973) <= a;
    layer1_outputs(2974) <= not b;
    layer1_outputs(2975) <= not b or a;
    layer1_outputs(2976) <= not (a and b);
    layer1_outputs(2977) <= a xor b;
    layer1_outputs(2978) <= not a or b;
    layer1_outputs(2979) <= not (a and b);
    layer1_outputs(2980) <= not a;
    layer1_outputs(2981) <= b;
    layer1_outputs(2982) <= a xor b;
    layer1_outputs(2983) <= a or b;
    layer1_outputs(2984) <= a and b;
    layer1_outputs(2985) <= not a;
    layer1_outputs(2986) <= not b or a;
    layer1_outputs(2987) <= not a;
    layer1_outputs(2988) <= not a;
    layer1_outputs(2989) <= not (a xor b);
    layer1_outputs(2990) <= not (a or b);
    layer1_outputs(2991) <= b;
    layer1_outputs(2992) <= not a;
    layer1_outputs(2993) <= b;
    layer1_outputs(2994) <= '0';
    layer1_outputs(2995) <= a xor b;
    layer1_outputs(2996) <= a xor b;
    layer1_outputs(2997) <= a xor b;
    layer1_outputs(2998) <= not a or b;
    layer1_outputs(2999) <= a;
    layer1_outputs(3000) <= b and not a;
    layer1_outputs(3001) <= a xor b;
    layer1_outputs(3002) <= a xor b;
    layer1_outputs(3003) <= a or b;
    layer1_outputs(3004) <= not (a and b);
    layer1_outputs(3005) <= a and not b;
    layer1_outputs(3006) <= a and not b;
    layer1_outputs(3007) <= not b;
    layer1_outputs(3008) <= b;
    layer1_outputs(3009) <= a and not b;
    layer1_outputs(3010) <= not a;
    layer1_outputs(3011) <= not b or a;
    layer1_outputs(3012) <= a and not b;
    layer1_outputs(3013) <= not (a and b);
    layer1_outputs(3014) <= not (a xor b);
    layer1_outputs(3015) <= not (a or b);
    layer1_outputs(3016) <= not (a and b);
    layer1_outputs(3017) <= not a or b;
    layer1_outputs(3018) <= not a;
    layer1_outputs(3019) <= a xor b;
    layer1_outputs(3020) <= b;
    layer1_outputs(3021) <= b and not a;
    layer1_outputs(3022) <= a;
    layer1_outputs(3023) <= not (a xor b);
    layer1_outputs(3024) <= not (a xor b);
    layer1_outputs(3025) <= not a or b;
    layer1_outputs(3026) <= b;
    layer1_outputs(3027) <= not a;
    layer1_outputs(3028) <= not (a or b);
    layer1_outputs(3029) <= not (a xor b);
    layer1_outputs(3030) <= not a;
    layer1_outputs(3031) <= not (a xor b);
    layer1_outputs(3032) <= a;
    layer1_outputs(3033) <= not (a or b);
    layer1_outputs(3034) <= a and b;
    layer1_outputs(3035) <= not b;
    layer1_outputs(3036) <= a;
    layer1_outputs(3037) <= not a or b;
    layer1_outputs(3038) <= not a;
    layer1_outputs(3039) <= a xor b;
    layer1_outputs(3040) <= not b or a;
    layer1_outputs(3041) <= not (a xor b);
    layer1_outputs(3042) <= a or b;
    layer1_outputs(3043) <= b;
    layer1_outputs(3044) <= a;
    layer1_outputs(3045) <= a;
    layer1_outputs(3046) <= a and b;
    layer1_outputs(3047) <= b;
    layer1_outputs(3048) <= not (a or b);
    layer1_outputs(3049) <= a;
    layer1_outputs(3050) <= not a or b;
    layer1_outputs(3051) <= not (a and b);
    layer1_outputs(3052) <= a and not b;
    layer1_outputs(3053) <= a and b;
    layer1_outputs(3054) <= '1';
    layer1_outputs(3055) <= not a;
    layer1_outputs(3056) <= a;
    layer1_outputs(3057) <= not a or b;
    layer1_outputs(3058) <= b;
    layer1_outputs(3059) <= not b or a;
    layer1_outputs(3060) <= not (a or b);
    layer1_outputs(3061) <= a xor b;
    layer1_outputs(3062) <= not a;
    layer1_outputs(3063) <= not (a and b);
    layer1_outputs(3064) <= not b or a;
    layer1_outputs(3065) <= not a or b;
    layer1_outputs(3066) <= not a;
    layer1_outputs(3067) <= a and b;
    layer1_outputs(3068) <= not (a xor b);
    layer1_outputs(3069) <= a and b;
    layer1_outputs(3070) <= a and not b;
    layer1_outputs(3071) <= a and b;
    layer1_outputs(3072) <= b and not a;
    layer1_outputs(3073) <= a xor b;
    layer1_outputs(3074) <= not b;
    layer1_outputs(3075) <= not b or a;
    layer1_outputs(3076) <= not (a xor b);
    layer1_outputs(3077) <= a and not b;
    layer1_outputs(3078) <= not b or a;
    layer1_outputs(3079) <= not (a or b);
    layer1_outputs(3080) <= a;
    layer1_outputs(3081) <= not b;
    layer1_outputs(3082) <= not b or a;
    layer1_outputs(3083) <= not b;
    layer1_outputs(3084) <= not (a and b);
    layer1_outputs(3085) <= '0';
    layer1_outputs(3086) <= not b;
    layer1_outputs(3087) <= '0';
    layer1_outputs(3088) <= a and b;
    layer1_outputs(3089) <= not b;
    layer1_outputs(3090) <= not b;
    layer1_outputs(3091) <= a and b;
    layer1_outputs(3092) <= a or b;
    layer1_outputs(3093) <= not a or b;
    layer1_outputs(3094) <= a or b;
    layer1_outputs(3095) <= a or b;
    layer1_outputs(3096) <= not a;
    layer1_outputs(3097) <= not a or b;
    layer1_outputs(3098) <= a or b;
    layer1_outputs(3099) <= not b;
    layer1_outputs(3100) <= not a;
    layer1_outputs(3101) <= '1';
    layer1_outputs(3102) <= b;
    layer1_outputs(3103) <= '1';
    layer1_outputs(3104) <= b;
    layer1_outputs(3105) <= not (a xor b);
    layer1_outputs(3106) <= not a;
    layer1_outputs(3107) <= a and not b;
    layer1_outputs(3108) <= not (a or b);
    layer1_outputs(3109) <= not (a or b);
    layer1_outputs(3110) <= not b;
    layer1_outputs(3111) <= not (a or b);
    layer1_outputs(3112) <= b;
    layer1_outputs(3113) <= a and b;
    layer1_outputs(3114) <= a or b;
    layer1_outputs(3115) <= b;
    layer1_outputs(3116) <= b and not a;
    layer1_outputs(3117) <= not (a and b);
    layer1_outputs(3118) <= a and not b;
    layer1_outputs(3119) <= '0';
    layer1_outputs(3120) <= a;
    layer1_outputs(3121) <= a or b;
    layer1_outputs(3122) <= a;
    layer1_outputs(3123) <= not a;
    layer1_outputs(3124) <= a and b;
    layer1_outputs(3125) <= a;
    layer1_outputs(3126) <= a;
    layer1_outputs(3127) <= a;
    layer1_outputs(3128) <= a and not b;
    layer1_outputs(3129) <= not (a xor b);
    layer1_outputs(3130) <= not a;
    layer1_outputs(3131) <= not (a xor b);
    layer1_outputs(3132) <= a;
    layer1_outputs(3133) <= not (a or b);
    layer1_outputs(3134) <= not (a or b);
    layer1_outputs(3135) <= not (a or b);
    layer1_outputs(3136) <= b;
    layer1_outputs(3137) <= a xor b;
    layer1_outputs(3138) <= not b;
    layer1_outputs(3139) <= a or b;
    layer1_outputs(3140) <= not a or b;
    layer1_outputs(3141) <= not b;
    layer1_outputs(3142) <= a xor b;
    layer1_outputs(3143) <= not b;
    layer1_outputs(3144) <= a xor b;
    layer1_outputs(3145) <= not (a or b);
    layer1_outputs(3146) <= not a or b;
    layer1_outputs(3147) <= not b;
    layer1_outputs(3148) <= not (a xor b);
    layer1_outputs(3149) <= not b;
    layer1_outputs(3150) <= not a or b;
    layer1_outputs(3151) <= a xor b;
    layer1_outputs(3152) <= not a;
    layer1_outputs(3153) <= b;
    layer1_outputs(3154) <= not a;
    layer1_outputs(3155) <= a;
    layer1_outputs(3156) <= not (a xor b);
    layer1_outputs(3157) <= not a or b;
    layer1_outputs(3158) <= a and not b;
    layer1_outputs(3159) <= a xor b;
    layer1_outputs(3160) <= a xor b;
    layer1_outputs(3161) <= a or b;
    layer1_outputs(3162) <= not b or a;
    layer1_outputs(3163) <= a;
    layer1_outputs(3164) <= not (a and b);
    layer1_outputs(3165) <= not (a xor b);
    layer1_outputs(3166) <= a or b;
    layer1_outputs(3167) <= a or b;
    layer1_outputs(3168) <= b and not a;
    layer1_outputs(3169) <= a or b;
    layer1_outputs(3170) <= '1';
    layer1_outputs(3171) <= a and b;
    layer1_outputs(3172) <= '1';
    layer1_outputs(3173) <= not b or a;
    layer1_outputs(3174) <= not (a and b);
    layer1_outputs(3175) <= not a or b;
    layer1_outputs(3176) <= a xor b;
    layer1_outputs(3177) <= b;
    layer1_outputs(3178) <= a and not b;
    layer1_outputs(3179) <= a and not b;
    layer1_outputs(3180) <= b and not a;
    layer1_outputs(3181) <= not (a or b);
    layer1_outputs(3182) <= b and not a;
    layer1_outputs(3183) <= not b or a;
    layer1_outputs(3184) <= not b or a;
    layer1_outputs(3185) <= not a or b;
    layer1_outputs(3186) <= not a;
    layer1_outputs(3187) <= a and b;
    layer1_outputs(3188) <= a xor b;
    layer1_outputs(3189) <= b and not a;
    layer1_outputs(3190) <= b;
    layer1_outputs(3191) <= a or b;
    layer1_outputs(3192) <= not a or b;
    layer1_outputs(3193) <= a;
    layer1_outputs(3194) <= not (a xor b);
    layer1_outputs(3195) <= a xor b;
    layer1_outputs(3196) <= not (a or b);
    layer1_outputs(3197) <= not (a or b);
    layer1_outputs(3198) <= not b;
    layer1_outputs(3199) <= a xor b;
    layer1_outputs(3200) <= a;
    layer1_outputs(3201) <= b;
    layer1_outputs(3202) <= not a or b;
    layer1_outputs(3203) <= a;
    layer1_outputs(3204) <= not b;
    layer1_outputs(3205) <= b;
    layer1_outputs(3206) <= b;
    layer1_outputs(3207) <= b;
    layer1_outputs(3208) <= b;
    layer1_outputs(3209) <= a;
    layer1_outputs(3210) <= not (a xor b);
    layer1_outputs(3211) <= '1';
    layer1_outputs(3212) <= b;
    layer1_outputs(3213) <= not b;
    layer1_outputs(3214) <= a;
    layer1_outputs(3215) <= not (a and b);
    layer1_outputs(3216) <= not a;
    layer1_outputs(3217) <= '0';
    layer1_outputs(3218) <= a;
    layer1_outputs(3219) <= a;
    layer1_outputs(3220) <= not b;
    layer1_outputs(3221) <= not a or b;
    layer1_outputs(3222) <= not b or a;
    layer1_outputs(3223) <= not a;
    layer1_outputs(3224) <= b and not a;
    layer1_outputs(3225) <= a;
    layer1_outputs(3226) <= not (a and b);
    layer1_outputs(3227) <= a;
    layer1_outputs(3228) <= not a or b;
    layer1_outputs(3229) <= not b or a;
    layer1_outputs(3230) <= not b or a;
    layer1_outputs(3231) <= a;
    layer1_outputs(3232) <= not b;
    layer1_outputs(3233) <= not (a xor b);
    layer1_outputs(3234) <= not a;
    layer1_outputs(3235) <= not b;
    layer1_outputs(3236) <= a xor b;
    layer1_outputs(3237) <= a and b;
    layer1_outputs(3238) <= b;
    layer1_outputs(3239) <= a;
    layer1_outputs(3240) <= not b or a;
    layer1_outputs(3241) <= a and not b;
    layer1_outputs(3242) <= not (a xor b);
    layer1_outputs(3243) <= not b;
    layer1_outputs(3244) <= not b;
    layer1_outputs(3245) <= a;
    layer1_outputs(3246) <= b;
    layer1_outputs(3247) <= not (a or b);
    layer1_outputs(3248) <= a and not b;
    layer1_outputs(3249) <= not (a and b);
    layer1_outputs(3250) <= not (a xor b);
    layer1_outputs(3251) <= b and not a;
    layer1_outputs(3252) <= b and not a;
    layer1_outputs(3253) <= a and not b;
    layer1_outputs(3254) <= a and not b;
    layer1_outputs(3255) <= not a or b;
    layer1_outputs(3256) <= b and not a;
    layer1_outputs(3257) <= a;
    layer1_outputs(3258) <= a and b;
    layer1_outputs(3259) <= b;
    layer1_outputs(3260) <= not b or a;
    layer1_outputs(3261) <= not a;
    layer1_outputs(3262) <= not a;
    layer1_outputs(3263) <= not b or a;
    layer1_outputs(3264) <= not b or a;
    layer1_outputs(3265) <= b and not a;
    layer1_outputs(3266) <= not (a or b);
    layer1_outputs(3267) <= a;
    layer1_outputs(3268) <= not (a xor b);
    layer1_outputs(3269) <= a;
    layer1_outputs(3270) <= b;
    layer1_outputs(3271) <= a and b;
    layer1_outputs(3272) <= not a;
    layer1_outputs(3273) <= a and not b;
    layer1_outputs(3274) <= b;
    layer1_outputs(3275) <= b;
    layer1_outputs(3276) <= a xor b;
    layer1_outputs(3277) <= b;
    layer1_outputs(3278) <= not a;
    layer1_outputs(3279) <= a xor b;
    layer1_outputs(3280) <= a and not b;
    layer1_outputs(3281) <= b and not a;
    layer1_outputs(3282) <= a and not b;
    layer1_outputs(3283) <= not b or a;
    layer1_outputs(3284) <= not (a xor b);
    layer1_outputs(3285) <= a xor b;
    layer1_outputs(3286) <= a;
    layer1_outputs(3287) <= not a or b;
    layer1_outputs(3288) <= a or b;
    layer1_outputs(3289) <= a xor b;
    layer1_outputs(3290) <= a or b;
    layer1_outputs(3291) <= not b;
    layer1_outputs(3292) <= not a or b;
    layer1_outputs(3293) <= not b or a;
    layer1_outputs(3294) <= not a;
    layer1_outputs(3295) <= not a or b;
    layer1_outputs(3296) <= a;
    layer1_outputs(3297) <= not (a or b);
    layer1_outputs(3298) <= not (a and b);
    layer1_outputs(3299) <= a and b;
    layer1_outputs(3300) <= a xor b;
    layer1_outputs(3301) <= not (a and b);
    layer1_outputs(3302) <= not a;
    layer1_outputs(3303) <= not b;
    layer1_outputs(3304) <= a or b;
    layer1_outputs(3305) <= b;
    layer1_outputs(3306) <= a or b;
    layer1_outputs(3307) <= b and not a;
    layer1_outputs(3308) <= b;
    layer1_outputs(3309) <= b;
    layer1_outputs(3310) <= not (a or b);
    layer1_outputs(3311) <= a xor b;
    layer1_outputs(3312) <= not b;
    layer1_outputs(3313) <= a xor b;
    layer1_outputs(3314) <= a or b;
    layer1_outputs(3315) <= a and b;
    layer1_outputs(3316) <= a xor b;
    layer1_outputs(3317) <= a and b;
    layer1_outputs(3318) <= not (a xor b);
    layer1_outputs(3319) <= a and b;
    layer1_outputs(3320) <= a;
    layer1_outputs(3321) <= not (a xor b);
    layer1_outputs(3322) <= not (a xor b);
    layer1_outputs(3323) <= not b or a;
    layer1_outputs(3324) <= b and not a;
    layer1_outputs(3325) <= a xor b;
    layer1_outputs(3326) <= not b;
    layer1_outputs(3327) <= '0';
    layer1_outputs(3328) <= a xor b;
    layer1_outputs(3329) <= a and b;
    layer1_outputs(3330) <= not b or a;
    layer1_outputs(3331) <= a xor b;
    layer1_outputs(3332) <= b and not a;
    layer1_outputs(3333) <= b and not a;
    layer1_outputs(3334) <= a xor b;
    layer1_outputs(3335) <= '0';
    layer1_outputs(3336) <= a and not b;
    layer1_outputs(3337) <= not a or b;
    layer1_outputs(3338) <= a and b;
    layer1_outputs(3339) <= not (a and b);
    layer1_outputs(3340) <= not a or b;
    layer1_outputs(3341) <= a and b;
    layer1_outputs(3342) <= b;
    layer1_outputs(3343) <= a;
    layer1_outputs(3344) <= not b or a;
    layer1_outputs(3345) <= not (a or b);
    layer1_outputs(3346) <= not b;
    layer1_outputs(3347) <= b;
    layer1_outputs(3348) <= not (a and b);
    layer1_outputs(3349) <= a;
    layer1_outputs(3350) <= a and b;
    layer1_outputs(3351) <= a;
    layer1_outputs(3352) <= not b;
    layer1_outputs(3353) <= a;
    layer1_outputs(3354) <= b;
    layer1_outputs(3355) <= not (a or b);
    layer1_outputs(3356) <= a and not b;
    layer1_outputs(3357) <= not (a and b);
    layer1_outputs(3358) <= a;
    layer1_outputs(3359) <= not a;
    layer1_outputs(3360) <= not b or a;
    layer1_outputs(3361) <= not (a or b);
    layer1_outputs(3362) <= a xor b;
    layer1_outputs(3363) <= not b;
    layer1_outputs(3364) <= not b;
    layer1_outputs(3365) <= a xor b;
    layer1_outputs(3366) <= not (a or b);
    layer1_outputs(3367) <= b;
    layer1_outputs(3368) <= not b;
    layer1_outputs(3369) <= b and not a;
    layer1_outputs(3370) <= a or b;
    layer1_outputs(3371) <= not (a xor b);
    layer1_outputs(3372) <= not b or a;
    layer1_outputs(3373) <= a xor b;
    layer1_outputs(3374) <= not b;
    layer1_outputs(3375) <= a and not b;
    layer1_outputs(3376) <= not b or a;
    layer1_outputs(3377) <= a and b;
    layer1_outputs(3378) <= b and not a;
    layer1_outputs(3379) <= a xor b;
    layer1_outputs(3380) <= a or b;
    layer1_outputs(3381) <= a;
    layer1_outputs(3382) <= b and not a;
    layer1_outputs(3383) <= b;
    layer1_outputs(3384) <= not a or b;
    layer1_outputs(3385) <= not (a xor b);
    layer1_outputs(3386) <= not b;
    layer1_outputs(3387) <= a and not b;
    layer1_outputs(3388) <= not (a or b);
    layer1_outputs(3389) <= not (a or b);
    layer1_outputs(3390) <= a and b;
    layer1_outputs(3391) <= not a;
    layer1_outputs(3392) <= a and b;
    layer1_outputs(3393) <= a or b;
    layer1_outputs(3394) <= a or b;
    layer1_outputs(3395) <= a and b;
    layer1_outputs(3396) <= not (a or b);
    layer1_outputs(3397) <= b;
    layer1_outputs(3398) <= not b;
    layer1_outputs(3399) <= a;
    layer1_outputs(3400) <= not a;
    layer1_outputs(3401) <= not (a xor b);
    layer1_outputs(3402) <= not (a or b);
    layer1_outputs(3403) <= a;
    layer1_outputs(3404) <= not a;
    layer1_outputs(3405) <= b;
    layer1_outputs(3406) <= a;
    layer1_outputs(3407) <= not (a and b);
    layer1_outputs(3408) <= not (a and b);
    layer1_outputs(3409) <= not a;
    layer1_outputs(3410) <= not (a xor b);
    layer1_outputs(3411) <= not b or a;
    layer1_outputs(3412) <= not a or b;
    layer1_outputs(3413) <= a;
    layer1_outputs(3414) <= not a or b;
    layer1_outputs(3415) <= a;
    layer1_outputs(3416) <= b and not a;
    layer1_outputs(3417) <= not a or b;
    layer1_outputs(3418) <= a or b;
    layer1_outputs(3419) <= b;
    layer1_outputs(3420) <= a and b;
    layer1_outputs(3421) <= not b;
    layer1_outputs(3422) <= not a;
    layer1_outputs(3423) <= b;
    layer1_outputs(3424) <= '0';
    layer1_outputs(3425) <= not a or b;
    layer1_outputs(3426) <= not (a xor b);
    layer1_outputs(3427) <= a;
    layer1_outputs(3428) <= b;
    layer1_outputs(3429) <= a or b;
    layer1_outputs(3430) <= a and b;
    layer1_outputs(3431) <= a;
    layer1_outputs(3432) <= a;
    layer1_outputs(3433) <= a or b;
    layer1_outputs(3434) <= b and not a;
    layer1_outputs(3435) <= not b or a;
    layer1_outputs(3436) <= not a or b;
    layer1_outputs(3437) <= a or b;
    layer1_outputs(3438) <= not b or a;
    layer1_outputs(3439) <= b and not a;
    layer1_outputs(3440) <= b;
    layer1_outputs(3441) <= not b;
    layer1_outputs(3442) <= b and not a;
    layer1_outputs(3443) <= a and not b;
    layer1_outputs(3444) <= not a;
    layer1_outputs(3445) <= not a;
    layer1_outputs(3446) <= a;
    layer1_outputs(3447) <= a and not b;
    layer1_outputs(3448) <= not b or a;
    layer1_outputs(3449) <= not a;
    layer1_outputs(3450) <= a;
    layer1_outputs(3451) <= '0';
    layer1_outputs(3452) <= a and not b;
    layer1_outputs(3453) <= not (a xor b);
    layer1_outputs(3454) <= not (a or b);
    layer1_outputs(3455) <= b;
    layer1_outputs(3456) <= a;
    layer1_outputs(3457) <= not a or b;
    layer1_outputs(3458) <= not (a and b);
    layer1_outputs(3459) <= a xor b;
    layer1_outputs(3460) <= not (a xor b);
    layer1_outputs(3461) <= not a;
    layer1_outputs(3462) <= not a or b;
    layer1_outputs(3463) <= not (a xor b);
    layer1_outputs(3464) <= a or b;
    layer1_outputs(3465) <= not (a xor b);
    layer1_outputs(3466) <= b;
    layer1_outputs(3467) <= not b;
    layer1_outputs(3468) <= not b;
    layer1_outputs(3469) <= not (a and b);
    layer1_outputs(3470) <= not b;
    layer1_outputs(3471) <= not b;
    layer1_outputs(3472) <= a xor b;
    layer1_outputs(3473) <= not a;
    layer1_outputs(3474) <= a and b;
    layer1_outputs(3475) <= a and not b;
    layer1_outputs(3476) <= not (a xor b);
    layer1_outputs(3477) <= not (a xor b);
    layer1_outputs(3478) <= not (a and b);
    layer1_outputs(3479) <= not a;
    layer1_outputs(3480) <= a xor b;
    layer1_outputs(3481) <= not (a and b);
    layer1_outputs(3482) <= a;
    layer1_outputs(3483) <= not a or b;
    layer1_outputs(3484) <= not a or b;
    layer1_outputs(3485) <= not b;
    layer1_outputs(3486) <= a xor b;
    layer1_outputs(3487) <= not (a or b);
    layer1_outputs(3488) <= not a;
    layer1_outputs(3489) <= a or b;
    layer1_outputs(3490) <= not b;
    layer1_outputs(3491) <= not a or b;
    layer1_outputs(3492) <= not (a and b);
    layer1_outputs(3493) <= not (a and b);
    layer1_outputs(3494) <= not (a xor b);
    layer1_outputs(3495) <= a and not b;
    layer1_outputs(3496) <= not (a or b);
    layer1_outputs(3497) <= not (a or b);
    layer1_outputs(3498) <= not (a or b);
    layer1_outputs(3499) <= a;
    layer1_outputs(3500) <= a xor b;
    layer1_outputs(3501) <= '1';
    layer1_outputs(3502) <= b and not a;
    layer1_outputs(3503) <= a;
    layer1_outputs(3504) <= a;
    layer1_outputs(3505) <= b;
    layer1_outputs(3506) <= a or b;
    layer1_outputs(3507) <= a;
    layer1_outputs(3508) <= a xor b;
    layer1_outputs(3509) <= b;
    layer1_outputs(3510) <= not b;
    layer1_outputs(3511) <= a or b;
    layer1_outputs(3512) <= a;
    layer1_outputs(3513) <= not b;
    layer1_outputs(3514) <= a or b;
    layer1_outputs(3515) <= b and not a;
    layer1_outputs(3516) <= not a;
    layer1_outputs(3517) <= not b;
    layer1_outputs(3518) <= a or b;
    layer1_outputs(3519) <= a and b;
    layer1_outputs(3520) <= a xor b;
    layer1_outputs(3521) <= a;
    layer1_outputs(3522) <= not b;
    layer1_outputs(3523) <= a;
    layer1_outputs(3524) <= a and b;
    layer1_outputs(3525) <= b;
    layer1_outputs(3526) <= '0';
    layer1_outputs(3527) <= not a or b;
    layer1_outputs(3528) <= not (a xor b);
    layer1_outputs(3529) <= '1';
    layer1_outputs(3530) <= not b;
    layer1_outputs(3531) <= not b;
    layer1_outputs(3532) <= a and not b;
    layer1_outputs(3533) <= a;
    layer1_outputs(3534) <= not a or b;
    layer1_outputs(3535) <= a and b;
    layer1_outputs(3536) <= not a or b;
    layer1_outputs(3537) <= a;
    layer1_outputs(3538) <= a;
    layer1_outputs(3539) <= a and not b;
    layer1_outputs(3540) <= not a or b;
    layer1_outputs(3541) <= a or b;
    layer1_outputs(3542) <= not a or b;
    layer1_outputs(3543) <= not b;
    layer1_outputs(3544) <= a;
    layer1_outputs(3545) <= a or b;
    layer1_outputs(3546) <= not b;
    layer1_outputs(3547) <= a and not b;
    layer1_outputs(3548) <= b;
    layer1_outputs(3549) <= a;
    layer1_outputs(3550) <= a or b;
    layer1_outputs(3551) <= not (a and b);
    layer1_outputs(3552) <= a or b;
    layer1_outputs(3553) <= a;
    layer1_outputs(3554) <= not b;
    layer1_outputs(3555) <= not a;
    layer1_outputs(3556) <= '0';
    layer1_outputs(3557) <= not a;
    layer1_outputs(3558) <= a;
    layer1_outputs(3559) <= not (a and b);
    layer1_outputs(3560) <= not a or b;
    layer1_outputs(3561) <= a or b;
    layer1_outputs(3562) <= not a;
    layer1_outputs(3563) <= not b;
    layer1_outputs(3564) <= not b;
    layer1_outputs(3565) <= a or b;
    layer1_outputs(3566) <= a and b;
    layer1_outputs(3567) <= not b or a;
    layer1_outputs(3568) <= b;
    layer1_outputs(3569) <= b and not a;
    layer1_outputs(3570) <= a xor b;
    layer1_outputs(3571) <= not (a xor b);
    layer1_outputs(3572) <= b;
    layer1_outputs(3573) <= not (a or b);
    layer1_outputs(3574) <= b;
    layer1_outputs(3575) <= not b;
    layer1_outputs(3576) <= a xor b;
    layer1_outputs(3577) <= b;
    layer1_outputs(3578) <= a;
    layer1_outputs(3579) <= not a or b;
    layer1_outputs(3580) <= not (a xor b);
    layer1_outputs(3581) <= b;
    layer1_outputs(3582) <= a xor b;
    layer1_outputs(3583) <= a and not b;
    layer1_outputs(3584) <= b;
    layer1_outputs(3585) <= not b or a;
    layer1_outputs(3586) <= a xor b;
    layer1_outputs(3587) <= not b or a;
    layer1_outputs(3588) <= not (a and b);
    layer1_outputs(3589) <= not a;
    layer1_outputs(3590) <= a and not b;
    layer1_outputs(3591) <= a;
    layer1_outputs(3592) <= not a;
    layer1_outputs(3593) <= a and not b;
    layer1_outputs(3594) <= not (a xor b);
    layer1_outputs(3595) <= not (a or b);
    layer1_outputs(3596) <= not (a or b);
    layer1_outputs(3597) <= a and not b;
    layer1_outputs(3598) <= b and not a;
    layer1_outputs(3599) <= a and not b;
    layer1_outputs(3600) <= a;
    layer1_outputs(3601) <= not a;
    layer1_outputs(3602) <= '0';
    layer1_outputs(3603) <= not (a and b);
    layer1_outputs(3604) <= not a;
    layer1_outputs(3605) <= not b or a;
    layer1_outputs(3606) <= b;
    layer1_outputs(3607) <= not b;
    layer1_outputs(3608) <= a and b;
    layer1_outputs(3609) <= a or b;
    layer1_outputs(3610) <= not a;
    layer1_outputs(3611) <= a and b;
    layer1_outputs(3612) <= b;
    layer1_outputs(3613) <= b and not a;
    layer1_outputs(3614) <= a or b;
    layer1_outputs(3615) <= not (a or b);
    layer1_outputs(3616) <= a xor b;
    layer1_outputs(3617) <= a or b;
    layer1_outputs(3618) <= b;
    layer1_outputs(3619) <= a;
    layer1_outputs(3620) <= b and not a;
    layer1_outputs(3621) <= not (a xor b);
    layer1_outputs(3622) <= b;
    layer1_outputs(3623) <= a;
    layer1_outputs(3624) <= a or b;
    layer1_outputs(3625) <= not b;
    layer1_outputs(3626) <= not a or b;
    layer1_outputs(3627) <= not (a or b);
    layer1_outputs(3628) <= b and not a;
    layer1_outputs(3629) <= not (a xor b);
    layer1_outputs(3630) <= not b or a;
    layer1_outputs(3631) <= a or b;
    layer1_outputs(3632) <= a xor b;
    layer1_outputs(3633) <= not a;
    layer1_outputs(3634) <= a;
    layer1_outputs(3635) <= not a or b;
    layer1_outputs(3636) <= not b;
    layer1_outputs(3637) <= b and not a;
    layer1_outputs(3638) <= b;
    layer1_outputs(3639) <= b and not a;
    layer1_outputs(3640) <= not (a or b);
    layer1_outputs(3641) <= not a or b;
    layer1_outputs(3642) <= not a or b;
    layer1_outputs(3643) <= a and b;
    layer1_outputs(3644) <= a xor b;
    layer1_outputs(3645) <= not a;
    layer1_outputs(3646) <= a or b;
    layer1_outputs(3647) <= a xor b;
    layer1_outputs(3648) <= not b;
    layer1_outputs(3649) <= a and b;
    layer1_outputs(3650) <= a;
    layer1_outputs(3651) <= not (a xor b);
    layer1_outputs(3652) <= b and not a;
    layer1_outputs(3653) <= not a or b;
    layer1_outputs(3654) <= b;
    layer1_outputs(3655) <= b;
    layer1_outputs(3656) <= b;
    layer1_outputs(3657) <= a or b;
    layer1_outputs(3658) <= not (a or b);
    layer1_outputs(3659) <= not (a and b);
    layer1_outputs(3660) <= b;
    layer1_outputs(3661) <= b and not a;
    layer1_outputs(3662) <= a and not b;
    layer1_outputs(3663) <= a and not b;
    layer1_outputs(3664) <= a or b;
    layer1_outputs(3665) <= b and not a;
    layer1_outputs(3666) <= not b or a;
    layer1_outputs(3667) <= not a;
    layer1_outputs(3668) <= b;
    layer1_outputs(3669) <= not (a or b);
    layer1_outputs(3670) <= b and not a;
    layer1_outputs(3671) <= not a;
    layer1_outputs(3672) <= not a;
    layer1_outputs(3673) <= b;
    layer1_outputs(3674) <= a or b;
    layer1_outputs(3675) <= a;
    layer1_outputs(3676) <= not a;
    layer1_outputs(3677) <= a;
    layer1_outputs(3678) <= not b;
    layer1_outputs(3679) <= a xor b;
    layer1_outputs(3680) <= not a;
    layer1_outputs(3681) <= a or b;
    layer1_outputs(3682) <= a xor b;
    layer1_outputs(3683) <= not a;
    layer1_outputs(3684) <= not a or b;
    layer1_outputs(3685) <= not a;
    layer1_outputs(3686) <= a and b;
    layer1_outputs(3687) <= not (a xor b);
    layer1_outputs(3688) <= a and not b;
    layer1_outputs(3689) <= not (a and b);
    layer1_outputs(3690) <= not a;
    layer1_outputs(3691) <= a and b;
    layer1_outputs(3692) <= b;
    layer1_outputs(3693) <= a and not b;
    layer1_outputs(3694) <= b and not a;
    layer1_outputs(3695) <= not b;
    layer1_outputs(3696) <= b and not a;
    layer1_outputs(3697) <= a;
    layer1_outputs(3698) <= b;
    layer1_outputs(3699) <= not (a xor b);
    layer1_outputs(3700) <= a;
    layer1_outputs(3701) <= not (a xor b);
    layer1_outputs(3702) <= b;
    layer1_outputs(3703) <= not a;
    layer1_outputs(3704) <= not (a and b);
    layer1_outputs(3705) <= not (a and b);
    layer1_outputs(3706) <= a or b;
    layer1_outputs(3707) <= not (a xor b);
    layer1_outputs(3708) <= not b or a;
    layer1_outputs(3709) <= b;
    layer1_outputs(3710) <= not a;
    layer1_outputs(3711) <= not (a and b);
    layer1_outputs(3712) <= a;
    layer1_outputs(3713) <= '0';
    layer1_outputs(3714) <= not a or b;
    layer1_outputs(3715) <= b and not a;
    layer1_outputs(3716) <= b;
    layer1_outputs(3717) <= '1';
    layer1_outputs(3718) <= b and not a;
    layer1_outputs(3719) <= b;
    layer1_outputs(3720) <= not b;
    layer1_outputs(3721) <= not b or a;
    layer1_outputs(3722) <= a and b;
    layer1_outputs(3723) <= a or b;
    layer1_outputs(3724) <= a or b;
    layer1_outputs(3725) <= not b;
    layer1_outputs(3726) <= not (a and b);
    layer1_outputs(3727) <= a or b;
    layer1_outputs(3728) <= not (a and b);
    layer1_outputs(3729) <= not a;
    layer1_outputs(3730) <= not a or b;
    layer1_outputs(3731) <= a and b;
    layer1_outputs(3732) <= '0';
    layer1_outputs(3733) <= a;
    layer1_outputs(3734) <= not (a xor b);
    layer1_outputs(3735) <= not (a and b);
    layer1_outputs(3736) <= a or b;
    layer1_outputs(3737) <= not (a xor b);
    layer1_outputs(3738) <= b and not a;
    layer1_outputs(3739) <= a;
    layer1_outputs(3740) <= not a;
    layer1_outputs(3741) <= '0';
    layer1_outputs(3742) <= not a;
    layer1_outputs(3743) <= a;
    layer1_outputs(3744) <= not (a and b);
    layer1_outputs(3745) <= b and not a;
    layer1_outputs(3746) <= not b or a;
    layer1_outputs(3747) <= a;
    layer1_outputs(3748) <= not a or b;
    layer1_outputs(3749) <= not b;
    layer1_outputs(3750) <= not (a xor b);
    layer1_outputs(3751) <= a and b;
    layer1_outputs(3752) <= b and not a;
    layer1_outputs(3753) <= a and b;
    layer1_outputs(3754) <= not a;
    layer1_outputs(3755) <= a and b;
    layer1_outputs(3756) <= b;
    layer1_outputs(3757) <= not (a xor b);
    layer1_outputs(3758) <= a and not b;
    layer1_outputs(3759) <= a and not b;
    layer1_outputs(3760) <= not (a and b);
    layer1_outputs(3761) <= not a;
    layer1_outputs(3762) <= a and b;
    layer1_outputs(3763) <= not a;
    layer1_outputs(3764) <= not a;
    layer1_outputs(3765) <= not (a or b);
    layer1_outputs(3766) <= not a;
    layer1_outputs(3767) <= a and b;
    layer1_outputs(3768) <= a;
    layer1_outputs(3769) <= b;
    layer1_outputs(3770) <= a and b;
    layer1_outputs(3771) <= a and not b;
    layer1_outputs(3772) <= a;
    layer1_outputs(3773) <= a or b;
    layer1_outputs(3774) <= a and b;
    layer1_outputs(3775) <= not (a xor b);
    layer1_outputs(3776) <= a xor b;
    layer1_outputs(3777) <= not (a xor b);
    layer1_outputs(3778) <= a and not b;
    layer1_outputs(3779) <= not b;
    layer1_outputs(3780) <= a;
    layer1_outputs(3781) <= a;
    layer1_outputs(3782) <= not (a xor b);
    layer1_outputs(3783) <= not (a and b);
    layer1_outputs(3784) <= a xor b;
    layer1_outputs(3785) <= not (a xor b);
    layer1_outputs(3786) <= a and not b;
    layer1_outputs(3787) <= not (a and b);
    layer1_outputs(3788) <= '1';
    layer1_outputs(3789) <= not b;
    layer1_outputs(3790) <= not (a or b);
    layer1_outputs(3791) <= b and not a;
    layer1_outputs(3792) <= not b;
    layer1_outputs(3793) <= a;
    layer1_outputs(3794) <= a and b;
    layer1_outputs(3795) <= not b;
    layer1_outputs(3796) <= not (a xor b);
    layer1_outputs(3797) <= not (a xor b);
    layer1_outputs(3798) <= not a;
    layer1_outputs(3799) <= not (a and b);
    layer1_outputs(3800) <= not b;
    layer1_outputs(3801) <= '1';
    layer1_outputs(3802) <= a or b;
    layer1_outputs(3803) <= not (a xor b);
    layer1_outputs(3804) <= a;
    layer1_outputs(3805) <= not (a or b);
    layer1_outputs(3806) <= a and not b;
    layer1_outputs(3807) <= a xor b;
    layer1_outputs(3808) <= not a or b;
    layer1_outputs(3809) <= not b;
    layer1_outputs(3810) <= a xor b;
    layer1_outputs(3811) <= not a;
    layer1_outputs(3812) <= not a;
    layer1_outputs(3813) <= not a;
    layer1_outputs(3814) <= not (a xor b);
    layer1_outputs(3815) <= b;
    layer1_outputs(3816) <= b;
    layer1_outputs(3817) <= not a;
    layer1_outputs(3818) <= not b or a;
    layer1_outputs(3819) <= not (a or b);
    layer1_outputs(3820) <= b;
    layer1_outputs(3821) <= b and not a;
    layer1_outputs(3822) <= a and b;
    layer1_outputs(3823) <= a and b;
    layer1_outputs(3824) <= not (a or b);
    layer1_outputs(3825) <= not b or a;
    layer1_outputs(3826) <= a and not b;
    layer1_outputs(3827) <= a;
    layer1_outputs(3828) <= a and b;
    layer1_outputs(3829) <= a xor b;
    layer1_outputs(3830) <= not b or a;
    layer1_outputs(3831) <= a xor b;
    layer1_outputs(3832) <= '1';
    layer1_outputs(3833) <= a xor b;
    layer1_outputs(3834) <= not (a and b);
    layer1_outputs(3835) <= not b;
    layer1_outputs(3836) <= a;
    layer1_outputs(3837) <= b;
    layer1_outputs(3838) <= not a or b;
    layer1_outputs(3839) <= not (a xor b);
    layer1_outputs(3840) <= not b or a;
    layer1_outputs(3841) <= a and not b;
    layer1_outputs(3842) <= not b;
    layer1_outputs(3843) <= a xor b;
    layer1_outputs(3844) <= not a or b;
    layer1_outputs(3845) <= b;
    layer1_outputs(3846) <= not b;
    layer1_outputs(3847) <= '1';
    layer1_outputs(3848) <= not a;
    layer1_outputs(3849) <= b;
    layer1_outputs(3850) <= b and not a;
    layer1_outputs(3851) <= a or b;
    layer1_outputs(3852) <= b and not a;
    layer1_outputs(3853) <= not a;
    layer1_outputs(3854) <= b and not a;
    layer1_outputs(3855) <= a and not b;
    layer1_outputs(3856) <= not a or b;
    layer1_outputs(3857) <= a xor b;
    layer1_outputs(3858) <= not (a xor b);
    layer1_outputs(3859) <= not (a xor b);
    layer1_outputs(3860) <= not (a xor b);
    layer1_outputs(3861) <= a xor b;
    layer1_outputs(3862) <= not (a and b);
    layer1_outputs(3863) <= not (a and b);
    layer1_outputs(3864) <= a;
    layer1_outputs(3865) <= a and not b;
    layer1_outputs(3866) <= not (a xor b);
    layer1_outputs(3867) <= not a or b;
    layer1_outputs(3868) <= not b;
    layer1_outputs(3869) <= not a;
    layer1_outputs(3870) <= not (a or b);
    layer1_outputs(3871) <= not a or b;
    layer1_outputs(3872) <= not (a and b);
    layer1_outputs(3873) <= not (a and b);
    layer1_outputs(3874) <= not b;
    layer1_outputs(3875) <= not a;
    layer1_outputs(3876) <= b;
    layer1_outputs(3877) <= a or b;
    layer1_outputs(3878) <= not (a and b);
    layer1_outputs(3879) <= a xor b;
    layer1_outputs(3880) <= a and not b;
    layer1_outputs(3881) <= not b;
    layer1_outputs(3882) <= a or b;
    layer1_outputs(3883) <= not a or b;
    layer1_outputs(3884) <= a xor b;
    layer1_outputs(3885) <= not b;
    layer1_outputs(3886) <= a;
    layer1_outputs(3887) <= a and b;
    layer1_outputs(3888) <= not (a or b);
    layer1_outputs(3889) <= a;
    layer1_outputs(3890) <= not b;
    layer1_outputs(3891) <= not (a xor b);
    layer1_outputs(3892) <= not b or a;
    layer1_outputs(3893) <= not (a or b);
    layer1_outputs(3894) <= a and b;
    layer1_outputs(3895) <= b;
    layer1_outputs(3896) <= not b;
    layer1_outputs(3897) <= not b;
    layer1_outputs(3898) <= b and not a;
    layer1_outputs(3899) <= not (a xor b);
    layer1_outputs(3900) <= not (a or b);
    layer1_outputs(3901) <= not a;
    layer1_outputs(3902) <= a xor b;
    layer1_outputs(3903) <= not b;
    layer1_outputs(3904) <= not (a xor b);
    layer1_outputs(3905) <= not a or b;
    layer1_outputs(3906) <= a and not b;
    layer1_outputs(3907) <= a and b;
    layer1_outputs(3908) <= not a;
    layer1_outputs(3909) <= not (a and b);
    layer1_outputs(3910) <= not (a xor b);
    layer1_outputs(3911) <= not b or a;
    layer1_outputs(3912) <= a and not b;
    layer1_outputs(3913) <= a and b;
    layer1_outputs(3914) <= a;
    layer1_outputs(3915) <= not (a xor b);
    layer1_outputs(3916) <= not a or b;
    layer1_outputs(3917) <= a xor b;
    layer1_outputs(3918) <= b and not a;
    layer1_outputs(3919) <= not b or a;
    layer1_outputs(3920) <= not (a xor b);
    layer1_outputs(3921) <= a or b;
    layer1_outputs(3922) <= a xor b;
    layer1_outputs(3923) <= not a or b;
    layer1_outputs(3924) <= not b;
    layer1_outputs(3925) <= not a;
    layer1_outputs(3926) <= '1';
    layer1_outputs(3927) <= not b;
    layer1_outputs(3928) <= a and not b;
    layer1_outputs(3929) <= a and b;
    layer1_outputs(3930) <= '1';
    layer1_outputs(3931) <= a or b;
    layer1_outputs(3932) <= not (a or b);
    layer1_outputs(3933) <= b;
    layer1_outputs(3934) <= not b;
    layer1_outputs(3935) <= a xor b;
    layer1_outputs(3936) <= not (a xor b);
    layer1_outputs(3937) <= not (a and b);
    layer1_outputs(3938) <= not b;
    layer1_outputs(3939) <= b and not a;
    layer1_outputs(3940) <= a and not b;
    layer1_outputs(3941) <= a or b;
    layer1_outputs(3942) <= a xor b;
    layer1_outputs(3943) <= b;
    layer1_outputs(3944) <= not (a xor b);
    layer1_outputs(3945) <= b;
    layer1_outputs(3946) <= b;
    layer1_outputs(3947) <= a or b;
    layer1_outputs(3948) <= a and b;
    layer1_outputs(3949) <= not (a and b);
    layer1_outputs(3950) <= not (a xor b);
    layer1_outputs(3951) <= not (a xor b);
    layer1_outputs(3952) <= not (a and b);
    layer1_outputs(3953) <= not a;
    layer1_outputs(3954) <= '1';
    layer1_outputs(3955) <= not b;
    layer1_outputs(3956) <= not (a or b);
    layer1_outputs(3957) <= a and not b;
    layer1_outputs(3958) <= not (a and b);
    layer1_outputs(3959) <= not b or a;
    layer1_outputs(3960) <= b;
    layer1_outputs(3961) <= a;
    layer1_outputs(3962) <= a and not b;
    layer1_outputs(3963) <= a and b;
    layer1_outputs(3964) <= a;
    layer1_outputs(3965) <= a and b;
    layer1_outputs(3966) <= b;
    layer1_outputs(3967) <= not (a xor b);
    layer1_outputs(3968) <= not a or b;
    layer1_outputs(3969) <= not (a and b);
    layer1_outputs(3970) <= not a;
    layer1_outputs(3971) <= not b;
    layer1_outputs(3972) <= b and not a;
    layer1_outputs(3973) <= not b;
    layer1_outputs(3974) <= not a;
    layer1_outputs(3975) <= a and not b;
    layer1_outputs(3976) <= a and not b;
    layer1_outputs(3977) <= not a;
    layer1_outputs(3978) <= '0';
    layer1_outputs(3979) <= not (a xor b);
    layer1_outputs(3980) <= a xor b;
    layer1_outputs(3981) <= not a;
    layer1_outputs(3982) <= a and b;
    layer1_outputs(3983) <= not (a or b);
    layer1_outputs(3984) <= a and b;
    layer1_outputs(3985) <= not a;
    layer1_outputs(3986) <= a xor b;
    layer1_outputs(3987) <= a;
    layer1_outputs(3988) <= not (a xor b);
    layer1_outputs(3989) <= a and b;
    layer1_outputs(3990) <= not b or a;
    layer1_outputs(3991) <= a;
    layer1_outputs(3992) <= not a or b;
    layer1_outputs(3993) <= a and b;
    layer1_outputs(3994) <= a or b;
    layer1_outputs(3995) <= not a;
    layer1_outputs(3996) <= not b or a;
    layer1_outputs(3997) <= a and not b;
    layer1_outputs(3998) <= not (a or b);
    layer1_outputs(3999) <= b and not a;
    layer1_outputs(4000) <= not a or b;
    layer1_outputs(4001) <= b;
    layer1_outputs(4002) <= not (a or b);
    layer1_outputs(4003) <= not a;
    layer1_outputs(4004) <= not b;
    layer1_outputs(4005) <= not b;
    layer1_outputs(4006) <= b;
    layer1_outputs(4007) <= not (a xor b);
    layer1_outputs(4008) <= not a or b;
    layer1_outputs(4009) <= not b or a;
    layer1_outputs(4010) <= a;
    layer1_outputs(4011) <= a;
    layer1_outputs(4012) <= not (a and b);
    layer1_outputs(4013) <= a or b;
    layer1_outputs(4014) <= not a;
    layer1_outputs(4015) <= a xor b;
    layer1_outputs(4016) <= not (a and b);
    layer1_outputs(4017) <= not b or a;
    layer1_outputs(4018) <= a or b;
    layer1_outputs(4019) <= not a;
    layer1_outputs(4020) <= a xor b;
    layer1_outputs(4021) <= not a or b;
    layer1_outputs(4022) <= a and not b;
    layer1_outputs(4023) <= a xor b;
    layer1_outputs(4024) <= a xor b;
    layer1_outputs(4025) <= a xor b;
    layer1_outputs(4026) <= a and not b;
    layer1_outputs(4027) <= b;
    layer1_outputs(4028) <= not a;
    layer1_outputs(4029) <= not (a and b);
    layer1_outputs(4030) <= not (a or b);
    layer1_outputs(4031) <= not (a and b);
    layer1_outputs(4032) <= '1';
    layer1_outputs(4033) <= not (a and b);
    layer1_outputs(4034) <= a and b;
    layer1_outputs(4035) <= not (a and b);
    layer1_outputs(4036) <= b and not a;
    layer1_outputs(4037) <= a xor b;
    layer1_outputs(4038) <= not a;
    layer1_outputs(4039) <= '0';
    layer1_outputs(4040) <= not (a xor b);
    layer1_outputs(4041) <= a xor b;
    layer1_outputs(4042) <= not (a or b);
    layer1_outputs(4043) <= a xor b;
    layer1_outputs(4044) <= not a;
    layer1_outputs(4045) <= a;
    layer1_outputs(4046) <= a and not b;
    layer1_outputs(4047) <= a and b;
    layer1_outputs(4048) <= a and not b;
    layer1_outputs(4049) <= not b;
    layer1_outputs(4050) <= a;
    layer1_outputs(4051) <= a xor b;
    layer1_outputs(4052) <= a;
    layer1_outputs(4053) <= not (a xor b);
    layer1_outputs(4054) <= a xor b;
    layer1_outputs(4055) <= not (a or b);
    layer1_outputs(4056) <= not a;
    layer1_outputs(4057) <= b and not a;
    layer1_outputs(4058) <= not b;
    layer1_outputs(4059) <= not (a and b);
    layer1_outputs(4060) <= not (a xor b);
    layer1_outputs(4061) <= b and not a;
    layer1_outputs(4062) <= not a or b;
    layer1_outputs(4063) <= a xor b;
    layer1_outputs(4064) <= not a;
    layer1_outputs(4065) <= not (a and b);
    layer1_outputs(4066) <= not (a or b);
    layer1_outputs(4067) <= a xor b;
    layer1_outputs(4068) <= not a or b;
    layer1_outputs(4069) <= b and not a;
    layer1_outputs(4070) <= not a;
    layer1_outputs(4071) <= a;
    layer1_outputs(4072) <= a and not b;
    layer1_outputs(4073) <= b;
    layer1_outputs(4074) <= '0';
    layer1_outputs(4075) <= a;
    layer1_outputs(4076) <= not a;
    layer1_outputs(4077) <= not a;
    layer1_outputs(4078) <= not a;
    layer1_outputs(4079) <= not (a xor b);
    layer1_outputs(4080) <= not b or a;
    layer1_outputs(4081) <= a and b;
    layer1_outputs(4082) <= b;
    layer1_outputs(4083) <= not (a xor b);
    layer1_outputs(4084) <= a xor b;
    layer1_outputs(4085) <= not a;
    layer1_outputs(4086) <= not b or a;
    layer1_outputs(4087) <= not a;
    layer1_outputs(4088) <= not (a and b);
    layer1_outputs(4089) <= not (a or b);
    layer1_outputs(4090) <= b;
    layer1_outputs(4091) <= not a;
    layer1_outputs(4092) <= not (a xor b);
    layer1_outputs(4093) <= not b;
    layer1_outputs(4094) <= b;
    layer1_outputs(4095) <= a or b;
    layer1_outputs(4096) <= not b;
    layer1_outputs(4097) <= not (a xor b);
    layer1_outputs(4098) <= not (a xor b);
    layer1_outputs(4099) <= not (a or b);
    layer1_outputs(4100) <= not a;
    layer1_outputs(4101) <= b;
    layer1_outputs(4102) <= not a or b;
    layer1_outputs(4103) <= not (a xor b);
    layer1_outputs(4104) <= not b;
    layer1_outputs(4105) <= b;
    layer1_outputs(4106) <= b;
    layer1_outputs(4107) <= not b;
    layer1_outputs(4108) <= not (a xor b);
    layer1_outputs(4109) <= a xor b;
    layer1_outputs(4110) <= not b or a;
    layer1_outputs(4111) <= not b;
    layer1_outputs(4112) <= a;
    layer1_outputs(4113) <= a;
    layer1_outputs(4114) <= b and not a;
    layer1_outputs(4115) <= a xor b;
    layer1_outputs(4116) <= not b;
    layer1_outputs(4117) <= a and b;
    layer1_outputs(4118) <= a or b;
    layer1_outputs(4119) <= b and not a;
    layer1_outputs(4120) <= b;
    layer1_outputs(4121) <= not (a xor b);
    layer1_outputs(4122) <= b and not a;
    layer1_outputs(4123) <= a;
    layer1_outputs(4124) <= a xor b;
    layer1_outputs(4125) <= not (a xor b);
    layer1_outputs(4126) <= a xor b;
    layer1_outputs(4127) <= a;
    layer1_outputs(4128) <= b;
    layer1_outputs(4129) <= not (a and b);
    layer1_outputs(4130) <= not b;
    layer1_outputs(4131) <= not (a xor b);
    layer1_outputs(4132) <= b;
    layer1_outputs(4133) <= '0';
    layer1_outputs(4134) <= a and b;
    layer1_outputs(4135) <= a or b;
    layer1_outputs(4136) <= not (a and b);
    layer1_outputs(4137) <= not b;
    layer1_outputs(4138) <= a and not b;
    layer1_outputs(4139) <= not b or a;
    layer1_outputs(4140) <= not b;
    layer1_outputs(4141) <= not b;
    layer1_outputs(4142) <= not b;
    layer1_outputs(4143) <= a and not b;
    layer1_outputs(4144) <= not (a or b);
    layer1_outputs(4145) <= a and not b;
    layer1_outputs(4146) <= a or b;
    layer1_outputs(4147) <= a and b;
    layer1_outputs(4148) <= '0';
    layer1_outputs(4149) <= a and not b;
    layer1_outputs(4150) <= not (a or b);
    layer1_outputs(4151) <= not a or b;
    layer1_outputs(4152) <= not (a and b);
    layer1_outputs(4153) <= a and not b;
    layer1_outputs(4154) <= a and b;
    layer1_outputs(4155) <= b;
    layer1_outputs(4156) <= not a or b;
    layer1_outputs(4157) <= b;
    layer1_outputs(4158) <= not (a xor b);
    layer1_outputs(4159) <= not b;
    layer1_outputs(4160) <= b and not a;
    layer1_outputs(4161) <= not b or a;
    layer1_outputs(4162) <= not b or a;
    layer1_outputs(4163) <= a or b;
    layer1_outputs(4164) <= not (a and b);
    layer1_outputs(4165) <= b;
    layer1_outputs(4166) <= b;
    layer1_outputs(4167) <= not b;
    layer1_outputs(4168) <= not (a or b);
    layer1_outputs(4169) <= a or b;
    layer1_outputs(4170) <= a and b;
    layer1_outputs(4171) <= a and b;
    layer1_outputs(4172) <= not a;
    layer1_outputs(4173) <= a;
    layer1_outputs(4174) <= not (a xor b);
    layer1_outputs(4175) <= not a;
    layer1_outputs(4176) <= b and not a;
    layer1_outputs(4177) <= a and b;
    layer1_outputs(4178) <= not b;
    layer1_outputs(4179) <= not a or b;
    layer1_outputs(4180) <= not b;
    layer1_outputs(4181) <= not (a and b);
    layer1_outputs(4182) <= not a;
    layer1_outputs(4183) <= not a;
    layer1_outputs(4184) <= a xor b;
    layer1_outputs(4185) <= not (a and b);
    layer1_outputs(4186) <= not (a or b);
    layer1_outputs(4187) <= not (a xor b);
    layer1_outputs(4188) <= not (a or b);
    layer1_outputs(4189) <= not b;
    layer1_outputs(4190) <= b;
    layer1_outputs(4191) <= '0';
    layer1_outputs(4192) <= not b or a;
    layer1_outputs(4193) <= not b or a;
    layer1_outputs(4194) <= a and b;
    layer1_outputs(4195) <= not b;
    layer1_outputs(4196) <= a and b;
    layer1_outputs(4197) <= a or b;
    layer1_outputs(4198) <= not a;
    layer1_outputs(4199) <= a and b;
    layer1_outputs(4200) <= not (a and b);
    layer1_outputs(4201) <= not a or b;
    layer1_outputs(4202) <= not b;
    layer1_outputs(4203) <= a and not b;
    layer1_outputs(4204) <= not a;
    layer1_outputs(4205) <= a and not b;
    layer1_outputs(4206) <= not (a and b);
    layer1_outputs(4207) <= not b;
    layer1_outputs(4208) <= b;
    layer1_outputs(4209) <= not a;
    layer1_outputs(4210) <= a xor b;
    layer1_outputs(4211) <= not b or a;
    layer1_outputs(4212) <= not b;
    layer1_outputs(4213) <= b;
    layer1_outputs(4214) <= not (a or b);
    layer1_outputs(4215) <= '0';
    layer1_outputs(4216) <= b;
    layer1_outputs(4217) <= not b or a;
    layer1_outputs(4218) <= a and not b;
    layer1_outputs(4219) <= not a;
    layer1_outputs(4220) <= not b or a;
    layer1_outputs(4221) <= not (a xor b);
    layer1_outputs(4222) <= not a or b;
    layer1_outputs(4223) <= a and b;
    layer1_outputs(4224) <= not b or a;
    layer1_outputs(4225) <= not (a and b);
    layer1_outputs(4226) <= not a;
    layer1_outputs(4227) <= not a;
    layer1_outputs(4228) <= b and not a;
    layer1_outputs(4229) <= not a or b;
    layer1_outputs(4230) <= a and not b;
    layer1_outputs(4231) <= not a or b;
    layer1_outputs(4232) <= b;
    layer1_outputs(4233) <= a or b;
    layer1_outputs(4234) <= not (a or b);
    layer1_outputs(4235) <= not b;
    layer1_outputs(4236) <= a and not b;
    layer1_outputs(4237) <= not (a xor b);
    layer1_outputs(4238) <= a or b;
    layer1_outputs(4239) <= not a or b;
    layer1_outputs(4240) <= not (a xor b);
    layer1_outputs(4241) <= not b;
    layer1_outputs(4242) <= b and not a;
    layer1_outputs(4243) <= not (a or b);
    layer1_outputs(4244) <= not b;
    layer1_outputs(4245) <= not b;
    layer1_outputs(4246) <= not a;
    layer1_outputs(4247) <= not (a xor b);
    layer1_outputs(4248) <= not a or b;
    layer1_outputs(4249) <= a xor b;
    layer1_outputs(4250) <= not b;
    layer1_outputs(4251) <= not b;
    layer1_outputs(4252) <= a and b;
    layer1_outputs(4253) <= b;
    layer1_outputs(4254) <= not b or a;
    layer1_outputs(4255) <= not b;
    layer1_outputs(4256) <= b;
    layer1_outputs(4257) <= a xor b;
    layer1_outputs(4258) <= not a or b;
    layer1_outputs(4259) <= a;
    layer1_outputs(4260) <= a or b;
    layer1_outputs(4261) <= a and b;
    layer1_outputs(4262) <= a and b;
    layer1_outputs(4263) <= not a;
    layer1_outputs(4264) <= a and not b;
    layer1_outputs(4265) <= b and not a;
    layer1_outputs(4266) <= b;
    layer1_outputs(4267) <= not (a or b);
    layer1_outputs(4268) <= b;
    layer1_outputs(4269) <= not a or b;
    layer1_outputs(4270) <= not a or b;
    layer1_outputs(4271) <= a xor b;
    layer1_outputs(4272) <= b;
    layer1_outputs(4273) <= a and not b;
    layer1_outputs(4274) <= a or b;
    layer1_outputs(4275) <= not a;
    layer1_outputs(4276) <= a xor b;
    layer1_outputs(4277) <= not a;
    layer1_outputs(4278) <= not a;
    layer1_outputs(4279) <= a and not b;
    layer1_outputs(4280) <= not a;
    layer1_outputs(4281) <= not (a xor b);
    layer1_outputs(4282) <= not a or b;
    layer1_outputs(4283) <= a;
    layer1_outputs(4284) <= not b or a;
    layer1_outputs(4285) <= not b;
    layer1_outputs(4286) <= a;
    layer1_outputs(4287) <= a or b;
    layer1_outputs(4288) <= a or b;
    layer1_outputs(4289) <= a;
    layer1_outputs(4290) <= not (a and b);
    layer1_outputs(4291) <= not b;
    layer1_outputs(4292) <= a xor b;
    layer1_outputs(4293) <= not a;
    layer1_outputs(4294) <= not b;
    layer1_outputs(4295) <= not a or b;
    layer1_outputs(4296) <= not a or b;
    layer1_outputs(4297) <= b and not a;
    layer1_outputs(4298) <= a xor b;
    layer1_outputs(4299) <= not (a or b);
    layer1_outputs(4300) <= not (a or b);
    layer1_outputs(4301) <= a and not b;
    layer1_outputs(4302) <= not (a or b);
    layer1_outputs(4303) <= a;
    layer1_outputs(4304) <= not b;
    layer1_outputs(4305) <= not b or a;
    layer1_outputs(4306) <= not b;
    layer1_outputs(4307) <= a;
    layer1_outputs(4308) <= a and not b;
    layer1_outputs(4309) <= a;
    layer1_outputs(4310) <= a;
    layer1_outputs(4311) <= b;
    layer1_outputs(4312) <= a;
    layer1_outputs(4313) <= not a or b;
    layer1_outputs(4314) <= a;
    layer1_outputs(4315) <= b;
    layer1_outputs(4316) <= not (a or b);
    layer1_outputs(4317) <= a;
    layer1_outputs(4318) <= not (a xor b);
    layer1_outputs(4319) <= a xor b;
    layer1_outputs(4320) <= not (a and b);
    layer1_outputs(4321) <= b;
    layer1_outputs(4322) <= a and b;
    layer1_outputs(4323) <= b and not a;
    layer1_outputs(4324) <= not (a xor b);
    layer1_outputs(4325) <= b;
    layer1_outputs(4326) <= a;
    layer1_outputs(4327) <= not b or a;
    layer1_outputs(4328) <= not b;
    layer1_outputs(4329) <= not b;
    layer1_outputs(4330) <= b;
    layer1_outputs(4331) <= not (a xor b);
    layer1_outputs(4332) <= b and not a;
    layer1_outputs(4333) <= a and b;
    layer1_outputs(4334) <= not (a or b);
    layer1_outputs(4335) <= b;
    layer1_outputs(4336) <= not b or a;
    layer1_outputs(4337) <= b and not a;
    layer1_outputs(4338) <= not b;
    layer1_outputs(4339) <= b;
    layer1_outputs(4340) <= b;
    layer1_outputs(4341) <= not b;
    layer1_outputs(4342) <= '0';
    layer1_outputs(4343) <= not (a xor b);
    layer1_outputs(4344) <= a and not b;
    layer1_outputs(4345) <= not b;
    layer1_outputs(4346) <= not a or b;
    layer1_outputs(4347) <= not (a or b);
    layer1_outputs(4348) <= b and not a;
    layer1_outputs(4349) <= not (a xor b);
    layer1_outputs(4350) <= b;
    layer1_outputs(4351) <= not a;
    layer1_outputs(4352) <= a or b;
    layer1_outputs(4353) <= not a;
    layer1_outputs(4354) <= a and not b;
    layer1_outputs(4355) <= not a;
    layer1_outputs(4356) <= not (a or b);
    layer1_outputs(4357) <= not (a xor b);
    layer1_outputs(4358) <= not b or a;
    layer1_outputs(4359) <= not a;
    layer1_outputs(4360) <= b;
    layer1_outputs(4361) <= not (a xor b);
    layer1_outputs(4362) <= not a;
    layer1_outputs(4363) <= a or b;
    layer1_outputs(4364) <= '1';
    layer1_outputs(4365) <= not b or a;
    layer1_outputs(4366) <= not (a and b);
    layer1_outputs(4367) <= not b;
    layer1_outputs(4368) <= not b;
    layer1_outputs(4369) <= '1';
    layer1_outputs(4370) <= '1';
    layer1_outputs(4371) <= not a;
    layer1_outputs(4372) <= not a or b;
    layer1_outputs(4373) <= not a;
    layer1_outputs(4374) <= not (a or b);
    layer1_outputs(4375) <= a and not b;
    layer1_outputs(4376) <= a and b;
    layer1_outputs(4377) <= not (a or b);
    layer1_outputs(4378) <= not (a and b);
    layer1_outputs(4379) <= '0';
    layer1_outputs(4380) <= not b;
    layer1_outputs(4381) <= a;
    layer1_outputs(4382) <= not (a or b);
    layer1_outputs(4383) <= not (a and b);
    layer1_outputs(4384) <= a or b;
    layer1_outputs(4385) <= not a or b;
    layer1_outputs(4386) <= a or b;
    layer1_outputs(4387) <= not b;
    layer1_outputs(4388) <= a;
    layer1_outputs(4389) <= not (a and b);
    layer1_outputs(4390) <= a xor b;
    layer1_outputs(4391) <= not b or a;
    layer1_outputs(4392) <= not b or a;
    layer1_outputs(4393) <= a and b;
    layer1_outputs(4394) <= a and not b;
    layer1_outputs(4395) <= b and not a;
    layer1_outputs(4396) <= a and b;
    layer1_outputs(4397) <= a and not b;
    layer1_outputs(4398) <= not (a and b);
    layer1_outputs(4399) <= b and not a;
    layer1_outputs(4400) <= a xor b;
    layer1_outputs(4401) <= not (a or b);
    layer1_outputs(4402) <= not b;
    layer1_outputs(4403) <= a;
    layer1_outputs(4404) <= b and not a;
    layer1_outputs(4405) <= a xor b;
    layer1_outputs(4406) <= a xor b;
    layer1_outputs(4407) <= a or b;
    layer1_outputs(4408) <= not b or a;
    layer1_outputs(4409) <= not b or a;
    layer1_outputs(4410) <= a and b;
    layer1_outputs(4411) <= a and not b;
    layer1_outputs(4412) <= not (a or b);
    layer1_outputs(4413) <= a;
    layer1_outputs(4414) <= not (a and b);
    layer1_outputs(4415) <= not a or b;
    layer1_outputs(4416) <= b and not a;
    layer1_outputs(4417) <= a and not b;
    layer1_outputs(4418) <= a and not b;
    layer1_outputs(4419) <= a xor b;
    layer1_outputs(4420) <= not a or b;
    layer1_outputs(4421) <= not (a or b);
    layer1_outputs(4422) <= '0';
    layer1_outputs(4423) <= not (a or b);
    layer1_outputs(4424) <= a;
    layer1_outputs(4425) <= not (a or b);
    layer1_outputs(4426) <= a and not b;
    layer1_outputs(4427) <= not a;
    layer1_outputs(4428) <= not (a or b);
    layer1_outputs(4429) <= a;
    layer1_outputs(4430) <= not b;
    layer1_outputs(4431) <= b;
    layer1_outputs(4432) <= a and not b;
    layer1_outputs(4433) <= b and not a;
    layer1_outputs(4434) <= not b or a;
    layer1_outputs(4435) <= a and b;
    layer1_outputs(4436) <= a or b;
    layer1_outputs(4437) <= a;
    layer1_outputs(4438) <= a xor b;
    layer1_outputs(4439) <= '0';
    layer1_outputs(4440) <= b and not a;
    layer1_outputs(4441) <= a xor b;
    layer1_outputs(4442) <= not a or b;
    layer1_outputs(4443) <= a;
    layer1_outputs(4444) <= b and not a;
    layer1_outputs(4445) <= a or b;
    layer1_outputs(4446) <= a and not b;
    layer1_outputs(4447) <= a;
    layer1_outputs(4448) <= not b;
    layer1_outputs(4449) <= not b;
    layer1_outputs(4450) <= a or b;
    layer1_outputs(4451) <= not b or a;
    layer1_outputs(4452) <= a;
    layer1_outputs(4453) <= not (a or b);
    layer1_outputs(4454) <= a xor b;
    layer1_outputs(4455) <= a xor b;
    layer1_outputs(4456) <= a;
    layer1_outputs(4457) <= a xor b;
    layer1_outputs(4458) <= b and not a;
    layer1_outputs(4459) <= a and not b;
    layer1_outputs(4460) <= not b;
    layer1_outputs(4461) <= '0';
    layer1_outputs(4462) <= not b;
    layer1_outputs(4463) <= b;
    layer1_outputs(4464) <= not a;
    layer1_outputs(4465) <= a;
    layer1_outputs(4466) <= a xor b;
    layer1_outputs(4467) <= b;
    layer1_outputs(4468) <= a;
    layer1_outputs(4469) <= not b;
    layer1_outputs(4470) <= not b;
    layer1_outputs(4471) <= not (a xor b);
    layer1_outputs(4472) <= not a;
    layer1_outputs(4473) <= not (a or b);
    layer1_outputs(4474) <= not a;
    layer1_outputs(4475) <= a and b;
    layer1_outputs(4476) <= a;
    layer1_outputs(4477) <= a or b;
    layer1_outputs(4478) <= not a or b;
    layer1_outputs(4479) <= a and not b;
    layer1_outputs(4480) <= b and not a;
    layer1_outputs(4481) <= not (a xor b);
    layer1_outputs(4482) <= not b;
    layer1_outputs(4483) <= b and not a;
    layer1_outputs(4484) <= '1';
    layer1_outputs(4485) <= b;
    layer1_outputs(4486) <= b;
    layer1_outputs(4487) <= not (a xor b);
    layer1_outputs(4488) <= a xor b;
    layer1_outputs(4489) <= not (a xor b);
    layer1_outputs(4490) <= a or b;
    layer1_outputs(4491) <= a;
    layer1_outputs(4492) <= a and not b;
    layer1_outputs(4493) <= not a or b;
    layer1_outputs(4494) <= not (a and b);
    layer1_outputs(4495) <= not (a and b);
    layer1_outputs(4496) <= not (a and b);
    layer1_outputs(4497) <= b and not a;
    layer1_outputs(4498) <= not a;
    layer1_outputs(4499) <= a;
    layer1_outputs(4500) <= not a;
    layer1_outputs(4501) <= a and b;
    layer1_outputs(4502) <= a xor b;
    layer1_outputs(4503) <= a;
    layer1_outputs(4504) <= a or b;
    layer1_outputs(4505) <= a;
    layer1_outputs(4506) <= a xor b;
    layer1_outputs(4507) <= not b or a;
    layer1_outputs(4508) <= a xor b;
    layer1_outputs(4509) <= a and b;
    layer1_outputs(4510) <= a;
    layer1_outputs(4511) <= not (a xor b);
    layer1_outputs(4512) <= a and not b;
    layer1_outputs(4513) <= a or b;
    layer1_outputs(4514) <= a and not b;
    layer1_outputs(4515) <= not a;
    layer1_outputs(4516) <= a;
    layer1_outputs(4517) <= a;
    layer1_outputs(4518) <= not b;
    layer1_outputs(4519) <= a or b;
    layer1_outputs(4520) <= not a or b;
    layer1_outputs(4521) <= a and not b;
    layer1_outputs(4522) <= not (a and b);
    layer1_outputs(4523) <= a;
    layer1_outputs(4524) <= a;
    layer1_outputs(4525) <= a;
    layer1_outputs(4526) <= not (a or b);
    layer1_outputs(4527) <= b and not a;
    layer1_outputs(4528) <= not b or a;
    layer1_outputs(4529) <= b and not a;
    layer1_outputs(4530) <= b;
    layer1_outputs(4531) <= b and not a;
    layer1_outputs(4532) <= a or b;
    layer1_outputs(4533) <= a;
    layer1_outputs(4534) <= not (a or b);
    layer1_outputs(4535) <= b and not a;
    layer1_outputs(4536) <= a and not b;
    layer1_outputs(4537) <= not b;
    layer1_outputs(4538) <= not a or b;
    layer1_outputs(4539) <= a and not b;
    layer1_outputs(4540) <= not a or b;
    layer1_outputs(4541) <= a and b;
    layer1_outputs(4542) <= a xor b;
    layer1_outputs(4543) <= not a or b;
    layer1_outputs(4544) <= a and not b;
    layer1_outputs(4545) <= a xor b;
    layer1_outputs(4546) <= a and not b;
    layer1_outputs(4547) <= not b;
    layer1_outputs(4548) <= not b;
    layer1_outputs(4549) <= a;
    layer1_outputs(4550) <= b;
    layer1_outputs(4551) <= not a or b;
    layer1_outputs(4552) <= not b or a;
    layer1_outputs(4553) <= not b or a;
    layer1_outputs(4554) <= not b or a;
    layer1_outputs(4555) <= a;
    layer1_outputs(4556) <= a;
    layer1_outputs(4557) <= a;
    layer1_outputs(4558) <= b;
    layer1_outputs(4559) <= not b or a;
    layer1_outputs(4560) <= '1';
    layer1_outputs(4561) <= a and not b;
    layer1_outputs(4562) <= not a;
    layer1_outputs(4563) <= a xor b;
    layer1_outputs(4564) <= not b;
    layer1_outputs(4565) <= a;
    layer1_outputs(4566) <= not b or a;
    layer1_outputs(4567) <= a xor b;
    layer1_outputs(4568) <= not a or b;
    layer1_outputs(4569) <= b and not a;
    layer1_outputs(4570) <= not b or a;
    layer1_outputs(4571) <= b;
    layer1_outputs(4572) <= not b;
    layer1_outputs(4573) <= a and not b;
    layer1_outputs(4574) <= a and not b;
    layer1_outputs(4575) <= not b or a;
    layer1_outputs(4576) <= not a or b;
    layer1_outputs(4577) <= not b;
    layer1_outputs(4578) <= a xor b;
    layer1_outputs(4579) <= not a or b;
    layer1_outputs(4580) <= b and not a;
    layer1_outputs(4581) <= b;
    layer1_outputs(4582) <= not a;
    layer1_outputs(4583) <= not (a xor b);
    layer1_outputs(4584) <= a and b;
    layer1_outputs(4585) <= not b or a;
    layer1_outputs(4586) <= not (a and b);
    layer1_outputs(4587) <= not (a or b);
    layer1_outputs(4588) <= not a or b;
    layer1_outputs(4589) <= a xor b;
    layer1_outputs(4590) <= a;
    layer1_outputs(4591) <= not (a and b);
    layer1_outputs(4592) <= b;
    layer1_outputs(4593) <= not a;
    layer1_outputs(4594) <= a and not b;
    layer1_outputs(4595) <= not a or b;
    layer1_outputs(4596) <= a and not b;
    layer1_outputs(4597) <= a;
    layer1_outputs(4598) <= not (a or b);
    layer1_outputs(4599) <= not a;
    layer1_outputs(4600) <= b;
    layer1_outputs(4601) <= b and not a;
    layer1_outputs(4602) <= not (a xor b);
    layer1_outputs(4603) <= b and not a;
    layer1_outputs(4604) <= not b or a;
    layer1_outputs(4605) <= a and not b;
    layer1_outputs(4606) <= b and not a;
    layer1_outputs(4607) <= not (a and b);
    layer1_outputs(4608) <= not b;
    layer1_outputs(4609) <= not b;
    layer1_outputs(4610) <= not (a xor b);
    layer1_outputs(4611) <= a and b;
    layer1_outputs(4612) <= b;
    layer1_outputs(4613) <= not a or b;
    layer1_outputs(4614) <= b;
    layer1_outputs(4615) <= b;
    layer1_outputs(4616) <= a and b;
    layer1_outputs(4617) <= not b;
    layer1_outputs(4618) <= a and not b;
    layer1_outputs(4619) <= not a;
    layer1_outputs(4620) <= a or b;
    layer1_outputs(4621) <= not (a and b);
    layer1_outputs(4622) <= a or b;
    layer1_outputs(4623) <= not (a or b);
    layer1_outputs(4624) <= not b;
    layer1_outputs(4625) <= not a or b;
    layer1_outputs(4626) <= not a;
    layer1_outputs(4627) <= not a or b;
    layer1_outputs(4628) <= not a;
    layer1_outputs(4629) <= '1';
    layer1_outputs(4630) <= a;
    layer1_outputs(4631) <= not a;
    layer1_outputs(4632) <= not (a xor b);
    layer1_outputs(4633) <= not a or b;
    layer1_outputs(4634) <= b and not a;
    layer1_outputs(4635) <= a;
    layer1_outputs(4636) <= a xor b;
    layer1_outputs(4637) <= b;
    layer1_outputs(4638) <= a and not b;
    layer1_outputs(4639) <= not (a xor b);
    layer1_outputs(4640) <= a and not b;
    layer1_outputs(4641) <= a xor b;
    layer1_outputs(4642) <= a;
    layer1_outputs(4643) <= a or b;
    layer1_outputs(4644) <= b;
    layer1_outputs(4645) <= a or b;
    layer1_outputs(4646) <= a and b;
    layer1_outputs(4647) <= a;
    layer1_outputs(4648) <= a and b;
    layer1_outputs(4649) <= not a or b;
    layer1_outputs(4650) <= not a or b;
    layer1_outputs(4651) <= a and b;
    layer1_outputs(4652) <= a or b;
    layer1_outputs(4653) <= a or b;
    layer1_outputs(4654) <= not a;
    layer1_outputs(4655) <= not (a and b);
    layer1_outputs(4656) <= not a or b;
    layer1_outputs(4657) <= not (a xor b);
    layer1_outputs(4658) <= not (a xor b);
    layer1_outputs(4659) <= not (a or b);
    layer1_outputs(4660) <= not (a and b);
    layer1_outputs(4661) <= b and not a;
    layer1_outputs(4662) <= b;
    layer1_outputs(4663) <= not (a xor b);
    layer1_outputs(4664) <= not b;
    layer1_outputs(4665) <= not b or a;
    layer1_outputs(4666) <= a;
    layer1_outputs(4667) <= not b;
    layer1_outputs(4668) <= not b;
    layer1_outputs(4669) <= b and not a;
    layer1_outputs(4670) <= not b;
    layer1_outputs(4671) <= not (a or b);
    layer1_outputs(4672) <= a;
    layer1_outputs(4673) <= not (a or b);
    layer1_outputs(4674) <= not a;
    layer1_outputs(4675) <= not (a or b);
    layer1_outputs(4676) <= b and not a;
    layer1_outputs(4677) <= a xor b;
    layer1_outputs(4678) <= not a;
    layer1_outputs(4679) <= not b;
    layer1_outputs(4680) <= not (a xor b);
    layer1_outputs(4681) <= b and not a;
    layer1_outputs(4682) <= a xor b;
    layer1_outputs(4683) <= not b;
    layer1_outputs(4684) <= b;
    layer1_outputs(4685) <= a xor b;
    layer1_outputs(4686) <= not b or a;
    layer1_outputs(4687) <= a xor b;
    layer1_outputs(4688) <= not (a xor b);
    layer1_outputs(4689) <= b and not a;
    layer1_outputs(4690) <= b and not a;
    layer1_outputs(4691) <= not a or b;
    layer1_outputs(4692) <= b and not a;
    layer1_outputs(4693) <= b;
    layer1_outputs(4694) <= a or b;
    layer1_outputs(4695) <= not b;
    layer1_outputs(4696) <= not a or b;
    layer1_outputs(4697) <= not (a and b);
    layer1_outputs(4698) <= a and b;
    layer1_outputs(4699) <= not a or b;
    layer1_outputs(4700) <= a;
    layer1_outputs(4701) <= b;
    layer1_outputs(4702) <= a and b;
    layer1_outputs(4703) <= a xor b;
    layer1_outputs(4704) <= a;
    layer1_outputs(4705) <= not a or b;
    layer1_outputs(4706) <= not a or b;
    layer1_outputs(4707) <= not (a xor b);
    layer1_outputs(4708) <= not b or a;
    layer1_outputs(4709) <= not a;
    layer1_outputs(4710) <= not (a or b);
    layer1_outputs(4711) <= a and not b;
    layer1_outputs(4712) <= b;
    layer1_outputs(4713) <= a;
    layer1_outputs(4714) <= a xor b;
    layer1_outputs(4715) <= b;
    layer1_outputs(4716) <= not a or b;
    layer1_outputs(4717) <= not b;
    layer1_outputs(4718) <= b;
    layer1_outputs(4719) <= not b;
    layer1_outputs(4720) <= a or b;
    layer1_outputs(4721) <= a xor b;
    layer1_outputs(4722) <= b;
    layer1_outputs(4723) <= a xor b;
    layer1_outputs(4724) <= '0';
    layer1_outputs(4725) <= a;
    layer1_outputs(4726) <= a or b;
    layer1_outputs(4727) <= '1';
    layer1_outputs(4728) <= b;
    layer1_outputs(4729) <= not a or b;
    layer1_outputs(4730) <= a xor b;
    layer1_outputs(4731) <= not b or a;
    layer1_outputs(4732) <= not a or b;
    layer1_outputs(4733) <= a or b;
    layer1_outputs(4734) <= not a;
    layer1_outputs(4735) <= not a or b;
    layer1_outputs(4736) <= not a or b;
    layer1_outputs(4737) <= a xor b;
    layer1_outputs(4738) <= not b;
    layer1_outputs(4739) <= not b or a;
    layer1_outputs(4740) <= b;
    layer1_outputs(4741) <= a;
    layer1_outputs(4742) <= a;
    layer1_outputs(4743) <= not b;
    layer1_outputs(4744) <= a xor b;
    layer1_outputs(4745) <= not (a xor b);
    layer1_outputs(4746) <= a;
    layer1_outputs(4747) <= a and b;
    layer1_outputs(4748) <= a xor b;
    layer1_outputs(4749) <= a and not b;
    layer1_outputs(4750) <= not b;
    layer1_outputs(4751) <= not b;
    layer1_outputs(4752) <= a or b;
    layer1_outputs(4753) <= b;
    layer1_outputs(4754) <= not (a xor b);
    layer1_outputs(4755) <= not (a and b);
    layer1_outputs(4756) <= a xor b;
    layer1_outputs(4757) <= not b;
    layer1_outputs(4758) <= a;
    layer1_outputs(4759) <= a and not b;
    layer1_outputs(4760) <= a and not b;
    layer1_outputs(4761) <= not a or b;
    layer1_outputs(4762) <= not (a or b);
    layer1_outputs(4763) <= b and not a;
    layer1_outputs(4764) <= b and not a;
    layer1_outputs(4765) <= a and b;
    layer1_outputs(4766) <= not a;
    layer1_outputs(4767) <= a and not b;
    layer1_outputs(4768) <= b;
    layer1_outputs(4769) <= a;
    layer1_outputs(4770) <= a xor b;
    layer1_outputs(4771) <= not (a xor b);
    layer1_outputs(4772) <= a and not b;
    layer1_outputs(4773) <= not a;
    layer1_outputs(4774) <= b and not a;
    layer1_outputs(4775) <= not a;
    layer1_outputs(4776) <= a xor b;
    layer1_outputs(4777) <= b and not a;
    layer1_outputs(4778) <= not b;
    layer1_outputs(4779) <= not (a xor b);
    layer1_outputs(4780) <= a and not b;
    layer1_outputs(4781) <= a or b;
    layer1_outputs(4782) <= a xor b;
    layer1_outputs(4783) <= a;
    layer1_outputs(4784) <= not b;
    layer1_outputs(4785) <= a and b;
    layer1_outputs(4786) <= b;
    layer1_outputs(4787) <= not (a xor b);
    layer1_outputs(4788) <= not a;
    layer1_outputs(4789) <= b;
    layer1_outputs(4790) <= a and b;
    layer1_outputs(4791) <= not a or b;
    layer1_outputs(4792) <= a and not b;
    layer1_outputs(4793) <= not b;
    layer1_outputs(4794) <= a xor b;
    layer1_outputs(4795) <= not b;
    layer1_outputs(4796) <= b;
    layer1_outputs(4797) <= not b or a;
    layer1_outputs(4798) <= not b or a;
    layer1_outputs(4799) <= not a;
    layer1_outputs(4800) <= a;
    layer1_outputs(4801) <= not b or a;
    layer1_outputs(4802) <= not b;
    layer1_outputs(4803) <= not b;
    layer1_outputs(4804) <= not (a xor b);
    layer1_outputs(4805) <= not a;
    layer1_outputs(4806) <= not a or b;
    layer1_outputs(4807) <= b;
    layer1_outputs(4808) <= not b;
    layer1_outputs(4809) <= not a;
    layer1_outputs(4810) <= b;
    layer1_outputs(4811) <= a or b;
    layer1_outputs(4812) <= not b;
    layer1_outputs(4813) <= '0';
    layer1_outputs(4814) <= '0';
    layer1_outputs(4815) <= b and not a;
    layer1_outputs(4816) <= b;
    layer1_outputs(4817) <= a or b;
    layer1_outputs(4818) <= a or b;
    layer1_outputs(4819) <= b and not a;
    layer1_outputs(4820) <= not (a and b);
    layer1_outputs(4821) <= a and not b;
    layer1_outputs(4822) <= not b;
    layer1_outputs(4823) <= not a or b;
    layer1_outputs(4824) <= not b;
    layer1_outputs(4825) <= not b or a;
    layer1_outputs(4826) <= a and not b;
    layer1_outputs(4827) <= a and not b;
    layer1_outputs(4828) <= not (a xor b);
    layer1_outputs(4829) <= not b or a;
    layer1_outputs(4830) <= a and b;
    layer1_outputs(4831) <= a;
    layer1_outputs(4832) <= not (a or b);
    layer1_outputs(4833) <= not b;
    layer1_outputs(4834) <= not (a xor b);
    layer1_outputs(4835) <= not b or a;
    layer1_outputs(4836) <= b;
    layer1_outputs(4837) <= a;
    layer1_outputs(4838) <= b;
    layer1_outputs(4839) <= not (a or b);
    layer1_outputs(4840) <= not b or a;
    layer1_outputs(4841) <= a or b;
    layer1_outputs(4842) <= b;
    layer1_outputs(4843) <= a xor b;
    layer1_outputs(4844) <= not a;
    layer1_outputs(4845) <= a or b;
    layer1_outputs(4846) <= not (a xor b);
    layer1_outputs(4847) <= a and b;
    layer1_outputs(4848) <= '1';
    layer1_outputs(4849) <= a and b;
    layer1_outputs(4850) <= not a or b;
    layer1_outputs(4851) <= not a;
    layer1_outputs(4852) <= b;
    layer1_outputs(4853) <= not b or a;
    layer1_outputs(4854) <= not a;
    layer1_outputs(4855) <= b and not a;
    layer1_outputs(4856) <= b;
    layer1_outputs(4857) <= not (a and b);
    layer1_outputs(4858) <= a xor b;
    layer1_outputs(4859) <= b and not a;
    layer1_outputs(4860) <= a and not b;
    layer1_outputs(4861) <= b and not a;
    layer1_outputs(4862) <= not b or a;
    layer1_outputs(4863) <= a and b;
    layer1_outputs(4864) <= a xor b;
    layer1_outputs(4865) <= a or b;
    layer1_outputs(4866) <= not a;
    layer1_outputs(4867) <= not b;
    layer1_outputs(4868) <= b;
    layer1_outputs(4869) <= a and not b;
    layer1_outputs(4870) <= a;
    layer1_outputs(4871) <= a;
    layer1_outputs(4872) <= a xor b;
    layer1_outputs(4873) <= not a;
    layer1_outputs(4874) <= not (a or b);
    layer1_outputs(4875) <= not (a or b);
    layer1_outputs(4876) <= b;
    layer1_outputs(4877) <= a;
    layer1_outputs(4878) <= not b;
    layer1_outputs(4879) <= a;
    layer1_outputs(4880) <= not b;
    layer1_outputs(4881) <= not a;
    layer1_outputs(4882) <= a and b;
    layer1_outputs(4883) <= a;
    layer1_outputs(4884) <= a;
    layer1_outputs(4885) <= a and not b;
    layer1_outputs(4886) <= a and not b;
    layer1_outputs(4887) <= not a or b;
    layer1_outputs(4888) <= a and not b;
    layer1_outputs(4889) <= not a or b;
    layer1_outputs(4890) <= '0';
    layer1_outputs(4891) <= a and not b;
    layer1_outputs(4892) <= a;
    layer1_outputs(4893) <= a xor b;
    layer1_outputs(4894) <= not b;
    layer1_outputs(4895) <= b and not a;
    layer1_outputs(4896) <= not a or b;
    layer1_outputs(4897) <= b and not a;
    layer1_outputs(4898) <= b;
    layer1_outputs(4899) <= not a or b;
    layer1_outputs(4900) <= b;
    layer1_outputs(4901) <= not a;
    layer1_outputs(4902) <= a xor b;
    layer1_outputs(4903) <= not (a and b);
    layer1_outputs(4904) <= a or b;
    layer1_outputs(4905) <= a;
    layer1_outputs(4906) <= a;
    layer1_outputs(4907) <= a;
    layer1_outputs(4908) <= a xor b;
    layer1_outputs(4909) <= not (a and b);
    layer1_outputs(4910) <= a and not b;
    layer1_outputs(4911) <= b;
    layer1_outputs(4912) <= not a;
    layer1_outputs(4913) <= not (a or b);
    layer1_outputs(4914) <= not (a xor b);
    layer1_outputs(4915) <= b;
    layer1_outputs(4916) <= a and b;
    layer1_outputs(4917) <= not (a xor b);
    layer1_outputs(4918) <= not (a xor b);
    layer1_outputs(4919) <= a and b;
    layer1_outputs(4920) <= not a;
    layer1_outputs(4921) <= a and not b;
    layer1_outputs(4922) <= a xor b;
    layer1_outputs(4923) <= not a or b;
    layer1_outputs(4924) <= a and b;
    layer1_outputs(4925) <= b and not a;
    layer1_outputs(4926) <= a;
    layer1_outputs(4927) <= not a or b;
    layer1_outputs(4928) <= not (a and b);
    layer1_outputs(4929) <= a xor b;
    layer1_outputs(4930) <= b and not a;
    layer1_outputs(4931) <= not a or b;
    layer1_outputs(4932) <= a;
    layer1_outputs(4933) <= b;
    layer1_outputs(4934) <= not a or b;
    layer1_outputs(4935) <= b;
    layer1_outputs(4936) <= not (a and b);
    layer1_outputs(4937) <= a and b;
    layer1_outputs(4938) <= a and not b;
    layer1_outputs(4939) <= not (a or b);
    layer1_outputs(4940) <= not a or b;
    layer1_outputs(4941) <= b and not a;
    layer1_outputs(4942) <= not a or b;
    layer1_outputs(4943) <= b and not a;
    layer1_outputs(4944) <= '0';
    layer1_outputs(4945) <= not a or b;
    layer1_outputs(4946) <= not (a xor b);
    layer1_outputs(4947) <= b and not a;
    layer1_outputs(4948) <= a and not b;
    layer1_outputs(4949) <= not (a and b);
    layer1_outputs(4950) <= b;
    layer1_outputs(4951) <= a or b;
    layer1_outputs(4952) <= not (a xor b);
    layer1_outputs(4953) <= a xor b;
    layer1_outputs(4954) <= b;
    layer1_outputs(4955) <= not a;
    layer1_outputs(4956) <= '1';
    layer1_outputs(4957) <= a and not b;
    layer1_outputs(4958) <= not (a and b);
    layer1_outputs(4959) <= a xor b;
    layer1_outputs(4960) <= a and not b;
    layer1_outputs(4961) <= not (a or b);
    layer1_outputs(4962) <= not b;
    layer1_outputs(4963) <= a;
    layer1_outputs(4964) <= not (a and b);
    layer1_outputs(4965) <= b and not a;
    layer1_outputs(4966) <= not b or a;
    layer1_outputs(4967) <= not a or b;
    layer1_outputs(4968) <= not (a and b);
    layer1_outputs(4969) <= not b;
    layer1_outputs(4970) <= b;
    layer1_outputs(4971) <= a or b;
    layer1_outputs(4972) <= a and b;
    layer1_outputs(4973) <= not a;
    layer1_outputs(4974) <= not a or b;
    layer1_outputs(4975) <= not (a and b);
    layer1_outputs(4976) <= a and not b;
    layer1_outputs(4977) <= not (a xor b);
    layer1_outputs(4978) <= not (a and b);
    layer1_outputs(4979) <= not b or a;
    layer1_outputs(4980) <= a or b;
    layer1_outputs(4981) <= b;
    layer1_outputs(4982) <= not (a or b);
    layer1_outputs(4983) <= not (a or b);
    layer1_outputs(4984) <= not b or a;
    layer1_outputs(4985) <= not a or b;
    layer1_outputs(4986) <= b;
    layer1_outputs(4987) <= not b;
    layer1_outputs(4988) <= not a;
    layer1_outputs(4989) <= a or b;
    layer1_outputs(4990) <= not b;
    layer1_outputs(4991) <= not a or b;
    layer1_outputs(4992) <= a or b;
    layer1_outputs(4993) <= b and not a;
    layer1_outputs(4994) <= not (a and b);
    layer1_outputs(4995) <= not a;
    layer1_outputs(4996) <= not a;
    layer1_outputs(4997) <= b;
    layer1_outputs(4998) <= a and b;
    layer1_outputs(4999) <= not (a xor b);
    layer1_outputs(5000) <= a xor b;
    layer1_outputs(5001) <= a and not b;
    layer1_outputs(5002) <= a or b;
    layer1_outputs(5003) <= not (a xor b);
    layer1_outputs(5004) <= b;
    layer1_outputs(5005) <= not (a xor b);
    layer1_outputs(5006) <= not (a and b);
    layer1_outputs(5007) <= b;
    layer1_outputs(5008) <= b;
    layer1_outputs(5009) <= a xor b;
    layer1_outputs(5010) <= not b;
    layer1_outputs(5011) <= not b;
    layer1_outputs(5012) <= not b;
    layer1_outputs(5013) <= not b or a;
    layer1_outputs(5014) <= not (a or b);
    layer1_outputs(5015) <= a xor b;
    layer1_outputs(5016) <= a xor b;
    layer1_outputs(5017) <= not b;
    layer1_outputs(5018) <= not (a and b);
    layer1_outputs(5019) <= b and not a;
    layer1_outputs(5020) <= a or b;
    layer1_outputs(5021) <= not (a and b);
    layer1_outputs(5022) <= not a or b;
    layer1_outputs(5023) <= a xor b;
    layer1_outputs(5024) <= b and not a;
    layer1_outputs(5025) <= b and not a;
    layer1_outputs(5026) <= a xor b;
    layer1_outputs(5027) <= not a;
    layer1_outputs(5028) <= not a;
    layer1_outputs(5029) <= a xor b;
    layer1_outputs(5030) <= b and not a;
    layer1_outputs(5031) <= b and not a;
    layer1_outputs(5032) <= a and b;
    layer1_outputs(5033) <= not a;
    layer1_outputs(5034) <= a xor b;
    layer1_outputs(5035) <= not b or a;
    layer1_outputs(5036) <= not (a and b);
    layer1_outputs(5037) <= not a;
    layer1_outputs(5038) <= a or b;
    layer1_outputs(5039) <= not b;
    layer1_outputs(5040) <= a and not b;
    layer1_outputs(5041) <= b;
    layer1_outputs(5042) <= not a;
    layer1_outputs(5043) <= not (a and b);
    layer1_outputs(5044) <= not a;
    layer1_outputs(5045) <= a and not b;
    layer1_outputs(5046) <= b;
    layer1_outputs(5047) <= a xor b;
    layer1_outputs(5048) <= b and not a;
    layer1_outputs(5049) <= not b;
    layer1_outputs(5050) <= a;
    layer1_outputs(5051) <= not (a or b);
    layer1_outputs(5052) <= b;
    layer1_outputs(5053) <= not b;
    layer1_outputs(5054) <= b;
    layer1_outputs(5055) <= not (a and b);
    layer1_outputs(5056) <= a and b;
    layer1_outputs(5057) <= b;
    layer1_outputs(5058) <= a;
    layer1_outputs(5059) <= not (a and b);
    layer1_outputs(5060) <= a xor b;
    layer1_outputs(5061) <= b;
    layer1_outputs(5062) <= b and not a;
    layer1_outputs(5063) <= a or b;
    layer1_outputs(5064) <= not b;
    layer1_outputs(5065) <= a or b;
    layer1_outputs(5066) <= a or b;
    layer1_outputs(5067) <= not a;
    layer1_outputs(5068) <= a and b;
    layer1_outputs(5069) <= a and not b;
    layer1_outputs(5070) <= a or b;
    layer1_outputs(5071) <= b and not a;
    layer1_outputs(5072) <= not a;
    layer1_outputs(5073) <= not a or b;
    layer1_outputs(5074) <= a and b;
    layer1_outputs(5075) <= a xor b;
    layer1_outputs(5076) <= b and not a;
    layer1_outputs(5077) <= not b;
    layer1_outputs(5078) <= not a;
    layer1_outputs(5079) <= not b or a;
    layer1_outputs(5080) <= b;
    layer1_outputs(5081) <= b;
    layer1_outputs(5082) <= not a;
    layer1_outputs(5083) <= a or b;
    layer1_outputs(5084) <= a and b;
    layer1_outputs(5085) <= '0';
    layer1_outputs(5086) <= not b;
    layer1_outputs(5087) <= not b or a;
    layer1_outputs(5088) <= not a;
    layer1_outputs(5089) <= not (a xor b);
    layer1_outputs(5090) <= not a or b;
    layer1_outputs(5091) <= not a or b;
    layer1_outputs(5092) <= not (a xor b);
    layer1_outputs(5093) <= not a;
    layer1_outputs(5094) <= not (a and b);
    layer1_outputs(5095) <= not b;
    layer1_outputs(5096) <= b and not a;
    layer1_outputs(5097) <= not b or a;
    layer1_outputs(5098) <= not b;
    layer1_outputs(5099) <= not (a or b);
    layer1_outputs(5100) <= a xor b;
    layer1_outputs(5101) <= not b or a;
    layer1_outputs(5102) <= a and b;
    layer1_outputs(5103) <= not (a xor b);
    layer1_outputs(5104) <= not b or a;
    layer1_outputs(5105) <= not b or a;
    layer1_outputs(5106) <= not b;
    layer1_outputs(5107) <= not (a or b);
    layer1_outputs(5108) <= not a;
    layer1_outputs(5109) <= not (a xor b);
    layer1_outputs(5110) <= a or b;
    layer1_outputs(5111) <= not a;
    layer1_outputs(5112) <= a;
    layer1_outputs(5113) <= a xor b;
    layer1_outputs(5114) <= a;
    layer1_outputs(5115) <= not (a xor b);
    layer1_outputs(5116) <= not (a and b);
    layer1_outputs(5117) <= not (a xor b);
    layer1_outputs(5118) <= not b or a;
    layer1_outputs(5119) <= a and b;
    layer1_outputs(5120) <= a xor b;
    layer1_outputs(5121) <= a xor b;
    layer1_outputs(5122) <= not a or b;
    layer1_outputs(5123) <= not (a or b);
    layer1_outputs(5124) <= a and b;
    layer1_outputs(5125) <= not b;
    layer1_outputs(5126) <= a and not b;
    layer1_outputs(5127) <= a;
    layer1_outputs(5128) <= not b or a;
    layer1_outputs(5129) <= a and not b;
    layer1_outputs(5130) <= a and not b;
    layer1_outputs(5131) <= not a;
    layer1_outputs(5132) <= b and not a;
    layer1_outputs(5133) <= a and not b;
    layer1_outputs(5134) <= a and b;
    layer1_outputs(5135) <= '0';
    layer1_outputs(5136) <= b;
    layer1_outputs(5137) <= not a;
    layer1_outputs(5138) <= a and not b;
    layer1_outputs(5139) <= not b;
    layer1_outputs(5140) <= not a;
    layer1_outputs(5141) <= not b or a;
    layer1_outputs(5142) <= b and not a;
    layer1_outputs(5143) <= not b or a;
    layer1_outputs(5144) <= b and not a;
    layer1_outputs(5145) <= b;
    layer1_outputs(5146) <= not a;
    layer1_outputs(5147) <= not (a and b);
    layer1_outputs(5148) <= b;
    layer1_outputs(5149) <= not a or b;
    layer1_outputs(5150) <= not (a and b);
    layer1_outputs(5151) <= not (a or b);
    layer1_outputs(5152) <= a xor b;
    layer1_outputs(5153) <= a and not b;
    layer1_outputs(5154) <= not a or b;
    layer1_outputs(5155) <= a;
    layer1_outputs(5156) <= a or b;
    layer1_outputs(5157) <= b and not a;
    layer1_outputs(5158) <= not b;
    layer1_outputs(5159) <= not a;
    layer1_outputs(5160) <= not (a and b);
    layer1_outputs(5161) <= not (a and b);
    layer1_outputs(5162) <= not a;
    layer1_outputs(5163) <= not b;
    layer1_outputs(5164) <= a and b;
    layer1_outputs(5165) <= not (a xor b);
    layer1_outputs(5166) <= a xor b;
    layer1_outputs(5167) <= not a;
    layer1_outputs(5168) <= not (a or b);
    layer1_outputs(5169) <= a xor b;
    layer1_outputs(5170) <= not (a and b);
    layer1_outputs(5171) <= a xor b;
    layer1_outputs(5172) <= a;
    layer1_outputs(5173) <= b;
    layer1_outputs(5174) <= not a;
    layer1_outputs(5175) <= not (a or b);
    layer1_outputs(5176) <= b and not a;
    layer1_outputs(5177) <= a and not b;
    layer1_outputs(5178) <= not b or a;
    layer1_outputs(5179) <= not a;
    layer1_outputs(5180) <= not a;
    layer1_outputs(5181) <= not b or a;
    layer1_outputs(5182) <= not (a xor b);
    layer1_outputs(5183) <= not b;
    layer1_outputs(5184) <= b;
    layer1_outputs(5185) <= b;
    layer1_outputs(5186) <= a and b;
    layer1_outputs(5187) <= b;
    layer1_outputs(5188) <= a and b;
    layer1_outputs(5189) <= b and not a;
    layer1_outputs(5190) <= a xor b;
    layer1_outputs(5191) <= not (a and b);
    layer1_outputs(5192) <= a and b;
    layer1_outputs(5193) <= '1';
    layer1_outputs(5194) <= a and b;
    layer1_outputs(5195) <= a and b;
    layer1_outputs(5196) <= a or b;
    layer1_outputs(5197) <= a or b;
    layer1_outputs(5198) <= not b;
    layer1_outputs(5199) <= b and not a;
    layer1_outputs(5200) <= a xor b;
    layer1_outputs(5201) <= not a;
    layer1_outputs(5202) <= a;
    layer1_outputs(5203) <= not b;
    layer1_outputs(5204) <= a and not b;
    layer1_outputs(5205) <= a xor b;
    layer1_outputs(5206) <= a and not b;
    layer1_outputs(5207) <= b;
    layer1_outputs(5208) <= not a or b;
    layer1_outputs(5209) <= a and not b;
    layer1_outputs(5210) <= not b or a;
    layer1_outputs(5211) <= b;
    layer1_outputs(5212) <= not b or a;
    layer1_outputs(5213) <= a;
    layer1_outputs(5214) <= a;
    layer1_outputs(5215) <= a;
    layer1_outputs(5216) <= not a or b;
    layer1_outputs(5217) <= not (a or b);
    layer1_outputs(5218) <= a;
    layer1_outputs(5219) <= not a or b;
    layer1_outputs(5220) <= not (a xor b);
    layer1_outputs(5221) <= not (a xor b);
    layer1_outputs(5222) <= not (a xor b);
    layer1_outputs(5223) <= not (a or b);
    layer1_outputs(5224) <= not (a and b);
    layer1_outputs(5225) <= a or b;
    layer1_outputs(5226) <= not a;
    layer1_outputs(5227) <= not b;
    layer1_outputs(5228) <= not (a xor b);
    layer1_outputs(5229) <= not (a or b);
    layer1_outputs(5230) <= a and not b;
    layer1_outputs(5231) <= b;
    layer1_outputs(5232) <= not (a xor b);
    layer1_outputs(5233) <= not (a or b);
    layer1_outputs(5234) <= b;
    layer1_outputs(5235) <= not (a or b);
    layer1_outputs(5236) <= not a or b;
    layer1_outputs(5237) <= not b or a;
    layer1_outputs(5238) <= not b or a;
    layer1_outputs(5239) <= b and not a;
    layer1_outputs(5240) <= not (a xor b);
    layer1_outputs(5241) <= b and not a;
    layer1_outputs(5242) <= a and not b;
    layer1_outputs(5243) <= a and b;
    layer1_outputs(5244) <= a and not b;
    layer1_outputs(5245) <= not a or b;
    layer1_outputs(5246) <= a xor b;
    layer1_outputs(5247) <= a and not b;
    layer1_outputs(5248) <= a and not b;
    layer1_outputs(5249) <= not a or b;
    layer1_outputs(5250) <= a and not b;
    layer1_outputs(5251) <= not (a and b);
    layer1_outputs(5252) <= not a or b;
    layer1_outputs(5253) <= not b;
    layer1_outputs(5254) <= a or b;
    layer1_outputs(5255) <= not (a xor b);
    layer1_outputs(5256) <= not (a or b);
    layer1_outputs(5257) <= not (a xor b);
    layer1_outputs(5258) <= not (a and b);
    layer1_outputs(5259) <= a or b;
    layer1_outputs(5260) <= a and not b;
    layer1_outputs(5261) <= not b;
    layer1_outputs(5262) <= a and b;
    layer1_outputs(5263) <= a or b;
    layer1_outputs(5264) <= not a or b;
    layer1_outputs(5265) <= a and not b;
    layer1_outputs(5266) <= b and not a;
    layer1_outputs(5267) <= not (a xor b);
    layer1_outputs(5268) <= not (a and b);
    layer1_outputs(5269) <= a and not b;
    layer1_outputs(5270) <= b;
    layer1_outputs(5271) <= a xor b;
    layer1_outputs(5272) <= not (a xor b);
    layer1_outputs(5273) <= not b;
    layer1_outputs(5274) <= not b;
    layer1_outputs(5275) <= not (a xor b);
    layer1_outputs(5276) <= b and not a;
    layer1_outputs(5277) <= not (a xor b);
    layer1_outputs(5278) <= not b;
    layer1_outputs(5279) <= not b;
    layer1_outputs(5280) <= not (a xor b);
    layer1_outputs(5281) <= b;
    layer1_outputs(5282) <= a and b;
    layer1_outputs(5283) <= a xor b;
    layer1_outputs(5284) <= not b or a;
    layer1_outputs(5285) <= not b or a;
    layer1_outputs(5286) <= b;
    layer1_outputs(5287) <= not a;
    layer1_outputs(5288) <= b and not a;
    layer1_outputs(5289) <= a or b;
    layer1_outputs(5290) <= not (a and b);
    layer1_outputs(5291) <= a and b;
    layer1_outputs(5292) <= '0';
    layer1_outputs(5293) <= not (a or b);
    layer1_outputs(5294) <= a and not b;
    layer1_outputs(5295) <= b;
    layer1_outputs(5296) <= a or b;
    layer1_outputs(5297) <= a xor b;
    layer1_outputs(5298) <= not (a and b);
    layer1_outputs(5299) <= a and b;
    layer1_outputs(5300) <= a and b;
    layer1_outputs(5301) <= a or b;
    layer1_outputs(5302) <= a and not b;
    layer1_outputs(5303) <= not (a xor b);
    layer1_outputs(5304) <= b;
    layer1_outputs(5305) <= b and not a;
    layer1_outputs(5306) <= not b or a;
    layer1_outputs(5307) <= a xor b;
    layer1_outputs(5308) <= a xor b;
    layer1_outputs(5309) <= a and not b;
    layer1_outputs(5310) <= not (a xor b);
    layer1_outputs(5311) <= not a;
    layer1_outputs(5312) <= not (a and b);
    layer1_outputs(5313) <= a xor b;
    layer1_outputs(5314) <= a;
    layer1_outputs(5315) <= a;
    layer1_outputs(5316) <= not a;
    layer1_outputs(5317) <= a;
    layer1_outputs(5318) <= a and b;
    layer1_outputs(5319) <= not (a or b);
    layer1_outputs(5320) <= a xor b;
    layer1_outputs(5321) <= a;
    layer1_outputs(5322) <= a and not b;
    layer1_outputs(5323) <= b and not a;
    layer1_outputs(5324) <= a;
    layer1_outputs(5325) <= a and not b;
    layer1_outputs(5326) <= not a;
    layer1_outputs(5327) <= a;
    layer1_outputs(5328) <= not (a or b);
    layer1_outputs(5329) <= a;
    layer1_outputs(5330) <= a and not b;
    layer1_outputs(5331) <= not a or b;
    layer1_outputs(5332) <= a xor b;
    layer1_outputs(5333) <= a or b;
    layer1_outputs(5334) <= b;
    layer1_outputs(5335) <= a xor b;
    layer1_outputs(5336) <= not b;
    layer1_outputs(5337) <= not b or a;
    layer1_outputs(5338) <= b;
    layer1_outputs(5339) <= b and not a;
    layer1_outputs(5340) <= b;
    layer1_outputs(5341) <= not a or b;
    layer1_outputs(5342) <= not a;
    layer1_outputs(5343) <= not (a and b);
    layer1_outputs(5344) <= not a;
    layer1_outputs(5345) <= b;
    layer1_outputs(5346) <= a xor b;
    layer1_outputs(5347) <= a or b;
    layer1_outputs(5348) <= a xor b;
    layer1_outputs(5349) <= b;
    layer1_outputs(5350) <= not (a and b);
    layer1_outputs(5351) <= not b;
    layer1_outputs(5352) <= not (a or b);
    layer1_outputs(5353) <= not (a or b);
    layer1_outputs(5354) <= a;
    layer1_outputs(5355) <= b;
    layer1_outputs(5356) <= a xor b;
    layer1_outputs(5357) <= not a;
    layer1_outputs(5358) <= a xor b;
    layer1_outputs(5359) <= b and not a;
    layer1_outputs(5360) <= a;
    layer1_outputs(5361) <= '0';
    layer1_outputs(5362) <= not a;
    layer1_outputs(5363) <= a;
    layer1_outputs(5364) <= a and b;
    layer1_outputs(5365) <= not (a and b);
    layer1_outputs(5366) <= a;
    layer1_outputs(5367) <= b and not a;
    layer1_outputs(5368) <= not b;
    layer1_outputs(5369) <= a;
    layer1_outputs(5370) <= not a or b;
    layer1_outputs(5371) <= b and not a;
    layer1_outputs(5372) <= not (a and b);
    layer1_outputs(5373) <= not b;
    layer1_outputs(5374) <= not (a xor b);
    layer1_outputs(5375) <= not a or b;
    layer1_outputs(5376) <= not a or b;
    layer1_outputs(5377) <= a;
    layer1_outputs(5378) <= not a or b;
    layer1_outputs(5379) <= a xor b;
    layer1_outputs(5380) <= a or b;
    layer1_outputs(5381) <= b;
    layer1_outputs(5382) <= a or b;
    layer1_outputs(5383) <= a and b;
    layer1_outputs(5384) <= not a or b;
    layer1_outputs(5385) <= a xor b;
    layer1_outputs(5386) <= not (a and b);
    layer1_outputs(5387) <= a;
    layer1_outputs(5388) <= b;
    layer1_outputs(5389) <= not (a xor b);
    layer1_outputs(5390) <= not (a xor b);
    layer1_outputs(5391) <= not b;
    layer1_outputs(5392) <= b;
    layer1_outputs(5393) <= not (a xor b);
    layer1_outputs(5394) <= not a or b;
    layer1_outputs(5395) <= a and b;
    layer1_outputs(5396) <= not a or b;
    layer1_outputs(5397) <= a and not b;
    layer1_outputs(5398) <= a;
    layer1_outputs(5399) <= not a;
    layer1_outputs(5400) <= not a or b;
    layer1_outputs(5401) <= not (a and b);
    layer1_outputs(5402) <= not a;
    layer1_outputs(5403) <= not (a xor b);
    layer1_outputs(5404) <= not a or b;
    layer1_outputs(5405) <= not (a or b);
    layer1_outputs(5406) <= not (a and b);
    layer1_outputs(5407) <= b;
    layer1_outputs(5408) <= not b;
    layer1_outputs(5409) <= not b;
    layer1_outputs(5410) <= a xor b;
    layer1_outputs(5411) <= a and b;
    layer1_outputs(5412) <= not (a xor b);
    layer1_outputs(5413) <= a and not b;
    layer1_outputs(5414) <= not a;
    layer1_outputs(5415) <= a and not b;
    layer1_outputs(5416) <= a and b;
    layer1_outputs(5417) <= a or b;
    layer1_outputs(5418) <= not a or b;
    layer1_outputs(5419) <= a;
    layer1_outputs(5420) <= b and not a;
    layer1_outputs(5421) <= not b;
    layer1_outputs(5422) <= a or b;
    layer1_outputs(5423) <= not a or b;
    layer1_outputs(5424) <= a and not b;
    layer1_outputs(5425) <= not (a or b);
    layer1_outputs(5426) <= a xor b;
    layer1_outputs(5427) <= not a;
    layer1_outputs(5428) <= not a or b;
    layer1_outputs(5429) <= not b;
    layer1_outputs(5430) <= not (a xor b);
    layer1_outputs(5431) <= a xor b;
    layer1_outputs(5432) <= a xor b;
    layer1_outputs(5433) <= not b;
    layer1_outputs(5434) <= not (a xor b);
    layer1_outputs(5435) <= a and b;
    layer1_outputs(5436) <= b and not a;
    layer1_outputs(5437) <= a or b;
    layer1_outputs(5438) <= not (a and b);
    layer1_outputs(5439) <= a and not b;
    layer1_outputs(5440) <= not a or b;
    layer1_outputs(5441) <= not b;
    layer1_outputs(5442) <= a or b;
    layer1_outputs(5443) <= b;
    layer1_outputs(5444) <= a;
    layer1_outputs(5445) <= a and not b;
    layer1_outputs(5446) <= not (a and b);
    layer1_outputs(5447) <= b and not a;
    layer1_outputs(5448) <= not (a and b);
    layer1_outputs(5449) <= a xor b;
    layer1_outputs(5450) <= not (a or b);
    layer1_outputs(5451) <= a or b;
    layer1_outputs(5452) <= not a;
    layer1_outputs(5453) <= not b;
    layer1_outputs(5454) <= not (a and b);
    layer1_outputs(5455) <= not b or a;
    layer1_outputs(5456) <= not b or a;
    layer1_outputs(5457) <= a and b;
    layer1_outputs(5458) <= not (a and b);
    layer1_outputs(5459) <= a or b;
    layer1_outputs(5460) <= a and b;
    layer1_outputs(5461) <= b;
    layer1_outputs(5462) <= b and not a;
    layer1_outputs(5463) <= a or b;
    layer1_outputs(5464) <= '0';
    layer1_outputs(5465) <= a or b;
    layer1_outputs(5466) <= not a or b;
    layer1_outputs(5467) <= a or b;
    layer1_outputs(5468) <= a and not b;
    layer1_outputs(5469) <= not (a xor b);
    layer1_outputs(5470) <= not b or a;
    layer1_outputs(5471) <= not (a or b);
    layer1_outputs(5472) <= a and not b;
    layer1_outputs(5473) <= '1';
    layer1_outputs(5474) <= not a or b;
    layer1_outputs(5475) <= b;
    layer1_outputs(5476) <= a xor b;
    layer1_outputs(5477) <= not (a and b);
    layer1_outputs(5478) <= a;
    layer1_outputs(5479) <= not b or a;
    layer1_outputs(5480) <= not b or a;
    layer1_outputs(5481) <= a and not b;
    layer1_outputs(5482) <= a;
    layer1_outputs(5483) <= not (a and b);
    layer1_outputs(5484) <= not a or b;
    layer1_outputs(5485) <= not (a or b);
    layer1_outputs(5486) <= not b;
    layer1_outputs(5487) <= a and not b;
    layer1_outputs(5488) <= not b or a;
    layer1_outputs(5489) <= not b or a;
    layer1_outputs(5490) <= b;
    layer1_outputs(5491) <= not b or a;
    layer1_outputs(5492) <= a;
    layer1_outputs(5493) <= not b or a;
    layer1_outputs(5494) <= a and b;
    layer1_outputs(5495) <= not b;
    layer1_outputs(5496) <= not (a or b);
    layer1_outputs(5497) <= not a;
    layer1_outputs(5498) <= b;
    layer1_outputs(5499) <= not a or b;
    layer1_outputs(5500) <= not b;
    layer1_outputs(5501) <= a and not b;
    layer1_outputs(5502) <= a or b;
    layer1_outputs(5503) <= not b;
    layer1_outputs(5504) <= b;
    layer1_outputs(5505) <= a or b;
    layer1_outputs(5506) <= not (a and b);
    layer1_outputs(5507) <= a and not b;
    layer1_outputs(5508) <= not b or a;
    layer1_outputs(5509) <= not a;
    layer1_outputs(5510) <= not (a or b);
    layer1_outputs(5511) <= not (a xor b);
    layer1_outputs(5512) <= not (a xor b);
    layer1_outputs(5513) <= not (a or b);
    layer1_outputs(5514) <= not b or a;
    layer1_outputs(5515) <= a and b;
    layer1_outputs(5516) <= not (a or b);
    layer1_outputs(5517) <= not a or b;
    layer1_outputs(5518) <= not (a xor b);
    layer1_outputs(5519) <= a xor b;
    layer1_outputs(5520) <= a and not b;
    layer1_outputs(5521) <= a or b;
    layer1_outputs(5522) <= not a;
    layer1_outputs(5523) <= a;
    layer1_outputs(5524) <= a and b;
    layer1_outputs(5525) <= a and b;
    layer1_outputs(5526) <= '0';
    layer1_outputs(5527) <= a and not b;
    layer1_outputs(5528) <= a;
    layer1_outputs(5529) <= b;
    layer1_outputs(5530) <= a;
    layer1_outputs(5531) <= b;
    layer1_outputs(5532) <= a and b;
    layer1_outputs(5533) <= a and b;
    layer1_outputs(5534) <= a and b;
    layer1_outputs(5535) <= a xor b;
    layer1_outputs(5536) <= a;
    layer1_outputs(5537) <= b;
    layer1_outputs(5538) <= not (a and b);
    layer1_outputs(5539) <= a and b;
    layer1_outputs(5540) <= not a;
    layer1_outputs(5541) <= not b;
    layer1_outputs(5542) <= not (a or b);
    layer1_outputs(5543) <= not a or b;
    layer1_outputs(5544) <= a xor b;
    layer1_outputs(5545) <= a;
    layer1_outputs(5546) <= not a;
    layer1_outputs(5547) <= not (a or b);
    layer1_outputs(5548) <= '0';
    layer1_outputs(5549) <= not a or b;
    layer1_outputs(5550) <= a;
    layer1_outputs(5551) <= not b or a;
    layer1_outputs(5552) <= b and not a;
    layer1_outputs(5553) <= b and not a;
    layer1_outputs(5554) <= a and not b;
    layer1_outputs(5555) <= not (a xor b);
    layer1_outputs(5556) <= not (a or b);
    layer1_outputs(5557) <= a;
    layer1_outputs(5558) <= not b or a;
    layer1_outputs(5559) <= not (a and b);
    layer1_outputs(5560) <= not b or a;
    layer1_outputs(5561) <= not a;
    layer1_outputs(5562) <= a and not b;
    layer1_outputs(5563) <= not (a xor b);
    layer1_outputs(5564) <= not (a and b);
    layer1_outputs(5565) <= a xor b;
    layer1_outputs(5566) <= a and b;
    layer1_outputs(5567) <= not (a or b);
    layer1_outputs(5568) <= a xor b;
    layer1_outputs(5569) <= not (a xor b);
    layer1_outputs(5570) <= not (a xor b);
    layer1_outputs(5571) <= not a;
    layer1_outputs(5572) <= a and not b;
    layer1_outputs(5573) <= not b;
    layer1_outputs(5574) <= b and not a;
    layer1_outputs(5575) <= a or b;
    layer1_outputs(5576) <= not a or b;
    layer1_outputs(5577) <= not a;
    layer1_outputs(5578) <= not b or a;
    layer1_outputs(5579) <= not (a or b);
    layer1_outputs(5580) <= a and b;
    layer1_outputs(5581) <= not b;
    layer1_outputs(5582) <= not (a or b);
    layer1_outputs(5583) <= b;
    layer1_outputs(5584) <= a and not b;
    layer1_outputs(5585) <= b;
    layer1_outputs(5586) <= b and not a;
    layer1_outputs(5587) <= not (a or b);
    layer1_outputs(5588) <= a and b;
    layer1_outputs(5589) <= b and not a;
    layer1_outputs(5590) <= not b;
    layer1_outputs(5591) <= b;
    layer1_outputs(5592) <= not b or a;
    layer1_outputs(5593) <= not a;
    layer1_outputs(5594) <= not a;
    layer1_outputs(5595) <= b;
    layer1_outputs(5596) <= b;
    layer1_outputs(5597) <= a and b;
    layer1_outputs(5598) <= not b;
    layer1_outputs(5599) <= b and not a;
    layer1_outputs(5600) <= a or b;
    layer1_outputs(5601) <= a;
    layer1_outputs(5602) <= not a;
    layer1_outputs(5603) <= not (a and b);
    layer1_outputs(5604) <= b;
    layer1_outputs(5605) <= not a or b;
    layer1_outputs(5606) <= b;
    layer1_outputs(5607) <= a;
    layer1_outputs(5608) <= b and not a;
    layer1_outputs(5609) <= not b;
    layer1_outputs(5610) <= b and not a;
    layer1_outputs(5611) <= not b;
    layer1_outputs(5612) <= a xor b;
    layer1_outputs(5613) <= a;
    layer1_outputs(5614) <= not b or a;
    layer1_outputs(5615) <= b and not a;
    layer1_outputs(5616) <= a;
    layer1_outputs(5617) <= b and not a;
    layer1_outputs(5618) <= b;
    layer1_outputs(5619) <= not b;
    layer1_outputs(5620) <= not (a or b);
    layer1_outputs(5621) <= not a;
    layer1_outputs(5622) <= a and b;
    layer1_outputs(5623) <= b;
    layer1_outputs(5624) <= not b;
    layer1_outputs(5625) <= a and not b;
    layer1_outputs(5626) <= not (a or b);
    layer1_outputs(5627) <= a;
    layer1_outputs(5628) <= not a or b;
    layer1_outputs(5629) <= a and b;
    layer1_outputs(5630) <= not a or b;
    layer1_outputs(5631) <= a and not b;
    layer1_outputs(5632) <= not (a and b);
    layer1_outputs(5633) <= a xor b;
    layer1_outputs(5634) <= b and not a;
    layer1_outputs(5635) <= not (a xor b);
    layer1_outputs(5636) <= a xor b;
    layer1_outputs(5637) <= a;
    layer1_outputs(5638) <= not (a and b);
    layer1_outputs(5639) <= not a or b;
    layer1_outputs(5640) <= a xor b;
    layer1_outputs(5641) <= not (a xor b);
    layer1_outputs(5642) <= a xor b;
    layer1_outputs(5643) <= a xor b;
    layer1_outputs(5644) <= not (a and b);
    layer1_outputs(5645) <= a or b;
    layer1_outputs(5646) <= not a;
    layer1_outputs(5647) <= not b;
    layer1_outputs(5648) <= a xor b;
    layer1_outputs(5649) <= not b;
    layer1_outputs(5650) <= not b or a;
    layer1_outputs(5651) <= not a;
    layer1_outputs(5652) <= not (a or b);
    layer1_outputs(5653) <= not (a and b);
    layer1_outputs(5654) <= a and not b;
    layer1_outputs(5655) <= a or b;
    layer1_outputs(5656) <= b;
    layer1_outputs(5657) <= b;
    layer1_outputs(5658) <= b;
    layer1_outputs(5659) <= not (a xor b);
    layer1_outputs(5660) <= b and not a;
    layer1_outputs(5661) <= not a;
    layer1_outputs(5662) <= a xor b;
    layer1_outputs(5663) <= a xor b;
    layer1_outputs(5664) <= a;
    layer1_outputs(5665) <= not b or a;
    layer1_outputs(5666) <= a xor b;
    layer1_outputs(5667) <= not a or b;
    layer1_outputs(5668) <= b and not a;
    layer1_outputs(5669) <= a xor b;
    layer1_outputs(5670) <= b and not a;
    layer1_outputs(5671) <= not (a xor b);
    layer1_outputs(5672) <= a;
    layer1_outputs(5673) <= not (a or b);
    layer1_outputs(5674) <= b and not a;
    layer1_outputs(5675) <= not (a or b);
    layer1_outputs(5676) <= a xor b;
    layer1_outputs(5677) <= a and b;
    layer1_outputs(5678) <= a;
    layer1_outputs(5679) <= a;
    layer1_outputs(5680) <= b;
    layer1_outputs(5681) <= not a;
    layer1_outputs(5682) <= a xor b;
    layer1_outputs(5683) <= not (a xor b);
    layer1_outputs(5684) <= not b;
    layer1_outputs(5685) <= not a or b;
    layer1_outputs(5686) <= a and b;
    layer1_outputs(5687) <= not a;
    layer1_outputs(5688) <= b and not a;
    layer1_outputs(5689) <= not (a and b);
    layer1_outputs(5690) <= a or b;
    layer1_outputs(5691) <= not a or b;
    layer1_outputs(5692) <= b and not a;
    layer1_outputs(5693) <= b;
    layer1_outputs(5694) <= not b or a;
    layer1_outputs(5695) <= b;
    layer1_outputs(5696) <= a xor b;
    layer1_outputs(5697) <= b;
    layer1_outputs(5698) <= not b;
    layer1_outputs(5699) <= not b or a;
    layer1_outputs(5700) <= b;
    layer1_outputs(5701) <= not (a xor b);
    layer1_outputs(5702) <= not (a xor b);
    layer1_outputs(5703) <= b and not a;
    layer1_outputs(5704) <= not a;
    layer1_outputs(5705) <= not (a or b);
    layer1_outputs(5706) <= a;
    layer1_outputs(5707) <= not (a xor b);
    layer1_outputs(5708) <= a and not b;
    layer1_outputs(5709) <= not (a xor b);
    layer1_outputs(5710) <= b;
    layer1_outputs(5711) <= not b;
    layer1_outputs(5712) <= a and not b;
    layer1_outputs(5713) <= not (a and b);
    layer1_outputs(5714) <= b;
    layer1_outputs(5715) <= not a or b;
    layer1_outputs(5716) <= a;
    layer1_outputs(5717) <= b;
    layer1_outputs(5718) <= a;
    layer1_outputs(5719) <= not (a or b);
    layer1_outputs(5720) <= not (a or b);
    layer1_outputs(5721) <= not b;
    layer1_outputs(5722) <= b;
    layer1_outputs(5723) <= b;
    layer1_outputs(5724) <= a xor b;
    layer1_outputs(5725) <= b;
    layer1_outputs(5726) <= a;
    layer1_outputs(5727) <= a and not b;
    layer1_outputs(5728) <= not (a or b);
    layer1_outputs(5729) <= not (a xor b);
    layer1_outputs(5730) <= '0';
    layer1_outputs(5731) <= a xor b;
    layer1_outputs(5732) <= a and not b;
    layer1_outputs(5733) <= not a;
    layer1_outputs(5734) <= a;
    layer1_outputs(5735) <= a and not b;
    layer1_outputs(5736) <= not a;
    layer1_outputs(5737) <= a and b;
    layer1_outputs(5738) <= a or b;
    layer1_outputs(5739) <= a xor b;
    layer1_outputs(5740) <= not (a xor b);
    layer1_outputs(5741) <= not (a xor b);
    layer1_outputs(5742) <= a;
    layer1_outputs(5743) <= a;
    layer1_outputs(5744) <= not a or b;
    layer1_outputs(5745) <= not (a xor b);
    layer1_outputs(5746) <= not b;
    layer1_outputs(5747) <= a or b;
    layer1_outputs(5748) <= not (a or b);
    layer1_outputs(5749) <= not b or a;
    layer1_outputs(5750) <= a;
    layer1_outputs(5751) <= a;
    layer1_outputs(5752) <= not b or a;
    layer1_outputs(5753) <= a;
    layer1_outputs(5754) <= b;
    layer1_outputs(5755) <= not a;
    layer1_outputs(5756) <= not b;
    layer1_outputs(5757) <= not (a or b);
    layer1_outputs(5758) <= a;
    layer1_outputs(5759) <= a or b;
    layer1_outputs(5760) <= a or b;
    layer1_outputs(5761) <= a or b;
    layer1_outputs(5762) <= not a or b;
    layer1_outputs(5763) <= not (a xor b);
    layer1_outputs(5764) <= not (a xor b);
    layer1_outputs(5765) <= b;
    layer1_outputs(5766) <= not (a and b);
    layer1_outputs(5767) <= not (a and b);
    layer1_outputs(5768) <= a and b;
    layer1_outputs(5769) <= not a;
    layer1_outputs(5770) <= not b;
    layer1_outputs(5771) <= a or b;
    layer1_outputs(5772) <= not a;
    layer1_outputs(5773) <= '1';
    layer1_outputs(5774) <= b;
    layer1_outputs(5775) <= '1';
    layer1_outputs(5776) <= not a;
    layer1_outputs(5777) <= b;
    layer1_outputs(5778) <= a or b;
    layer1_outputs(5779) <= b;
    layer1_outputs(5780) <= not b or a;
    layer1_outputs(5781) <= not a or b;
    layer1_outputs(5782) <= a and not b;
    layer1_outputs(5783) <= a xor b;
    layer1_outputs(5784) <= not (a or b);
    layer1_outputs(5785) <= not b or a;
    layer1_outputs(5786) <= not (a xor b);
    layer1_outputs(5787) <= not a;
    layer1_outputs(5788) <= not b;
    layer1_outputs(5789) <= b;
    layer1_outputs(5790) <= b and not a;
    layer1_outputs(5791) <= a;
    layer1_outputs(5792) <= a xor b;
    layer1_outputs(5793) <= not (a and b);
    layer1_outputs(5794) <= not (a xor b);
    layer1_outputs(5795) <= a xor b;
    layer1_outputs(5796) <= not (a or b);
    layer1_outputs(5797) <= b;
    layer1_outputs(5798) <= b and not a;
    layer1_outputs(5799) <= a and not b;
    layer1_outputs(5800) <= not a or b;
    layer1_outputs(5801) <= a or b;
    layer1_outputs(5802) <= a xor b;
    layer1_outputs(5803) <= b;
    layer1_outputs(5804) <= b and not a;
    layer1_outputs(5805) <= b and not a;
    layer1_outputs(5806) <= not b or a;
    layer1_outputs(5807) <= not (a xor b);
    layer1_outputs(5808) <= a and not b;
    layer1_outputs(5809) <= a;
    layer1_outputs(5810) <= not (a and b);
    layer1_outputs(5811) <= not a;
    layer1_outputs(5812) <= not (a xor b);
    layer1_outputs(5813) <= not (a or b);
    layer1_outputs(5814) <= not (a or b);
    layer1_outputs(5815) <= b;
    layer1_outputs(5816) <= a;
    layer1_outputs(5817) <= not (a and b);
    layer1_outputs(5818) <= not b;
    layer1_outputs(5819) <= a;
    layer1_outputs(5820) <= not a or b;
    layer1_outputs(5821) <= not (a or b);
    layer1_outputs(5822) <= a and b;
    layer1_outputs(5823) <= a xor b;
    layer1_outputs(5824) <= a or b;
    layer1_outputs(5825) <= b;
    layer1_outputs(5826) <= a;
    layer1_outputs(5827) <= a and not b;
    layer1_outputs(5828) <= not a or b;
    layer1_outputs(5829) <= b;
    layer1_outputs(5830) <= not b;
    layer1_outputs(5831) <= not b or a;
    layer1_outputs(5832) <= b and not a;
    layer1_outputs(5833) <= b;
    layer1_outputs(5834) <= not a;
    layer1_outputs(5835) <= a and b;
    layer1_outputs(5836) <= a;
    layer1_outputs(5837) <= b and not a;
    layer1_outputs(5838) <= b;
    layer1_outputs(5839) <= a;
    layer1_outputs(5840) <= a xor b;
    layer1_outputs(5841) <= not (a or b);
    layer1_outputs(5842) <= b and not a;
    layer1_outputs(5843) <= b;
    layer1_outputs(5844) <= a or b;
    layer1_outputs(5845) <= not (a xor b);
    layer1_outputs(5846) <= a;
    layer1_outputs(5847) <= a or b;
    layer1_outputs(5848) <= not a;
    layer1_outputs(5849) <= b and not a;
    layer1_outputs(5850) <= not (a or b);
    layer1_outputs(5851) <= not b or a;
    layer1_outputs(5852) <= a and b;
    layer1_outputs(5853) <= a or b;
    layer1_outputs(5854) <= not (a and b);
    layer1_outputs(5855) <= b and not a;
    layer1_outputs(5856) <= not a or b;
    layer1_outputs(5857) <= b and not a;
    layer1_outputs(5858) <= b;
    layer1_outputs(5859) <= not a or b;
    layer1_outputs(5860) <= not (a and b);
    layer1_outputs(5861) <= not b;
    layer1_outputs(5862) <= not b;
    layer1_outputs(5863) <= not (a xor b);
    layer1_outputs(5864) <= not b or a;
    layer1_outputs(5865) <= a and b;
    layer1_outputs(5866) <= b and not a;
    layer1_outputs(5867) <= a or b;
    layer1_outputs(5868) <= a and not b;
    layer1_outputs(5869) <= not a or b;
    layer1_outputs(5870) <= a and not b;
    layer1_outputs(5871) <= a and b;
    layer1_outputs(5872) <= '0';
    layer1_outputs(5873) <= a and b;
    layer1_outputs(5874) <= not a;
    layer1_outputs(5875) <= not (a and b);
    layer1_outputs(5876) <= not (a or b);
    layer1_outputs(5877) <= not a or b;
    layer1_outputs(5878) <= a;
    layer1_outputs(5879) <= not (a or b);
    layer1_outputs(5880) <= a and b;
    layer1_outputs(5881) <= not b;
    layer1_outputs(5882) <= not b or a;
    layer1_outputs(5883) <= not b;
    layer1_outputs(5884) <= not b;
    layer1_outputs(5885) <= a and b;
    layer1_outputs(5886) <= not b;
    layer1_outputs(5887) <= not b;
    layer1_outputs(5888) <= a or b;
    layer1_outputs(5889) <= a;
    layer1_outputs(5890) <= not b;
    layer1_outputs(5891) <= not a;
    layer1_outputs(5892) <= not (a or b);
    layer1_outputs(5893) <= a and b;
    layer1_outputs(5894) <= not a or b;
    layer1_outputs(5895) <= b;
    layer1_outputs(5896) <= not b;
    layer1_outputs(5897) <= a and b;
    layer1_outputs(5898) <= not b;
    layer1_outputs(5899) <= b;
    layer1_outputs(5900) <= b;
    layer1_outputs(5901) <= a and b;
    layer1_outputs(5902) <= a xor b;
    layer1_outputs(5903) <= not (a xor b);
    layer1_outputs(5904) <= b;
    layer1_outputs(5905) <= a;
    layer1_outputs(5906) <= not b;
    layer1_outputs(5907) <= a and b;
    layer1_outputs(5908) <= b and not a;
    layer1_outputs(5909) <= b and not a;
    layer1_outputs(5910) <= b;
    layer1_outputs(5911) <= not (a and b);
    layer1_outputs(5912) <= not b;
    layer1_outputs(5913) <= not a;
    layer1_outputs(5914) <= a and b;
    layer1_outputs(5915) <= a;
    layer1_outputs(5916) <= a and not b;
    layer1_outputs(5917) <= b;
    layer1_outputs(5918) <= not (a or b);
    layer1_outputs(5919) <= not (a or b);
    layer1_outputs(5920) <= a;
    layer1_outputs(5921) <= not (a xor b);
    layer1_outputs(5922) <= a and b;
    layer1_outputs(5923) <= a and b;
    layer1_outputs(5924) <= not a;
    layer1_outputs(5925) <= a;
    layer1_outputs(5926) <= not b;
    layer1_outputs(5927) <= '0';
    layer1_outputs(5928) <= a or b;
    layer1_outputs(5929) <= not a;
    layer1_outputs(5930) <= not b or a;
    layer1_outputs(5931) <= a or b;
    layer1_outputs(5932) <= b;
    layer1_outputs(5933) <= not b;
    layer1_outputs(5934) <= b;
    layer1_outputs(5935) <= not (a xor b);
    layer1_outputs(5936) <= not b or a;
    layer1_outputs(5937) <= a and b;
    layer1_outputs(5938) <= a and not b;
    layer1_outputs(5939) <= a xor b;
    layer1_outputs(5940) <= not a;
    layer1_outputs(5941) <= a xor b;
    layer1_outputs(5942) <= b and not a;
    layer1_outputs(5943) <= not a;
    layer1_outputs(5944) <= not a;
    layer1_outputs(5945) <= a xor b;
    layer1_outputs(5946) <= a or b;
    layer1_outputs(5947) <= a xor b;
    layer1_outputs(5948) <= not (a and b);
    layer1_outputs(5949) <= b and not a;
    layer1_outputs(5950) <= not a or b;
    layer1_outputs(5951) <= a or b;
    layer1_outputs(5952) <= not b;
    layer1_outputs(5953) <= not a or b;
    layer1_outputs(5954) <= not b or a;
    layer1_outputs(5955) <= b and not a;
    layer1_outputs(5956) <= a and not b;
    layer1_outputs(5957) <= not a or b;
    layer1_outputs(5958) <= a and not b;
    layer1_outputs(5959) <= not b or a;
    layer1_outputs(5960) <= a and b;
    layer1_outputs(5961) <= a xor b;
    layer1_outputs(5962) <= not a or b;
    layer1_outputs(5963) <= b;
    layer1_outputs(5964) <= a xor b;
    layer1_outputs(5965) <= not a;
    layer1_outputs(5966) <= b and not a;
    layer1_outputs(5967) <= not a;
    layer1_outputs(5968) <= a;
    layer1_outputs(5969) <= a xor b;
    layer1_outputs(5970) <= not a;
    layer1_outputs(5971) <= a and b;
    layer1_outputs(5972) <= a and b;
    layer1_outputs(5973) <= b and not a;
    layer1_outputs(5974) <= a and b;
    layer1_outputs(5975) <= a and not b;
    layer1_outputs(5976) <= a or b;
    layer1_outputs(5977) <= b and not a;
    layer1_outputs(5978) <= a and not b;
    layer1_outputs(5979) <= b and not a;
    layer1_outputs(5980) <= a and b;
    layer1_outputs(5981) <= a xor b;
    layer1_outputs(5982) <= not (a xor b);
    layer1_outputs(5983) <= b and not a;
    layer1_outputs(5984) <= not b or a;
    layer1_outputs(5985) <= a or b;
    layer1_outputs(5986) <= a and b;
    layer1_outputs(5987) <= not (a and b);
    layer1_outputs(5988) <= '1';
    layer1_outputs(5989) <= a;
    layer1_outputs(5990) <= not a;
    layer1_outputs(5991) <= not a;
    layer1_outputs(5992) <= a and not b;
    layer1_outputs(5993) <= not a or b;
    layer1_outputs(5994) <= b;
    layer1_outputs(5995) <= not a;
    layer1_outputs(5996) <= not (a or b);
    layer1_outputs(5997) <= not a;
    layer1_outputs(5998) <= a xor b;
    layer1_outputs(5999) <= not b;
    layer1_outputs(6000) <= a and b;
    layer1_outputs(6001) <= '0';
    layer1_outputs(6002) <= not (a and b);
    layer1_outputs(6003) <= not b;
    layer1_outputs(6004) <= a;
    layer1_outputs(6005) <= b and not a;
    layer1_outputs(6006) <= not a;
    layer1_outputs(6007) <= b and not a;
    layer1_outputs(6008) <= a and not b;
    layer1_outputs(6009) <= not b or a;
    layer1_outputs(6010) <= a xor b;
    layer1_outputs(6011) <= a or b;
    layer1_outputs(6012) <= a and b;
    layer1_outputs(6013) <= a and not b;
    layer1_outputs(6014) <= b and not a;
    layer1_outputs(6015) <= not b;
    layer1_outputs(6016) <= a;
    layer1_outputs(6017) <= a or b;
    layer1_outputs(6018) <= not (a xor b);
    layer1_outputs(6019) <= a xor b;
    layer1_outputs(6020) <= a;
    layer1_outputs(6021) <= not (a or b);
    layer1_outputs(6022) <= b;
    layer1_outputs(6023) <= not a;
    layer1_outputs(6024) <= b;
    layer1_outputs(6025) <= b;
    layer1_outputs(6026) <= not (a or b);
    layer1_outputs(6027) <= not b;
    layer1_outputs(6028) <= not b or a;
    layer1_outputs(6029) <= a;
    layer1_outputs(6030) <= a;
    layer1_outputs(6031) <= b;
    layer1_outputs(6032) <= not (a xor b);
    layer1_outputs(6033) <= not a or b;
    layer1_outputs(6034) <= not a;
    layer1_outputs(6035) <= a or b;
    layer1_outputs(6036) <= not (a xor b);
    layer1_outputs(6037) <= a and b;
    layer1_outputs(6038) <= not (a and b);
    layer1_outputs(6039) <= b and not a;
    layer1_outputs(6040) <= not b or a;
    layer1_outputs(6041) <= not a;
    layer1_outputs(6042) <= not b;
    layer1_outputs(6043) <= not b;
    layer1_outputs(6044) <= a and b;
    layer1_outputs(6045) <= a or b;
    layer1_outputs(6046) <= a and not b;
    layer1_outputs(6047) <= not a or b;
    layer1_outputs(6048) <= a xor b;
    layer1_outputs(6049) <= '1';
    layer1_outputs(6050) <= b;
    layer1_outputs(6051) <= b;
    layer1_outputs(6052) <= a and b;
    layer1_outputs(6053) <= '1';
    layer1_outputs(6054) <= not b;
    layer1_outputs(6055) <= not a;
    layer1_outputs(6056) <= a and b;
    layer1_outputs(6057) <= not b;
    layer1_outputs(6058) <= b;
    layer1_outputs(6059) <= a xor b;
    layer1_outputs(6060) <= '0';
    layer1_outputs(6061) <= a xor b;
    layer1_outputs(6062) <= not b;
    layer1_outputs(6063) <= a;
    layer1_outputs(6064) <= a xor b;
    layer1_outputs(6065) <= not a or b;
    layer1_outputs(6066) <= a or b;
    layer1_outputs(6067) <= not (a xor b);
    layer1_outputs(6068) <= a or b;
    layer1_outputs(6069) <= not b;
    layer1_outputs(6070) <= '1';
    layer1_outputs(6071) <= not a or b;
    layer1_outputs(6072) <= a and b;
    layer1_outputs(6073) <= not b;
    layer1_outputs(6074) <= not (a xor b);
    layer1_outputs(6075) <= not b or a;
    layer1_outputs(6076) <= a and not b;
    layer1_outputs(6077) <= not a;
    layer1_outputs(6078) <= '0';
    layer1_outputs(6079) <= b;
    layer1_outputs(6080) <= not a;
    layer1_outputs(6081) <= a xor b;
    layer1_outputs(6082) <= a;
    layer1_outputs(6083) <= not b;
    layer1_outputs(6084) <= not (a and b);
    layer1_outputs(6085) <= not (a xor b);
    layer1_outputs(6086) <= not (a or b);
    layer1_outputs(6087) <= b and not a;
    layer1_outputs(6088) <= not b;
    layer1_outputs(6089) <= not a;
    layer1_outputs(6090) <= a xor b;
    layer1_outputs(6091) <= not b or a;
    layer1_outputs(6092) <= not (a and b);
    layer1_outputs(6093) <= a or b;
    layer1_outputs(6094) <= a xor b;
    layer1_outputs(6095) <= b;
    layer1_outputs(6096) <= not (a and b);
    layer1_outputs(6097) <= not a;
    layer1_outputs(6098) <= b and not a;
    layer1_outputs(6099) <= a;
    layer1_outputs(6100) <= b;
    layer1_outputs(6101) <= b;
    layer1_outputs(6102) <= not b;
    layer1_outputs(6103) <= a xor b;
    layer1_outputs(6104) <= not b;
    layer1_outputs(6105) <= not a;
    layer1_outputs(6106) <= b;
    layer1_outputs(6107) <= not (a or b);
    layer1_outputs(6108) <= b;
    layer1_outputs(6109) <= a and not b;
    layer1_outputs(6110) <= a or b;
    layer1_outputs(6111) <= b;
    layer1_outputs(6112) <= a xor b;
    layer1_outputs(6113) <= not b;
    layer1_outputs(6114) <= not (a xor b);
    layer1_outputs(6115) <= '0';
    layer1_outputs(6116) <= not (a and b);
    layer1_outputs(6117) <= a and b;
    layer1_outputs(6118) <= not a or b;
    layer1_outputs(6119) <= not (a xor b);
    layer1_outputs(6120) <= a or b;
    layer1_outputs(6121) <= b;
    layer1_outputs(6122) <= b;
    layer1_outputs(6123) <= not a;
    layer1_outputs(6124) <= not b or a;
    layer1_outputs(6125) <= not (a and b);
    layer1_outputs(6126) <= b;
    layer1_outputs(6127) <= a and not b;
    layer1_outputs(6128) <= not b;
    layer1_outputs(6129) <= a or b;
    layer1_outputs(6130) <= a;
    layer1_outputs(6131) <= not a;
    layer1_outputs(6132) <= b;
    layer1_outputs(6133) <= not b;
    layer1_outputs(6134) <= not (a xor b);
    layer1_outputs(6135) <= not (a or b);
    layer1_outputs(6136) <= a xor b;
    layer1_outputs(6137) <= not b or a;
    layer1_outputs(6138) <= a;
    layer1_outputs(6139) <= not a or b;
    layer1_outputs(6140) <= a;
    layer1_outputs(6141) <= not a;
    layer1_outputs(6142) <= not (a or b);
    layer1_outputs(6143) <= not a or b;
    layer1_outputs(6144) <= a and b;
    layer1_outputs(6145) <= not (a or b);
    layer1_outputs(6146) <= not (a or b);
    layer1_outputs(6147) <= not (a and b);
    layer1_outputs(6148) <= a and not b;
    layer1_outputs(6149) <= not a or b;
    layer1_outputs(6150) <= a xor b;
    layer1_outputs(6151) <= a;
    layer1_outputs(6152) <= not a or b;
    layer1_outputs(6153) <= a xor b;
    layer1_outputs(6154) <= not (a xor b);
    layer1_outputs(6155) <= not (a xor b);
    layer1_outputs(6156) <= a;
    layer1_outputs(6157) <= not (a or b);
    layer1_outputs(6158) <= a or b;
    layer1_outputs(6159) <= not a;
    layer1_outputs(6160) <= b;
    layer1_outputs(6161) <= b and not a;
    layer1_outputs(6162) <= not a;
    layer1_outputs(6163) <= a xor b;
    layer1_outputs(6164) <= a xor b;
    layer1_outputs(6165) <= not a;
    layer1_outputs(6166) <= a and not b;
    layer1_outputs(6167) <= not a or b;
    layer1_outputs(6168) <= not b or a;
    layer1_outputs(6169) <= not b;
    layer1_outputs(6170) <= b and not a;
    layer1_outputs(6171) <= not a or b;
    layer1_outputs(6172) <= not (a xor b);
    layer1_outputs(6173) <= a;
    layer1_outputs(6174) <= not (a xor b);
    layer1_outputs(6175) <= a xor b;
    layer1_outputs(6176) <= a xor b;
    layer1_outputs(6177) <= a or b;
    layer1_outputs(6178) <= not (a and b);
    layer1_outputs(6179) <= not (a xor b);
    layer1_outputs(6180) <= not b;
    layer1_outputs(6181) <= a;
    layer1_outputs(6182) <= b and not a;
    layer1_outputs(6183) <= not a or b;
    layer1_outputs(6184) <= a;
    layer1_outputs(6185) <= a or b;
    layer1_outputs(6186) <= not a;
    layer1_outputs(6187) <= not a or b;
    layer1_outputs(6188) <= a xor b;
    layer1_outputs(6189) <= a xor b;
    layer1_outputs(6190) <= not a or b;
    layer1_outputs(6191) <= not b;
    layer1_outputs(6192) <= not b or a;
    layer1_outputs(6193) <= a xor b;
    layer1_outputs(6194) <= a;
    layer1_outputs(6195) <= a or b;
    layer1_outputs(6196) <= a;
    layer1_outputs(6197) <= a and b;
    layer1_outputs(6198) <= not (a and b);
    layer1_outputs(6199) <= not (a xor b);
    layer1_outputs(6200) <= not b or a;
    layer1_outputs(6201) <= a and b;
    layer1_outputs(6202) <= a xor b;
    layer1_outputs(6203) <= a and not b;
    layer1_outputs(6204) <= not b;
    layer1_outputs(6205) <= '1';
    layer1_outputs(6206) <= a and b;
    layer1_outputs(6207) <= not a or b;
    layer1_outputs(6208) <= b and not a;
    layer1_outputs(6209) <= a or b;
    layer1_outputs(6210) <= a or b;
    layer1_outputs(6211) <= b;
    layer1_outputs(6212) <= not (a xor b);
    layer1_outputs(6213) <= not a or b;
    layer1_outputs(6214) <= not (a xor b);
    layer1_outputs(6215) <= a and b;
    layer1_outputs(6216) <= not a or b;
    layer1_outputs(6217) <= b;
    layer1_outputs(6218) <= a or b;
    layer1_outputs(6219) <= not b;
    layer1_outputs(6220) <= not a or b;
    layer1_outputs(6221) <= not a or b;
    layer1_outputs(6222) <= a and b;
    layer1_outputs(6223) <= a and not b;
    layer1_outputs(6224) <= b;
    layer1_outputs(6225) <= not b or a;
    layer1_outputs(6226) <= a and b;
    layer1_outputs(6227) <= not a;
    layer1_outputs(6228) <= not (a and b);
    layer1_outputs(6229) <= a or b;
    layer1_outputs(6230) <= a;
    layer1_outputs(6231) <= not a;
    layer1_outputs(6232) <= not a or b;
    layer1_outputs(6233) <= not b or a;
    layer1_outputs(6234) <= not (a xor b);
    layer1_outputs(6235) <= '0';
    layer1_outputs(6236) <= not b;
    layer1_outputs(6237) <= not a;
    layer1_outputs(6238) <= b;
    layer1_outputs(6239) <= a and b;
    layer1_outputs(6240) <= a or b;
    layer1_outputs(6241) <= not (a xor b);
    layer1_outputs(6242) <= a or b;
    layer1_outputs(6243) <= a;
    layer1_outputs(6244) <= not (a or b);
    layer1_outputs(6245) <= not a;
    layer1_outputs(6246) <= not (a xor b);
    layer1_outputs(6247) <= not (a and b);
    layer1_outputs(6248) <= not b;
    layer1_outputs(6249) <= not a;
    layer1_outputs(6250) <= not a or b;
    layer1_outputs(6251) <= not b;
    layer1_outputs(6252) <= not b;
    layer1_outputs(6253) <= a;
    layer1_outputs(6254) <= a and not b;
    layer1_outputs(6255) <= b and not a;
    layer1_outputs(6256) <= b;
    layer1_outputs(6257) <= not b;
    layer1_outputs(6258) <= not a;
    layer1_outputs(6259) <= b and not a;
    layer1_outputs(6260) <= not b or a;
    layer1_outputs(6261) <= not (a xor b);
    layer1_outputs(6262) <= not (a or b);
    layer1_outputs(6263) <= b;
    layer1_outputs(6264) <= not b or a;
    layer1_outputs(6265) <= b;
    layer1_outputs(6266) <= b and not a;
    layer1_outputs(6267) <= not a;
    layer1_outputs(6268) <= a xor b;
    layer1_outputs(6269) <= a and not b;
    layer1_outputs(6270) <= not b or a;
    layer1_outputs(6271) <= a;
    layer1_outputs(6272) <= b;
    layer1_outputs(6273) <= a;
    layer1_outputs(6274) <= b and not a;
    layer1_outputs(6275) <= not (a or b);
    layer1_outputs(6276) <= not a;
    layer1_outputs(6277) <= not (a and b);
    layer1_outputs(6278) <= a and b;
    layer1_outputs(6279) <= not b or a;
    layer1_outputs(6280) <= not a;
    layer1_outputs(6281) <= a xor b;
    layer1_outputs(6282) <= not (a and b);
    layer1_outputs(6283) <= a;
    layer1_outputs(6284) <= not b or a;
    layer1_outputs(6285) <= a and b;
    layer1_outputs(6286) <= a or b;
    layer1_outputs(6287) <= not (a xor b);
    layer1_outputs(6288) <= a and b;
    layer1_outputs(6289) <= not (a and b);
    layer1_outputs(6290) <= not b or a;
    layer1_outputs(6291) <= not a;
    layer1_outputs(6292) <= b and not a;
    layer1_outputs(6293) <= not a or b;
    layer1_outputs(6294) <= a;
    layer1_outputs(6295) <= a or b;
    layer1_outputs(6296) <= a;
    layer1_outputs(6297) <= a;
    layer1_outputs(6298) <= a and b;
    layer1_outputs(6299) <= not b or a;
    layer1_outputs(6300) <= a or b;
    layer1_outputs(6301) <= a or b;
    layer1_outputs(6302) <= not (a or b);
    layer1_outputs(6303) <= not (a xor b);
    layer1_outputs(6304) <= a or b;
    layer1_outputs(6305) <= not b or a;
    layer1_outputs(6306) <= not (a and b);
    layer1_outputs(6307) <= a and not b;
    layer1_outputs(6308) <= not (a or b);
    layer1_outputs(6309) <= not (a or b);
    layer1_outputs(6310) <= a xor b;
    layer1_outputs(6311) <= not b;
    layer1_outputs(6312) <= a and not b;
    layer1_outputs(6313) <= a xor b;
    layer1_outputs(6314) <= a and not b;
    layer1_outputs(6315) <= a or b;
    layer1_outputs(6316) <= a or b;
    layer1_outputs(6317) <= '1';
    layer1_outputs(6318) <= a and b;
    layer1_outputs(6319) <= b and not a;
    layer1_outputs(6320) <= not (a or b);
    layer1_outputs(6321) <= not (a or b);
    layer1_outputs(6322) <= a xor b;
    layer1_outputs(6323) <= b;
    layer1_outputs(6324) <= a and b;
    layer1_outputs(6325) <= a and not b;
    layer1_outputs(6326) <= a;
    layer1_outputs(6327) <= not b or a;
    layer1_outputs(6328) <= not a or b;
    layer1_outputs(6329) <= a or b;
    layer1_outputs(6330) <= a;
    layer1_outputs(6331) <= not (a xor b);
    layer1_outputs(6332) <= not a;
    layer1_outputs(6333) <= '0';
    layer1_outputs(6334) <= a or b;
    layer1_outputs(6335) <= a;
    layer1_outputs(6336) <= not b or a;
    layer1_outputs(6337) <= not a;
    layer1_outputs(6338) <= a;
    layer1_outputs(6339) <= b;
    layer1_outputs(6340) <= a and b;
    layer1_outputs(6341) <= b;
    layer1_outputs(6342) <= b and not a;
    layer1_outputs(6343) <= not a;
    layer1_outputs(6344) <= not (a and b);
    layer1_outputs(6345) <= not a;
    layer1_outputs(6346) <= a xor b;
    layer1_outputs(6347) <= not (a or b);
    layer1_outputs(6348) <= not a;
    layer1_outputs(6349) <= not (a or b);
    layer1_outputs(6350) <= not a or b;
    layer1_outputs(6351) <= a or b;
    layer1_outputs(6352) <= not a;
    layer1_outputs(6353) <= a;
    layer1_outputs(6354) <= not b;
    layer1_outputs(6355) <= not (a or b);
    layer1_outputs(6356) <= b and not a;
    layer1_outputs(6357) <= b and not a;
    layer1_outputs(6358) <= not (a xor b);
    layer1_outputs(6359) <= not b or a;
    layer1_outputs(6360) <= a;
    layer1_outputs(6361) <= not b;
    layer1_outputs(6362) <= not a or b;
    layer1_outputs(6363) <= not a or b;
    layer1_outputs(6364) <= not a or b;
    layer1_outputs(6365) <= a and not b;
    layer1_outputs(6366) <= not (a xor b);
    layer1_outputs(6367) <= a;
    layer1_outputs(6368) <= not a;
    layer1_outputs(6369) <= b;
    layer1_outputs(6370) <= b and not a;
    layer1_outputs(6371) <= a and not b;
    layer1_outputs(6372) <= a xor b;
    layer1_outputs(6373) <= not (a or b);
    layer1_outputs(6374) <= b;
    layer1_outputs(6375) <= not a or b;
    layer1_outputs(6376) <= b;
    layer1_outputs(6377) <= a and b;
    layer1_outputs(6378) <= b and not a;
    layer1_outputs(6379) <= a;
    layer1_outputs(6380) <= not a or b;
    layer1_outputs(6381) <= b;
    layer1_outputs(6382) <= not b or a;
    layer1_outputs(6383) <= b and not a;
    layer1_outputs(6384) <= a xor b;
    layer1_outputs(6385) <= not b or a;
    layer1_outputs(6386) <= a;
    layer1_outputs(6387) <= not (a xor b);
    layer1_outputs(6388) <= a xor b;
    layer1_outputs(6389) <= a;
    layer1_outputs(6390) <= a;
    layer1_outputs(6391) <= not (a xor b);
    layer1_outputs(6392) <= not a or b;
    layer1_outputs(6393) <= a or b;
    layer1_outputs(6394) <= b and not a;
    layer1_outputs(6395) <= not b;
    layer1_outputs(6396) <= b;
    layer1_outputs(6397) <= b;
    layer1_outputs(6398) <= not a;
    layer1_outputs(6399) <= a and not b;
    layer1_outputs(6400) <= a;
    layer1_outputs(6401) <= not (a and b);
    layer1_outputs(6402) <= not (a or b);
    layer1_outputs(6403) <= a and not b;
    layer1_outputs(6404) <= not a or b;
    layer1_outputs(6405) <= not b or a;
    layer1_outputs(6406) <= not (a xor b);
    layer1_outputs(6407) <= a;
    layer1_outputs(6408) <= not (a xor b);
    layer1_outputs(6409) <= not a;
    layer1_outputs(6410) <= not (a or b);
    layer1_outputs(6411) <= not b;
    layer1_outputs(6412) <= not b or a;
    layer1_outputs(6413) <= b;
    layer1_outputs(6414) <= a;
    layer1_outputs(6415) <= b;
    layer1_outputs(6416) <= b and not a;
    layer1_outputs(6417) <= a and not b;
    layer1_outputs(6418) <= not b or a;
    layer1_outputs(6419) <= not b;
    layer1_outputs(6420) <= not a or b;
    layer1_outputs(6421) <= a or b;
    layer1_outputs(6422) <= a and not b;
    layer1_outputs(6423) <= a;
    layer1_outputs(6424) <= a;
    layer1_outputs(6425) <= not (a or b);
    layer1_outputs(6426) <= not (a xor b);
    layer1_outputs(6427) <= not a;
    layer1_outputs(6428) <= b and not a;
    layer1_outputs(6429) <= not (a and b);
    layer1_outputs(6430) <= not (a xor b);
    layer1_outputs(6431) <= a and not b;
    layer1_outputs(6432) <= '1';
    layer1_outputs(6433) <= not (a or b);
    layer1_outputs(6434) <= a xor b;
    layer1_outputs(6435) <= not (a and b);
    layer1_outputs(6436) <= not (a or b);
    layer1_outputs(6437) <= not a;
    layer1_outputs(6438) <= not (a and b);
    layer1_outputs(6439) <= not b;
    layer1_outputs(6440) <= a and b;
    layer1_outputs(6441) <= a and not b;
    layer1_outputs(6442) <= b and not a;
    layer1_outputs(6443) <= not a;
    layer1_outputs(6444) <= not b or a;
    layer1_outputs(6445) <= not b or a;
    layer1_outputs(6446) <= b and not a;
    layer1_outputs(6447) <= not a;
    layer1_outputs(6448) <= not b or a;
    layer1_outputs(6449) <= not a or b;
    layer1_outputs(6450) <= not b;
    layer1_outputs(6451) <= not a;
    layer1_outputs(6452) <= not a;
    layer1_outputs(6453) <= a;
    layer1_outputs(6454) <= not (a xor b);
    layer1_outputs(6455) <= b and not a;
    layer1_outputs(6456) <= b;
    layer1_outputs(6457) <= not (a xor b);
    layer1_outputs(6458) <= b;
    layer1_outputs(6459) <= not b;
    layer1_outputs(6460) <= not (a and b);
    layer1_outputs(6461) <= not a;
    layer1_outputs(6462) <= b;
    layer1_outputs(6463) <= not (a xor b);
    layer1_outputs(6464) <= a and b;
    layer1_outputs(6465) <= a or b;
    layer1_outputs(6466) <= b and not a;
    layer1_outputs(6467) <= b;
    layer1_outputs(6468) <= a;
    layer1_outputs(6469) <= '0';
    layer1_outputs(6470) <= a and not b;
    layer1_outputs(6471) <= not (a or b);
    layer1_outputs(6472) <= a or b;
    layer1_outputs(6473) <= not a;
    layer1_outputs(6474) <= a;
    layer1_outputs(6475) <= not (a and b);
    layer1_outputs(6476) <= not b;
    layer1_outputs(6477) <= not b;
    layer1_outputs(6478) <= not b or a;
    layer1_outputs(6479) <= a xor b;
    layer1_outputs(6480) <= a;
    layer1_outputs(6481) <= a;
    layer1_outputs(6482) <= a;
    layer1_outputs(6483) <= a and b;
    layer1_outputs(6484) <= not (a or b);
    layer1_outputs(6485) <= not a or b;
    layer1_outputs(6486) <= b;
    layer1_outputs(6487) <= not b;
    layer1_outputs(6488) <= not b;
    layer1_outputs(6489) <= not b;
    layer1_outputs(6490) <= b and not a;
    layer1_outputs(6491) <= a;
    layer1_outputs(6492) <= a and b;
    layer1_outputs(6493) <= b;
    layer1_outputs(6494) <= '0';
    layer1_outputs(6495) <= not b;
    layer1_outputs(6496) <= b;
    layer1_outputs(6497) <= b and not a;
    layer1_outputs(6498) <= not (a and b);
    layer1_outputs(6499) <= not (a xor b);
    layer1_outputs(6500) <= not (a and b);
    layer1_outputs(6501) <= a;
    layer1_outputs(6502) <= not a or b;
    layer1_outputs(6503) <= a;
    layer1_outputs(6504) <= b;
    layer1_outputs(6505) <= a and not b;
    layer1_outputs(6506) <= b and not a;
    layer1_outputs(6507) <= b and not a;
    layer1_outputs(6508) <= not (a or b);
    layer1_outputs(6509) <= not (a or b);
    layer1_outputs(6510) <= not b;
    layer1_outputs(6511) <= a or b;
    layer1_outputs(6512) <= a or b;
    layer1_outputs(6513) <= not b;
    layer1_outputs(6514) <= a;
    layer1_outputs(6515) <= not (a or b);
    layer1_outputs(6516) <= a and not b;
    layer1_outputs(6517) <= a and b;
    layer1_outputs(6518) <= a and not b;
    layer1_outputs(6519) <= a;
    layer1_outputs(6520) <= a;
    layer1_outputs(6521) <= a xor b;
    layer1_outputs(6522) <= not a;
    layer1_outputs(6523) <= a;
    layer1_outputs(6524) <= a xor b;
    layer1_outputs(6525) <= a xor b;
    layer1_outputs(6526) <= not b;
    layer1_outputs(6527) <= b;
    layer1_outputs(6528) <= a xor b;
    layer1_outputs(6529) <= a;
    layer1_outputs(6530) <= a;
    layer1_outputs(6531) <= b;
    layer1_outputs(6532) <= b and not a;
    layer1_outputs(6533) <= not a or b;
    layer1_outputs(6534) <= not a or b;
    layer1_outputs(6535) <= a;
    layer1_outputs(6536) <= not b;
    layer1_outputs(6537) <= not b;
    layer1_outputs(6538) <= not (a and b);
    layer1_outputs(6539) <= '0';
    layer1_outputs(6540) <= not (a or b);
    layer1_outputs(6541) <= not b or a;
    layer1_outputs(6542) <= not b;
    layer1_outputs(6543) <= not a or b;
    layer1_outputs(6544) <= not b or a;
    layer1_outputs(6545) <= a or b;
    layer1_outputs(6546) <= a;
    layer1_outputs(6547) <= a;
    layer1_outputs(6548) <= a or b;
    layer1_outputs(6549) <= not a or b;
    layer1_outputs(6550) <= b and not a;
    layer1_outputs(6551) <= not b;
    layer1_outputs(6552) <= not (a and b);
    layer1_outputs(6553) <= '1';
    layer1_outputs(6554) <= a and not b;
    layer1_outputs(6555) <= not (a and b);
    layer1_outputs(6556) <= not b or a;
    layer1_outputs(6557) <= b;
    layer1_outputs(6558) <= a xor b;
    layer1_outputs(6559) <= not (a and b);
    layer1_outputs(6560) <= a and not b;
    layer1_outputs(6561) <= a or b;
    layer1_outputs(6562) <= a;
    layer1_outputs(6563) <= a;
    layer1_outputs(6564) <= b and not a;
    layer1_outputs(6565) <= not a or b;
    layer1_outputs(6566) <= a;
    layer1_outputs(6567) <= a xor b;
    layer1_outputs(6568) <= not (a and b);
    layer1_outputs(6569) <= not a;
    layer1_outputs(6570) <= a and b;
    layer1_outputs(6571) <= a;
    layer1_outputs(6572) <= a and b;
    layer1_outputs(6573) <= not (a or b);
    layer1_outputs(6574) <= not a;
    layer1_outputs(6575) <= a and b;
    layer1_outputs(6576) <= b;
    layer1_outputs(6577) <= b;
    layer1_outputs(6578) <= not b;
    layer1_outputs(6579) <= a and b;
    layer1_outputs(6580) <= a and not b;
    layer1_outputs(6581) <= a;
    layer1_outputs(6582) <= a and not b;
    layer1_outputs(6583) <= a;
    layer1_outputs(6584) <= a and not b;
    layer1_outputs(6585) <= not a;
    layer1_outputs(6586) <= not a;
    layer1_outputs(6587) <= not a;
    layer1_outputs(6588) <= not (a or b);
    layer1_outputs(6589) <= not (a or b);
    layer1_outputs(6590) <= not b or a;
    layer1_outputs(6591) <= a;
    layer1_outputs(6592) <= a xor b;
    layer1_outputs(6593) <= not (a xor b);
    layer1_outputs(6594) <= a and not b;
    layer1_outputs(6595) <= not a or b;
    layer1_outputs(6596) <= '0';
    layer1_outputs(6597) <= not b or a;
    layer1_outputs(6598) <= b;
    layer1_outputs(6599) <= a and b;
    layer1_outputs(6600) <= a;
    layer1_outputs(6601) <= not a or b;
    layer1_outputs(6602) <= b and not a;
    layer1_outputs(6603) <= a;
    layer1_outputs(6604) <= a;
    layer1_outputs(6605) <= not (a xor b);
    layer1_outputs(6606) <= not (a and b);
    layer1_outputs(6607) <= not a;
    layer1_outputs(6608) <= a and b;
    layer1_outputs(6609) <= b;
    layer1_outputs(6610) <= b and not a;
    layer1_outputs(6611) <= a xor b;
    layer1_outputs(6612) <= b;
    layer1_outputs(6613) <= b and not a;
    layer1_outputs(6614) <= a;
    layer1_outputs(6615) <= b and not a;
    layer1_outputs(6616) <= b and not a;
    layer1_outputs(6617) <= not (a xor b);
    layer1_outputs(6618) <= a;
    layer1_outputs(6619) <= not (a xor b);
    layer1_outputs(6620) <= not (a xor b);
    layer1_outputs(6621) <= not a or b;
    layer1_outputs(6622) <= a or b;
    layer1_outputs(6623) <= a and not b;
    layer1_outputs(6624) <= b;
    layer1_outputs(6625) <= not (a xor b);
    layer1_outputs(6626) <= a or b;
    layer1_outputs(6627) <= not a;
    layer1_outputs(6628) <= not a or b;
    layer1_outputs(6629) <= not a;
    layer1_outputs(6630) <= not b;
    layer1_outputs(6631) <= a and not b;
    layer1_outputs(6632) <= a;
    layer1_outputs(6633) <= not (a xor b);
    layer1_outputs(6634) <= b and not a;
    layer1_outputs(6635) <= not (a and b);
    layer1_outputs(6636) <= not b;
    layer1_outputs(6637) <= a and not b;
    layer1_outputs(6638) <= not (a and b);
    layer1_outputs(6639) <= a and b;
    layer1_outputs(6640) <= a xor b;
    layer1_outputs(6641) <= not a or b;
    layer1_outputs(6642) <= b;
    layer1_outputs(6643) <= b;
    layer1_outputs(6644) <= a xor b;
    layer1_outputs(6645) <= b and not a;
    layer1_outputs(6646) <= b;
    layer1_outputs(6647) <= not (a or b);
    layer1_outputs(6648) <= a or b;
    layer1_outputs(6649) <= a or b;
    layer1_outputs(6650) <= a xor b;
    layer1_outputs(6651) <= a xor b;
    layer1_outputs(6652) <= not b or a;
    layer1_outputs(6653) <= not a;
    layer1_outputs(6654) <= a and b;
    layer1_outputs(6655) <= not (a xor b);
    layer1_outputs(6656) <= a;
    layer1_outputs(6657) <= a;
    layer1_outputs(6658) <= a xor b;
    layer1_outputs(6659) <= '0';
    layer1_outputs(6660) <= not a;
    layer1_outputs(6661) <= not a;
    layer1_outputs(6662) <= a or b;
    layer1_outputs(6663) <= not a;
    layer1_outputs(6664) <= not b;
    layer1_outputs(6665) <= b;
    layer1_outputs(6666) <= not (a or b);
    layer1_outputs(6667) <= not (a or b);
    layer1_outputs(6668) <= not (a and b);
    layer1_outputs(6669) <= b;
    layer1_outputs(6670) <= a and not b;
    layer1_outputs(6671) <= a and b;
    layer1_outputs(6672) <= not a;
    layer1_outputs(6673) <= a;
    layer1_outputs(6674) <= not b or a;
    layer1_outputs(6675) <= not b;
    layer1_outputs(6676) <= a xor b;
    layer1_outputs(6677) <= not (a xor b);
    layer1_outputs(6678) <= a and not b;
    layer1_outputs(6679) <= b;
    layer1_outputs(6680) <= not (a and b);
    layer1_outputs(6681) <= not b;
    layer1_outputs(6682) <= not a or b;
    layer1_outputs(6683) <= b;
    layer1_outputs(6684) <= b;
    layer1_outputs(6685) <= not (a xor b);
    layer1_outputs(6686) <= a or b;
    layer1_outputs(6687) <= not a;
    layer1_outputs(6688) <= b;
    layer1_outputs(6689) <= a;
    layer1_outputs(6690) <= a;
    layer1_outputs(6691) <= not (a and b);
    layer1_outputs(6692) <= b;
    layer1_outputs(6693) <= not (a xor b);
    layer1_outputs(6694) <= not (a xor b);
    layer1_outputs(6695) <= a;
    layer1_outputs(6696) <= not (a or b);
    layer1_outputs(6697) <= b and not a;
    layer1_outputs(6698) <= not a;
    layer1_outputs(6699) <= b and not a;
    layer1_outputs(6700) <= a;
    layer1_outputs(6701) <= a;
    layer1_outputs(6702) <= not a;
    layer1_outputs(6703) <= not (a xor b);
    layer1_outputs(6704) <= not (a xor b);
    layer1_outputs(6705) <= a or b;
    layer1_outputs(6706) <= b and not a;
    layer1_outputs(6707) <= not (a xor b);
    layer1_outputs(6708) <= not b;
    layer1_outputs(6709) <= not (a xor b);
    layer1_outputs(6710) <= a xor b;
    layer1_outputs(6711) <= b;
    layer1_outputs(6712) <= not b;
    layer1_outputs(6713) <= not (a xor b);
    layer1_outputs(6714) <= not (a or b);
    layer1_outputs(6715) <= a xor b;
    layer1_outputs(6716) <= a and not b;
    layer1_outputs(6717) <= not b;
    layer1_outputs(6718) <= b and not a;
    layer1_outputs(6719) <= a;
    layer1_outputs(6720) <= b and not a;
    layer1_outputs(6721) <= a;
    layer1_outputs(6722) <= b and not a;
    layer1_outputs(6723) <= a or b;
    layer1_outputs(6724) <= not a or b;
    layer1_outputs(6725) <= '1';
    layer1_outputs(6726) <= not (a or b);
    layer1_outputs(6727) <= a xor b;
    layer1_outputs(6728) <= a xor b;
    layer1_outputs(6729) <= not (a and b);
    layer1_outputs(6730) <= a and b;
    layer1_outputs(6731) <= not a or b;
    layer1_outputs(6732) <= a;
    layer1_outputs(6733) <= a or b;
    layer1_outputs(6734) <= a xor b;
    layer1_outputs(6735) <= not (a and b);
    layer1_outputs(6736) <= a xor b;
    layer1_outputs(6737) <= '1';
    layer1_outputs(6738) <= not (a or b);
    layer1_outputs(6739) <= b and not a;
    layer1_outputs(6740) <= not a;
    layer1_outputs(6741) <= '0';
    layer1_outputs(6742) <= a or b;
    layer1_outputs(6743) <= not a;
    layer1_outputs(6744) <= a;
    layer1_outputs(6745) <= a;
    layer1_outputs(6746) <= not b;
    layer1_outputs(6747) <= a;
    layer1_outputs(6748) <= a;
    layer1_outputs(6749) <= not b;
    layer1_outputs(6750) <= b;
    layer1_outputs(6751) <= a;
    layer1_outputs(6752) <= not a;
    layer1_outputs(6753) <= not (a and b);
    layer1_outputs(6754) <= a and b;
    layer1_outputs(6755) <= not b;
    layer1_outputs(6756) <= not a or b;
    layer1_outputs(6757) <= a and not b;
    layer1_outputs(6758) <= b and not a;
    layer1_outputs(6759) <= not b or a;
    layer1_outputs(6760) <= not a;
    layer1_outputs(6761) <= a or b;
    layer1_outputs(6762) <= '1';
    layer1_outputs(6763) <= not b;
    layer1_outputs(6764) <= a and not b;
    layer1_outputs(6765) <= not (a xor b);
    layer1_outputs(6766) <= not (a xor b);
    layer1_outputs(6767) <= not b or a;
    layer1_outputs(6768) <= a;
    layer1_outputs(6769) <= a xor b;
    layer1_outputs(6770) <= not (a or b);
    layer1_outputs(6771) <= a xor b;
    layer1_outputs(6772) <= b and not a;
    layer1_outputs(6773) <= b;
    layer1_outputs(6774) <= not b;
    layer1_outputs(6775) <= b and not a;
    layer1_outputs(6776) <= a and not b;
    layer1_outputs(6777) <= not b;
    layer1_outputs(6778) <= not b;
    layer1_outputs(6779) <= not (a xor b);
    layer1_outputs(6780) <= not b;
    layer1_outputs(6781) <= a;
    layer1_outputs(6782) <= not b;
    layer1_outputs(6783) <= a or b;
    layer1_outputs(6784) <= not (a xor b);
    layer1_outputs(6785) <= not b or a;
    layer1_outputs(6786) <= not (a and b);
    layer1_outputs(6787) <= not a or b;
    layer1_outputs(6788) <= a or b;
    layer1_outputs(6789) <= not (a and b);
    layer1_outputs(6790) <= b and not a;
    layer1_outputs(6791) <= a and b;
    layer1_outputs(6792) <= a and not b;
    layer1_outputs(6793) <= not (a and b);
    layer1_outputs(6794) <= a and b;
    layer1_outputs(6795) <= b and not a;
    layer1_outputs(6796) <= not (a xor b);
    layer1_outputs(6797) <= a or b;
    layer1_outputs(6798) <= a;
    layer1_outputs(6799) <= not b or a;
    layer1_outputs(6800) <= a or b;
    layer1_outputs(6801) <= not a or b;
    layer1_outputs(6802) <= a xor b;
    layer1_outputs(6803) <= '0';
    layer1_outputs(6804) <= not (a or b);
    layer1_outputs(6805) <= not a;
    layer1_outputs(6806) <= a and not b;
    layer1_outputs(6807) <= a and b;
    layer1_outputs(6808) <= a xor b;
    layer1_outputs(6809) <= not a or b;
    layer1_outputs(6810) <= not (a and b);
    layer1_outputs(6811) <= not a or b;
    layer1_outputs(6812) <= b;
    layer1_outputs(6813) <= not (a xor b);
    layer1_outputs(6814) <= a and b;
    layer1_outputs(6815) <= a and not b;
    layer1_outputs(6816) <= a and b;
    layer1_outputs(6817) <= a;
    layer1_outputs(6818) <= a xor b;
    layer1_outputs(6819) <= b and not a;
    layer1_outputs(6820) <= a or b;
    layer1_outputs(6821) <= b and not a;
    layer1_outputs(6822) <= not a or b;
    layer1_outputs(6823) <= not a or b;
    layer1_outputs(6824) <= not a or b;
    layer1_outputs(6825) <= not a or b;
    layer1_outputs(6826) <= not (a xor b);
    layer1_outputs(6827) <= a;
    layer1_outputs(6828) <= not a;
    layer1_outputs(6829) <= b and not a;
    layer1_outputs(6830) <= not b or a;
    layer1_outputs(6831) <= a xor b;
    layer1_outputs(6832) <= b;
    layer1_outputs(6833) <= not b;
    layer1_outputs(6834) <= not b or a;
    layer1_outputs(6835) <= a and b;
    layer1_outputs(6836) <= not (a or b);
    layer1_outputs(6837) <= b;
    layer1_outputs(6838) <= a or b;
    layer1_outputs(6839) <= a;
    layer1_outputs(6840) <= b;
    layer1_outputs(6841) <= not (a xor b);
    layer1_outputs(6842) <= b;
    layer1_outputs(6843) <= b and not a;
    layer1_outputs(6844) <= not a;
    layer1_outputs(6845) <= not (a or b);
    layer1_outputs(6846) <= a and b;
    layer1_outputs(6847) <= not (a and b);
    layer1_outputs(6848) <= a or b;
    layer1_outputs(6849) <= b;
    layer1_outputs(6850) <= b;
    layer1_outputs(6851) <= not b;
    layer1_outputs(6852) <= a;
    layer1_outputs(6853) <= a and b;
    layer1_outputs(6854) <= a and not b;
    layer1_outputs(6855) <= b;
    layer1_outputs(6856) <= a;
    layer1_outputs(6857) <= not b;
    layer1_outputs(6858) <= not (a or b);
    layer1_outputs(6859) <= not b;
    layer1_outputs(6860) <= not b or a;
    layer1_outputs(6861) <= '1';
    layer1_outputs(6862) <= not b;
    layer1_outputs(6863) <= a;
    layer1_outputs(6864) <= not (a or b);
    layer1_outputs(6865) <= a xor b;
    layer1_outputs(6866) <= b;
    layer1_outputs(6867) <= b;
    layer1_outputs(6868) <= not (a or b);
    layer1_outputs(6869) <= a xor b;
    layer1_outputs(6870) <= not a or b;
    layer1_outputs(6871) <= not (a xor b);
    layer1_outputs(6872) <= not a;
    layer1_outputs(6873) <= not a or b;
    layer1_outputs(6874) <= not (a or b);
    layer1_outputs(6875) <= not (a and b);
    layer1_outputs(6876) <= a or b;
    layer1_outputs(6877) <= not (a or b);
    layer1_outputs(6878) <= a;
    layer1_outputs(6879) <= a and not b;
    layer1_outputs(6880) <= a and b;
    layer1_outputs(6881) <= not a;
    layer1_outputs(6882) <= a;
    layer1_outputs(6883) <= not (a and b);
    layer1_outputs(6884) <= not (a xor b);
    layer1_outputs(6885) <= a and b;
    layer1_outputs(6886) <= not a;
    layer1_outputs(6887) <= not (a xor b);
    layer1_outputs(6888) <= not b;
    layer1_outputs(6889) <= not (a xor b);
    layer1_outputs(6890) <= not (a or b);
    layer1_outputs(6891) <= not (a xor b);
    layer1_outputs(6892) <= b and not a;
    layer1_outputs(6893) <= not (a and b);
    layer1_outputs(6894) <= not (a xor b);
    layer1_outputs(6895) <= b;
    layer1_outputs(6896) <= not (a xor b);
    layer1_outputs(6897) <= a;
    layer1_outputs(6898) <= not a;
    layer1_outputs(6899) <= b and not a;
    layer1_outputs(6900) <= b;
    layer1_outputs(6901) <= a or b;
    layer1_outputs(6902) <= not (a xor b);
    layer1_outputs(6903) <= b and not a;
    layer1_outputs(6904) <= a;
    layer1_outputs(6905) <= b and not a;
    layer1_outputs(6906) <= not a;
    layer1_outputs(6907) <= a xor b;
    layer1_outputs(6908) <= not a or b;
    layer1_outputs(6909) <= b;
    layer1_outputs(6910) <= not a or b;
    layer1_outputs(6911) <= not a;
    layer1_outputs(6912) <= a;
    layer1_outputs(6913) <= not b or a;
    layer1_outputs(6914) <= b;
    layer1_outputs(6915) <= a and not b;
    layer1_outputs(6916) <= a or b;
    layer1_outputs(6917) <= not a;
    layer1_outputs(6918) <= not (a and b);
    layer1_outputs(6919) <= not b;
    layer1_outputs(6920) <= a and b;
    layer1_outputs(6921) <= a;
    layer1_outputs(6922) <= not (a xor b);
    layer1_outputs(6923) <= not a or b;
    layer1_outputs(6924) <= not b;
    layer1_outputs(6925) <= b;
    layer1_outputs(6926) <= not (a or b);
    layer1_outputs(6927) <= b and not a;
    layer1_outputs(6928) <= not a or b;
    layer1_outputs(6929) <= b;
    layer1_outputs(6930) <= b and not a;
    layer1_outputs(6931) <= not a;
    layer1_outputs(6932) <= a or b;
    layer1_outputs(6933) <= not b or a;
    layer1_outputs(6934) <= not a;
    layer1_outputs(6935) <= not b or a;
    layer1_outputs(6936) <= b;
    layer1_outputs(6937) <= not a or b;
    layer1_outputs(6938) <= a and not b;
    layer1_outputs(6939) <= b;
    layer1_outputs(6940) <= not b;
    layer1_outputs(6941) <= not a or b;
    layer1_outputs(6942) <= b;
    layer1_outputs(6943) <= a;
    layer1_outputs(6944) <= not a;
    layer1_outputs(6945) <= not (a xor b);
    layer1_outputs(6946) <= not (a or b);
    layer1_outputs(6947) <= b and not a;
    layer1_outputs(6948) <= a and not b;
    layer1_outputs(6949) <= b and not a;
    layer1_outputs(6950) <= not a or b;
    layer1_outputs(6951) <= a;
    layer1_outputs(6952) <= a xor b;
    layer1_outputs(6953) <= not b;
    layer1_outputs(6954) <= not (a or b);
    layer1_outputs(6955) <= a and b;
    layer1_outputs(6956) <= not b or a;
    layer1_outputs(6957) <= a xor b;
    layer1_outputs(6958) <= not b or a;
    layer1_outputs(6959) <= not a;
    layer1_outputs(6960) <= b;
    layer1_outputs(6961) <= a;
    layer1_outputs(6962) <= a and not b;
    layer1_outputs(6963) <= not b;
    layer1_outputs(6964) <= not b;
    layer1_outputs(6965) <= b and not a;
    layer1_outputs(6966) <= not a or b;
    layer1_outputs(6967) <= '0';
    layer1_outputs(6968) <= a xor b;
    layer1_outputs(6969) <= b and not a;
    layer1_outputs(6970) <= b;
    layer1_outputs(6971) <= b and not a;
    layer1_outputs(6972) <= not b;
    layer1_outputs(6973) <= a xor b;
    layer1_outputs(6974) <= b;
    layer1_outputs(6975) <= not b or a;
    layer1_outputs(6976) <= a and not b;
    layer1_outputs(6977) <= not (a xor b);
    layer1_outputs(6978) <= not b;
    layer1_outputs(6979) <= b;
    layer1_outputs(6980) <= a xor b;
    layer1_outputs(6981) <= not (a and b);
    layer1_outputs(6982) <= not b;
    layer1_outputs(6983) <= a and b;
    layer1_outputs(6984) <= a or b;
    layer1_outputs(6985) <= a;
    layer1_outputs(6986) <= a xor b;
    layer1_outputs(6987) <= not (a and b);
    layer1_outputs(6988) <= not b or a;
    layer1_outputs(6989) <= not (a or b);
    layer1_outputs(6990) <= not b;
    layer1_outputs(6991) <= not b;
    layer1_outputs(6992) <= not b;
    layer1_outputs(6993) <= a and not b;
    layer1_outputs(6994) <= not (a and b);
    layer1_outputs(6995) <= a;
    layer1_outputs(6996) <= not b;
    layer1_outputs(6997) <= not (a or b);
    layer1_outputs(6998) <= a and b;
    layer1_outputs(6999) <= a xor b;
    layer1_outputs(7000) <= not b;
    layer1_outputs(7001) <= not a;
    layer1_outputs(7002) <= not b;
    layer1_outputs(7003) <= b;
    layer1_outputs(7004) <= b;
    layer1_outputs(7005) <= not b;
    layer1_outputs(7006) <= a;
    layer1_outputs(7007) <= b and not a;
    layer1_outputs(7008) <= not a or b;
    layer1_outputs(7009) <= b and not a;
    layer1_outputs(7010) <= not a;
    layer1_outputs(7011) <= a or b;
    layer1_outputs(7012) <= a and not b;
    layer1_outputs(7013) <= not (a xor b);
    layer1_outputs(7014) <= b;
    layer1_outputs(7015) <= b and not a;
    layer1_outputs(7016) <= not (a or b);
    layer1_outputs(7017) <= not (a and b);
    layer1_outputs(7018) <= b and not a;
    layer1_outputs(7019) <= a xor b;
    layer1_outputs(7020) <= not a or b;
    layer1_outputs(7021) <= not b or a;
    layer1_outputs(7022) <= not a or b;
    layer1_outputs(7023) <= not (a xor b);
    layer1_outputs(7024) <= not (a or b);
    layer1_outputs(7025) <= not a;
    layer1_outputs(7026) <= a;
    layer1_outputs(7027) <= not (a xor b);
    layer1_outputs(7028) <= b and not a;
    layer1_outputs(7029) <= not b;
    layer1_outputs(7030) <= not a or b;
    layer1_outputs(7031) <= a and b;
    layer1_outputs(7032) <= a and b;
    layer1_outputs(7033) <= a and not b;
    layer1_outputs(7034) <= a;
    layer1_outputs(7035) <= b;
    layer1_outputs(7036) <= not a or b;
    layer1_outputs(7037) <= b and not a;
    layer1_outputs(7038) <= a and not b;
    layer1_outputs(7039) <= a and not b;
    layer1_outputs(7040) <= a;
    layer1_outputs(7041) <= not b or a;
    layer1_outputs(7042) <= a and b;
    layer1_outputs(7043) <= not b or a;
    layer1_outputs(7044) <= b;
    layer1_outputs(7045) <= a xor b;
    layer1_outputs(7046) <= not b;
    layer1_outputs(7047) <= a xor b;
    layer1_outputs(7048) <= not (a xor b);
    layer1_outputs(7049) <= not (a xor b);
    layer1_outputs(7050) <= not a;
    layer1_outputs(7051) <= not (a xor b);
    layer1_outputs(7052) <= not b;
    layer1_outputs(7053) <= not b or a;
    layer1_outputs(7054) <= not a or b;
    layer1_outputs(7055) <= a and b;
    layer1_outputs(7056) <= b;
    layer1_outputs(7057) <= a;
    layer1_outputs(7058) <= not (a xor b);
    layer1_outputs(7059) <= a or b;
    layer1_outputs(7060) <= a and not b;
    layer1_outputs(7061) <= not a;
    layer1_outputs(7062) <= b;
    layer1_outputs(7063) <= not a or b;
    layer1_outputs(7064) <= a xor b;
    layer1_outputs(7065) <= not (a xor b);
    layer1_outputs(7066) <= not a;
    layer1_outputs(7067) <= a;
    layer1_outputs(7068) <= a xor b;
    layer1_outputs(7069) <= not b;
    layer1_outputs(7070) <= a xor b;
    layer1_outputs(7071) <= a xor b;
    layer1_outputs(7072) <= not b;
    layer1_outputs(7073) <= not b;
    layer1_outputs(7074) <= a xor b;
    layer1_outputs(7075) <= not a or b;
    layer1_outputs(7076) <= a and not b;
    layer1_outputs(7077) <= b and not a;
    layer1_outputs(7078) <= '1';
    layer1_outputs(7079) <= not (a xor b);
    layer1_outputs(7080) <= not (a and b);
    layer1_outputs(7081) <= '1';
    layer1_outputs(7082) <= not (a and b);
    layer1_outputs(7083) <= not b or a;
    layer1_outputs(7084) <= b;
    layer1_outputs(7085) <= b;
    layer1_outputs(7086) <= not b;
    layer1_outputs(7087) <= not a or b;
    layer1_outputs(7088) <= not a;
    layer1_outputs(7089) <= a;
    layer1_outputs(7090) <= '1';
    layer1_outputs(7091) <= not b;
    layer1_outputs(7092) <= b and not a;
    layer1_outputs(7093) <= b;
    layer1_outputs(7094) <= a and not b;
    layer1_outputs(7095) <= a;
    layer1_outputs(7096) <= a;
    layer1_outputs(7097) <= a;
    layer1_outputs(7098) <= not (a xor b);
    layer1_outputs(7099) <= b;
    layer1_outputs(7100) <= a;
    layer1_outputs(7101) <= a or b;
    layer1_outputs(7102) <= b;
    layer1_outputs(7103) <= not b;
    layer1_outputs(7104) <= not (a xor b);
    layer1_outputs(7105) <= a and b;
    layer1_outputs(7106) <= a and not b;
    layer1_outputs(7107) <= a and b;
    layer1_outputs(7108) <= not a;
    layer1_outputs(7109) <= a or b;
    layer1_outputs(7110) <= a;
    layer1_outputs(7111) <= not (a xor b);
    layer1_outputs(7112) <= b;
    layer1_outputs(7113) <= not a;
    layer1_outputs(7114) <= a;
    layer1_outputs(7115) <= b;
    layer1_outputs(7116) <= a or b;
    layer1_outputs(7117) <= a or b;
    layer1_outputs(7118) <= b and not a;
    layer1_outputs(7119) <= not b;
    layer1_outputs(7120) <= a and not b;
    layer1_outputs(7121) <= a xor b;
    layer1_outputs(7122) <= a or b;
    layer1_outputs(7123) <= not b;
    layer1_outputs(7124) <= a or b;
    layer1_outputs(7125) <= not (a or b);
    layer1_outputs(7126) <= not a;
    layer1_outputs(7127) <= not (a and b);
    layer1_outputs(7128) <= b;
    layer1_outputs(7129) <= a xor b;
    layer1_outputs(7130) <= b;
    layer1_outputs(7131) <= a;
    layer1_outputs(7132) <= a and b;
    layer1_outputs(7133) <= not a or b;
    layer1_outputs(7134) <= not b or a;
    layer1_outputs(7135) <= not (a xor b);
    layer1_outputs(7136) <= b and not a;
    layer1_outputs(7137) <= a and b;
    layer1_outputs(7138) <= a;
    layer1_outputs(7139) <= not a;
    layer1_outputs(7140) <= b;
    layer1_outputs(7141) <= not b;
    layer1_outputs(7142) <= not a;
    layer1_outputs(7143) <= a;
    layer1_outputs(7144) <= not (a and b);
    layer1_outputs(7145) <= not (a or b);
    layer1_outputs(7146) <= not a or b;
    layer1_outputs(7147) <= not (a and b);
    layer1_outputs(7148) <= '1';
    layer1_outputs(7149) <= a or b;
    layer1_outputs(7150) <= b and not a;
    layer1_outputs(7151) <= not (a xor b);
    layer1_outputs(7152) <= a and not b;
    layer1_outputs(7153) <= a or b;
    layer1_outputs(7154) <= a and not b;
    layer1_outputs(7155) <= '0';
    layer1_outputs(7156) <= not b;
    layer1_outputs(7157) <= b;
    layer1_outputs(7158) <= a xor b;
    layer1_outputs(7159) <= not (a and b);
    layer1_outputs(7160) <= not a or b;
    layer1_outputs(7161) <= a xor b;
    layer1_outputs(7162) <= not (a and b);
    layer1_outputs(7163) <= a and not b;
    layer1_outputs(7164) <= not a or b;
    layer1_outputs(7165) <= b and not a;
    layer1_outputs(7166) <= not b or a;
    layer1_outputs(7167) <= a or b;
    layer1_outputs(7168) <= '1';
    layer1_outputs(7169) <= a and b;
    layer1_outputs(7170) <= not (a or b);
    layer1_outputs(7171) <= a;
    layer1_outputs(7172) <= not b;
    layer1_outputs(7173) <= b;
    layer1_outputs(7174) <= b;
    layer1_outputs(7175) <= a or b;
    layer1_outputs(7176) <= not (a xor b);
    layer1_outputs(7177) <= not (a and b);
    layer1_outputs(7178) <= not b;
    layer1_outputs(7179) <= not a;
    layer1_outputs(7180) <= not (a or b);
    layer1_outputs(7181) <= b and not a;
    layer1_outputs(7182) <= '1';
    layer1_outputs(7183) <= not b or a;
    layer1_outputs(7184) <= b;
    layer1_outputs(7185) <= not (a xor b);
    layer1_outputs(7186) <= a and not b;
    layer1_outputs(7187) <= not b;
    layer1_outputs(7188) <= a;
    layer1_outputs(7189) <= a and b;
    layer1_outputs(7190) <= b;
    layer1_outputs(7191) <= a and not b;
    layer1_outputs(7192) <= a or b;
    layer1_outputs(7193) <= a and b;
    layer1_outputs(7194) <= a;
    layer1_outputs(7195) <= b;
    layer1_outputs(7196) <= a and b;
    layer1_outputs(7197) <= not (a or b);
    layer1_outputs(7198) <= '1';
    layer1_outputs(7199) <= not b;
    layer1_outputs(7200) <= a;
    layer1_outputs(7201) <= not (a or b);
    layer1_outputs(7202) <= a;
    layer1_outputs(7203) <= not a or b;
    layer1_outputs(7204) <= a xor b;
    layer1_outputs(7205) <= b;
    layer1_outputs(7206) <= not b;
    layer1_outputs(7207) <= not a or b;
    layer1_outputs(7208) <= a;
    layer1_outputs(7209) <= not (a xor b);
    layer1_outputs(7210) <= not b;
    layer1_outputs(7211) <= '1';
    layer1_outputs(7212) <= b;
    layer1_outputs(7213) <= b;
    layer1_outputs(7214) <= not a or b;
    layer1_outputs(7215) <= a;
    layer1_outputs(7216) <= not a;
    layer1_outputs(7217) <= not a;
    layer1_outputs(7218) <= not b;
    layer1_outputs(7219) <= not (a and b);
    layer1_outputs(7220) <= not (a or b);
    layer1_outputs(7221) <= a or b;
    layer1_outputs(7222) <= not a;
    layer1_outputs(7223) <= a and not b;
    layer1_outputs(7224) <= b and not a;
    layer1_outputs(7225) <= b;
    layer1_outputs(7226) <= a or b;
    layer1_outputs(7227) <= not b;
    layer1_outputs(7228) <= not (a xor b);
    layer1_outputs(7229) <= a;
    layer1_outputs(7230) <= a and not b;
    layer1_outputs(7231) <= not a;
    layer1_outputs(7232) <= '1';
    layer1_outputs(7233) <= a xor b;
    layer1_outputs(7234) <= not b;
    layer1_outputs(7235) <= not (a or b);
    layer1_outputs(7236) <= not a or b;
    layer1_outputs(7237) <= not (a or b);
    layer1_outputs(7238) <= not b or a;
    layer1_outputs(7239) <= not b or a;
    layer1_outputs(7240) <= not (a xor b);
    layer1_outputs(7241) <= a or b;
    layer1_outputs(7242) <= a and b;
    layer1_outputs(7243) <= a xor b;
    layer1_outputs(7244) <= not a;
    layer1_outputs(7245) <= not b or a;
    layer1_outputs(7246) <= b;
    layer1_outputs(7247) <= a and not b;
    layer1_outputs(7248) <= a and b;
    layer1_outputs(7249) <= b;
    layer1_outputs(7250) <= b and not a;
    layer1_outputs(7251) <= not (a or b);
    layer1_outputs(7252) <= a;
    layer1_outputs(7253) <= not (a and b);
    layer1_outputs(7254) <= '0';
    layer1_outputs(7255) <= not (a xor b);
    layer1_outputs(7256) <= a xor b;
    layer1_outputs(7257) <= b and not a;
    layer1_outputs(7258) <= not b or a;
    layer1_outputs(7259) <= b and not a;
    layer1_outputs(7260) <= a or b;
    layer1_outputs(7261) <= not a;
    layer1_outputs(7262) <= not (a and b);
    layer1_outputs(7263) <= not b;
    layer1_outputs(7264) <= a;
    layer1_outputs(7265) <= a;
    layer1_outputs(7266) <= not b;
    layer1_outputs(7267) <= a and not b;
    layer1_outputs(7268) <= b and not a;
    layer1_outputs(7269) <= b and not a;
    layer1_outputs(7270) <= a;
    layer1_outputs(7271) <= b;
    layer1_outputs(7272) <= a;
    layer1_outputs(7273) <= b and not a;
    layer1_outputs(7274) <= a and not b;
    layer1_outputs(7275) <= not b;
    layer1_outputs(7276) <= a xor b;
    layer1_outputs(7277) <= a;
    layer1_outputs(7278) <= b;
    layer1_outputs(7279) <= not a;
    layer1_outputs(7280) <= a;
    layer1_outputs(7281) <= b and not a;
    layer1_outputs(7282) <= not (a xor b);
    layer1_outputs(7283) <= a;
    layer1_outputs(7284) <= '1';
    layer1_outputs(7285) <= not b or a;
    layer1_outputs(7286) <= not b;
    layer1_outputs(7287) <= b and not a;
    layer1_outputs(7288) <= not a or b;
    layer1_outputs(7289) <= not a;
    layer1_outputs(7290) <= not (a and b);
    layer1_outputs(7291) <= not b;
    layer1_outputs(7292) <= b;
    layer1_outputs(7293) <= a and not b;
    layer1_outputs(7294) <= not b or a;
    layer1_outputs(7295) <= b and not a;
    layer1_outputs(7296) <= a;
    layer1_outputs(7297) <= a xor b;
    layer1_outputs(7298) <= b and not a;
    layer1_outputs(7299) <= '0';
    layer1_outputs(7300) <= not b;
    layer1_outputs(7301) <= not b or a;
    layer1_outputs(7302) <= not a;
    layer1_outputs(7303) <= not a;
    layer1_outputs(7304) <= b;
    layer1_outputs(7305) <= b;
    layer1_outputs(7306) <= not (a or b);
    layer1_outputs(7307) <= a and b;
    layer1_outputs(7308) <= a xor b;
    layer1_outputs(7309) <= b;
    layer1_outputs(7310) <= a or b;
    layer1_outputs(7311) <= not a;
    layer1_outputs(7312) <= b;
    layer1_outputs(7313) <= b;
    layer1_outputs(7314) <= not a;
    layer1_outputs(7315) <= a;
    layer1_outputs(7316) <= not (a or b);
    layer1_outputs(7317) <= b;
    layer1_outputs(7318) <= b;
    layer1_outputs(7319) <= not b;
    layer1_outputs(7320) <= b and not a;
    layer1_outputs(7321) <= not a;
    layer1_outputs(7322) <= not b;
    layer1_outputs(7323) <= not (a xor b);
    layer1_outputs(7324) <= not (a xor b);
    layer1_outputs(7325) <= not b;
    layer1_outputs(7326) <= a;
    layer1_outputs(7327) <= a and b;
    layer1_outputs(7328) <= a;
    layer1_outputs(7329) <= not (a and b);
    layer1_outputs(7330) <= not (a or b);
    layer1_outputs(7331) <= a;
    layer1_outputs(7332) <= b and not a;
    layer1_outputs(7333) <= not b or a;
    layer1_outputs(7334) <= b;
    layer1_outputs(7335) <= b;
    layer1_outputs(7336) <= not (a or b);
    layer1_outputs(7337) <= a and b;
    layer1_outputs(7338) <= not b;
    layer1_outputs(7339) <= a xor b;
    layer1_outputs(7340) <= not (a and b);
    layer1_outputs(7341) <= b;
    layer1_outputs(7342) <= not (a xor b);
    layer1_outputs(7343) <= not a or b;
    layer1_outputs(7344) <= a and not b;
    layer1_outputs(7345) <= b;
    layer1_outputs(7346) <= not (a and b);
    layer1_outputs(7347) <= b;
    layer1_outputs(7348) <= not (a or b);
    layer1_outputs(7349) <= not (a or b);
    layer1_outputs(7350) <= a xor b;
    layer1_outputs(7351) <= a xor b;
    layer1_outputs(7352) <= a or b;
    layer1_outputs(7353) <= not (a xor b);
    layer1_outputs(7354) <= b and not a;
    layer1_outputs(7355) <= a or b;
    layer1_outputs(7356) <= a and b;
    layer1_outputs(7357) <= a or b;
    layer1_outputs(7358) <= a;
    layer1_outputs(7359) <= a or b;
    layer1_outputs(7360) <= '1';
    layer1_outputs(7361) <= not a or b;
    layer1_outputs(7362) <= not (a or b);
    layer1_outputs(7363) <= not (a and b);
    layer1_outputs(7364) <= not b or a;
    layer1_outputs(7365) <= a and not b;
    layer1_outputs(7366) <= b;
    layer1_outputs(7367) <= a;
    layer1_outputs(7368) <= b;
    layer1_outputs(7369) <= b;
    layer1_outputs(7370) <= a;
    layer1_outputs(7371) <= not (a and b);
    layer1_outputs(7372) <= b;
    layer1_outputs(7373) <= a and not b;
    layer1_outputs(7374) <= a xor b;
    layer1_outputs(7375) <= a or b;
    layer1_outputs(7376) <= b;
    layer1_outputs(7377) <= not b;
    layer1_outputs(7378) <= a and not b;
    layer1_outputs(7379) <= b;
    layer1_outputs(7380) <= not a;
    layer1_outputs(7381) <= b and not a;
    layer1_outputs(7382) <= b;
    layer1_outputs(7383) <= not a or b;
    layer1_outputs(7384) <= b and not a;
    layer1_outputs(7385) <= not b;
    layer1_outputs(7386) <= a or b;
    layer1_outputs(7387) <= not (a xor b);
    layer1_outputs(7388) <= not b;
    layer1_outputs(7389) <= a and not b;
    layer1_outputs(7390) <= not (a and b);
    layer1_outputs(7391) <= not b or a;
    layer1_outputs(7392) <= a xor b;
    layer1_outputs(7393) <= a xor b;
    layer1_outputs(7394) <= not (a xor b);
    layer1_outputs(7395) <= a and not b;
    layer1_outputs(7396) <= a and not b;
    layer1_outputs(7397) <= a or b;
    layer1_outputs(7398) <= a and not b;
    layer1_outputs(7399) <= b;
    layer1_outputs(7400) <= not (a and b);
    layer1_outputs(7401) <= not (a and b);
    layer1_outputs(7402) <= a or b;
    layer1_outputs(7403) <= not (a xor b);
    layer1_outputs(7404) <= a and b;
    layer1_outputs(7405) <= not a;
    layer1_outputs(7406) <= b and not a;
    layer1_outputs(7407) <= not (a xor b);
    layer1_outputs(7408) <= not a;
    layer1_outputs(7409) <= a;
    layer1_outputs(7410) <= not a or b;
    layer1_outputs(7411) <= not (a or b);
    layer1_outputs(7412) <= b and not a;
    layer1_outputs(7413) <= not (a or b);
    layer1_outputs(7414) <= a or b;
    layer1_outputs(7415) <= not a;
    layer1_outputs(7416) <= not (a xor b);
    layer1_outputs(7417) <= a or b;
    layer1_outputs(7418) <= a xor b;
    layer1_outputs(7419) <= not (a or b);
    layer1_outputs(7420) <= a and b;
    layer1_outputs(7421) <= b;
    layer1_outputs(7422) <= b;
    layer1_outputs(7423) <= a and b;
    layer1_outputs(7424) <= a and not b;
    layer1_outputs(7425) <= a;
    layer1_outputs(7426) <= a or b;
    layer1_outputs(7427) <= a;
    layer1_outputs(7428) <= not b or a;
    layer1_outputs(7429) <= b;
    layer1_outputs(7430) <= a xor b;
    layer1_outputs(7431) <= not (a and b);
    layer1_outputs(7432) <= not a or b;
    layer1_outputs(7433) <= not (a and b);
    layer1_outputs(7434) <= not b or a;
    layer1_outputs(7435) <= a;
    layer1_outputs(7436) <= not (a or b);
    layer1_outputs(7437) <= a and b;
    layer1_outputs(7438) <= a xor b;
    layer1_outputs(7439) <= not a;
    layer1_outputs(7440) <= '1';
    layer1_outputs(7441) <= a;
    layer1_outputs(7442) <= a and not b;
    layer1_outputs(7443) <= a and b;
    layer1_outputs(7444) <= not a or b;
    layer1_outputs(7445) <= a and b;
    layer1_outputs(7446) <= not a;
    layer1_outputs(7447) <= a;
    layer1_outputs(7448) <= not a or b;
    layer1_outputs(7449) <= b;
    layer1_outputs(7450) <= b and not a;
    layer1_outputs(7451) <= a;
    layer1_outputs(7452) <= not a;
    layer1_outputs(7453) <= a and b;
    layer1_outputs(7454) <= b and not a;
    layer1_outputs(7455) <= not (a or b);
    layer1_outputs(7456) <= a or b;
    layer1_outputs(7457) <= not a;
    layer1_outputs(7458) <= not a or b;
    layer1_outputs(7459) <= b;
    layer1_outputs(7460) <= not (a or b);
    layer1_outputs(7461) <= b and not a;
    layer1_outputs(7462) <= not b or a;
    layer1_outputs(7463) <= not a;
    layer1_outputs(7464) <= not a or b;
    layer1_outputs(7465) <= not b;
    layer1_outputs(7466) <= '1';
    layer1_outputs(7467) <= a and b;
    layer1_outputs(7468) <= not (a and b);
    layer1_outputs(7469) <= b and not a;
    layer1_outputs(7470) <= not b;
    layer1_outputs(7471) <= a and b;
    layer1_outputs(7472) <= b;
    layer1_outputs(7473) <= not a or b;
    layer1_outputs(7474) <= a;
    layer1_outputs(7475) <= a or b;
    layer1_outputs(7476) <= not (a xor b);
    layer1_outputs(7477) <= not a;
    layer1_outputs(7478) <= a;
    layer1_outputs(7479) <= a and b;
    layer1_outputs(7480) <= not (a and b);
    layer1_outputs(7481) <= b;
    layer1_outputs(7482) <= a xor b;
    layer1_outputs(7483) <= not a;
    layer1_outputs(7484) <= not a or b;
    layer1_outputs(7485) <= a xor b;
    layer1_outputs(7486) <= not (a or b);
    layer1_outputs(7487) <= b and not a;
    layer1_outputs(7488) <= not b;
    layer1_outputs(7489) <= not b or a;
    layer1_outputs(7490) <= not a or b;
    layer1_outputs(7491) <= not a or b;
    layer1_outputs(7492) <= a or b;
    layer1_outputs(7493) <= not (a xor b);
    layer1_outputs(7494) <= not a or b;
    layer1_outputs(7495) <= not a or b;
    layer1_outputs(7496) <= a and not b;
    layer1_outputs(7497) <= not a;
    layer1_outputs(7498) <= not b or a;
    layer1_outputs(7499) <= b;
    layer1_outputs(7500) <= a and b;
    layer1_outputs(7501) <= not b;
    layer1_outputs(7502) <= a and b;
    layer1_outputs(7503) <= a;
    layer1_outputs(7504) <= a and not b;
    layer1_outputs(7505) <= not a;
    layer1_outputs(7506) <= not b or a;
    layer1_outputs(7507) <= a;
    layer1_outputs(7508) <= a and b;
    layer1_outputs(7509) <= not (a and b);
    layer1_outputs(7510) <= not (a or b);
    layer1_outputs(7511) <= not a;
    layer1_outputs(7512) <= b and not a;
    layer1_outputs(7513) <= b and not a;
    layer1_outputs(7514) <= not b;
    layer1_outputs(7515) <= a and b;
    layer1_outputs(7516) <= not a or b;
    layer1_outputs(7517) <= not (a or b);
    layer1_outputs(7518) <= not a;
    layer1_outputs(7519) <= not (a or b);
    layer1_outputs(7520) <= b and not a;
    layer1_outputs(7521) <= b;
    layer1_outputs(7522) <= a and not b;
    layer1_outputs(7523) <= a;
    layer1_outputs(7524) <= not a or b;
    layer1_outputs(7525) <= a;
    layer1_outputs(7526) <= not (a xor b);
    layer1_outputs(7527) <= a and b;
    layer1_outputs(7528) <= not b or a;
    layer1_outputs(7529) <= a and not b;
    layer1_outputs(7530) <= a xor b;
    layer1_outputs(7531) <= b;
    layer1_outputs(7532) <= a and b;
    layer1_outputs(7533) <= not a or b;
    layer1_outputs(7534) <= a xor b;
    layer1_outputs(7535) <= a;
    layer1_outputs(7536) <= not (a and b);
    layer1_outputs(7537) <= a xor b;
    layer1_outputs(7538) <= not b or a;
    layer1_outputs(7539) <= not b or a;
    layer1_outputs(7540) <= a and not b;
    layer1_outputs(7541) <= a or b;
    layer1_outputs(7542) <= a or b;
    layer1_outputs(7543) <= a and b;
    layer1_outputs(7544) <= a;
    layer1_outputs(7545) <= a;
    layer1_outputs(7546) <= a xor b;
    layer1_outputs(7547) <= not a;
    layer1_outputs(7548) <= not a or b;
    layer1_outputs(7549) <= not a or b;
    layer1_outputs(7550) <= a or b;
    layer1_outputs(7551) <= not b;
    layer1_outputs(7552) <= not (a or b);
    layer1_outputs(7553) <= a;
    layer1_outputs(7554) <= not b;
    layer1_outputs(7555) <= a or b;
    layer1_outputs(7556) <= a or b;
    layer1_outputs(7557) <= a xor b;
    layer1_outputs(7558) <= not b or a;
    layer1_outputs(7559) <= b and not a;
    layer1_outputs(7560) <= a xor b;
    layer1_outputs(7561) <= b;
    layer1_outputs(7562) <= b;
    layer1_outputs(7563) <= not b or a;
    layer1_outputs(7564) <= not (a and b);
    layer1_outputs(7565) <= not b;
    layer1_outputs(7566) <= not a or b;
    layer1_outputs(7567) <= not b;
    layer1_outputs(7568) <= not a;
    layer1_outputs(7569) <= a and not b;
    layer1_outputs(7570) <= not (a xor b);
    layer1_outputs(7571) <= b and not a;
    layer1_outputs(7572) <= not (a or b);
    layer1_outputs(7573) <= a;
    layer1_outputs(7574) <= a;
    layer1_outputs(7575) <= not (a or b);
    layer1_outputs(7576) <= not b;
    layer1_outputs(7577) <= b and not a;
    layer1_outputs(7578) <= not (a and b);
    layer1_outputs(7579) <= b;
    layer1_outputs(7580) <= a and not b;
    layer1_outputs(7581) <= a;
    layer1_outputs(7582) <= a;
    layer1_outputs(7583) <= a;
    layer1_outputs(7584) <= not b;
    layer1_outputs(7585) <= not b;
    layer1_outputs(7586) <= a;
    layer1_outputs(7587) <= a and not b;
    layer1_outputs(7588) <= b and not a;
    layer1_outputs(7589) <= b;
    layer1_outputs(7590) <= not (a or b);
    layer1_outputs(7591) <= not a;
    layer1_outputs(7592) <= a or b;
    layer1_outputs(7593) <= b;
    layer1_outputs(7594) <= b;
    layer1_outputs(7595) <= not (a or b);
    layer1_outputs(7596) <= a xor b;
    layer1_outputs(7597) <= a or b;
    layer1_outputs(7598) <= not (a and b);
    layer1_outputs(7599) <= not (a xor b);
    layer1_outputs(7600) <= not b;
    layer1_outputs(7601) <= not b;
    layer1_outputs(7602) <= a or b;
    layer1_outputs(7603) <= a and b;
    layer1_outputs(7604) <= not (a and b);
    layer1_outputs(7605) <= not (a xor b);
    layer1_outputs(7606) <= not (a xor b);
    layer1_outputs(7607) <= not b;
    layer1_outputs(7608) <= a or b;
    layer1_outputs(7609) <= not (a xor b);
    layer1_outputs(7610) <= not (a or b);
    layer1_outputs(7611) <= a and not b;
    layer1_outputs(7612) <= b and not a;
    layer1_outputs(7613) <= a;
    layer1_outputs(7614) <= a and not b;
    layer1_outputs(7615) <= a;
    layer1_outputs(7616) <= b;
    layer1_outputs(7617) <= b and not a;
    layer1_outputs(7618) <= a and b;
    layer1_outputs(7619) <= a and b;
    layer1_outputs(7620) <= b;
    layer1_outputs(7621) <= b and not a;
    layer1_outputs(7622) <= not (a xor b);
    layer1_outputs(7623) <= b;
    layer1_outputs(7624) <= a;
    layer1_outputs(7625) <= b and not a;
    layer1_outputs(7626) <= not a;
    layer1_outputs(7627) <= not (a or b);
    layer1_outputs(7628) <= b;
    layer1_outputs(7629) <= a and b;
    layer1_outputs(7630) <= not b or a;
    layer1_outputs(7631) <= not (a or b);
    layer1_outputs(7632) <= a or b;
    layer1_outputs(7633) <= not (a and b);
    layer1_outputs(7634) <= a;
    layer1_outputs(7635) <= not a;
    layer1_outputs(7636) <= a;
    layer1_outputs(7637) <= not (a and b);
    layer1_outputs(7638) <= not b or a;
    layer1_outputs(7639) <= b;
    layer1_outputs(7640) <= b;
    layer1_outputs(7641) <= not (a and b);
    layer1_outputs(7642) <= a;
    layer1_outputs(7643) <= a and b;
    layer1_outputs(7644) <= b and not a;
    layer1_outputs(7645) <= not b;
    layer1_outputs(7646) <= a or b;
    layer1_outputs(7647) <= b and not a;
    layer1_outputs(7648) <= not (a xor b);
    layer1_outputs(7649) <= a and not b;
    layer1_outputs(7650) <= b;
    layer1_outputs(7651) <= b and not a;
    layer1_outputs(7652) <= not a or b;
    layer1_outputs(7653) <= not (a and b);
    layer1_outputs(7654) <= b;
    layer1_outputs(7655) <= not a;
    layer1_outputs(7656) <= not b;
    layer1_outputs(7657) <= a xor b;
    layer1_outputs(7658) <= not (a or b);
    layer1_outputs(7659) <= a xor b;
    layer1_outputs(7660) <= b and not a;
    layer1_outputs(7661) <= a and not b;
    layer1_outputs(7662) <= b and not a;
    layer1_outputs(7663) <= a and b;
    layer1_outputs(7664) <= b;
    layer1_outputs(7665) <= b and not a;
    layer1_outputs(7666) <= not (a or b);
    layer1_outputs(7667) <= a;
    layer1_outputs(7668) <= not a;
    layer1_outputs(7669) <= not a or b;
    layer1_outputs(7670) <= not a;
    layer1_outputs(7671) <= b;
    layer1_outputs(7672) <= a xor b;
    layer1_outputs(7673) <= not (a or b);
    layer1_outputs(7674) <= not b;
    layer1_outputs(7675) <= b and not a;
    layer1_outputs(7676) <= a and not b;
    layer1_outputs(7677) <= not (a and b);
    layer1_outputs(7678) <= a;
    layer1_outputs(7679) <= a xor b;
    layer1_outputs(7680) <= a or b;
    layer1_outputs(7681) <= not b or a;
    layer1_outputs(7682) <= not b;
    layer1_outputs(7683) <= not (a xor b);
    layer1_outputs(7684) <= a xor b;
    layer1_outputs(7685) <= a and not b;
    layer1_outputs(7686) <= not (a and b);
    layer1_outputs(7687) <= a;
    layer1_outputs(7688) <= a and b;
    layer1_outputs(7689) <= not (a or b);
    layer1_outputs(7690) <= a;
    layer1_outputs(7691) <= a xor b;
    layer1_outputs(7692) <= a and b;
    layer1_outputs(7693) <= b and not a;
    layer1_outputs(7694) <= not (a xor b);
    layer1_outputs(7695) <= a or b;
    layer1_outputs(7696) <= not b or a;
    layer1_outputs(7697) <= not (a and b);
    layer1_outputs(7698) <= a and not b;
    layer1_outputs(7699) <= a;
    layer1_outputs(7700) <= b and not a;
    layer1_outputs(7701) <= a xor b;
    layer1_outputs(7702) <= not a or b;
    layer1_outputs(7703) <= a;
    layer1_outputs(7704) <= not (a xor b);
    layer1_outputs(7705) <= not b;
    layer1_outputs(7706) <= not a;
    layer1_outputs(7707) <= a and not b;
    layer1_outputs(7708) <= not b or a;
    layer1_outputs(7709) <= not b or a;
    layer1_outputs(7710) <= not (a xor b);
    layer1_outputs(7711) <= not a;
    layer1_outputs(7712) <= b;
    layer1_outputs(7713) <= '0';
    layer1_outputs(7714) <= not (a or b);
    layer1_outputs(7715) <= '1';
    layer1_outputs(7716) <= a;
    layer1_outputs(7717) <= not a;
    layer1_outputs(7718) <= not (a xor b);
    layer1_outputs(7719) <= not (a xor b);
    layer1_outputs(7720) <= b;
    layer1_outputs(7721) <= a;
    layer1_outputs(7722) <= a or b;
    layer1_outputs(7723) <= not b or a;
    layer1_outputs(7724) <= a and not b;
    layer1_outputs(7725) <= a;
    layer1_outputs(7726) <= not (a or b);
    layer1_outputs(7727) <= not a or b;
    layer1_outputs(7728) <= a xor b;
    layer1_outputs(7729) <= not (a xor b);
    layer1_outputs(7730) <= a or b;
    layer1_outputs(7731) <= not b;
    layer1_outputs(7732) <= not b;
    layer1_outputs(7733) <= not b or a;
    layer1_outputs(7734) <= not (a or b);
    layer1_outputs(7735) <= b and not a;
    layer1_outputs(7736) <= a and b;
    layer1_outputs(7737) <= b;
    layer1_outputs(7738) <= not (a and b);
    layer1_outputs(7739) <= not a;
    layer1_outputs(7740) <= a and not b;
    layer1_outputs(7741) <= not (a xor b);
    layer1_outputs(7742) <= a or b;
    layer1_outputs(7743) <= a;
    layer1_outputs(7744) <= a and b;
    layer1_outputs(7745) <= not b;
    layer1_outputs(7746) <= b;
    layer1_outputs(7747) <= a xor b;
    layer1_outputs(7748) <= not b;
    layer1_outputs(7749) <= b;
    layer1_outputs(7750) <= b;
    layer1_outputs(7751) <= not b;
    layer1_outputs(7752) <= a and not b;
    layer1_outputs(7753) <= a and b;
    layer1_outputs(7754) <= b and not a;
    layer1_outputs(7755) <= a and b;
    layer1_outputs(7756) <= a;
    layer1_outputs(7757) <= not a or b;
    layer1_outputs(7758) <= b;
    layer1_outputs(7759) <= not b;
    layer1_outputs(7760) <= not b;
    layer1_outputs(7761) <= not a;
    layer1_outputs(7762) <= not a;
    layer1_outputs(7763) <= not b;
    layer1_outputs(7764) <= a and b;
    layer1_outputs(7765) <= not (a and b);
    layer1_outputs(7766) <= not (a or b);
    layer1_outputs(7767) <= not b;
    layer1_outputs(7768) <= a or b;
    layer1_outputs(7769) <= not (a xor b);
    layer1_outputs(7770) <= a and b;
    layer1_outputs(7771) <= b;
    layer1_outputs(7772) <= not a;
    layer1_outputs(7773) <= b;
    layer1_outputs(7774) <= a or b;
    layer1_outputs(7775) <= not a;
    layer1_outputs(7776) <= a and b;
    layer1_outputs(7777) <= not a;
    layer1_outputs(7778) <= a and b;
    layer1_outputs(7779) <= b and not a;
    layer1_outputs(7780) <= not (a xor b);
    layer1_outputs(7781) <= a;
    layer1_outputs(7782) <= not b;
    layer1_outputs(7783) <= not a or b;
    layer1_outputs(7784) <= not a;
    layer1_outputs(7785) <= not (a and b);
    layer1_outputs(7786) <= not a;
    layer1_outputs(7787) <= a and not b;
    layer1_outputs(7788) <= b;
    layer1_outputs(7789) <= a;
    layer1_outputs(7790) <= b;
    layer1_outputs(7791) <= b;
    layer1_outputs(7792) <= not (a xor b);
    layer1_outputs(7793) <= not b;
    layer1_outputs(7794) <= a and b;
    layer1_outputs(7795) <= a;
    layer1_outputs(7796) <= not a;
    layer1_outputs(7797) <= a;
    layer1_outputs(7798) <= b and not a;
    layer1_outputs(7799) <= a;
    layer1_outputs(7800) <= '0';
    layer1_outputs(7801) <= a;
    layer1_outputs(7802) <= b and not a;
    layer1_outputs(7803) <= a;
    layer1_outputs(7804) <= not b;
    layer1_outputs(7805) <= b and not a;
    layer1_outputs(7806) <= not b;
    layer1_outputs(7807) <= a and b;
    layer1_outputs(7808) <= b;
    layer1_outputs(7809) <= b;
    layer1_outputs(7810) <= not (a or b);
    layer1_outputs(7811) <= a and not b;
    layer1_outputs(7812) <= a or b;
    layer1_outputs(7813) <= not (a xor b);
    layer1_outputs(7814) <= a;
    layer1_outputs(7815) <= a xor b;
    layer1_outputs(7816) <= a and not b;
    layer1_outputs(7817) <= not a;
    layer1_outputs(7818) <= not a;
    layer1_outputs(7819) <= a and b;
    layer1_outputs(7820) <= not (a xor b);
    layer1_outputs(7821) <= b and not a;
    layer1_outputs(7822) <= b;
    layer1_outputs(7823) <= not (a or b);
    layer1_outputs(7824) <= not a;
    layer1_outputs(7825) <= a or b;
    layer1_outputs(7826) <= b;
    layer1_outputs(7827) <= not b or a;
    layer1_outputs(7828) <= a and b;
    layer1_outputs(7829) <= not a or b;
    layer1_outputs(7830) <= not a;
    layer1_outputs(7831) <= not b or a;
    layer1_outputs(7832) <= a and not b;
    layer1_outputs(7833) <= not a;
    layer1_outputs(7834) <= not a;
    layer1_outputs(7835) <= a;
    layer1_outputs(7836) <= not b or a;
    layer1_outputs(7837) <= a and b;
    layer1_outputs(7838) <= not (a or b);
    layer1_outputs(7839) <= not (a xor b);
    layer1_outputs(7840) <= not (a xor b);
    layer1_outputs(7841) <= a and b;
    layer1_outputs(7842) <= not b;
    layer1_outputs(7843) <= a;
    layer1_outputs(7844) <= not a or b;
    layer1_outputs(7845) <= a or b;
    layer1_outputs(7846) <= not b;
    layer1_outputs(7847) <= a or b;
    layer1_outputs(7848) <= not a or b;
    layer1_outputs(7849) <= not b;
    layer1_outputs(7850) <= not a or b;
    layer1_outputs(7851) <= not (a xor b);
    layer1_outputs(7852) <= a and b;
    layer1_outputs(7853) <= not b or a;
    layer1_outputs(7854) <= not (a xor b);
    layer1_outputs(7855) <= not a;
    layer1_outputs(7856) <= not b;
    layer1_outputs(7857) <= not a;
    layer1_outputs(7858) <= not b;
    layer1_outputs(7859) <= not a;
    layer1_outputs(7860) <= not (a or b);
    layer1_outputs(7861) <= not a;
    layer1_outputs(7862) <= not a or b;
    layer1_outputs(7863) <= not (a xor b);
    layer1_outputs(7864) <= a;
    layer1_outputs(7865) <= not (a xor b);
    layer1_outputs(7866) <= not b or a;
    layer1_outputs(7867) <= b;
    layer1_outputs(7868) <= not a;
    layer1_outputs(7869) <= b and not a;
    layer1_outputs(7870) <= not (a or b);
    layer1_outputs(7871) <= not (a and b);
    layer1_outputs(7872) <= not (a or b);
    layer1_outputs(7873) <= not (a xor b);
    layer1_outputs(7874) <= b;
    layer1_outputs(7875) <= b;
    layer1_outputs(7876) <= not b;
    layer1_outputs(7877) <= not a;
    layer1_outputs(7878) <= b;
    layer1_outputs(7879) <= not (a or b);
    layer1_outputs(7880) <= not b or a;
    layer1_outputs(7881) <= not (a and b);
    layer1_outputs(7882) <= not a or b;
    layer1_outputs(7883) <= b;
    layer1_outputs(7884) <= a xor b;
    layer1_outputs(7885) <= b;
    layer1_outputs(7886) <= not a or b;
    layer1_outputs(7887) <= not b or a;
    layer1_outputs(7888) <= '0';
    layer1_outputs(7889) <= not b;
    layer1_outputs(7890) <= not (a xor b);
    layer1_outputs(7891) <= not b;
    layer1_outputs(7892) <= a and not b;
    layer1_outputs(7893) <= not (a and b);
    layer1_outputs(7894) <= b and not a;
    layer1_outputs(7895) <= not a;
    layer1_outputs(7896) <= a and b;
    layer1_outputs(7897) <= not (a or b);
    layer1_outputs(7898) <= not a;
    layer1_outputs(7899) <= a or b;
    layer1_outputs(7900) <= b;
    layer1_outputs(7901) <= b and not a;
    layer1_outputs(7902) <= not (a xor b);
    layer1_outputs(7903) <= a xor b;
    layer1_outputs(7904) <= not (a and b);
    layer1_outputs(7905) <= not a;
    layer1_outputs(7906) <= not a or b;
    layer1_outputs(7907) <= a or b;
    layer1_outputs(7908) <= not a or b;
    layer1_outputs(7909) <= not b;
    layer1_outputs(7910) <= a xor b;
    layer1_outputs(7911) <= a;
    layer1_outputs(7912) <= not a or b;
    layer1_outputs(7913) <= not (a and b);
    layer1_outputs(7914) <= a or b;
    layer1_outputs(7915) <= not b;
    layer1_outputs(7916) <= a xor b;
    layer1_outputs(7917) <= b;
    layer1_outputs(7918) <= a;
    layer1_outputs(7919) <= not a;
    layer1_outputs(7920) <= a;
    layer1_outputs(7921) <= not (a and b);
    layer1_outputs(7922) <= not (a xor b);
    layer1_outputs(7923) <= not b;
    layer1_outputs(7924) <= not a;
    layer1_outputs(7925) <= b;
    layer1_outputs(7926) <= not (a or b);
    layer1_outputs(7927) <= b;
    layer1_outputs(7928) <= b and not a;
    layer1_outputs(7929) <= not (a xor b);
    layer1_outputs(7930) <= not a or b;
    layer1_outputs(7931) <= a;
    layer1_outputs(7932) <= not a;
    layer1_outputs(7933) <= not b;
    layer1_outputs(7934) <= not b or a;
    layer1_outputs(7935) <= a xor b;
    layer1_outputs(7936) <= a or b;
    layer1_outputs(7937) <= not (a or b);
    layer1_outputs(7938) <= b;
    layer1_outputs(7939) <= not b;
    layer1_outputs(7940) <= a and not b;
    layer1_outputs(7941) <= not a or b;
    layer1_outputs(7942) <= a xor b;
    layer1_outputs(7943) <= not b;
    layer1_outputs(7944) <= a;
    layer1_outputs(7945) <= a;
    layer1_outputs(7946) <= not (a xor b);
    layer1_outputs(7947) <= not (a and b);
    layer1_outputs(7948) <= a;
    layer1_outputs(7949) <= not a or b;
    layer1_outputs(7950) <= not (a or b);
    layer1_outputs(7951) <= a or b;
    layer1_outputs(7952) <= not (a or b);
    layer1_outputs(7953) <= not (a and b);
    layer1_outputs(7954) <= not b;
    layer1_outputs(7955) <= not a;
    layer1_outputs(7956) <= not b or a;
    layer1_outputs(7957) <= not b or a;
    layer1_outputs(7958) <= not a or b;
    layer1_outputs(7959) <= a;
    layer1_outputs(7960) <= b and not a;
    layer1_outputs(7961) <= a xor b;
    layer1_outputs(7962) <= b;
    layer1_outputs(7963) <= a and not b;
    layer1_outputs(7964) <= '1';
    layer1_outputs(7965) <= a;
    layer1_outputs(7966) <= not (a xor b);
    layer1_outputs(7967) <= a and not b;
    layer1_outputs(7968) <= '1';
    layer1_outputs(7969) <= a or b;
    layer1_outputs(7970) <= b and not a;
    layer1_outputs(7971) <= b and not a;
    layer1_outputs(7972) <= a;
    layer1_outputs(7973) <= b;
    layer1_outputs(7974) <= not (a or b);
    layer1_outputs(7975) <= not (a xor b);
    layer1_outputs(7976) <= not a;
    layer1_outputs(7977) <= a;
    layer1_outputs(7978) <= not (a xor b);
    layer1_outputs(7979) <= b;
    layer1_outputs(7980) <= not (a xor b);
    layer1_outputs(7981) <= b and not a;
    layer1_outputs(7982) <= not b;
    layer1_outputs(7983) <= b;
    layer1_outputs(7984) <= not b or a;
    layer1_outputs(7985) <= not a or b;
    layer1_outputs(7986) <= a and not b;
    layer1_outputs(7987) <= a;
    layer1_outputs(7988) <= not a or b;
    layer1_outputs(7989) <= a and not b;
    layer1_outputs(7990) <= '0';
    layer1_outputs(7991) <= a and b;
    layer1_outputs(7992) <= a;
    layer1_outputs(7993) <= not a;
    layer1_outputs(7994) <= not (a or b);
    layer1_outputs(7995) <= not (a or b);
    layer1_outputs(7996) <= a or b;
    layer1_outputs(7997) <= b and not a;
    layer1_outputs(7998) <= a and not b;
    layer1_outputs(7999) <= '1';
    layer1_outputs(8000) <= '1';
    layer1_outputs(8001) <= not b;
    layer1_outputs(8002) <= a and not b;
    layer1_outputs(8003) <= not b or a;
    layer1_outputs(8004) <= a;
    layer1_outputs(8005) <= not b or a;
    layer1_outputs(8006) <= not (a xor b);
    layer1_outputs(8007) <= b;
    layer1_outputs(8008) <= '1';
    layer1_outputs(8009) <= a and b;
    layer1_outputs(8010) <= b and not a;
    layer1_outputs(8011) <= not (a xor b);
    layer1_outputs(8012) <= not b or a;
    layer1_outputs(8013) <= not (a xor b);
    layer1_outputs(8014) <= b;
    layer1_outputs(8015) <= not b;
    layer1_outputs(8016) <= not a or b;
    layer1_outputs(8017) <= a;
    layer1_outputs(8018) <= not (a or b);
    layer1_outputs(8019) <= not b;
    layer1_outputs(8020) <= a;
    layer1_outputs(8021) <= b;
    layer1_outputs(8022) <= a or b;
    layer1_outputs(8023) <= not (a or b);
    layer1_outputs(8024) <= not a;
    layer1_outputs(8025) <= not a;
    layer1_outputs(8026) <= not (a or b);
    layer1_outputs(8027) <= not b or a;
    layer1_outputs(8028) <= not (a or b);
    layer1_outputs(8029) <= not (a or b);
    layer1_outputs(8030) <= a or b;
    layer1_outputs(8031) <= a and not b;
    layer1_outputs(8032) <= not (a or b);
    layer1_outputs(8033) <= not a or b;
    layer1_outputs(8034) <= not (a and b);
    layer1_outputs(8035) <= not (a xor b);
    layer1_outputs(8036) <= not (a or b);
    layer1_outputs(8037) <= a;
    layer1_outputs(8038) <= not b or a;
    layer1_outputs(8039) <= not b or a;
    layer1_outputs(8040) <= a xor b;
    layer1_outputs(8041) <= not (a and b);
    layer1_outputs(8042) <= not a;
    layer1_outputs(8043) <= b and not a;
    layer1_outputs(8044) <= b;
    layer1_outputs(8045) <= not (a xor b);
    layer1_outputs(8046) <= a and not b;
    layer1_outputs(8047) <= b;
    layer1_outputs(8048) <= b and not a;
    layer1_outputs(8049) <= not b or a;
    layer1_outputs(8050) <= a or b;
    layer1_outputs(8051) <= b;
    layer1_outputs(8052) <= a;
    layer1_outputs(8053) <= not (a xor b);
    layer1_outputs(8054) <= not (a and b);
    layer1_outputs(8055) <= not b;
    layer1_outputs(8056) <= a and not b;
    layer1_outputs(8057) <= not (a and b);
    layer1_outputs(8058) <= not a or b;
    layer1_outputs(8059) <= a;
    layer1_outputs(8060) <= a and not b;
    layer1_outputs(8061) <= '0';
    layer1_outputs(8062) <= b and not a;
    layer1_outputs(8063) <= not b or a;
    layer1_outputs(8064) <= a;
    layer1_outputs(8065) <= b;
    layer1_outputs(8066) <= not (a and b);
    layer1_outputs(8067) <= not (a and b);
    layer1_outputs(8068) <= not (a or b);
    layer1_outputs(8069) <= b;
    layer1_outputs(8070) <= a and not b;
    layer1_outputs(8071) <= '1';
    layer1_outputs(8072) <= not a or b;
    layer1_outputs(8073) <= not b;
    layer1_outputs(8074) <= b;
    layer1_outputs(8075) <= a or b;
    layer1_outputs(8076) <= not (a xor b);
    layer1_outputs(8077) <= not b;
    layer1_outputs(8078) <= not (a or b);
    layer1_outputs(8079) <= b and not a;
    layer1_outputs(8080) <= a and b;
    layer1_outputs(8081) <= b and not a;
    layer1_outputs(8082) <= not (a or b);
    layer1_outputs(8083) <= a or b;
    layer1_outputs(8084) <= a or b;
    layer1_outputs(8085) <= a and not b;
    layer1_outputs(8086) <= not a or b;
    layer1_outputs(8087) <= not a;
    layer1_outputs(8088) <= not b;
    layer1_outputs(8089) <= a or b;
    layer1_outputs(8090) <= not b;
    layer1_outputs(8091) <= b;
    layer1_outputs(8092) <= b;
    layer1_outputs(8093) <= b;
    layer1_outputs(8094) <= a or b;
    layer1_outputs(8095) <= a;
    layer1_outputs(8096) <= b;
    layer1_outputs(8097) <= not a or b;
    layer1_outputs(8098) <= not a or b;
    layer1_outputs(8099) <= a xor b;
    layer1_outputs(8100) <= a and b;
    layer1_outputs(8101) <= not (a or b);
    layer1_outputs(8102) <= not a;
    layer1_outputs(8103) <= a and b;
    layer1_outputs(8104) <= a xor b;
    layer1_outputs(8105) <= b;
    layer1_outputs(8106) <= b and not a;
    layer1_outputs(8107) <= a;
    layer1_outputs(8108) <= not a or b;
    layer1_outputs(8109) <= b and not a;
    layer1_outputs(8110) <= b;
    layer1_outputs(8111) <= a and b;
    layer1_outputs(8112) <= not (a xor b);
    layer1_outputs(8113) <= not (a or b);
    layer1_outputs(8114) <= not (a xor b);
    layer1_outputs(8115) <= not (a xor b);
    layer1_outputs(8116) <= a and not b;
    layer1_outputs(8117) <= b and not a;
    layer1_outputs(8118) <= a or b;
    layer1_outputs(8119) <= not b;
    layer1_outputs(8120) <= a and not b;
    layer1_outputs(8121) <= not (a and b);
    layer1_outputs(8122) <= not (a xor b);
    layer1_outputs(8123) <= not b;
    layer1_outputs(8124) <= b;
    layer1_outputs(8125) <= not a or b;
    layer1_outputs(8126) <= not a;
    layer1_outputs(8127) <= not (a or b);
    layer1_outputs(8128) <= not a or b;
    layer1_outputs(8129) <= not b;
    layer1_outputs(8130) <= not b;
    layer1_outputs(8131) <= b;
    layer1_outputs(8132) <= a;
    layer1_outputs(8133) <= not a;
    layer1_outputs(8134) <= not (a or b);
    layer1_outputs(8135) <= a and not b;
    layer1_outputs(8136) <= a;
    layer1_outputs(8137) <= not a;
    layer1_outputs(8138) <= a xor b;
    layer1_outputs(8139) <= not b or a;
    layer1_outputs(8140) <= '1';
    layer1_outputs(8141) <= a xor b;
    layer1_outputs(8142) <= a;
    layer1_outputs(8143) <= a;
    layer1_outputs(8144) <= b and not a;
    layer1_outputs(8145) <= not (a xor b);
    layer1_outputs(8146) <= b;
    layer1_outputs(8147) <= a and b;
    layer1_outputs(8148) <= not a or b;
    layer1_outputs(8149) <= not (a or b);
    layer1_outputs(8150) <= not b;
    layer1_outputs(8151) <= b;
    layer1_outputs(8152) <= a xor b;
    layer1_outputs(8153) <= not b or a;
    layer1_outputs(8154) <= not a;
    layer1_outputs(8155) <= not a or b;
    layer1_outputs(8156) <= not b;
    layer1_outputs(8157) <= '0';
    layer1_outputs(8158) <= not (a and b);
    layer1_outputs(8159) <= not b;
    layer1_outputs(8160) <= not b;
    layer1_outputs(8161) <= a and b;
    layer1_outputs(8162) <= not b;
    layer1_outputs(8163) <= a;
    layer1_outputs(8164) <= a;
    layer1_outputs(8165) <= not b;
    layer1_outputs(8166) <= not (a xor b);
    layer1_outputs(8167) <= a and not b;
    layer1_outputs(8168) <= not b;
    layer1_outputs(8169) <= not a;
    layer1_outputs(8170) <= not b;
    layer1_outputs(8171) <= not (a or b);
    layer1_outputs(8172) <= a;
    layer1_outputs(8173) <= a and b;
    layer1_outputs(8174) <= not a or b;
    layer1_outputs(8175) <= a and not b;
    layer1_outputs(8176) <= a or b;
    layer1_outputs(8177) <= a or b;
    layer1_outputs(8178) <= not a or b;
    layer1_outputs(8179) <= not a or b;
    layer1_outputs(8180) <= not b;
    layer1_outputs(8181) <= a and not b;
    layer1_outputs(8182) <= not a;
    layer1_outputs(8183) <= not a;
    layer1_outputs(8184) <= not a or b;
    layer1_outputs(8185) <= not (a xor b);
    layer1_outputs(8186) <= not b or a;
    layer1_outputs(8187) <= b;
    layer1_outputs(8188) <= not (a and b);
    layer1_outputs(8189) <= b;
    layer1_outputs(8190) <= a and not b;
    layer1_outputs(8191) <= a and not b;
    layer1_outputs(8192) <= a xor b;
    layer1_outputs(8193) <= not a;
    layer1_outputs(8194) <= a;
    layer1_outputs(8195) <= b and not a;
    layer1_outputs(8196) <= b and not a;
    layer1_outputs(8197) <= not a;
    layer1_outputs(8198) <= not a or b;
    layer1_outputs(8199) <= not b or a;
    layer1_outputs(8200) <= not (a or b);
    layer1_outputs(8201) <= a xor b;
    layer1_outputs(8202) <= a and not b;
    layer1_outputs(8203) <= not b or a;
    layer1_outputs(8204) <= not (a or b);
    layer1_outputs(8205) <= not (a and b);
    layer1_outputs(8206) <= b;
    layer1_outputs(8207) <= not (a or b);
    layer1_outputs(8208) <= not (a or b);
    layer1_outputs(8209) <= a;
    layer1_outputs(8210) <= not a or b;
    layer1_outputs(8211) <= '0';
    layer1_outputs(8212) <= a;
    layer1_outputs(8213) <= not a;
    layer1_outputs(8214) <= a;
    layer1_outputs(8215) <= not a or b;
    layer1_outputs(8216) <= a and not b;
    layer1_outputs(8217) <= not b or a;
    layer1_outputs(8218) <= a xor b;
    layer1_outputs(8219) <= a;
    layer1_outputs(8220) <= a;
    layer1_outputs(8221) <= not (a and b);
    layer1_outputs(8222) <= a;
    layer1_outputs(8223) <= not (a xor b);
    layer1_outputs(8224) <= not b or a;
    layer1_outputs(8225) <= not a;
    layer1_outputs(8226) <= not b;
    layer1_outputs(8227) <= b;
    layer1_outputs(8228) <= not a or b;
    layer1_outputs(8229) <= not a or b;
    layer1_outputs(8230) <= '0';
    layer1_outputs(8231) <= a and b;
    layer1_outputs(8232) <= a;
    layer1_outputs(8233) <= not (a or b);
    layer1_outputs(8234) <= not a or b;
    layer1_outputs(8235) <= a;
    layer1_outputs(8236) <= not (a and b);
    layer1_outputs(8237) <= a or b;
    layer1_outputs(8238) <= b;
    layer1_outputs(8239) <= not a;
    layer1_outputs(8240) <= not b or a;
    layer1_outputs(8241) <= a xor b;
    layer1_outputs(8242) <= a or b;
    layer1_outputs(8243) <= b and not a;
    layer1_outputs(8244) <= a xor b;
    layer1_outputs(8245) <= not b or a;
    layer1_outputs(8246) <= not a;
    layer1_outputs(8247) <= not b;
    layer1_outputs(8248) <= a xor b;
    layer1_outputs(8249) <= b;
    layer1_outputs(8250) <= not (a and b);
    layer1_outputs(8251) <= not a or b;
    layer1_outputs(8252) <= a and b;
    layer1_outputs(8253) <= a and not b;
    layer1_outputs(8254) <= a and not b;
    layer1_outputs(8255) <= not b or a;
    layer1_outputs(8256) <= b;
    layer1_outputs(8257) <= not (a or b);
    layer1_outputs(8258) <= b;
    layer1_outputs(8259) <= not (a and b);
    layer1_outputs(8260) <= '0';
    layer1_outputs(8261) <= not a;
    layer1_outputs(8262) <= a xor b;
    layer1_outputs(8263) <= a;
    layer1_outputs(8264) <= not a;
    layer1_outputs(8265) <= a and not b;
    layer1_outputs(8266) <= a;
    layer1_outputs(8267) <= a;
    layer1_outputs(8268) <= b;
    layer1_outputs(8269) <= a and not b;
    layer1_outputs(8270) <= a;
    layer1_outputs(8271) <= not (a or b);
    layer1_outputs(8272) <= a xor b;
    layer1_outputs(8273) <= b;
    layer1_outputs(8274) <= not a or b;
    layer1_outputs(8275) <= a and not b;
    layer1_outputs(8276) <= not b;
    layer1_outputs(8277) <= not (a xor b);
    layer1_outputs(8278) <= b;
    layer1_outputs(8279) <= a;
    layer1_outputs(8280) <= not (a xor b);
    layer1_outputs(8281) <= b and not a;
    layer1_outputs(8282) <= not b;
    layer1_outputs(8283) <= not (a or b);
    layer1_outputs(8284) <= not b;
    layer1_outputs(8285) <= not a or b;
    layer1_outputs(8286) <= not b;
    layer1_outputs(8287) <= a and not b;
    layer1_outputs(8288) <= not (a or b);
    layer1_outputs(8289) <= not b;
    layer1_outputs(8290) <= not a;
    layer1_outputs(8291) <= not b or a;
    layer1_outputs(8292) <= not a;
    layer1_outputs(8293) <= b and not a;
    layer1_outputs(8294) <= not b or a;
    layer1_outputs(8295) <= not b or a;
    layer1_outputs(8296) <= not a;
    layer1_outputs(8297) <= not a or b;
    layer1_outputs(8298) <= not b;
    layer1_outputs(8299) <= a xor b;
    layer1_outputs(8300) <= a;
    layer1_outputs(8301) <= not a or b;
    layer1_outputs(8302) <= a xor b;
    layer1_outputs(8303) <= not a;
    layer1_outputs(8304) <= not a;
    layer1_outputs(8305) <= '1';
    layer1_outputs(8306) <= a or b;
    layer1_outputs(8307) <= a xor b;
    layer1_outputs(8308) <= a;
    layer1_outputs(8309) <= not a or b;
    layer1_outputs(8310) <= b;
    layer1_outputs(8311) <= not b or a;
    layer1_outputs(8312) <= a and not b;
    layer1_outputs(8313) <= not (a and b);
    layer1_outputs(8314) <= not b;
    layer1_outputs(8315) <= not a;
    layer1_outputs(8316) <= not (a or b);
    layer1_outputs(8317) <= not (a or b);
    layer1_outputs(8318) <= not (a or b);
    layer1_outputs(8319) <= not a;
    layer1_outputs(8320) <= not b;
    layer1_outputs(8321) <= not (a xor b);
    layer1_outputs(8322) <= b;
    layer1_outputs(8323) <= not b;
    layer1_outputs(8324) <= a xor b;
    layer1_outputs(8325) <= a;
    layer1_outputs(8326) <= not (a and b);
    layer1_outputs(8327) <= not b or a;
    layer1_outputs(8328) <= not (a and b);
    layer1_outputs(8329) <= not b or a;
    layer1_outputs(8330) <= not (a and b);
    layer1_outputs(8331) <= a xor b;
    layer1_outputs(8332) <= not a;
    layer1_outputs(8333) <= not b;
    layer1_outputs(8334) <= a or b;
    layer1_outputs(8335) <= a and not b;
    layer1_outputs(8336) <= b;
    layer1_outputs(8337) <= a;
    layer1_outputs(8338) <= not (a xor b);
    layer1_outputs(8339) <= not (a xor b);
    layer1_outputs(8340) <= b;
    layer1_outputs(8341) <= a xor b;
    layer1_outputs(8342) <= '1';
    layer1_outputs(8343) <= b;
    layer1_outputs(8344) <= not b or a;
    layer1_outputs(8345) <= a or b;
    layer1_outputs(8346) <= a and not b;
    layer1_outputs(8347) <= a and b;
    layer1_outputs(8348) <= b;
    layer1_outputs(8349) <= not (a or b);
    layer1_outputs(8350) <= not (a and b);
    layer1_outputs(8351) <= b;
    layer1_outputs(8352) <= b;
    layer1_outputs(8353) <= not (a xor b);
    layer1_outputs(8354) <= not (a or b);
    layer1_outputs(8355) <= not b or a;
    layer1_outputs(8356) <= a xor b;
    layer1_outputs(8357) <= not a or b;
    layer1_outputs(8358) <= a or b;
    layer1_outputs(8359) <= not (a xor b);
    layer1_outputs(8360) <= b;
    layer1_outputs(8361) <= a and not b;
    layer1_outputs(8362) <= b and not a;
    layer1_outputs(8363) <= not a or b;
    layer1_outputs(8364) <= not (a xor b);
    layer1_outputs(8365) <= not a;
    layer1_outputs(8366) <= '1';
    layer1_outputs(8367) <= b;
    layer1_outputs(8368) <= not b or a;
    layer1_outputs(8369) <= not (a or b);
    layer1_outputs(8370) <= not (a xor b);
    layer1_outputs(8371) <= not (a and b);
    layer1_outputs(8372) <= not b;
    layer1_outputs(8373) <= not (a or b);
    layer1_outputs(8374) <= a xor b;
    layer1_outputs(8375) <= a xor b;
    layer1_outputs(8376) <= not a;
    layer1_outputs(8377) <= a xor b;
    layer1_outputs(8378) <= not a;
    layer1_outputs(8379) <= not (a or b);
    layer1_outputs(8380) <= not a or b;
    layer1_outputs(8381) <= not a or b;
    layer1_outputs(8382) <= not b;
    layer1_outputs(8383) <= not (a xor b);
    layer1_outputs(8384) <= a xor b;
    layer1_outputs(8385) <= b;
    layer1_outputs(8386) <= not (a or b);
    layer1_outputs(8387) <= not b;
    layer1_outputs(8388) <= not (a and b);
    layer1_outputs(8389) <= a;
    layer1_outputs(8390) <= not b or a;
    layer1_outputs(8391) <= not a;
    layer1_outputs(8392) <= not a;
    layer1_outputs(8393) <= '1';
    layer1_outputs(8394) <= b;
    layer1_outputs(8395) <= not (a or b);
    layer1_outputs(8396) <= not b;
    layer1_outputs(8397) <= not (a xor b);
    layer1_outputs(8398) <= a and b;
    layer1_outputs(8399) <= not b;
    layer1_outputs(8400) <= b and not a;
    layer1_outputs(8401) <= a;
    layer1_outputs(8402) <= not (a or b);
    layer1_outputs(8403) <= a xor b;
    layer1_outputs(8404) <= not b or a;
    layer1_outputs(8405) <= a and not b;
    layer1_outputs(8406) <= a xor b;
    layer1_outputs(8407) <= not a;
    layer1_outputs(8408) <= b;
    layer1_outputs(8409) <= not (a or b);
    layer1_outputs(8410) <= a and not b;
    layer1_outputs(8411) <= b and not a;
    layer1_outputs(8412) <= not (a xor b);
    layer1_outputs(8413) <= a and b;
    layer1_outputs(8414) <= a or b;
    layer1_outputs(8415) <= not a or b;
    layer1_outputs(8416) <= not b;
    layer1_outputs(8417) <= not (a xor b);
    layer1_outputs(8418) <= a or b;
    layer1_outputs(8419) <= not b or a;
    layer1_outputs(8420) <= not (a and b);
    layer1_outputs(8421) <= not b;
    layer1_outputs(8422) <= a;
    layer1_outputs(8423) <= a and not b;
    layer1_outputs(8424) <= not b or a;
    layer1_outputs(8425) <= not a or b;
    layer1_outputs(8426) <= not (a and b);
    layer1_outputs(8427) <= a and b;
    layer1_outputs(8428) <= not b;
    layer1_outputs(8429) <= a;
    layer1_outputs(8430) <= not b;
    layer1_outputs(8431) <= a xor b;
    layer1_outputs(8432) <= a;
    layer1_outputs(8433) <= not b;
    layer1_outputs(8434) <= not a;
    layer1_outputs(8435) <= a;
    layer1_outputs(8436) <= not b;
    layer1_outputs(8437) <= not (a xor b);
    layer1_outputs(8438) <= a and not b;
    layer1_outputs(8439) <= b;
    layer1_outputs(8440) <= not (a and b);
    layer1_outputs(8441) <= not (a and b);
    layer1_outputs(8442) <= a and b;
    layer1_outputs(8443) <= not a;
    layer1_outputs(8444) <= a and b;
    layer1_outputs(8445) <= b;
    layer1_outputs(8446) <= not b;
    layer1_outputs(8447) <= a or b;
    layer1_outputs(8448) <= not b;
    layer1_outputs(8449) <= a and not b;
    layer1_outputs(8450) <= a and not b;
    layer1_outputs(8451) <= not b;
    layer1_outputs(8452) <= not (a and b);
    layer1_outputs(8453) <= not b;
    layer1_outputs(8454) <= not a;
    layer1_outputs(8455) <= not a or b;
    layer1_outputs(8456) <= not (a or b);
    layer1_outputs(8457) <= a and not b;
    layer1_outputs(8458) <= a xor b;
    layer1_outputs(8459) <= not a or b;
    layer1_outputs(8460) <= not (a xor b);
    layer1_outputs(8461) <= a and not b;
    layer1_outputs(8462) <= a xor b;
    layer1_outputs(8463) <= not b or a;
    layer1_outputs(8464) <= not b;
    layer1_outputs(8465) <= a or b;
    layer1_outputs(8466) <= a xor b;
    layer1_outputs(8467) <= not a;
    layer1_outputs(8468) <= b and not a;
    layer1_outputs(8469) <= b and not a;
    layer1_outputs(8470) <= a or b;
    layer1_outputs(8471) <= a and not b;
    layer1_outputs(8472) <= a and b;
    layer1_outputs(8473) <= b;
    layer1_outputs(8474) <= b and not a;
    layer1_outputs(8475) <= not a or b;
    layer1_outputs(8476) <= not a or b;
    layer1_outputs(8477) <= a or b;
    layer1_outputs(8478) <= not (a xor b);
    layer1_outputs(8479) <= b;
    layer1_outputs(8480) <= not (a and b);
    layer1_outputs(8481) <= a and b;
    layer1_outputs(8482) <= b and not a;
    layer1_outputs(8483) <= not b or a;
    layer1_outputs(8484) <= b and not a;
    layer1_outputs(8485) <= not a;
    layer1_outputs(8486) <= a and b;
    layer1_outputs(8487) <= a xor b;
    layer1_outputs(8488) <= a and b;
    layer1_outputs(8489) <= not b;
    layer1_outputs(8490) <= b and not a;
    layer1_outputs(8491) <= b and not a;
    layer1_outputs(8492) <= a xor b;
    layer1_outputs(8493) <= a and not b;
    layer1_outputs(8494) <= a or b;
    layer1_outputs(8495) <= not (a or b);
    layer1_outputs(8496) <= a;
    layer1_outputs(8497) <= not b;
    layer1_outputs(8498) <= a;
    layer1_outputs(8499) <= a or b;
    layer1_outputs(8500) <= not (a and b);
    layer1_outputs(8501) <= not a or b;
    layer1_outputs(8502) <= not b;
    layer1_outputs(8503) <= not a or b;
    layer1_outputs(8504) <= not a;
    layer1_outputs(8505) <= a;
    layer1_outputs(8506) <= a;
    layer1_outputs(8507) <= not a;
    layer1_outputs(8508) <= a xor b;
    layer1_outputs(8509) <= not a or b;
    layer1_outputs(8510) <= b;
    layer1_outputs(8511) <= not (a xor b);
    layer1_outputs(8512) <= not (a xor b);
    layer1_outputs(8513) <= a xor b;
    layer1_outputs(8514) <= not b;
    layer1_outputs(8515) <= not (a and b);
    layer1_outputs(8516) <= not a or b;
    layer1_outputs(8517) <= a or b;
    layer1_outputs(8518) <= a;
    layer1_outputs(8519) <= not (a or b);
    layer1_outputs(8520) <= not a;
    layer1_outputs(8521) <= b and not a;
    layer1_outputs(8522) <= not (a xor b);
    layer1_outputs(8523) <= a;
    layer1_outputs(8524) <= not b;
    layer1_outputs(8525) <= b and not a;
    layer1_outputs(8526) <= not (a xor b);
    layer1_outputs(8527) <= a;
    layer1_outputs(8528) <= a and b;
    layer1_outputs(8529) <= not (a and b);
    layer1_outputs(8530) <= a;
    layer1_outputs(8531) <= a or b;
    layer1_outputs(8532) <= not (a or b);
    layer1_outputs(8533) <= a;
    layer1_outputs(8534) <= not b;
    layer1_outputs(8535) <= not b;
    layer1_outputs(8536) <= b and not a;
    layer1_outputs(8537) <= not b;
    layer1_outputs(8538) <= not (a and b);
    layer1_outputs(8539) <= not a;
    layer1_outputs(8540) <= '1';
    layer1_outputs(8541) <= a or b;
    layer1_outputs(8542) <= b;
    layer1_outputs(8543) <= a and b;
    layer1_outputs(8544) <= not a or b;
    layer1_outputs(8545) <= not (a or b);
    layer1_outputs(8546) <= not (a xor b);
    layer1_outputs(8547) <= not (a and b);
    layer1_outputs(8548) <= not b;
    layer1_outputs(8549) <= '0';
    layer1_outputs(8550) <= a xor b;
    layer1_outputs(8551) <= not (a xor b);
    layer1_outputs(8552) <= not b;
    layer1_outputs(8553) <= not (a xor b);
    layer1_outputs(8554) <= not a;
    layer1_outputs(8555) <= not b or a;
    layer1_outputs(8556) <= not (a and b);
    layer1_outputs(8557) <= a and not b;
    layer1_outputs(8558) <= b and not a;
    layer1_outputs(8559) <= b;
    layer1_outputs(8560) <= not b;
    layer1_outputs(8561) <= a xor b;
    layer1_outputs(8562) <= not a;
    layer1_outputs(8563) <= a or b;
    layer1_outputs(8564) <= not (a and b);
    layer1_outputs(8565) <= a;
    layer1_outputs(8566) <= '0';
    layer1_outputs(8567) <= b;
    layer1_outputs(8568) <= not a;
    layer1_outputs(8569) <= b and not a;
    layer1_outputs(8570) <= not (a and b);
    layer1_outputs(8571) <= not b;
    layer1_outputs(8572) <= a and not b;
    layer1_outputs(8573) <= b;
    layer1_outputs(8574) <= not (a xor b);
    layer1_outputs(8575) <= '1';
    layer1_outputs(8576) <= not a;
    layer1_outputs(8577) <= a xor b;
    layer1_outputs(8578) <= not (a or b);
    layer1_outputs(8579) <= not (a or b);
    layer1_outputs(8580) <= a xor b;
    layer1_outputs(8581) <= a and b;
    layer1_outputs(8582) <= a;
    layer1_outputs(8583) <= not b or a;
    layer1_outputs(8584) <= a and not b;
    layer1_outputs(8585) <= not b;
    layer1_outputs(8586) <= a xor b;
    layer1_outputs(8587) <= not (a and b);
    layer1_outputs(8588) <= a;
    layer1_outputs(8589) <= b and not a;
    layer1_outputs(8590) <= '1';
    layer1_outputs(8591) <= b;
    layer1_outputs(8592) <= a xor b;
    layer1_outputs(8593) <= a xor b;
    layer1_outputs(8594) <= a;
    layer1_outputs(8595) <= a xor b;
    layer1_outputs(8596) <= not b or a;
    layer1_outputs(8597) <= a xor b;
    layer1_outputs(8598) <= b;
    layer1_outputs(8599) <= not a;
    layer1_outputs(8600) <= not a;
    layer1_outputs(8601) <= not b or a;
    layer1_outputs(8602) <= not b;
    layer1_outputs(8603) <= b and not a;
    layer1_outputs(8604) <= not b or a;
    layer1_outputs(8605) <= a and b;
    layer1_outputs(8606) <= not (a xor b);
    layer1_outputs(8607) <= a and b;
    layer1_outputs(8608) <= a or b;
    layer1_outputs(8609) <= not b;
    layer1_outputs(8610) <= a;
    layer1_outputs(8611) <= not (a and b);
    layer1_outputs(8612) <= not (a or b);
    layer1_outputs(8613) <= not a or b;
    layer1_outputs(8614) <= a or b;
    layer1_outputs(8615) <= b;
    layer1_outputs(8616) <= a xor b;
    layer1_outputs(8617) <= not b;
    layer1_outputs(8618) <= a and b;
    layer1_outputs(8619) <= b and not a;
    layer1_outputs(8620) <= not b;
    layer1_outputs(8621) <= a;
    layer1_outputs(8622) <= not b or a;
    layer1_outputs(8623) <= not (a and b);
    layer1_outputs(8624) <= a;
    layer1_outputs(8625) <= not b;
    layer1_outputs(8626) <= not a or b;
    layer1_outputs(8627) <= not b;
    layer1_outputs(8628) <= a;
    layer1_outputs(8629) <= not (a xor b);
    layer1_outputs(8630) <= a xor b;
    layer1_outputs(8631) <= not a or b;
    layer1_outputs(8632) <= not b;
    layer1_outputs(8633) <= not a;
    layer1_outputs(8634) <= not (a and b);
    layer1_outputs(8635) <= a or b;
    layer1_outputs(8636) <= a and b;
    layer1_outputs(8637) <= not (a and b);
    layer1_outputs(8638) <= b;
    layer1_outputs(8639) <= a;
    layer1_outputs(8640) <= not (a xor b);
    layer1_outputs(8641) <= not b;
    layer1_outputs(8642) <= not a;
    layer1_outputs(8643) <= a and not b;
    layer1_outputs(8644) <= not a;
    layer1_outputs(8645) <= b and not a;
    layer1_outputs(8646) <= not (a xor b);
    layer1_outputs(8647) <= a or b;
    layer1_outputs(8648) <= b and not a;
    layer1_outputs(8649) <= not (a xor b);
    layer1_outputs(8650) <= a and not b;
    layer1_outputs(8651) <= not (a and b);
    layer1_outputs(8652) <= not a;
    layer1_outputs(8653) <= not b;
    layer1_outputs(8654) <= b;
    layer1_outputs(8655) <= a and b;
    layer1_outputs(8656) <= not b or a;
    layer1_outputs(8657) <= b;
    layer1_outputs(8658) <= not (a xor b);
    layer1_outputs(8659) <= a;
    layer1_outputs(8660) <= b;
    layer1_outputs(8661) <= not b or a;
    layer1_outputs(8662) <= not (a xor b);
    layer1_outputs(8663) <= not a;
    layer1_outputs(8664) <= a and not b;
    layer1_outputs(8665) <= not (a xor b);
    layer1_outputs(8666) <= a and b;
    layer1_outputs(8667) <= not (a and b);
    layer1_outputs(8668) <= not b;
    layer1_outputs(8669) <= not (a or b);
    layer1_outputs(8670) <= b;
    layer1_outputs(8671) <= not b;
    layer1_outputs(8672) <= a and not b;
    layer1_outputs(8673) <= not b;
    layer1_outputs(8674) <= not b;
    layer1_outputs(8675) <= not a;
    layer1_outputs(8676) <= a;
    layer1_outputs(8677) <= not a;
    layer1_outputs(8678) <= not (a xor b);
    layer1_outputs(8679) <= a and not b;
    layer1_outputs(8680) <= '0';
    layer1_outputs(8681) <= not b;
    layer1_outputs(8682) <= a xor b;
    layer1_outputs(8683) <= '0';
    layer1_outputs(8684) <= a and b;
    layer1_outputs(8685) <= not b;
    layer1_outputs(8686) <= not (a or b);
    layer1_outputs(8687) <= not a;
    layer1_outputs(8688) <= a and b;
    layer1_outputs(8689) <= not a;
    layer1_outputs(8690) <= b and not a;
    layer1_outputs(8691) <= b and not a;
    layer1_outputs(8692) <= not b or a;
    layer1_outputs(8693) <= not (a or b);
    layer1_outputs(8694) <= not (a and b);
    layer1_outputs(8695) <= a;
    layer1_outputs(8696) <= b and not a;
    layer1_outputs(8697) <= b and not a;
    layer1_outputs(8698) <= not (a xor b);
    layer1_outputs(8699) <= not b;
    layer1_outputs(8700) <= not b;
    layer1_outputs(8701) <= a;
    layer1_outputs(8702) <= not b;
    layer1_outputs(8703) <= not a;
    layer1_outputs(8704) <= a or b;
    layer1_outputs(8705) <= not (a and b);
    layer1_outputs(8706) <= not a;
    layer1_outputs(8707) <= not b or a;
    layer1_outputs(8708) <= a;
    layer1_outputs(8709) <= a;
    layer1_outputs(8710) <= not b or a;
    layer1_outputs(8711) <= b and not a;
    layer1_outputs(8712) <= b and not a;
    layer1_outputs(8713) <= not (a and b);
    layer1_outputs(8714) <= not b;
    layer1_outputs(8715) <= a xor b;
    layer1_outputs(8716) <= not a;
    layer1_outputs(8717) <= a or b;
    layer1_outputs(8718) <= a or b;
    layer1_outputs(8719) <= a;
    layer1_outputs(8720) <= not a;
    layer1_outputs(8721) <= a and b;
    layer1_outputs(8722) <= a xor b;
    layer1_outputs(8723) <= not a;
    layer1_outputs(8724) <= not (a xor b);
    layer1_outputs(8725) <= b and not a;
    layer1_outputs(8726) <= not a or b;
    layer1_outputs(8727) <= not (a xor b);
    layer1_outputs(8728) <= not (a or b);
    layer1_outputs(8729) <= a;
    layer1_outputs(8730) <= a xor b;
    layer1_outputs(8731) <= a and not b;
    layer1_outputs(8732) <= a and b;
    layer1_outputs(8733) <= not b or a;
    layer1_outputs(8734) <= not (a or b);
    layer1_outputs(8735) <= b and not a;
    layer1_outputs(8736) <= a and not b;
    layer1_outputs(8737) <= a or b;
    layer1_outputs(8738) <= not b;
    layer1_outputs(8739) <= not b;
    layer1_outputs(8740) <= not (a xor b);
    layer1_outputs(8741) <= b and not a;
    layer1_outputs(8742) <= '0';
    layer1_outputs(8743) <= a xor b;
    layer1_outputs(8744) <= not b or a;
    layer1_outputs(8745) <= a or b;
    layer1_outputs(8746) <= not (a and b);
    layer1_outputs(8747) <= a xor b;
    layer1_outputs(8748) <= '0';
    layer1_outputs(8749) <= a;
    layer1_outputs(8750) <= a or b;
    layer1_outputs(8751) <= b;
    layer1_outputs(8752) <= a;
    layer1_outputs(8753) <= not (a xor b);
    layer1_outputs(8754) <= a;
    layer1_outputs(8755) <= a and b;
    layer1_outputs(8756) <= b and not a;
    layer1_outputs(8757) <= not (a and b);
    layer1_outputs(8758) <= a and not b;
    layer1_outputs(8759) <= not a;
    layer1_outputs(8760) <= a xor b;
    layer1_outputs(8761) <= not b or a;
    layer1_outputs(8762) <= not (a and b);
    layer1_outputs(8763) <= not a;
    layer1_outputs(8764) <= a xor b;
    layer1_outputs(8765) <= not (a and b);
    layer1_outputs(8766) <= not (a and b);
    layer1_outputs(8767) <= b;
    layer1_outputs(8768) <= a;
    layer1_outputs(8769) <= not a;
    layer1_outputs(8770) <= not a;
    layer1_outputs(8771) <= a and not b;
    layer1_outputs(8772) <= b and not a;
    layer1_outputs(8773) <= not b;
    layer1_outputs(8774) <= not a or b;
    layer1_outputs(8775) <= not b;
    layer1_outputs(8776) <= a and not b;
    layer1_outputs(8777) <= a and not b;
    layer1_outputs(8778) <= a xor b;
    layer1_outputs(8779) <= a;
    layer1_outputs(8780) <= a and b;
    layer1_outputs(8781) <= not (a and b);
    layer1_outputs(8782) <= b and not a;
    layer1_outputs(8783) <= not a;
    layer1_outputs(8784) <= b;
    layer1_outputs(8785) <= b;
    layer1_outputs(8786) <= not a;
    layer1_outputs(8787) <= not (a or b);
    layer1_outputs(8788) <= a xor b;
    layer1_outputs(8789) <= not b or a;
    layer1_outputs(8790) <= not b or a;
    layer1_outputs(8791) <= a xor b;
    layer1_outputs(8792) <= a and b;
    layer1_outputs(8793) <= not a or b;
    layer1_outputs(8794) <= not a or b;
    layer1_outputs(8795) <= not (a and b);
    layer1_outputs(8796) <= '0';
    layer1_outputs(8797) <= a or b;
    layer1_outputs(8798) <= not a;
    layer1_outputs(8799) <= a and b;
    layer1_outputs(8800) <= not a;
    layer1_outputs(8801) <= a or b;
    layer1_outputs(8802) <= not b;
    layer1_outputs(8803) <= not a;
    layer1_outputs(8804) <= not a;
    layer1_outputs(8805) <= not (a or b);
    layer1_outputs(8806) <= not (a and b);
    layer1_outputs(8807) <= a xor b;
    layer1_outputs(8808) <= a or b;
    layer1_outputs(8809) <= a and not b;
    layer1_outputs(8810) <= b and not a;
    layer1_outputs(8811) <= b and not a;
    layer1_outputs(8812) <= not b or a;
    layer1_outputs(8813) <= a and b;
    layer1_outputs(8814) <= a;
    layer1_outputs(8815) <= a and b;
    layer1_outputs(8816) <= a xor b;
    layer1_outputs(8817) <= not b or a;
    layer1_outputs(8818) <= not (a xor b);
    layer1_outputs(8819) <= not b or a;
    layer1_outputs(8820) <= not (a xor b);
    layer1_outputs(8821) <= not b or a;
    layer1_outputs(8822) <= not b;
    layer1_outputs(8823) <= a xor b;
    layer1_outputs(8824) <= '0';
    layer1_outputs(8825) <= b;
    layer1_outputs(8826) <= a xor b;
    layer1_outputs(8827) <= a or b;
    layer1_outputs(8828) <= a;
    layer1_outputs(8829) <= not (a or b);
    layer1_outputs(8830) <= not a or b;
    layer1_outputs(8831) <= not (a xor b);
    layer1_outputs(8832) <= not (a and b);
    layer1_outputs(8833) <= a and not b;
    layer1_outputs(8834) <= b and not a;
    layer1_outputs(8835) <= a;
    layer1_outputs(8836) <= not a;
    layer1_outputs(8837) <= b;
    layer1_outputs(8838) <= not (a and b);
    layer1_outputs(8839) <= not a;
    layer1_outputs(8840) <= not (a or b);
    layer1_outputs(8841) <= a;
    layer1_outputs(8842) <= a and b;
    layer1_outputs(8843) <= not (a and b);
    layer1_outputs(8844) <= a and b;
    layer1_outputs(8845) <= not (a and b);
    layer1_outputs(8846) <= not b or a;
    layer1_outputs(8847) <= b and not a;
    layer1_outputs(8848) <= b and not a;
    layer1_outputs(8849) <= a and b;
    layer1_outputs(8850) <= not b or a;
    layer1_outputs(8851) <= a and b;
    layer1_outputs(8852) <= a and not b;
    layer1_outputs(8853) <= a or b;
    layer1_outputs(8854) <= not a;
    layer1_outputs(8855) <= not b;
    layer1_outputs(8856) <= a or b;
    layer1_outputs(8857) <= not b or a;
    layer1_outputs(8858) <= a;
    layer1_outputs(8859) <= a and b;
    layer1_outputs(8860) <= b;
    layer1_outputs(8861) <= not (a xor b);
    layer1_outputs(8862) <= a;
    layer1_outputs(8863) <= not a;
    layer1_outputs(8864) <= b;
    layer1_outputs(8865) <= not (a xor b);
    layer1_outputs(8866) <= not b;
    layer1_outputs(8867) <= not (a or b);
    layer1_outputs(8868) <= a;
    layer1_outputs(8869) <= not a;
    layer1_outputs(8870) <= not b;
    layer1_outputs(8871) <= not b or a;
    layer1_outputs(8872) <= not b;
    layer1_outputs(8873) <= a or b;
    layer1_outputs(8874) <= not b;
    layer1_outputs(8875) <= b;
    layer1_outputs(8876) <= a;
    layer1_outputs(8877) <= not (a and b);
    layer1_outputs(8878) <= not b or a;
    layer1_outputs(8879) <= not b;
    layer1_outputs(8880) <= a and not b;
    layer1_outputs(8881) <= not (a and b);
    layer1_outputs(8882) <= not b;
    layer1_outputs(8883) <= a or b;
    layer1_outputs(8884) <= b;
    layer1_outputs(8885) <= '0';
    layer1_outputs(8886) <= b;
    layer1_outputs(8887) <= not b;
    layer1_outputs(8888) <= a and not b;
    layer1_outputs(8889) <= a or b;
    layer1_outputs(8890) <= not a;
    layer1_outputs(8891) <= not a;
    layer1_outputs(8892) <= not b or a;
    layer1_outputs(8893) <= a;
    layer1_outputs(8894) <= not (a or b);
    layer1_outputs(8895) <= b;
    layer1_outputs(8896) <= not (a xor b);
    layer1_outputs(8897) <= a and b;
    layer1_outputs(8898) <= not b or a;
    layer1_outputs(8899) <= a and not b;
    layer1_outputs(8900) <= not a;
    layer1_outputs(8901) <= b;
    layer1_outputs(8902) <= not a;
    layer1_outputs(8903) <= a and b;
    layer1_outputs(8904) <= not b;
    layer1_outputs(8905) <= b and not a;
    layer1_outputs(8906) <= not b;
    layer1_outputs(8907) <= not b;
    layer1_outputs(8908) <= not a or b;
    layer1_outputs(8909) <= b;
    layer1_outputs(8910) <= not b;
    layer1_outputs(8911) <= not (a and b);
    layer1_outputs(8912) <= not (a and b);
    layer1_outputs(8913) <= a;
    layer1_outputs(8914) <= not a or b;
    layer1_outputs(8915) <= a and not b;
    layer1_outputs(8916) <= not (a or b);
    layer1_outputs(8917) <= a and b;
    layer1_outputs(8918) <= b;
    layer1_outputs(8919) <= not a or b;
    layer1_outputs(8920) <= not b or a;
    layer1_outputs(8921) <= b and not a;
    layer1_outputs(8922) <= a or b;
    layer1_outputs(8923) <= b and not a;
    layer1_outputs(8924) <= not b;
    layer1_outputs(8925) <= a and not b;
    layer1_outputs(8926) <= a and b;
    layer1_outputs(8927) <= a;
    layer1_outputs(8928) <= b;
    layer1_outputs(8929) <= not b;
    layer1_outputs(8930) <= b;
    layer1_outputs(8931) <= a;
    layer1_outputs(8932) <= not (a xor b);
    layer1_outputs(8933) <= a and not b;
    layer1_outputs(8934) <= b;
    layer1_outputs(8935) <= b;
    layer1_outputs(8936) <= not a or b;
    layer1_outputs(8937) <= not (a and b);
    layer1_outputs(8938) <= b and not a;
    layer1_outputs(8939) <= not (a xor b);
    layer1_outputs(8940) <= a and not b;
    layer1_outputs(8941) <= b and not a;
    layer1_outputs(8942) <= a or b;
    layer1_outputs(8943) <= a or b;
    layer1_outputs(8944) <= not (a and b);
    layer1_outputs(8945) <= a or b;
    layer1_outputs(8946) <= a xor b;
    layer1_outputs(8947) <= not (a xor b);
    layer1_outputs(8948) <= a xor b;
    layer1_outputs(8949) <= not a;
    layer1_outputs(8950) <= a or b;
    layer1_outputs(8951) <= a xor b;
    layer1_outputs(8952) <= not (a or b);
    layer1_outputs(8953) <= a;
    layer1_outputs(8954) <= not b;
    layer1_outputs(8955) <= not (a xor b);
    layer1_outputs(8956) <= not (a and b);
    layer1_outputs(8957) <= not (a xor b);
    layer1_outputs(8958) <= not (a and b);
    layer1_outputs(8959) <= b and not a;
    layer1_outputs(8960) <= not a;
    layer1_outputs(8961) <= not a or b;
    layer1_outputs(8962) <= a and not b;
    layer1_outputs(8963) <= a or b;
    layer1_outputs(8964) <= b and not a;
    layer1_outputs(8965) <= '0';
    layer1_outputs(8966) <= not (a or b);
    layer1_outputs(8967) <= a;
    layer1_outputs(8968) <= a;
    layer1_outputs(8969) <= not (a or b);
    layer1_outputs(8970) <= not a or b;
    layer1_outputs(8971) <= b;
    layer1_outputs(8972) <= a and not b;
    layer1_outputs(8973) <= not a or b;
    layer1_outputs(8974) <= '1';
    layer1_outputs(8975) <= a and b;
    layer1_outputs(8976) <= not b;
    layer1_outputs(8977) <= not a or b;
    layer1_outputs(8978) <= not b or a;
    layer1_outputs(8979) <= not b;
    layer1_outputs(8980) <= b;
    layer1_outputs(8981) <= '1';
    layer1_outputs(8982) <= a or b;
    layer1_outputs(8983) <= a and b;
    layer1_outputs(8984) <= b;
    layer1_outputs(8985) <= not a or b;
    layer1_outputs(8986) <= not b;
    layer1_outputs(8987) <= a and not b;
    layer1_outputs(8988) <= not (a and b);
    layer1_outputs(8989) <= not a or b;
    layer1_outputs(8990) <= a or b;
    layer1_outputs(8991) <= not b;
    layer1_outputs(8992) <= a or b;
    layer1_outputs(8993) <= b;
    layer1_outputs(8994) <= not a;
    layer1_outputs(8995) <= not b;
    layer1_outputs(8996) <= a;
    layer1_outputs(8997) <= b;
    layer1_outputs(8998) <= b and not a;
    layer1_outputs(8999) <= b;
    layer1_outputs(9000) <= not a;
    layer1_outputs(9001) <= b;
    layer1_outputs(9002) <= not (a xor b);
    layer1_outputs(9003) <= not b;
    layer1_outputs(9004) <= not (a xor b);
    layer1_outputs(9005) <= not b or a;
    layer1_outputs(9006) <= b;
    layer1_outputs(9007) <= not (a or b);
    layer1_outputs(9008) <= not (a and b);
    layer1_outputs(9009) <= b and not a;
    layer1_outputs(9010) <= '0';
    layer1_outputs(9011) <= a or b;
    layer1_outputs(9012) <= not a;
    layer1_outputs(9013) <= not b or a;
    layer1_outputs(9014) <= not a;
    layer1_outputs(9015) <= a;
    layer1_outputs(9016) <= a;
    layer1_outputs(9017) <= not (a or b);
    layer1_outputs(9018) <= a and b;
    layer1_outputs(9019) <= a;
    layer1_outputs(9020) <= not (a and b);
    layer1_outputs(9021) <= not (a xor b);
    layer1_outputs(9022) <= not a;
    layer1_outputs(9023) <= a or b;
    layer1_outputs(9024) <= not (a and b);
    layer1_outputs(9025) <= not a or b;
    layer1_outputs(9026) <= a or b;
    layer1_outputs(9027) <= a xor b;
    layer1_outputs(9028) <= not a;
    layer1_outputs(9029) <= not b or a;
    layer1_outputs(9030) <= a xor b;
    layer1_outputs(9031) <= b and not a;
    layer1_outputs(9032) <= a;
    layer1_outputs(9033) <= not (a and b);
    layer1_outputs(9034) <= b and not a;
    layer1_outputs(9035) <= not (a or b);
    layer1_outputs(9036) <= b;
    layer1_outputs(9037) <= not b;
    layer1_outputs(9038) <= not (a and b);
    layer1_outputs(9039) <= not b;
    layer1_outputs(9040) <= not b;
    layer1_outputs(9041) <= b;
    layer1_outputs(9042) <= not b;
    layer1_outputs(9043) <= not b;
    layer1_outputs(9044) <= not a;
    layer1_outputs(9045) <= not a or b;
    layer1_outputs(9046) <= b and not a;
    layer1_outputs(9047) <= a xor b;
    layer1_outputs(9048) <= not b;
    layer1_outputs(9049) <= a and not b;
    layer1_outputs(9050) <= b;
    layer1_outputs(9051) <= a;
    layer1_outputs(9052) <= not (a and b);
    layer1_outputs(9053) <= a;
    layer1_outputs(9054) <= not (a and b);
    layer1_outputs(9055) <= b and not a;
    layer1_outputs(9056) <= not a;
    layer1_outputs(9057) <= a and b;
    layer1_outputs(9058) <= not a;
    layer1_outputs(9059) <= a xor b;
    layer1_outputs(9060) <= a and b;
    layer1_outputs(9061) <= not b;
    layer1_outputs(9062) <= a xor b;
    layer1_outputs(9063) <= not (a xor b);
    layer1_outputs(9064) <= a xor b;
    layer1_outputs(9065) <= a and not b;
    layer1_outputs(9066) <= not (a or b);
    layer1_outputs(9067) <= a or b;
    layer1_outputs(9068) <= a and not b;
    layer1_outputs(9069) <= not b;
    layer1_outputs(9070) <= a xor b;
    layer1_outputs(9071) <= a xor b;
    layer1_outputs(9072) <= a or b;
    layer1_outputs(9073) <= a and b;
    layer1_outputs(9074) <= not (a xor b);
    layer1_outputs(9075) <= not (a or b);
    layer1_outputs(9076) <= b and not a;
    layer1_outputs(9077) <= not b or a;
    layer1_outputs(9078) <= a and b;
    layer1_outputs(9079) <= not (a and b);
    layer1_outputs(9080) <= a xor b;
    layer1_outputs(9081) <= b and not a;
    layer1_outputs(9082) <= not a;
    layer1_outputs(9083) <= not b or a;
    layer1_outputs(9084) <= b;
    layer1_outputs(9085) <= not a or b;
    layer1_outputs(9086) <= not (a xor b);
    layer1_outputs(9087) <= a xor b;
    layer1_outputs(9088) <= b and not a;
    layer1_outputs(9089) <= b and not a;
    layer1_outputs(9090) <= not (a or b);
    layer1_outputs(9091) <= b and not a;
    layer1_outputs(9092) <= not b or a;
    layer1_outputs(9093) <= not b or a;
    layer1_outputs(9094) <= '1';
    layer1_outputs(9095) <= not (a xor b);
    layer1_outputs(9096) <= b and not a;
    layer1_outputs(9097) <= not b;
    layer1_outputs(9098) <= not (a and b);
    layer1_outputs(9099) <= b;
    layer1_outputs(9100) <= '0';
    layer1_outputs(9101) <= not b or a;
    layer1_outputs(9102) <= not b;
    layer1_outputs(9103) <= a;
    layer1_outputs(9104) <= not b or a;
    layer1_outputs(9105) <= a;
    layer1_outputs(9106) <= b;
    layer1_outputs(9107) <= not b;
    layer1_outputs(9108) <= not b;
    layer1_outputs(9109) <= not b;
    layer1_outputs(9110) <= not (a and b);
    layer1_outputs(9111) <= not (a xor b);
    layer1_outputs(9112) <= not a;
    layer1_outputs(9113) <= '0';
    layer1_outputs(9114) <= not b or a;
    layer1_outputs(9115) <= not a;
    layer1_outputs(9116) <= not (a xor b);
    layer1_outputs(9117) <= not b;
    layer1_outputs(9118) <= a xor b;
    layer1_outputs(9119) <= not b or a;
    layer1_outputs(9120) <= not (a xor b);
    layer1_outputs(9121) <= a and b;
    layer1_outputs(9122) <= not b;
    layer1_outputs(9123) <= b and not a;
    layer1_outputs(9124) <= not (a xor b);
    layer1_outputs(9125) <= b;
    layer1_outputs(9126) <= a and b;
    layer1_outputs(9127) <= b;
    layer1_outputs(9128) <= not b;
    layer1_outputs(9129) <= b;
    layer1_outputs(9130) <= a or b;
    layer1_outputs(9131) <= not a or b;
    layer1_outputs(9132) <= not a;
    layer1_outputs(9133) <= not (a and b);
    layer1_outputs(9134) <= a;
    layer1_outputs(9135) <= a and not b;
    layer1_outputs(9136) <= not (a xor b);
    layer1_outputs(9137) <= not a or b;
    layer1_outputs(9138) <= a and not b;
    layer1_outputs(9139) <= a or b;
    layer1_outputs(9140) <= not (a and b);
    layer1_outputs(9141) <= not b or a;
    layer1_outputs(9142) <= not a or b;
    layer1_outputs(9143) <= not a;
    layer1_outputs(9144) <= a and not b;
    layer1_outputs(9145) <= b;
    layer1_outputs(9146) <= b and not a;
    layer1_outputs(9147) <= b;
    layer1_outputs(9148) <= not a;
    layer1_outputs(9149) <= not b;
    layer1_outputs(9150) <= a and not b;
    layer1_outputs(9151) <= not (a xor b);
    layer1_outputs(9152) <= a and not b;
    layer1_outputs(9153) <= not (a or b);
    layer1_outputs(9154) <= b;
    layer1_outputs(9155) <= a xor b;
    layer1_outputs(9156) <= b;
    layer1_outputs(9157) <= a or b;
    layer1_outputs(9158) <= not b;
    layer1_outputs(9159) <= not a;
    layer1_outputs(9160) <= not a or b;
    layer1_outputs(9161) <= not (a and b);
    layer1_outputs(9162) <= not (a or b);
    layer1_outputs(9163) <= a;
    layer1_outputs(9164) <= a and b;
    layer1_outputs(9165) <= not b;
    layer1_outputs(9166) <= not a;
    layer1_outputs(9167) <= a or b;
    layer1_outputs(9168) <= a or b;
    layer1_outputs(9169) <= a xor b;
    layer1_outputs(9170) <= not (a xor b);
    layer1_outputs(9171) <= not (a or b);
    layer1_outputs(9172) <= b;
    layer1_outputs(9173) <= not (a and b);
    layer1_outputs(9174) <= not (a xor b);
    layer1_outputs(9175) <= not b;
    layer1_outputs(9176) <= a xor b;
    layer1_outputs(9177) <= a xor b;
    layer1_outputs(9178) <= not a or b;
    layer1_outputs(9179) <= not b;
    layer1_outputs(9180) <= a and b;
    layer1_outputs(9181) <= not (a and b);
    layer1_outputs(9182) <= not (a xor b);
    layer1_outputs(9183) <= not (a xor b);
    layer1_outputs(9184) <= a or b;
    layer1_outputs(9185) <= not b or a;
    layer1_outputs(9186) <= '0';
    layer1_outputs(9187) <= b and not a;
    layer1_outputs(9188) <= a xor b;
    layer1_outputs(9189) <= a and not b;
    layer1_outputs(9190) <= not b or a;
    layer1_outputs(9191) <= not b or a;
    layer1_outputs(9192) <= not a;
    layer1_outputs(9193) <= a and b;
    layer1_outputs(9194) <= not (a and b);
    layer1_outputs(9195) <= a;
    layer1_outputs(9196) <= not (a xor b);
    layer1_outputs(9197) <= not (a or b);
    layer1_outputs(9198) <= not (a xor b);
    layer1_outputs(9199) <= a and b;
    layer1_outputs(9200) <= not b or a;
    layer1_outputs(9201) <= a xor b;
    layer1_outputs(9202) <= a xor b;
    layer1_outputs(9203) <= a and b;
    layer1_outputs(9204) <= a;
    layer1_outputs(9205) <= b;
    layer1_outputs(9206) <= not a or b;
    layer1_outputs(9207) <= a or b;
    layer1_outputs(9208) <= not b or a;
    layer1_outputs(9209) <= not a;
    layer1_outputs(9210) <= a or b;
    layer1_outputs(9211) <= not (a xor b);
    layer1_outputs(9212) <= not (a xor b);
    layer1_outputs(9213) <= a;
    layer1_outputs(9214) <= b;
    layer1_outputs(9215) <= a;
    layer1_outputs(9216) <= a and not b;
    layer1_outputs(9217) <= not a or b;
    layer1_outputs(9218) <= a or b;
    layer1_outputs(9219) <= a and b;
    layer1_outputs(9220) <= a;
    layer1_outputs(9221) <= a and not b;
    layer1_outputs(9222) <= a;
    layer1_outputs(9223) <= not b;
    layer1_outputs(9224) <= not a or b;
    layer1_outputs(9225) <= not a;
    layer1_outputs(9226) <= b;
    layer1_outputs(9227) <= a;
    layer1_outputs(9228) <= a and b;
    layer1_outputs(9229) <= a;
    layer1_outputs(9230) <= a and b;
    layer1_outputs(9231) <= not a or b;
    layer1_outputs(9232) <= a or b;
    layer1_outputs(9233) <= not a;
    layer1_outputs(9234) <= not a;
    layer1_outputs(9235) <= not a;
    layer1_outputs(9236) <= not b or a;
    layer1_outputs(9237) <= not a;
    layer1_outputs(9238) <= not b;
    layer1_outputs(9239) <= not b;
    layer1_outputs(9240) <= not (a or b);
    layer1_outputs(9241) <= not (a or b);
    layer1_outputs(9242) <= a and b;
    layer1_outputs(9243) <= not a;
    layer1_outputs(9244) <= a and not b;
    layer1_outputs(9245) <= not (a and b);
    layer1_outputs(9246) <= '1';
    layer1_outputs(9247) <= a xor b;
    layer1_outputs(9248) <= not a;
    layer1_outputs(9249) <= a xor b;
    layer1_outputs(9250) <= b and not a;
    layer1_outputs(9251) <= not a;
    layer1_outputs(9252) <= b;
    layer1_outputs(9253) <= not (a or b);
    layer1_outputs(9254) <= not (a and b);
    layer1_outputs(9255) <= not b;
    layer1_outputs(9256) <= b;
    layer1_outputs(9257) <= b and not a;
    layer1_outputs(9258) <= b and not a;
    layer1_outputs(9259) <= not a;
    layer1_outputs(9260) <= not a;
    layer1_outputs(9261) <= not (a or b);
    layer1_outputs(9262) <= b;
    layer1_outputs(9263) <= not b;
    layer1_outputs(9264) <= not b;
    layer1_outputs(9265) <= a;
    layer1_outputs(9266) <= not (a and b);
    layer1_outputs(9267) <= b;
    layer1_outputs(9268) <= b and not a;
    layer1_outputs(9269) <= a or b;
    layer1_outputs(9270) <= not a;
    layer1_outputs(9271) <= not (a and b);
    layer1_outputs(9272) <= not (a or b);
    layer1_outputs(9273) <= not a or b;
    layer1_outputs(9274) <= b;
    layer1_outputs(9275) <= a;
    layer1_outputs(9276) <= a;
    layer1_outputs(9277) <= a xor b;
    layer1_outputs(9278) <= '0';
    layer1_outputs(9279) <= a and not b;
    layer1_outputs(9280) <= not b;
    layer1_outputs(9281) <= not (a and b);
    layer1_outputs(9282) <= a and b;
    layer1_outputs(9283) <= not (a xor b);
    layer1_outputs(9284) <= a xor b;
    layer1_outputs(9285) <= not (a or b);
    layer1_outputs(9286) <= not a;
    layer1_outputs(9287) <= a;
    layer1_outputs(9288) <= not a or b;
    layer1_outputs(9289) <= a;
    layer1_outputs(9290) <= a and not b;
    layer1_outputs(9291) <= '1';
    layer1_outputs(9292) <= not a;
    layer1_outputs(9293) <= b;
    layer1_outputs(9294) <= a and b;
    layer1_outputs(9295) <= not (a or b);
    layer1_outputs(9296) <= not a or b;
    layer1_outputs(9297) <= a or b;
    layer1_outputs(9298) <= a xor b;
    layer1_outputs(9299) <= a;
    layer1_outputs(9300) <= not (a xor b);
    layer1_outputs(9301) <= a or b;
    layer1_outputs(9302) <= a;
    layer1_outputs(9303) <= not a or b;
    layer1_outputs(9304) <= a and not b;
    layer1_outputs(9305) <= not (a xor b);
    layer1_outputs(9306) <= a and b;
    layer1_outputs(9307) <= b and not a;
    layer1_outputs(9308) <= a or b;
    layer1_outputs(9309) <= a or b;
    layer1_outputs(9310) <= a;
    layer1_outputs(9311) <= not b;
    layer1_outputs(9312) <= not (a xor b);
    layer1_outputs(9313) <= b;
    layer1_outputs(9314) <= b;
    layer1_outputs(9315) <= not (a and b);
    layer1_outputs(9316) <= b and not a;
    layer1_outputs(9317) <= not b;
    layer1_outputs(9318) <= not b;
    layer1_outputs(9319) <= not (a or b);
    layer1_outputs(9320) <= not b or a;
    layer1_outputs(9321) <= '1';
    layer1_outputs(9322) <= a and b;
    layer1_outputs(9323) <= not a or b;
    layer1_outputs(9324) <= not b or a;
    layer1_outputs(9325) <= a or b;
    layer1_outputs(9326) <= not (a xor b);
    layer1_outputs(9327) <= a and not b;
    layer1_outputs(9328) <= b;
    layer1_outputs(9329) <= not (a and b);
    layer1_outputs(9330) <= not (a xor b);
    layer1_outputs(9331) <= not a or b;
    layer1_outputs(9332) <= not a;
    layer1_outputs(9333) <= a or b;
    layer1_outputs(9334) <= b;
    layer1_outputs(9335) <= a xor b;
    layer1_outputs(9336) <= not b;
    layer1_outputs(9337) <= not b or a;
    layer1_outputs(9338) <= not b or a;
    layer1_outputs(9339) <= a and b;
    layer1_outputs(9340) <= a and b;
    layer1_outputs(9341) <= a and not b;
    layer1_outputs(9342) <= not a;
    layer1_outputs(9343) <= a and not b;
    layer1_outputs(9344) <= b;
    layer1_outputs(9345) <= not (a xor b);
    layer1_outputs(9346) <= not (a or b);
    layer1_outputs(9347) <= not a or b;
    layer1_outputs(9348) <= b and not a;
    layer1_outputs(9349) <= a;
    layer1_outputs(9350) <= a xor b;
    layer1_outputs(9351) <= a;
    layer1_outputs(9352) <= a and not b;
    layer1_outputs(9353) <= not (a xor b);
    layer1_outputs(9354) <= a xor b;
    layer1_outputs(9355) <= '0';
    layer1_outputs(9356) <= not (a and b);
    layer1_outputs(9357) <= a and not b;
    layer1_outputs(9358) <= not a;
    layer1_outputs(9359) <= not b;
    layer1_outputs(9360) <= not b or a;
    layer1_outputs(9361) <= b;
    layer1_outputs(9362) <= a;
    layer1_outputs(9363) <= b and not a;
    layer1_outputs(9364) <= '0';
    layer1_outputs(9365) <= not (a or b);
    layer1_outputs(9366) <= a or b;
    layer1_outputs(9367) <= a and b;
    layer1_outputs(9368) <= b and not a;
    layer1_outputs(9369) <= not a;
    layer1_outputs(9370) <= b;
    layer1_outputs(9371) <= a;
    layer1_outputs(9372) <= not b;
    layer1_outputs(9373) <= a and b;
    layer1_outputs(9374) <= a;
    layer1_outputs(9375) <= not (a or b);
    layer1_outputs(9376) <= a xor b;
    layer1_outputs(9377) <= a;
    layer1_outputs(9378) <= not (a xor b);
    layer1_outputs(9379) <= not (a and b);
    layer1_outputs(9380) <= not (a xor b);
    layer1_outputs(9381) <= not a;
    layer1_outputs(9382) <= a;
    layer1_outputs(9383) <= not a or b;
    layer1_outputs(9384) <= a and b;
    layer1_outputs(9385) <= a and not b;
    layer1_outputs(9386) <= not b;
    layer1_outputs(9387) <= not b or a;
    layer1_outputs(9388) <= not (a xor b);
    layer1_outputs(9389) <= b and not a;
    layer1_outputs(9390) <= not (a and b);
    layer1_outputs(9391) <= b;
    layer1_outputs(9392) <= a and b;
    layer1_outputs(9393) <= not b;
    layer1_outputs(9394) <= not (a xor b);
    layer1_outputs(9395) <= not (a and b);
    layer1_outputs(9396) <= not a;
    layer1_outputs(9397) <= a xor b;
    layer1_outputs(9398) <= b;
    layer1_outputs(9399) <= b;
    layer1_outputs(9400) <= not a;
    layer1_outputs(9401) <= a and not b;
    layer1_outputs(9402) <= a and b;
    layer1_outputs(9403) <= b;
    layer1_outputs(9404) <= not (a xor b);
    layer1_outputs(9405) <= not a or b;
    layer1_outputs(9406) <= not b;
    layer1_outputs(9407) <= not (a or b);
    layer1_outputs(9408) <= a xor b;
    layer1_outputs(9409) <= not a or b;
    layer1_outputs(9410) <= not (a or b);
    layer1_outputs(9411) <= b;
    layer1_outputs(9412) <= '0';
    layer1_outputs(9413) <= b;
    layer1_outputs(9414) <= not (a or b);
    layer1_outputs(9415) <= a;
    layer1_outputs(9416) <= a;
    layer1_outputs(9417) <= a and b;
    layer1_outputs(9418) <= not (a or b);
    layer1_outputs(9419) <= not (a xor b);
    layer1_outputs(9420) <= not (a xor b);
    layer1_outputs(9421) <= a;
    layer1_outputs(9422) <= a xor b;
    layer1_outputs(9423) <= not b or a;
    layer1_outputs(9424) <= not a;
    layer1_outputs(9425) <= not (a and b);
    layer1_outputs(9426) <= a;
    layer1_outputs(9427) <= a and not b;
    layer1_outputs(9428) <= not b;
    layer1_outputs(9429) <= not (a and b);
    layer1_outputs(9430) <= not a or b;
    layer1_outputs(9431) <= not (a and b);
    layer1_outputs(9432) <= not b;
    layer1_outputs(9433) <= not a;
    layer1_outputs(9434) <= b;
    layer1_outputs(9435) <= a;
    layer1_outputs(9436) <= a xor b;
    layer1_outputs(9437) <= a and b;
    layer1_outputs(9438) <= not a;
    layer1_outputs(9439) <= a or b;
    layer1_outputs(9440) <= not b or a;
    layer1_outputs(9441) <= not a;
    layer1_outputs(9442) <= a;
    layer1_outputs(9443) <= not (a and b);
    layer1_outputs(9444) <= not b;
    layer1_outputs(9445) <= not a or b;
    layer1_outputs(9446) <= not b or a;
    layer1_outputs(9447) <= not (a xor b);
    layer1_outputs(9448) <= not a;
    layer1_outputs(9449) <= not (a or b);
    layer1_outputs(9450) <= a;
    layer1_outputs(9451) <= not b;
    layer1_outputs(9452) <= a and not b;
    layer1_outputs(9453) <= not (a or b);
    layer1_outputs(9454) <= not (a and b);
    layer1_outputs(9455) <= not (a or b);
    layer1_outputs(9456) <= b;
    layer1_outputs(9457) <= b;
    layer1_outputs(9458) <= a xor b;
    layer1_outputs(9459) <= '0';
    layer1_outputs(9460) <= b;
    layer1_outputs(9461) <= not b;
    layer1_outputs(9462) <= not (a xor b);
    layer1_outputs(9463) <= b;
    layer1_outputs(9464) <= a xor b;
    layer1_outputs(9465) <= not (a and b);
    layer1_outputs(9466) <= a and b;
    layer1_outputs(9467) <= a;
    layer1_outputs(9468) <= not (a and b);
    layer1_outputs(9469) <= a xor b;
    layer1_outputs(9470) <= a xor b;
    layer1_outputs(9471) <= a;
    layer1_outputs(9472) <= b and not a;
    layer1_outputs(9473) <= b and not a;
    layer1_outputs(9474) <= a;
    layer1_outputs(9475) <= b and not a;
    layer1_outputs(9476) <= not a;
    layer1_outputs(9477) <= b and not a;
    layer1_outputs(9478) <= a xor b;
    layer1_outputs(9479) <= a and b;
    layer1_outputs(9480) <= a and b;
    layer1_outputs(9481) <= a or b;
    layer1_outputs(9482) <= not a or b;
    layer1_outputs(9483) <= a and b;
    layer1_outputs(9484) <= a;
    layer1_outputs(9485) <= not b or a;
    layer1_outputs(9486) <= not b;
    layer1_outputs(9487) <= not (a and b);
    layer1_outputs(9488) <= b;
    layer1_outputs(9489) <= not (a xor b);
    layer1_outputs(9490) <= a xor b;
    layer1_outputs(9491) <= a xor b;
    layer1_outputs(9492) <= not (a and b);
    layer1_outputs(9493) <= not (a xor b);
    layer1_outputs(9494) <= not a;
    layer1_outputs(9495) <= a xor b;
    layer1_outputs(9496) <= not (a xor b);
    layer1_outputs(9497) <= a xor b;
    layer1_outputs(9498) <= not b or a;
    layer1_outputs(9499) <= a or b;
    layer1_outputs(9500) <= b;
    layer1_outputs(9501) <= a;
    layer1_outputs(9502) <= a and not b;
    layer1_outputs(9503) <= not b or a;
    layer1_outputs(9504) <= a and not b;
    layer1_outputs(9505) <= not b;
    layer1_outputs(9506) <= a or b;
    layer1_outputs(9507) <= not a;
    layer1_outputs(9508) <= a;
    layer1_outputs(9509) <= not b;
    layer1_outputs(9510) <= b;
    layer1_outputs(9511) <= a and b;
    layer1_outputs(9512) <= '0';
    layer1_outputs(9513) <= not (a and b);
    layer1_outputs(9514) <= not a or b;
    layer1_outputs(9515) <= not a;
    layer1_outputs(9516) <= a and b;
    layer1_outputs(9517) <= a and not b;
    layer1_outputs(9518) <= not (a or b);
    layer1_outputs(9519) <= not (a and b);
    layer1_outputs(9520) <= not (a or b);
    layer1_outputs(9521) <= a;
    layer1_outputs(9522) <= not (a and b);
    layer1_outputs(9523) <= not a or b;
    layer1_outputs(9524) <= not (a and b);
    layer1_outputs(9525) <= not a;
    layer1_outputs(9526) <= not (a xor b);
    layer1_outputs(9527) <= a xor b;
    layer1_outputs(9528) <= not (a or b);
    layer1_outputs(9529) <= b;
    layer1_outputs(9530) <= not b;
    layer1_outputs(9531) <= b and not a;
    layer1_outputs(9532) <= a and b;
    layer1_outputs(9533) <= not (a or b);
    layer1_outputs(9534) <= a;
    layer1_outputs(9535) <= a or b;
    layer1_outputs(9536) <= not b;
    layer1_outputs(9537) <= a and b;
    layer1_outputs(9538) <= a or b;
    layer1_outputs(9539) <= not a;
    layer1_outputs(9540) <= not a or b;
    layer1_outputs(9541) <= not b;
    layer1_outputs(9542) <= a xor b;
    layer1_outputs(9543) <= not (a or b);
    layer1_outputs(9544) <= a xor b;
    layer1_outputs(9545) <= not (a xor b);
    layer1_outputs(9546) <= not a or b;
    layer1_outputs(9547) <= a and not b;
    layer1_outputs(9548) <= a;
    layer1_outputs(9549) <= b;
    layer1_outputs(9550) <= not (a or b);
    layer1_outputs(9551) <= not a or b;
    layer1_outputs(9552) <= not (a xor b);
    layer1_outputs(9553) <= a xor b;
    layer1_outputs(9554) <= a;
    layer1_outputs(9555) <= not b or a;
    layer1_outputs(9556) <= b;
    layer1_outputs(9557) <= b and not a;
    layer1_outputs(9558) <= not b or a;
    layer1_outputs(9559) <= b and not a;
    layer1_outputs(9560) <= not b or a;
    layer1_outputs(9561) <= b;
    layer1_outputs(9562) <= a and not b;
    layer1_outputs(9563) <= a;
    layer1_outputs(9564) <= a and not b;
    layer1_outputs(9565) <= not b;
    layer1_outputs(9566) <= not b or a;
    layer1_outputs(9567) <= b and not a;
    layer1_outputs(9568) <= not b;
    layer1_outputs(9569) <= not a;
    layer1_outputs(9570) <= not (a or b);
    layer1_outputs(9571) <= b and not a;
    layer1_outputs(9572) <= not a;
    layer1_outputs(9573) <= not a or b;
    layer1_outputs(9574) <= not b;
    layer1_outputs(9575) <= not b or a;
    layer1_outputs(9576) <= not (a or b);
    layer1_outputs(9577) <= a and b;
    layer1_outputs(9578) <= a and not b;
    layer1_outputs(9579) <= not (a and b);
    layer1_outputs(9580) <= not (a xor b);
    layer1_outputs(9581) <= not a or b;
    layer1_outputs(9582) <= not b or a;
    layer1_outputs(9583) <= not b or a;
    layer1_outputs(9584) <= not a;
    layer1_outputs(9585) <= not b;
    layer1_outputs(9586) <= not (a xor b);
    layer1_outputs(9587) <= not a;
    layer1_outputs(9588) <= not (a or b);
    layer1_outputs(9589) <= not (a or b);
    layer1_outputs(9590) <= not a;
    layer1_outputs(9591) <= not (a xor b);
    layer1_outputs(9592) <= a and b;
    layer1_outputs(9593) <= b;
    layer1_outputs(9594) <= b;
    layer1_outputs(9595) <= a and not b;
    layer1_outputs(9596) <= not (a or b);
    layer1_outputs(9597) <= not b or a;
    layer1_outputs(9598) <= not a;
    layer1_outputs(9599) <= not (a and b);
    layer1_outputs(9600) <= b and not a;
    layer1_outputs(9601) <= b and not a;
    layer1_outputs(9602) <= not b or a;
    layer1_outputs(9603) <= a;
    layer1_outputs(9604) <= not (a or b);
    layer1_outputs(9605) <= not a or b;
    layer1_outputs(9606) <= not a or b;
    layer1_outputs(9607) <= a or b;
    layer1_outputs(9608) <= b;
    layer1_outputs(9609) <= b;
    layer1_outputs(9610) <= b and not a;
    layer1_outputs(9611) <= a or b;
    layer1_outputs(9612) <= a;
    layer1_outputs(9613) <= a or b;
    layer1_outputs(9614) <= not a;
    layer1_outputs(9615) <= a or b;
    layer1_outputs(9616) <= a and not b;
    layer1_outputs(9617) <= not a;
    layer1_outputs(9618) <= not (a or b);
    layer1_outputs(9619) <= a and not b;
    layer1_outputs(9620) <= a and not b;
    layer1_outputs(9621) <= not b;
    layer1_outputs(9622) <= not b or a;
    layer1_outputs(9623) <= a and not b;
    layer1_outputs(9624) <= not (a xor b);
    layer1_outputs(9625) <= not a;
    layer1_outputs(9626) <= a or b;
    layer1_outputs(9627) <= a xor b;
    layer1_outputs(9628) <= a xor b;
    layer1_outputs(9629) <= a;
    layer1_outputs(9630) <= b and not a;
    layer1_outputs(9631) <= not b;
    layer1_outputs(9632) <= a xor b;
    layer1_outputs(9633) <= a or b;
    layer1_outputs(9634) <= a xor b;
    layer1_outputs(9635) <= a and b;
    layer1_outputs(9636) <= not (a or b);
    layer1_outputs(9637) <= not a;
    layer1_outputs(9638) <= not a or b;
    layer1_outputs(9639) <= not a;
    layer1_outputs(9640) <= a;
    layer1_outputs(9641) <= not a;
    layer1_outputs(9642) <= a or b;
    layer1_outputs(9643) <= a xor b;
    layer1_outputs(9644) <= not (a xor b);
    layer1_outputs(9645) <= not a;
    layer1_outputs(9646) <= not b or a;
    layer1_outputs(9647) <= not a;
    layer1_outputs(9648) <= a xor b;
    layer1_outputs(9649) <= b;
    layer1_outputs(9650) <= not b or a;
    layer1_outputs(9651) <= not (a and b);
    layer1_outputs(9652) <= a;
    layer1_outputs(9653) <= not a;
    layer1_outputs(9654) <= a or b;
    layer1_outputs(9655) <= a or b;
    layer1_outputs(9656) <= not a;
    layer1_outputs(9657) <= a;
    layer1_outputs(9658) <= a or b;
    layer1_outputs(9659) <= a and not b;
    layer1_outputs(9660) <= not a or b;
    layer1_outputs(9661) <= not b;
    layer1_outputs(9662) <= a and not b;
    layer1_outputs(9663) <= a or b;
    layer1_outputs(9664) <= not (a xor b);
    layer1_outputs(9665) <= not b or a;
    layer1_outputs(9666) <= a;
    layer1_outputs(9667) <= b and not a;
    layer1_outputs(9668) <= b;
    layer1_outputs(9669) <= b;
    layer1_outputs(9670) <= not (a xor b);
    layer1_outputs(9671) <= not a or b;
    layer1_outputs(9672) <= a or b;
    layer1_outputs(9673) <= a or b;
    layer1_outputs(9674) <= b;
    layer1_outputs(9675) <= a or b;
    layer1_outputs(9676) <= a;
    layer1_outputs(9677) <= not b;
    layer1_outputs(9678) <= not (a or b);
    layer1_outputs(9679) <= a and not b;
    layer1_outputs(9680) <= not (a xor b);
    layer1_outputs(9681) <= not (a xor b);
    layer1_outputs(9682) <= a xor b;
    layer1_outputs(9683) <= not (a xor b);
    layer1_outputs(9684) <= not b or a;
    layer1_outputs(9685) <= a;
    layer1_outputs(9686) <= not a;
    layer1_outputs(9687) <= b and not a;
    layer1_outputs(9688) <= a or b;
    layer1_outputs(9689) <= b and not a;
    layer1_outputs(9690) <= a or b;
    layer1_outputs(9691) <= not (a xor b);
    layer1_outputs(9692) <= not (a xor b);
    layer1_outputs(9693) <= not a or b;
    layer1_outputs(9694) <= not a;
    layer1_outputs(9695) <= not a;
    layer1_outputs(9696) <= not (a and b);
    layer1_outputs(9697) <= b and not a;
    layer1_outputs(9698) <= not (a and b);
    layer1_outputs(9699) <= b;
    layer1_outputs(9700) <= a and not b;
    layer1_outputs(9701) <= not (a and b);
    layer1_outputs(9702) <= a and b;
    layer1_outputs(9703) <= a xor b;
    layer1_outputs(9704) <= a and not b;
    layer1_outputs(9705) <= not (a or b);
    layer1_outputs(9706) <= not a or b;
    layer1_outputs(9707) <= not b or a;
    layer1_outputs(9708) <= not (a xor b);
    layer1_outputs(9709) <= not a or b;
    layer1_outputs(9710) <= not b;
    layer1_outputs(9711) <= not a or b;
    layer1_outputs(9712) <= not (a xor b);
    layer1_outputs(9713) <= a xor b;
    layer1_outputs(9714) <= not (a or b);
    layer1_outputs(9715) <= a and not b;
    layer1_outputs(9716) <= a and not b;
    layer1_outputs(9717) <= not (a and b);
    layer1_outputs(9718) <= not (a and b);
    layer1_outputs(9719) <= not a;
    layer1_outputs(9720) <= not (a and b);
    layer1_outputs(9721) <= not b;
    layer1_outputs(9722) <= not b or a;
    layer1_outputs(9723) <= not b or a;
    layer1_outputs(9724) <= a;
    layer1_outputs(9725) <= a;
    layer1_outputs(9726) <= a;
    layer1_outputs(9727) <= not (a and b);
    layer1_outputs(9728) <= a and not b;
    layer1_outputs(9729) <= a or b;
    layer1_outputs(9730) <= not (a and b);
    layer1_outputs(9731) <= a and not b;
    layer1_outputs(9732) <= not b;
    layer1_outputs(9733) <= not (a and b);
    layer1_outputs(9734) <= a xor b;
    layer1_outputs(9735) <= a or b;
    layer1_outputs(9736) <= not b;
    layer1_outputs(9737) <= b and not a;
    layer1_outputs(9738) <= not a;
    layer1_outputs(9739) <= not (a or b);
    layer1_outputs(9740) <= not b or a;
    layer1_outputs(9741) <= a;
    layer1_outputs(9742) <= b and not a;
    layer1_outputs(9743) <= b;
    layer1_outputs(9744) <= b;
    layer1_outputs(9745) <= not a or b;
    layer1_outputs(9746) <= not (a xor b);
    layer1_outputs(9747) <= not b;
    layer1_outputs(9748) <= b and not a;
    layer1_outputs(9749) <= a and b;
    layer1_outputs(9750) <= a;
    layer1_outputs(9751) <= not b;
    layer1_outputs(9752) <= not a or b;
    layer1_outputs(9753) <= not b;
    layer1_outputs(9754) <= not a or b;
    layer1_outputs(9755) <= a;
    layer1_outputs(9756) <= not a;
    layer1_outputs(9757) <= not (a or b);
    layer1_outputs(9758) <= a;
    layer1_outputs(9759) <= a;
    layer1_outputs(9760) <= a and b;
    layer1_outputs(9761) <= a or b;
    layer1_outputs(9762) <= not (a and b);
    layer1_outputs(9763) <= a xor b;
    layer1_outputs(9764) <= not (a or b);
    layer1_outputs(9765) <= a;
    layer1_outputs(9766) <= a or b;
    layer1_outputs(9767) <= b;
    layer1_outputs(9768) <= not (a xor b);
    layer1_outputs(9769) <= not b or a;
    layer1_outputs(9770) <= not a;
    layer1_outputs(9771) <= not (a xor b);
    layer1_outputs(9772) <= a xor b;
    layer1_outputs(9773) <= not (a or b);
    layer1_outputs(9774) <= not (a xor b);
    layer1_outputs(9775) <= not a or b;
    layer1_outputs(9776) <= b and not a;
    layer1_outputs(9777) <= not b or a;
    layer1_outputs(9778) <= b and not a;
    layer1_outputs(9779) <= not (a and b);
    layer1_outputs(9780) <= a xor b;
    layer1_outputs(9781) <= not (a xor b);
    layer1_outputs(9782) <= a xor b;
    layer1_outputs(9783) <= '0';
    layer1_outputs(9784) <= not (a xor b);
    layer1_outputs(9785) <= not (a xor b);
    layer1_outputs(9786) <= not b;
    layer1_outputs(9787) <= '0';
    layer1_outputs(9788) <= not (a xor b);
    layer1_outputs(9789) <= not b;
    layer1_outputs(9790) <= a or b;
    layer1_outputs(9791) <= a and not b;
    layer1_outputs(9792) <= a;
    layer1_outputs(9793) <= a and b;
    layer1_outputs(9794) <= not (a or b);
    layer1_outputs(9795) <= a and not b;
    layer1_outputs(9796) <= b and not a;
    layer1_outputs(9797) <= a and not b;
    layer1_outputs(9798) <= not (a or b);
    layer1_outputs(9799) <= not b or a;
    layer1_outputs(9800) <= not b or a;
    layer1_outputs(9801) <= not (a and b);
    layer1_outputs(9802) <= a;
    layer1_outputs(9803) <= not b;
    layer1_outputs(9804) <= not (a and b);
    layer1_outputs(9805) <= not (a and b);
    layer1_outputs(9806) <= b;
    layer1_outputs(9807) <= not b;
    layer1_outputs(9808) <= not b or a;
    layer1_outputs(9809) <= a or b;
    layer1_outputs(9810) <= b and not a;
    layer1_outputs(9811) <= not a;
    layer1_outputs(9812) <= b and not a;
    layer1_outputs(9813) <= a xor b;
    layer1_outputs(9814) <= b and not a;
    layer1_outputs(9815) <= not b;
    layer1_outputs(9816) <= a;
    layer1_outputs(9817) <= not (a xor b);
    layer1_outputs(9818) <= a or b;
    layer1_outputs(9819) <= a;
    layer1_outputs(9820) <= not (a xor b);
    layer1_outputs(9821) <= not a;
    layer1_outputs(9822) <= not b or a;
    layer1_outputs(9823) <= b;
    layer1_outputs(9824) <= not a;
    layer1_outputs(9825) <= not (a xor b);
    layer1_outputs(9826) <= not a;
    layer1_outputs(9827) <= not a or b;
    layer1_outputs(9828) <= a xor b;
    layer1_outputs(9829) <= not (a or b);
    layer1_outputs(9830) <= b;
    layer1_outputs(9831) <= not b;
    layer1_outputs(9832) <= a;
    layer1_outputs(9833) <= a and b;
    layer1_outputs(9834) <= not (a or b);
    layer1_outputs(9835) <= not a;
    layer1_outputs(9836) <= not a;
    layer1_outputs(9837) <= not (a xor b);
    layer1_outputs(9838) <= not a;
    layer1_outputs(9839) <= not b or a;
    layer1_outputs(9840) <= a or b;
    layer1_outputs(9841) <= a and b;
    layer1_outputs(9842) <= a xor b;
    layer1_outputs(9843) <= b;
    layer1_outputs(9844) <= b;
    layer1_outputs(9845) <= not (a xor b);
    layer1_outputs(9846) <= not (a xor b);
    layer1_outputs(9847) <= a xor b;
    layer1_outputs(9848) <= '0';
    layer1_outputs(9849) <= not a or b;
    layer1_outputs(9850) <= a or b;
    layer1_outputs(9851) <= '0';
    layer1_outputs(9852) <= a;
    layer1_outputs(9853) <= not (a or b);
    layer1_outputs(9854) <= a xor b;
    layer1_outputs(9855) <= a or b;
    layer1_outputs(9856) <= not b;
    layer1_outputs(9857) <= not a;
    layer1_outputs(9858) <= not (a or b);
    layer1_outputs(9859) <= a and not b;
    layer1_outputs(9860) <= b;
    layer1_outputs(9861) <= not b;
    layer1_outputs(9862) <= b and not a;
    layer1_outputs(9863) <= not b or a;
    layer1_outputs(9864) <= not b;
    layer1_outputs(9865) <= a;
    layer1_outputs(9866) <= b and not a;
    layer1_outputs(9867) <= not b;
    layer1_outputs(9868) <= a and b;
    layer1_outputs(9869) <= a;
    layer1_outputs(9870) <= a;
    layer1_outputs(9871) <= a;
    layer1_outputs(9872) <= not a;
    layer1_outputs(9873) <= b;
    layer1_outputs(9874) <= a and b;
    layer1_outputs(9875) <= not (a xor b);
    layer1_outputs(9876) <= not (a and b);
    layer1_outputs(9877) <= a;
    layer1_outputs(9878) <= b;
    layer1_outputs(9879) <= a and b;
    layer1_outputs(9880) <= not b or a;
    layer1_outputs(9881) <= a xor b;
    layer1_outputs(9882) <= b and not a;
    layer1_outputs(9883) <= b and not a;
    layer1_outputs(9884) <= a or b;
    layer1_outputs(9885) <= not (a or b);
    layer1_outputs(9886) <= not a or b;
    layer1_outputs(9887) <= not (a xor b);
    layer1_outputs(9888) <= a and b;
    layer1_outputs(9889) <= a and b;
    layer1_outputs(9890) <= a;
    layer1_outputs(9891) <= a or b;
    layer1_outputs(9892) <= b;
    layer1_outputs(9893) <= b;
    layer1_outputs(9894) <= a or b;
    layer1_outputs(9895) <= a and b;
    layer1_outputs(9896) <= not b;
    layer1_outputs(9897) <= a xor b;
    layer1_outputs(9898) <= not b;
    layer1_outputs(9899) <= a and b;
    layer1_outputs(9900) <= b;
    layer1_outputs(9901) <= b;
    layer1_outputs(9902) <= a;
    layer1_outputs(9903) <= not a;
    layer1_outputs(9904) <= not (a xor b);
    layer1_outputs(9905) <= a;
    layer1_outputs(9906) <= not a;
    layer1_outputs(9907) <= not b;
    layer1_outputs(9908) <= b and not a;
    layer1_outputs(9909) <= not (a and b);
    layer1_outputs(9910) <= '1';
    layer1_outputs(9911) <= not b;
    layer1_outputs(9912) <= not b;
    layer1_outputs(9913) <= a;
    layer1_outputs(9914) <= a;
    layer1_outputs(9915) <= not (a xor b);
    layer1_outputs(9916) <= not b;
    layer1_outputs(9917) <= not b or a;
    layer1_outputs(9918) <= a xor b;
    layer1_outputs(9919) <= a and not b;
    layer1_outputs(9920) <= not a or b;
    layer1_outputs(9921) <= b and not a;
    layer1_outputs(9922) <= not b or a;
    layer1_outputs(9923) <= a;
    layer1_outputs(9924) <= not b or a;
    layer1_outputs(9925) <= b;
    layer1_outputs(9926) <= a;
    layer1_outputs(9927) <= not a or b;
    layer1_outputs(9928) <= not b;
    layer1_outputs(9929) <= a;
    layer1_outputs(9930) <= b;
    layer1_outputs(9931) <= a xor b;
    layer1_outputs(9932) <= a and not b;
    layer1_outputs(9933) <= b;
    layer1_outputs(9934) <= not (a and b);
    layer1_outputs(9935) <= a and not b;
    layer1_outputs(9936) <= not (a xor b);
    layer1_outputs(9937) <= a or b;
    layer1_outputs(9938) <= not (a xor b);
    layer1_outputs(9939) <= a xor b;
    layer1_outputs(9940) <= not a;
    layer1_outputs(9941) <= not (a xor b);
    layer1_outputs(9942) <= not b or a;
    layer1_outputs(9943) <= a;
    layer1_outputs(9944) <= not (a and b);
    layer1_outputs(9945) <= not (a or b);
    layer1_outputs(9946) <= not (a or b);
    layer1_outputs(9947) <= a xor b;
    layer1_outputs(9948) <= a and b;
    layer1_outputs(9949) <= not a;
    layer1_outputs(9950) <= not (a xor b);
    layer1_outputs(9951) <= b and not a;
    layer1_outputs(9952) <= not a;
    layer1_outputs(9953) <= not (a and b);
    layer1_outputs(9954) <= not (a and b);
    layer1_outputs(9955) <= not b or a;
    layer1_outputs(9956) <= a;
    layer1_outputs(9957) <= a or b;
    layer1_outputs(9958) <= not b or a;
    layer1_outputs(9959) <= not (a or b);
    layer1_outputs(9960) <= not (a xor b);
    layer1_outputs(9961) <= not b;
    layer1_outputs(9962) <= a;
    layer1_outputs(9963) <= a;
    layer1_outputs(9964) <= not a;
    layer1_outputs(9965) <= a xor b;
    layer1_outputs(9966) <= a or b;
    layer1_outputs(9967) <= not a;
    layer1_outputs(9968) <= not b or a;
    layer1_outputs(9969) <= not (a xor b);
    layer1_outputs(9970) <= a xor b;
    layer1_outputs(9971) <= not a or b;
    layer1_outputs(9972) <= not (a and b);
    layer1_outputs(9973) <= a;
    layer1_outputs(9974) <= not a;
    layer1_outputs(9975) <= a;
    layer1_outputs(9976) <= not a;
    layer1_outputs(9977) <= a and b;
    layer1_outputs(9978) <= a and b;
    layer1_outputs(9979) <= b and not a;
    layer1_outputs(9980) <= not (a xor b);
    layer1_outputs(9981) <= not (a and b);
    layer1_outputs(9982) <= not b;
    layer1_outputs(9983) <= not b;
    layer1_outputs(9984) <= b and not a;
    layer1_outputs(9985) <= not (a xor b);
    layer1_outputs(9986) <= not b or a;
    layer1_outputs(9987) <= not b or a;
    layer1_outputs(9988) <= a;
    layer1_outputs(9989) <= a and not b;
    layer1_outputs(9990) <= not (a xor b);
    layer1_outputs(9991) <= a xor b;
    layer1_outputs(9992) <= not b;
    layer1_outputs(9993) <= not (a or b);
    layer1_outputs(9994) <= a and not b;
    layer1_outputs(9995) <= not b or a;
    layer1_outputs(9996) <= a xor b;
    layer1_outputs(9997) <= not (a and b);
    layer1_outputs(9998) <= not (a xor b);
    layer1_outputs(9999) <= b and not a;
    layer1_outputs(10000) <= a;
    layer1_outputs(10001) <= not a;
    layer1_outputs(10002) <= not a;
    layer1_outputs(10003) <= not b;
    layer1_outputs(10004) <= b;
    layer1_outputs(10005) <= not a;
    layer1_outputs(10006) <= b and not a;
    layer1_outputs(10007) <= not (a or b);
    layer1_outputs(10008) <= a;
    layer1_outputs(10009) <= a;
    layer1_outputs(10010) <= not a;
    layer1_outputs(10011) <= not (a and b);
    layer1_outputs(10012) <= a and not b;
    layer1_outputs(10013) <= '0';
    layer1_outputs(10014) <= not (a or b);
    layer1_outputs(10015) <= not (a xor b);
    layer1_outputs(10016) <= a xor b;
    layer1_outputs(10017) <= not a;
    layer1_outputs(10018) <= not a;
    layer1_outputs(10019) <= a or b;
    layer1_outputs(10020) <= not (a and b);
    layer1_outputs(10021) <= not (a xor b);
    layer1_outputs(10022) <= a or b;
    layer1_outputs(10023) <= not a;
    layer1_outputs(10024) <= a and not b;
    layer1_outputs(10025) <= not (a and b);
    layer1_outputs(10026) <= a xor b;
    layer1_outputs(10027) <= not b or a;
    layer1_outputs(10028) <= b;
    layer1_outputs(10029) <= not a;
    layer1_outputs(10030) <= not (a or b);
    layer1_outputs(10031) <= not b or a;
    layer1_outputs(10032) <= not b or a;
    layer1_outputs(10033) <= a;
    layer1_outputs(10034) <= b;
    layer1_outputs(10035) <= not a;
    layer1_outputs(10036) <= not b;
    layer1_outputs(10037) <= not (a xor b);
    layer1_outputs(10038) <= a and not b;
    layer1_outputs(10039) <= a;
    layer1_outputs(10040) <= a;
    layer1_outputs(10041) <= not b;
    layer1_outputs(10042) <= b;
    layer1_outputs(10043) <= b;
    layer1_outputs(10044) <= '1';
    layer1_outputs(10045) <= not a;
    layer1_outputs(10046) <= not b;
    layer1_outputs(10047) <= a or b;
    layer1_outputs(10048) <= a;
    layer1_outputs(10049) <= not b or a;
    layer1_outputs(10050) <= not a;
    layer1_outputs(10051) <= not a;
    layer1_outputs(10052) <= not b;
    layer1_outputs(10053) <= a;
    layer1_outputs(10054) <= not b or a;
    layer1_outputs(10055) <= not (a xor b);
    layer1_outputs(10056) <= a and not b;
    layer1_outputs(10057) <= a or b;
    layer1_outputs(10058) <= not (a and b);
    layer1_outputs(10059) <= not b;
    layer1_outputs(10060) <= not (a or b);
    layer1_outputs(10061) <= not a;
    layer1_outputs(10062) <= not (a and b);
    layer1_outputs(10063) <= a and b;
    layer1_outputs(10064) <= a xor b;
    layer1_outputs(10065) <= not (a or b);
    layer1_outputs(10066) <= '0';
    layer1_outputs(10067) <= a and not b;
    layer1_outputs(10068) <= a;
    layer1_outputs(10069) <= not a or b;
    layer1_outputs(10070) <= not a or b;
    layer1_outputs(10071) <= a and b;
    layer1_outputs(10072) <= not a or b;
    layer1_outputs(10073) <= a and b;
    layer1_outputs(10074) <= not b;
    layer1_outputs(10075) <= not (a xor b);
    layer1_outputs(10076) <= not a or b;
    layer1_outputs(10077) <= a;
    layer1_outputs(10078) <= not a;
    layer1_outputs(10079) <= not a;
    layer1_outputs(10080) <= not a or b;
    layer1_outputs(10081) <= not a;
    layer1_outputs(10082) <= not b;
    layer1_outputs(10083) <= not b or a;
    layer1_outputs(10084) <= not a;
    layer1_outputs(10085) <= not a;
    layer1_outputs(10086) <= not b or a;
    layer1_outputs(10087) <= a or b;
    layer1_outputs(10088) <= a;
    layer1_outputs(10089) <= a and b;
    layer1_outputs(10090) <= a and b;
    layer1_outputs(10091) <= b and not a;
    layer1_outputs(10092) <= b;
    layer1_outputs(10093) <= a and not b;
    layer1_outputs(10094) <= a or b;
    layer1_outputs(10095) <= not b;
    layer1_outputs(10096) <= b;
    layer1_outputs(10097) <= a xor b;
    layer1_outputs(10098) <= not (a xor b);
    layer1_outputs(10099) <= a xor b;
    layer1_outputs(10100) <= a xor b;
    layer1_outputs(10101) <= a and b;
    layer1_outputs(10102) <= b and not a;
    layer1_outputs(10103) <= not b;
    layer1_outputs(10104) <= a and not b;
    layer1_outputs(10105) <= not (a xor b);
    layer1_outputs(10106) <= not b;
    layer1_outputs(10107) <= not b;
    layer1_outputs(10108) <= b;
    layer1_outputs(10109) <= a or b;
    layer1_outputs(10110) <= a and b;
    layer1_outputs(10111) <= not a;
    layer1_outputs(10112) <= not a;
    layer1_outputs(10113) <= a and b;
    layer1_outputs(10114) <= a xor b;
    layer1_outputs(10115) <= '0';
    layer1_outputs(10116) <= b;
    layer1_outputs(10117) <= not (a xor b);
    layer1_outputs(10118) <= a and b;
    layer1_outputs(10119) <= b;
    layer1_outputs(10120) <= a;
    layer1_outputs(10121) <= b;
    layer1_outputs(10122) <= not a;
    layer1_outputs(10123) <= a and b;
    layer1_outputs(10124) <= not a or b;
    layer1_outputs(10125) <= not (a xor b);
    layer1_outputs(10126) <= not b;
    layer1_outputs(10127) <= a and b;
    layer1_outputs(10128) <= not a;
    layer1_outputs(10129) <= not a;
    layer1_outputs(10130) <= not a or b;
    layer1_outputs(10131) <= a and b;
    layer1_outputs(10132) <= not a;
    layer1_outputs(10133) <= not (a and b);
    layer1_outputs(10134) <= b;
    layer1_outputs(10135) <= b;
    layer1_outputs(10136) <= a xor b;
    layer1_outputs(10137) <= a;
    layer1_outputs(10138) <= a xor b;
    layer1_outputs(10139) <= b;
    layer1_outputs(10140) <= not b;
    layer1_outputs(10141) <= not (a and b);
    layer1_outputs(10142) <= a;
    layer1_outputs(10143) <= not (a xor b);
    layer1_outputs(10144) <= not (a xor b);
    layer1_outputs(10145) <= not b;
    layer1_outputs(10146) <= a and b;
    layer1_outputs(10147) <= a xor b;
    layer1_outputs(10148) <= not (a xor b);
    layer1_outputs(10149) <= not b;
    layer1_outputs(10150) <= a or b;
    layer1_outputs(10151) <= not a or b;
    layer1_outputs(10152) <= not (a xor b);
    layer1_outputs(10153) <= not a;
    layer1_outputs(10154) <= not b or a;
    layer1_outputs(10155) <= a;
    layer1_outputs(10156) <= not b or a;
    layer1_outputs(10157) <= a and not b;
    layer1_outputs(10158) <= a and not b;
    layer1_outputs(10159) <= a and b;
    layer1_outputs(10160) <= a xor b;
    layer1_outputs(10161) <= a xor b;
    layer1_outputs(10162) <= not a or b;
    layer1_outputs(10163) <= not (a or b);
    layer1_outputs(10164) <= a and b;
    layer1_outputs(10165) <= not a or b;
    layer1_outputs(10166) <= a xor b;
    layer1_outputs(10167) <= not a;
    layer1_outputs(10168) <= a;
    layer1_outputs(10169) <= a and b;
    layer1_outputs(10170) <= b;
    layer1_outputs(10171) <= not (a or b);
    layer1_outputs(10172) <= a xor b;
    layer1_outputs(10173) <= b;
    layer1_outputs(10174) <= not a;
    layer1_outputs(10175) <= not (a or b);
    layer1_outputs(10176) <= a xor b;
    layer1_outputs(10177) <= a or b;
    layer1_outputs(10178) <= not a;
    layer1_outputs(10179) <= a xor b;
    layer1_outputs(10180) <= not a or b;
    layer1_outputs(10181) <= a and not b;
    layer1_outputs(10182) <= a and not b;
    layer1_outputs(10183) <= not (a or b);
    layer1_outputs(10184) <= not a;
    layer1_outputs(10185) <= not b or a;
    layer1_outputs(10186) <= a or b;
    layer1_outputs(10187) <= a and b;
    layer1_outputs(10188) <= b and not a;
    layer1_outputs(10189) <= not a or b;
    layer1_outputs(10190) <= a or b;
    layer1_outputs(10191) <= not (a or b);
    layer1_outputs(10192) <= not b;
    layer1_outputs(10193) <= not a;
    layer1_outputs(10194) <= b and not a;
    layer1_outputs(10195) <= b;
    layer1_outputs(10196) <= a and b;
    layer1_outputs(10197) <= not a;
    layer1_outputs(10198) <= not (a xor b);
    layer1_outputs(10199) <= not (a xor b);
    layer1_outputs(10200) <= not a or b;
    layer1_outputs(10201) <= not (a or b);
    layer1_outputs(10202) <= a xor b;
    layer1_outputs(10203) <= a and not b;
    layer1_outputs(10204) <= a and not b;
    layer1_outputs(10205) <= not (a and b);
    layer1_outputs(10206) <= a and b;
    layer1_outputs(10207) <= b;
    layer1_outputs(10208) <= not (a and b);
    layer1_outputs(10209) <= a or b;
    layer1_outputs(10210) <= b and not a;
    layer1_outputs(10211) <= a and b;
    layer1_outputs(10212) <= not b or a;
    layer1_outputs(10213) <= not (a or b);
    layer1_outputs(10214) <= not (a or b);
    layer1_outputs(10215) <= not b;
    layer1_outputs(10216) <= a and not b;
    layer1_outputs(10217) <= not a or b;
    layer1_outputs(10218) <= not (a xor b);
    layer1_outputs(10219) <= not b or a;
    layer1_outputs(10220) <= a and not b;
    layer1_outputs(10221) <= not (a and b);
    layer1_outputs(10222) <= not b;
    layer1_outputs(10223) <= a and b;
    layer1_outputs(10224) <= a or b;
    layer1_outputs(10225) <= not (a and b);
    layer1_outputs(10226) <= not b or a;
    layer1_outputs(10227) <= a or b;
    layer1_outputs(10228) <= '0';
    layer1_outputs(10229) <= '1';
    layer1_outputs(10230) <= not (a xor b);
    layer1_outputs(10231) <= not (a xor b);
    layer1_outputs(10232) <= not b;
    layer1_outputs(10233) <= not (a xor b);
    layer1_outputs(10234) <= b;
    layer1_outputs(10235) <= a and not b;
    layer1_outputs(10236) <= not a or b;
    layer1_outputs(10237) <= not a;
    layer1_outputs(10238) <= a and b;
    layer1_outputs(10239) <= not (a xor b);
    layer2_outputs(0) <= not b;
    layer2_outputs(1) <= not (a xor b);
    layer2_outputs(2) <= not a or b;
    layer2_outputs(3) <= a;
    layer2_outputs(4) <= b and not a;
    layer2_outputs(5) <= not (a xor b);
    layer2_outputs(6) <= a or b;
    layer2_outputs(7) <= not (a xor b);
    layer2_outputs(8) <= b;
    layer2_outputs(9) <= a;
    layer2_outputs(10) <= not (a xor b);
    layer2_outputs(11) <= b and not a;
    layer2_outputs(12) <= a;
    layer2_outputs(13) <= not a;
    layer2_outputs(14) <= not (a or b);
    layer2_outputs(15) <= not a;
    layer2_outputs(16) <= not b or a;
    layer2_outputs(17) <= not (a or b);
    layer2_outputs(18) <= not a or b;
    layer2_outputs(19) <= not (a and b);
    layer2_outputs(20) <= not a;
    layer2_outputs(21) <= not a;
    layer2_outputs(22) <= not b;
    layer2_outputs(23) <= not b;
    layer2_outputs(24) <= not (a xor b);
    layer2_outputs(25) <= not b;
    layer2_outputs(26) <= a;
    layer2_outputs(27) <= a and not b;
    layer2_outputs(28) <= a and not b;
    layer2_outputs(29) <= not (a and b);
    layer2_outputs(30) <= a;
    layer2_outputs(31) <= not a;
    layer2_outputs(32) <= b;
    layer2_outputs(33) <= not a;
    layer2_outputs(34) <= a;
    layer2_outputs(35) <= b and not a;
    layer2_outputs(36) <= a;
    layer2_outputs(37) <= b;
    layer2_outputs(38) <= not a;
    layer2_outputs(39) <= a;
    layer2_outputs(40) <= a and not b;
    layer2_outputs(41) <= not a;
    layer2_outputs(42) <= not b;
    layer2_outputs(43) <= not b;
    layer2_outputs(44) <= '0';
    layer2_outputs(45) <= not (a xor b);
    layer2_outputs(46) <= b;
    layer2_outputs(47) <= not a;
    layer2_outputs(48) <= a xor b;
    layer2_outputs(49) <= b;
    layer2_outputs(50) <= a and not b;
    layer2_outputs(51) <= b;
    layer2_outputs(52) <= b and not a;
    layer2_outputs(53) <= a;
    layer2_outputs(54) <= not a;
    layer2_outputs(55) <= not (a xor b);
    layer2_outputs(56) <= not (a or b);
    layer2_outputs(57) <= a;
    layer2_outputs(58) <= b;
    layer2_outputs(59) <= a xor b;
    layer2_outputs(60) <= b and not a;
    layer2_outputs(61) <= b;
    layer2_outputs(62) <= b;
    layer2_outputs(63) <= not (a xor b);
    layer2_outputs(64) <= a and not b;
    layer2_outputs(65) <= b and not a;
    layer2_outputs(66) <= a;
    layer2_outputs(67) <= b;
    layer2_outputs(68) <= a xor b;
    layer2_outputs(69) <= not a;
    layer2_outputs(70) <= not b or a;
    layer2_outputs(71) <= b;
    layer2_outputs(72) <= not (a or b);
    layer2_outputs(73) <= a or b;
    layer2_outputs(74) <= a;
    layer2_outputs(75) <= not a or b;
    layer2_outputs(76) <= '1';
    layer2_outputs(77) <= b and not a;
    layer2_outputs(78) <= not (a xor b);
    layer2_outputs(79) <= not a;
    layer2_outputs(80) <= a;
    layer2_outputs(81) <= not (a or b);
    layer2_outputs(82) <= a xor b;
    layer2_outputs(83) <= b;
    layer2_outputs(84) <= a xor b;
    layer2_outputs(85) <= not (a or b);
    layer2_outputs(86) <= a or b;
    layer2_outputs(87) <= a and b;
    layer2_outputs(88) <= a or b;
    layer2_outputs(89) <= a or b;
    layer2_outputs(90) <= a and not b;
    layer2_outputs(91) <= not b;
    layer2_outputs(92) <= b;
    layer2_outputs(93) <= a xor b;
    layer2_outputs(94) <= not (a and b);
    layer2_outputs(95) <= not b;
    layer2_outputs(96) <= b;
    layer2_outputs(97) <= not (a or b);
    layer2_outputs(98) <= not b or a;
    layer2_outputs(99) <= not a;
    layer2_outputs(100) <= a xor b;
    layer2_outputs(101) <= a xor b;
    layer2_outputs(102) <= b and not a;
    layer2_outputs(103) <= not a;
    layer2_outputs(104) <= a xor b;
    layer2_outputs(105) <= a and b;
    layer2_outputs(106) <= a and not b;
    layer2_outputs(107) <= a or b;
    layer2_outputs(108) <= not b or a;
    layer2_outputs(109) <= a xor b;
    layer2_outputs(110) <= not (a or b);
    layer2_outputs(111) <= not (a or b);
    layer2_outputs(112) <= a and b;
    layer2_outputs(113) <= a;
    layer2_outputs(114) <= not b or a;
    layer2_outputs(115) <= a or b;
    layer2_outputs(116) <= not b or a;
    layer2_outputs(117) <= not a or b;
    layer2_outputs(118) <= not b;
    layer2_outputs(119) <= not a;
    layer2_outputs(120) <= not (a and b);
    layer2_outputs(121) <= a and b;
    layer2_outputs(122) <= b;
    layer2_outputs(123) <= not a;
    layer2_outputs(124) <= b;
    layer2_outputs(125) <= not (a xor b);
    layer2_outputs(126) <= a;
    layer2_outputs(127) <= not (a and b);
    layer2_outputs(128) <= not (a and b);
    layer2_outputs(129) <= not (a xor b);
    layer2_outputs(130) <= not b;
    layer2_outputs(131) <= not (a xor b);
    layer2_outputs(132) <= b and not a;
    layer2_outputs(133) <= not (a xor b);
    layer2_outputs(134) <= b;
    layer2_outputs(135) <= not a;
    layer2_outputs(136) <= not b;
    layer2_outputs(137) <= not (a or b);
    layer2_outputs(138) <= not a;
    layer2_outputs(139) <= a xor b;
    layer2_outputs(140) <= a xor b;
    layer2_outputs(141) <= a and not b;
    layer2_outputs(142) <= not a;
    layer2_outputs(143) <= not a;
    layer2_outputs(144) <= not (a or b);
    layer2_outputs(145) <= b;
    layer2_outputs(146) <= a and not b;
    layer2_outputs(147) <= a and not b;
    layer2_outputs(148) <= a xor b;
    layer2_outputs(149) <= b;
    layer2_outputs(150) <= not (a or b);
    layer2_outputs(151) <= not a;
    layer2_outputs(152) <= a;
    layer2_outputs(153) <= not b;
    layer2_outputs(154) <= b;
    layer2_outputs(155) <= not b;
    layer2_outputs(156) <= a;
    layer2_outputs(157) <= a;
    layer2_outputs(158) <= not b;
    layer2_outputs(159) <= a xor b;
    layer2_outputs(160) <= b;
    layer2_outputs(161) <= not (a or b);
    layer2_outputs(162) <= not (a xor b);
    layer2_outputs(163) <= a and not b;
    layer2_outputs(164) <= not b or a;
    layer2_outputs(165) <= b and not a;
    layer2_outputs(166) <= a;
    layer2_outputs(167) <= not b or a;
    layer2_outputs(168) <= a xor b;
    layer2_outputs(169) <= not (a xor b);
    layer2_outputs(170) <= b;
    layer2_outputs(171) <= a or b;
    layer2_outputs(172) <= a and not b;
    layer2_outputs(173) <= not b;
    layer2_outputs(174) <= a;
    layer2_outputs(175) <= not b or a;
    layer2_outputs(176) <= not b or a;
    layer2_outputs(177) <= a xor b;
    layer2_outputs(178) <= not (a and b);
    layer2_outputs(179) <= b;
    layer2_outputs(180) <= a and b;
    layer2_outputs(181) <= b and not a;
    layer2_outputs(182) <= not b or a;
    layer2_outputs(183) <= a;
    layer2_outputs(184) <= a or b;
    layer2_outputs(185) <= '0';
    layer2_outputs(186) <= a or b;
    layer2_outputs(187) <= a and not b;
    layer2_outputs(188) <= a xor b;
    layer2_outputs(189) <= not (a xor b);
    layer2_outputs(190) <= a;
    layer2_outputs(191) <= a;
    layer2_outputs(192) <= a xor b;
    layer2_outputs(193) <= not b or a;
    layer2_outputs(194) <= not (a xor b);
    layer2_outputs(195) <= not b;
    layer2_outputs(196) <= not a;
    layer2_outputs(197) <= not (a and b);
    layer2_outputs(198) <= b and not a;
    layer2_outputs(199) <= b;
    layer2_outputs(200) <= a xor b;
    layer2_outputs(201) <= not b or a;
    layer2_outputs(202) <= a xor b;
    layer2_outputs(203) <= a;
    layer2_outputs(204) <= not a;
    layer2_outputs(205) <= not (a and b);
    layer2_outputs(206) <= not (a xor b);
    layer2_outputs(207) <= not (a and b);
    layer2_outputs(208) <= a xor b;
    layer2_outputs(209) <= not (a or b);
    layer2_outputs(210) <= a or b;
    layer2_outputs(211) <= not (a and b);
    layer2_outputs(212) <= a xor b;
    layer2_outputs(213) <= not b;
    layer2_outputs(214) <= a or b;
    layer2_outputs(215) <= not b;
    layer2_outputs(216) <= not (a xor b);
    layer2_outputs(217) <= not b or a;
    layer2_outputs(218) <= a or b;
    layer2_outputs(219) <= a and not b;
    layer2_outputs(220) <= a xor b;
    layer2_outputs(221) <= a and b;
    layer2_outputs(222) <= not b or a;
    layer2_outputs(223) <= b;
    layer2_outputs(224) <= not b or a;
    layer2_outputs(225) <= b and not a;
    layer2_outputs(226) <= a and b;
    layer2_outputs(227) <= a;
    layer2_outputs(228) <= a;
    layer2_outputs(229) <= not (a or b);
    layer2_outputs(230) <= '1';
    layer2_outputs(231) <= b;
    layer2_outputs(232) <= not a;
    layer2_outputs(233) <= a xor b;
    layer2_outputs(234) <= b;
    layer2_outputs(235) <= not b or a;
    layer2_outputs(236) <= not a;
    layer2_outputs(237) <= not b;
    layer2_outputs(238) <= not a;
    layer2_outputs(239) <= not (a xor b);
    layer2_outputs(240) <= a or b;
    layer2_outputs(241) <= a xor b;
    layer2_outputs(242) <= not a or b;
    layer2_outputs(243) <= not a or b;
    layer2_outputs(244) <= not (a xor b);
    layer2_outputs(245) <= not b;
    layer2_outputs(246) <= not a or b;
    layer2_outputs(247) <= a or b;
    layer2_outputs(248) <= not a or b;
    layer2_outputs(249) <= not b;
    layer2_outputs(250) <= a and not b;
    layer2_outputs(251) <= not a;
    layer2_outputs(252) <= a;
    layer2_outputs(253) <= not (a or b);
    layer2_outputs(254) <= not (a and b);
    layer2_outputs(255) <= not a;
    layer2_outputs(256) <= not (a xor b);
    layer2_outputs(257) <= a or b;
    layer2_outputs(258) <= b and not a;
    layer2_outputs(259) <= not a or b;
    layer2_outputs(260) <= b and not a;
    layer2_outputs(261) <= not (a xor b);
    layer2_outputs(262) <= a;
    layer2_outputs(263) <= a or b;
    layer2_outputs(264) <= not b;
    layer2_outputs(265) <= not (a or b);
    layer2_outputs(266) <= a;
    layer2_outputs(267) <= a xor b;
    layer2_outputs(268) <= not b;
    layer2_outputs(269) <= a;
    layer2_outputs(270) <= not b;
    layer2_outputs(271) <= a xor b;
    layer2_outputs(272) <= a xor b;
    layer2_outputs(273) <= not b;
    layer2_outputs(274) <= a and not b;
    layer2_outputs(275) <= not a or b;
    layer2_outputs(276) <= not a;
    layer2_outputs(277) <= not b or a;
    layer2_outputs(278) <= not (a xor b);
    layer2_outputs(279) <= a;
    layer2_outputs(280) <= not b;
    layer2_outputs(281) <= not (a xor b);
    layer2_outputs(282) <= not (a or b);
    layer2_outputs(283) <= not (a and b);
    layer2_outputs(284) <= a or b;
    layer2_outputs(285) <= not b or a;
    layer2_outputs(286) <= not (a or b);
    layer2_outputs(287) <= a;
    layer2_outputs(288) <= b;
    layer2_outputs(289) <= b;
    layer2_outputs(290) <= not a;
    layer2_outputs(291) <= not (a and b);
    layer2_outputs(292) <= b;
    layer2_outputs(293) <= not (a xor b);
    layer2_outputs(294) <= not b;
    layer2_outputs(295) <= not (a xor b);
    layer2_outputs(296) <= not (a and b);
    layer2_outputs(297) <= a xor b;
    layer2_outputs(298) <= b;
    layer2_outputs(299) <= not a or b;
    layer2_outputs(300) <= not a;
    layer2_outputs(301) <= a or b;
    layer2_outputs(302) <= a and not b;
    layer2_outputs(303) <= b;
    layer2_outputs(304) <= b;
    layer2_outputs(305) <= a;
    layer2_outputs(306) <= a xor b;
    layer2_outputs(307) <= not b or a;
    layer2_outputs(308) <= b;
    layer2_outputs(309) <= b;
    layer2_outputs(310) <= not a;
    layer2_outputs(311) <= b and not a;
    layer2_outputs(312) <= b;
    layer2_outputs(313) <= not (a and b);
    layer2_outputs(314) <= a;
    layer2_outputs(315) <= a;
    layer2_outputs(316) <= not (a and b);
    layer2_outputs(317) <= not (a xor b);
    layer2_outputs(318) <= b;
    layer2_outputs(319) <= not (a xor b);
    layer2_outputs(320) <= not (a xor b);
    layer2_outputs(321) <= b;
    layer2_outputs(322) <= b;
    layer2_outputs(323) <= not b;
    layer2_outputs(324) <= a;
    layer2_outputs(325) <= not (a and b);
    layer2_outputs(326) <= not a;
    layer2_outputs(327) <= a;
    layer2_outputs(328) <= not b;
    layer2_outputs(329) <= a;
    layer2_outputs(330) <= not b;
    layer2_outputs(331) <= b and not a;
    layer2_outputs(332) <= a;
    layer2_outputs(333) <= b;
    layer2_outputs(334) <= not (a or b);
    layer2_outputs(335) <= not b;
    layer2_outputs(336) <= not a;
    layer2_outputs(337) <= not (a xor b);
    layer2_outputs(338) <= a or b;
    layer2_outputs(339) <= not (a or b);
    layer2_outputs(340) <= a or b;
    layer2_outputs(341) <= not (a or b);
    layer2_outputs(342) <= b and not a;
    layer2_outputs(343) <= not b;
    layer2_outputs(344) <= not b or a;
    layer2_outputs(345) <= a xor b;
    layer2_outputs(346) <= not a or b;
    layer2_outputs(347) <= not (a xor b);
    layer2_outputs(348) <= a xor b;
    layer2_outputs(349) <= b;
    layer2_outputs(350) <= not a;
    layer2_outputs(351) <= b;
    layer2_outputs(352) <= a xor b;
    layer2_outputs(353) <= not (a xor b);
    layer2_outputs(354) <= a and not b;
    layer2_outputs(355) <= not b;
    layer2_outputs(356) <= a and b;
    layer2_outputs(357) <= a xor b;
    layer2_outputs(358) <= not b or a;
    layer2_outputs(359) <= b;
    layer2_outputs(360) <= not (a xor b);
    layer2_outputs(361) <= not b;
    layer2_outputs(362) <= not a;
    layer2_outputs(363) <= a;
    layer2_outputs(364) <= not (a xor b);
    layer2_outputs(365) <= not (a xor b);
    layer2_outputs(366) <= a;
    layer2_outputs(367) <= not (a xor b);
    layer2_outputs(368) <= a xor b;
    layer2_outputs(369) <= a;
    layer2_outputs(370) <= not a or b;
    layer2_outputs(371) <= not (a and b);
    layer2_outputs(372) <= not a or b;
    layer2_outputs(373) <= not (a xor b);
    layer2_outputs(374) <= a;
    layer2_outputs(375) <= b;
    layer2_outputs(376) <= b;
    layer2_outputs(377) <= b;
    layer2_outputs(378) <= a and not b;
    layer2_outputs(379) <= not (a or b);
    layer2_outputs(380) <= not (a xor b);
    layer2_outputs(381) <= not a or b;
    layer2_outputs(382) <= b and not a;
    layer2_outputs(383) <= not b;
    layer2_outputs(384) <= not b or a;
    layer2_outputs(385) <= not b;
    layer2_outputs(386) <= not (a xor b);
    layer2_outputs(387) <= not (a or b);
    layer2_outputs(388) <= a xor b;
    layer2_outputs(389) <= a;
    layer2_outputs(390) <= not b;
    layer2_outputs(391) <= not (a or b);
    layer2_outputs(392) <= not a or b;
    layer2_outputs(393) <= not b or a;
    layer2_outputs(394) <= a and not b;
    layer2_outputs(395) <= not (a xor b);
    layer2_outputs(396) <= not b or a;
    layer2_outputs(397) <= not (a xor b);
    layer2_outputs(398) <= not (a and b);
    layer2_outputs(399) <= a and not b;
    layer2_outputs(400) <= a xor b;
    layer2_outputs(401) <= not (a or b);
    layer2_outputs(402) <= a xor b;
    layer2_outputs(403) <= b;
    layer2_outputs(404) <= a xor b;
    layer2_outputs(405) <= b;
    layer2_outputs(406) <= a or b;
    layer2_outputs(407) <= not a;
    layer2_outputs(408) <= not b;
    layer2_outputs(409) <= not a or b;
    layer2_outputs(410) <= not (a or b);
    layer2_outputs(411) <= a and not b;
    layer2_outputs(412) <= not b;
    layer2_outputs(413) <= a xor b;
    layer2_outputs(414) <= not a;
    layer2_outputs(415) <= a xor b;
    layer2_outputs(416) <= b and not a;
    layer2_outputs(417) <= a and not b;
    layer2_outputs(418) <= a and b;
    layer2_outputs(419) <= a and not b;
    layer2_outputs(420) <= a;
    layer2_outputs(421) <= b;
    layer2_outputs(422) <= b;
    layer2_outputs(423) <= not b or a;
    layer2_outputs(424) <= not a or b;
    layer2_outputs(425) <= b;
    layer2_outputs(426) <= a or b;
    layer2_outputs(427) <= a;
    layer2_outputs(428) <= not b;
    layer2_outputs(429) <= not b or a;
    layer2_outputs(430) <= not (a or b);
    layer2_outputs(431) <= not b or a;
    layer2_outputs(432) <= not (a xor b);
    layer2_outputs(433) <= not (a xor b);
    layer2_outputs(434) <= not a or b;
    layer2_outputs(435) <= a;
    layer2_outputs(436) <= not a or b;
    layer2_outputs(437) <= b;
    layer2_outputs(438) <= b and not a;
    layer2_outputs(439) <= a and b;
    layer2_outputs(440) <= not b or a;
    layer2_outputs(441) <= a or b;
    layer2_outputs(442) <= not (a xor b);
    layer2_outputs(443) <= not b or a;
    layer2_outputs(444) <= not (a xor b);
    layer2_outputs(445) <= b and not a;
    layer2_outputs(446) <= a and not b;
    layer2_outputs(447) <= a;
    layer2_outputs(448) <= not b;
    layer2_outputs(449) <= a;
    layer2_outputs(450) <= not a;
    layer2_outputs(451) <= a or b;
    layer2_outputs(452) <= a xor b;
    layer2_outputs(453) <= a and not b;
    layer2_outputs(454) <= a and b;
    layer2_outputs(455) <= a;
    layer2_outputs(456) <= a and not b;
    layer2_outputs(457) <= not b;
    layer2_outputs(458) <= not (a xor b);
    layer2_outputs(459) <= not (a and b);
    layer2_outputs(460) <= a and not b;
    layer2_outputs(461) <= b;
    layer2_outputs(462) <= a or b;
    layer2_outputs(463) <= not b;
    layer2_outputs(464) <= b;
    layer2_outputs(465) <= not (a or b);
    layer2_outputs(466) <= not b;
    layer2_outputs(467) <= not b;
    layer2_outputs(468) <= b;
    layer2_outputs(469) <= a;
    layer2_outputs(470) <= a xor b;
    layer2_outputs(471) <= b and not a;
    layer2_outputs(472) <= not a;
    layer2_outputs(473) <= not (a xor b);
    layer2_outputs(474) <= b;
    layer2_outputs(475) <= not b;
    layer2_outputs(476) <= b;
    layer2_outputs(477) <= not b;
    layer2_outputs(478) <= b and not a;
    layer2_outputs(479) <= not (a xor b);
    layer2_outputs(480) <= not (a and b);
    layer2_outputs(481) <= b;
    layer2_outputs(482) <= a and b;
    layer2_outputs(483) <= not (a and b);
    layer2_outputs(484) <= b;
    layer2_outputs(485) <= b;
    layer2_outputs(486) <= a and not b;
    layer2_outputs(487) <= not (a xor b);
    layer2_outputs(488) <= not b;
    layer2_outputs(489) <= b;
    layer2_outputs(490) <= not (a and b);
    layer2_outputs(491) <= not (a or b);
    layer2_outputs(492) <= not a;
    layer2_outputs(493) <= a xor b;
    layer2_outputs(494) <= not a;
    layer2_outputs(495) <= a;
    layer2_outputs(496) <= not (a and b);
    layer2_outputs(497) <= not a or b;
    layer2_outputs(498) <= not (a and b);
    layer2_outputs(499) <= b;
    layer2_outputs(500) <= not a or b;
    layer2_outputs(501) <= not (a and b);
    layer2_outputs(502) <= a or b;
    layer2_outputs(503) <= a;
    layer2_outputs(504) <= not b or a;
    layer2_outputs(505) <= a and not b;
    layer2_outputs(506) <= not (a and b);
    layer2_outputs(507) <= b;
    layer2_outputs(508) <= a xor b;
    layer2_outputs(509) <= not (a and b);
    layer2_outputs(510) <= a and b;
    layer2_outputs(511) <= not a or b;
    layer2_outputs(512) <= a;
    layer2_outputs(513) <= not (a and b);
    layer2_outputs(514) <= a or b;
    layer2_outputs(515) <= a xor b;
    layer2_outputs(516) <= not a;
    layer2_outputs(517) <= not (a xor b);
    layer2_outputs(518) <= a and b;
    layer2_outputs(519) <= not (a and b);
    layer2_outputs(520) <= a and not b;
    layer2_outputs(521) <= a xor b;
    layer2_outputs(522) <= b;
    layer2_outputs(523) <= b;
    layer2_outputs(524) <= not b;
    layer2_outputs(525) <= a;
    layer2_outputs(526) <= not b;
    layer2_outputs(527) <= a and not b;
    layer2_outputs(528) <= not (a or b);
    layer2_outputs(529) <= a and b;
    layer2_outputs(530) <= not a;
    layer2_outputs(531) <= a and b;
    layer2_outputs(532) <= not (a xor b);
    layer2_outputs(533) <= b and not a;
    layer2_outputs(534) <= a and not b;
    layer2_outputs(535) <= b and not a;
    layer2_outputs(536) <= a or b;
    layer2_outputs(537) <= a and not b;
    layer2_outputs(538) <= not b;
    layer2_outputs(539) <= b;
    layer2_outputs(540) <= not (a xor b);
    layer2_outputs(541) <= a;
    layer2_outputs(542) <= a and b;
    layer2_outputs(543) <= a;
    layer2_outputs(544) <= not (a and b);
    layer2_outputs(545) <= not (a xor b);
    layer2_outputs(546) <= a and not b;
    layer2_outputs(547) <= not a;
    layer2_outputs(548) <= b;
    layer2_outputs(549) <= b;
    layer2_outputs(550) <= a;
    layer2_outputs(551) <= not b;
    layer2_outputs(552) <= a and b;
    layer2_outputs(553) <= not b;
    layer2_outputs(554) <= b;
    layer2_outputs(555) <= b;
    layer2_outputs(556) <= a xor b;
    layer2_outputs(557) <= not a or b;
    layer2_outputs(558) <= '1';
    layer2_outputs(559) <= not b or a;
    layer2_outputs(560) <= a and not b;
    layer2_outputs(561) <= b and not a;
    layer2_outputs(562) <= not (a xor b);
    layer2_outputs(563) <= a and b;
    layer2_outputs(564) <= not (a xor b);
    layer2_outputs(565) <= not (a xor b);
    layer2_outputs(566) <= not b;
    layer2_outputs(567) <= not b or a;
    layer2_outputs(568) <= b and not a;
    layer2_outputs(569) <= a xor b;
    layer2_outputs(570) <= a or b;
    layer2_outputs(571) <= not (a or b);
    layer2_outputs(572) <= b;
    layer2_outputs(573) <= not (a xor b);
    layer2_outputs(574) <= a and b;
    layer2_outputs(575) <= not a;
    layer2_outputs(576) <= not b;
    layer2_outputs(577) <= not b;
    layer2_outputs(578) <= a xor b;
    layer2_outputs(579) <= a and not b;
    layer2_outputs(580) <= not a or b;
    layer2_outputs(581) <= not (a xor b);
    layer2_outputs(582) <= a;
    layer2_outputs(583) <= not b or a;
    layer2_outputs(584) <= not a;
    layer2_outputs(585) <= a or b;
    layer2_outputs(586) <= not a or b;
    layer2_outputs(587) <= not a;
    layer2_outputs(588) <= not (a and b);
    layer2_outputs(589) <= a and not b;
    layer2_outputs(590) <= b and not a;
    layer2_outputs(591) <= not a;
    layer2_outputs(592) <= not b;
    layer2_outputs(593) <= b;
    layer2_outputs(594) <= a xor b;
    layer2_outputs(595) <= b;
    layer2_outputs(596) <= b;
    layer2_outputs(597) <= not b or a;
    layer2_outputs(598) <= b;
    layer2_outputs(599) <= not (a xor b);
    layer2_outputs(600) <= a and b;
    layer2_outputs(601) <= a xor b;
    layer2_outputs(602) <= b;
    layer2_outputs(603) <= a;
    layer2_outputs(604) <= b;
    layer2_outputs(605) <= a xor b;
    layer2_outputs(606) <= not a;
    layer2_outputs(607) <= not a;
    layer2_outputs(608) <= a;
    layer2_outputs(609) <= not (a xor b);
    layer2_outputs(610) <= not (a and b);
    layer2_outputs(611) <= a xor b;
    layer2_outputs(612) <= a xor b;
    layer2_outputs(613) <= not (a or b);
    layer2_outputs(614) <= not a;
    layer2_outputs(615) <= not (a or b);
    layer2_outputs(616) <= a xor b;
    layer2_outputs(617) <= not b;
    layer2_outputs(618) <= not (a and b);
    layer2_outputs(619) <= b;
    layer2_outputs(620) <= b;
    layer2_outputs(621) <= not (a and b);
    layer2_outputs(622) <= a or b;
    layer2_outputs(623) <= a and b;
    layer2_outputs(624) <= not (a xor b);
    layer2_outputs(625) <= not a;
    layer2_outputs(626) <= a and b;
    layer2_outputs(627) <= b;
    layer2_outputs(628) <= a;
    layer2_outputs(629) <= not (a and b);
    layer2_outputs(630) <= not (a xor b);
    layer2_outputs(631) <= not (a and b);
    layer2_outputs(632) <= a xor b;
    layer2_outputs(633) <= a;
    layer2_outputs(634) <= a;
    layer2_outputs(635) <= not b;
    layer2_outputs(636) <= b;
    layer2_outputs(637) <= not a or b;
    layer2_outputs(638) <= a xor b;
    layer2_outputs(639) <= not a or b;
    layer2_outputs(640) <= not a;
    layer2_outputs(641) <= not (a and b);
    layer2_outputs(642) <= not a;
    layer2_outputs(643) <= not (a or b);
    layer2_outputs(644) <= not a or b;
    layer2_outputs(645) <= not b or a;
    layer2_outputs(646) <= a and not b;
    layer2_outputs(647) <= not b;
    layer2_outputs(648) <= b;
    layer2_outputs(649) <= a and b;
    layer2_outputs(650) <= a xor b;
    layer2_outputs(651) <= b;
    layer2_outputs(652) <= not b or a;
    layer2_outputs(653) <= b;
    layer2_outputs(654) <= not a or b;
    layer2_outputs(655) <= a or b;
    layer2_outputs(656) <= b;
    layer2_outputs(657) <= not b;
    layer2_outputs(658) <= not (a and b);
    layer2_outputs(659) <= b;
    layer2_outputs(660) <= not b;
    layer2_outputs(661) <= not (a or b);
    layer2_outputs(662) <= a or b;
    layer2_outputs(663) <= not a or b;
    layer2_outputs(664) <= not b;
    layer2_outputs(665) <= b;
    layer2_outputs(666) <= b and not a;
    layer2_outputs(667) <= b and not a;
    layer2_outputs(668) <= not (a or b);
    layer2_outputs(669) <= b;
    layer2_outputs(670) <= a and not b;
    layer2_outputs(671) <= b and not a;
    layer2_outputs(672) <= not (a and b);
    layer2_outputs(673) <= b and not a;
    layer2_outputs(674) <= not (a xor b);
    layer2_outputs(675) <= not a or b;
    layer2_outputs(676) <= not b or a;
    layer2_outputs(677) <= not (a and b);
    layer2_outputs(678) <= not (a and b);
    layer2_outputs(679) <= b and not a;
    layer2_outputs(680) <= not b;
    layer2_outputs(681) <= not b or a;
    layer2_outputs(682) <= b;
    layer2_outputs(683) <= b;
    layer2_outputs(684) <= not (a or b);
    layer2_outputs(685) <= a and b;
    layer2_outputs(686) <= not b or a;
    layer2_outputs(687) <= a and b;
    layer2_outputs(688) <= a and b;
    layer2_outputs(689) <= a and not b;
    layer2_outputs(690) <= b and not a;
    layer2_outputs(691) <= not (a xor b);
    layer2_outputs(692) <= b and not a;
    layer2_outputs(693) <= a xor b;
    layer2_outputs(694) <= not b;
    layer2_outputs(695) <= b;
    layer2_outputs(696) <= not a or b;
    layer2_outputs(697) <= not b or a;
    layer2_outputs(698) <= not b;
    layer2_outputs(699) <= not a;
    layer2_outputs(700) <= a or b;
    layer2_outputs(701) <= not (a xor b);
    layer2_outputs(702) <= a and not b;
    layer2_outputs(703) <= not (a xor b);
    layer2_outputs(704) <= not b or a;
    layer2_outputs(705) <= not a or b;
    layer2_outputs(706) <= a xor b;
    layer2_outputs(707) <= a xor b;
    layer2_outputs(708) <= not b or a;
    layer2_outputs(709) <= not a;
    layer2_outputs(710) <= not (a xor b);
    layer2_outputs(711) <= not (a xor b);
    layer2_outputs(712) <= not b;
    layer2_outputs(713) <= not b;
    layer2_outputs(714) <= a or b;
    layer2_outputs(715) <= not (a xor b);
    layer2_outputs(716) <= a and b;
    layer2_outputs(717) <= not (a xor b);
    layer2_outputs(718) <= '1';
    layer2_outputs(719) <= a xor b;
    layer2_outputs(720) <= not a or b;
    layer2_outputs(721) <= not a;
    layer2_outputs(722) <= b and not a;
    layer2_outputs(723) <= a xor b;
    layer2_outputs(724) <= not b or a;
    layer2_outputs(725) <= not b;
    layer2_outputs(726) <= not b;
    layer2_outputs(727) <= not b;
    layer2_outputs(728) <= b and not a;
    layer2_outputs(729) <= b;
    layer2_outputs(730) <= not (a or b);
    layer2_outputs(731) <= a xor b;
    layer2_outputs(732) <= not a;
    layer2_outputs(733) <= not b;
    layer2_outputs(734) <= a xor b;
    layer2_outputs(735) <= not (a and b);
    layer2_outputs(736) <= a and not b;
    layer2_outputs(737) <= a;
    layer2_outputs(738) <= not a;
    layer2_outputs(739) <= not b;
    layer2_outputs(740) <= a;
    layer2_outputs(741) <= not (a xor b);
    layer2_outputs(742) <= not a or b;
    layer2_outputs(743) <= not (a xor b);
    layer2_outputs(744) <= not a;
    layer2_outputs(745) <= b and not a;
    layer2_outputs(746) <= not (a xor b);
    layer2_outputs(747) <= a;
    layer2_outputs(748) <= a xor b;
    layer2_outputs(749) <= not a;
    layer2_outputs(750) <= not (a and b);
    layer2_outputs(751) <= not (a and b);
    layer2_outputs(752) <= not a or b;
    layer2_outputs(753) <= not b;
    layer2_outputs(754) <= b;
    layer2_outputs(755) <= not a or b;
    layer2_outputs(756) <= not a or b;
    layer2_outputs(757) <= a xor b;
    layer2_outputs(758) <= not (a xor b);
    layer2_outputs(759) <= a and b;
    layer2_outputs(760) <= not (a or b);
    layer2_outputs(761) <= not (a or b);
    layer2_outputs(762) <= a or b;
    layer2_outputs(763) <= a or b;
    layer2_outputs(764) <= a and not b;
    layer2_outputs(765) <= a;
    layer2_outputs(766) <= a;
    layer2_outputs(767) <= not (a and b);
    layer2_outputs(768) <= a xor b;
    layer2_outputs(769) <= not a;
    layer2_outputs(770) <= a;
    layer2_outputs(771) <= not a;
    layer2_outputs(772) <= not b or a;
    layer2_outputs(773) <= not b;
    layer2_outputs(774) <= not (a xor b);
    layer2_outputs(775) <= not b or a;
    layer2_outputs(776) <= b and not a;
    layer2_outputs(777) <= a;
    layer2_outputs(778) <= b;
    layer2_outputs(779) <= a or b;
    layer2_outputs(780) <= a and b;
    layer2_outputs(781) <= not (a xor b);
    layer2_outputs(782) <= a xor b;
    layer2_outputs(783) <= a and not b;
    layer2_outputs(784) <= not a;
    layer2_outputs(785) <= not (a xor b);
    layer2_outputs(786) <= a;
    layer2_outputs(787) <= a;
    layer2_outputs(788) <= not b;
    layer2_outputs(789) <= b and not a;
    layer2_outputs(790) <= not (a or b);
    layer2_outputs(791) <= a;
    layer2_outputs(792) <= not (a and b);
    layer2_outputs(793) <= not a or b;
    layer2_outputs(794) <= a;
    layer2_outputs(795) <= not b or a;
    layer2_outputs(796) <= not (a xor b);
    layer2_outputs(797) <= not (a or b);
    layer2_outputs(798) <= a xor b;
    layer2_outputs(799) <= not a;
    layer2_outputs(800) <= a and b;
    layer2_outputs(801) <= not b or a;
    layer2_outputs(802) <= not b;
    layer2_outputs(803) <= a and b;
    layer2_outputs(804) <= not a;
    layer2_outputs(805) <= a xor b;
    layer2_outputs(806) <= not a or b;
    layer2_outputs(807) <= a xor b;
    layer2_outputs(808) <= not a;
    layer2_outputs(809) <= not b or a;
    layer2_outputs(810) <= a;
    layer2_outputs(811) <= '0';
    layer2_outputs(812) <= not (a xor b);
    layer2_outputs(813) <= not b or a;
    layer2_outputs(814) <= a;
    layer2_outputs(815) <= not b or a;
    layer2_outputs(816) <= not a;
    layer2_outputs(817) <= not b;
    layer2_outputs(818) <= not a;
    layer2_outputs(819) <= a and not b;
    layer2_outputs(820) <= a or b;
    layer2_outputs(821) <= a and b;
    layer2_outputs(822) <= b and not a;
    layer2_outputs(823) <= a or b;
    layer2_outputs(824) <= not (a and b);
    layer2_outputs(825) <= not b;
    layer2_outputs(826) <= b and not a;
    layer2_outputs(827) <= not (a and b);
    layer2_outputs(828) <= b;
    layer2_outputs(829) <= b;
    layer2_outputs(830) <= not a or b;
    layer2_outputs(831) <= a;
    layer2_outputs(832) <= a or b;
    layer2_outputs(833) <= b and not a;
    layer2_outputs(834) <= a or b;
    layer2_outputs(835) <= not a;
    layer2_outputs(836) <= b;
    layer2_outputs(837) <= not a;
    layer2_outputs(838) <= a xor b;
    layer2_outputs(839) <= not (a xor b);
    layer2_outputs(840) <= not a;
    layer2_outputs(841) <= a;
    layer2_outputs(842) <= not a;
    layer2_outputs(843) <= not a;
    layer2_outputs(844) <= a and not b;
    layer2_outputs(845) <= not (a or b);
    layer2_outputs(846) <= a;
    layer2_outputs(847) <= not b;
    layer2_outputs(848) <= b;
    layer2_outputs(849) <= not a or b;
    layer2_outputs(850) <= a xor b;
    layer2_outputs(851) <= a xor b;
    layer2_outputs(852) <= a;
    layer2_outputs(853) <= not a;
    layer2_outputs(854) <= a xor b;
    layer2_outputs(855) <= not a;
    layer2_outputs(856) <= a and not b;
    layer2_outputs(857) <= a and not b;
    layer2_outputs(858) <= a and b;
    layer2_outputs(859) <= not b;
    layer2_outputs(860) <= a and b;
    layer2_outputs(861) <= not b;
    layer2_outputs(862) <= b;
    layer2_outputs(863) <= a xor b;
    layer2_outputs(864) <= not (a xor b);
    layer2_outputs(865) <= b;
    layer2_outputs(866) <= a;
    layer2_outputs(867) <= not (a and b);
    layer2_outputs(868) <= not (a xor b);
    layer2_outputs(869) <= not a or b;
    layer2_outputs(870) <= not b;
    layer2_outputs(871) <= a or b;
    layer2_outputs(872) <= not (a or b);
    layer2_outputs(873) <= not (a and b);
    layer2_outputs(874) <= a;
    layer2_outputs(875) <= b;
    layer2_outputs(876) <= a;
    layer2_outputs(877) <= a and b;
    layer2_outputs(878) <= not a or b;
    layer2_outputs(879) <= a and b;
    layer2_outputs(880) <= b;
    layer2_outputs(881) <= a xor b;
    layer2_outputs(882) <= not b or a;
    layer2_outputs(883) <= not (a xor b);
    layer2_outputs(884) <= b and not a;
    layer2_outputs(885) <= not b or a;
    layer2_outputs(886) <= a and not b;
    layer2_outputs(887) <= not (a or b);
    layer2_outputs(888) <= a;
    layer2_outputs(889) <= a;
    layer2_outputs(890) <= a or b;
    layer2_outputs(891) <= not b;
    layer2_outputs(892) <= not b;
    layer2_outputs(893) <= not a or b;
    layer2_outputs(894) <= '1';
    layer2_outputs(895) <= not b;
    layer2_outputs(896) <= b;
    layer2_outputs(897) <= not b;
    layer2_outputs(898) <= b and not a;
    layer2_outputs(899) <= a;
    layer2_outputs(900) <= not b or a;
    layer2_outputs(901) <= not b or a;
    layer2_outputs(902) <= b;
    layer2_outputs(903) <= not b;
    layer2_outputs(904) <= b;
    layer2_outputs(905) <= a or b;
    layer2_outputs(906) <= not (a xor b);
    layer2_outputs(907) <= a and b;
    layer2_outputs(908) <= not a or b;
    layer2_outputs(909) <= a;
    layer2_outputs(910) <= b;
    layer2_outputs(911) <= not (a xor b);
    layer2_outputs(912) <= a;
    layer2_outputs(913) <= a xor b;
    layer2_outputs(914) <= not (a xor b);
    layer2_outputs(915) <= not (a xor b);
    layer2_outputs(916) <= a;
    layer2_outputs(917) <= b;
    layer2_outputs(918) <= not a or b;
    layer2_outputs(919) <= a xor b;
    layer2_outputs(920) <= not (a xor b);
    layer2_outputs(921) <= not b;
    layer2_outputs(922) <= not (a or b);
    layer2_outputs(923) <= a and not b;
    layer2_outputs(924) <= a and b;
    layer2_outputs(925) <= not b or a;
    layer2_outputs(926) <= b;
    layer2_outputs(927) <= not (a xor b);
    layer2_outputs(928) <= a and not b;
    layer2_outputs(929) <= a xor b;
    layer2_outputs(930) <= a and b;
    layer2_outputs(931) <= not (a or b);
    layer2_outputs(932) <= a;
    layer2_outputs(933) <= not a;
    layer2_outputs(934) <= not a;
    layer2_outputs(935) <= a;
    layer2_outputs(936) <= a;
    layer2_outputs(937) <= b and not a;
    layer2_outputs(938) <= a and b;
    layer2_outputs(939) <= b and not a;
    layer2_outputs(940) <= a;
    layer2_outputs(941) <= a and b;
    layer2_outputs(942) <= a and b;
    layer2_outputs(943) <= b;
    layer2_outputs(944) <= not a;
    layer2_outputs(945) <= not (a or b);
    layer2_outputs(946) <= not (a xor b);
    layer2_outputs(947) <= b and not a;
    layer2_outputs(948) <= '1';
    layer2_outputs(949) <= not b or a;
    layer2_outputs(950) <= not b;
    layer2_outputs(951) <= not a;
    layer2_outputs(952) <= not b;
    layer2_outputs(953) <= a;
    layer2_outputs(954) <= b;
    layer2_outputs(955) <= a xor b;
    layer2_outputs(956) <= not a;
    layer2_outputs(957) <= not (a and b);
    layer2_outputs(958) <= b;
    layer2_outputs(959) <= a and b;
    layer2_outputs(960) <= not b or a;
    layer2_outputs(961) <= not (a or b);
    layer2_outputs(962) <= not (a or b);
    layer2_outputs(963) <= a and b;
    layer2_outputs(964) <= not (a xor b);
    layer2_outputs(965) <= a xor b;
    layer2_outputs(966) <= a and not b;
    layer2_outputs(967) <= a xor b;
    layer2_outputs(968) <= not a;
    layer2_outputs(969) <= a xor b;
    layer2_outputs(970) <= not a;
    layer2_outputs(971) <= a or b;
    layer2_outputs(972) <= not b;
    layer2_outputs(973) <= not a;
    layer2_outputs(974) <= not a;
    layer2_outputs(975) <= b;
    layer2_outputs(976) <= a and not b;
    layer2_outputs(977) <= not (a xor b);
    layer2_outputs(978) <= not b;
    layer2_outputs(979) <= b and not a;
    layer2_outputs(980) <= not (a and b);
    layer2_outputs(981) <= a xor b;
    layer2_outputs(982) <= not b or a;
    layer2_outputs(983) <= a;
    layer2_outputs(984) <= a or b;
    layer2_outputs(985) <= not (a or b);
    layer2_outputs(986) <= not b or a;
    layer2_outputs(987) <= '1';
    layer2_outputs(988) <= not a or b;
    layer2_outputs(989) <= b and not a;
    layer2_outputs(990) <= b;
    layer2_outputs(991) <= not a;
    layer2_outputs(992) <= a and not b;
    layer2_outputs(993) <= not (a or b);
    layer2_outputs(994) <= not (a or b);
    layer2_outputs(995) <= b and not a;
    layer2_outputs(996) <= b;
    layer2_outputs(997) <= not b or a;
    layer2_outputs(998) <= a or b;
    layer2_outputs(999) <= a;
    layer2_outputs(1000) <= not (a and b);
    layer2_outputs(1001) <= a and b;
    layer2_outputs(1002) <= '0';
    layer2_outputs(1003) <= a and not b;
    layer2_outputs(1004) <= not a;
    layer2_outputs(1005) <= not b;
    layer2_outputs(1006) <= b and not a;
    layer2_outputs(1007) <= not (a and b);
    layer2_outputs(1008) <= b and not a;
    layer2_outputs(1009) <= '1';
    layer2_outputs(1010) <= a xor b;
    layer2_outputs(1011) <= b;
    layer2_outputs(1012) <= a xor b;
    layer2_outputs(1013) <= b;
    layer2_outputs(1014) <= b;
    layer2_outputs(1015) <= not (a or b);
    layer2_outputs(1016) <= not a;
    layer2_outputs(1017) <= not b;
    layer2_outputs(1018) <= a;
    layer2_outputs(1019) <= not a;
    layer2_outputs(1020) <= a xor b;
    layer2_outputs(1021) <= a or b;
    layer2_outputs(1022) <= not a or b;
    layer2_outputs(1023) <= not b;
    layer2_outputs(1024) <= b;
    layer2_outputs(1025) <= a and not b;
    layer2_outputs(1026) <= a xor b;
    layer2_outputs(1027) <= a;
    layer2_outputs(1028) <= not b;
    layer2_outputs(1029) <= a xor b;
    layer2_outputs(1030) <= not (a and b);
    layer2_outputs(1031) <= a xor b;
    layer2_outputs(1032) <= not (a or b);
    layer2_outputs(1033) <= b and not a;
    layer2_outputs(1034) <= b;
    layer2_outputs(1035) <= b;
    layer2_outputs(1036) <= a;
    layer2_outputs(1037) <= not (a or b);
    layer2_outputs(1038) <= not (a and b);
    layer2_outputs(1039) <= a;
    layer2_outputs(1040) <= not (a or b);
    layer2_outputs(1041) <= not a;
    layer2_outputs(1042) <= a xor b;
    layer2_outputs(1043) <= a or b;
    layer2_outputs(1044) <= not (a or b);
    layer2_outputs(1045) <= not a;
    layer2_outputs(1046) <= b;
    layer2_outputs(1047) <= not (a and b);
    layer2_outputs(1048) <= a;
    layer2_outputs(1049) <= not b;
    layer2_outputs(1050) <= a;
    layer2_outputs(1051) <= not (a and b);
    layer2_outputs(1052) <= a and b;
    layer2_outputs(1053) <= a and not b;
    layer2_outputs(1054) <= a and b;
    layer2_outputs(1055) <= a and not b;
    layer2_outputs(1056) <= a and not b;
    layer2_outputs(1057) <= a and not b;
    layer2_outputs(1058) <= not (a xor b);
    layer2_outputs(1059) <= not (a xor b);
    layer2_outputs(1060) <= b;
    layer2_outputs(1061) <= not b or a;
    layer2_outputs(1062) <= b;
    layer2_outputs(1063) <= not (a xor b);
    layer2_outputs(1064) <= not a;
    layer2_outputs(1065) <= a and not b;
    layer2_outputs(1066) <= not a;
    layer2_outputs(1067) <= a and not b;
    layer2_outputs(1068) <= b;
    layer2_outputs(1069) <= a and b;
    layer2_outputs(1070) <= a xor b;
    layer2_outputs(1071) <= not (a xor b);
    layer2_outputs(1072) <= not b or a;
    layer2_outputs(1073) <= a or b;
    layer2_outputs(1074) <= not (a and b);
    layer2_outputs(1075) <= b;
    layer2_outputs(1076) <= not a;
    layer2_outputs(1077) <= not (a and b);
    layer2_outputs(1078) <= not (a or b);
    layer2_outputs(1079) <= not a or b;
    layer2_outputs(1080) <= not b;
    layer2_outputs(1081) <= a or b;
    layer2_outputs(1082) <= b and not a;
    layer2_outputs(1083) <= not (a xor b);
    layer2_outputs(1084) <= not (a and b);
    layer2_outputs(1085) <= a and not b;
    layer2_outputs(1086) <= a;
    layer2_outputs(1087) <= not a;
    layer2_outputs(1088) <= a xor b;
    layer2_outputs(1089) <= not b;
    layer2_outputs(1090) <= not (a and b);
    layer2_outputs(1091) <= not (a or b);
    layer2_outputs(1092) <= a;
    layer2_outputs(1093) <= b;
    layer2_outputs(1094) <= not a;
    layer2_outputs(1095) <= a and b;
    layer2_outputs(1096) <= not a;
    layer2_outputs(1097) <= a or b;
    layer2_outputs(1098) <= a;
    layer2_outputs(1099) <= not b;
    layer2_outputs(1100) <= not b or a;
    layer2_outputs(1101) <= a and b;
    layer2_outputs(1102) <= not b;
    layer2_outputs(1103) <= a and b;
    layer2_outputs(1104) <= not (a and b);
    layer2_outputs(1105) <= b;
    layer2_outputs(1106) <= not a;
    layer2_outputs(1107) <= a xor b;
    layer2_outputs(1108) <= not a;
    layer2_outputs(1109) <= a and not b;
    layer2_outputs(1110) <= a;
    layer2_outputs(1111) <= b;
    layer2_outputs(1112) <= b and not a;
    layer2_outputs(1113) <= not a or b;
    layer2_outputs(1114) <= not b;
    layer2_outputs(1115) <= a and b;
    layer2_outputs(1116) <= a;
    layer2_outputs(1117) <= a;
    layer2_outputs(1118) <= not a or b;
    layer2_outputs(1119) <= not a or b;
    layer2_outputs(1120) <= a xor b;
    layer2_outputs(1121) <= a and not b;
    layer2_outputs(1122) <= not (a and b);
    layer2_outputs(1123) <= a or b;
    layer2_outputs(1124) <= a and b;
    layer2_outputs(1125) <= not b;
    layer2_outputs(1126) <= b and not a;
    layer2_outputs(1127) <= a;
    layer2_outputs(1128) <= b;
    layer2_outputs(1129) <= a or b;
    layer2_outputs(1130) <= a and not b;
    layer2_outputs(1131) <= not a or b;
    layer2_outputs(1132) <= not (a and b);
    layer2_outputs(1133) <= not b;
    layer2_outputs(1134) <= a xor b;
    layer2_outputs(1135) <= not (a or b);
    layer2_outputs(1136) <= not (a xor b);
    layer2_outputs(1137) <= not b or a;
    layer2_outputs(1138) <= a xor b;
    layer2_outputs(1139) <= a;
    layer2_outputs(1140) <= not b;
    layer2_outputs(1141) <= not (a or b);
    layer2_outputs(1142) <= not (a or b);
    layer2_outputs(1143) <= not (a xor b);
    layer2_outputs(1144) <= a;
    layer2_outputs(1145) <= not b;
    layer2_outputs(1146) <= not a;
    layer2_outputs(1147) <= a and not b;
    layer2_outputs(1148) <= not b or a;
    layer2_outputs(1149) <= a and b;
    layer2_outputs(1150) <= a xor b;
    layer2_outputs(1151) <= not a or b;
    layer2_outputs(1152) <= not (a xor b);
    layer2_outputs(1153) <= a or b;
    layer2_outputs(1154) <= not (a xor b);
    layer2_outputs(1155) <= a xor b;
    layer2_outputs(1156) <= not (a and b);
    layer2_outputs(1157) <= a and not b;
    layer2_outputs(1158) <= a and not b;
    layer2_outputs(1159) <= not a;
    layer2_outputs(1160) <= a;
    layer2_outputs(1161) <= b;
    layer2_outputs(1162) <= a and b;
    layer2_outputs(1163) <= not (a xor b);
    layer2_outputs(1164) <= not a;
    layer2_outputs(1165) <= not (a or b);
    layer2_outputs(1166) <= b;
    layer2_outputs(1167) <= a and not b;
    layer2_outputs(1168) <= a and b;
    layer2_outputs(1169) <= a;
    layer2_outputs(1170) <= a;
    layer2_outputs(1171) <= not b;
    layer2_outputs(1172) <= not a or b;
    layer2_outputs(1173) <= a;
    layer2_outputs(1174) <= a and not b;
    layer2_outputs(1175) <= a;
    layer2_outputs(1176) <= a;
    layer2_outputs(1177) <= not a;
    layer2_outputs(1178) <= not a or b;
    layer2_outputs(1179) <= a and not b;
    layer2_outputs(1180) <= a xor b;
    layer2_outputs(1181) <= not a;
    layer2_outputs(1182) <= b;
    layer2_outputs(1183) <= a and not b;
    layer2_outputs(1184) <= not (a and b);
    layer2_outputs(1185) <= a and b;
    layer2_outputs(1186) <= a;
    layer2_outputs(1187) <= not b;
    layer2_outputs(1188) <= b and not a;
    layer2_outputs(1189) <= b;
    layer2_outputs(1190) <= not (a or b);
    layer2_outputs(1191) <= a;
    layer2_outputs(1192) <= not b or a;
    layer2_outputs(1193) <= b and not a;
    layer2_outputs(1194) <= a xor b;
    layer2_outputs(1195) <= a xor b;
    layer2_outputs(1196) <= a or b;
    layer2_outputs(1197) <= not (a xor b);
    layer2_outputs(1198) <= a and not b;
    layer2_outputs(1199) <= not b;
    layer2_outputs(1200) <= not (a and b);
    layer2_outputs(1201) <= not a or b;
    layer2_outputs(1202) <= a xor b;
    layer2_outputs(1203) <= a or b;
    layer2_outputs(1204) <= b;
    layer2_outputs(1205) <= a xor b;
    layer2_outputs(1206) <= not (a xor b);
    layer2_outputs(1207) <= not (a xor b);
    layer2_outputs(1208) <= not a;
    layer2_outputs(1209) <= not a;
    layer2_outputs(1210) <= a xor b;
    layer2_outputs(1211) <= a xor b;
    layer2_outputs(1212) <= a xor b;
    layer2_outputs(1213) <= b;
    layer2_outputs(1214) <= not b;
    layer2_outputs(1215) <= not a;
    layer2_outputs(1216) <= not a;
    layer2_outputs(1217) <= b;
    layer2_outputs(1218) <= a xor b;
    layer2_outputs(1219) <= a;
    layer2_outputs(1220) <= b and not a;
    layer2_outputs(1221) <= b;
    layer2_outputs(1222) <= a or b;
    layer2_outputs(1223) <= not (a and b);
    layer2_outputs(1224) <= not b;
    layer2_outputs(1225) <= not a;
    layer2_outputs(1226) <= not (a xor b);
    layer2_outputs(1227) <= not a or b;
    layer2_outputs(1228) <= a or b;
    layer2_outputs(1229) <= b and not a;
    layer2_outputs(1230) <= b;
    layer2_outputs(1231) <= not a;
    layer2_outputs(1232) <= a;
    layer2_outputs(1233) <= not a;
    layer2_outputs(1234) <= a xor b;
    layer2_outputs(1235) <= b and not a;
    layer2_outputs(1236) <= not b;
    layer2_outputs(1237) <= b;
    layer2_outputs(1238) <= not (a or b);
    layer2_outputs(1239) <= not (a xor b);
    layer2_outputs(1240) <= not a or b;
    layer2_outputs(1241) <= not (a or b);
    layer2_outputs(1242) <= a and b;
    layer2_outputs(1243) <= not (a xor b);
    layer2_outputs(1244) <= b;
    layer2_outputs(1245) <= b and not a;
    layer2_outputs(1246) <= not (a and b);
    layer2_outputs(1247) <= b and not a;
    layer2_outputs(1248) <= not a;
    layer2_outputs(1249) <= a;
    layer2_outputs(1250) <= not a or b;
    layer2_outputs(1251) <= a;
    layer2_outputs(1252) <= a;
    layer2_outputs(1253) <= a or b;
    layer2_outputs(1254) <= not b;
    layer2_outputs(1255) <= a and not b;
    layer2_outputs(1256) <= not b or a;
    layer2_outputs(1257) <= a;
    layer2_outputs(1258) <= not a;
    layer2_outputs(1259) <= a xor b;
    layer2_outputs(1260) <= not b;
    layer2_outputs(1261) <= not (a or b);
    layer2_outputs(1262) <= a;
    layer2_outputs(1263) <= a or b;
    layer2_outputs(1264) <= a or b;
    layer2_outputs(1265) <= not a;
    layer2_outputs(1266) <= a;
    layer2_outputs(1267) <= a;
    layer2_outputs(1268) <= not a;
    layer2_outputs(1269) <= b and not a;
    layer2_outputs(1270) <= not b;
    layer2_outputs(1271) <= not a;
    layer2_outputs(1272) <= b;
    layer2_outputs(1273) <= a;
    layer2_outputs(1274) <= b and not a;
    layer2_outputs(1275) <= not a;
    layer2_outputs(1276) <= a and b;
    layer2_outputs(1277) <= a or b;
    layer2_outputs(1278) <= a;
    layer2_outputs(1279) <= not (a and b);
    layer2_outputs(1280) <= not a;
    layer2_outputs(1281) <= a and b;
    layer2_outputs(1282) <= not a;
    layer2_outputs(1283) <= a xor b;
    layer2_outputs(1284) <= not b;
    layer2_outputs(1285) <= not b;
    layer2_outputs(1286) <= not (a or b);
    layer2_outputs(1287) <= a xor b;
    layer2_outputs(1288) <= a;
    layer2_outputs(1289) <= b;
    layer2_outputs(1290) <= a and b;
    layer2_outputs(1291) <= not a;
    layer2_outputs(1292) <= not a or b;
    layer2_outputs(1293) <= b;
    layer2_outputs(1294) <= a xor b;
    layer2_outputs(1295) <= a or b;
    layer2_outputs(1296) <= not a;
    layer2_outputs(1297) <= b;
    layer2_outputs(1298) <= not a;
    layer2_outputs(1299) <= a xor b;
    layer2_outputs(1300) <= a;
    layer2_outputs(1301) <= a xor b;
    layer2_outputs(1302) <= b and not a;
    layer2_outputs(1303) <= not a;
    layer2_outputs(1304) <= a xor b;
    layer2_outputs(1305) <= not b or a;
    layer2_outputs(1306) <= not a or b;
    layer2_outputs(1307) <= a;
    layer2_outputs(1308) <= b;
    layer2_outputs(1309) <= not (a xor b);
    layer2_outputs(1310) <= not a;
    layer2_outputs(1311) <= not b;
    layer2_outputs(1312) <= a xor b;
    layer2_outputs(1313) <= a;
    layer2_outputs(1314) <= a xor b;
    layer2_outputs(1315) <= not a;
    layer2_outputs(1316) <= b;
    layer2_outputs(1317) <= a;
    layer2_outputs(1318) <= not b;
    layer2_outputs(1319) <= not (a and b);
    layer2_outputs(1320) <= a and b;
    layer2_outputs(1321) <= a xor b;
    layer2_outputs(1322) <= a and not b;
    layer2_outputs(1323) <= a xor b;
    layer2_outputs(1324) <= a;
    layer2_outputs(1325) <= not b;
    layer2_outputs(1326) <= not a;
    layer2_outputs(1327) <= b and not a;
    layer2_outputs(1328) <= not (a xor b);
    layer2_outputs(1329) <= b;
    layer2_outputs(1330) <= a xor b;
    layer2_outputs(1331) <= not (a xor b);
    layer2_outputs(1332) <= a and not b;
    layer2_outputs(1333) <= a xor b;
    layer2_outputs(1334) <= b and not a;
    layer2_outputs(1335) <= not b;
    layer2_outputs(1336) <= not b;
    layer2_outputs(1337) <= not b;
    layer2_outputs(1338) <= a and not b;
    layer2_outputs(1339) <= a and b;
    layer2_outputs(1340) <= b;
    layer2_outputs(1341) <= '0';
    layer2_outputs(1342) <= not b;
    layer2_outputs(1343) <= not a;
    layer2_outputs(1344) <= not b;
    layer2_outputs(1345) <= a;
    layer2_outputs(1346) <= not b;
    layer2_outputs(1347) <= not b;
    layer2_outputs(1348) <= b and not a;
    layer2_outputs(1349) <= not (a or b);
    layer2_outputs(1350) <= not b or a;
    layer2_outputs(1351) <= a or b;
    layer2_outputs(1352) <= a and not b;
    layer2_outputs(1353) <= a or b;
    layer2_outputs(1354) <= a;
    layer2_outputs(1355) <= not b;
    layer2_outputs(1356) <= a and b;
    layer2_outputs(1357) <= not a;
    layer2_outputs(1358) <= a and b;
    layer2_outputs(1359) <= a and b;
    layer2_outputs(1360) <= not (a xor b);
    layer2_outputs(1361) <= a;
    layer2_outputs(1362) <= b;
    layer2_outputs(1363) <= a and not b;
    layer2_outputs(1364) <= b and not a;
    layer2_outputs(1365) <= a xor b;
    layer2_outputs(1366) <= a;
    layer2_outputs(1367) <= not (a and b);
    layer2_outputs(1368) <= a;
    layer2_outputs(1369) <= not a or b;
    layer2_outputs(1370) <= not (a xor b);
    layer2_outputs(1371) <= not b;
    layer2_outputs(1372) <= a and b;
    layer2_outputs(1373) <= a;
    layer2_outputs(1374) <= not b;
    layer2_outputs(1375) <= a and not b;
    layer2_outputs(1376) <= not a;
    layer2_outputs(1377) <= b;
    layer2_outputs(1378) <= b;
    layer2_outputs(1379) <= not (a xor b);
    layer2_outputs(1380) <= not b or a;
    layer2_outputs(1381) <= not (a xor b);
    layer2_outputs(1382) <= a;
    layer2_outputs(1383) <= not (a xor b);
    layer2_outputs(1384) <= a xor b;
    layer2_outputs(1385) <= not (a xor b);
    layer2_outputs(1386) <= a xor b;
    layer2_outputs(1387) <= b and not a;
    layer2_outputs(1388) <= not b;
    layer2_outputs(1389) <= not (a xor b);
    layer2_outputs(1390) <= not b or a;
    layer2_outputs(1391) <= a xor b;
    layer2_outputs(1392) <= not (a xor b);
    layer2_outputs(1393) <= not a;
    layer2_outputs(1394) <= not b or a;
    layer2_outputs(1395) <= not a;
    layer2_outputs(1396) <= not a or b;
    layer2_outputs(1397) <= not (a xor b);
    layer2_outputs(1398) <= b and not a;
    layer2_outputs(1399) <= not b or a;
    layer2_outputs(1400) <= not (a and b);
    layer2_outputs(1401) <= not (a xor b);
    layer2_outputs(1402) <= not b or a;
    layer2_outputs(1403) <= not b;
    layer2_outputs(1404) <= not a or b;
    layer2_outputs(1405) <= not a;
    layer2_outputs(1406) <= not a;
    layer2_outputs(1407) <= not b or a;
    layer2_outputs(1408) <= b;
    layer2_outputs(1409) <= a and not b;
    layer2_outputs(1410) <= b;
    layer2_outputs(1411) <= a and b;
    layer2_outputs(1412) <= a and b;
    layer2_outputs(1413) <= not (a xor b);
    layer2_outputs(1414) <= not a or b;
    layer2_outputs(1415) <= b and not a;
    layer2_outputs(1416) <= not a;
    layer2_outputs(1417) <= b;
    layer2_outputs(1418) <= not b or a;
    layer2_outputs(1419) <= a xor b;
    layer2_outputs(1420) <= a xor b;
    layer2_outputs(1421) <= b;
    layer2_outputs(1422) <= a xor b;
    layer2_outputs(1423) <= not b;
    layer2_outputs(1424) <= not a;
    layer2_outputs(1425) <= a;
    layer2_outputs(1426) <= not a;
    layer2_outputs(1427) <= a;
    layer2_outputs(1428) <= a and not b;
    layer2_outputs(1429) <= a or b;
    layer2_outputs(1430) <= not (a xor b);
    layer2_outputs(1431) <= a;
    layer2_outputs(1432) <= not (a xor b);
    layer2_outputs(1433) <= not b or a;
    layer2_outputs(1434) <= b and not a;
    layer2_outputs(1435) <= a or b;
    layer2_outputs(1436) <= a;
    layer2_outputs(1437) <= a and b;
    layer2_outputs(1438) <= a;
    layer2_outputs(1439) <= not (a and b);
    layer2_outputs(1440) <= not (a xor b);
    layer2_outputs(1441) <= not b;
    layer2_outputs(1442) <= a xor b;
    layer2_outputs(1443) <= a xor b;
    layer2_outputs(1444) <= b and not a;
    layer2_outputs(1445) <= not b;
    layer2_outputs(1446) <= not (a and b);
    layer2_outputs(1447) <= not (a and b);
    layer2_outputs(1448) <= a or b;
    layer2_outputs(1449) <= not (a and b);
    layer2_outputs(1450) <= not (a and b);
    layer2_outputs(1451) <= not (a and b);
    layer2_outputs(1452) <= b;
    layer2_outputs(1453) <= not (a or b);
    layer2_outputs(1454) <= b;
    layer2_outputs(1455) <= a or b;
    layer2_outputs(1456) <= a;
    layer2_outputs(1457) <= not a;
    layer2_outputs(1458) <= not (a or b);
    layer2_outputs(1459) <= b and not a;
    layer2_outputs(1460) <= not b;
    layer2_outputs(1461) <= not b;
    layer2_outputs(1462) <= not b;
    layer2_outputs(1463) <= not a;
    layer2_outputs(1464) <= not a or b;
    layer2_outputs(1465) <= a;
    layer2_outputs(1466) <= not a or b;
    layer2_outputs(1467) <= not (a xor b);
    layer2_outputs(1468) <= not a or b;
    layer2_outputs(1469) <= not b or a;
    layer2_outputs(1470) <= not b;
    layer2_outputs(1471) <= a xor b;
    layer2_outputs(1472) <= a xor b;
    layer2_outputs(1473) <= a or b;
    layer2_outputs(1474) <= not b;
    layer2_outputs(1475) <= not b;
    layer2_outputs(1476) <= a and not b;
    layer2_outputs(1477) <= a xor b;
    layer2_outputs(1478) <= a;
    layer2_outputs(1479) <= not a;
    layer2_outputs(1480) <= a and not b;
    layer2_outputs(1481) <= a xor b;
    layer2_outputs(1482) <= a and b;
    layer2_outputs(1483) <= not b;
    layer2_outputs(1484) <= not b or a;
    layer2_outputs(1485) <= b;
    layer2_outputs(1486) <= not (a or b);
    layer2_outputs(1487) <= not a or b;
    layer2_outputs(1488) <= not (a and b);
    layer2_outputs(1489) <= a and b;
    layer2_outputs(1490) <= a and not b;
    layer2_outputs(1491) <= b and not a;
    layer2_outputs(1492) <= not (a xor b);
    layer2_outputs(1493) <= not b;
    layer2_outputs(1494) <= not a;
    layer2_outputs(1495) <= not (a and b);
    layer2_outputs(1496) <= not (a xor b);
    layer2_outputs(1497) <= a xor b;
    layer2_outputs(1498) <= not b or a;
    layer2_outputs(1499) <= a;
    layer2_outputs(1500) <= b;
    layer2_outputs(1501) <= not a or b;
    layer2_outputs(1502) <= not (a and b);
    layer2_outputs(1503) <= b;
    layer2_outputs(1504) <= not (a xor b);
    layer2_outputs(1505) <= a xor b;
    layer2_outputs(1506) <= not (a or b);
    layer2_outputs(1507) <= b;
    layer2_outputs(1508) <= a;
    layer2_outputs(1509) <= a;
    layer2_outputs(1510) <= not b;
    layer2_outputs(1511) <= not b;
    layer2_outputs(1512) <= not a;
    layer2_outputs(1513) <= b;
    layer2_outputs(1514) <= not b or a;
    layer2_outputs(1515) <= b;
    layer2_outputs(1516) <= not (a xor b);
    layer2_outputs(1517) <= a and b;
    layer2_outputs(1518) <= a;
    layer2_outputs(1519) <= a or b;
    layer2_outputs(1520) <= a xor b;
    layer2_outputs(1521) <= a;
    layer2_outputs(1522) <= a and b;
    layer2_outputs(1523) <= '0';
    layer2_outputs(1524) <= not (a xor b);
    layer2_outputs(1525) <= not (a xor b);
    layer2_outputs(1526) <= a xor b;
    layer2_outputs(1527) <= b and not a;
    layer2_outputs(1528) <= not a or b;
    layer2_outputs(1529) <= not (a xor b);
    layer2_outputs(1530) <= a xor b;
    layer2_outputs(1531) <= a xor b;
    layer2_outputs(1532) <= a;
    layer2_outputs(1533) <= '0';
    layer2_outputs(1534) <= b;
    layer2_outputs(1535) <= not (a and b);
    layer2_outputs(1536) <= a or b;
    layer2_outputs(1537) <= not (a xor b);
    layer2_outputs(1538) <= not (a and b);
    layer2_outputs(1539) <= a xor b;
    layer2_outputs(1540) <= a and b;
    layer2_outputs(1541) <= b;
    layer2_outputs(1542) <= not a;
    layer2_outputs(1543) <= a;
    layer2_outputs(1544) <= not (a xor b);
    layer2_outputs(1545) <= a xor b;
    layer2_outputs(1546) <= not b;
    layer2_outputs(1547) <= not a;
    layer2_outputs(1548) <= a or b;
    layer2_outputs(1549) <= not b;
    layer2_outputs(1550) <= not (a and b);
    layer2_outputs(1551) <= a xor b;
    layer2_outputs(1552) <= a xor b;
    layer2_outputs(1553) <= a and b;
    layer2_outputs(1554) <= a xor b;
    layer2_outputs(1555) <= not (a or b);
    layer2_outputs(1556) <= a;
    layer2_outputs(1557) <= a or b;
    layer2_outputs(1558) <= not b;
    layer2_outputs(1559) <= not (a or b);
    layer2_outputs(1560) <= b;
    layer2_outputs(1561) <= not (a or b);
    layer2_outputs(1562) <= a;
    layer2_outputs(1563) <= a or b;
    layer2_outputs(1564) <= a;
    layer2_outputs(1565) <= a xor b;
    layer2_outputs(1566) <= a or b;
    layer2_outputs(1567) <= not a;
    layer2_outputs(1568) <= a;
    layer2_outputs(1569) <= a xor b;
    layer2_outputs(1570) <= a and not b;
    layer2_outputs(1571) <= not b;
    layer2_outputs(1572) <= a;
    layer2_outputs(1573) <= not (a xor b);
    layer2_outputs(1574) <= a xor b;
    layer2_outputs(1575) <= not a;
    layer2_outputs(1576) <= not a or b;
    layer2_outputs(1577) <= b and not a;
    layer2_outputs(1578) <= a and b;
    layer2_outputs(1579) <= a and b;
    layer2_outputs(1580) <= not a;
    layer2_outputs(1581) <= not a;
    layer2_outputs(1582) <= a or b;
    layer2_outputs(1583) <= not a or b;
    layer2_outputs(1584) <= a xor b;
    layer2_outputs(1585) <= b and not a;
    layer2_outputs(1586) <= not b or a;
    layer2_outputs(1587) <= not a or b;
    layer2_outputs(1588) <= a xor b;
    layer2_outputs(1589) <= not a;
    layer2_outputs(1590) <= b;
    layer2_outputs(1591) <= a and b;
    layer2_outputs(1592) <= a;
    layer2_outputs(1593) <= b and not a;
    layer2_outputs(1594) <= not a;
    layer2_outputs(1595) <= b and not a;
    layer2_outputs(1596) <= not b;
    layer2_outputs(1597) <= b;
    layer2_outputs(1598) <= a xor b;
    layer2_outputs(1599) <= not (a xor b);
    layer2_outputs(1600) <= not (a xor b);
    layer2_outputs(1601) <= a and not b;
    layer2_outputs(1602) <= b;
    layer2_outputs(1603) <= not b;
    layer2_outputs(1604) <= not (a or b);
    layer2_outputs(1605) <= not a;
    layer2_outputs(1606) <= not (a xor b);
    layer2_outputs(1607) <= not a or b;
    layer2_outputs(1608) <= a and not b;
    layer2_outputs(1609) <= a;
    layer2_outputs(1610) <= a and not b;
    layer2_outputs(1611) <= '0';
    layer2_outputs(1612) <= a;
    layer2_outputs(1613) <= a and not b;
    layer2_outputs(1614) <= not b;
    layer2_outputs(1615) <= not (a or b);
    layer2_outputs(1616) <= b and not a;
    layer2_outputs(1617) <= not a;
    layer2_outputs(1618) <= not a;
    layer2_outputs(1619) <= a xor b;
    layer2_outputs(1620) <= b;
    layer2_outputs(1621) <= not a;
    layer2_outputs(1622) <= b and not a;
    layer2_outputs(1623) <= b;
    layer2_outputs(1624) <= a and b;
    layer2_outputs(1625) <= not (a or b);
    layer2_outputs(1626) <= not b;
    layer2_outputs(1627) <= a xor b;
    layer2_outputs(1628) <= b;
    layer2_outputs(1629) <= a xor b;
    layer2_outputs(1630) <= a;
    layer2_outputs(1631) <= a;
    layer2_outputs(1632) <= b and not a;
    layer2_outputs(1633) <= a and b;
    layer2_outputs(1634) <= a;
    layer2_outputs(1635) <= a xor b;
    layer2_outputs(1636) <= a;
    layer2_outputs(1637) <= b and not a;
    layer2_outputs(1638) <= a xor b;
    layer2_outputs(1639) <= b;
    layer2_outputs(1640) <= not b or a;
    layer2_outputs(1641) <= not b or a;
    layer2_outputs(1642) <= not b;
    layer2_outputs(1643) <= b;
    layer2_outputs(1644) <= a and not b;
    layer2_outputs(1645) <= not (a or b);
    layer2_outputs(1646) <= not b;
    layer2_outputs(1647) <= not a;
    layer2_outputs(1648) <= not a;
    layer2_outputs(1649) <= not (a or b);
    layer2_outputs(1650) <= not (a or b);
    layer2_outputs(1651) <= a;
    layer2_outputs(1652) <= b;
    layer2_outputs(1653) <= not b;
    layer2_outputs(1654) <= a and not b;
    layer2_outputs(1655) <= a and not b;
    layer2_outputs(1656) <= not (a or b);
    layer2_outputs(1657) <= b and not a;
    layer2_outputs(1658) <= not a;
    layer2_outputs(1659) <= not (a xor b);
    layer2_outputs(1660) <= b;
    layer2_outputs(1661) <= a;
    layer2_outputs(1662) <= not (a xor b);
    layer2_outputs(1663) <= not (a xor b);
    layer2_outputs(1664) <= a;
    layer2_outputs(1665) <= not b;
    layer2_outputs(1666) <= not a;
    layer2_outputs(1667) <= not a or b;
    layer2_outputs(1668) <= not b;
    layer2_outputs(1669) <= not (a and b);
    layer2_outputs(1670) <= not a;
    layer2_outputs(1671) <= a;
    layer2_outputs(1672) <= a and b;
    layer2_outputs(1673) <= a;
    layer2_outputs(1674) <= not b;
    layer2_outputs(1675) <= a xor b;
    layer2_outputs(1676) <= not (a and b);
    layer2_outputs(1677) <= a or b;
    layer2_outputs(1678) <= b and not a;
    layer2_outputs(1679) <= a and b;
    layer2_outputs(1680) <= not a or b;
    layer2_outputs(1681) <= not b or a;
    layer2_outputs(1682) <= not (a xor b);
    layer2_outputs(1683) <= not (a and b);
    layer2_outputs(1684) <= not (a xor b);
    layer2_outputs(1685) <= not (a and b);
    layer2_outputs(1686) <= not a;
    layer2_outputs(1687) <= a;
    layer2_outputs(1688) <= a and b;
    layer2_outputs(1689) <= not (a or b);
    layer2_outputs(1690) <= a;
    layer2_outputs(1691) <= a;
    layer2_outputs(1692) <= not a;
    layer2_outputs(1693) <= b;
    layer2_outputs(1694) <= not (a xor b);
    layer2_outputs(1695) <= not b or a;
    layer2_outputs(1696) <= a;
    layer2_outputs(1697) <= b and not a;
    layer2_outputs(1698) <= not a;
    layer2_outputs(1699) <= not (a and b);
    layer2_outputs(1700) <= not (a or b);
    layer2_outputs(1701) <= not (a xor b);
    layer2_outputs(1702) <= not (a xor b);
    layer2_outputs(1703) <= not (a xor b);
    layer2_outputs(1704) <= a;
    layer2_outputs(1705) <= not (a xor b);
    layer2_outputs(1706) <= b;
    layer2_outputs(1707) <= not b or a;
    layer2_outputs(1708) <= not a;
    layer2_outputs(1709) <= not a;
    layer2_outputs(1710) <= not (a xor b);
    layer2_outputs(1711) <= not b;
    layer2_outputs(1712) <= b and not a;
    layer2_outputs(1713) <= not b or a;
    layer2_outputs(1714) <= b and not a;
    layer2_outputs(1715) <= a xor b;
    layer2_outputs(1716) <= not (a xor b);
    layer2_outputs(1717) <= not b;
    layer2_outputs(1718) <= b;
    layer2_outputs(1719) <= '1';
    layer2_outputs(1720) <= not (a and b);
    layer2_outputs(1721) <= not (a xor b);
    layer2_outputs(1722) <= a;
    layer2_outputs(1723) <= not (a or b);
    layer2_outputs(1724) <= not b;
    layer2_outputs(1725) <= b;
    layer2_outputs(1726) <= not a or b;
    layer2_outputs(1727) <= a and not b;
    layer2_outputs(1728) <= not a;
    layer2_outputs(1729) <= a;
    layer2_outputs(1730) <= a and b;
    layer2_outputs(1731) <= a and not b;
    layer2_outputs(1732) <= not b;
    layer2_outputs(1733) <= not (a and b);
    layer2_outputs(1734) <= a;
    layer2_outputs(1735) <= '0';
    layer2_outputs(1736) <= a;
    layer2_outputs(1737) <= not (a xor b);
    layer2_outputs(1738) <= not (a xor b);
    layer2_outputs(1739) <= not b or a;
    layer2_outputs(1740) <= not (a xor b);
    layer2_outputs(1741) <= not a;
    layer2_outputs(1742) <= a xor b;
    layer2_outputs(1743) <= b;
    layer2_outputs(1744) <= not a or b;
    layer2_outputs(1745) <= not (a or b);
    layer2_outputs(1746) <= not (a xor b);
    layer2_outputs(1747) <= not b;
    layer2_outputs(1748) <= a;
    layer2_outputs(1749) <= not a;
    layer2_outputs(1750) <= a xor b;
    layer2_outputs(1751) <= not (a and b);
    layer2_outputs(1752) <= not a or b;
    layer2_outputs(1753) <= not (a or b);
    layer2_outputs(1754) <= not (a and b);
    layer2_outputs(1755) <= not (a or b);
    layer2_outputs(1756) <= not a or b;
    layer2_outputs(1757) <= a xor b;
    layer2_outputs(1758) <= not b;
    layer2_outputs(1759) <= not a;
    layer2_outputs(1760) <= a or b;
    layer2_outputs(1761) <= not b;
    layer2_outputs(1762) <= a and b;
    layer2_outputs(1763) <= not a or b;
    layer2_outputs(1764) <= not (a xor b);
    layer2_outputs(1765) <= a xor b;
    layer2_outputs(1766) <= not (a or b);
    layer2_outputs(1767) <= not (a xor b);
    layer2_outputs(1768) <= not (a xor b);
    layer2_outputs(1769) <= a;
    layer2_outputs(1770) <= a;
    layer2_outputs(1771) <= not (a or b);
    layer2_outputs(1772) <= not b;
    layer2_outputs(1773) <= b;
    layer2_outputs(1774) <= a;
    layer2_outputs(1775) <= not a;
    layer2_outputs(1776) <= b and not a;
    layer2_outputs(1777) <= not (a or b);
    layer2_outputs(1778) <= not (a xor b);
    layer2_outputs(1779) <= not (a or b);
    layer2_outputs(1780) <= not (a and b);
    layer2_outputs(1781) <= not b;
    layer2_outputs(1782) <= a xor b;
    layer2_outputs(1783) <= not b;
    layer2_outputs(1784) <= b and not a;
    layer2_outputs(1785) <= a xor b;
    layer2_outputs(1786) <= a xor b;
    layer2_outputs(1787) <= not (a or b);
    layer2_outputs(1788) <= '0';
    layer2_outputs(1789) <= '1';
    layer2_outputs(1790) <= a and b;
    layer2_outputs(1791) <= not (a xor b);
    layer2_outputs(1792) <= not (a xor b);
    layer2_outputs(1793) <= b and not a;
    layer2_outputs(1794) <= a;
    layer2_outputs(1795) <= not (a xor b);
    layer2_outputs(1796) <= a;
    layer2_outputs(1797) <= b;
    layer2_outputs(1798) <= a;
    layer2_outputs(1799) <= not (a and b);
    layer2_outputs(1800) <= a and not b;
    layer2_outputs(1801) <= not a;
    layer2_outputs(1802) <= a;
    layer2_outputs(1803) <= not a;
    layer2_outputs(1804) <= b and not a;
    layer2_outputs(1805) <= a and not b;
    layer2_outputs(1806) <= not a;
    layer2_outputs(1807) <= b;
    layer2_outputs(1808) <= b;
    layer2_outputs(1809) <= a or b;
    layer2_outputs(1810) <= b;
    layer2_outputs(1811) <= not a;
    layer2_outputs(1812) <= a xor b;
    layer2_outputs(1813) <= b and not a;
    layer2_outputs(1814) <= not (a and b);
    layer2_outputs(1815) <= a or b;
    layer2_outputs(1816) <= not b or a;
    layer2_outputs(1817) <= a or b;
    layer2_outputs(1818) <= a or b;
    layer2_outputs(1819) <= a;
    layer2_outputs(1820) <= a xor b;
    layer2_outputs(1821) <= b and not a;
    layer2_outputs(1822) <= not (a and b);
    layer2_outputs(1823) <= not (a xor b);
    layer2_outputs(1824) <= not b;
    layer2_outputs(1825) <= b;
    layer2_outputs(1826) <= a and b;
    layer2_outputs(1827) <= b and not a;
    layer2_outputs(1828) <= not a;
    layer2_outputs(1829) <= not b;
    layer2_outputs(1830) <= a and b;
    layer2_outputs(1831) <= not (a xor b);
    layer2_outputs(1832) <= not b;
    layer2_outputs(1833) <= not a;
    layer2_outputs(1834) <= a;
    layer2_outputs(1835) <= not b;
    layer2_outputs(1836) <= a and not b;
    layer2_outputs(1837) <= b;
    layer2_outputs(1838) <= not a;
    layer2_outputs(1839) <= b;
    layer2_outputs(1840) <= not a or b;
    layer2_outputs(1841) <= not b;
    layer2_outputs(1842) <= not a;
    layer2_outputs(1843) <= a xor b;
    layer2_outputs(1844) <= b;
    layer2_outputs(1845) <= a;
    layer2_outputs(1846) <= not (a xor b);
    layer2_outputs(1847) <= not (a xor b);
    layer2_outputs(1848) <= not a;
    layer2_outputs(1849) <= a and b;
    layer2_outputs(1850) <= not (a or b);
    layer2_outputs(1851) <= not (a or b);
    layer2_outputs(1852) <= b;
    layer2_outputs(1853) <= a and b;
    layer2_outputs(1854) <= a and not b;
    layer2_outputs(1855) <= not a or b;
    layer2_outputs(1856) <= not (a or b);
    layer2_outputs(1857) <= b;
    layer2_outputs(1858) <= not b;
    layer2_outputs(1859) <= not a;
    layer2_outputs(1860) <= not a or b;
    layer2_outputs(1861) <= b;
    layer2_outputs(1862) <= not b or a;
    layer2_outputs(1863) <= not b;
    layer2_outputs(1864) <= not a;
    layer2_outputs(1865) <= not b or a;
    layer2_outputs(1866) <= not a;
    layer2_outputs(1867) <= not a;
    layer2_outputs(1868) <= not b;
    layer2_outputs(1869) <= b;
    layer2_outputs(1870) <= '0';
    layer2_outputs(1871) <= not (a and b);
    layer2_outputs(1872) <= not (a xor b);
    layer2_outputs(1873) <= not (a or b);
    layer2_outputs(1874) <= b and not a;
    layer2_outputs(1875) <= not b;
    layer2_outputs(1876) <= a;
    layer2_outputs(1877) <= a;
    layer2_outputs(1878) <= not b;
    layer2_outputs(1879) <= '1';
    layer2_outputs(1880) <= not b or a;
    layer2_outputs(1881) <= not a;
    layer2_outputs(1882) <= not (a and b);
    layer2_outputs(1883) <= a xor b;
    layer2_outputs(1884) <= a xor b;
    layer2_outputs(1885) <= not (a and b);
    layer2_outputs(1886) <= not a or b;
    layer2_outputs(1887) <= not (a xor b);
    layer2_outputs(1888) <= b;
    layer2_outputs(1889) <= not (a or b);
    layer2_outputs(1890) <= b;
    layer2_outputs(1891) <= not b;
    layer2_outputs(1892) <= not b;
    layer2_outputs(1893) <= not (a and b);
    layer2_outputs(1894) <= a and b;
    layer2_outputs(1895) <= b;
    layer2_outputs(1896) <= a and b;
    layer2_outputs(1897) <= a or b;
    layer2_outputs(1898) <= a xor b;
    layer2_outputs(1899) <= b and not a;
    layer2_outputs(1900) <= a and not b;
    layer2_outputs(1901) <= not (a and b);
    layer2_outputs(1902) <= not b or a;
    layer2_outputs(1903) <= not a;
    layer2_outputs(1904) <= a;
    layer2_outputs(1905) <= not b or a;
    layer2_outputs(1906) <= not (a xor b);
    layer2_outputs(1907) <= not (a and b);
    layer2_outputs(1908) <= not b;
    layer2_outputs(1909) <= a;
    layer2_outputs(1910) <= not (a or b);
    layer2_outputs(1911) <= a xor b;
    layer2_outputs(1912) <= a or b;
    layer2_outputs(1913) <= a and not b;
    layer2_outputs(1914) <= not (a xor b);
    layer2_outputs(1915) <= not (a xor b);
    layer2_outputs(1916) <= a;
    layer2_outputs(1917) <= not (a xor b);
    layer2_outputs(1918) <= not (a xor b);
    layer2_outputs(1919) <= not a;
    layer2_outputs(1920) <= a xor b;
    layer2_outputs(1921) <= not (a xor b);
    layer2_outputs(1922) <= not a or b;
    layer2_outputs(1923) <= not (a xor b);
    layer2_outputs(1924) <= a and not b;
    layer2_outputs(1925) <= a xor b;
    layer2_outputs(1926) <= a or b;
    layer2_outputs(1927) <= b and not a;
    layer2_outputs(1928) <= not a or b;
    layer2_outputs(1929) <= not (a xor b);
    layer2_outputs(1930) <= not (a xor b);
    layer2_outputs(1931) <= not (a xor b);
    layer2_outputs(1932) <= a and b;
    layer2_outputs(1933) <= a;
    layer2_outputs(1934) <= a or b;
    layer2_outputs(1935) <= not a;
    layer2_outputs(1936) <= b;
    layer2_outputs(1937) <= a;
    layer2_outputs(1938) <= not a;
    layer2_outputs(1939) <= a;
    layer2_outputs(1940) <= a or b;
    layer2_outputs(1941) <= a xor b;
    layer2_outputs(1942) <= a xor b;
    layer2_outputs(1943) <= a xor b;
    layer2_outputs(1944) <= not a;
    layer2_outputs(1945) <= not (a xor b);
    layer2_outputs(1946) <= not b or a;
    layer2_outputs(1947) <= not b;
    layer2_outputs(1948) <= not b;
    layer2_outputs(1949) <= a;
    layer2_outputs(1950) <= a xor b;
    layer2_outputs(1951) <= not a;
    layer2_outputs(1952) <= a or b;
    layer2_outputs(1953) <= not b or a;
    layer2_outputs(1954) <= a;
    layer2_outputs(1955) <= not a;
    layer2_outputs(1956) <= a and b;
    layer2_outputs(1957) <= a and b;
    layer2_outputs(1958) <= not b;
    layer2_outputs(1959) <= not (a xor b);
    layer2_outputs(1960) <= not (a or b);
    layer2_outputs(1961) <= not a;
    layer2_outputs(1962) <= not (a xor b);
    layer2_outputs(1963) <= not b;
    layer2_outputs(1964) <= not b;
    layer2_outputs(1965) <= not a;
    layer2_outputs(1966) <= not (a xor b);
    layer2_outputs(1967) <= b;
    layer2_outputs(1968) <= not a;
    layer2_outputs(1969) <= not (a or b);
    layer2_outputs(1970) <= a and not b;
    layer2_outputs(1971) <= b and not a;
    layer2_outputs(1972) <= not (a or b);
    layer2_outputs(1973) <= a and not b;
    layer2_outputs(1974) <= not b;
    layer2_outputs(1975) <= a or b;
    layer2_outputs(1976) <= not b;
    layer2_outputs(1977) <= not (a or b);
    layer2_outputs(1978) <= not b;
    layer2_outputs(1979) <= not a;
    layer2_outputs(1980) <= not a;
    layer2_outputs(1981) <= '1';
    layer2_outputs(1982) <= not a;
    layer2_outputs(1983) <= a and not b;
    layer2_outputs(1984) <= not a;
    layer2_outputs(1985) <= not (a and b);
    layer2_outputs(1986) <= not a;
    layer2_outputs(1987) <= not (a or b);
    layer2_outputs(1988) <= not a;
    layer2_outputs(1989) <= not (a xor b);
    layer2_outputs(1990) <= b;
    layer2_outputs(1991) <= b;
    layer2_outputs(1992) <= b and not a;
    layer2_outputs(1993) <= a and b;
    layer2_outputs(1994) <= not (a and b);
    layer2_outputs(1995) <= not (a or b);
    layer2_outputs(1996) <= not (a xor b);
    layer2_outputs(1997) <= a xor b;
    layer2_outputs(1998) <= b;
    layer2_outputs(1999) <= a xor b;
    layer2_outputs(2000) <= a and b;
    layer2_outputs(2001) <= not a;
    layer2_outputs(2002) <= not b;
    layer2_outputs(2003) <= b;
    layer2_outputs(2004) <= not a;
    layer2_outputs(2005) <= not (a xor b);
    layer2_outputs(2006) <= a or b;
    layer2_outputs(2007) <= a xor b;
    layer2_outputs(2008) <= b and not a;
    layer2_outputs(2009) <= a xor b;
    layer2_outputs(2010) <= not a;
    layer2_outputs(2011) <= a xor b;
    layer2_outputs(2012) <= a;
    layer2_outputs(2013) <= b and not a;
    layer2_outputs(2014) <= a and b;
    layer2_outputs(2015) <= not a;
    layer2_outputs(2016) <= a xor b;
    layer2_outputs(2017) <= not (a xor b);
    layer2_outputs(2018) <= a xor b;
    layer2_outputs(2019) <= not (a xor b);
    layer2_outputs(2020) <= not (a xor b);
    layer2_outputs(2021) <= not (a xor b);
    layer2_outputs(2022) <= a xor b;
    layer2_outputs(2023) <= b and not a;
    layer2_outputs(2024) <= not b;
    layer2_outputs(2025) <= not b;
    layer2_outputs(2026) <= not b;
    layer2_outputs(2027) <= a;
    layer2_outputs(2028) <= b and not a;
    layer2_outputs(2029) <= not b;
    layer2_outputs(2030) <= not b;
    layer2_outputs(2031) <= not b;
    layer2_outputs(2032) <= not b or a;
    layer2_outputs(2033) <= b;
    layer2_outputs(2034) <= b;
    layer2_outputs(2035) <= not a or b;
    layer2_outputs(2036) <= not b or a;
    layer2_outputs(2037) <= not a;
    layer2_outputs(2038) <= not a or b;
    layer2_outputs(2039) <= not b;
    layer2_outputs(2040) <= a xor b;
    layer2_outputs(2041) <= a xor b;
    layer2_outputs(2042) <= a or b;
    layer2_outputs(2043) <= not (a xor b);
    layer2_outputs(2044) <= a;
    layer2_outputs(2045) <= a and b;
    layer2_outputs(2046) <= not (a xor b);
    layer2_outputs(2047) <= not (a or b);
    layer2_outputs(2048) <= b and not a;
    layer2_outputs(2049) <= not (a xor b);
    layer2_outputs(2050) <= not (a xor b);
    layer2_outputs(2051) <= b and not a;
    layer2_outputs(2052) <= not a or b;
    layer2_outputs(2053) <= b;
    layer2_outputs(2054) <= not b;
    layer2_outputs(2055) <= a or b;
    layer2_outputs(2056) <= b;
    layer2_outputs(2057) <= not a;
    layer2_outputs(2058) <= a and b;
    layer2_outputs(2059) <= '0';
    layer2_outputs(2060) <= a xor b;
    layer2_outputs(2061) <= '1';
    layer2_outputs(2062) <= not (a xor b);
    layer2_outputs(2063) <= b;
    layer2_outputs(2064) <= a and not b;
    layer2_outputs(2065) <= a;
    layer2_outputs(2066) <= not (a and b);
    layer2_outputs(2067) <= a xor b;
    layer2_outputs(2068) <= b and not a;
    layer2_outputs(2069) <= a xor b;
    layer2_outputs(2070) <= b;
    layer2_outputs(2071) <= not a;
    layer2_outputs(2072) <= not a or b;
    layer2_outputs(2073) <= '1';
    layer2_outputs(2074) <= not (a xor b);
    layer2_outputs(2075) <= not a;
    layer2_outputs(2076) <= b and not a;
    layer2_outputs(2077) <= not a;
    layer2_outputs(2078) <= a and b;
    layer2_outputs(2079) <= a and not b;
    layer2_outputs(2080) <= a;
    layer2_outputs(2081) <= a;
    layer2_outputs(2082) <= a;
    layer2_outputs(2083) <= a and b;
    layer2_outputs(2084) <= a and not b;
    layer2_outputs(2085) <= not a or b;
    layer2_outputs(2086) <= not a;
    layer2_outputs(2087) <= a;
    layer2_outputs(2088) <= a;
    layer2_outputs(2089) <= not a or b;
    layer2_outputs(2090) <= b and not a;
    layer2_outputs(2091) <= not a;
    layer2_outputs(2092) <= a;
    layer2_outputs(2093) <= a xor b;
    layer2_outputs(2094) <= b;
    layer2_outputs(2095) <= not b;
    layer2_outputs(2096) <= b;
    layer2_outputs(2097) <= not a;
    layer2_outputs(2098) <= not (a xor b);
    layer2_outputs(2099) <= a xor b;
    layer2_outputs(2100) <= not b;
    layer2_outputs(2101) <= not a or b;
    layer2_outputs(2102) <= not a or b;
    layer2_outputs(2103) <= not a;
    layer2_outputs(2104) <= a;
    layer2_outputs(2105) <= a;
    layer2_outputs(2106) <= not (a or b);
    layer2_outputs(2107) <= b;
    layer2_outputs(2108) <= a;
    layer2_outputs(2109) <= not (a and b);
    layer2_outputs(2110) <= not b or a;
    layer2_outputs(2111) <= not (a xor b);
    layer2_outputs(2112) <= not a or b;
    layer2_outputs(2113) <= not (a and b);
    layer2_outputs(2114) <= a and not b;
    layer2_outputs(2115) <= a and not b;
    layer2_outputs(2116) <= not b or a;
    layer2_outputs(2117) <= a;
    layer2_outputs(2118) <= not (a xor b);
    layer2_outputs(2119) <= not (a and b);
    layer2_outputs(2120) <= not a;
    layer2_outputs(2121) <= not (a xor b);
    layer2_outputs(2122) <= not a or b;
    layer2_outputs(2123) <= a and not b;
    layer2_outputs(2124) <= a and b;
    layer2_outputs(2125) <= not (a and b);
    layer2_outputs(2126) <= not b;
    layer2_outputs(2127) <= not (a or b);
    layer2_outputs(2128) <= not b;
    layer2_outputs(2129) <= a;
    layer2_outputs(2130) <= not (a and b);
    layer2_outputs(2131) <= not a;
    layer2_outputs(2132) <= a or b;
    layer2_outputs(2133) <= not b or a;
    layer2_outputs(2134) <= not (a or b);
    layer2_outputs(2135) <= not (a or b);
    layer2_outputs(2136) <= a or b;
    layer2_outputs(2137) <= a and b;
    layer2_outputs(2138) <= b;
    layer2_outputs(2139) <= not a or b;
    layer2_outputs(2140) <= a;
    layer2_outputs(2141) <= not b or a;
    layer2_outputs(2142) <= b and not a;
    layer2_outputs(2143) <= b and not a;
    layer2_outputs(2144) <= b and not a;
    layer2_outputs(2145) <= b;
    layer2_outputs(2146) <= a xor b;
    layer2_outputs(2147) <= not (a or b);
    layer2_outputs(2148) <= b;
    layer2_outputs(2149) <= a xor b;
    layer2_outputs(2150) <= not (a xor b);
    layer2_outputs(2151) <= not b;
    layer2_outputs(2152) <= b and not a;
    layer2_outputs(2153) <= b;
    layer2_outputs(2154) <= a or b;
    layer2_outputs(2155) <= a or b;
    layer2_outputs(2156) <= not (a or b);
    layer2_outputs(2157) <= not (a xor b);
    layer2_outputs(2158) <= not b;
    layer2_outputs(2159) <= b and not a;
    layer2_outputs(2160) <= not b;
    layer2_outputs(2161) <= not a;
    layer2_outputs(2162) <= not a;
    layer2_outputs(2163) <= b;
    layer2_outputs(2164) <= b;
    layer2_outputs(2165) <= not (a xor b);
    layer2_outputs(2166) <= b;
    layer2_outputs(2167) <= not a;
    layer2_outputs(2168) <= a and b;
    layer2_outputs(2169) <= a and not b;
    layer2_outputs(2170) <= not a or b;
    layer2_outputs(2171) <= a;
    layer2_outputs(2172) <= a and b;
    layer2_outputs(2173) <= not a;
    layer2_outputs(2174) <= b;
    layer2_outputs(2175) <= not (a xor b);
    layer2_outputs(2176) <= not b;
    layer2_outputs(2177) <= a and b;
    layer2_outputs(2178) <= a;
    layer2_outputs(2179) <= not b or a;
    layer2_outputs(2180) <= a and not b;
    layer2_outputs(2181) <= not a or b;
    layer2_outputs(2182) <= not (a xor b);
    layer2_outputs(2183) <= b;
    layer2_outputs(2184) <= a xor b;
    layer2_outputs(2185) <= b and not a;
    layer2_outputs(2186) <= b;
    layer2_outputs(2187) <= a and b;
    layer2_outputs(2188) <= a or b;
    layer2_outputs(2189) <= b;
    layer2_outputs(2190) <= not b;
    layer2_outputs(2191) <= a xor b;
    layer2_outputs(2192) <= not (a xor b);
    layer2_outputs(2193) <= not (a and b);
    layer2_outputs(2194) <= a and not b;
    layer2_outputs(2195) <= a;
    layer2_outputs(2196) <= b;
    layer2_outputs(2197) <= a and b;
    layer2_outputs(2198) <= a and not b;
    layer2_outputs(2199) <= b and not a;
    layer2_outputs(2200) <= not a or b;
    layer2_outputs(2201) <= a and b;
    layer2_outputs(2202) <= a xor b;
    layer2_outputs(2203) <= a;
    layer2_outputs(2204) <= not b;
    layer2_outputs(2205) <= not a;
    layer2_outputs(2206) <= b;
    layer2_outputs(2207) <= not (a and b);
    layer2_outputs(2208) <= b;
    layer2_outputs(2209) <= not (a or b);
    layer2_outputs(2210) <= not (a xor b);
    layer2_outputs(2211) <= a or b;
    layer2_outputs(2212) <= not (a or b);
    layer2_outputs(2213) <= b;
    layer2_outputs(2214) <= not a;
    layer2_outputs(2215) <= a or b;
    layer2_outputs(2216) <= not b;
    layer2_outputs(2217) <= not (a xor b);
    layer2_outputs(2218) <= a;
    layer2_outputs(2219) <= a or b;
    layer2_outputs(2220) <= not (a and b);
    layer2_outputs(2221) <= not b;
    layer2_outputs(2222) <= b;
    layer2_outputs(2223) <= a or b;
    layer2_outputs(2224) <= not (a and b);
    layer2_outputs(2225) <= not a;
    layer2_outputs(2226) <= b;
    layer2_outputs(2227) <= a and b;
    layer2_outputs(2228) <= not (a or b);
    layer2_outputs(2229) <= not (a and b);
    layer2_outputs(2230) <= b and not a;
    layer2_outputs(2231) <= not b or a;
    layer2_outputs(2232) <= not (a and b);
    layer2_outputs(2233) <= a;
    layer2_outputs(2234) <= a xor b;
    layer2_outputs(2235) <= not a;
    layer2_outputs(2236) <= a;
    layer2_outputs(2237) <= not (a xor b);
    layer2_outputs(2238) <= b;
    layer2_outputs(2239) <= not (a or b);
    layer2_outputs(2240) <= a and b;
    layer2_outputs(2241) <= not (a xor b);
    layer2_outputs(2242) <= a xor b;
    layer2_outputs(2243) <= not a or b;
    layer2_outputs(2244) <= not b;
    layer2_outputs(2245) <= a xor b;
    layer2_outputs(2246) <= not b;
    layer2_outputs(2247) <= not b or a;
    layer2_outputs(2248) <= a xor b;
    layer2_outputs(2249) <= not b or a;
    layer2_outputs(2250) <= b;
    layer2_outputs(2251) <= not a;
    layer2_outputs(2252) <= a and not b;
    layer2_outputs(2253) <= b and not a;
    layer2_outputs(2254) <= a xor b;
    layer2_outputs(2255) <= not a;
    layer2_outputs(2256) <= not (a or b);
    layer2_outputs(2257) <= a and not b;
    layer2_outputs(2258) <= a;
    layer2_outputs(2259) <= b;
    layer2_outputs(2260) <= not a or b;
    layer2_outputs(2261) <= not a;
    layer2_outputs(2262) <= a;
    layer2_outputs(2263) <= not b;
    layer2_outputs(2264) <= not (a xor b);
    layer2_outputs(2265) <= not (a or b);
    layer2_outputs(2266) <= a and not b;
    layer2_outputs(2267) <= a xor b;
    layer2_outputs(2268) <= not (a and b);
    layer2_outputs(2269) <= not b;
    layer2_outputs(2270) <= a xor b;
    layer2_outputs(2271) <= not b or a;
    layer2_outputs(2272) <= not a;
    layer2_outputs(2273) <= not a;
    layer2_outputs(2274) <= not (a and b);
    layer2_outputs(2275) <= not (a or b);
    layer2_outputs(2276) <= not (a xor b);
    layer2_outputs(2277) <= not a;
    layer2_outputs(2278) <= not b;
    layer2_outputs(2279) <= not (a or b);
    layer2_outputs(2280) <= not (a xor b);
    layer2_outputs(2281) <= not b or a;
    layer2_outputs(2282) <= not (a or b);
    layer2_outputs(2283) <= not a;
    layer2_outputs(2284) <= not (a or b);
    layer2_outputs(2285) <= not b;
    layer2_outputs(2286) <= b and not a;
    layer2_outputs(2287) <= a;
    layer2_outputs(2288) <= not (a or b);
    layer2_outputs(2289) <= not (a xor b);
    layer2_outputs(2290) <= not a;
    layer2_outputs(2291) <= not a;
    layer2_outputs(2292) <= a;
    layer2_outputs(2293) <= a and b;
    layer2_outputs(2294) <= not b or a;
    layer2_outputs(2295) <= not (a xor b);
    layer2_outputs(2296) <= a or b;
    layer2_outputs(2297) <= not (a and b);
    layer2_outputs(2298) <= a and b;
    layer2_outputs(2299) <= not a or b;
    layer2_outputs(2300) <= a and b;
    layer2_outputs(2301) <= not a;
    layer2_outputs(2302) <= a and b;
    layer2_outputs(2303) <= not (a or b);
    layer2_outputs(2304) <= not (a and b);
    layer2_outputs(2305) <= not a or b;
    layer2_outputs(2306) <= a xor b;
    layer2_outputs(2307) <= not (a xor b);
    layer2_outputs(2308) <= not (a and b);
    layer2_outputs(2309) <= b and not a;
    layer2_outputs(2310) <= b and not a;
    layer2_outputs(2311) <= not (a xor b);
    layer2_outputs(2312) <= a and b;
    layer2_outputs(2313) <= not b;
    layer2_outputs(2314) <= a xor b;
    layer2_outputs(2315) <= not (a and b);
    layer2_outputs(2316) <= b and not a;
    layer2_outputs(2317) <= a and not b;
    layer2_outputs(2318) <= b;
    layer2_outputs(2319) <= b;
    layer2_outputs(2320) <= not (a and b);
    layer2_outputs(2321) <= a;
    layer2_outputs(2322) <= not a or b;
    layer2_outputs(2323) <= not b or a;
    layer2_outputs(2324) <= a or b;
    layer2_outputs(2325) <= a xor b;
    layer2_outputs(2326) <= not b or a;
    layer2_outputs(2327) <= not (a xor b);
    layer2_outputs(2328) <= a;
    layer2_outputs(2329) <= not a;
    layer2_outputs(2330) <= a and b;
    layer2_outputs(2331) <= a or b;
    layer2_outputs(2332) <= not b;
    layer2_outputs(2333) <= a xor b;
    layer2_outputs(2334) <= a;
    layer2_outputs(2335) <= not (a xor b);
    layer2_outputs(2336) <= a and not b;
    layer2_outputs(2337) <= b and not a;
    layer2_outputs(2338) <= a;
    layer2_outputs(2339) <= a;
    layer2_outputs(2340) <= not b or a;
    layer2_outputs(2341) <= a xor b;
    layer2_outputs(2342) <= not a;
    layer2_outputs(2343) <= not b;
    layer2_outputs(2344) <= not a;
    layer2_outputs(2345) <= a;
    layer2_outputs(2346) <= not (a or b);
    layer2_outputs(2347) <= a and not b;
    layer2_outputs(2348) <= a and not b;
    layer2_outputs(2349) <= a;
    layer2_outputs(2350) <= not a;
    layer2_outputs(2351) <= not a;
    layer2_outputs(2352) <= a and not b;
    layer2_outputs(2353) <= a;
    layer2_outputs(2354) <= not b;
    layer2_outputs(2355) <= a and b;
    layer2_outputs(2356) <= b and not a;
    layer2_outputs(2357) <= not (a xor b);
    layer2_outputs(2358) <= not b;
    layer2_outputs(2359) <= not (a and b);
    layer2_outputs(2360) <= a;
    layer2_outputs(2361) <= not (a xor b);
    layer2_outputs(2362) <= not (a or b);
    layer2_outputs(2363) <= not b or a;
    layer2_outputs(2364) <= not (a or b);
    layer2_outputs(2365) <= a and not b;
    layer2_outputs(2366) <= b;
    layer2_outputs(2367) <= a and not b;
    layer2_outputs(2368) <= a and b;
    layer2_outputs(2369) <= not (a and b);
    layer2_outputs(2370) <= not a;
    layer2_outputs(2371) <= not (a xor b);
    layer2_outputs(2372) <= a and b;
    layer2_outputs(2373) <= a and not b;
    layer2_outputs(2374) <= not b or a;
    layer2_outputs(2375) <= not (a xor b);
    layer2_outputs(2376) <= b;
    layer2_outputs(2377) <= not (a xor b);
    layer2_outputs(2378) <= not a or b;
    layer2_outputs(2379) <= not (a xor b);
    layer2_outputs(2380) <= a;
    layer2_outputs(2381) <= not (a or b);
    layer2_outputs(2382) <= not (a and b);
    layer2_outputs(2383) <= a and b;
    layer2_outputs(2384) <= not (a and b);
    layer2_outputs(2385) <= a and not b;
    layer2_outputs(2386) <= not b or a;
    layer2_outputs(2387) <= a xor b;
    layer2_outputs(2388) <= not (a xor b);
    layer2_outputs(2389) <= a xor b;
    layer2_outputs(2390) <= a or b;
    layer2_outputs(2391) <= a and b;
    layer2_outputs(2392) <= not (a xor b);
    layer2_outputs(2393) <= b;
    layer2_outputs(2394) <= a xor b;
    layer2_outputs(2395) <= b;
    layer2_outputs(2396) <= not b;
    layer2_outputs(2397) <= not (a and b);
    layer2_outputs(2398) <= not a or b;
    layer2_outputs(2399) <= not b or a;
    layer2_outputs(2400) <= b and not a;
    layer2_outputs(2401) <= not (a xor b);
    layer2_outputs(2402) <= not (a xor b);
    layer2_outputs(2403) <= not a;
    layer2_outputs(2404) <= b and not a;
    layer2_outputs(2405) <= not b or a;
    layer2_outputs(2406) <= not b or a;
    layer2_outputs(2407) <= not a or b;
    layer2_outputs(2408) <= not b or a;
    layer2_outputs(2409) <= not b;
    layer2_outputs(2410) <= not (a xor b);
    layer2_outputs(2411) <= a;
    layer2_outputs(2412) <= not a;
    layer2_outputs(2413) <= not b;
    layer2_outputs(2414) <= b;
    layer2_outputs(2415) <= a;
    layer2_outputs(2416) <= not b or a;
    layer2_outputs(2417) <= b;
    layer2_outputs(2418) <= not a;
    layer2_outputs(2419) <= a and not b;
    layer2_outputs(2420) <= not a;
    layer2_outputs(2421) <= not a;
    layer2_outputs(2422) <= a and not b;
    layer2_outputs(2423) <= not (a xor b);
    layer2_outputs(2424) <= not b or a;
    layer2_outputs(2425) <= a and b;
    layer2_outputs(2426) <= b;
    layer2_outputs(2427) <= b;
    layer2_outputs(2428) <= not a or b;
    layer2_outputs(2429) <= a and b;
    layer2_outputs(2430) <= not a;
    layer2_outputs(2431) <= not (a or b);
    layer2_outputs(2432) <= a xor b;
    layer2_outputs(2433) <= not a;
    layer2_outputs(2434) <= not a or b;
    layer2_outputs(2435) <= not a;
    layer2_outputs(2436) <= b;
    layer2_outputs(2437) <= a or b;
    layer2_outputs(2438) <= a or b;
    layer2_outputs(2439) <= not b;
    layer2_outputs(2440) <= not (a xor b);
    layer2_outputs(2441) <= not b or a;
    layer2_outputs(2442) <= a and not b;
    layer2_outputs(2443) <= a;
    layer2_outputs(2444) <= not (a or b);
    layer2_outputs(2445) <= not b or a;
    layer2_outputs(2446) <= not (a xor b);
    layer2_outputs(2447) <= not (a xor b);
    layer2_outputs(2448) <= not (a and b);
    layer2_outputs(2449) <= not b;
    layer2_outputs(2450) <= not b or a;
    layer2_outputs(2451) <= not b or a;
    layer2_outputs(2452) <= a;
    layer2_outputs(2453) <= a xor b;
    layer2_outputs(2454) <= a;
    layer2_outputs(2455) <= a and b;
    layer2_outputs(2456) <= not (a or b);
    layer2_outputs(2457) <= a or b;
    layer2_outputs(2458) <= b;
    layer2_outputs(2459) <= a and not b;
    layer2_outputs(2460) <= not (a and b);
    layer2_outputs(2461) <= not a;
    layer2_outputs(2462) <= a;
    layer2_outputs(2463) <= not b or a;
    layer2_outputs(2464) <= a and not b;
    layer2_outputs(2465) <= a;
    layer2_outputs(2466) <= not b or a;
    layer2_outputs(2467) <= not (a xor b);
    layer2_outputs(2468) <= a;
    layer2_outputs(2469) <= '0';
    layer2_outputs(2470) <= not a or b;
    layer2_outputs(2471) <= a xor b;
    layer2_outputs(2472) <= not (a or b);
    layer2_outputs(2473) <= b and not a;
    layer2_outputs(2474) <= not (a and b);
    layer2_outputs(2475) <= not a;
    layer2_outputs(2476) <= b and not a;
    layer2_outputs(2477) <= not b;
    layer2_outputs(2478) <= b;
    layer2_outputs(2479) <= a and not b;
    layer2_outputs(2480) <= not (a and b);
    layer2_outputs(2481) <= a xor b;
    layer2_outputs(2482) <= b;
    layer2_outputs(2483) <= b and not a;
    layer2_outputs(2484) <= a;
    layer2_outputs(2485) <= a;
    layer2_outputs(2486) <= a and b;
    layer2_outputs(2487) <= not (a or b);
    layer2_outputs(2488) <= not (a or b);
    layer2_outputs(2489) <= a and b;
    layer2_outputs(2490) <= a;
    layer2_outputs(2491) <= not b;
    layer2_outputs(2492) <= not (a or b);
    layer2_outputs(2493) <= not a;
    layer2_outputs(2494) <= not (a xor b);
    layer2_outputs(2495) <= not b or a;
    layer2_outputs(2496) <= a xor b;
    layer2_outputs(2497) <= a;
    layer2_outputs(2498) <= not a;
    layer2_outputs(2499) <= a and b;
    layer2_outputs(2500) <= not a;
    layer2_outputs(2501) <= b and not a;
    layer2_outputs(2502) <= not a;
    layer2_outputs(2503) <= b;
    layer2_outputs(2504) <= a;
    layer2_outputs(2505) <= not (a and b);
    layer2_outputs(2506) <= not a or b;
    layer2_outputs(2507) <= not b;
    layer2_outputs(2508) <= b;
    layer2_outputs(2509) <= not b;
    layer2_outputs(2510) <= a or b;
    layer2_outputs(2511) <= a or b;
    layer2_outputs(2512) <= not a;
    layer2_outputs(2513) <= not a;
    layer2_outputs(2514) <= not (a or b);
    layer2_outputs(2515) <= not (a or b);
    layer2_outputs(2516) <= not (a xor b);
    layer2_outputs(2517) <= not (a xor b);
    layer2_outputs(2518) <= not b;
    layer2_outputs(2519) <= not b;
    layer2_outputs(2520) <= not b;
    layer2_outputs(2521) <= not (a xor b);
    layer2_outputs(2522) <= a xor b;
    layer2_outputs(2523) <= b and not a;
    layer2_outputs(2524) <= b and not a;
    layer2_outputs(2525) <= a xor b;
    layer2_outputs(2526) <= not (a and b);
    layer2_outputs(2527) <= a and b;
    layer2_outputs(2528) <= not a;
    layer2_outputs(2529) <= a or b;
    layer2_outputs(2530) <= not (a xor b);
    layer2_outputs(2531) <= not b or a;
    layer2_outputs(2532) <= b;
    layer2_outputs(2533) <= a and not b;
    layer2_outputs(2534) <= a xor b;
    layer2_outputs(2535) <= b and not a;
    layer2_outputs(2536) <= not a;
    layer2_outputs(2537) <= a and b;
    layer2_outputs(2538) <= a;
    layer2_outputs(2539) <= a and not b;
    layer2_outputs(2540) <= not (a and b);
    layer2_outputs(2541) <= a or b;
    layer2_outputs(2542) <= '0';
    layer2_outputs(2543) <= b;
    layer2_outputs(2544) <= a;
    layer2_outputs(2545) <= a and not b;
    layer2_outputs(2546) <= b and not a;
    layer2_outputs(2547) <= not a;
    layer2_outputs(2548) <= a and b;
    layer2_outputs(2549) <= not a;
    layer2_outputs(2550) <= not b;
    layer2_outputs(2551) <= not a or b;
    layer2_outputs(2552) <= not b or a;
    layer2_outputs(2553) <= not b or a;
    layer2_outputs(2554) <= a and not b;
    layer2_outputs(2555) <= not (a xor b);
    layer2_outputs(2556) <= a;
    layer2_outputs(2557) <= b;
    layer2_outputs(2558) <= not a;
    layer2_outputs(2559) <= not a;
    layer2_outputs(2560) <= a and b;
    layer2_outputs(2561) <= a;
    layer2_outputs(2562) <= b and not a;
    layer2_outputs(2563) <= not b;
    layer2_outputs(2564) <= not a;
    layer2_outputs(2565) <= b;
    layer2_outputs(2566) <= not a or b;
    layer2_outputs(2567) <= b and not a;
    layer2_outputs(2568) <= not b or a;
    layer2_outputs(2569) <= b and not a;
    layer2_outputs(2570) <= not (a and b);
    layer2_outputs(2571) <= a xor b;
    layer2_outputs(2572) <= a;
    layer2_outputs(2573) <= a;
    layer2_outputs(2574) <= not (a or b);
    layer2_outputs(2575) <= a xor b;
    layer2_outputs(2576) <= a;
    layer2_outputs(2577) <= not (a or b);
    layer2_outputs(2578) <= a;
    layer2_outputs(2579) <= not b;
    layer2_outputs(2580) <= not (a and b);
    layer2_outputs(2581) <= not (a xor b);
    layer2_outputs(2582) <= a or b;
    layer2_outputs(2583) <= not a;
    layer2_outputs(2584) <= not (a or b);
    layer2_outputs(2585) <= a;
    layer2_outputs(2586) <= b and not a;
    layer2_outputs(2587) <= a xor b;
    layer2_outputs(2588) <= a xor b;
    layer2_outputs(2589) <= not a or b;
    layer2_outputs(2590) <= not a or b;
    layer2_outputs(2591) <= not a;
    layer2_outputs(2592) <= b;
    layer2_outputs(2593) <= a and b;
    layer2_outputs(2594) <= not a;
    layer2_outputs(2595) <= a or b;
    layer2_outputs(2596) <= not b or a;
    layer2_outputs(2597) <= not (a xor b);
    layer2_outputs(2598) <= b and not a;
    layer2_outputs(2599) <= not a or b;
    layer2_outputs(2600) <= a;
    layer2_outputs(2601) <= not b or a;
    layer2_outputs(2602) <= a and not b;
    layer2_outputs(2603) <= a;
    layer2_outputs(2604) <= not a or b;
    layer2_outputs(2605) <= a and b;
    layer2_outputs(2606) <= b and not a;
    layer2_outputs(2607) <= not a;
    layer2_outputs(2608) <= a or b;
    layer2_outputs(2609) <= not b;
    layer2_outputs(2610) <= not a or b;
    layer2_outputs(2611) <= not a;
    layer2_outputs(2612) <= not a;
    layer2_outputs(2613) <= not (a or b);
    layer2_outputs(2614) <= a or b;
    layer2_outputs(2615) <= not (a or b);
    layer2_outputs(2616) <= not b or a;
    layer2_outputs(2617) <= not b;
    layer2_outputs(2618) <= not b or a;
    layer2_outputs(2619) <= a;
    layer2_outputs(2620) <= a xor b;
    layer2_outputs(2621) <= not b or a;
    layer2_outputs(2622) <= not (a and b);
    layer2_outputs(2623) <= b;
    layer2_outputs(2624) <= not (a and b);
    layer2_outputs(2625) <= a or b;
    layer2_outputs(2626) <= not b or a;
    layer2_outputs(2627) <= a xor b;
    layer2_outputs(2628) <= a and b;
    layer2_outputs(2629) <= a or b;
    layer2_outputs(2630) <= b;
    layer2_outputs(2631) <= not a;
    layer2_outputs(2632) <= not (a and b);
    layer2_outputs(2633) <= a and not b;
    layer2_outputs(2634) <= a and b;
    layer2_outputs(2635) <= not b;
    layer2_outputs(2636) <= not a or b;
    layer2_outputs(2637) <= b and not a;
    layer2_outputs(2638) <= not b;
    layer2_outputs(2639) <= a;
    layer2_outputs(2640) <= b and not a;
    layer2_outputs(2641) <= not (a xor b);
    layer2_outputs(2642) <= a;
    layer2_outputs(2643) <= not (a and b);
    layer2_outputs(2644) <= a;
    layer2_outputs(2645) <= not (a and b);
    layer2_outputs(2646) <= a xor b;
    layer2_outputs(2647) <= not a or b;
    layer2_outputs(2648) <= a and not b;
    layer2_outputs(2649) <= a;
    layer2_outputs(2650) <= not a;
    layer2_outputs(2651) <= a;
    layer2_outputs(2652) <= a and not b;
    layer2_outputs(2653) <= a and b;
    layer2_outputs(2654) <= not b or a;
    layer2_outputs(2655) <= not a or b;
    layer2_outputs(2656) <= b and not a;
    layer2_outputs(2657) <= b;
    layer2_outputs(2658) <= not b;
    layer2_outputs(2659) <= a;
    layer2_outputs(2660) <= b;
    layer2_outputs(2661) <= not (a xor b);
    layer2_outputs(2662) <= b;
    layer2_outputs(2663) <= a and b;
    layer2_outputs(2664) <= a xor b;
    layer2_outputs(2665) <= a xor b;
    layer2_outputs(2666) <= a xor b;
    layer2_outputs(2667) <= not a;
    layer2_outputs(2668) <= not (a xor b);
    layer2_outputs(2669) <= a;
    layer2_outputs(2670) <= not b;
    layer2_outputs(2671) <= not (a and b);
    layer2_outputs(2672) <= not b or a;
    layer2_outputs(2673) <= not (a xor b);
    layer2_outputs(2674) <= a or b;
    layer2_outputs(2675) <= not b or a;
    layer2_outputs(2676) <= a;
    layer2_outputs(2677) <= a;
    layer2_outputs(2678) <= a and not b;
    layer2_outputs(2679) <= a or b;
    layer2_outputs(2680) <= b and not a;
    layer2_outputs(2681) <= not a;
    layer2_outputs(2682) <= not b;
    layer2_outputs(2683) <= b;
    layer2_outputs(2684) <= not a;
    layer2_outputs(2685) <= a xor b;
    layer2_outputs(2686) <= a or b;
    layer2_outputs(2687) <= a xor b;
    layer2_outputs(2688) <= not (a or b);
    layer2_outputs(2689) <= a;
    layer2_outputs(2690) <= b;
    layer2_outputs(2691) <= not a;
    layer2_outputs(2692) <= not (a and b);
    layer2_outputs(2693) <= a or b;
    layer2_outputs(2694) <= a;
    layer2_outputs(2695) <= b and not a;
    layer2_outputs(2696) <= a and b;
    layer2_outputs(2697) <= a and not b;
    layer2_outputs(2698) <= not b or a;
    layer2_outputs(2699) <= a;
    layer2_outputs(2700) <= b;
    layer2_outputs(2701) <= not a or b;
    layer2_outputs(2702) <= b and not a;
    layer2_outputs(2703) <= a or b;
    layer2_outputs(2704) <= a;
    layer2_outputs(2705) <= not b;
    layer2_outputs(2706) <= not a or b;
    layer2_outputs(2707) <= a and b;
    layer2_outputs(2708) <= a xor b;
    layer2_outputs(2709) <= not b;
    layer2_outputs(2710) <= not (a and b);
    layer2_outputs(2711) <= not a or b;
    layer2_outputs(2712) <= b;
    layer2_outputs(2713) <= a or b;
    layer2_outputs(2714) <= b;
    layer2_outputs(2715) <= not a;
    layer2_outputs(2716) <= not b or a;
    layer2_outputs(2717) <= a xor b;
    layer2_outputs(2718) <= not a;
    layer2_outputs(2719) <= not b;
    layer2_outputs(2720) <= b and not a;
    layer2_outputs(2721) <= not (a and b);
    layer2_outputs(2722) <= b;
    layer2_outputs(2723) <= a;
    layer2_outputs(2724) <= not b;
    layer2_outputs(2725) <= not a;
    layer2_outputs(2726) <= b;
    layer2_outputs(2727) <= not a;
    layer2_outputs(2728) <= b and not a;
    layer2_outputs(2729) <= b and not a;
    layer2_outputs(2730) <= not (a and b);
    layer2_outputs(2731) <= not (a xor b);
    layer2_outputs(2732) <= a;
    layer2_outputs(2733) <= not b;
    layer2_outputs(2734) <= not (a and b);
    layer2_outputs(2735) <= not (a xor b);
    layer2_outputs(2736) <= b and not a;
    layer2_outputs(2737) <= not b;
    layer2_outputs(2738) <= not a or b;
    layer2_outputs(2739) <= not (a xor b);
    layer2_outputs(2740) <= not a;
    layer2_outputs(2741) <= not a;
    layer2_outputs(2742) <= not a or b;
    layer2_outputs(2743) <= a;
    layer2_outputs(2744) <= not (a xor b);
    layer2_outputs(2745) <= a and not b;
    layer2_outputs(2746) <= not (a or b);
    layer2_outputs(2747) <= not b;
    layer2_outputs(2748) <= b and not a;
    layer2_outputs(2749) <= not a;
    layer2_outputs(2750) <= a xor b;
    layer2_outputs(2751) <= a;
    layer2_outputs(2752) <= not a;
    layer2_outputs(2753) <= a;
    layer2_outputs(2754) <= b;
    layer2_outputs(2755) <= not b;
    layer2_outputs(2756) <= b;
    layer2_outputs(2757) <= a and not b;
    layer2_outputs(2758) <= not a;
    layer2_outputs(2759) <= not b;
    layer2_outputs(2760) <= b;
    layer2_outputs(2761) <= not (a xor b);
    layer2_outputs(2762) <= a and b;
    layer2_outputs(2763) <= not (a or b);
    layer2_outputs(2764) <= not a or b;
    layer2_outputs(2765) <= a xor b;
    layer2_outputs(2766) <= b;
    layer2_outputs(2767) <= b;
    layer2_outputs(2768) <= not (a or b);
    layer2_outputs(2769) <= not (a xor b);
    layer2_outputs(2770) <= not a;
    layer2_outputs(2771) <= a and b;
    layer2_outputs(2772) <= not a or b;
    layer2_outputs(2773) <= not a;
    layer2_outputs(2774) <= not (a and b);
    layer2_outputs(2775) <= a and b;
    layer2_outputs(2776) <= b;
    layer2_outputs(2777) <= not (a xor b);
    layer2_outputs(2778) <= not b or a;
    layer2_outputs(2779) <= a and b;
    layer2_outputs(2780) <= a or b;
    layer2_outputs(2781) <= not b;
    layer2_outputs(2782) <= not (a xor b);
    layer2_outputs(2783) <= b;
    layer2_outputs(2784) <= not (a xor b);
    layer2_outputs(2785) <= not (a or b);
    layer2_outputs(2786) <= b and not a;
    layer2_outputs(2787) <= b;
    layer2_outputs(2788) <= not a;
    layer2_outputs(2789) <= a and b;
    layer2_outputs(2790) <= not (a or b);
    layer2_outputs(2791) <= b and not a;
    layer2_outputs(2792) <= not a;
    layer2_outputs(2793) <= not a;
    layer2_outputs(2794) <= a xor b;
    layer2_outputs(2795) <= not b or a;
    layer2_outputs(2796) <= not a;
    layer2_outputs(2797) <= a xor b;
    layer2_outputs(2798) <= not (a and b);
    layer2_outputs(2799) <= a xor b;
    layer2_outputs(2800) <= not a;
    layer2_outputs(2801) <= a or b;
    layer2_outputs(2802) <= a and not b;
    layer2_outputs(2803) <= not a or b;
    layer2_outputs(2804) <= not a;
    layer2_outputs(2805) <= not a or b;
    layer2_outputs(2806) <= a;
    layer2_outputs(2807) <= not (a xor b);
    layer2_outputs(2808) <= not b or a;
    layer2_outputs(2809) <= not b or a;
    layer2_outputs(2810) <= b and not a;
    layer2_outputs(2811) <= not a;
    layer2_outputs(2812) <= not b;
    layer2_outputs(2813) <= a and b;
    layer2_outputs(2814) <= not a or b;
    layer2_outputs(2815) <= not a or b;
    layer2_outputs(2816) <= a;
    layer2_outputs(2817) <= a and b;
    layer2_outputs(2818) <= not a or b;
    layer2_outputs(2819) <= not (a or b);
    layer2_outputs(2820) <= b and not a;
    layer2_outputs(2821) <= not (a xor b);
    layer2_outputs(2822) <= not a or b;
    layer2_outputs(2823) <= not b;
    layer2_outputs(2824) <= not (a xor b);
    layer2_outputs(2825) <= not b;
    layer2_outputs(2826) <= not a;
    layer2_outputs(2827) <= not (a xor b);
    layer2_outputs(2828) <= a or b;
    layer2_outputs(2829) <= '0';
    layer2_outputs(2830) <= b and not a;
    layer2_outputs(2831) <= a;
    layer2_outputs(2832) <= not b;
    layer2_outputs(2833) <= b and not a;
    layer2_outputs(2834) <= not b or a;
    layer2_outputs(2835) <= not (a xor b);
    layer2_outputs(2836) <= a xor b;
    layer2_outputs(2837) <= not a;
    layer2_outputs(2838) <= a or b;
    layer2_outputs(2839) <= a;
    layer2_outputs(2840) <= not a or b;
    layer2_outputs(2841) <= a xor b;
    layer2_outputs(2842) <= not (a or b);
    layer2_outputs(2843) <= not (a and b);
    layer2_outputs(2844) <= not (a xor b);
    layer2_outputs(2845) <= a xor b;
    layer2_outputs(2846) <= a and b;
    layer2_outputs(2847) <= not (a and b);
    layer2_outputs(2848) <= a or b;
    layer2_outputs(2849) <= a xor b;
    layer2_outputs(2850) <= a and not b;
    layer2_outputs(2851) <= not b;
    layer2_outputs(2852) <= not b or a;
    layer2_outputs(2853) <= not (a and b);
    layer2_outputs(2854) <= a xor b;
    layer2_outputs(2855) <= not a or b;
    layer2_outputs(2856) <= a and not b;
    layer2_outputs(2857) <= not a;
    layer2_outputs(2858) <= a;
    layer2_outputs(2859) <= not (a or b);
    layer2_outputs(2860) <= not a;
    layer2_outputs(2861) <= a xor b;
    layer2_outputs(2862) <= not b or a;
    layer2_outputs(2863) <= not (a xor b);
    layer2_outputs(2864) <= not (a xor b);
    layer2_outputs(2865) <= a;
    layer2_outputs(2866) <= a or b;
    layer2_outputs(2867) <= not a;
    layer2_outputs(2868) <= a;
    layer2_outputs(2869) <= a xor b;
    layer2_outputs(2870) <= not a;
    layer2_outputs(2871) <= not b;
    layer2_outputs(2872) <= not (a xor b);
    layer2_outputs(2873) <= not (a xor b);
    layer2_outputs(2874) <= a or b;
    layer2_outputs(2875) <= a and b;
    layer2_outputs(2876) <= not b;
    layer2_outputs(2877) <= not b or a;
    layer2_outputs(2878) <= a or b;
    layer2_outputs(2879) <= not b or a;
    layer2_outputs(2880) <= a xor b;
    layer2_outputs(2881) <= not a;
    layer2_outputs(2882) <= b;
    layer2_outputs(2883) <= a and b;
    layer2_outputs(2884) <= not a;
    layer2_outputs(2885) <= b and not a;
    layer2_outputs(2886) <= b;
    layer2_outputs(2887) <= not (a xor b);
    layer2_outputs(2888) <= a xor b;
    layer2_outputs(2889) <= a and b;
    layer2_outputs(2890) <= not (a and b);
    layer2_outputs(2891) <= a xor b;
    layer2_outputs(2892) <= not a;
    layer2_outputs(2893) <= not a;
    layer2_outputs(2894) <= a xor b;
    layer2_outputs(2895) <= not (a xor b);
    layer2_outputs(2896) <= a or b;
    layer2_outputs(2897) <= not a or b;
    layer2_outputs(2898) <= a and b;
    layer2_outputs(2899) <= a and b;
    layer2_outputs(2900) <= not b;
    layer2_outputs(2901) <= a and b;
    layer2_outputs(2902) <= not (a xor b);
    layer2_outputs(2903) <= b;
    layer2_outputs(2904) <= b and not a;
    layer2_outputs(2905) <= not b;
    layer2_outputs(2906) <= not (a xor b);
    layer2_outputs(2907) <= not (a or b);
    layer2_outputs(2908) <= b;
    layer2_outputs(2909) <= not b or a;
    layer2_outputs(2910) <= a and not b;
    layer2_outputs(2911) <= not b;
    layer2_outputs(2912) <= not a or b;
    layer2_outputs(2913) <= b;
    layer2_outputs(2914) <= a and not b;
    layer2_outputs(2915) <= not a;
    layer2_outputs(2916) <= a and b;
    layer2_outputs(2917) <= b;
    layer2_outputs(2918) <= b and not a;
    layer2_outputs(2919) <= not (a xor b);
    layer2_outputs(2920) <= a or b;
    layer2_outputs(2921) <= not b;
    layer2_outputs(2922) <= not b or a;
    layer2_outputs(2923) <= a and not b;
    layer2_outputs(2924) <= not (a xor b);
    layer2_outputs(2925) <= not a;
    layer2_outputs(2926) <= not a;
    layer2_outputs(2927) <= a xor b;
    layer2_outputs(2928) <= a and not b;
    layer2_outputs(2929) <= not (a and b);
    layer2_outputs(2930) <= not b;
    layer2_outputs(2931) <= a;
    layer2_outputs(2932) <= not b;
    layer2_outputs(2933) <= b and not a;
    layer2_outputs(2934) <= not b or a;
    layer2_outputs(2935) <= a and b;
    layer2_outputs(2936) <= a;
    layer2_outputs(2937) <= b;
    layer2_outputs(2938) <= a and not b;
    layer2_outputs(2939) <= not b or a;
    layer2_outputs(2940) <= not (a xor b);
    layer2_outputs(2941) <= b and not a;
    layer2_outputs(2942) <= not a;
    layer2_outputs(2943) <= not a;
    layer2_outputs(2944) <= a and b;
    layer2_outputs(2945) <= not a;
    layer2_outputs(2946) <= not (a xor b);
    layer2_outputs(2947) <= a xor b;
    layer2_outputs(2948) <= a or b;
    layer2_outputs(2949) <= not b or a;
    layer2_outputs(2950) <= not b;
    layer2_outputs(2951) <= a and b;
    layer2_outputs(2952) <= not b;
    layer2_outputs(2953) <= not (a or b);
    layer2_outputs(2954) <= b;
    layer2_outputs(2955) <= a xor b;
    layer2_outputs(2956) <= a and not b;
    layer2_outputs(2957) <= a xor b;
    layer2_outputs(2958) <= not b;
    layer2_outputs(2959) <= b and not a;
    layer2_outputs(2960) <= a or b;
    layer2_outputs(2961) <= a;
    layer2_outputs(2962) <= a;
    layer2_outputs(2963) <= b;
    layer2_outputs(2964) <= a;
    layer2_outputs(2965) <= a;
    layer2_outputs(2966) <= a xor b;
    layer2_outputs(2967) <= not b;
    layer2_outputs(2968) <= a;
    layer2_outputs(2969) <= not a;
    layer2_outputs(2970) <= not a;
    layer2_outputs(2971) <= not a or b;
    layer2_outputs(2972) <= a;
    layer2_outputs(2973) <= not (a xor b);
    layer2_outputs(2974) <= not b;
    layer2_outputs(2975) <= not b;
    layer2_outputs(2976) <= a;
    layer2_outputs(2977) <= not b;
    layer2_outputs(2978) <= not (a xor b);
    layer2_outputs(2979) <= a;
    layer2_outputs(2980) <= not (a xor b);
    layer2_outputs(2981) <= b;
    layer2_outputs(2982) <= a xor b;
    layer2_outputs(2983) <= not b;
    layer2_outputs(2984) <= a;
    layer2_outputs(2985) <= not b;
    layer2_outputs(2986) <= b;
    layer2_outputs(2987) <= b;
    layer2_outputs(2988) <= not b;
    layer2_outputs(2989) <= a xor b;
    layer2_outputs(2990) <= b;
    layer2_outputs(2991) <= a and b;
    layer2_outputs(2992) <= not (a xor b);
    layer2_outputs(2993) <= a;
    layer2_outputs(2994) <= a and b;
    layer2_outputs(2995) <= not (a and b);
    layer2_outputs(2996) <= a;
    layer2_outputs(2997) <= a or b;
    layer2_outputs(2998) <= not b;
    layer2_outputs(2999) <= not (a and b);
    layer2_outputs(3000) <= a or b;
    layer2_outputs(3001) <= b;
    layer2_outputs(3002) <= not (a xor b);
    layer2_outputs(3003) <= a or b;
    layer2_outputs(3004) <= b and not a;
    layer2_outputs(3005) <= not (a or b);
    layer2_outputs(3006) <= b;
    layer2_outputs(3007) <= a xor b;
    layer2_outputs(3008) <= a and b;
    layer2_outputs(3009) <= b;
    layer2_outputs(3010) <= not (a and b);
    layer2_outputs(3011) <= not a or b;
    layer2_outputs(3012) <= b;
    layer2_outputs(3013) <= not a;
    layer2_outputs(3014) <= a;
    layer2_outputs(3015) <= b;
    layer2_outputs(3016) <= not a;
    layer2_outputs(3017) <= a and b;
    layer2_outputs(3018) <= not b;
    layer2_outputs(3019) <= b;
    layer2_outputs(3020) <= not a or b;
    layer2_outputs(3021) <= a xor b;
    layer2_outputs(3022) <= not b;
    layer2_outputs(3023) <= not a or b;
    layer2_outputs(3024) <= a;
    layer2_outputs(3025) <= not (a and b);
    layer2_outputs(3026) <= not b;
    layer2_outputs(3027) <= a;
    layer2_outputs(3028) <= not (a and b);
    layer2_outputs(3029) <= not (a and b);
    layer2_outputs(3030) <= a and b;
    layer2_outputs(3031) <= b and not a;
    layer2_outputs(3032) <= b;
    layer2_outputs(3033) <= a or b;
    layer2_outputs(3034) <= not a;
    layer2_outputs(3035) <= not (a or b);
    layer2_outputs(3036) <= not a;
    layer2_outputs(3037) <= b and not a;
    layer2_outputs(3038) <= not (a xor b);
    layer2_outputs(3039) <= b and not a;
    layer2_outputs(3040) <= not (a xor b);
    layer2_outputs(3041) <= not a;
    layer2_outputs(3042) <= not (a and b);
    layer2_outputs(3043) <= not a or b;
    layer2_outputs(3044) <= a and not b;
    layer2_outputs(3045) <= a and not b;
    layer2_outputs(3046) <= a;
    layer2_outputs(3047) <= not b or a;
    layer2_outputs(3048) <= a or b;
    layer2_outputs(3049) <= not a;
    layer2_outputs(3050) <= not a or b;
    layer2_outputs(3051) <= a or b;
    layer2_outputs(3052) <= not a or b;
    layer2_outputs(3053) <= a and not b;
    layer2_outputs(3054) <= not a;
    layer2_outputs(3055) <= not a;
    layer2_outputs(3056) <= a and b;
    layer2_outputs(3057) <= b and not a;
    layer2_outputs(3058) <= not b;
    layer2_outputs(3059) <= not (a xor b);
    layer2_outputs(3060) <= '1';
    layer2_outputs(3061) <= a xor b;
    layer2_outputs(3062) <= not b or a;
    layer2_outputs(3063) <= b;
    layer2_outputs(3064) <= not b;
    layer2_outputs(3065) <= not (a or b);
    layer2_outputs(3066) <= not a or b;
    layer2_outputs(3067) <= not b or a;
    layer2_outputs(3068) <= a xor b;
    layer2_outputs(3069) <= not (a and b);
    layer2_outputs(3070) <= not b;
    layer2_outputs(3071) <= not (a xor b);
    layer2_outputs(3072) <= a;
    layer2_outputs(3073) <= not a or b;
    layer2_outputs(3074) <= a xor b;
    layer2_outputs(3075) <= not b or a;
    layer2_outputs(3076) <= a and b;
    layer2_outputs(3077) <= not (a or b);
    layer2_outputs(3078) <= a;
    layer2_outputs(3079) <= a;
    layer2_outputs(3080) <= not (a and b);
    layer2_outputs(3081) <= a and not b;
    layer2_outputs(3082) <= not (a or b);
    layer2_outputs(3083) <= b and not a;
    layer2_outputs(3084) <= a;
    layer2_outputs(3085) <= not (a or b);
    layer2_outputs(3086) <= a and b;
    layer2_outputs(3087) <= a and b;
    layer2_outputs(3088) <= a xor b;
    layer2_outputs(3089) <= b;
    layer2_outputs(3090) <= not b;
    layer2_outputs(3091) <= a;
    layer2_outputs(3092) <= not a;
    layer2_outputs(3093) <= a;
    layer2_outputs(3094) <= not b;
    layer2_outputs(3095) <= b;
    layer2_outputs(3096) <= not (a xor b);
    layer2_outputs(3097) <= not a or b;
    layer2_outputs(3098) <= not b or a;
    layer2_outputs(3099) <= a and not b;
    layer2_outputs(3100) <= not (a xor b);
    layer2_outputs(3101) <= a and b;
    layer2_outputs(3102) <= not a;
    layer2_outputs(3103) <= a;
    layer2_outputs(3104) <= not a or b;
    layer2_outputs(3105) <= b and not a;
    layer2_outputs(3106) <= b;
    layer2_outputs(3107) <= not a;
    layer2_outputs(3108) <= b;
    layer2_outputs(3109) <= a xor b;
    layer2_outputs(3110) <= b and not a;
    layer2_outputs(3111) <= b;
    layer2_outputs(3112) <= not b;
    layer2_outputs(3113) <= not a or b;
    layer2_outputs(3114) <= a and b;
    layer2_outputs(3115) <= a and b;
    layer2_outputs(3116) <= b and not a;
    layer2_outputs(3117) <= a and not b;
    layer2_outputs(3118) <= not b or a;
    layer2_outputs(3119) <= not (a or b);
    layer2_outputs(3120) <= a xor b;
    layer2_outputs(3121) <= not a;
    layer2_outputs(3122) <= a and not b;
    layer2_outputs(3123) <= not a;
    layer2_outputs(3124) <= not (a and b);
    layer2_outputs(3125) <= '1';
    layer2_outputs(3126) <= a and b;
    layer2_outputs(3127) <= a;
    layer2_outputs(3128) <= a;
    layer2_outputs(3129) <= a;
    layer2_outputs(3130) <= not b;
    layer2_outputs(3131) <= not a;
    layer2_outputs(3132) <= not (a and b);
    layer2_outputs(3133) <= not b;
    layer2_outputs(3134) <= not a or b;
    layer2_outputs(3135) <= not (a and b);
    layer2_outputs(3136) <= a xor b;
    layer2_outputs(3137) <= a and not b;
    layer2_outputs(3138) <= a or b;
    layer2_outputs(3139) <= a and not b;
    layer2_outputs(3140) <= not (a xor b);
    layer2_outputs(3141) <= a and b;
    layer2_outputs(3142) <= not a;
    layer2_outputs(3143) <= a xor b;
    layer2_outputs(3144) <= b;
    layer2_outputs(3145) <= a xor b;
    layer2_outputs(3146) <= a;
    layer2_outputs(3147) <= not (a xor b);
    layer2_outputs(3148) <= not b;
    layer2_outputs(3149) <= not b;
    layer2_outputs(3150) <= not (a xor b);
    layer2_outputs(3151) <= a and not b;
    layer2_outputs(3152) <= b;
    layer2_outputs(3153) <= a or b;
    layer2_outputs(3154) <= a xor b;
    layer2_outputs(3155) <= not (a or b);
    layer2_outputs(3156) <= a and not b;
    layer2_outputs(3157) <= not (a and b);
    layer2_outputs(3158) <= a or b;
    layer2_outputs(3159) <= a;
    layer2_outputs(3160) <= a or b;
    layer2_outputs(3161) <= not a;
    layer2_outputs(3162) <= not (a xor b);
    layer2_outputs(3163) <= b;
    layer2_outputs(3164) <= a;
    layer2_outputs(3165) <= not a or b;
    layer2_outputs(3166) <= not a;
    layer2_outputs(3167) <= a;
    layer2_outputs(3168) <= not (a xor b);
    layer2_outputs(3169) <= a xor b;
    layer2_outputs(3170) <= a and not b;
    layer2_outputs(3171) <= a and b;
    layer2_outputs(3172) <= b and not a;
    layer2_outputs(3173) <= b;
    layer2_outputs(3174) <= a and not b;
    layer2_outputs(3175) <= not a;
    layer2_outputs(3176) <= a;
    layer2_outputs(3177) <= not (a and b);
    layer2_outputs(3178) <= a or b;
    layer2_outputs(3179) <= a xor b;
    layer2_outputs(3180) <= a and not b;
    layer2_outputs(3181) <= a or b;
    layer2_outputs(3182) <= a or b;
    layer2_outputs(3183) <= not (a or b);
    layer2_outputs(3184) <= not b;
    layer2_outputs(3185) <= b;
    layer2_outputs(3186) <= a;
    layer2_outputs(3187) <= a xor b;
    layer2_outputs(3188) <= not b or a;
    layer2_outputs(3189) <= a xor b;
    layer2_outputs(3190) <= a;
    layer2_outputs(3191) <= a and not b;
    layer2_outputs(3192) <= a or b;
    layer2_outputs(3193) <= not (a xor b);
    layer2_outputs(3194) <= a and b;
    layer2_outputs(3195) <= b and not a;
    layer2_outputs(3196) <= not a;
    layer2_outputs(3197) <= b;
    layer2_outputs(3198) <= b;
    layer2_outputs(3199) <= a or b;
    layer2_outputs(3200) <= not a or b;
    layer2_outputs(3201) <= not a or b;
    layer2_outputs(3202) <= a;
    layer2_outputs(3203) <= not (a and b);
    layer2_outputs(3204) <= not (a xor b);
    layer2_outputs(3205) <= not b;
    layer2_outputs(3206) <= a and b;
    layer2_outputs(3207) <= not b;
    layer2_outputs(3208) <= not b;
    layer2_outputs(3209) <= b;
    layer2_outputs(3210) <= not (a xor b);
    layer2_outputs(3211) <= not a;
    layer2_outputs(3212) <= b;
    layer2_outputs(3213) <= not (a or b);
    layer2_outputs(3214) <= not b or a;
    layer2_outputs(3215) <= a and b;
    layer2_outputs(3216) <= a and not b;
    layer2_outputs(3217) <= a;
    layer2_outputs(3218) <= not a;
    layer2_outputs(3219) <= not (a or b);
    layer2_outputs(3220) <= a;
    layer2_outputs(3221) <= b;
    layer2_outputs(3222) <= a or b;
    layer2_outputs(3223) <= a and not b;
    layer2_outputs(3224) <= not (a and b);
    layer2_outputs(3225) <= a or b;
    layer2_outputs(3226) <= not b;
    layer2_outputs(3227) <= b and not a;
    layer2_outputs(3228) <= not a;
    layer2_outputs(3229) <= not (a xor b);
    layer2_outputs(3230) <= not b;
    layer2_outputs(3231) <= b and not a;
    layer2_outputs(3232) <= not (a xor b);
    layer2_outputs(3233) <= a xor b;
    layer2_outputs(3234) <= not b;
    layer2_outputs(3235) <= not a;
    layer2_outputs(3236) <= a and b;
    layer2_outputs(3237) <= not a;
    layer2_outputs(3238) <= a;
    layer2_outputs(3239) <= b;
    layer2_outputs(3240) <= a xor b;
    layer2_outputs(3241) <= a and b;
    layer2_outputs(3242) <= not (a or b);
    layer2_outputs(3243) <= not (a xor b);
    layer2_outputs(3244) <= not (a xor b);
    layer2_outputs(3245) <= a and b;
    layer2_outputs(3246) <= a xor b;
    layer2_outputs(3247) <= a and b;
    layer2_outputs(3248) <= not a;
    layer2_outputs(3249) <= a;
    layer2_outputs(3250) <= not (a xor b);
    layer2_outputs(3251) <= a or b;
    layer2_outputs(3252) <= not (a and b);
    layer2_outputs(3253) <= a and not b;
    layer2_outputs(3254) <= b and not a;
    layer2_outputs(3255) <= a and not b;
    layer2_outputs(3256) <= b;
    layer2_outputs(3257) <= not (a and b);
    layer2_outputs(3258) <= not a or b;
    layer2_outputs(3259) <= not b;
    layer2_outputs(3260) <= not a;
    layer2_outputs(3261) <= a xor b;
    layer2_outputs(3262) <= b;
    layer2_outputs(3263) <= not (a xor b);
    layer2_outputs(3264) <= a or b;
    layer2_outputs(3265) <= not (a xor b);
    layer2_outputs(3266) <= a xor b;
    layer2_outputs(3267) <= b;
    layer2_outputs(3268) <= not (a xor b);
    layer2_outputs(3269) <= not (a or b);
    layer2_outputs(3270) <= a and b;
    layer2_outputs(3271) <= a xor b;
    layer2_outputs(3272) <= a xor b;
    layer2_outputs(3273) <= a;
    layer2_outputs(3274) <= a or b;
    layer2_outputs(3275) <= a and not b;
    layer2_outputs(3276) <= not (a and b);
    layer2_outputs(3277) <= a;
    layer2_outputs(3278) <= a and not b;
    layer2_outputs(3279) <= a;
    layer2_outputs(3280) <= not a or b;
    layer2_outputs(3281) <= not (a xor b);
    layer2_outputs(3282) <= b and not a;
    layer2_outputs(3283) <= b;
    layer2_outputs(3284) <= not a or b;
    layer2_outputs(3285) <= not (a or b);
    layer2_outputs(3286) <= not b;
    layer2_outputs(3287) <= b;
    layer2_outputs(3288) <= not a or b;
    layer2_outputs(3289) <= not a;
    layer2_outputs(3290) <= a;
    layer2_outputs(3291) <= not (a or b);
    layer2_outputs(3292) <= not b or a;
    layer2_outputs(3293) <= a and not b;
    layer2_outputs(3294) <= not (a xor b);
    layer2_outputs(3295) <= not (a or b);
    layer2_outputs(3296) <= not b;
    layer2_outputs(3297) <= a;
    layer2_outputs(3298) <= a;
    layer2_outputs(3299) <= not b;
    layer2_outputs(3300) <= not a;
    layer2_outputs(3301) <= b and not a;
    layer2_outputs(3302) <= not a or b;
    layer2_outputs(3303) <= a and not b;
    layer2_outputs(3304) <= a and b;
    layer2_outputs(3305) <= not (a and b);
    layer2_outputs(3306) <= not a or b;
    layer2_outputs(3307) <= not (a or b);
    layer2_outputs(3308) <= b;
    layer2_outputs(3309) <= not (a and b);
    layer2_outputs(3310) <= b;
    layer2_outputs(3311) <= a xor b;
    layer2_outputs(3312) <= not a;
    layer2_outputs(3313) <= a xor b;
    layer2_outputs(3314) <= not a;
    layer2_outputs(3315) <= a and b;
    layer2_outputs(3316) <= a or b;
    layer2_outputs(3317) <= not (a or b);
    layer2_outputs(3318) <= a;
    layer2_outputs(3319) <= not b;
    layer2_outputs(3320) <= a xor b;
    layer2_outputs(3321) <= not (a or b);
    layer2_outputs(3322) <= not a;
    layer2_outputs(3323) <= b and not a;
    layer2_outputs(3324) <= b;
    layer2_outputs(3325) <= b;
    layer2_outputs(3326) <= a or b;
    layer2_outputs(3327) <= not (a xor b);
    layer2_outputs(3328) <= not (a and b);
    layer2_outputs(3329) <= a;
    layer2_outputs(3330) <= not a or b;
    layer2_outputs(3331) <= not (a and b);
    layer2_outputs(3332) <= not a or b;
    layer2_outputs(3333) <= not (a and b);
    layer2_outputs(3334) <= a and not b;
    layer2_outputs(3335) <= a and not b;
    layer2_outputs(3336) <= not b;
    layer2_outputs(3337) <= not (a xor b);
    layer2_outputs(3338) <= not a;
    layer2_outputs(3339) <= not a;
    layer2_outputs(3340) <= a;
    layer2_outputs(3341) <= not a;
    layer2_outputs(3342) <= a;
    layer2_outputs(3343) <= not a;
    layer2_outputs(3344) <= not (a and b);
    layer2_outputs(3345) <= a and not b;
    layer2_outputs(3346) <= not b or a;
    layer2_outputs(3347) <= a and b;
    layer2_outputs(3348) <= not b;
    layer2_outputs(3349) <= not a;
    layer2_outputs(3350) <= a xor b;
    layer2_outputs(3351) <= a and b;
    layer2_outputs(3352) <= a;
    layer2_outputs(3353) <= a;
    layer2_outputs(3354) <= not a;
    layer2_outputs(3355) <= not (a and b);
    layer2_outputs(3356) <= a xor b;
    layer2_outputs(3357) <= a and not b;
    layer2_outputs(3358) <= a;
    layer2_outputs(3359) <= not (a xor b);
    layer2_outputs(3360) <= a and b;
    layer2_outputs(3361) <= not (a and b);
    layer2_outputs(3362) <= a xor b;
    layer2_outputs(3363) <= not b;
    layer2_outputs(3364) <= b;
    layer2_outputs(3365) <= not (a and b);
    layer2_outputs(3366) <= not (a or b);
    layer2_outputs(3367) <= a or b;
    layer2_outputs(3368) <= a and not b;
    layer2_outputs(3369) <= a and not b;
    layer2_outputs(3370) <= a or b;
    layer2_outputs(3371) <= a and not b;
    layer2_outputs(3372) <= a xor b;
    layer2_outputs(3373) <= not (a or b);
    layer2_outputs(3374) <= b and not a;
    layer2_outputs(3375) <= not b or a;
    layer2_outputs(3376) <= not a;
    layer2_outputs(3377) <= not b;
    layer2_outputs(3378) <= '0';
    layer2_outputs(3379) <= a;
    layer2_outputs(3380) <= a and b;
    layer2_outputs(3381) <= b;
    layer2_outputs(3382) <= not b or a;
    layer2_outputs(3383) <= not (a xor b);
    layer2_outputs(3384) <= not b;
    layer2_outputs(3385) <= a or b;
    layer2_outputs(3386) <= not a or b;
    layer2_outputs(3387) <= not (a or b);
    layer2_outputs(3388) <= a xor b;
    layer2_outputs(3389) <= not (a and b);
    layer2_outputs(3390) <= a;
    layer2_outputs(3391) <= a and not b;
    layer2_outputs(3392) <= not b;
    layer2_outputs(3393) <= b;
    layer2_outputs(3394) <= not (a or b);
    layer2_outputs(3395) <= not a or b;
    layer2_outputs(3396) <= a and b;
    layer2_outputs(3397) <= b;
    layer2_outputs(3398) <= a xor b;
    layer2_outputs(3399) <= a and b;
    layer2_outputs(3400) <= not a;
    layer2_outputs(3401) <= not (a xor b);
    layer2_outputs(3402) <= not a;
    layer2_outputs(3403) <= b;
    layer2_outputs(3404) <= not a;
    layer2_outputs(3405) <= not a;
    layer2_outputs(3406) <= not b;
    layer2_outputs(3407) <= not a;
    layer2_outputs(3408) <= a xor b;
    layer2_outputs(3409) <= a xor b;
    layer2_outputs(3410) <= not a;
    layer2_outputs(3411) <= not b;
    layer2_outputs(3412) <= not b or a;
    layer2_outputs(3413) <= not b;
    layer2_outputs(3414) <= a xor b;
    layer2_outputs(3415) <= b and not a;
    layer2_outputs(3416) <= a and b;
    layer2_outputs(3417) <= not (a or b);
    layer2_outputs(3418) <= not b or a;
    layer2_outputs(3419) <= a;
    layer2_outputs(3420) <= not a or b;
    layer2_outputs(3421) <= not b or a;
    layer2_outputs(3422) <= a xor b;
    layer2_outputs(3423) <= a or b;
    layer2_outputs(3424) <= a;
    layer2_outputs(3425) <= not (a and b);
    layer2_outputs(3426) <= not a or b;
    layer2_outputs(3427) <= not b;
    layer2_outputs(3428) <= a xor b;
    layer2_outputs(3429) <= a xor b;
    layer2_outputs(3430) <= not a;
    layer2_outputs(3431) <= '1';
    layer2_outputs(3432) <= not (a xor b);
    layer2_outputs(3433) <= b and not a;
    layer2_outputs(3434) <= not a;
    layer2_outputs(3435) <= not b or a;
    layer2_outputs(3436) <= not (a and b);
    layer2_outputs(3437) <= a xor b;
    layer2_outputs(3438) <= a;
    layer2_outputs(3439) <= b;
    layer2_outputs(3440) <= b;
    layer2_outputs(3441) <= not a;
    layer2_outputs(3442) <= b;
    layer2_outputs(3443) <= b and not a;
    layer2_outputs(3444) <= a and b;
    layer2_outputs(3445) <= not (a and b);
    layer2_outputs(3446) <= not a;
    layer2_outputs(3447) <= not a or b;
    layer2_outputs(3448) <= not b;
    layer2_outputs(3449) <= a xor b;
    layer2_outputs(3450) <= not a;
    layer2_outputs(3451) <= not a or b;
    layer2_outputs(3452) <= not a or b;
    layer2_outputs(3453) <= not (a or b);
    layer2_outputs(3454) <= not (a xor b);
    layer2_outputs(3455) <= not b or a;
    layer2_outputs(3456) <= b;
    layer2_outputs(3457) <= a or b;
    layer2_outputs(3458) <= not b or a;
    layer2_outputs(3459) <= not (a and b);
    layer2_outputs(3460) <= b and not a;
    layer2_outputs(3461) <= not (a and b);
    layer2_outputs(3462) <= not b or a;
    layer2_outputs(3463) <= b and not a;
    layer2_outputs(3464) <= not a;
    layer2_outputs(3465) <= not a;
    layer2_outputs(3466) <= not b;
    layer2_outputs(3467) <= not a;
    layer2_outputs(3468) <= a;
    layer2_outputs(3469) <= a and not b;
    layer2_outputs(3470) <= a xor b;
    layer2_outputs(3471) <= not b;
    layer2_outputs(3472) <= a xor b;
    layer2_outputs(3473) <= a;
    layer2_outputs(3474) <= not (a xor b);
    layer2_outputs(3475) <= not (a and b);
    layer2_outputs(3476) <= not a;
    layer2_outputs(3477) <= a xor b;
    layer2_outputs(3478) <= b and not a;
    layer2_outputs(3479) <= b;
    layer2_outputs(3480) <= a or b;
    layer2_outputs(3481) <= not a;
    layer2_outputs(3482) <= not b;
    layer2_outputs(3483) <= not b or a;
    layer2_outputs(3484) <= not a;
    layer2_outputs(3485) <= a and not b;
    layer2_outputs(3486) <= not b or a;
    layer2_outputs(3487) <= a xor b;
    layer2_outputs(3488) <= a;
    layer2_outputs(3489) <= b;
    layer2_outputs(3490) <= not (a xor b);
    layer2_outputs(3491) <= not (a xor b);
    layer2_outputs(3492) <= not (a xor b);
    layer2_outputs(3493) <= a;
    layer2_outputs(3494) <= not (a xor b);
    layer2_outputs(3495) <= a and not b;
    layer2_outputs(3496) <= not b;
    layer2_outputs(3497) <= a xor b;
    layer2_outputs(3498) <= a or b;
    layer2_outputs(3499) <= not (a and b);
    layer2_outputs(3500) <= b;
    layer2_outputs(3501) <= not b;
    layer2_outputs(3502) <= a xor b;
    layer2_outputs(3503) <= not b;
    layer2_outputs(3504) <= a and not b;
    layer2_outputs(3505) <= not (a or b);
    layer2_outputs(3506) <= a or b;
    layer2_outputs(3507) <= a;
    layer2_outputs(3508) <= not a or b;
    layer2_outputs(3509) <= a and not b;
    layer2_outputs(3510) <= b and not a;
    layer2_outputs(3511) <= a xor b;
    layer2_outputs(3512) <= a xor b;
    layer2_outputs(3513) <= not b;
    layer2_outputs(3514) <= b;
    layer2_outputs(3515) <= a and not b;
    layer2_outputs(3516) <= not (a or b);
    layer2_outputs(3517) <= not b or a;
    layer2_outputs(3518) <= not b;
    layer2_outputs(3519) <= not b;
    layer2_outputs(3520) <= not b;
    layer2_outputs(3521) <= not b or a;
    layer2_outputs(3522) <= not a;
    layer2_outputs(3523) <= a xor b;
    layer2_outputs(3524) <= a xor b;
    layer2_outputs(3525) <= not (a and b);
    layer2_outputs(3526) <= not b or a;
    layer2_outputs(3527) <= a or b;
    layer2_outputs(3528) <= not a;
    layer2_outputs(3529) <= b and not a;
    layer2_outputs(3530) <= not (a or b);
    layer2_outputs(3531) <= a;
    layer2_outputs(3532) <= b;
    layer2_outputs(3533) <= not (a or b);
    layer2_outputs(3534) <= not (a xor b);
    layer2_outputs(3535) <= not b or a;
    layer2_outputs(3536) <= a;
    layer2_outputs(3537) <= not a;
    layer2_outputs(3538) <= not b;
    layer2_outputs(3539) <= not a;
    layer2_outputs(3540) <= b;
    layer2_outputs(3541) <= b and not a;
    layer2_outputs(3542) <= a and b;
    layer2_outputs(3543) <= not a;
    layer2_outputs(3544) <= not a;
    layer2_outputs(3545) <= b;
    layer2_outputs(3546) <= not b;
    layer2_outputs(3547) <= b and not a;
    layer2_outputs(3548) <= not (a or b);
    layer2_outputs(3549) <= not (a and b);
    layer2_outputs(3550) <= a or b;
    layer2_outputs(3551) <= not b or a;
    layer2_outputs(3552) <= b;
    layer2_outputs(3553) <= not (a and b);
    layer2_outputs(3554) <= a and b;
    layer2_outputs(3555) <= a;
    layer2_outputs(3556) <= not b or a;
    layer2_outputs(3557) <= not (a xor b);
    layer2_outputs(3558) <= not b;
    layer2_outputs(3559) <= not a;
    layer2_outputs(3560) <= a and not b;
    layer2_outputs(3561) <= not a;
    layer2_outputs(3562) <= a and b;
    layer2_outputs(3563) <= a xor b;
    layer2_outputs(3564) <= b;
    layer2_outputs(3565) <= not a;
    layer2_outputs(3566) <= a xor b;
    layer2_outputs(3567) <= not a;
    layer2_outputs(3568) <= a xor b;
    layer2_outputs(3569) <= not a;
    layer2_outputs(3570) <= not a;
    layer2_outputs(3571) <= not (a xor b);
    layer2_outputs(3572) <= b;
    layer2_outputs(3573) <= a xor b;
    layer2_outputs(3574) <= a or b;
    layer2_outputs(3575) <= not (a or b);
    layer2_outputs(3576) <= not b;
    layer2_outputs(3577) <= not (a or b);
    layer2_outputs(3578) <= not a;
    layer2_outputs(3579) <= a xor b;
    layer2_outputs(3580) <= a or b;
    layer2_outputs(3581) <= b;
    layer2_outputs(3582) <= a and b;
    layer2_outputs(3583) <= not b;
    layer2_outputs(3584) <= not (a xor b);
    layer2_outputs(3585) <= not (a or b);
    layer2_outputs(3586) <= not b or a;
    layer2_outputs(3587) <= '1';
    layer2_outputs(3588) <= a and not b;
    layer2_outputs(3589) <= a;
    layer2_outputs(3590) <= a xor b;
    layer2_outputs(3591) <= not a;
    layer2_outputs(3592) <= a and not b;
    layer2_outputs(3593) <= not a;
    layer2_outputs(3594) <= not a;
    layer2_outputs(3595) <= a and not b;
    layer2_outputs(3596) <= a or b;
    layer2_outputs(3597) <= a and not b;
    layer2_outputs(3598) <= not a;
    layer2_outputs(3599) <= not (a xor b);
    layer2_outputs(3600) <= not b;
    layer2_outputs(3601) <= a or b;
    layer2_outputs(3602) <= '1';
    layer2_outputs(3603) <= b and not a;
    layer2_outputs(3604) <= not a;
    layer2_outputs(3605) <= a xor b;
    layer2_outputs(3606) <= a and b;
    layer2_outputs(3607) <= a xor b;
    layer2_outputs(3608) <= not b or a;
    layer2_outputs(3609) <= b;
    layer2_outputs(3610) <= a and b;
    layer2_outputs(3611) <= b and not a;
    layer2_outputs(3612) <= not (a xor b);
    layer2_outputs(3613) <= a and b;
    layer2_outputs(3614) <= not a;
    layer2_outputs(3615) <= not (a or b);
    layer2_outputs(3616) <= a xor b;
    layer2_outputs(3617) <= b;
    layer2_outputs(3618) <= not (a xor b);
    layer2_outputs(3619) <= not (a xor b);
    layer2_outputs(3620) <= not (a and b);
    layer2_outputs(3621) <= not (a xor b);
    layer2_outputs(3622) <= a;
    layer2_outputs(3623) <= not a;
    layer2_outputs(3624) <= a;
    layer2_outputs(3625) <= not (a or b);
    layer2_outputs(3626) <= a and b;
    layer2_outputs(3627) <= a or b;
    layer2_outputs(3628) <= not b;
    layer2_outputs(3629) <= not b or a;
    layer2_outputs(3630) <= b;
    layer2_outputs(3631) <= not b or a;
    layer2_outputs(3632) <= b;
    layer2_outputs(3633) <= a and not b;
    layer2_outputs(3634) <= not b;
    layer2_outputs(3635) <= a and not b;
    layer2_outputs(3636) <= b and not a;
    layer2_outputs(3637) <= not b;
    layer2_outputs(3638) <= not a;
    layer2_outputs(3639) <= not (a xor b);
    layer2_outputs(3640) <= a or b;
    layer2_outputs(3641) <= a or b;
    layer2_outputs(3642) <= '0';
    layer2_outputs(3643) <= not (a or b);
    layer2_outputs(3644) <= not (a or b);
    layer2_outputs(3645) <= a and not b;
    layer2_outputs(3646) <= a xor b;
    layer2_outputs(3647) <= not b or a;
    layer2_outputs(3648) <= not a;
    layer2_outputs(3649) <= not b;
    layer2_outputs(3650) <= a xor b;
    layer2_outputs(3651) <= b;
    layer2_outputs(3652) <= b;
    layer2_outputs(3653) <= not (a and b);
    layer2_outputs(3654) <= not a;
    layer2_outputs(3655) <= not b;
    layer2_outputs(3656) <= b;
    layer2_outputs(3657) <= a and b;
    layer2_outputs(3658) <= a or b;
    layer2_outputs(3659) <= not (a and b);
    layer2_outputs(3660) <= not a or b;
    layer2_outputs(3661) <= not (a or b);
    layer2_outputs(3662) <= not b;
    layer2_outputs(3663) <= not (a and b);
    layer2_outputs(3664) <= a;
    layer2_outputs(3665) <= a;
    layer2_outputs(3666) <= a or b;
    layer2_outputs(3667) <= a xor b;
    layer2_outputs(3668) <= not (a or b);
    layer2_outputs(3669) <= b;
    layer2_outputs(3670) <= not b;
    layer2_outputs(3671) <= a;
    layer2_outputs(3672) <= not b;
    layer2_outputs(3673) <= not b;
    layer2_outputs(3674) <= b and not a;
    layer2_outputs(3675) <= not (a or b);
    layer2_outputs(3676) <= not (a xor b);
    layer2_outputs(3677) <= not a;
    layer2_outputs(3678) <= not (a or b);
    layer2_outputs(3679) <= a xor b;
    layer2_outputs(3680) <= b and not a;
    layer2_outputs(3681) <= not b;
    layer2_outputs(3682) <= not a;
    layer2_outputs(3683) <= a and b;
    layer2_outputs(3684) <= not (a xor b);
    layer2_outputs(3685) <= not (a and b);
    layer2_outputs(3686) <= a or b;
    layer2_outputs(3687) <= not a;
    layer2_outputs(3688) <= not b;
    layer2_outputs(3689) <= a and not b;
    layer2_outputs(3690) <= a;
    layer2_outputs(3691) <= a xor b;
    layer2_outputs(3692) <= not (a or b);
    layer2_outputs(3693) <= b;
    layer2_outputs(3694) <= b;
    layer2_outputs(3695) <= not (a xor b);
    layer2_outputs(3696) <= not a;
    layer2_outputs(3697) <= not b;
    layer2_outputs(3698) <= not (a and b);
    layer2_outputs(3699) <= not b or a;
    layer2_outputs(3700) <= b and not a;
    layer2_outputs(3701) <= a xor b;
    layer2_outputs(3702) <= a or b;
    layer2_outputs(3703) <= not b or a;
    layer2_outputs(3704) <= not a or b;
    layer2_outputs(3705) <= not a or b;
    layer2_outputs(3706) <= b and not a;
    layer2_outputs(3707) <= a xor b;
    layer2_outputs(3708) <= not b or a;
    layer2_outputs(3709) <= not a;
    layer2_outputs(3710) <= not a;
    layer2_outputs(3711) <= not (a or b);
    layer2_outputs(3712) <= not (a or b);
    layer2_outputs(3713) <= not b;
    layer2_outputs(3714) <= not (a and b);
    layer2_outputs(3715) <= not a;
    layer2_outputs(3716) <= not a;
    layer2_outputs(3717) <= not b;
    layer2_outputs(3718) <= b;
    layer2_outputs(3719) <= not (a and b);
    layer2_outputs(3720) <= not a or b;
    layer2_outputs(3721) <= not a;
    layer2_outputs(3722) <= not (a xor b);
    layer2_outputs(3723) <= a;
    layer2_outputs(3724) <= not (a xor b);
    layer2_outputs(3725) <= b;
    layer2_outputs(3726) <= a xor b;
    layer2_outputs(3727) <= a;
    layer2_outputs(3728) <= a or b;
    layer2_outputs(3729) <= not b or a;
    layer2_outputs(3730) <= b and not a;
    layer2_outputs(3731) <= a and not b;
    layer2_outputs(3732) <= a;
    layer2_outputs(3733) <= b;
    layer2_outputs(3734) <= not a;
    layer2_outputs(3735) <= not (a and b);
    layer2_outputs(3736) <= not a;
    layer2_outputs(3737) <= not a or b;
    layer2_outputs(3738) <= not a;
    layer2_outputs(3739) <= a;
    layer2_outputs(3740) <= not (a or b);
    layer2_outputs(3741) <= not b;
    layer2_outputs(3742) <= not (a or b);
    layer2_outputs(3743) <= b;
    layer2_outputs(3744) <= not b;
    layer2_outputs(3745) <= not (a or b);
    layer2_outputs(3746) <= a and b;
    layer2_outputs(3747) <= b;
    layer2_outputs(3748) <= not b;
    layer2_outputs(3749) <= a or b;
    layer2_outputs(3750) <= not b;
    layer2_outputs(3751) <= not b;
    layer2_outputs(3752) <= not b;
    layer2_outputs(3753) <= a xor b;
    layer2_outputs(3754) <= a or b;
    layer2_outputs(3755) <= not (a xor b);
    layer2_outputs(3756) <= a;
    layer2_outputs(3757) <= not (a xor b);
    layer2_outputs(3758) <= not a;
    layer2_outputs(3759) <= a and not b;
    layer2_outputs(3760) <= a;
    layer2_outputs(3761) <= not b;
    layer2_outputs(3762) <= not b;
    layer2_outputs(3763) <= not (a xor b);
    layer2_outputs(3764) <= a;
    layer2_outputs(3765) <= b and not a;
    layer2_outputs(3766) <= not (a or b);
    layer2_outputs(3767) <= not b;
    layer2_outputs(3768) <= b;
    layer2_outputs(3769) <= a and b;
    layer2_outputs(3770) <= a xor b;
    layer2_outputs(3771) <= a;
    layer2_outputs(3772) <= b;
    layer2_outputs(3773) <= not b or a;
    layer2_outputs(3774) <= not (a and b);
    layer2_outputs(3775) <= a xor b;
    layer2_outputs(3776) <= a xor b;
    layer2_outputs(3777) <= not (a and b);
    layer2_outputs(3778) <= not a;
    layer2_outputs(3779) <= not b;
    layer2_outputs(3780) <= a xor b;
    layer2_outputs(3781) <= a;
    layer2_outputs(3782) <= a and b;
    layer2_outputs(3783) <= not (a xor b);
    layer2_outputs(3784) <= a xor b;
    layer2_outputs(3785) <= not (a or b);
    layer2_outputs(3786) <= a and b;
    layer2_outputs(3787) <= a xor b;
    layer2_outputs(3788) <= a xor b;
    layer2_outputs(3789) <= not b or a;
    layer2_outputs(3790) <= not b;
    layer2_outputs(3791) <= b;
    layer2_outputs(3792) <= b;
    layer2_outputs(3793) <= '0';
    layer2_outputs(3794) <= not a;
    layer2_outputs(3795) <= not b;
    layer2_outputs(3796) <= not (a and b);
    layer2_outputs(3797) <= not (a and b);
    layer2_outputs(3798) <= a;
    layer2_outputs(3799) <= not a or b;
    layer2_outputs(3800) <= a;
    layer2_outputs(3801) <= a xor b;
    layer2_outputs(3802) <= not b or a;
    layer2_outputs(3803) <= not a;
    layer2_outputs(3804) <= not b;
    layer2_outputs(3805) <= not a;
    layer2_outputs(3806) <= a and not b;
    layer2_outputs(3807) <= b;
    layer2_outputs(3808) <= b;
    layer2_outputs(3809) <= a;
    layer2_outputs(3810) <= not (a or b);
    layer2_outputs(3811) <= not (a or b);
    layer2_outputs(3812) <= not (a xor b);
    layer2_outputs(3813) <= a xor b;
    layer2_outputs(3814) <= a;
    layer2_outputs(3815) <= not a or b;
    layer2_outputs(3816) <= not a;
    layer2_outputs(3817) <= not a;
    layer2_outputs(3818) <= b;
    layer2_outputs(3819) <= a;
    layer2_outputs(3820) <= a xor b;
    layer2_outputs(3821) <= b;
    layer2_outputs(3822) <= a and b;
    layer2_outputs(3823) <= a and not b;
    layer2_outputs(3824) <= not b;
    layer2_outputs(3825) <= '1';
    layer2_outputs(3826) <= not a;
    layer2_outputs(3827) <= b;
    layer2_outputs(3828) <= not a or b;
    layer2_outputs(3829) <= not a;
    layer2_outputs(3830) <= '0';
    layer2_outputs(3831) <= not (a xor b);
    layer2_outputs(3832) <= not b;
    layer2_outputs(3833) <= b;
    layer2_outputs(3834) <= not a;
    layer2_outputs(3835) <= not b or a;
    layer2_outputs(3836) <= not b;
    layer2_outputs(3837) <= a;
    layer2_outputs(3838) <= a;
    layer2_outputs(3839) <= not (a or b);
    layer2_outputs(3840) <= not (a xor b);
    layer2_outputs(3841) <= a xor b;
    layer2_outputs(3842) <= b and not a;
    layer2_outputs(3843) <= a xor b;
    layer2_outputs(3844) <= not b;
    layer2_outputs(3845) <= a xor b;
    layer2_outputs(3846) <= not a;
    layer2_outputs(3847) <= not a;
    layer2_outputs(3848) <= not a;
    layer2_outputs(3849) <= not b;
    layer2_outputs(3850) <= not a;
    layer2_outputs(3851) <= not a;
    layer2_outputs(3852) <= not a or b;
    layer2_outputs(3853) <= not (a or b);
    layer2_outputs(3854) <= a xor b;
    layer2_outputs(3855) <= not (a and b);
    layer2_outputs(3856) <= a and not b;
    layer2_outputs(3857) <= b;
    layer2_outputs(3858) <= not a;
    layer2_outputs(3859) <= b and not a;
    layer2_outputs(3860) <= b;
    layer2_outputs(3861) <= not a;
    layer2_outputs(3862) <= not (a and b);
    layer2_outputs(3863) <= not (a xor b);
    layer2_outputs(3864) <= a or b;
    layer2_outputs(3865) <= not (a or b);
    layer2_outputs(3866) <= not b;
    layer2_outputs(3867) <= not b or a;
    layer2_outputs(3868) <= a xor b;
    layer2_outputs(3869) <= a;
    layer2_outputs(3870) <= '1';
    layer2_outputs(3871) <= not b;
    layer2_outputs(3872) <= a;
    layer2_outputs(3873) <= not b;
    layer2_outputs(3874) <= not a;
    layer2_outputs(3875) <= a and b;
    layer2_outputs(3876) <= not (a or b);
    layer2_outputs(3877) <= a and not b;
    layer2_outputs(3878) <= a;
    layer2_outputs(3879) <= not (a xor b);
    layer2_outputs(3880) <= not b;
    layer2_outputs(3881) <= not b or a;
    layer2_outputs(3882) <= not a;
    layer2_outputs(3883) <= not b;
    layer2_outputs(3884) <= not (a and b);
    layer2_outputs(3885) <= b;
    layer2_outputs(3886) <= a xor b;
    layer2_outputs(3887) <= not (a or b);
    layer2_outputs(3888) <= not a or b;
    layer2_outputs(3889) <= not (a or b);
    layer2_outputs(3890) <= not (a xor b);
    layer2_outputs(3891) <= not a;
    layer2_outputs(3892) <= not a;
    layer2_outputs(3893) <= b;
    layer2_outputs(3894) <= a xor b;
    layer2_outputs(3895) <= not (a xor b);
    layer2_outputs(3896) <= a xor b;
    layer2_outputs(3897) <= a and b;
    layer2_outputs(3898) <= a or b;
    layer2_outputs(3899) <= a;
    layer2_outputs(3900) <= not b;
    layer2_outputs(3901) <= a;
    layer2_outputs(3902) <= a xor b;
    layer2_outputs(3903) <= not (a xor b);
    layer2_outputs(3904) <= b and not a;
    layer2_outputs(3905) <= not b;
    layer2_outputs(3906) <= not a;
    layer2_outputs(3907) <= b and not a;
    layer2_outputs(3908) <= not (a xor b);
    layer2_outputs(3909) <= not a or b;
    layer2_outputs(3910) <= not (a or b);
    layer2_outputs(3911) <= not b;
    layer2_outputs(3912) <= not (a or b);
    layer2_outputs(3913) <= a and b;
    layer2_outputs(3914) <= a or b;
    layer2_outputs(3915) <= a;
    layer2_outputs(3916) <= not a;
    layer2_outputs(3917) <= not b;
    layer2_outputs(3918) <= not (a xor b);
    layer2_outputs(3919) <= not (a and b);
    layer2_outputs(3920) <= not (a xor b);
    layer2_outputs(3921) <= not (a xor b);
    layer2_outputs(3922) <= a xor b;
    layer2_outputs(3923) <= not (a xor b);
    layer2_outputs(3924) <= b;
    layer2_outputs(3925) <= not b;
    layer2_outputs(3926) <= b;
    layer2_outputs(3927) <= b;
    layer2_outputs(3928) <= not a;
    layer2_outputs(3929) <= not b or a;
    layer2_outputs(3930) <= not (a xor b);
    layer2_outputs(3931) <= not b or a;
    layer2_outputs(3932) <= a;
    layer2_outputs(3933) <= not a;
    layer2_outputs(3934) <= a;
    layer2_outputs(3935) <= a and not b;
    layer2_outputs(3936) <= a;
    layer2_outputs(3937) <= a or b;
    layer2_outputs(3938) <= a and b;
    layer2_outputs(3939) <= not a;
    layer2_outputs(3940) <= b and not a;
    layer2_outputs(3941) <= a xor b;
    layer2_outputs(3942) <= not a;
    layer2_outputs(3943) <= not (a xor b);
    layer2_outputs(3944) <= not (a or b);
    layer2_outputs(3945) <= b;
    layer2_outputs(3946) <= b;
    layer2_outputs(3947) <= b;
    layer2_outputs(3948) <= b and not a;
    layer2_outputs(3949) <= a;
    layer2_outputs(3950) <= a xor b;
    layer2_outputs(3951) <= not (a xor b);
    layer2_outputs(3952) <= not (a or b);
    layer2_outputs(3953) <= not (a and b);
    layer2_outputs(3954) <= not b or a;
    layer2_outputs(3955) <= a and b;
    layer2_outputs(3956) <= a xor b;
    layer2_outputs(3957) <= b;
    layer2_outputs(3958) <= not (a or b);
    layer2_outputs(3959) <= b;
    layer2_outputs(3960) <= not b or a;
    layer2_outputs(3961) <= not b or a;
    layer2_outputs(3962) <= not a or b;
    layer2_outputs(3963) <= a xor b;
    layer2_outputs(3964) <= a and b;
    layer2_outputs(3965) <= b;
    layer2_outputs(3966) <= b;
    layer2_outputs(3967) <= not (a xor b);
    layer2_outputs(3968) <= not (a xor b);
    layer2_outputs(3969) <= not (a and b);
    layer2_outputs(3970) <= a and not b;
    layer2_outputs(3971) <= a and b;
    layer2_outputs(3972) <= b;
    layer2_outputs(3973) <= a and b;
    layer2_outputs(3974) <= b and not a;
    layer2_outputs(3975) <= not b;
    layer2_outputs(3976) <= a;
    layer2_outputs(3977) <= not b or a;
    layer2_outputs(3978) <= a or b;
    layer2_outputs(3979) <= not b;
    layer2_outputs(3980) <= not b;
    layer2_outputs(3981) <= a;
    layer2_outputs(3982) <= a;
    layer2_outputs(3983) <= a;
    layer2_outputs(3984) <= not (a xor b);
    layer2_outputs(3985) <= not a;
    layer2_outputs(3986) <= not a;
    layer2_outputs(3987) <= not (a and b);
    layer2_outputs(3988) <= not b;
    layer2_outputs(3989) <= not b;
    layer2_outputs(3990) <= a;
    layer2_outputs(3991) <= a;
    layer2_outputs(3992) <= not (a xor b);
    layer2_outputs(3993) <= a and not b;
    layer2_outputs(3994) <= not b;
    layer2_outputs(3995) <= not a;
    layer2_outputs(3996) <= a or b;
    layer2_outputs(3997) <= b;
    layer2_outputs(3998) <= a and not b;
    layer2_outputs(3999) <= not a;
    layer2_outputs(4000) <= a xor b;
    layer2_outputs(4001) <= b;
    layer2_outputs(4002) <= not b;
    layer2_outputs(4003) <= not a or b;
    layer2_outputs(4004) <= not (a or b);
    layer2_outputs(4005) <= a xor b;
    layer2_outputs(4006) <= '0';
    layer2_outputs(4007) <= not b;
    layer2_outputs(4008) <= b;
    layer2_outputs(4009) <= a xor b;
    layer2_outputs(4010) <= b and not a;
    layer2_outputs(4011) <= a and not b;
    layer2_outputs(4012) <= a;
    layer2_outputs(4013) <= not (a xor b);
    layer2_outputs(4014) <= a and not b;
    layer2_outputs(4015) <= not b;
    layer2_outputs(4016) <= not b or a;
    layer2_outputs(4017) <= a or b;
    layer2_outputs(4018) <= b;
    layer2_outputs(4019) <= b and not a;
    layer2_outputs(4020) <= b;
    layer2_outputs(4021) <= not b;
    layer2_outputs(4022) <= b;
    layer2_outputs(4023) <= not b;
    layer2_outputs(4024) <= a;
    layer2_outputs(4025) <= not (a xor b);
    layer2_outputs(4026) <= not a or b;
    layer2_outputs(4027) <= not a or b;
    layer2_outputs(4028) <= b;
    layer2_outputs(4029) <= not (a and b);
    layer2_outputs(4030) <= a;
    layer2_outputs(4031) <= not (a xor b);
    layer2_outputs(4032) <= a or b;
    layer2_outputs(4033) <= b;
    layer2_outputs(4034) <= a or b;
    layer2_outputs(4035) <= not (a xor b);
    layer2_outputs(4036) <= a xor b;
    layer2_outputs(4037) <= not b or a;
    layer2_outputs(4038) <= not (a and b);
    layer2_outputs(4039) <= not b or a;
    layer2_outputs(4040) <= not b or a;
    layer2_outputs(4041) <= not b;
    layer2_outputs(4042) <= not b;
    layer2_outputs(4043) <= a and b;
    layer2_outputs(4044) <= a or b;
    layer2_outputs(4045) <= a;
    layer2_outputs(4046) <= not (a xor b);
    layer2_outputs(4047) <= not b or a;
    layer2_outputs(4048) <= not a;
    layer2_outputs(4049) <= not a or b;
    layer2_outputs(4050) <= b and not a;
    layer2_outputs(4051) <= a xor b;
    layer2_outputs(4052) <= a;
    layer2_outputs(4053) <= a;
    layer2_outputs(4054) <= not (a xor b);
    layer2_outputs(4055) <= a and b;
    layer2_outputs(4056) <= a xor b;
    layer2_outputs(4057) <= a xor b;
    layer2_outputs(4058) <= not a;
    layer2_outputs(4059) <= not (a xor b);
    layer2_outputs(4060) <= b;
    layer2_outputs(4061) <= a;
    layer2_outputs(4062) <= not a;
    layer2_outputs(4063) <= b;
    layer2_outputs(4064) <= a or b;
    layer2_outputs(4065) <= b;
    layer2_outputs(4066) <= b;
    layer2_outputs(4067) <= b;
    layer2_outputs(4068) <= a and b;
    layer2_outputs(4069) <= not b or a;
    layer2_outputs(4070) <= not (a xor b);
    layer2_outputs(4071) <= a and b;
    layer2_outputs(4072) <= not b or a;
    layer2_outputs(4073) <= a xor b;
    layer2_outputs(4074) <= b;
    layer2_outputs(4075) <= not b;
    layer2_outputs(4076) <= not b or a;
    layer2_outputs(4077) <= not b or a;
    layer2_outputs(4078) <= not a;
    layer2_outputs(4079) <= not b;
    layer2_outputs(4080) <= not a or b;
    layer2_outputs(4081) <= not a or b;
    layer2_outputs(4082) <= not a or b;
    layer2_outputs(4083) <= a or b;
    layer2_outputs(4084) <= a;
    layer2_outputs(4085) <= not (a and b);
    layer2_outputs(4086) <= not (a xor b);
    layer2_outputs(4087) <= not a;
    layer2_outputs(4088) <= b and not a;
    layer2_outputs(4089) <= '0';
    layer2_outputs(4090) <= b;
    layer2_outputs(4091) <= not b;
    layer2_outputs(4092) <= not (a or b);
    layer2_outputs(4093) <= b;
    layer2_outputs(4094) <= a or b;
    layer2_outputs(4095) <= not b;
    layer2_outputs(4096) <= b and not a;
    layer2_outputs(4097) <= not b or a;
    layer2_outputs(4098) <= a or b;
    layer2_outputs(4099) <= a xor b;
    layer2_outputs(4100) <= not (a or b);
    layer2_outputs(4101) <= not (a xor b);
    layer2_outputs(4102) <= not (a and b);
    layer2_outputs(4103) <= b;
    layer2_outputs(4104) <= not (a or b);
    layer2_outputs(4105) <= not a;
    layer2_outputs(4106) <= b;
    layer2_outputs(4107) <= a;
    layer2_outputs(4108) <= a xor b;
    layer2_outputs(4109) <= not a;
    layer2_outputs(4110) <= a and b;
    layer2_outputs(4111) <= a and not b;
    layer2_outputs(4112) <= a and b;
    layer2_outputs(4113) <= a xor b;
    layer2_outputs(4114) <= a xor b;
    layer2_outputs(4115) <= not b;
    layer2_outputs(4116) <= a xor b;
    layer2_outputs(4117) <= a or b;
    layer2_outputs(4118) <= a;
    layer2_outputs(4119) <= a xor b;
    layer2_outputs(4120) <= not b or a;
    layer2_outputs(4121) <= a xor b;
    layer2_outputs(4122) <= a;
    layer2_outputs(4123) <= not a;
    layer2_outputs(4124) <= a;
    layer2_outputs(4125) <= not (a and b);
    layer2_outputs(4126) <= a and not b;
    layer2_outputs(4127) <= b and not a;
    layer2_outputs(4128) <= not (a and b);
    layer2_outputs(4129) <= a and b;
    layer2_outputs(4130) <= not a or b;
    layer2_outputs(4131) <= not b;
    layer2_outputs(4132) <= not (a and b);
    layer2_outputs(4133) <= not a;
    layer2_outputs(4134) <= not a or b;
    layer2_outputs(4135) <= a xor b;
    layer2_outputs(4136) <= b and not a;
    layer2_outputs(4137) <= not a;
    layer2_outputs(4138) <= a xor b;
    layer2_outputs(4139) <= not (a and b);
    layer2_outputs(4140) <= a;
    layer2_outputs(4141) <= not b;
    layer2_outputs(4142) <= not a or b;
    layer2_outputs(4143) <= not (a or b);
    layer2_outputs(4144) <= not b;
    layer2_outputs(4145) <= not (a or b);
    layer2_outputs(4146) <= not b;
    layer2_outputs(4147) <= not (a and b);
    layer2_outputs(4148) <= not (a or b);
    layer2_outputs(4149) <= a;
    layer2_outputs(4150) <= a and b;
    layer2_outputs(4151) <= not (a xor b);
    layer2_outputs(4152) <= a xor b;
    layer2_outputs(4153) <= a or b;
    layer2_outputs(4154) <= not b;
    layer2_outputs(4155) <= not (a or b);
    layer2_outputs(4156) <= not b;
    layer2_outputs(4157) <= not a;
    layer2_outputs(4158) <= a and b;
    layer2_outputs(4159) <= not a;
    layer2_outputs(4160) <= b;
    layer2_outputs(4161) <= not (a or b);
    layer2_outputs(4162) <= a or b;
    layer2_outputs(4163) <= not b;
    layer2_outputs(4164) <= not (a or b);
    layer2_outputs(4165) <= a xor b;
    layer2_outputs(4166) <= not a;
    layer2_outputs(4167) <= not a;
    layer2_outputs(4168) <= not (a or b);
    layer2_outputs(4169) <= a xor b;
    layer2_outputs(4170) <= b;
    layer2_outputs(4171) <= a xor b;
    layer2_outputs(4172) <= b and not a;
    layer2_outputs(4173) <= a or b;
    layer2_outputs(4174) <= not a;
    layer2_outputs(4175) <= b and not a;
    layer2_outputs(4176) <= not b;
    layer2_outputs(4177) <= a xor b;
    layer2_outputs(4178) <= b;
    layer2_outputs(4179) <= a and not b;
    layer2_outputs(4180) <= not (a and b);
    layer2_outputs(4181) <= a;
    layer2_outputs(4182) <= not a or b;
    layer2_outputs(4183) <= a and not b;
    layer2_outputs(4184) <= a and not b;
    layer2_outputs(4185) <= b;
    layer2_outputs(4186) <= not a or b;
    layer2_outputs(4187) <= not a;
    layer2_outputs(4188) <= '0';
    layer2_outputs(4189) <= not (a or b);
    layer2_outputs(4190) <= a xor b;
    layer2_outputs(4191) <= not (a or b);
    layer2_outputs(4192) <= not (a or b);
    layer2_outputs(4193) <= not (a xor b);
    layer2_outputs(4194) <= not (a or b);
    layer2_outputs(4195) <= b and not a;
    layer2_outputs(4196) <= a xor b;
    layer2_outputs(4197) <= not (a xor b);
    layer2_outputs(4198) <= b and not a;
    layer2_outputs(4199) <= a;
    layer2_outputs(4200) <= b;
    layer2_outputs(4201) <= b;
    layer2_outputs(4202) <= not a;
    layer2_outputs(4203) <= b;
    layer2_outputs(4204) <= a and b;
    layer2_outputs(4205) <= not (a or b);
    layer2_outputs(4206) <= not (a xor b);
    layer2_outputs(4207) <= a or b;
    layer2_outputs(4208) <= not b;
    layer2_outputs(4209) <= a and b;
    layer2_outputs(4210) <= not a;
    layer2_outputs(4211) <= a xor b;
    layer2_outputs(4212) <= not b or a;
    layer2_outputs(4213) <= not a;
    layer2_outputs(4214) <= a;
    layer2_outputs(4215) <= a xor b;
    layer2_outputs(4216) <= not b;
    layer2_outputs(4217) <= b;
    layer2_outputs(4218) <= b and not a;
    layer2_outputs(4219) <= not b;
    layer2_outputs(4220) <= not (a xor b);
    layer2_outputs(4221) <= not b or a;
    layer2_outputs(4222) <= a and not b;
    layer2_outputs(4223) <= not (a or b);
    layer2_outputs(4224) <= b;
    layer2_outputs(4225) <= not a;
    layer2_outputs(4226) <= a and not b;
    layer2_outputs(4227) <= not b or a;
    layer2_outputs(4228) <= a;
    layer2_outputs(4229) <= not a;
    layer2_outputs(4230) <= not (a xor b);
    layer2_outputs(4231) <= not (a xor b);
    layer2_outputs(4232) <= not (a or b);
    layer2_outputs(4233) <= not a or b;
    layer2_outputs(4234) <= not a or b;
    layer2_outputs(4235) <= not a;
    layer2_outputs(4236) <= b and not a;
    layer2_outputs(4237) <= not (a xor b);
    layer2_outputs(4238) <= a and not b;
    layer2_outputs(4239) <= a and not b;
    layer2_outputs(4240) <= a;
    layer2_outputs(4241) <= not (a or b);
    layer2_outputs(4242) <= not (a or b);
    layer2_outputs(4243) <= a;
    layer2_outputs(4244) <= not a or b;
    layer2_outputs(4245) <= a and not b;
    layer2_outputs(4246) <= not a;
    layer2_outputs(4247) <= a;
    layer2_outputs(4248) <= a and b;
    layer2_outputs(4249) <= b;
    layer2_outputs(4250) <= not (a xor b);
    layer2_outputs(4251) <= not a;
    layer2_outputs(4252) <= not a or b;
    layer2_outputs(4253) <= not a or b;
    layer2_outputs(4254) <= not a or b;
    layer2_outputs(4255) <= not (a and b);
    layer2_outputs(4256) <= not a;
    layer2_outputs(4257) <= not (a or b);
    layer2_outputs(4258) <= a;
    layer2_outputs(4259) <= not a;
    layer2_outputs(4260) <= not b;
    layer2_outputs(4261) <= a;
    layer2_outputs(4262) <= not (a xor b);
    layer2_outputs(4263) <= a;
    layer2_outputs(4264) <= not a;
    layer2_outputs(4265) <= not (a xor b);
    layer2_outputs(4266) <= not b;
    layer2_outputs(4267) <= not b;
    layer2_outputs(4268) <= not (a and b);
    layer2_outputs(4269) <= a xor b;
    layer2_outputs(4270) <= not b;
    layer2_outputs(4271) <= a xor b;
    layer2_outputs(4272) <= b;
    layer2_outputs(4273) <= b and not a;
    layer2_outputs(4274) <= not a;
    layer2_outputs(4275) <= not (a and b);
    layer2_outputs(4276) <= a and b;
    layer2_outputs(4277) <= not (a xor b);
    layer2_outputs(4278) <= not b or a;
    layer2_outputs(4279) <= a and b;
    layer2_outputs(4280) <= not b;
    layer2_outputs(4281) <= a and not b;
    layer2_outputs(4282) <= not a;
    layer2_outputs(4283) <= not (a xor b);
    layer2_outputs(4284) <= not a;
    layer2_outputs(4285) <= a xor b;
    layer2_outputs(4286) <= '1';
    layer2_outputs(4287) <= not (a and b);
    layer2_outputs(4288) <= not b;
    layer2_outputs(4289) <= a xor b;
    layer2_outputs(4290) <= b;
    layer2_outputs(4291) <= a xor b;
    layer2_outputs(4292) <= not b;
    layer2_outputs(4293) <= not b or a;
    layer2_outputs(4294) <= b and not a;
    layer2_outputs(4295) <= not a;
    layer2_outputs(4296) <= not (a xor b);
    layer2_outputs(4297) <= not (a or b);
    layer2_outputs(4298) <= not b;
    layer2_outputs(4299) <= not a;
    layer2_outputs(4300) <= b;
    layer2_outputs(4301) <= a;
    layer2_outputs(4302) <= a;
    layer2_outputs(4303) <= a and b;
    layer2_outputs(4304) <= not (a or b);
    layer2_outputs(4305) <= not (a or b);
    layer2_outputs(4306) <= not (a or b);
    layer2_outputs(4307) <= a and not b;
    layer2_outputs(4308) <= not b;
    layer2_outputs(4309) <= not b;
    layer2_outputs(4310) <= b;
    layer2_outputs(4311) <= a;
    layer2_outputs(4312) <= not (a xor b);
    layer2_outputs(4313) <= a and not b;
    layer2_outputs(4314) <= a;
    layer2_outputs(4315) <= not b or a;
    layer2_outputs(4316) <= b;
    layer2_outputs(4317) <= not a or b;
    layer2_outputs(4318) <= b and not a;
    layer2_outputs(4319) <= b;
    layer2_outputs(4320) <= not (a and b);
    layer2_outputs(4321) <= b and not a;
    layer2_outputs(4322) <= a;
    layer2_outputs(4323) <= a and b;
    layer2_outputs(4324) <= a xor b;
    layer2_outputs(4325) <= b;
    layer2_outputs(4326) <= not b;
    layer2_outputs(4327) <= a xor b;
    layer2_outputs(4328) <= a xor b;
    layer2_outputs(4329) <= not a or b;
    layer2_outputs(4330) <= a;
    layer2_outputs(4331) <= a and b;
    layer2_outputs(4332) <= a or b;
    layer2_outputs(4333) <= not (a xor b);
    layer2_outputs(4334) <= not a;
    layer2_outputs(4335) <= not b;
    layer2_outputs(4336) <= a xor b;
    layer2_outputs(4337) <= a xor b;
    layer2_outputs(4338) <= not b or a;
    layer2_outputs(4339) <= not b or a;
    layer2_outputs(4340) <= a;
    layer2_outputs(4341) <= b and not a;
    layer2_outputs(4342) <= not b or a;
    layer2_outputs(4343) <= a or b;
    layer2_outputs(4344) <= b and not a;
    layer2_outputs(4345) <= not (a or b);
    layer2_outputs(4346) <= not a;
    layer2_outputs(4347) <= b and not a;
    layer2_outputs(4348) <= not b;
    layer2_outputs(4349) <= a;
    layer2_outputs(4350) <= not a;
    layer2_outputs(4351) <= not b or a;
    layer2_outputs(4352) <= a xor b;
    layer2_outputs(4353) <= not b;
    layer2_outputs(4354) <= not a;
    layer2_outputs(4355) <= not (a and b);
    layer2_outputs(4356) <= not (a xor b);
    layer2_outputs(4357) <= b;
    layer2_outputs(4358) <= not (a or b);
    layer2_outputs(4359) <= not (a or b);
    layer2_outputs(4360) <= b;
    layer2_outputs(4361) <= not a;
    layer2_outputs(4362) <= a and not b;
    layer2_outputs(4363) <= not a or b;
    layer2_outputs(4364) <= not b;
    layer2_outputs(4365) <= b;
    layer2_outputs(4366) <= a xor b;
    layer2_outputs(4367) <= a;
    layer2_outputs(4368) <= b;
    layer2_outputs(4369) <= b and not a;
    layer2_outputs(4370) <= a xor b;
    layer2_outputs(4371) <= not (a xor b);
    layer2_outputs(4372) <= a and not b;
    layer2_outputs(4373) <= not b;
    layer2_outputs(4374) <= not b;
    layer2_outputs(4375) <= a and not b;
    layer2_outputs(4376) <= a and b;
    layer2_outputs(4377) <= b;
    layer2_outputs(4378) <= b and not a;
    layer2_outputs(4379) <= not a;
    layer2_outputs(4380) <= not a or b;
    layer2_outputs(4381) <= not (a xor b);
    layer2_outputs(4382) <= a;
    layer2_outputs(4383) <= a;
    layer2_outputs(4384) <= not a;
    layer2_outputs(4385) <= not a;
    layer2_outputs(4386) <= not (a and b);
    layer2_outputs(4387) <= not b or a;
    layer2_outputs(4388) <= b and not a;
    layer2_outputs(4389) <= not a;
    layer2_outputs(4390) <= not (a and b);
    layer2_outputs(4391) <= b;
    layer2_outputs(4392) <= a;
    layer2_outputs(4393) <= not (a xor b);
    layer2_outputs(4394) <= not b;
    layer2_outputs(4395) <= not (a or b);
    layer2_outputs(4396) <= a and not b;
    layer2_outputs(4397) <= b;
    layer2_outputs(4398) <= not (a and b);
    layer2_outputs(4399) <= b and not a;
    layer2_outputs(4400) <= a xor b;
    layer2_outputs(4401) <= a and not b;
    layer2_outputs(4402) <= not b;
    layer2_outputs(4403) <= a;
    layer2_outputs(4404) <= a;
    layer2_outputs(4405) <= a and b;
    layer2_outputs(4406) <= not b;
    layer2_outputs(4407) <= b;
    layer2_outputs(4408) <= b;
    layer2_outputs(4409) <= not a or b;
    layer2_outputs(4410) <= not a;
    layer2_outputs(4411) <= not b or a;
    layer2_outputs(4412) <= a xor b;
    layer2_outputs(4413) <= a and not b;
    layer2_outputs(4414) <= '1';
    layer2_outputs(4415) <= b;
    layer2_outputs(4416) <= not a;
    layer2_outputs(4417) <= not a;
    layer2_outputs(4418) <= b and not a;
    layer2_outputs(4419) <= not a or b;
    layer2_outputs(4420) <= a xor b;
    layer2_outputs(4421) <= b;
    layer2_outputs(4422) <= a and b;
    layer2_outputs(4423) <= a;
    layer2_outputs(4424) <= not (a xor b);
    layer2_outputs(4425) <= not (a and b);
    layer2_outputs(4426) <= a and not b;
    layer2_outputs(4427) <= a and not b;
    layer2_outputs(4428) <= not b or a;
    layer2_outputs(4429) <= a xor b;
    layer2_outputs(4430) <= b and not a;
    layer2_outputs(4431) <= a and b;
    layer2_outputs(4432) <= a;
    layer2_outputs(4433) <= a xor b;
    layer2_outputs(4434) <= '1';
    layer2_outputs(4435) <= not (a and b);
    layer2_outputs(4436) <= not a;
    layer2_outputs(4437) <= a or b;
    layer2_outputs(4438) <= a;
    layer2_outputs(4439) <= a and not b;
    layer2_outputs(4440) <= a;
    layer2_outputs(4441) <= b and not a;
    layer2_outputs(4442) <= a or b;
    layer2_outputs(4443) <= not b or a;
    layer2_outputs(4444) <= not a or b;
    layer2_outputs(4445) <= a xor b;
    layer2_outputs(4446) <= not a;
    layer2_outputs(4447) <= not a;
    layer2_outputs(4448) <= b;
    layer2_outputs(4449) <= not a;
    layer2_outputs(4450) <= b;
    layer2_outputs(4451) <= a;
    layer2_outputs(4452) <= b and not a;
    layer2_outputs(4453) <= not (a xor b);
    layer2_outputs(4454) <= not b or a;
    layer2_outputs(4455) <= not a or b;
    layer2_outputs(4456) <= not (a or b);
    layer2_outputs(4457) <= not b;
    layer2_outputs(4458) <= a or b;
    layer2_outputs(4459) <= a xor b;
    layer2_outputs(4460) <= b and not a;
    layer2_outputs(4461) <= not b;
    layer2_outputs(4462) <= not (a xor b);
    layer2_outputs(4463) <= not b;
    layer2_outputs(4464) <= b and not a;
    layer2_outputs(4465) <= not (a xor b);
    layer2_outputs(4466) <= not (a xor b);
    layer2_outputs(4467) <= a;
    layer2_outputs(4468) <= a;
    layer2_outputs(4469) <= not b;
    layer2_outputs(4470) <= not a or b;
    layer2_outputs(4471) <= not b or a;
    layer2_outputs(4472) <= a;
    layer2_outputs(4473) <= not (a or b);
    layer2_outputs(4474) <= a xor b;
    layer2_outputs(4475) <= not (a xor b);
    layer2_outputs(4476) <= not (a and b);
    layer2_outputs(4477) <= b;
    layer2_outputs(4478) <= b;
    layer2_outputs(4479) <= not a;
    layer2_outputs(4480) <= a;
    layer2_outputs(4481) <= not a;
    layer2_outputs(4482) <= not (a and b);
    layer2_outputs(4483) <= not a;
    layer2_outputs(4484) <= not (a and b);
    layer2_outputs(4485) <= a xor b;
    layer2_outputs(4486) <= not (a xor b);
    layer2_outputs(4487) <= not b;
    layer2_outputs(4488) <= not a;
    layer2_outputs(4489) <= not a;
    layer2_outputs(4490) <= a and b;
    layer2_outputs(4491) <= b;
    layer2_outputs(4492) <= a xor b;
    layer2_outputs(4493) <= not a;
    layer2_outputs(4494) <= not b;
    layer2_outputs(4495) <= not (a or b);
    layer2_outputs(4496) <= a or b;
    layer2_outputs(4497) <= b;
    layer2_outputs(4498) <= a;
    layer2_outputs(4499) <= a;
    layer2_outputs(4500) <= not (a xor b);
    layer2_outputs(4501) <= '1';
    layer2_outputs(4502) <= b and not a;
    layer2_outputs(4503) <= not (a xor b);
    layer2_outputs(4504) <= not (a and b);
    layer2_outputs(4505) <= not a;
    layer2_outputs(4506) <= a and not b;
    layer2_outputs(4507) <= a xor b;
    layer2_outputs(4508) <= not a;
    layer2_outputs(4509) <= not a;
    layer2_outputs(4510) <= not b;
    layer2_outputs(4511) <= not b;
    layer2_outputs(4512) <= a and not b;
    layer2_outputs(4513) <= b and not a;
    layer2_outputs(4514) <= a;
    layer2_outputs(4515) <= a xor b;
    layer2_outputs(4516) <= not b or a;
    layer2_outputs(4517) <= not b;
    layer2_outputs(4518) <= b;
    layer2_outputs(4519) <= a or b;
    layer2_outputs(4520) <= b and not a;
    layer2_outputs(4521) <= not a;
    layer2_outputs(4522) <= not b or a;
    layer2_outputs(4523) <= '0';
    layer2_outputs(4524) <= a and not b;
    layer2_outputs(4525) <= a or b;
    layer2_outputs(4526) <= b;
    layer2_outputs(4527) <= not a;
    layer2_outputs(4528) <= b;
    layer2_outputs(4529) <= a or b;
    layer2_outputs(4530) <= not (a and b);
    layer2_outputs(4531) <= not a or b;
    layer2_outputs(4532) <= a;
    layer2_outputs(4533) <= not a or b;
    layer2_outputs(4534) <= not (a xor b);
    layer2_outputs(4535) <= a and b;
    layer2_outputs(4536) <= not (a and b);
    layer2_outputs(4537) <= not b;
    layer2_outputs(4538) <= a xor b;
    layer2_outputs(4539) <= not (a xor b);
    layer2_outputs(4540) <= not b or a;
    layer2_outputs(4541) <= b;
    layer2_outputs(4542) <= a and not b;
    layer2_outputs(4543) <= not (a and b);
    layer2_outputs(4544) <= not (a xor b);
    layer2_outputs(4545) <= not (a and b);
    layer2_outputs(4546) <= a or b;
    layer2_outputs(4547) <= not b;
    layer2_outputs(4548) <= a and b;
    layer2_outputs(4549) <= b;
    layer2_outputs(4550) <= not b;
    layer2_outputs(4551) <= b and not a;
    layer2_outputs(4552) <= a;
    layer2_outputs(4553) <= a;
    layer2_outputs(4554) <= a and not b;
    layer2_outputs(4555) <= b;
    layer2_outputs(4556) <= a and b;
    layer2_outputs(4557) <= a;
    layer2_outputs(4558) <= b and not a;
    layer2_outputs(4559) <= not a or b;
    layer2_outputs(4560) <= not a;
    layer2_outputs(4561) <= a;
    layer2_outputs(4562) <= not a;
    layer2_outputs(4563) <= not (a or b);
    layer2_outputs(4564) <= not a;
    layer2_outputs(4565) <= not (a and b);
    layer2_outputs(4566) <= a;
    layer2_outputs(4567) <= not a;
    layer2_outputs(4568) <= a and b;
    layer2_outputs(4569) <= not a;
    layer2_outputs(4570) <= b;
    layer2_outputs(4571) <= not a;
    layer2_outputs(4572) <= not (a or b);
    layer2_outputs(4573) <= a;
    layer2_outputs(4574) <= '0';
    layer2_outputs(4575) <= not b;
    layer2_outputs(4576) <= not (a xor b);
    layer2_outputs(4577) <= not (a xor b);
    layer2_outputs(4578) <= not a or b;
    layer2_outputs(4579) <= a;
    layer2_outputs(4580) <= a xor b;
    layer2_outputs(4581) <= not (a xor b);
    layer2_outputs(4582) <= a or b;
    layer2_outputs(4583) <= not b;
    layer2_outputs(4584) <= not (a or b);
    layer2_outputs(4585) <= not (a xor b);
    layer2_outputs(4586) <= not a or b;
    layer2_outputs(4587) <= not b or a;
    layer2_outputs(4588) <= a and b;
    layer2_outputs(4589) <= not b or a;
    layer2_outputs(4590) <= not a;
    layer2_outputs(4591) <= a;
    layer2_outputs(4592) <= not b;
    layer2_outputs(4593) <= not a or b;
    layer2_outputs(4594) <= a;
    layer2_outputs(4595) <= not a;
    layer2_outputs(4596) <= not a;
    layer2_outputs(4597) <= b and not a;
    layer2_outputs(4598) <= b;
    layer2_outputs(4599) <= a and b;
    layer2_outputs(4600) <= not b or a;
    layer2_outputs(4601) <= a;
    layer2_outputs(4602) <= b;
    layer2_outputs(4603) <= a and b;
    layer2_outputs(4604) <= not (a and b);
    layer2_outputs(4605) <= a and not b;
    layer2_outputs(4606) <= not a;
    layer2_outputs(4607) <= not b;
    layer2_outputs(4608) <= b;
    layer2_outputs(4609) <= b;
    layer2_outputs(4610) <= b and not a;
    layer2_outputs(4611) <= a;
    layer2_outputs(4612) <= not a;
    layer2_outputs(4613) <= a;
    layer2_outputs(4614) <= a;
    layer2_outputs(4615) <= not a;
    layer2_outputs(4616) <= a and b;
    layer2_outputs(4617) <= not b or a;
    layer2_outputs(4618) <= not b or a;
    layer2_outputs(4619) <= not b;
    layer2_outputs(4620) <= not b or a;
    layer2_outputs(4621) <= not (a and b);
    layer2_outputs(4622) <= a;
    layer2_outputs(4623) <= b and not a;
    layer2_outputs(4624) <= b;
    layer2_outputs(4625) <= a;
    layer2_outputs(4626) <= a and b;
    layer2_outputs(4627) <= not b;
    layer2_outputs(4628) <= not b;
    layer2_outputs(4629) <= a xor b;
    layer2_outputs(4630) <= not a;
    layer2_outputs(4631) <= a xor b;
    layer2_outputs(4632) <= a xor b;
    layer2_outputs(4633) <= a or b;
    layer2_outputs(4634) <= a xor b;
    layer2_outputs(4635) <= not a or b;
    layer2_outputs(4636) <= a xor b;
    layer2_outputs(4637) <= a or b;
    layer2_outputs(4638) <= a or b;
    layer2_outputs(4639) <= not b;
    layer2_outputs(4640) <= a or b;
    layer2_outputs(4641) <= a or b;
    layer2_outputs(4642) <= not (a xor b);
    layer2_outputs(4643) <= not a;
    layer2_outputs(4644) <= not (a xor b);
    layer2_outputs(4645) <= a;
    layer2_outputs(4646) <= not a or b;
    layer2_outputs(4647) <= not a;
    layer2_outputs(4648) <= b and not a;
    layer2_outputs(4649) <= a and not b;
    layer2_outputs(4650) <= not (a xor b);
    layer2_outputs(4651) <= a and b;
    layer2_outputs(4652) <= a and b;
    layer2_outputs(4653) <= not a or b;
    layer2_outputs(4654) <= a xor b;
    layer2_outputs(4655) <= not a or b;
    layer2_outputs(4656) <= b and not a;
    layer2_outputs(4657) <= a or b;
    layer2_outputs(4658) <= a and not b;
    layer2_outputs(4659) <= not a;
    layer2_outputs(4660) <= a and not b;
    layer2_outputs(4661) <= a and b;
    layer2_outputs(4662) <= not a;
    layer2_outputs(4663) <= not a;
    layer2_outputs(4664) <= a and not b;
    layer2_outputs(4665) <= a and not b;
    layer2_outputs(4666) <= not (a xor b);
    layer2_outputs(4667) <= a;
    layer2_outputs(4668) <= b;
    layer2_outputs(4669) <= not a or b;
    layer2_outputs(4670) <= not b;
    layer2_outputs(4671) <= not (a xor b);
    layer2_outputs(4672) <= not a or b;
    layer2_outputs(4673) <= not a;
    layer2_outputs(4674) <= a xor b;
    layer2_outputs(4675) <= not a;
    layer2_outputs(4676) <= not (a or b);
    layer2_outputs(4677) <= not (a and b);
    layer2_outputs(4678) <= a;
    layer2_outputs(4679) <= a xor b;
    layer2_outputs(4680) <= a;
    layer2_outputs(4681) <= not (a xor b);
    layer2_outputs(4682) <= b;
    layer2_outputs(4683) <= a or b;
    layer2_outputs(4684) <= b and not a;
    layer2_outputs(4685) <= not (a and b);
    layer2_outputs(4686) <= a and not b;
    layer2_outputs(4687) <= b;
    layer2_outputs(4688) <= not (a and b);
    layer2_outputs(4689) <= a xor b;
    layer2_outputs(4690) <= b;
    layer2_outputs(4691) <= a;
    layer2_outputs(4692) <= not (a or b);
    layer2_outputs(4693) <= not (a or b);
    layer2_outputs(4694) <= a xor b;
    layer2_outputs(4695) <= a and b;
    layer2_outputs(4696) <= b;
    layer2_outputs(4697) <= a or b;
    layer2_outputs(4698) <= not a;
    layer2_outputs(4699) <= a;
    layer2_outputs(4700) <= not b or a;
    layer2_outputs(4701) <= not b;
    layer2_outputs(4702) <= not b;
    layer2_outputs(4703) <= not b or a;
    layer2_outputs(4704) <= a and not b;
    layer2_outputs(4705) <= not b or a;
    layer2_outputs(4706) <= not a;
    layer2_outputs(4707) <= not b;
    layer2_outputs(4708) <= not a;
    layer2_outputs(4709) <= not (a xor b);
    layer2_outputs(4710) <= not (a xor b);
    layer2_outputs(4711) <= not (a xor b);
    layer2_outputs(4712) <= a;
    layer2_outputs(4713) <= a;
    layer2_outputs(4714) <= not a;
    layer2_outputs(4715) <= b;
    layer2_outputs(4716) <= b;
    layer2_outputs(4717) <= a;
    layer2_outputs(4718) <= not a;
    layer2_outputs(4719) <= not (a xor b);
    layer2_outputs(4720) <= a and b;
    layer2_outputs(4721) <= a xor b;
    layer2_outputs(4722) <= not b or a;
    layer2_outputs(4723) <= not (a and b);
    layer2_outputs(4724) <= not a;
    layer2_outputs(4725) <= b;
    layer2_outputs(4726) <= not (a xor b);
    layer2_outputs(4727) <= b;
    layer2_outputs(4728) <= not (a or b);
    layer2_outputs(4729) <= not a or b;
    layer2_outputs(4730) <= a xor b;
    layer2_outputs(4731) <= not a;
    layer2_outputs(4732) <= b and not a;
    layer2_outputs(4733) <= b;
    layer2_outputs(4734) <= b;
    layer2_outputs(4735) <= a xor b;
    layer2_outputs(4736) <= a xor b;
    layer2_outputs(4737) <= b;
    layer2_outputs(4738) <= '1';
    layer2_outputs(4739) <= not (a xor b);
    layer2_outputs(4740) <= not a;
    layer2_outputs(4741) <= a xor b;
    layer2_outputs(4742) <= not b or a;
    layer2_outputs(4743) <= not a;
    layer2_outputs(4744) <= not b;
    layer2_outputs(4745) <= b;
    layer2_outputs(4746) <= a or b;
    layer2_outputs(4747) <= not (a xor b);
    layer2_outputs(4748) <= not b;
    layer2_outputs(4749) <= a;
    layer2_outputs(4750) <= not b;
    layer2_outputs(4751) <= not (a or b);
    layer2_outputs(4752) <= not a;
    layer2_outputs(4753) <= not a;
    layer2_outputs(4754) <= a or b;
    layer2_outputs(4755) <= a and b;
    layer2_outputs(4756) <= a xor b;
    layer2_outputs(4757) <= a;
    layer2_outputs(4758) <= b;
    layer2_outputs(4759) <= not b;
    layer2_outputs(4760) <= a and b;
    layer2_outputs(4761) <= not a;
    layer2_outputs(4762) <= not a;
    layer2_outputs(4763) <= not (a xor b);
    layer2_outputs(4764) <= b;
    layer2_outputs(4765) <= a;
    layer2_outputs(4766) <= a;
    layer2_outputs(4767) <= not (a xor b);
    layer2_outputs(4768) <= b;
    layer2_outputs(4769) <= b;
    layer2_outputs(4770) <= a;
    layer2_outputs(4771) <= not (a and b);
    layer2_outputs(4772) <= not b;
    layer2_outputs(4773) <= a;
    layer2_outputs(4774) <= not (a or b);
    layer2_outputs(4775) <= a xor b;
    layer2_outputs(4776) <= not b;
    layer2_outputs(4777) <= a and not b;
    layer2_outputs(4778) <= not (a xor b);
    layer2_outputs(4779) <= a xor b;
    layer2_outputs(4780) <= a;
    layer2_outputs(4781) <= b and not a;
    layer2_outputs(4782) <= a and not b;
    layer2_outputs(4783) <= not b or a;
    layer2_outputs(4784) <= b;
    layer2_outputs(4785) <= b and not a;
    layer2_outputs(4786) <= not a or b;
    layer2_outputs(4787) <= not a;
    layer2_outputs(4788) <= not a or b;
    layer2_outputs(4789) <= a xor b;
    layer2_outputs(4790) <= not (a xor b);
    layer2_outputs(4791) <= not (a or b);
    layer2_outputs(4792) <= a or b;
    layer2_outputs(4793) <= not b;
    layer2_outputs(4794) <= not b or a;
    layer2_outputs(4795) <= not b or a;
    layer2_outputs(4796) <= b and not a;
    layer2_outputs(4797) <= not (a or b);
    layer2_outputs(4798) <= a and b;
    layer2_outputs(4799) <= a xor b;
    layer2_outputs(4800) <= a and b;
    layer2_outputs(4801) <= not a or b;
    layer2_outputs(4802) <= a or b;
    layer2_outputs(4803) <= not b;
    layer2_outputs(4804) <= b and not a;
    layer2_outputs(4805) <= not a;
    layer2_outputs(4806) <= a xor b;
    layer2_outputs(4807) <= not b;
    layer2_outputs(4808) <= not a;
    layer2_outputs(4809) <= a;
    layer2_outputs(4810) <= a or b;
    layer2_outputs(4811) <= b;
    layer2_outputs(4812) <= a;
    layer2_outputs(4813) <= b;
    layer2_outputs(4814) <= a;
    layer2_outputs(4815) <= a;
    layer2_outputs(4816) <= a and b;
    layer2_outputs(4817) <= a xor b;
    layer2_outputs(4818) <= a or b;
    layer2_outputs(4819) <= not b;
    layer2_outputs(4820) <= b;
    layer2_outputs(4821) <= not b;
    layer2_outputs(4822) <= not a;
    layer2_outputs(4823) <= not b;
    layer2_outputs(4824) <= a;
    layer2_outputs(4825) <= not a;
    layer2_outputs(4826) <= a xor b;
    layer2_outputs(4827) <= b;
    layer2_outputs(4828) <= not a;
    layer2_outputs(4829) <= b;
    layer2_outputs(4830) <= not (a or b);
    layer2_outputs(4831) <= a xor b;
    layer2_outputs(4832) <= a;
    layer2_outputs(4833) <= a and b;
    layer2_outputs(4834) <= not a or b;
    layer2_outputs(4835) <= a and not b;
    layer2_outputs(4836) <= not (a xor b);
    layer2_outputs(4837) <= a and not b;
    layer2_outputs(4838) <= not b or a;
    layer2_outputs(4839) <= not b or a;
    layer2_outputs(4840) <= not b;
    layer2_outputs(4841) <= a xor b;
    layer2_outputs(4842) <= not b or a;
    layer2_outputs(4843) <= a;
    layer2_outputs(4844) <= not a or b;
    layer2_outputs(4845) <= b and not a;
    layer2_outputs(4846) <= not b or a;
    layer2_outputs(4847) <= not (a or b);
    layer2_outputs(4848) <= b and not a;
    layer2_outputs(4849) <= not b or a;
    layer2_outputs(4850) <= not (a xor b);
    layer2_outputs(4851) <= not (a or b);
    layer2_outputs(4852) <= not a or b;
    layer2_outputs(4853) <= b;
    layer2_outputs(4854) <= a xor b;
    layer2_outputs(4855) <= not a;
    layer2_outputs(4856) <= not a or b;
    layer2_outputs(4857) <= b;
    layer2_outputs(4858) <= not (a xor b);
    layer2_outputs(4859) <= not (a xor b);
    layer2_outputs(4860) <= a and b;
    layer2_outputs(4861) <= not b;
    layer2_outputs(4862) <= not (a and b);
    layer2_outputs(4863) <= not a;
    layer2_outputs(4864) <= a or b;
    layer2_outputs(4865) <= not a;
    layer2_outputs(4866) <= b and not a;
    layer2_outputs(4867) <= not b or a;
    layer2_outputs(4868) <= a or b;
    layer2_outputs(4869) <= a;
    layer2_outputs(4870) <= a or b;
    layer2_outputs(4871) <= a and b;
    layer2_outputs(4872) <= not (a and b);
    layer2_outputs(4873) <= a and not b;
    layer2_outputs(4874) <= a;
    layer2_outputs(4875) <= b and not a;
    layer2_outputs(4876) <= not (a xor b);
    layer2_outputs(4877) <= not (a and b);
    layer2_outputs(4878) <= b;
    layer2_outputs(4879) <= a;
    layer2_outputs(4880) <= b and not a;
    layer2_outputs(4881) <= not b or a;
    layer2_outputs(4882) <= b and not a;
    layer2_outputs(4883) <= b;
    layer2_outputs(4884) <= not a;
    layer2_outputs(4885) <= not (a and b);
    layer2_outputs(4886) <= not b;
    layer2_outputs(4887) <= b and not a;
    layer2_outputs(4888) <= not a;
    layer2_outputs(4889) <= not (a xor b);
    layer2_outputs(4890) <= b;
    layer2_outputs(4891) <= not a;
    layer2_outputs(4892) <= a and b;
    layer2_outputs(4893) <= not b;
    layer2_outputs(4894) <= not (a xor b);
    layer2_outputs(4895) <= '1';
    layer2_outputs(4896) <= a;
    layer2_outputs(4897) <= not (a or b);
    layer2_outputs(4898) <= not (a xor b);
    layer2_outputs(4899) <= not a or b;
    layer2_outputs(4900) <= not (a and b);
    layer2_outputs(4901) <= b;
    layer2_outputs(4902) <= a and not b;
    layer2_outputs(4903) <= not (a or b);
    layer2_outputs(4904) <= a;
    layer2_outputs(4905) <= not (a xor b);
    layer2_outputs(4906) <= not a;
    layer2_outputs(4907) <= not a;
    layer2_outputs(4908) <= not (a and b);
    layer2_outputs(4909) <= a xor b;
    layer2_outputs(4910) <= not (a and b);
    layer2_outputs(4911) <= b;
    layer2_outputs(4912) <= a or b;
    layer2_outputs(4913) <= not b;
    layer2_outputs(4914) <= not (a or b);
    layer2_outputs(4915) <= not (a and b);
    layer2_outputs(4916) <= b and not a;
    layer2_outputs(4917) <= a;
    layer2_outputs(4918) <= b;
    layer2_outputs(4919) <= b;
    layer2_outputs(4920) <= a and b;
    layer2_outputs(4921) <= not (a and b);
    layer2_outputs(4922) <= not b;
    layer2_outputs(4923) <= not a;
    layer2_outputs(4924) <= b;
    layer2_outputs(4925) <= '1';
    layer2_outputs(4926) <= not (a xor b);
    layer2_outputs(4927) <= a or b;
    layer2_outputs(4928) <= a;
    layer2_outputs(4929) <= not (a and b);
    layer2_outputs(4930) <= not (a xor b);
    layer2_outputs(4931) <= b;
    layer2_outputs(4932) <= not a;
    layer2_outputs(4933) <= not (a and b);
    layer2_outputs(4934) <= a and not b;
    layer2_outputs(4935) <= a;
    layer2_outputs(4936) <= not a;
    layer2_outputs(4937) <= b and not a;
    layer2_outputs(4938) <= not a or b;
    layer2_outputs(4939) <= a;
    layer2_outputs(4940) <= a and b;
    layer2_outputs(4941) <= b;
    layer2_outputs(4942) <= not a;
    layer2_outputs(4943) <= a and not b;
    layer2_outputs(4944) <= a xor b;
    layer2_outputs(4945) <= not a or b;
    layer2_outputs(4946) <= not (a xor b);
    layer2_outputs(4947) <= b;
    layer2_outputs(4948) <= a and b;
    layer2_outputs(4949) <= a xor b;
    layer2_outputs(4950) <= a and b;
    layer2_outputs(4951) <= a and not b;
    layer2_outputs(4952) <= a;
    layer2_outputs(4953) <= b;
    layer2_outputs(4954) <= not a;
    layer2_outputs(4955) <= not b;
    layer2_outputs(4956) <= not b or a;
    layer2_outputs(4957) <= not b;
    layer2_outputs(4958) <= '0';
    layer2_outputs(4959) <= a or b;
    layer2_outputs(4960) <= not (a xor b);
    layer2_outputs(4961) <= a xor b;
    layer2_outputs(4962) <= not b;
    layer2_outputs(4963) <= b and not a;
    layer2_outputs(4964) <= b and not a;
    layer2_outputs(4965) <= b;
    layer2_outputs(4966) <= not a;
    layer2_outputs(4967) <= a and b;
    layer2_outputs(4968) <= a and not b;
    layer2_outputs(4969) <= not (a and b);
    layer2_outputs(4970) <= a or b;
    layer2_outputs(4971) <= a and b;
    layer2_outputs(4972) <= not b;
    layer2_outputs(4973) <= b;
    layer2_outputs(4974) <= not (a xor b);
    layer2_outputs(4975) <= not a;
    layer2_outputs(4976) <= a or b;
    layer2_outputs(4977) <= not b;
    layer2_outputs(4978) <= a;
    layer2_outputs(4979) <= '0';
    layer2_outputs(4980) <= not b;
    layer2_outputs(4981) <= a;
    layer2_outputs(4982) <= not (a xor b);
    layer2_outputs(4983) <= not a;
    layer2_outputs(4984) <= a xor b;
    layer2_outputs(4985) <= not (a or b);
    layer2_outputs(4986) <= not a;
    layer2_outputs(4987) <= a;
    layer2_outputs(4988) <= not (a xor b);
    layer2_outputs(4989) <= not (a or b);
    layer2_outputs(4990) <= not b;
    layer2_outputs(4991) <= not a;
    layer2_outputs(4992) <= not (a xor b);
    layer2_outputs(4993) <= a;
    layer2_outputs(4994) <= a;
    layer2_outputs(4995) <= not b;
    layer2_outputs(4996) <= not b;
    layer2_outputs(4997) <= b and not a;
    layer2_outputs(4998) <= a xor b;
    layer2_outputs(4999) <= b;
    layer2_outputs(5000) <= not b;
    layer2_outputs(5001) <= not a;
    layer2_outputs(5002) <= a;
    layer2_outputs(5003) <= a;
    layer2_outputs(5004) <= '0';
    layer2_outputs(5005) <= a;
    layer2_outputs(5006) <= a xor b;
    layer2_outputs(5007) <= not (a xor b);
    layer2_outputs(5008) <= a;
    layer2_outputs(5009) <= not (a and b);
    layer2_outputs(5010) <= not (a or b);
    layer2_outputs(5011) <= not (a xor b);
    layer2_outputs(5012) <= not (a xor b);
    layer2_outputs(5013) <= b;
    layer2_outputs(5014) <= not (a xor b);
    layer2_outputs(5015) <= a and not b;
    layer2_outputs(5016) <= not (a xor b);
    layer2_outputs(5017) <= b;
    layer2_outputs(5018) <= not b;
    layer2_outputs(5019) <= a xor b;
    layer2_outputs(5020) <= a;
    layer2_outputs(5021) <= b;
    layer2_outputs(5022) <= not b;
    layer2_outputs(5023) <= a and b;
    layer2_outputs(5024) <= a and b;
    layer2_outputs(5025) <= a and b;
    layer2_outputs(5026) <= not b;
    layer2_outputs(5027) <= not a;
    layer2_outputs(5028) <= not (a and b);
    layer2_outputs(5029) <= a xor b;
    layer2_outputs(5030) <= not a or b;
    layer2_outputs(5031) <= not a;
    layer2_outputs(5032) <= a;
    layer2_outputs(5033) <= not a or b;
    layer2_outputs(5034) <= not a;
    layer2_outputs(5035) <= a xor b;
    layer2_outputs(5036) <= not (a xor b);
    layer2_outputs(5037) <= a and not b;
    layer2_outputs(5038) <= not b;
    layer2_outputs(5039) <= '0';
    layer2_outputs(5040) <= a and not b;
    layer2_outputs(5041) <= not (a xor b);
    layer2_outputs(5042) <= a;
    layer2_outputs(5043) <= not (a xor b);
    layer2_outputs(5044) <= b and not a;
    layer2_outputs(5045) <= b;
    layer2_outputs(5046) <= '1';
    layer2_outputs(5047) <= not (a xor b);
    layer2_outputs(5048) <= a or b;
    layer2_outputs(5049) <= not a;
    layer2_outputs(5050) <= '1';
    layer2_outputs(5051) <= not (a xor b);
    layer2_outputs(5052) <= a xor b;
    layer2_outputs(5053) <= a;
    layer2_outputs(5054) <= not (a and b);
    layer2_outputs(5055) <= a;
    layer2_outputs(5056) <= not b;
    layer2_outputs(5057) <= b and not a;
    layer2_outputs(5058) <= not (a xor b);
    layer2_outputs(5059) <= b;
    layer2_outputs(5060) <= not (a or b);
    layer2_outputs(5061) <= not b;
    layer2_outputs(5062) <= not (a xor b);
    layer2_outputs(5063) <= a and b;
    layer2_outputs(5064) <= a xor b;
    layer2_outputs(5065) <= not (a or b);
    layer2_outputs(5066) <= b and not a;
    layer2_outputs(5067) <= not (a or b);
    layer2_outputs(5068) <= not b or a;
    layer2_outputs(5069) <= not (a xor b);
    layer2_outputs(5070) <= not (a xor b);
    layer2_outputs(5071) <= not b or a;
    layer2_outputs(5072) <= not b;
    layer2_outputs(5073) <= not b or a;
    layer2_outputs(5074) <= not b;
    layer2_outputs(5075) <= b;
    layer2_outputs(5076) <= a xor b;
    layer2_outputs(5077) <= a;
    layer2_outputs(5078) <= a;
    layer2_outputs(5079) <= a;
    layer2_outputs(5080) <= b;
    layer2_outputs(5081) <= a and b;
    layer2_outputs(5082) <= a and not b;
    layer2_outputs(5083) <= a or b;
    layer2_outputs(5084) <= not (a or b);
    layer2_outputs(5085) <= a;
    layer2_outputs(5086) <= not (a or b);
    layer2_outputs(5087) <= not a;
    layer2_outputs(5088) <= not (a or b);
    layer2_outputs(5089) <= a xor b;
    layer2_outputs(5090) <= a xor b;
    layer2_outputs(5091) <= not b;
    layer2_outputs(5092) <= a and b;
    layer2_outputs(5093) <= a xor b;
    layer2_outputs(5094) <= a and b;
    layer2_outputs(5095) <= not (a or b);
    layer2_outputs(5096) <= not b;
    layer2_outputs(5097) <= not a;
    layer2_outputs(5098) <= not (a xor b);
    layer2_outputs(5099) <= a;
    layer2_outputs(5100) <= not b;
    layer2_outputs(5101) <= a and not b;
    layer2_outputs(5102) <= not (a xor b);
    layer2_outputs(5103) <= not b or a;
    layer2_outputs(5104) <= not b;
    layer2_outputs(5105) <= a;
    layer2_outputs(5106) <= a xor b;
    layer2_outputs(5107) <= not (a and b);
    layer2_outputs(5108) <= not b;
    layer2_outputs(5109) <= b;
    layer2_outputs(5110) <= a and not b;
    layer2_outputs(5111) <= not (a xor b);
    layer2_outputs(5112) <= a xor b;
    layer2_outputs(5113) <= not a or b;
    layer2_outputs(5114) <= a xor b;
    layer2_outputs(5115) <= a;
    layer2_outputs(5116) <= a;
    layer2_outputs(5117) <= a or b;
    layer2_outputs(5118) <= not a;
    layer2_outputs(5119) <= a and not b;
    layer2_outputs(5120) <= a;
    layer2_outputs(5121) <= a;
    layer2_outputs(5122) <= b;
    layer2_outputs(5123) <= b and not a;
    layer2_outputs(5124) <= a xor b;
    layer2_outputs(5125) <= a and not b;
    layer2_outputs(5126) <= a;
    layer2_outputs(5127) <= a and not b;
    layer2_outputs(5128) <= not (a or b);
    layer2_outputs(5129) <= not b or a;
    layer2_outputs(5130) <= not (a or b);
    layer2_outputs(5131) <= a and b;
    layer2_outputs(5132) <= a xor b;
    layer2_outputs(5133) <= b;
    layer2_outputs(5134) <= not b or a;
    layer2_outputs(5135) <= b;
    layer2_outputs(5136) <= a xor b;
    layer2_outputs(5137) <= not (a and b);
    layer2_outputs(5138) <= b;
    layer2_outputs(5139) <= not b;
    layer2_outputs(5140) <= b;
    layer2_outputs(5141) <= b;
    layer2_outputs(5142) <= a xor b;
    layer2_outputs(5143) <= a;
    layer2_outputs(5144) <= a and not b;
    layer2_outputs(5145) <= not b or a;
    layer2_outputs(5146) <= not (a xor b);
    layer2_outputs(5147) <= not (a or b);
    layer2_outputs(5148) <= not (a xor b);
    layer2_outputs(5149) <= a;
    layer2_outputs(5150) <= not b;
    layer2_outputs(5151) <= b and not a;
    layer2_outputs(5152) <= not b;
    layer2_outputs(5153) <= not (a xor b);
    layer2_outputs(5154) <= not a;
    layer2_outputs(5155) <= not b;
    layer2_outputs(5156) <= not a;
    layer2_outputs(5157) <= a and b;
    layer2_outputs(5158) <= not a;
    layer2_outputs(5159) <= a xor b;
    layer2_outputs(5160) <= not b or a;
    layer2_outputs(5161) <= not a or b;
    layer2_outputs(5162) <= not a;
    layer2_outputs(5163) <= not a;
    layer2_outputs(5164) <= b;
    layer2_outputs(5165) <= a;
    layer2_outputs(5166) <= b;
    layer2_outputs(5167) <= a xor b;
    layer2_outputs(5168) <= b and not a;
    layer2_outputs(5169) <= a xor b;
    layer2_outputs(5170) <= not (a xor b);
    layer2_outputs(5171) <= not (a or b);
    layer2_outputs(5172) <= not a;
    layer2_outputs(5173) <= not b;
    layer2_outputs(5174) <= not b or a;
    layer2_outputs(5175) <= a xor b;
    layer2_outputs(5176) <= b and not a;
    layer2_outputs(5177) <= not b;
    layer2_outputs(5178) <= a and b;
    layer2_outputs(5179) <= not b;
    layer2_outputs(5180) <= not (a and b);
    layer2_outputs(5181) <= not b;
    layer2_outputs(5182) <= a xor b;
    layer2_outputs(5183) <= b;
    layer2_outputs(5184) <= not (a xor b);
    layer2_outputs(5185) <= b and not a;
    layer2_outputs(5186) <= b and not a;
    layer2_outputs(5187) <= not a;
    layer2_outputs(5188) <= not a;
    layer2_outputs(5189) <= not (a xor b);
    layer2_outputs(5190) <= b;
    layer2_outputs(5191) <= b;
    layer2_outputs(5192) <= b;
    layer2_outputs(5193) <= '0';
    layer2_outputs(5194) <= a xor b;
    layer2_outputs(5195) <= not a;
    layer2_outputs(5196) <= a and not b;
    layer2_outputs(5197) <= not a;
    layer2_outputs(5198) <= not (a xor b);
    layer2_outputs(5199) <= not (a and b);
    layer2_outputs(5200) <= a and not b;
    layer2_outputs(5201) <= not (a xor b);
    layer2_outputs(5202) <= not a or b;
    layer2_outputs(5203) <= a or b;
    layer2_outputs(5204) <= not b;
    layer2_outputs(5205) <= a;
    layer2_outputs(5206) <= not a or b;
    layer2_outputs(5207) <= not b or a;
    layer2_outputs(5208) <= not b;
    layer2_outputs(5209) <= a xor b;
    layer2_outputs(5210) <= b;
    layer2_outputs(5211) <= not a or b;
    layer2_outputs(5212) <= not a or b;
    layer2_outputs(5213) <= not (a or b);
    layer2_outputs(5214) <= not (a xor b);
    layer2_outputs(5215) <= b and not a;
    layer2_outputs(5216) <= not a;
    layer2_outputs(5217) <= not b;
    layer2_outputs(5218) <= not (a and b);
    layer2_outputs(5219) <= b;
    layer2_outputs(5220) <= not b;
    layer2_outputs(5221) <= not (a and b);
    layer2_outputs(5222) <= not (a or b);
    layer2_outputs(5223) <= not (a and b);
    layer2_outputs(5224) <= not (a xor b);
    layer2_outputs(5225) <= not a;
    layer2_outputs(5226) <= not (a or b);
    layer2_outputs(5227) <= not (a or b);
    layer2_outputs(5228) <= not b;
    layer2_outputs(5229) <= b and not a;
    layer2_outputs(5230) <= not b;
    layer2_outputs(5231) <= a and b;
    layer2_outputs(5232) <= b and not a;
    layer2_outputs(5233) <= not (a or b);
    layer2_outputs(5234) <= not (a and b);
    layer2_outputs(5235) <= not (a xor b);
    layer2_outputs(5236) <= not b;
    layer2_outputs(5237) <= not (a or b);
    layer2_outputs(5238) <= not (a and b);
    layer2_outputs(5239) <= not (a or b);
    layer2_outputs(5240) <= b;
    layer2_outputs(5241) <= not b;
    layer2_outputs(5242) <= a;
    layer2_outputs(5243) <= a or b;
    layer2_outputs(5244) <= not a;
    layer2_outputs(5245) <= b;
    layer2_outputs(5246) <= not b or a;
    layer2_outputs(5247) <= not a or b;
    layer2_outputs(5248) <= not b or a;
    layer2_outputs(5249) <= not b or a;
    layer2_outputs(5250) <= a;
    layer2_outputs(5251) <= not a;
    layer2_outputs(5252) <= not b or a;
    layer2_outputs(5253) <= a and b;
    layer2_outputs(5254) <= not b;
    layer2_outputs(5255) <= b;
    layer2_outputs(5256) <= not (a and b);
    layer2_outputs(5257) <= not a;
    layer2_outputs(5258) <= b;
    layer2_outputs(5259) <= a;
    layer2_outputs(5260) <= not a;
    layer2_outputs(5261) <= a or b;
    layer2_outputs(5262) <= not (a or b);
    layer2_outputs(5263) <= a;
    layer2_outputs(5264) <= a xor b;
    layer2_outputs(5265) <= not b;
    layer2_outputs(5266) <= not (a and b);
    layer2_outputs(5267) <= not a;
    layer2_outputs(5268) <= not (a xor b);
    layer2_outputs(5269) <= a and b;
    layer2_outputs(5270) <= not b;
    layer2_outputs(5271) <= not b or a;
    layer2_outputs(5272) <= b;
    layer2_outputs(5273) <= not (a xor b);
    layer2_outputs(5274) <= not (a or b);
    layer2_outputs(5275) <= b;
    layer2_outputs(5276) <= b and not a;
    layer2_outputs(5277) <= not b or a;
    layer2_outputs(5278) <= not (a xor b);
    layer2_outputs(5279) <= a xor b;
    layer2_outputs(5280) <= a xor b;
    layer2_outputs(5281) <= not b;
    layer2_outputs(5282) <= not b;
    layer2_outputs(5283) <= not b or a;
    layer2_outputs(5284) <= a;
    layer2_outputs(5285) <= not a or b;
    layer2_outputs(5286) <= not (a and b);
    layer2_outputs(5287) <= not b;
    layer2_outputs(5288) <= not (a xor b);
    layer2_outputs(5289) <= not b;
    layer2_outputs(5290) <= b;
    layer2_outputs(5291) <= not a;
    layer2_outputs(5292) <= not (a and b);
    layer2_outputs(5293) <= a or b;
    layer2_outputs(5294) <= not a or b;
    layer2_outputs(5295) <= b;
    layer2_outputs(5296) <= b and not a;
    layer2_outputs(5297) <= a and b;
    layer2_outputs(5298) <= not b;
    layer2_outputs(5299) <= a;
    layer2_outputs(5300) <= not (a xor b);
    layer2_outputs(5301) <= not b or a;
    layer2_outputs(5302) <= a;
    layer2_outputs(5303) <= not (a xor b);
    layer2_outputs(5304) <= a;
    layer2_outputs(5305) <= not a or b;
    layer2_outputs(5306) <= not a or b;
    layer2_outputs(5307) <= not b;
    layer2_outputs(5308) <= not b or a;
    layer2_outputs(5309) <= not b or a;
    layer2_outputs(5310) <= a and not b;
    layer2_outputs(5311) <= not b;
    layer2_outputs(5312) <= not b;
    layer2_outputs(5313) <= b;
    layer2_outputs(5314) <= not (a xor b);
    layer2_outputs(5315) <= not (a xor b);
    layer2_outputs(5316) <= a or b;
    layer2_outputs(5317) <= not a;
    layer2_outputs(5318) <= not b or a;
    layer2_outputs(5319) <= not b;
    layer2_outputs(5320) <= a;
    layer2_outputs(5321) <= not b;
    layer2_outputs(5322) <= not b or a;
    layer2_outputs(5323) <= a and b;
    layer2_outputs(5324) <= not (a xor b);
    layer2_outputs(5325) <= not a;
    layer2_outputs(5326) <= a xor b;
    layer2_outputs(5327) <= a or b;
    layer2_outputs(5328) <= not (a xor b);
    layer2_outputs(5329) <= not (a xor b);
    layer2_outputs(5330) <= not a;
    layer2_outputs(5331) <= not b;
    layer2_outputs(5332) <= a;
    layer2_outputs(5333) <= a or b;
    layer2_outputs(5334) <= not (a xor b);
    layer2_outputs(5335) <= not b;
    layer2_outputs(5336) <= '1';
    layer2_outputs(5337) <= a and not b;
    layer2_outputs(5338) <= a and not b;
    layer2_outputs(5339) <= not (a and b);
    layer2_outputs(5340) <= a;
    layer2_outputs(5341) <= a xor b;
    layer2_outputs(5342) <= b;
    layer2_outputs(5343) <= not b or a;
    layer2_outputs(5344) <= b;
    layer2_outputs(5345) <= a;
    layer2_outputs(5346) <= b and not a;
    layer2_outputs(5347) <= a or b;
    layer2_outputs(5348) <= a xor b;
    layer2_outputs(5349) <= a;
    layer2_outputs(5350) <= not (a or b);
    layer2_outputs(5351) <= not b;
    layer2_outputs(5352) <= a;
    layer2_outputs(5353) <= not a or b;
    layer2_outputs(5354) <= not a;
    layer2_outputs(5355) <= not (a or b);
    layer2_outputs(5356) <= b;
    layer2_outputs(5357) <= a or b;
    layer2_outputs(5358) <= a or b;
    layer2_outputs(5359) <= a;
    layer2_outputs(5360) <= a or b;
    layer2_outputs(5361) <= not (a and b);
    layer2_outputs(5362) <= not a or b;
    layer2_outputs(5363) <= not (a or b);
    layer2_outputs(5364) <= b and not a;
    layer2_outputs(5365) <= not a or b;
    layer2_outputs(5366) <= a and b;
    layer2_outputs(5367) <= b and not a;
    layer2_outputs(5368) <= not a;
    layer2_outputs(5369) <= not (a or b);
    layer2_outputs(5370) <= a;
    layer2_outputs(5371) <= not b or a;
    layer2_outputs(5372) <= not (a xor b);
    layer2_outputs(5373) <= a or b;
    layer2_outputs(5374) <= a and b;
    layer2_outputs(5375) <= not a;
    layer2_outputs(5376) <= not (a or b);
    layer2_outputs(5377) <= a or b;
    layer2_outputs(5378) <= a and not b;
    layer2_outputs(5379) <= b;
    layer2_outputs(5380) <= not (a xor b);
    layer2_outputs(5381) <= a or b;
    layer2_outputs(5382) <= a;
    layer2_outputs(5383) <= not b or a;
    layer2_outputs(5384) <= not a;
    layer2_outputs(5385) <= a or b;
    layer2_outputs(5386) <= a and not b;
    layer2_outputs(5387) <= a and not b;
    layer2_outputs(5388) <= not a;
    layer2_outputs(5389) <= a or b;
    layer2_outputs(5390) <= not (a or b);
    layer2_outputs(5391) <= a and b;
    layer2_outputs(5392) <= not a;
    layer2_outputs(5393) <= not b or a;
    layer2_outputs(5394) <= a;
    layer2_outputs(5395) <= not b;
    layer2_outputs(5396) <= a and b;
    layer2_outputs(5397) <= not (a or b);
    layer2_outputs(5398) <= b and not a;
    layer2_outputs(5399) <= not (a xor b);
    layer2_outputs(5400) <= a;
    layer2_outputs(5401) <= not (a xor b);
    layer2_outputs(5402) <= not a or b;
    layer2_outputs(5403) <= a or b;
    layer2_outputs(5404) <= b and not a;
    layer2_outputs(5405) <= not b or a;
    layer2_outputs(5406) <= not (a or b);
    layer2_outputs(5407) <= a and b;
    layer2_outputs(5408) <= b;
    layer2_outputs(5409) <= not b or a;
    layer2_outputs(5410) <= a and b;
    layer2_outputs(5411) <= a xor b;
    layer2_outputs(5412) <= not b;
    layer2_outputs(5413) <= a;
    layer2_outputs(5414) <= a and not b;
    layer2_outputs(5415) <= not (a xor b);
    layer2_outputs(5416) <= a or b;
    layer2_outputs(5417) <= a;
    layer2_outputs(5418) <= a and b;
    layer2_outputs(5419) <= a;
    layer2_outputs(5420) <= not (a xor b);
    layer2_outputs(5421) <= not (a and b);
    layer2_outputs(5422) <= not b;
    layer2_outputs(5423) <= not a or b;
    layer2_outputs(5424) <= not b or a;
    layer2_outputs(5425) <= a or b;
    layer2_outputs(5426) <= not (a xor b);
    layer2_outputs(5427) <= a;
    layer2_outputs(5428) <= b;
    layer2_outputs(5429) <= not (a xor b);
    layer2_outputs(5430) <= b;
    layer2_outputs(5431) <= not (a and b);
    layer2_outputs(5432) <= b;
    layer2_outputs(5433) <= not b;
    layer2_outputs(5434) <= not (a or b);
    layer2_outputs(5435) <= b and not a;
    layer2_outputs(5436) <= a xor b;
    layer2_outputs(5437) <= a and b;
    layer2_outputs(5438) <= a xor b;
    layer2_outputs(5439) <= a xor b;
    layer2_outputs(5440) <= not (a and b);
    layer2_outputs(5441) <= not b;
    layer2_outputs(5442) <= not (a or b);
    layer2_outputs(5443) <= a and not b;
    layer2_outputs(5444) <= not b;
    layer2_outputs(5445) <= a xor b;
    layer2_outputs(5446) <= a;
    layer2_outputs(5447) <= a xor b;
    layer2_outputs(5448) <= not b;
    layer2_outputs(5449) <= a;
    layer2_outputs(5450) <= b;
    layer2_outputs(5451) <= not (a or b);
    layer2_outputs(5452) <= a and b;
    layer2_outputs(5453) <= b and not a;
    layer2_outputs(5454) <= not (a or b);
    layer2_outputs(5455) <= b and not a;
    layer2_outputs(5456) <= b;
    layer2_outputs(5457) <= not a;
    layer2_outputs(5458) <= not (a or b);
    layer2_outputs(5459) <= not b;
    layer2_outputs(5460) <= a;
    layer2_outputs(5461) <= a or b;
    layer2_outputs(5462) <= not a;
    layer2_outputs(5463) <= a;
    layer2_outputs(5464) <= not (a xor b);
    layer2_outputs(5465) <= b;
    layer2_outputs(5466) <= b and not a;
    layer2_outputs(5467) <= a and b;
    layer2_outputs(5468) <= a xor b;
    layer2_outputs(5469) <= not a;
    layer2_outputs(5470) <= not a;
    layer2_outputs(5471) <= a or b;
    layer2_outputs(5472) <= not (a or b);
    layer2_outputs(5473) <= not a;
    layer2_outputs(5474) <= not (a or b);
    layer2_outputs(5475) <= not (a and b);
    layer2_outputs(5476) <= a xor b;
    layer2_outputs(5477) <= not (a xor b);
    layer2_outputs(5478) <= a;
    layer2_outputs(5479) <= not a;
    layer2_outputs(5480) <= not b or a;
    layer2_outputs(5481) <= b and not a;
    layer2_outputs(5482) <= not a;
    layer2_outputs(5483) <= a and b;
    layer2_outputs(5484) <= b;
    layer2_outputs(5485) <= not (a xor b);
    layer2_outputs(5486) <= b and not a;
    layer2_outputs(5487) <= not a or b;
    layer2_outputs(5488) <= not (a and b);
    layer2_outputs(5489) <= not (a xor b);
    layer2_outputs(5490) <= a and not b;
    layer2_outputs(5491) <= not b;
    layer2_outputs(5492) <= a;
    layer2_outputs(5493) <= b and not a;
    layer2_outputs(5494) <= not a;
    layer2_outputs(5495) <= a and not b;
    layer2_outputs(5496) <= not (a and b);
    layer2_outputs(5497) <= not (a xor b);
    layer2_outputs(5498) <= not b or a;
    layer2_outputs(5499) <= not b;
    layer2_outputs(5500) <= a xor b;
    layer2_outputs(5501) <= b and not a;
    layer2_outputs(5502) <= not (a xor b);
    layer2_outputs(5503) <= not (a xor b);
    layer2_outputs(5504) <= a;
    layer2_outputs(5505) <= a;
    layer2_outputs(5506) <= not a;
    layer2_outputs(5507) <= not (a or b);
    layer2_outputs(5508) <= not (a or b);
    layer2_outputs(5509) <= not a;
    layer2_outputs(5510) <= a and b;
    layer2_outputs(5511) <= b;
    layer2_outputs(5512) <= not (a or b);
    layer2_outputs(5513) <= not a;
    layer2_outputs(5514) <= not (a or b);
    layer2_outputs(5515) <= a;
    layer2_outputs(5516) <= not b;
    layer2_outputs(5517) <= a or b;
    layer2_outputs(5518) <= not (a xor b);
    layer2_outputs(5519) <= a;
    layer2_outputs(5520) <= b;
    layer2_outputs(5521) <= a xor b;
    layer2_outputs(5522) <= a;
    layer2_outputs(5523) <= not (a or b);
    layer2_outputs(5524) <= a and not b;
    layer2_outputs(5525) <= b and not a;
    layer2_outputs(5526) <= not a;
    layer2_outputs(5527) <= a;
    layer2_outputs(5528) <= not a;
    layer2_outputs(5529) <= not (a or b);
    layer2_outputs(5530) <= not a or b;
    layer2_outputs(5531) <= a and b;
    layer2_outputs(5532) <= b;
    layer2_outputs(5533) <= a;
    layer2_outputs(5534) <= a and not b;
    layer2_outputs(5535) <= b and not a;
    layer2_outputs(5536) <= not b;
    layer2_outputs(5537) <= b and not a;
    layer2_outputs(5538) <= a xor b;
    layer2_outputs(5539) <= not (a or b);
    layer2_outputs(5540) <= a or b;
    layer2_outputs(5541) <= not (a or b);
    layer2_outputs(5542) <= b and not a;
    layer2_outputs(5543) <= not b;
    layer2_outputs(5544) <= a;
    layer2_outputs(5545) <= not b or a;
    layer2_outputs(5546) <= not b;
    layer2_outputs(5547) <= b and not a;
    layer2_outputs(5548) <= not (a or b);
    layer2_outputs(5549) <= b;
    layer2_outputs(5550) <= not a;
    layer2_outputs(5551) <= b;
    layer2_outputs(5552) <= a;
    layer2_outputs(5553) <= a;
    layer2_outputs(5554) <= not b;
    layer2_outputs(5555) <= not a or b;
    layer2_outputs(5556) <= a and not b;
    layer2_outputs(5557) <= not (a and b);
    layer2_outputs(5558) <= not b;
    layer2_outputs(5559) <= not (a and b);
    layer2_outputs(5560) <= not (a xor b);
    layer2_outputs(5561) <= a or b;
    layer2_outputs(5562) <= a xor b;
    layer2_outputs(5563) <= b and not a;
    layer2_outputs(5564) <= not b or a;
    layer2_outputs(5565) <= a xor b;
    layer2_outputs(5566) <= not (a xor b);
    layer2_outputs(5567) <= a;
    layer2_outputs(5568) <= a and b;
    layer2_outputs(5569) <= b;
    layer2_outputs(5570) <= not b;
    layer2_outputs(5571) <= a;
    layer2_outputs(5572) <= b and not a;
    layer2_outputs(5573) <= b;
    layer2_outputs(5574) <= a;
    layer2_outputs(5575) <= a;
    layer2_outputs(5576) <= '0';
    layer2_outputs(5577) <= not a;
    layer2_outputs(5578) <= not b;
    layer2_outputs(5579) <= not b or a;
    layer2_outputs(5580) <= b;
    layer2_outputs(5581) <= a or b;
    layer2_outputs(5582) <= not b;
    layer2_outputs(5583) <= '1';
    layer2_outputs(5584) <= not b;
    layer2_outputs(5585) <= not a;
    layer2_outputs(5586) <= not a or b;
    layer2_outputs(5587) <= not b;
    layer2_outputs(5588) <= not b;
    layer2_outputs(5589) <= not (a xor b);
    layer2_outputs(5590) <= not (a xor b);
    layer2_outputs(5591) <= a xor b;
    layer2_outputs(5592) <= not (a and b);
    layer2_outputs(5593) <= a or b;
    layer2_outputs(5594) <= not (a or b);
    layer2_outputs(5595) <= b and not a;
    layer2_outputs(5596) <= not a or b;
    layer2_outputs(5597) <= not a;
    layer2_outputs(5598) <= not (a xor b);
    layer2_outputs(5599) <= not (a xor b);
    layer2_outputs(5600) <= not a;
    layer2_outputs(5601) <= not a or b;
    layer2_outputs(5602) <= not a;
    layer2_outputs(5603) <= a and b;
    layer2_outputs(5604) <= not a;
    layer2_outputs(5605) <= b;
    layer2_outputs(5606) <= a;
    layer2_outputs(5607) <= not b or a;
    layer2_outputs(5608) <= a xor b;
    layer2_outputs(5609) <= not a or b;
    layer2_outputs(5610) <= not b;
    layer2_outputs(5611) <= a and b;
    layer2_outputs(5612) <= a and not b;
    layer2_outputs(5613) <= a xor b;
    layer2_outputs(5614) <= not a or b;
    layer2_outputs(5615) <= not (a and b);
    layer2_outputs(5616) <= not (a and b);
    layer2_outputs(5617) <= b and not a;
    layer2_outputs(5618) <= a;
    layer2_outputs(5619) <= a or b;
    layer2_outputs(5620) <= a or b;
    layer2_outputs(5621) <= a and b;
    layer2_outputs(5622) <= not b or a;
    layer2_outputs(5623) <= a;
    layer2_outputs(5624) <= not a;
    layer2_outputs(5625) <= a or b;
    layer2_outputs(5626) <= a and not b;
    layer2_outputs(5627) <= b;
    layer2_outputs(5628) <= a;
    layer2_outputs(5629) <= a or b;
    layer2_outputs(5630) <= a and b;
    layer2_outputs(5631) <= a;
    layer2_outputs(5632) <= a xor b;
    layer2_outputs(5633) <= a xor b;
    layer2_outputs(5634) <= not (a or b);
    layer2_outputs(5635) <= not (a and b);
    layer2_outputs(5636) <= not b or a;
    layer2_outputs(5637) <= a xor b;
    layer2_outputs(5638) <= not b;
    layer2_outputs(5639) <= a or b;
    layer2_outputs(5640) <= not b;
    layer2_outputs(5641) <= not a;
    layer2_outputs(5642) <= a xor b;
    layer2_outputs(5643) <= not (a and b);
    layer2_outputs(5644) <= not a or b;
    layer2_outputs(5645) <= b;
    layer2_outputs(5646) <= not a or b;
    layer2_outputs(5647) <= not (a and b);
    layer2_outputs(5648) <= not (a or b);
    layer2_outputs(5649) <= a;
    layer2_outputs(5650) <= not (a or b);
    layer2_outputs(5651) <= a and b;
    layer2_outputs(5652) <= not a;
    layer2_outputs(5653) <= a and not b;
    layer2_outputs(5654) <= not a;
    layer2_outputs(5655) <= not a;
    layer2_outputs(5656) <= a;
    layer2_outputs(5657) <= not b or a;
    layer2_outputs(5658) <= not (a xor b);
    layer2_outputs(5659) <= '0';
    layer2_outputs(5660) <= a xor b;
    layer2_outputs(5661) <= not a or b;
    layer2_outputs(5662) <= a or b;
    layer2_outputs(5663) <= not (a xor b);
    layer2_outputs(5664) <= a and not b;
    layer2_outputs(5665) <= not (a or b);
    layer2_outputs(5666) <= not b;
    layer2_outputs(5667) <= a;
    layer2_outputs(5668) <= not b or a;
    layer2_outputs(5669) <= a;
    layer2_outputs(5670) <= not b;
    layer2_outputs(5671) <= not (a xor b);
    layer2_outputs(5672) <= b;
    layer2_outputs(5673) <= a and b;
    layer2_outputs(5674) <= not b;
    layer2_outputs(5675) <= not a or b;
    layer2_outputs(5676) <= a and b;
    layer2_outputs(5677) <= a or b;
    layer2_outputs(5678) <= a;
    layer2_outputs(5679) <= a and not b;
    layer2_outputs(5680) <= not (a xor b);
    layer2_outputs(5681) <= not a;
    layer2_outputs(5682) <= a;
    layer2_outputs(5683) <= not (a xor b);
    layer2_outputs(5684) <= a;
    layer2_outputs(5685) <= a;
    layer2_outputs(5686) <= not (a xor b);
    layer2_outputs(5687) <= not a;
    layer2_outputs(5688) <= b;
    layer2_outputs(5689) <= not a or b;
    layer2_outputs(5690) <= not a;
    layer2_outputs(5691) <= b;
    layer2_outputs(5692) <= not (a or b);
    layer2_outputs(5693) <= a;
    layer2_outputs(5694) <= not b or a;
    layer2_outputs(5695) <= not a or b;
    layer2_outputs(5696) <= not (a xor b);
    layer2_outputs(5697) <= not b or a;
    layer2_outputs(5698) <= a and not b;
    layer2_outputs(5699) <= not b;
    layer2_outputs(5700) <= not (a or b);
    layer2_outputs(5701) <= a and not b;
    layer2_outputs(5702) <= a;
    layer2_outputs(5703) <= a xor b;
    layer2_outputs(5704) <= a xor b;
    layer2_outputs(5705) <= a;
    layer2_outputs(5706) <= not b;
    layer2_outputs(5707) <= not b or a;
    layer2_outputs(5708) <= a;
    layer2_outputs(5709) <= a;
    layer2_outputs(5710) <= not (a or b);
    layer2_outputs(5711) <= not (a xor b);
    layer2_outputs(5712) <= a or b;
    layer2_outputs(5713) <= a;
    layer2_outputs(5714) <= not (a or b);
    layer2_outputs(5715) <= b;
    layer2_outputs(5716) <= b;
    layer2_outputs(5717) <= a or b;
    layer2_outputs(5718) <= not b or a;
    layer2_outputs(5719) <= a and not b;
    layer2_outputs(5720) <= not (a or b);
    layer2_outputs(5721) <= b and not a;
    layer2_outputs(5722) <= a xor b;
    layer2_outputs(5723) <= a xor b;
    layer2_outputs(5724) <= not (a or b);
    layer2_outputs(5725) <= '0';
    layer2_outputs(5726) <= not a;
    layer2_outputs(5727) <= not (a or b);
    layer2_outputs(5728) <= not (a or b);
    layer2_outputs(5729) <= a and b;
    layer2_outputs(5730) <= not b;
    layer2_outputs(5731) <= b;
    layer2_outputs(5732) <= a and not b;
    layer2_outputs(5733) <= a xor b;
    layer2_outputs(5734) <= not (a and b);
    layer2_outputs(5735) <= not b or a;
    layer2_outputs(5736) <= a;
    layer2_outputs(5737) <= not b or a;
    layer2_outputs(5738) <= b and not a;
    layer2_outputs(5739) <= a xor b;
    layer2_outputs(5740) <= b and not a;
    layer2_outputs(5741) <= a and not b;
    layer2_outputs(5742) <= b and not a;
    layer2_outputs(5743) <= b;
    layer2_outputs(5744) <= a;
    layer2_outputs(5745) <= a and b;
    layer2_outputs(5746) <= not a;
    layer2_outputs(5747) <= a xor b;
    layer2_outputs(5748) <= not a or b;
    layer2_outputs(5749) <= a xor b;
    layer2_outputs(5750) <= not (a and b);
    layer2_outputs(5751) <= a;
    layer2_outputs(5752) <= a and b;
    layer2_outputs(5753) <= not a;
    layer2_outputs(5754) <= not a;
    layer2_outputs(5755) <= b;
    layer2_outputs(5756) <= a;
    layer2_outputs(5757) <= not (a xor b);
    layer2_outputs(5758) <= a and not b;
    layer2_outputs(5759) <= a xor b;
    layer2_outputs(5760) <= not (a or b);
    layer2_outputs(5761) <= a and not b;
    layer2_outputs(5762) <= not (a xor b);
    layer2_outputs(5763) <= not b or a;
    layer2_outputs(5764) <= not a;
    layer2_outputs(5765) <= not (a or b);
    layer2_outputs(5766) <= not a;
    layer2_outputs(5767) <= a;
    layer2_outputs(5768) <= not a;
    layer2_outputs(5769) <= a and b;
    layer2_outputs(5770) <= a and b;
    layer2_outputs(5771) <= not (a and b);
    layer2_outputs(5772) <= not (a xor b);
    layer2_outputs(5773) <= not b or a;
    layer2_outputs(5774) <= a xor b;
    layer2_outputs(5775) <= a and b;
    layer2_outputs(5776) <= a;
    layer2_outputs(5777) <= not a;
    layer2_outputs(5778) <= a and not b;
    layer2_outputs(5779) <= not b;
    layer2_outputs(5780) <= b and not a;
    layer2_outputs(5781) <= b;
    layer2_outputs(5782) <= not b;
    layer2_outputs(5783) <= not b;
    layer2_outputs(5784) <= not b;
    layer2_outputs(5785) <= b and not a;
    layer2_outputs(5786) <= not (a and b);
    layer2_outputs(5787) <= b and not a;
    layer2_outputs(5788) <= b;
    layer2_outputs(5789) <= not a;
    layer2_outputs(5790) <= not a;
    layer2_outputs(5791) <= a;
    layer2_outputs(5792) <= not (a and b);
    layer2_outputs(5793) <= not a or b;
    layer2_outputs(5794) <= not b;
    layer2_outputs(5795) <= not b;
    layer2_outputs(5796) <= a or b;
    layer2_outputs(5797) <= b;
    layer2_outputs(5798) <= not (a xor b);
    layer2_outputs(5799) <= not a;
    layer2_outputs(5800) <= not b;
    layer2_outputs(5801) <= b;
    layer2_outputs(5802) <= b;
    layer2_outputs(5803) <= not (a xor b);
    layer2_outputs(5804) <= b and not a;
    layer2_outputs(5805) <= not a;
    layer2_outputs(5806) <= not b or a;
    layer2_outputs(5807) <= not a;
    layer2_outputs(5808) <= b and not a;
    layer2_outputs(5809) <= not b or a;
    layer2_outputs(5810) <= not a or b;
    layer2_outputs(5811) <= a xor b;
    layer2_outputs(5812) <= a and b;
    layer2_outputs(5813) <= not b;
    layer2_outputs(5814) <= a xor b;
    layer2_outputs(5815) <= not (a xor b);
    layer2_outputs(5816) <= not b or a;
    layer2_outputs(5817) <= not (a xor b);
    layer2_outputs(5818) <= not a;
    layer2_outputs(5819) <= not b;
    layer2_outputs(5820) <= not a or b;
    layer2_outputs(5821) <= b and not a;
    layer2_outputs(5822) <= a xor b;
    layer2_outputs(5823) <= b;
    layer2_outputs(5824) <= not a;
    layer2_outputs(5825) <= not (a and b);
    layer2_outputs(5826) <= not a;
    layer2_outputs(5827) <= not b or a;
    layer2_outputs(5828) <= b;
    layer2_outputs(5829) <= b and not a;
    layer2_outputs(5830) <= not (a xor b);
    layer2_outputs(5831) <= a or b;
    layer2_outputs(5832) <= not (a and b);
    layer2_outputs(5833) <= not a;
    layer2_outputs(5834) <= a and not b;
    layer2_outputs(5835) <= not b or a;
    layer2_outputs(5836) <= not (a xor b);
    layer2_outputs(5837) <= not (a or b);
    layer2_outputs(5838) <= a or b;
    layer2_outputs(5839) <= not b or a;
    layer2_outputs(5840) <= not (a xor b);
    layer2_outputs(5841) <= a;
    layer2_outputs(5842) <= a;
    layer2_outputs(5843) <= not a;
    layer2_outputs(5844) <= a and b;
    layer2_outputs(5845) <= not a;
    layer2_outputs(5846) <= a xor b;
    layer2_outputs(5847) <= a and b;
    layer2_outputs(5848) <= not a;
    layer2_outputs(5849) <= not (a xor b);
    layer2_outputs(5850) <= b;
    layer2_outputs(5851) <= a;
    layer2_outputs(5852) <= a;
    layer2_outputs(5853) <= not (a xor b);
    layer2_outputs(5854) <= a xor b;
    layer2_outputs(5855) <= not b;
    layer2_outputs(5856) <= not a or b;
    layer2_outputs(5857) <= b;
    layer2_outputs(5858) <= not b;
    layer2_outputs(5859) <= not (a and b);
    layer2_outputs(5860) <= not (a xor b);
    layer2_outputs(5861) <= not (a xor b);
    layer2_outputs(5862) <= not a or b;
    layer2_outputs(5863) <= b;
    layer2_outputs(5864) <= a and b;
    layer2_outputs(5865) <= not b;
    layer2_outputs(5866) <= b and not a;
    layer2_outputs(5867) <= not (a and b);
    layer2_outputs(5868) <= not a;
    layer2_outputs(5869) <= not (a xor b);
    layer2_outputs(5870) <= not a;
    layer2_outputs(5871) <= b and not a;
    layer2_outputs(5872) <= a;
    layer2_outputs(5873) <= not a;
    layer2_outputs(5874) <= '1';
    layer2_outputs(5875) <= a and b;
    layer2_outputs(5876) <= not (a xor b);
    layer2_outputs(5877) <= b;
    layer2_outputs(5878) <= not (a and b);
    layer2_outputs(5879) <= not (a xor b);
    layer2_outputs(5880) <= b;
    layer2_outputs(5881) <= not b;
    layer2_outputs(5882) <= a and b;
    layer2_outputs(5883) <= not a;
    layer2_outputs(5884) <= b;
    layer2_outputs(5885) <= a xor b;
    layer2_outputs(5886) <= b;
    layer2_outputs(5887) <= a and not b;
    layer2_outputs(5888) <= not a or b;
    layer2_outputs(5889) <= not b or a;
    layer2_outputs(5890) <= b and not a;
    layer2_outputs(5891) <= not a;
    layer2_outputs(5892) <= a and not b;
    layer2_outputs(5893) <= not (a xor b);
    layer2_outputs(5894) <= a xor b;
    layer2_outputs(5895) <= not (a xor b);
    layer2_outputs(5896) <= not a;
    layer2_outputs(5897) <= a;
    layer2_outputs(5898) <= a xor b;
    layer2_outputs(5899) <= not a;
    layer2_outputs(5900) <= a or b;
    layer2_outputs(5901) <= b;
    layer2_outputs(5902) <= not (a and b);
    layer2_outputs(5903) <= a and b;
    layer2_outputs(5904) <= not (a or b);
    layer2_outputs(5905) <= not (a or b);
    layer2_outputs(5906) <= a and b;
    layer2_outputs(5907) <= b and not a;
    layer2_outputs(5908) <= not (a and b);
    layer2_outputs(5909) <= b and not a;
    layer2_outputs(5910) <= a;
    layer2_outputs(5911) <= a xor b;
    layer2_outputs(5912) <= b;
    layer2_outputs(5913) <= a and b;
    layer2_outputs(5914) <= a xor b;
    layer2_outputs(5915) <= a or b;
    layer2_outputs(5916) <= not (a or b);
    layer2_outputs(5917) <= a;
    layer2_outputs(5918) <= b and not a;
    layer2_outputs(5919) <= a;
    layer2_outputs(5920) <= not (a xor b);
    layer2_outputs(5921) <= a xor b;
    layer2_outputs(5922) <= '1';
    layer2_outputs(5923) <= a;
    layer2_outputs(5924) <= b;
    layer2_outputs(5925) <= b;
    layer2_outputs(5926) <= not (a or b);
    layer2_outputs(5927) <= not b;
    layer2_outputs(5928) <= a and b;
    layer2_outputs(5929) <= not b or a;
    layer2_outputs(5930) <= not (a or b);
    layer2_outputs(5931) <= not (a xor b);
    layer2_outputs(5932) <= not b;
    layer2_outputs(5933) <= a and b;
    layer2_outputs(5934) <= not (a or b);
    layer2_outputs(5935) <= not (a and b);
    layer2_outputs(5936) <= not a;
    layer2_outputs(5937) <= not (a and b);
    layer2_outputs(5938) <= not (a xor b);
    layer2_outputs(5939) <= not (a xor b);
    layer2_outputs(5940) <= not b;
    layer2_outputs(5941) <= a and not b;
    layer2_outputs(5942) <= not b;
    layer2_outputs(5943) <= not (a and b);
    layer2_outputs(5944) <= a;
    layer2_outputs(5945) <= not b;
    layer2_outputs(5946) <= not b or a;
    layer2_outputs(5947) <= a;
    layer2_outputs(5948) <= not (a and b);
    layer2_outputs(5949) <= a or b;
    layer2_outputs(5950) <= not b or a;
    layer2_outputs(5951) <= not b or a;
    layer2_outputs(5952) <= not a;
    layer2_outputs(5953) <= not b;
    layer2_outputs(5954) <= not b;
    layer2_outputs(5955) <= not (a or b);
    layer2_outputs(5956) <= a;
    layer2_outputs(5957) <= b and not a;
    layer2_outputs(5958) <= a and not b;
    layer2_outputs(5959) <= a or b;
    layer2_outputs(5960) <= not (a xor b);
    layer2_outputs(5961) <= not a;
    layer2_outputs(5962) <= not b or a;
    layer2_outputs(5963) <= not (a xor b);
    layer2_outputs(5964) <= a xor b;
    layer2_outputs(5965) <= not a;
    layer2_outputs(5966) <= not b;
    layer2_outputs(5967) <= not a;
    layer2_outputs(5968) <= b and not a;
    layer2_outputs(5969) <= not (a and b);
    layer2_outputs(5970) <= not (a or b);
    layer2_outputs(5971) <= not (a and b);
    layer2_outputs(5972) <= not a or b;
    layer2_outputs(5973) <= '1';
    layer2_outputs(5974) <= not a;
    layer2_outputs(5975) <= a;
    layer2_outputs(5976) <= not a or b;
    layer2_outputs(5977) <= a and not b;
    layer2_outputs(5978) <= a xor b;
    layer2_outputs(5979) <= not b;
    layer2_outputs(5980) <= a xor b;
    layer2_outputs(5981) <= not (a xor b);
    layer2_outputs(5982) <= a;
    layer2_outputs(5983) <= a;
    layer2_outputs(5984) <= a and not b;
    layer2_outputs(5985) <= a and not b;
    layer2_outputs(5986) <= b;
    layer2_outputs(5987) <= not a;
    layer2_outputs(5988) <= b and not a;
    layer2_outputs(5989) <= not a;
    layer2_outputs(5990) <= b;
    layer2_outputs(5991) <= not a;
    layer2_outputs(5992) <= not a;
    layer2_outputs(5993) <= not (a xor b);
    layer2_outputs(5994) <= a and not b;
    layer2_outputs(5995) <= a;
    layer2_outputs(5996) <= b;
    layer2_outputs(5997) <= a;
    layer2_outputs(5998) <= not (a xor b);
    layer2_outputs(5999) <= not b;
    layer2_outputs(6000) <= not a or b;
    layer2_outputs(6001) <= not b or a;
    layer2_outputs(6002) <= not a;
    layer2_outputs(6003) <= not b;
    layer2_outputs(6004) <= b and not a;
    layer2_outputs(6005) <= a xor b;
    layer2_outputs(6006) <= not a;
    layer2_outputs(6007) <= not a;
    layer2_outputs(6008) <= a and not b;
    layer2_outputs(6009) <= not a or b;
    layer2_outputs(6010) <= '1';
    layer2_outputs(6011) <= not b;
    layer2_outputs(6012) <= a xor b;
    layer2_outputs(6013) <= not b;
    layer2_outputs(6014) <= not b;
    layer2_outputs(6015) <= not a or b;
    layer2_outputs(6016) <= not a or b;
    layer2_outputs(6017) <= a xor b;
    layer2_outputs(6018) <= a or b;
    layer2_outputs(6019) <= a xor b;
    layer2_outputs(6020) <= a xor b;
    layer2_outputs(6021) <= not b;
    layer2_outputs(6022) <= a xor b;
    layer2_outputs(6023) <= b;
    layer2_outputs(6024) <= b;
    layer2_outputs(6025) <= a and not b;
    layer2_outputs(6026) <= not b;
    layer2_outputs(6027) <= not (a or b);
    layer2_outputs(6028) <= not a;
    layer2_outputs(6029) <= not a;
    layer2_outputs(6030) <= not (a xor b);
    layer2_outputs(6031) <= not b or a;
    layer2_outputs(6032) <= a xor b;
    layer2_outputs(6033) <= a xor b;
    layer2_outputs(6034) <= a and not b;
    layer2_outputs(6035) <= a and not b;
    layer2_outputs(6036) <= not (a and b);
    layer2_outputs(6037) <= a;
    layer2_outputs(6038) <= not (a or b);
    layer2_outputs(6039) <= b;
    layer2_outputs(6040) <= a;
    layer2_outputs(6041) <= a xor b;
    layer2_outputs(6042) <= a xor b;
    layer2_outputs(6043) <= not b;
    layer2_outputs(6044) <= b and not a;
    layer2_outputs(6045) <= a;
    layer2_outputs(6046) <= not (a xor b);
    layer2_outputs(6047) <= a or b;
    layer2_outputs(6048) <= not a or b;
    layer2_outputs(6049) <= a;
    layer2_outputs(6050) <= a xor b;
    layer2_outputs(6051) <= not (a or b);
    layer2_outputs(6052) <= not (a xor b);
    layer2_outputs(6053) <= not (a xor b);
    layer2_outputs(6054) <= not a;
    layer2_outputs(6055) <= not a;
    layer2_outputs(6056) <= not b;
    layer2_outputs(6057) <= b;
    layer2_outputs(6058) <= not b;
    layer2_outputs(6059) <= not a or b;
    layer2_outputs(6060) <= not a;
    layer2_outputs(6061) <= not a;
    layer2_outputs(6062) <= not a;
    layer2_outputs(6063) <= not b or a;
    layer2_outputs(6064) <= a and b;
    layer2_outputs(6065) <= not a or b;
    layer2_outputs(6066) <= a and b;
    layer2_outputs(6067) <= not b;
    layer2_outputs(6068) <= a and b;
    layer2_outputs(6069) <= b and not a;
    layer2_outputs(6070) <= not (a xor b);
    layer2_outputs(6071) <= a xor b;
    layer2_outputs(6072) <= not a;
    layer2_outputs(6073) <= not b;
    layer2_outputs(6074) <= not (a xor b);
    layer2_outputs(6075) <= a and b;
    layer2_outputs(6076) <= not (a xor b);
    layer2_outputs(6077) <= not a;
    layer2_outputs(6078) <= not b;
    layer2_outputs(6079) <= not b;
    layer2_outputs(6080) <= not a;
    layer2_outputs(6081) <= not (a and b);
    layer2_outputs(6082) <= a or b;
    layer2_outputs(6083) <= b and not a;
    layer2_outputs(6084) <= not (a or b);
    layer2_outputs(6085) <= not a or b;
    layer2_outputs(6086) <= not (a and b);
    layer2_outputs(6087) <= not (a or b);
    layer2_outputs(6088) <= not (a xor b);
    layer2_outputs(6089) <= a and not b;
    layer2_outputs(6090) <= not b or a;
    layer2_outputs(6091) <= a and b;
    layer2_outputs(6092) <= not a or b;
    layer2_outputs(6093) <= not b or a;
    layer2_outputs(6094) <= not a or b;
    layer2_outputs(6095) <= not a;
    layer2_outputs(6096) <= not a;
    layer2_outputs(6097) <= not b or a;
    layer2_outputs(6098) <= a;
    layer2_outputs(6099) <= not (a and b);
    layer2_outputs(6100) <= a;
    layer2_outputs(6101) <= not (a xor b);
    layer2_outputs(6102) <= not b or a;
    layer2_outputs(6103) <= a xor b;
    layer2_outputs(6104) <= a;
    layer2_outputs(6105) <= not (a xor b);
    layer2_outputs(6106) <= a xor b;
    layer2_outputs(6107) <= a or b;
    layer2_outputs(6108) <= not (a xor b);
    layer2_outputs(6109) <= a;
    layer2_outputs(6110) <= a or b;
    layer2_outputs(6111) <= not (a or b);
    layer2_outputs(6112) <= not a;
    layer2_outputs(6113) <= not b;
    layer2_outputs(6114) <= not (a xor b);
    layer2_outputs(6115) <= not b;
    layer2_outputs(6116) <= a xor b;
    layer2_outputs(6117) <= b;
    layer2_outputs(6118) <= not a;
    layer2_outputs(6119) <= not b;
    layer2_outputs(6120) <= not (a xor b);
    layer2_outputs(6121) <= not (a or b);
    layer2_outputs(6122) <= not a;
    layer2_outputs(6123) <= a and b;
    layer2_outputs(6124) <= b and not a;
    layer2_outputs(6125) <= a xor b;
    layer2_outputs(6126) <= not (a xor b);
    layer2_outputs(6127) <= not (a and b);
    layer2_outputs(6128) <= b;
    layer2_outputs(6129) <= not b or a;
    layer2_outputs(6130) <= a;
    layer2_outputs(6131) <= not b;
    layer2_outputs(6132) <= a or b;
    layer2_outputs(6133) <= not b or a;
    layer2_outputs(6134) <= b;
    layer2_outputs(6135) <= a and b;
    layer2_outputs(6136) <= not (a xor b);
    layer2_outputs(6137) <= a xor b;
    layer2_outputs(6138) <= not (a xor b);
    layer2_outputs(6139) <= not b;
    layer2_outputs(6140) <= b;
    layer2_outputs(6141) <= not a;
    layer2_outputs(6142) <= not a;
    layer2_outputs(6143) <= b;
    layer2_outputs(6144) <= not b or a;
    layer2_outputs(6145) <= b;
    layer2_outputs(6146) <= b;
    layer2_outputs(6147) <= not (a or b);
    layer2_outputs(6148) <= b;
    layer2_outputs(6149) <= not b or a;
    layer2_outputs(6150) <= a;
    layer2_outputs(6151) <= not (a and b);
    layer2_outputs(6152) <= not a;
    layer2_outputs(6153) <= not a;
    layer2_outputs(6154) <= not (a xor b);
    layer2_outputs(6155) <= b;
    layer2_outputs(6156) <= a or b;
    layer2_outputs(6157) <= not (a xor b);
    layer2_outputs(6158) <= b;
    layer2_outputs(6159) <= a;
    layer2_outputs(6160) <= not b;
    layer2_outputs(6161) <= not (a and b);
    layer2_outputs(6162) <= not (a xor b);
    layer2_outputs(6163) <= not (a xor b);
    layer2_outputs(6164) <= not (a and b);
    layer2_outputs(6165) <= b and not a;
    layer2_outputs(6166) <= a;
    layer2_outputs(6167) <= not a;
    layer2_outputs(6168) <= a and b;
    layer2_outputs(6169) <= not a;
    layer2_outputs(6170) <= a and not b;
    layer2_outputs(6171) <= not a or b;
    layer2_outputs(6172) <= a xor b;
    layer2_outputs(6173) <= a and b;
    layer2_outputs(6174) <= not (a xor b);
    layer2_outputs(6175) <= a and not b;
    layer2_outputs(6176) <= b;
    layer2_outputs(6177) <= not b;
    layer2_outputs(6178) <= a xor b;
    layer2_outputs(6179) <= not a or b;
    layer2_outputs(6180) <= a xor b;
    layer2_outputs(6181) <= a;
    layer2_outputs(6182) <= b;
    layer2_outputs(6183) <= not b or a;
    layer2_outputs(6184) <= a or b;
    layer2_outputs(6185) <= not a;
    layer2_outputs(6186) <= not (a and b);
    layer2_outputs(6187) <= a or b;
    layer2_outputs(6188) <= a and b;
    layer2_outputs(6189) <= b and not a;
    layer2_outputs(6190) <= not a;
    layer2_outputs(6191) <= b;
    layer2_outputs(6192) <= not (a xor b);
    layer2_outputs(6193) <= b and not a;
    layer2_outputs(6194) <= not b;
    layer2_outputs(6195) <= a and not b;
    layer2_outputs(6196) <= a xor b;
    layer2_outputs(6197) <= not b;
    layer2_outputs(6198) <= b;
    layer2_outputs(6199) <= b;
    layer2_outputs(6200) <= a xor b;
    layer2_outputs(6201) <= a and not b;
    layer2_outputs(6202) <= a and not b;
    layer2_outputs(6203) <= b;
    layer2_outputs(6204) <= not a or b;
    layer2_outputs(6205) <= not (a or b);
    layer2_outputs(6206) <= a xor b;
    layer2_outputs(6207) <= not b or a;
    layer2_outputs(6208) <= not (a or b);
    layer2_outputs(6209) <= not b;
    layer2_outputs(6210) <= a and not b;
    layer2_outputs(6211) <= not (a and b);
    layer2_outputs(6212) <= b;
    layer2_outputs(6213) <= not b;
    layer2_outputs(6214) <= not (a and b);
    layer2_outputs(6215) <= not (a and b);
    layer2_outputs(6216) <= not (a and b);
    layer2_outputs(6217) <= a or b;
    layer2_outputs(6218) <= not (a xor b);
    layer2_outputs(6219) <= b;
    layer2_outputs(6220) <= not (a and b);
    layer2_outputs(6221) <= not a;
    layer2_outputs(6222) <= not b;
    layer2_outputs(6223) <= b;
    layer2_outputs(6224) <= not b;
    layer2_outputs(6225) <= b and not a;
    layer2_outputs(6226) <= not a;
    layer2_outputs(6227) <= a and not b;
    layer2_outputs(6228) <= not a;
    layer2_outputs(6229) <= b;
    layer2_outputs(6230) <= a;
    layer2_outputs(6231) <= a;
    layer2_outputs(6232) <= not (a and b);
    layer2_outputs(6233) <= not (a and b);
    layer2_outputs(6234) <= not a;
    layer2_outputs(6235) <= not a;
    layer2_outputs(6236) <= not b;
    layer2_outputs(6237) <= a;
    layer2_outputs(6238) <= a and b;
    layer2_outputs(6239) <= not (a xor b);
    layer2_outputs(6240) <= a;
    layer2_outputs(6241) <= b;
    layer2_outputs(6242) <= a xor b;
    layer2_outputs(6243) <= not a;
    layer2_outputs(6244) <= a or b;
    layer2_outputs(6245) <= a or b;
    layer2_outputs(6246) <= not (a xor b);
    layer2_outputs(6247) <= not a or b;
    layer2_outputs(6248) <= a;
    layer2_outputs(6249) <= b and not a;
    layer2_outputs(6250) <= not (a and b);
    layer2_outputs(6251) <= a xor b;
    layer2_outputs(6252) <= not a;
    layer2_outputs(6253) <= not a or b;
    layer2_outputs(6254) <= b;
    layer2_outputs(6255) <= a and b;
    layer2_outputs(6256) <= a or b;
    layer2_outputs(6257) <= a;
    layer2_outputs(6258) <= b;
    layer2_outputs(6259) <= not a;
    layer2_outputs(6260) <= not b;
    layer2_outputs(6261) <= '0';
    layer2_outputs(6262) <= not (a xor b);
    layer2_outputs(6263) <= '0';
    layer2_outputs(6264) <= not b;
    layer2_outputs(6265) <= not a or b;
    layer2_outputs(6266) <= a;
    layer2_outputs(6267) <= a or b;
    layer2_outputs(6268) <= not (a and b);
    layer2_outputs(6269) <= not (a xor b);
    layer2_outputs(6270) <= a and b;
    layer2_outputs(6271) <= a and not b;
    layer2_outputs(6272) <= a or b;
    layer2_outputs(6273) <= b;
    layer2_outputs(6274) <= not b;
    layer2_outputs(6275) <= a xor b;
    layer2_outputs(6276) <= a;
    layer2_outputs(6277) <= not a or b;
    layer2_outputs(6278) <= b;
    layer2_outputs(6279) <= not a;
    layer2_outputs(6280) <= a;
    layer2_outputs(6281) <= b and not a;
    layer2_outputs(6282) <= not a;
    layer2_outputs(6283) <= b;
    layer2_outputs(6284) <= not (a or b);
    layer2_outputs(6285) <= not b;
    layer2_outputs(6286) <= a and not b;
    layer2_outputs(6287) <= not (a and b);
    layer2_outputs(6288) <= b;
    layer2_outputs(6289) <= b;
    layer2_outputs(6290) <= '1';
    layer2_outputs(6291) <= b;
    layer2_outputs(6292) <= not b or a;
    layer2_outputs(6293) <= not a;
    layer2_outputs(6294) <= not b or a;
    layer2_outputs(6295) <= not (a xor b);
    layer2_outputs(6296) <= not a;
    layer2_outputs(6297) <= not (a or b);
    layer2_outputs(6298) <= a;
    layer2_outputs(6299) <= b;
    layer2_outputs(6300) <= not (a or b);
    layer2_outputs(6301) <= b;
    layer2_outputs(6302) <= not b or a;
    layer2_outputs(6303) <= not b;
    layer2_outputs(6304) <= not b;
    layer2_outputs(6305) <= not (a xor b);
    layer2_outputs(6306) <= a xor b;
    layer2_outputs(6307) <= a and b;
    layer2_outputs(6308) <= a and not b;
    layer2_outputs(6309) <= a and not b;
    layer2_outputs(6310) <= not (a and b);
    layer2_outputs(6311) <= not (a or b);
    layer2_outputs(6312) <= not (a xor b);
    layer2_outputs(6313) <= a xor b;
    layer2_outputs(6314) <= not a;
    layer2_outputs(6315) <= a xor b;
    layer2_outputs(6316) <= not a;
    layer2_outputs(6317) <= a and b;
    layer2_outputs(6318) <= not b;
    layer2_outputs(6319) <= a or b;
    layer2_outputs(6320) <= not a;
    layer2_outputs(6321) <= a and b;
    layer2_outputs(6322) <= a or b;
    layer2_outputs(6323) <= not b;
    layer2_outputs(6324) <= not b;
    layer2_outputs(6325) <= not b or a;
    layer2_outputs(6326) <= a xor b;
    layer2_outputs(6327) <= not b or a;
    layer2_outputs(6328) <= not b;
    layer2_outputs(6329) <= not b or a;
    layer2_outputs(6330) <= not a;
    layer2_outputs(6331) <= b;
    layer2_outputs(6332) <= a and not b;
    layer2_outputs(6333) <= a xor b;
    layer2_outputs(6334) <= not a;
    layer2_outputs(6335) <= not (a xor b);
    layer2_outputs(6336) <= not b or a;
    layer2_outputs(6337) <= a;
    layer2_outputs(6338) <= not a or b;
    layer2_outputs(6339) <= not (a xor b);
    layer2_outputs(6340) <= not a or b;
    layer2_outputs(6341) <= not (a and b);
    layer2_outputs(6342) <= b;
    layer2_outputs(6343) <= a;
    layer2_outputs(6344) <= not (a and b);
    layer2_outputs(6345) <= b;
    layer2_outputs(6346) <= a and not b;
    layer2_outputs(6347) <= not a or b;
    layer2_outputs(6348) <= a xor b;
    layer2_outputs(6349) <= a;
    layer2_outputs(6350) <= b;
    layer2_outputs(6351) <= b;
    layer2_outputs(6352) <= not (a xor b);
    layer2_outputs(6353) <= not (a xor b);
    layer2_outputs(6354) <= not (a or b);
    layer2_outputs(6355) <= a;
    layer2_outputs(6356) <= a and not b;
    layer2_outputs(6357) <= a and not b;
    layer2_outputs(6358) <= b;
    layer2_outputs(6359) <= a or b;
    layer2_outputs(6360) <= b and not a;
    layer2_outputs(6361) <= not b;
    layer2_outputs(6362) <= a xor b;
    layer2_outputs(6363) <= not (a xor b);
    layer2_outputs(6364) <= not (a or b);
    layer2_outputs(6365) <= not (a and b);
    layer2_outputs(6366) <= a;
    layer2_outputs(6367) <= not (a or b);
    layer2_outputs(6368) <= not (a and b);
    layer2_outputs(6369) <= not a;
    layer2_outputs(6370) <= b and not a;
    layer2_outputs(6371) <= a and not b;
    layer2_outputs(6372) <= a;
    layer2_outputs(6373) <= not b;
    layer2_outputs(6374) <= a and b;
    layer2_outputs(6375) <= not b or a;
    layer2_outputs(6376) <= b and not a;
    layer2_outputs(6377) <= a;
    layer2_outputs(6378) <= b;
    layer2_outputs(6379) <= a xor b;
    layer2_outputs(6380) <= not b or a;
    layer2_outputs(6381) <= not a or b;
    layer2_outputs(6382) <= not b or a;
    layer2_outputs(6383) <= not (a xor b);
    layer2_outputs(6384) <= not (a xor b);
    layer2_outputs(6385) <= not b;
    layer2_outputs(6386) <= not a or b;
    layer2_outputs(6387) <= not b;
    layer2_outputs(6388) <= a or b;
    layer2_outputs(6389) <= b;
    layer2_outputs(6390) <= b and not a;
    layer2_outputs(6391) <= a xor b;
    layer2_outputs(6392) <= a and not b;
    layer2_outputs(6393) <= not a;
    layer2_outputs(6394) <= not b;
    layer2_outputs(6395) <= not (a xor b);
    layer2_outputs(6396) <= a;
    layer2_outputs(6397) <= not (a or b);
    layer2_outputs(6398) <= not a;
    layer2_outputs(6399) <= a xor b;
    layer2_outputs(6400) <= not b;
    layer2_outputs(6401) <= '0';
    layer2_outputs(6402) <= not (a xor b);
    layer2_outputs(6403) <= a xor b;
    layer2_outputs(6404) <= not (a xor b);
    layer2_outputs(6405) <= a;
    layer2_outputs(6406) <= b;
    layer2_outputs(6407) <= not (a or b);
    layer2_outputs(6408) <= not b;
    layer2_outputs(6409) <= not (a and b);
    layer2_outputs(6410) <= a;
    layer2_outputs(6411) <= '1';
    layer2_outputs(6412) <= not (a and b);
    layer2_outputs(6413) <= not b;
    layer2_outputs(6414) <= not (a xor b);
    layer2_outputs(6415) <= b and not a;
    layer2_outputs(6416) <= not (a or b);
    layer2_outputs(6417) <= a and b;
    layer2_outputs(6418) <= a or b;
    layer2_outputs(6419) <= not (a and b);
    layer2_outputs(6420) <= a and not b;
    layer2_outputs(6421) <= not (a xor b);
    layer2_outputs(6422) <= not b;
    layer2_outputs(6423) <= a;
    layer2_outputs(6424) <= a;
    layer2_outputs(6425) <= a;
    layer2_outputs(6426) <= not a;
    layer2_outputs(6427) <= not a;
    layer2_outputs(6428) <= not (a or b);
    layer2_outputs(6429) <= not a;
    layer2_outputs(6430) <= a and not b;
    layer2_outputs(6431) <= not a;
    layer2_outputs(6432) <= not (a and b);
    layer2_outputs(6433) <= not (a xor b);
    layer2_outputs(6434) <= not b;
    layer2_outputs(6435) <= not (a or b);
    layer2_outputs(6436) <= not b;
    layer2_outputs(6437) <= not a;
    layer2_outputs(6438) <= not a;
    layer2_outputs(6439) <= not b;
    layer2_outputs(6440) <= not b;
    layer2_outputs(6441) <= not (a xor b);
    layer2_outputs(6442) <= b;
    layer2_outputs(6443) <= a and not b;
    layer2_outputs(6444) <= b;
    layer2_outputs(6445) <= b;
    layer2_outputs(6446) <= a and b;
    layer2_outputs(6447) <= b;
    layer2_outputs(6448) <= a;
    layer2_outputs(6449) <= b and not a;
    layer2_outputs(6450) <= a xor b;
    layer2_outputs(6451) <= a;
    layer2_outputs(6452) <= a and b;
    layer2_outputs(6453) <= not a;
    layer2_outputs(6454) <= not b;
    layer2_outputs(6455) <= not (a xor b);
    layer2_outputs(6456) <= not a or b;
    layer2_outputs(6457) <= a and not b;
    layer2_outputs(6458) <= not a;
    layer2_outputs(6459) <= a and not b;
    layer2_outputs(6460) <= a or b;
    layer2_outputs(6461) <= not a;
    layer2_outputs(6462) <= not (a xor b);
    layer2_outputs(6463) <= b and not a;
    layer2_outputs(6464) <= b and not a;
    layer2_outputs(6465) <= b;
    layer2_outputs(6466) <= not (a xor b);
    layer2_outputs(6467) <= not (a and b);
    layer2_outputs(6468) <= a xor b;
    layer2_outputs(6469) <= not (a and b);
    layer2_outputs(6470) <= a and b;
    layer2_outputs(6471) <= a or b;
    layer2_outputs(6472) <= not (a xor b);
    layer2_outputs(6473) <= '0';
    layer2_outputs(6474) <= not a;
    layer2_outputs(6475) <= not a;
    layer2_outputs(6476) <= a or b;
    layer2_outputs(6477) <= not b or a;
    layer2_outputs(6478) <= b and not a;
    layer2_outputs(6479) <= a;
    layer2_outputs(6480) <= not a;
    layer2_outputs(6481) <= not (a xor b);
    layer2_outputs(6482) <= a;
    layer2_outputs(6483) <= not a;
    layer2_outputs(6484) <= not (a xor b);
    layer2_outputs(6485) <= a;
    layer2_outputs(6486) <= a and not b;
    layer2_outputs(6487) <= not a;
    layer2_outputs(6488) <= a;
    layer2_outputs(6489) <= a;
    layer2_outputs(6490) <= b;
    layer2_outputs(6491) <= not (a or b);
    layer2_outputs(6492) <= a and b;
    layer2_outputs(6493) <= not a;
    layer2_outputs(6494) <= not a or b;
    layer2_outputs(6495) <= not b;
    layer2_outputs(6496) <= not a;
    layer2_outputs(6497) <= not b or a;
    layer2_outputs(6498) <= a xor b;
    layer2_outputs(6499) <= not (a xor b);
    layer2_outputs(6500) <= a xor b;
    layer2_outputs(6501) <= a and b;
    layer2_outputs(6502) <= a xor b;
    layer2_outputs(6503) <= not (a xor b);
    layer2_outputs(6504) <= not a or b;
    layer2_outputs(6505) <= b and not a;
    layer2_outputs(6506) <= not a;
    layer2_outputs(6507) <= a xor b;
    layer2_outputs(6508) <= not (a and b);
    layer2_outputs(6509) <= b and not a;
    layer2_outputs(6510) <= b and not a;
    layer2_outputs(6511) <= not a or b;
    layer2_outputs(6512) <= b;
    layer2_outputs(6513) <= not (a or b);
    layer2_outputs(6514) <= b and not a;
    layer2_outputs(6515) <= not a;
    layer2_outputs(6516) <= not b;
    layer2_outputs(6517) <= not a;
    layer2_outputs(6518) <= a;
    layer2_outputs(6519) <= not (a xor b);
    layer2_outputs(6520) <= not b;
    layer2_outputs(6521) <= not (a xor b);
    layer2_outputs(6522) <= not a or b;
    layer2_outputs(6523) <= b;
    layer2_outputs(6524) <= a xor b;
    layer2_outputs(6525) <= b and not a;
    layer2_outputs(6526) <= not (a and b);
    layer2_outputs(6527) <= b and not a;
    layer2_outputs(6528) <= not (a and b);
    layer2_outputs(6529) <= not a;
    layer2_outputs(6530) <= not (a and b);
    layer2_outputs(6531) <= a;
    layer2_outputs(6532) <= not (a xor b);
    layer2_outputs(6533) <= a;
    layer2_outputs(6534) <= not b;
    layer2_outputs(6535) <= not (a xor b);
    layer2_outputs(6536) <= b;
    layer2_outputs(6537) <= a and b;
    layer2_outputs(6538) <= b;
    layer2_outputs(6539) <= not b or a;
    layer2_outputs(6540) <= a;
    layer2_outputs(6541) <= not (a and b);
    layer2_outputs(6542) <= a and not b;
    layer2_outputs(6543) <= not b;
    layer2_outputs(6544) <= a and not b;
    layer2_outputs(6545) <= b;
    layer2_outputs(6546) <= not a;
    layer2_outputs(6547) <= a xor b;
    layer2_outputs(6548) <= not (a xor b);
    layer2_outputs(6549) <= a and not b;
    layer2_outputs(6550) <= not b;
    layer2_outputs(6551) <= a and not b;
    layer2_outputs(6552) <= not (a and b);
    layer2_outputs(6553) <= '1';
    layer2_outputs(6554) <= a;
    layer2_outputs(6555) <= b and not a;
    layer2_outputs(6556) <= a xor b;
    layer2_outputs(6557) <= a or b;
    layer2_outputs(6558) <= not a;
    layer2_outputs(6559) <= b and not a;
    layer2_outputs(6560) <= a and not b;
    layer2_outputs(6561) <= not (a or b);
    layer2_outputs(6562) <= not b or a;
    layer2_outputs(6563) <= a and not b;
    layer2_outputs(6564) <= not b;
    layer2_outputs(6565) <= a and not b;
    layer2_outputs(6566) <= not b;
    layer2_outputs(6567) <= not (a or b);
    layer2_outputs(6568) <= a xor b;
    layer2_outputs(6569) <= a xor b;
    layer2_outputs(6570) <= a and not b;
    layer2_outputs(6571) <= not (a and b);
    layer2_outputs(6572) <= b;
    layer2_outputs(6573) <= not (a or b);
    layer2_outputs(6574) <= not (a and b);
    layer2_outputs(6575) <= a and not b;
    layer2_outputs(6576) <= not b or a;
    layer2_outputs(6577) <= not (a xor b);
    layer2_outputs(6578) <= not b;
    layer2_outputs(6579) <= b;
    layer2_outputs(6580) <= not b;
    layer2_outputs(6581) <= not b;
    layer2_outputs(6582) <= not b or a;
    layer2_outputs(6583) <= a;
    layer2_outputs(6584) <= a and not b;
    layer2_outputs(6585) <= a and b;
    layer2_outputs(6586) <= not (a or b);
    layer2_outputs(6587) <= not a or b;
    layer2_outputs(6588) <= a and not b;
    layer2_outputs(6589) <= a;
    layer2_outputs(6590) <= not a;
    layer2_outputs(6591) <= not (a xor b);
    layer2_outputs(6592) <= b and not a;
    layer2_outputs(6593) <= b and not a;
    layer2_outputs(6594) <= a xor b;
    layer2_outputs(6595) <= b;
    layer2_outputs(6596) <= not a or b;
    layer2_outputs(6597) <= a and b;
    layer2_outputs(6598) <= b;
    layer2_outputs(6599) <= a;
    layer2_outputs(6600) <= a or b;
    layer2_outputs(6601) <= a;
    layer2_outputs(6602) <= a xor b;
    layer2_outputs(6603) <= a or b;
    layer2_outputs(6604) <= not b;
    layer2_outputs(6605) <= b and not a;
    layer2_outputs(6606) <= a and not b;
    layer2_outputs(6607) <= a;
    layer2_outputs(6608) <= b;
    layer2_outputs(6609) <= a;
    layer2_outputs(6610) <= not (a xor b);
    layer2_outputs(6611) <= b and not a;
    layer2_outputs(6612) <= a xor b;
    layer2_outputs(6613) <= not a;
    layer2_outputs(6614) <= not b;
    layer2_outputs(6615) <= not a;
    layer2_outputs(6616) <= b;
    layer2_outputs(6617) <= b;
    layer2_outputs(6618) <= not a;
    layer2_outputs(6619) <= not a;
    layer2_outputs(6620) <= not a;
    layer2_outputs(6621) <= a;
    layer2_outputs(6622) <= not (a or b);
    layer2_outputs(6623) <= not (a xor b);
    layer2_outputs(6624) <= b;
    layer2_outputs(6625) <= not (a xor b);
    layer2_outputs(6626) <= not (a xor b);
    layer2_outputs(6627) <= a;
    layer2_outputs(6628) <= not (a xor b);
    layer2_outputs(6629) <= a xor b;
    layer2_outputs(6630) <= a and not b;
    layer2_outputs(6631) <= not a;
    layer2_outputs(6632) <= not (a or b);
    layer2_outputs(6633) <= not b;
    layer2_outputs(6634) <= not b;
    layer2_outputs(6635) <= not a or b;
    layer2_outputs(6636) <= not b;
    layer2_outputs(6637) <= a xor b;
    layer2_outputs(6638) <= not a or b;
    layer2_outputs(6639) <= not (a or b);
    layer2_outputs(6640) <= b and not a;
    layer2_outputs(6641) <= a;
    layer2_outputs(6642) <= not (a xor b);
    layer2_outputs(6643) <= not (a xor b);
    layer2_outputs(6644) <= a;
    layer2_outputs(6645) <= not b;
    layer2_outputs(6646) <= b;
    layer2_outputs(6647) <= a and b;
    layer2_outputs(6648) <= a and not b;
    layer2_outputs(6649) <= not b or a;
    layer2_outputs(6650) <= a and b;
    layer2_outputs(6651) <= not a;
    layer2_outputs(6652) <= a xor b;
    layer2_outputs(6653) <= b;
    layer2_outputs(6654) <= not (a and b);
    layer2_outputs(6655) <= a and b;
    layer2_outputs(6656) <= not b;
    layer2_outputs(6657) <= b;
    layer2_outputs(6658) <= a xor b;
    layer2_outputs(6659) <= '1';
    layer2_outputs(6660) <= a and not b;
    layer2_outputs(6661) <= a;
    layer2_outputs(6662) <= not a or b;
    layer2_outputs(6663) <= a xor b;
    layer2_outputs(6664) <= a xor b;
    layer2_outputs(6665) <= b and not a;
    layer2_outputs(6666) <= b;
    layer2_outputs(6667) <= a or b;
    layer2_outputs(6668) <= b;
    layer2_outputs(6669) <= not b or a;
    layer2_outputs(6670) <= not (a or b);
    layer2_outputs(6671) <= not (a xor b);
    layer2_outputs(6672) <= not b;
    layer2_outputs(6673) <= not (a xor b);
    layer2_outputs(6674) <= not a;
    layer2_outputs(6675) <= a and b;
    layer2_outputs(6676) <= not a;
    layer2_outputs(6677) <= not b;
    layer2_outputs(6678) <= a;
    layer2_outputs(6679) <= not a;
    layer2_outputs(6680) <= not (a or b);
    layer2_outputs(6681) <= not b;
    layer2_outputs(6682) <= not (a and b);
    layer2_outputs(6683) <= a;
    layer2_outputs(6684) <= not a or b;
    layer2_outputs(6685) <= b;
    layer2_outputs(6686) <= a xor b;
    layer2_outputs(6687) <= a;
    layer2_outputs(6688) <= not a;
    layer2_outputs(6689) <= a;
    layer2_outputs(6690) <= a;
    layer2_outputs(6691) <= a;
    layer2_outputs(6692) <= b and not a;
    layer2_outputs(6693) <= not (a xor b);
    layer2_outputs(6694) <= not a;
    layer2_outputs(6695) <= not (a xor b);
    layer2_outputs(6696) <= a xor b;
    layer2_outputs(6697) <= b;
    layer2_outputs(6698) <= a xor b;
    layer2_outputs(6699) <= a xor b;
    layer2_outputs(6700) <= a;
    layer2_outputs(6701) <= b;
    layer2_outputs(6702) <= b;
    layer2_outputs(6703) <= a or b;
    layer2_outputs(6704) <= not (a or b);
    layer2_outputs(6705) <= not a;
    layer2_outputs(6706) <= not (a xor b);
    layer2_outputs(6707) <= not (a or b);
    layer2_outputs(6708) <= a xor b;
    layer2_outputs(6709) <= not b;
    layer2_outputs(6710) <= a;
    layer2_outputs(6711) <= a xor b;
    layer2_outputs(6712) <= not a;
    layer2_outputs(6713) <= not b or a;
    layer2_outputs(6714) <= b;
    layer2_outputs(6715) <= a and not b;
    layer2_outputs(6716) <= a and b;
    layer2_outputs(6717) <= not a or b;
    layer2_outputs(6718) <= a;
    layer2_outputs(6719) <= not a;
    layer2_outputs(6720) <= a and b;
    layer2_outputs(6721) <= not b;
    layer2_outputs(6722) <= not (a and b);
    layer2_outputs(6723) <= a xor b;
    layer2_outputs(6724) <= not b or a;
    layer2_outputs(6725) <= a;
    layer2_outputs(6726) <= a and not b;
    layer2_outputs(6727) <= not b or a;
    layer2_outputs(6728) <= a;
    layer2_outputs(6729) <= not a;
    layer2_outputs(6730) <= not (a xor b);
    layer2_outputs(6731) <= not (a xor b);
    layer2_outputs(6732) <= not (a xor b);
    layer2_outputs(6733) <= a and not b;
    layer2_outputs(6734) <= not b;
    layer2_outputs(6735) <= a xor b;
    layer2_outputs(6736) <= a;
    layer2_outputs(6737) <= a and b;
    layer2_outputs(6738) <= a and b;
    layer2_outputs(6739) <= not a or b;
    layer2_outputs(6740) <= a and not b;
    layer2_outputs(6741) <= not b;
    layer2_outputs(6742) <= a and not b;
    layer2_outputs(6743) <= not (a and b);
    layer2_outputs(6744) <= not b or a;
    layer2_outputs(6745) <= a;
    layer2_outputs(6746) <= a or b;
    layer2_outputs(6747) <= not b;
    layer2_outputs(6748) <= not b;
    layer2_outputs(6749) <= b and not a;
    layer2_outputs(6750) <= a;
    layer2_outputs(6751) <= not a or b;
    layer2_outputs(6752) <= not (a xor b);
    layer2_outputs(6753) <= a or b;
    layer2_outputs(6754) <= a xor b;
    layer2_outputs(6755) <= not b;
    layer2_outputs(6756) <= b;
    layer2_outputs(6757) <= not (a and b);
    layer2_outputs(6758) <= a;
    layer2_outputs(6759) <= b and not a;
    layer2_outputs(6760) <= a and b;
    layer2_outputs(6761) <= not (a xor b);
    layer2_outputs(6762) <= a and not b;
    layer2_outputs(6763) <= a xor b;
    layer2_outputs(6764) <= not b or a;
    layer2_outputs(6765) <= a and b;
    layer2_outputs(6766) <= a;
    layer2_outputs(6767) <= b and not a;
    layer2_outputs(6768) <= not b;
    layer2_outputs(6769) <= not (a xor b);
    layer2_outputs(6770) <= not a;
    layer2_outputs(6771) <= not (a or b);
    layer2_outputs(6772) <= a or b;
    layer2_outputs(6773) <= b;
    layer2_outputs(6774) <= a or b;
    layer2_outputs(6775) <= not a;
    layer2_outputs(6776) <= a and b;
    layer2_outputs(6777) <= a;
    layer2_outputs(6778) <= not b;
    layer2_outputs(6779) <= not (a or b);
    layer2_outputs(6780) <= not b;
    layer2_outputs(6781) <= a;
    layer2_outputs(6782) <= a and b;
    layer2_outputs(6783) <= a;
    layer2_outputs(6784) <= not (a or b);
    layer2_outputs(6785) <= not a;
    layer2_outputs(6786) <= a and b;
    layer2_outputs(6787) <= not b;
    layer2_outputs(6788) <= not (a xor b);
    layer2_outputs(6789) <= a xor b;
    layer2_outputs(6790) <= b;
    layer2_outputs(6791) <= not a;
    layer2_outputs(6792) <= a;
    layer2_outputs(6793) <= a and b;
    layer2_outputs(6794) <= not b;
    layer2_outputs(6795) <= b;
    layer2_outputs(6796) <= not a;
    layer2_outputs(6797) <= a and b;
    layer2_outputs(6798) <= not (a xor b);
    layer2_outputs(6799) <= a xor b;
    layer2_outputs(6800) <= not b or a;
    layer2_outputs(6801) <= b;
    layer2_outputs(6802) <= b and not a;
    layer2_outputs(6803) <= not a;
    layer2_outputs(6804) <= '1';
    layer2_outputs(6805) <= not a;
    layer2_outputs(6806) <= b;
    layer2_outputs(6807) <= not (a xor b);
    layer2_outputs(6808) <= not a;
    layer2_outputs(6809) <= a or b;
    layer2_outputs(6810) <= b;
    layer2_outputs(6811) <= not b;
    layer2_outputs(6812) <= a or b;
    layer2_outputs(6813) <= a;
    layer2_outputs(6814) <= not b or a;
    layer2_outputs(6815) <= not b;
    layer2_outputs(6816) <= not a;
    layer2_outputs(6817) <= b;
    layer2_outputs(6818) <= a;
    layer2_outputs(6819) <= a;
    layer2_outputs(6820) <= not (a and b);
    layer2_outputs(6821) <= a and not b;
    layer2_outputs(6822) <= not a or b;
    layer2_outputs(6823) <= b;
    layer2_outputs(6824) <= a and b;
    layer2_outputs(6825) <= not a or b;
    layer2_outputs(6826) <= not a or b;
    layer2_outputs(6827) <= not b;
    layer2_outputs(6828) <= b;
    layer2_outputs(6829) <= '0';
    layer2_outputs(6830) <= b;
    layer2_outputs(6831) <= not (a or b);
    layer2_outputs(6832) <= not b;
    layer2_outputs(6833) <= not a;
    layer2_outputs(6834) <= a xor b;
    layer2_outputs(6835) <= a;
    layer2_outputs(6836) <= not b;
    layer2_outputs(6837) <= not b;
    layer2_outputs(6838) <= a;
    layer2_outputs(6839) <= a;
    layer2_outputs(6840) <= not a;
    layer2_outputs(6841) <= b;
    layer2_outputs(6842) <= not b;
    layer2_outputs(6843) <= not (a and b);
    layer2_outputs(6844) <= b;
    layer2_outputs(6845) <= a;
    layer2_outputs(6846) <= a and b;
    layer2_outputs(6847) <= not a;
    layer2_outputs(6848) <= not a or b;
    layer2_outputs(6849) <= b and not a;
    layer2_outputs(6850) <= not (a and b);
    layer2_outputs(6851) <= not b;
    layer2_outputs(6852) <= b and not a;
    layer2_outputs(6853) <= a;
    layer2_outputs(6854) <= '0';
    layer2_outputs(6855) <= a xor b;
    layer2_outputs(6856) <= not (a or b);
    layer2_outputs(6857) <= b;
    layer2_outputs(6858) <= b;
    layer2_outputs(6859) <= a or b;
    layer2_outputs(6860) <= not a or b;
    layer2_outputs(6861) <= not a;
    layer2_outputs(6862) <= not (a or b);
    layer2_outputs(6863) <= b;
    layer2_outputs(6864) <= not b;
    layer2_outputs(6865) <= not (a xor b);
    layer2_outputs(6866) <= b and not a;
    layer2_outputs(6867) <= a and b;
    layer2_outputs(6868) <= a;
    layer2_outputs(6869) <= a or b;
    layer2_outputs(6870) <= a and not b;
    layer2_outputs(6871) <= not a;
    layer2_outputs(6872) <= a and not b;
    layer2_outputs(6873) <= a xor b;
    layer2_outputs(6874) <= not a or b;
    layer2_outputs(6875) <= a;
    layer2_outputs(6876) <= a and b;
    layer2_outputs(6877) <= b and not a;
    layer2_outputs(6878) <= not (a xor b);
    layer2_outputs(6879) <= not (a xor b);
    layer2_outputs(6880) <= a or b;
    layer2_outputs(6881) <= a and not b;
    layer2_outputs(6882) <= '1';
    layer2_outputs(6883) <= not (a and b);
    layer2_outputs(6884) <= not (a or b);
    layer2_outputs(6885) <= not b or a;
    layer2_outputs(6886) <= a and b;
    layer2_outputs(6887) <= not a;
    layer2_outputs(6888) <= b;
    layer2_outputs(6889) <= not b or a;
    layer2_outputs(6890) <= a and not b;
    layer2_outputs(6891) <= not (a and b);
    layer2_outputs(6892) <= not a or b;
    layer2_outputs(6893) <= not (a xor b);
    layer2_outputs(6894) <= not (a and b);
    layer2_outputs(6895) <= b and not a;
    layer2_outputs(6896) <= a xor b;
    layer2_outputs(6897) <= not b or a;
    layer2_outputs(6898) <= a or b;
    layer2_outputs(6899) <= b;
    layer2_outputs(6900) <= a and b;
    layer2_outputs(6901) <= a and b;
    layer2_outputs(6902) <= not (a xor b);
    layer2_outputs(6903) <= a xor b;
    layer2_outputs(6904) <= a;
    layer2_outputs(6905) <= b;
    layer2_outputs(6906) <= not b;
    layer2_outputs(6907) <= a xor b;
    layer2_outputs(6908) <= not b;
    layer2_outputs(6909) <= not b;
    layer2_outputs(6910) <= not (a or b);
    layer2_outputs(6911) <= not a;
    layer2_outputs(6912) <= a xor b;
    layer2_outputs(6913) <= not a or b;
    layer2_outputs(6914) <= a xor b;
    layer2_outputs(6915) <= a and b;
    layer2_outputs(6916) <= a;
    layer2_outputs(6917) <= a xor b;
    layer2_outputs(6918) <= not a or b;
    layer2_outputs(6919) <= a and b;
    layer2_outputs(6920) <= not a;
    layer2_outputs(6921) <= not (a or b);
    layer2_outputs(6922) <= b;
    layer2_outputs(6923) <= a and not b;
    layer2_outputs(6924) <= not b or a;
    layer2_outputs(6925) <= not a or b;
    layer2_outputs(6926) <= a and not b;
    layer2_outputs(6927) <= not (a and b);
    layer2_outputs(6928) <= a xor b;
    layer2_outputs(6929) <= a xor b;
    layer2_outputs(6930) <= a or b;
    layer2_outputs(6931) <= not a;
    layer2_outputs(6932) <= a and b;
    layer2_outputs(6933) <= a;
    layer2_outputs(6934) <= a xor b;
    layer2_outputs(6935) <= a and not b;
    layer2_outputs(6936) <= b;
    layer2_outputs(6937) <= a and b;
    layer2_outputs(6938) <= not (a xor b);
    layer2_outputs(6939) <= not b;
    layer2_outputs(6940) <= a and b;
    layer2_outputs(6941) <= a xor b;
    layer2_outputs(6942) <= a and not b;
    layer2_outputs(6943) <= not b;
    layer2_outputs(6944) <= a or b;
    layer2_outputs(6945) <= a and b;
    layer2_outputs(6946) <= b;
    layer2_outputs(6947) <= not b;
    layer2_outputs(6948) <= b and not a;
    layer2_outputs(6949) <= not b or a;
    layer2_outputs(6950) <= b;
    layer2_outputs(6951) <= not b;
    layer2_outputs(6952) <= a;
    layer2_outputs(6953) <= a;
    layer2_outputs(6954) <= b;
    layer2_outputs(6955) <= not (a or b);
    layer2_outputs(6956) <= not b;
    layer2_outputs(6957) <= not a;
    layer2_outputs(6958) <= not b or a;
    layer2_outputs(6959) <= not a;
    layer2_outputs(6960) <= a and b;
    layer2_outputs(6961) <= a xor b;
    layer2_outputs(6962) <= a and not b;
    layer2_outputs(6963) <= a and not b;
    layer2_outputs(6964) <= not b or a;
    layer2_outputs(6965) <= a;
    layer2_outputs(6966) <= b;
    layer2_outputs(6967) <= a;
    layer2_outputs(6968) <= a and not b;
    layer2_outputs(6969) <= a and b;
    layer2_outputs(6970) <= not a or b;
    layer2_outputs(6971) <= not a;
    layer2_outputs(6972) <= a;
    layer2_outputs(6973) <= not (a and b);
    layer2_outputs(6974) <= not b or a;
    layer2_outputs(6975) <= not b;
    layer2_outputs(6976) <= b;
    layer2_outputs(6977) <= a and not b;
    layer2_outputs(6978) <= not a;
    layer2_outputs(6979) <= not b;
    layer2_outputs(6980) <= not b;
    layer2_outputs(6981) <= b;
    layer2_outputs(6982) <= b;
    layer2_outputs(6983) <= a xor b;
    layer2_outputs(6984) <= a xor b;
    layer2_outputs(6985) <= a xor b;
    layer2_outputs(6986) <= a and not b;
    layer2_outputs(6987) <= a or b;
    layer2_outputs(6988) <= not b;
    layer2_outputs(6989) <= b;
    layer2_outputs(6990) <= not a or b;
    layer2_outputs(6991) <= a xor b;
    layer2_outputs(6992) <= a and not b;
    layer2_outputs(6993) <= a or b;
    layer2_outputs(6994) <= a and b;
    layer2_outputs(6995) <= '1';
    layer2_outputs(6996) <= a xor b;
    layer2_outputs(6997) <= not (a and b);
    layer2_outputs(6998) <= b;
    layer2_outputs(6999) <= a and b;
    layer2_outputs(7000) <= not (a xor b);
    layer2_outputs(7001) <= a or b;
    layer2_outputs(7002) <= not a or b;
    layer2_outputs(7003) <= a xor b;
    layer2_outputs(7004) <= not (a and b);
    layer2_outputs(7005) <= not b;
    layer2_outputs(7006) <= b and not a;
    layer2_outputs(7007) <= b;
    layer2_outputs(7008) <= not a;
    layer2_outputs(7009) <= not (a or b);
    layer2_outputs(7010) <= a and b;
    layer2_outputs(7011) <= a xor b;
    layer2_outputs(7012) <= b and not a;
    layer2_outputs(7013) <= not (a xor b);
    layer2_outputs(7014) <= a and not b;
    layer2_outputs(7015) <= not (a xor b);
    layer2_outputs(7016) <= a and not b;
    layer2_outputs(7017) <= not a;
    layer2_outputs(7018) <= a;
    layer2_outputs(7019) <= b;
    layer2_outputs(7020) <= not a;
    layer2_outputs(7021) <= a xor b;
    layer2_outputs(7022) <= not (a or b);
    layer2_outputs(7023) <= not b or a;
    layer2_outputs(7024) <= a;
    layer2_outputs(7025) <= not a;
    layer2_outputs(7026) <= a xor b;
    layer2_outputs(7027) <= b;
    layer2_outputs(7028) <= a xor b;
    layer2_outputs(7029) <= not (a xor b);
    layer2_outputs(7030) <= a or b;
    layer2_outputs(7031) <= not (a or b);
    layer2_outputs(7032) <= a and not b;
    layer2_outputs(7033) <= not (a or b);
    layer2_outputs(7034) <= not b;
    layer2_outputs(7035) <= a xor b;
    layer2_outputs(7036) <= not (a and b);
    layer2_outputs(7037) <= not (a or b);
    layer2_outputs(7038) <= not a;
    layer2_outputs(7039) <= not b;
    layer2_outputs(7040) <= not a;
    layer2_outputs(7041) <= a xor b;
    layer2_outputs(7042) <= a;
    layer2_outputs(7043) <= not b or a;
    layer2_outputs(7044) <= not (a xor b);
    layer2_outputs(7045) <= not (a and b);
    layer2_outputs(7046) <= not (a or b);
    layer2_outputs(7047) <= a and b;
    layer2_outputs(7048) <= a and not b;
    layer2_outputs(7049) <= b;
    layer2_outputs(7050) <= a;
    layer2_outputs(7051) <= not (a or b);
    layer2_outputs(7052) <= a or b;
    layer2_outputs(7053) <= a and not b;
    layer2_outputs(7054) <= not b;
    layer2_outputs(7055) <= a xor b;
    layer2_outputs(7056) <= not (a xor b);
    layer2_outputs(7057) <= a;
    layer2_outputs(7058) <= not (a or b);
    layer2_outputs(7059) <= b;
    layer2_outputs(7060) <= a xor b;
    layer2_outputs(7061) <= a xor b;
    layer2_outputs(7062) <= not (a xor b);
    layer2_outputs(7063) <= b;
    layer2_outputs(7064) <= not b or a;
    layer2_outputs(7065) <= not (a or b);
    layer2_outputs(7066) <= a and not b;
    layer2_outputs(7067) <= a;
    layer2_outputs(7068) <= not b;
    layer2_outputs(7069) <= a;
    layer2_outputs(7070) <= not b or a;
    layer2_outputs(7071) <= not (a and b);
    layer2_outputs(7072) <= a and not b;
    layer2_outputs(7073) <= not b or a;
    layer2_outputs(7074) <= not a or b;
    layer2_outputs(7075) <= a and not b;
    layer2_outputs(7076) <= a;
    layer2_outputs(7077) <= a;
    layer2_outputs(7078) <= a;
    layer2_outputs(7079) <= not a;
    layer2_outputs(7080) <= a and not b;
    layer2_outputs(7081) <= not b;
    layer2_outputs(7082) <= not (a xor b);
    layer2_outputs(7083) <= not (a xor b);
    layer2_outputs(7084) <= b;
    layer2_outputs(7085) <= b and not a;
    layer2_outputs(7086) <= not b or a;
    layer2_outputs(7087) <= not a or b;
    layer2_outputs(7088) <= b;
    layer2_outputs(7089) <= not b;
    layer2_outputs(7090) <= not a;
    layer2_outputs(7091) <= not (a or b);
    layer2_outputs(7092) <= a xor b;
    layer2_outputs(7093) <= not (a and b);
    layer2_outputs(7094) <= not (a or b);
    layer2_outputs(7095) <= not a;
    layer2_outputs(7096) <= b;
    layer2_outputs(7097) <= b and not a;
    layer2_outputs(7098) <= not b;
    layer2_outputs(7099) <= not a;
    layer2_outputs(7100) <= a and b;
    layer2_outputs(7101) <= not (a and b);
    layer2_outputs(7102) <= not b;
    layer2_outputs(7103) <= not b;
    layer2_outputs(7104) <= b;
    layer2_outputs(7105) <= not b or a;
    layer2_outputs(7106) <= a or b;
    layer2_outputs(7107) <= not a or b;
    layer2_outputs(7108) <= b;
    layer2_outputs(7109) <= not b or a;
    layer2_outputs(7110) <= not (a and b);
    layer2_outputs(7111) <= not (a and b);
    layer2_outputs(7112) <= not b;
    layer2_outputs(7113) <= not (a xor b);
    layer2_outputs(7114) <= b;
    layer2_outputs(7115) <= a xor b;
    layer2_outputs(7116) <= not (a or b);
    layer2_outputs(7117) <= not a;
    layer2_outputs(7118) <= a and b;
    layer2_outputs(7119) <= a and not b;
    layer2_outputs(7120) <= not b or a;
    layer2_outputs(7121) <= not a;
    layer2_outputs(7122) <= a and b;
    layer2_outputs(7123) <= a and b;
    layer2_outputs(7124) <= a or b;
    layer2_outputs(7125) <= a or b;
    layer2_outputs(7126) <= a xor b;
    layer2_outputs(7127) <= a and b;
    layer2_outputs(7128) <= not a;
    layer2_outputs(7129) <= not (a or b);
    layer2_outputs(7130) <= not (a and b);
    layer2_outputs(7131) <= b;
    layer2_outputs(7132) <= a and not b;
    layer2_outputs(7133) <= a;
    layer2_outputs(7134) <= not b or a;
    layer2_outputs(7135) <= a;
    layer2_outputs(7136) <= not a;
    layer2_outputs(7137) <= b;
    layer2_outputs(7138) <= not b;
    layer2_outputs(7139) <= not (a or b);
    layer2_outputs(7140) <= a xor b;
    layer2_outputs(7141) <= b;
    layer2_outputs(7142) <= not (a xor b);
    layer2_outputs(7143) <= not (a or b);
    layer2_outputs(7144) <= not a;
    layer2_outputs(7145) <= not (a or b);
    layer2_outputs(7146) <= not (a xor b);
    layer2_outputs(7147) <= not b;
    layer2_outputs(7148) <= not (a and b);
    layer2_outputs(7149) <= b;
    layer2_outputs(7150) <= a xor b;
    layer2_outputs(7151) <= not (a and b);
    layer2_outputs(7152) <= not (a and b);
    layer2_outputs(7153) <= not b;
    layer2_outputs(7154) <= a;
    layer2_outputs(7155) <= b;
    layer2_outputs(7156) <= b;
    layer2_outputs(7157) <= not b or a;
    layer2_outputs(7158) <= not (a xor b);
    layer2_outputs(7159) <= '0';
    layer2_outputs(7160) <= not (a and b);
    layer2_outputs(7161) <= b and not a;
    layer2_outputs(7162) <= not (a or b);
    layer2_outputs(7163) <= not a;
    layer2_outputs(7164) <= a;
    layer2_outputs(7165) <= a or b;
    layer2_outputs(7166) <= a;
    layer2_outputs(7167) <= not b or a;
    layer2_outputs(7168) <= not b;
    layer2_outputs(7169) <= not b;
    layer2_outputs(7170) <= b;
    layer2_outputs(7171) <= not a;
    layer2_outputs(7172) <= b;
    layer2_outputs(7173) <= not (a or b);
    layer2_outputs(7174) <= b;
    layer2_outputs(7175) <= not (a xor b);
    layer2_outputs(7176) <= not (a or b);
    layer2_outputs(7177) <= b and not a;
    layer2_outputs(7178) <= a or b;
    layer2_outputs(7179) <= a;
    layer2_outputs(7180) <= not (a xor b);
    layer2_outputs(7181) <= not (a xor b);
    layer2_outputs(7182) <= not b;
    layer2_outputs(7183) <= b and not a;
    layer2_outputs(7184) <= not b;
    layer2_outputs(7185) <= b;
    layer2_outputs(7186) <= not (a and b);
    layer2_outputs(7187) <= a;
    layer2_outputs(7188) <= a;
    layer2_outputs(7189) <= not a;
    layer2_outputs(7190) <= b;
    layer2_outputs(7191) <= a and not b;
    layer2_outputs(7192) <= b and not a;
    layer2_outputs(7193) <= not a;
    layer2_outputs(7194) <= b;
    layer2_outputs(7195) <= b and not a;
    layer2_outputs(7196) <= not b or a;
    layer2_outputs(7197) <= not b;
    layer2_outputs(7198) <= not b;
    layer2_outputs(7199) <= a or b;
    layer2_outputs(7200) <= a and b;
    layer2_outputs(7201) <= a or b;
    layer2_outputs(7202) <= not a;
    layer2_outputs(7203) <= not b;
    layer2_outputs(7204) <= a;
    layer2_outputs(7205) <= not a;
    layer2_outputs(7206) <= not b;
    layer2_outputs(7207) <= not b;
    layer2_outputs(7208) <= not (a and b);
    layer2_outputs(7209) <= b;
    layer2_outputs(7210) <= a;
    layer2_outputs(7211) <= a or b;
    layer2_outputs(7212) <= not b or a;
    layer2_outputs(7213) <= not b;
    layer2_outputs(7214) <= a and not b;
    layer2_outputs(7215) <= not b or a;
    layer2_outputs(7216) <= not (a and b);
    layer2_outputs(7217) <= not a;
    layer2_outputs(7218) <= not b or a;
    layer2_outputs(7219) <= a xor b;
    layer2_outputs(7220) <= b;
    layer2_outputs(7221) <= not (a or b);
    layer2_outputs(7222) <= not b or a;
    layer2_outputs(7223) <= not a;
    layer2_outputs(7224) <= a and not b;
    layer2_outputs(7225) <= not (a or b);
    layer2_outputs(7226) <= a;
    layer2_outputs(7227) <= not (a xor b);
    layer2_outputs(7228) <= not (a or b);
    layer2_outputs(7229) <= a and not b;
    layer2_outputs(7230) <= a and b;
    layer2_outputs(7231) <= not (a xor b);
    layer2_outputs(7232) <= not a or b;
    layer2_outputs(7233) <= not a;
    layer2_outputs(7234) <= a and not b;
    layer2_outputs(7235) <= not a or b;
    layer2_outputs(7236) <= not a or b;
    layer2_outputs(7237) <= a or b;
    layer2_outputs(7238) <= not a or b;
    layer2_outputs(7239) <= b;
    layer2_outputs(7240) <= a xor b;
    layer2_outputs(7241) <= not a;
    layer2_outputs(7242) <= '1';
    layer2_outputs(7243) <= a;
    layer2_outputs(7244) <= not a;
    layer2_outputs(7245) <= not (a and b);
    layer2_outputs(7246) <= a or b;
    layer2_outputs(7247) <= not b or a;
    layer2_outputs(7248) <= b and not a;
    layer2_outputs(7249) <= b and not a;
    layer2_outputs(7250) <= not b or a;
    layer2_outputs(7251) <= not a;
    layer2_outputs(7252) <= not a;
    layer2_outputs(7253) <= b;
    layer2_outputs(7254) <= not (a and b);
    layer2_outputs(7255) <= not a;
    layer2_outputs(7256) <= a and b;
    layer2_outputs(7257) <= a and b;
    layer2_outputs(7258) <= not b or a;
    layer2_outputs(7259) <= a and b;
    layer2_outputs(7260) <= not b;
    layer2_outputs(7261) <= a and not b;
    layer2_outputs(7262) <= not (a or b);
    layer2_outputs(7263) <= not a;
    layer2_outputs(7264) <= a or b;
    layer2_outputs(7265) <= not (a and b);
    layer2_outputs(7266) <= a and b;
    layer2_outputs(7267) <= a or b;
    layer2_outputs(7268) <= not (a xor b);
    layer2_outputs(7269) <= '0';
    layer2_outputs(7270) <= b;
    layer2_outputs(7271) <= b and not a;
    layer2_outputs(7272) <= not a;
    layer2_outputs(7273) <= a and not b;
    layer2_outputs(7274) <= not b;
    layer2_outputs(7275) <= not (a or b);
    layer2_outputs(7276) <= not a;
    layer2_outputs(7277) <= b;
    layer2_outputs(7278) <= a;
    layer2_outputs(7279) <= not a;
    layer2_outputs(7280) <= b;
    layer2_outputs(7281) <= not a or b;
    layer2_outputs(7282) <= b and not a;
    layer2_outputs(7283) <= a xor b;
    layer2_outputs(7284) <= a;
    layer2_outputs(7285) <= a or b;
    layer2_outputs(7286) <= not (a or b);
    layer2_outputs(7287) <= not (a and b);
    layer2_outputs(7288) <= not a;
    layer2_outputs(7289) <= not (a and b);
    layer2_outputs(7290) <= b;
    layer2_outputs(7291) <= not b or a;
    layer2_outputs(7292) <= a and not b;
    layer2_outputs(7293) <= not (a xor b);
    layer2_outputs(7294) <= a and not b;
    layer2_outputs(7295) <= a and b;
    layer2_outputs(7296) <= a xor b;
    layer2_outputs(7297) <= a or b;
    layer2_outputs(7298) <= not a;
    layer2_outputs(7299) <= a and not b;
    layer2_outputs(7300) <= a;
    layer2_outputs(7301) <= a;
    layer2_outputs(7302) <= b and not a;
    layer2_outputs(7303) <= a;
    layer2_outputs(7304) <= not (a or b);
    layer2_outputs(7305) <= a or b;
    layer2_outputs(7306) <= not a;
    layer2_outputs(7307) <= not b or a;
    layer2_outputs(7308) <= not b;
    layer2_outputs(7309) <= not a or b;
    layer2_outputs(7310) <= b;
    layer2_outputs(7311) <= not (a xor b);
    layer2_outputs(7312) <= a;
    layer2_outputs(7313) <= a;
    layer2_outputs(7314) <= a and b;
    layer2_outputs(7315) <= a;
    layer2_outputs(7316) <= not (a or b);
    layer2_outputs(7317) <= not b or a;
    layer2_outputs(7318) <= a;
    layer2_outputs(7319) <= a;
    layer2_outputs(7320) <= b and not a;
    layer2_outputs(7321) <= not (a and b);
    layer2_outputs(7322) <= b and not a;
    layer2_outputs(7323) <= not (a and b);
    layer2_outputs(7324) <= a and not b;
    layer2_outputs(7325) <= not a;
    layer2_outputs(7326) <= not (a and b);
    layer2_outputs(7327) <= a xor b;
    layer2_outputs(7328) <= a;
    layer2_outputs(7329) <= not a or b;
    layer2_outputs(7330) <= a or b;
    layer2_outputs(7331) <= not a or b;
    layer2_outputs(7332) <= not (a xor b);
    layer2_outputs(7333) <= a or b;
    layer2_outputs(7334) <= not b;
    layer2_outputs(7335) <= '0';
    layer2_outputs(7336) <= not a or b;
    layer2_outputs(7337) <= not a or b;
    layer2_outputs(7338) <= a xor b;
    layer2_outputs(7339) <= not b;
    layer2_outputs(7340) <= a;
    layer2_outputs(7341) <= b and not a;
    layer2_outputs(7342) <= not a;
    layer2_outputs(7343) <= not (a or b);
    layer2_outputs(7344) <= a;
    layer2_outputs(7345) <= not (a or b);
    layer2_outputs(7346) <= not b;
    layer2_outputs(7347) <= not (a xor b);
    layer2_outputs(7348) <= not b;
    layer2_outputs(7349) <= not b;
    layer2_outputs(7350) <= not a or b;
    layer2_outputs(7351) <= not b or a;
    layer2_outputs(7352) <= a;
    layer2_outputs(7353) <= a;
    layer2_outputs(7354) <= a;
    layer2_outputs(7355) <= not b or a;
    layer2_outputs(7356) <= b;
    layer2_outputs(7357) <= a xor b;
    layer2_outputs(7358) <= '1';
    layer2_outputs(7359) <= not b;
    layer2_outputs(7360) <= a xor b;
    layer2_outputs(7361) <= not a;
    layer2_outputs(7362) <= not a;
    layer2_outputs(7363) <= not b;
    layer2_outputs(7364) <= not a or b;
    layer2_outputs(7365) <= not a;
    layer2_outputs(7366) <= not a;
    layer2_outputs(7367) <= not b or a;
    layer2_outputs(7368) <= b;
    layer2_outputs(7369) <= b;
    layer2_outputs(7370) <= b and not a;
    layer2_outputs(7371) <= not a;
    layer2_outputs(7372) <= not b or a;
    layer2_outputs(7373) <= a and b;
    layer2_outputs(7374) <= a xor b;
    layer2_outputs(7375) <= b and not a;
    layer2_outputs(7376) <= a and not b;
    layer2_outputs(7377) <= not a or b;
    layer2_outputs(7378) <= b;
    layer2_outputs(7379) <= b and not a;
    layer2_outputs(7380) <= a and not b;
    layer2_outputs(7381) <= a xor b;
    layer2_outputs(7382) <= a;
    layer2_outputs(7383) <= a and not b;
    layer2_outputs(7384) <= not (a or b);
    layer2_outputs(7385) <= a;
    layer2_outputs(7386) <= b;
    layer2_outputs(7387) <= not (a and b);
    layer2_outputs(7388) <= b and not a;
    layer2_outputs(7389) <= a xor b;
    layer2_outputs(7390) <= not b;
    layer2_outputs(7391) <= not a;
    layer2_outputs(7392) <= not (a xor b);
    layer2_outputs(7393) <= b;
    layer2_outputs(7394) <= not a or b;
    layer2_outputs(7395) <= not b;
    layer2_outputs(7396) <= not (a xor b);
    layer2_outputs(7397) <= not a;
    layer2_outputs(7398) <= a xor b;
    layer2_outputs(7399) <= a and b;
    layer2_outputs(7400) <= not a or b;
    layer2_outputs(7401) <= not a or b;
    layer2_outputs(7402) <= not a or b;
    layer2_outputs(7403) <= not b;
    layer2_outputs(7404) <= not (a and b);
    layer2_outputs(7405) <= a;
    layer2_outputs(7406) <= a xor b;
    layer2_outputs(7407) <= not b;
    layer2_outputs(7408) <= a or b;
    layer2_outputs(7409) <= not (a xor b);
    layer2_outputs(7410) <= not (a xor b);
    layer2_outputs(7411) <= not (a xor b);
    layer2_outputs(7412) <= b;
    layer2_outputs(7413) <= not (a and b);
    layer2_outputs(7414) <= not b;
    layer2_outputs(7415) <= not (a or b);
    layer2_outputs(7416) <= not (a and b);
    layer2_outputs(7417) <= not (a xor b);
    layer2_outputs(7418) <= a or b;
    layer2_outputs(7419) <= a;
    layer2_outputs(7420) <= a and not b;
    layer2_outputs(7421) <= not b or a;
    layer2_outputs(7422) <= '1';
    layer2_outputs(7423) <= a or b;
    layer2_outputs(7424) <= not (a xor b);
    layer2_outputs(7425) <= not a;
    layer2_outputs(7426) <= b and not a;
    layer2_outputs(7427) <= not a;
    layer2_outputs(7428) <= not (a xor b);
    layer2_outputs(7429) <= not (a xor b);
    layer2_outputs(7430) <= not a;
    layer2_outputs(7431) <= a;
    layer2_outputs(7432) <= not (a or b);
    layer2_outputs(7433) <= a xor b;
    layer2_outputs(7434) <= a xor b;
    layer2_outputs(7435) <= a xor b;
    layer2_outputs(7436) <= a;
    layer2_outputs(7437) <= not b;
    layer2_outputs(7438) <= b;
    layer2_outputs(7439) <= not (a or b);
    layer2_outputs(7440) <= a xor b;
    layer2_outputs(7441) <= b and not a;
    layer2_outputs(7442) <= not (a and b);
    layer2_outputs(7443) <= not b;
    layer2_outputs(7444) <= a xor b;
    layer2_outputs(7445) <= a and not b;
    layer2_outputs(7446) <= not a;
    layer2_outputs(7447) <= not a or b;
    layer2_outputs(7448) <= not a or b;
    layer2_outputs(7449) <= not b;
    layer2_outputs(7450) <= not b;
    layer2_outputs(7451) <= b;
    layer2_outputs(7452) <= a and b;
    layer2_outputs(7453) <= not b;
    layer2_outputs(7454) <= a xor b;
    layer2_outputs(7455) <= not (a or b);
    layer2_outputs(7456) <= not b;
    layer2_outputs(7457) <= a xor b;
    layer2_outputs(7458) <= not (a and b);
    layer2_outputs(7459) <= b;
    layer2_outputs(7460) <= not b or a;
    layer2_outputs(7461) <= not (a xor b);
    layer2_outputs(7462) <= a;
    layer2_outputs(7463) <= a xor b;
    layer2_outputs(7464) <= not a;
    layer2_outputs(7465) <= not a or b;
    layer2_outputs(7466) <= b and not a;
    layer2_outputs(7467) <= not a or b;
    layer2_outputs(7468) <= a;
    layer2_outputs(7469) <= not b;
    layer2_outputs(7470) <= not a;
    layer2_outputs(7471) <= not (a and b);
    layer2_outputs(7472) <= not a or b;
    layer2_outputs(7473) <= not b;
    layer2_outputs(7474) <= not a or b;
    layer2_outputs(7475) <= not (a and b);
    layer2_outputs(7476) <= a or b;
    layer2_outputs(7477) <= b;
    layer2_outputs(7478) <= a;
    layer2_outputs(7479) <= a;
    layer2_outputs(7480) <= a;
    layer2_outputs(7481) <= not a;
    layer2_outputs(7482) <= not b or a;
    layer2_outputs(7483) <= not (a and b);
    layer2_outputs(7484) <= a xor b;
    layer2_outputs(7485) <= a and not b;
    layer2_outputs(7486) <= a xor b;
    layer2_outputs(7487) <= not a;
    layer2_outputs(7488) <= not a or b;
    layer2_outputs(7489) <= a and not b;
    layer2_outputs(7490) <= not (a and b);
    layer2_outputs(7491) <= not a;
    layer2_outputs(7492) <= b and not a;
    layer2_outputs(7493) <= not a;
    layer2_outputs(7494) <= not b or a;
    layer2_outputs(7495) <= a and not b;
    layer2_outputs(7496) <= not a;
    layer2_outputs(7497) <= not a or b;
    layer2_outputs(7498) <= not (a xor b);
    layer2_outputs(7499) <= a xor b;
    layer2_outputs(7500) <= not (a and b);
    layer2_outputs(7501) <= not (a xor b);
    layer2_outputs(7502) <= a xor b;
    layer2_outputs(7503) <= a;
    layer2_outputs(7504) <= not b;
    layer2_outputs(7505) <= a and b;
    layer2_outputs(7506) <= b;
    layer2_outputs(7507) <= a;
    layer2_outputs(7508) <= not b;
    layer2_outputs(7509) <= not (a or b);
    layer2_outputs(7510) <= a and not b;
    layer2_outputs(7511) <= a and b;
    layer2_outputs(7512) <= a xor b;
    layer2_outputs(7513) <= not a;
    layer2_outputs(7514) <= not a or b;
    layer2_outputs(7515) <= not (a xor b);
    layer2_outputs(7516) <= a xor b;
    layer2_outputs(7517) <= a xor b;
    layer2_outputs(7518) <= not a;
    layer2_outputs(7519) <= not a;
    layer2_outputs(7520) <= not a or b;
    layer2_outputs(7521) <= a;
    layer2_outputs(7522) <= not b;
    layer2_outputs(7523) <= b;
    layer2_outputs(7524) <= not (a or b);
    layer2_outputs(7525) <= b;
    layer2_outputs(7526) <= b and not a;
    layer2_outputs(7527) <= a;
    layer2_outputs(7528) <= a and not b;
    layer2_outputs(7529) <= not (a and b);
    layer2_outputs(7530) <= not a;
    layer2_outputs(7531) <= not (a xor b);
    layer2_outputs(7532) <= not (a xor b);
    layer2_outputs(7533) <= not (a xor b);
    layer2_outputs(7534) <= b and not a;
    layer2_outputs(7535) <= not a or b;
    layer2_outputs(7536) <= b;
    layer2_outputs(7537) <= not (a or b);
    layer2_outputs(7538) <= not (a xor b);
    layer2_outputs(7539) <= b;
    layer2_outputs(7540) <= not (a or b);
    layer2_outputs(7541) <= not b;
    layer2_outputs(7542) <= not a;
    layer2_outputs(7543) <= a;
    layer2_outputs(7544) <= b;
    layer2_outputs(7545) <= not b or a;
    layer2_outputs(7546) <= not a;
    layer2_outputs(7547) <= not b;
    layer2_outputs(7548) <= a or b;
    layer2_outputs(7549) <= not (a xor b);
    layer2_outputs(7550) <= not (a or b);
    layer2_outputs(7551) <= a and not b;
    layer2_outputs(7552) <= not b;
    layer2_outputs(7553) <= a or b;
    layer2_outputs(7554) <= b;
    layer2_outputs(7555) <= not (a xor b);
    layer2_outputs(7556) <= a and not b;
    layer2_outputs(7557) <= not (a xor b);
    layer2_outputs(7558) <= not a;
    layer2_outputs(7559) <= not b;
    layer2_outputs(7560) <= not (a or b);
    layer2_outputs(7561) <= not b;
    layer2_outputs(7562) <= b;
    layer2_outputs(7563) <= not b;
    layer2_outputs(7564) <= not a or b;
    layer2_outputs(7565) <= not a or b;
    layer2_outputs(7566) <= not a;
    layer2_outputs(7567) <= not b;
    layer2_outputs(7568) <= not b;
    layer2_outputs(7569) <= not a;
    layer2_outputs(7570) <= b;
    layer2_outputs(7571) <= a and not b;
    layer2_outputs(7572) <= a xor b;
    layer2_outputs(7573) <= not (a xor b);
    layer2_outputs(7574) <= b;
    layer2_outputs(7575) <= b;
    layer2_outputs(7576) <= a xor b;
    layer2_outputs(7577) <= b and not a;
    layer2_outputs(7578) <= not (a xor b);
    layer2_outputs(7579) <= not (a xor b);
    layer2_outputs(7580) <= not (a xor b);
    layer2_outputs(7581) <= not b or a;
    layer2_outputs(7582) <= a and not b;
    layer2_outputs(7583) <= a xor b;
    layer2_outputs(7584) <= b and not a;
    layer2_outputs(7585) <= not b;
    layer2_outputs(7586) <= not (a and b);
    layer2_outputs(7587) <= not (a xor b);
    layer2_outputs(7588) <= b;
    layer2_outputs(7589) <= b;
    layer2_outputs(7590) <= b;
    layer2_outputs(7591) <= not (a xor b);
    layer2_outputs(7592) <= a or b;
    layer2_outputs(7593) <= a and not b;
    layer2_outputs(7594) <= not (a xor b);
    layer2_outputs(7595) <= b and not a;
    layer2_outputs(7596) <= not a;
    layer2_outputs(7597) <= a;
    layer2_outputs(7598) <= a and b;
    layer2_outputs(7599) <= not (a xor b);
    layer2_outputs(7600) <= a;
    layer2_outputs(7601) <= not a;
    layer2_outputs(7602) <= not b;
    layer2_outputs(7603) <= not b;
    layer2_outputs(7604) <= a;
    layer2_outputs(7605) <= not (a or b);
    layer2_outputs(7606) <= a xor b;
    layer2_outputs(7607) <= not a;
    layer2_outputs(7608) <= a and not b;
    layer2_outputs(7609) <= a;
    layer2_outputs(7610) <= not (a and b);
    layer2_outputs(7611) <= a;
    layer2_outputs(7612) <= a and not b;
    layer2_outputs(7613) <= a and b;
    layer2_outputs(7614) <= not (a and b);
    layer2_outputs(7615) <= not b;
    layer2_outputs(7616) <= not (a or b);
    layer2_outputs(7617) <= b and not a;
    layer2_outputs(7618) <= not b;
    layer2_outputs(7619) <= not (a or b);
    layer2_outputs(7620) <= a and b;
    layer2_outputs(7621) <= not a;
    layer2_outputs(7622) <= b and not a;
    layer2_outputs(7623) <= not b or a;
    layer2_outputs(7624) <= '0';
    layer2_outputs(7625) <= a and not b;
    layer2_outputs(7626) <= not a;
    layer2_outputs(7627) <= not a;
    layer2_outputs(7628) <= not (a xor b);
    layer2_outputs(7629) <= a xor b;
    layer2_outputs(7630) <= not (a xor b);
    layer2_outputs(7631) <= a and not b;
    layer2_outputs(7632) <= not a;
    layer2_outputs(7633) <= not a;
    layer2_outputs(7634) <= a xor b;
    layer2_outputs(7635) <= not b;
    layer2_outputs(7636) <= not b or a;
    layer2_outputs(7637) <= b;
    layer2_outputs(7638) <= a or b;
    layer2_outputs(7639) <= a and not b;
    layer2_outputs(7640) <= not b or a;
    layer2_outputs(7641) <= a xor b;
    layer2_outputs(7642) <= '1';
    layer2_outputs(7643) <= a and b;
    layer2_outputs(7644) <= not (a and b);
    layer2_outputs(7645) <= not (a and b);
    layer2_outputs(7646) <= not (a and b);
    layer2_outputs(7647) <= b;
    layer2_outputs(7648) <= a and not b;
    layer2_outputs(7649) <= a and not b;
    layer2_outputs(7650) <= not a;
    layer2_outputs(7651) <= a;
    layer2_outputs(7652) <= a or b;
    layer2_outputs(7653) <= not (a and b);
    layer2_outputs(7654) <= b;
    layer2_outputs(7655) <= not (a or b);
    layer2_outputs(7656) <= b;
    layer2_outputs(7657) <= a or b;
    layer2_outputs(7658) <= not b;
    layer2_outputs(7659) <= not (a and b);
    layer2_outputs(7660) <= a xor b;
    layer2_outputs(7661) <= b;
    layer2_outputs(7662) <= not a or b;
    layer2_outputs(7663) <= b;
    layer2_outputs(7664) <= not (a and b);
    layer2_outputs(7665) <= a and not b;
    layer2_outputs(7666) <= not b;
    layer2_outputs(7667) <= a xor b;
    layer2_outputs(7668) <= not a;
    layer2_outputs(7669) <= not b or a;
    layer2_outputs(7670) <= a and b;
    layer2_outputs(7671) <= a xor b;
    layer2_outputs(7672) <= not a;
    layer2_outputs(7673) <= a;
    layer2_outputs(7674) <= not (a and b);
    layer2_outputs(7675) <= a and b;
    layer2_outputs(7676) <= a or b;
    layer2_outputs(7677) <= b and not a;
    layer2_outputs(7678) <= a or b;
    layer2_outputs(7679) <= a;
    layer2_outputs(7680) <= a or b;
    layer2_outputs(7681) <= not b;
    layer2_outputs(7682) <= b and not a;
    layer2_outputs(7683) <= not (a xor b);
    layer2_outputs(7684) <= not a;
    layer2_outputs(7685) <= not (a and b);
    layer2_outputs(7686) <= a or b;
    layer2_outputs(7687) <= b and not a;
    layer2_outputs(7688) <= not a;
    layer2_outputs(7689) <= a xor b;
    layer2_outputs(7690) <= b;
    layer2_outputs(7691) <= not a or b;
    layer2_outputs(7692) <= not b or a;
    layer2_outputs(7693) <= not a or b;
    layer2_outputs(7694) <= a xor b;
    layer2_outputs(7695) <= b;
    layer2_outputs(7696) <= a xor b;
    layer2_outputs(7697) <= not (a xor b);
    layer2_outputs(7698) <= not (a xor b);
    layer2_outputs(7699) <= a xor b;
    layer2_outputs(7700) <= a;
    layer2_outputs(7701) <= a and not b;
    layer2_outputs(7702) <= not a;
    layer2_outputs(7703) <= not (a and b);
    layer2_outputs(7704) <= a and not b;
    layer2_outputs(7705) <= a;
    layer2_outputs(7706) <= not b or a;
    layer2_outputs(7707) <= b;
    layer2_outputs(7708) <= a or b;
    layer2_outputs(7709) <= b;
    layer2_outputs(7710) <= a;
    layer2_outputs(7711) <= not b;
    layer2_outputs(7712) <= a and b;
    layer2_outputs(7713) <= a xor b;
    layer2_outputs(7714) <= b;
    layer2_outputs(7715) <= not (a or b);
    layer2_outputs(7716) <= not a or b;
    layer2_outputs(7717) <= not b;
    layer2_outputs(7718) <= b and not a;
    layer2_outputs(7719) <= not a;
    layer2_outputs(7720) <= a xor b;
    layer2_outputs(7721) <= not b;
    layer2_outputs(7722) <= not a;
    layer2_outputs(7723) <= a;
    layer2_outputs(7724) <= not a or b;
    layer2_outputs(7725) <= not b;
    layer2_outputs(7726) <= not (a xor b);
    layer2_outputs(7727) <= b;
    layer2_outputs(7728) <= a and not b;
    layer2_outputs(7729) <= a xor b;
    layer2_outputs(7730) <= not a or b;
    layer2_outputs(7731) <= not b;
    layer2_outputs(7732) <= not (a or b);
    layer2_outputs(7733) <= not b;
    layer2_outputs(7734) <= a xor b;
    layer2_outputs(7735) <= a or b;
    layer2_outputs(7736) <= a and not b;
    layer2_outputs(7737) <= not a;
    layer2_outputs(7738) <= not b;
    layer2_outputs(7739) <= b;
    layer2_outputs(7740) <= not a;
    layer2_outputs(7741) <= not (a or b);
    layer2_outputs(7742) <= a;
    layer2_outputs(7743) <= not (a and b);
    layer2_outputs(7744) <= a and b;
    layer2_outputs(7745) <= a xor b;
    layer2_outputs(7746) <= a xor b;
    layer2_outputs(7747) <= a and not b;
    layer2_outputs(7748) <= not (a or b);
    layer2_outputs(7749) <= not b or a;
    layer2_outputs(7750) <= a xor b;
    layer2_outputs(7751) <= b;
    layer2_outputs(7752) <= b;
    layer2_outputs(7753) <= a xor b;
    layer2_outputs(7754) <= b;
    layer2_outputs(7755) <= a;
    layer2_outputs(7756) <= a and not b;
    layer2_outputs(7757) <= a xor b;
    layer2_outputs(7758) <= a;
    layer2_outputs(7759) <= not (a or b);
    layer2_outputs(7760) <= not (a or b);
    layer2_outputs(7761) <= a and not b;
    layer2_outputs(7762) <= a and b;
    layer2_outputs(7763) <= a;
    layer2_outputs(7764) <= a xor b;
    layer2_outputs(7765) <= a and b;
    layer2_outputs(7766) <= a;
    layer2_outputs(7767) <= a and not b;
    layer2_outputs(7768) <= a and not b;
    layer2_outputs(7769) <= not a;
    layer2_outputs(7770) <= not b;
    layer2_outputs(7771) <= not (a xor b);
    layer2_outputs(7772) <= a or b;
    layer2_outputs(7773) <= a xor b;
    layer2_outputs(7774) <= a or b;
    layer2_outputs(7775) <= not b or a;
    layer2_outputs(7776) <= not (a or b);
    layer2_outputs(7777) <= a;
    layer2_outputs(7778) <= not (a or b);
    layer2_outputs(7779) <= not b;
    layer2_outputs(7780) <= not a;
    layer2_outputs(7781) <= a xor b;
    layer2_outputs(7782) <= not (a and b);
    layer2_outputs(7783) <= not (a xor b);
    layer2_outputs(7784) <= b and not a;
    layer2_outputs(7785) <= not b;
    layer2_outputs(7786) <= a or b;
    layer2_outputs(7787) <= b;
    layer2_outputs(7788) <= a xor b;
    layer2_outputs(7789) <= not b;
    layer2_outputs(7790) <= not b or a;
    layer2_outputs(7791) <= a xor b;
    layer2_outputs(7792) <= not a;
    layer2_outputs(7793) <= a and b;
    layer2_outputs(7794) <= b and not a;
    layer2_outputs(7795) <= a;
    layer2_outputs(7796) <= not b;
    layer2_outputs(7797) <= not b or a;
    layer2_outputs(7798) <= a;
    layer2_outputs(7799) <= a and not b;
    layer2_outputs(7800) <= a xor b;
    layer2_outputs(7801) <= a xor b;
    layer2_outputs(7802) <= a xor b;
    layer2_outputs(7803) <= not (a xor b);
    layer2_outputs(7804) <= a xor b;
    layer2_outputs(7805) <= b;
    layer2_outputs(7806) <= not a;
    layer2_outputs(7807) <= not (a and b);
    layer2_outputs(7808) <= not a;
    layer2_outputs(7809) <= not (a xor b);
    layer2_outputs(7810) <= not (a xor b);
    layer2_outputs(7811) <= '0';
    layer2_outputs(7812) <= a and b;
    layer2_outputs(7813) <= not a;
    layer2_outputs(7814) <= a and b;
    layer2_outputs(7815) <= not a;
    layer2_outputs(7816) <= not b or a;
    layer2_outputs(7817) <= a and b;
    layer2_outputs(7818) <= not (a xor b);
    layer2_outputs(7819) <= not a;
    layer2_outputs(7820) <= not (a xor b);
    layer2_outputs(7821) <= b;
    layer2_outputs(7822) <= not a or b;
    layer2_outputs(7823) <= not a;
    layer2_outputs(7824) <= a;
    layer2_outputs(7825) <= a and b;
    layer2_outputs(7826) <= a xor b;
    layer2_outputs(7827) <= not a or b;
    layer2_outputs(7828) <= not b;
    layer2_outputs(7829) <= b and not a;
    layer2_outputs(7830) <= not b;
    layer2_outputs(7831) <= not a;
    layer2_outputs(7832) <= not (a xor b);
    layer2_outputs(7833) <= a or b;
    layer2_outputs(7834) <= not b;
    layer2_outputs(7835) <= not b;
    layer2_outputs(7836) <= b;
    layer2_outputs(7837) <= a xor b;
    layer2_outputs(7838) <= not b;
    layer2_outputs(7839) <= a xor b;
    layer2_outputs(7840) <= not b;
    layer2_outputs(7841) <= a;
    layer2_outputs(7842) <= not a;
    layer2_outputs(7843) <= not b;
    layer2_outputs(7844) <= not (a and b);
    layer2_outputs(7845) <= not b;
    layer2_outputs(7846) <= not a;
    layer2_outputs(7847) <= a;
    layer2_outputs(7848) <= a xor b;
    layer2_outputs(7849) <= b and not a;
    layer2_outputs(7850) <= a or b;
    layer2_outputs(7851) <= b;
    layer2_outputs(7852) <= a;
    layer2_outputs(7853) <= a and b;
    layer2_outputs(7854) <= a;
    layer2_outputs(7855) <= not b;
    layer2_outputs(7856) <= b and not a;
    layer2_outputs(7857) <= b;
    layer2_outputs(7858) <= not a;
    layer2_outputs(7859) <= a and b;
    layer2_outputs(7860) <= a xor b;
    layer2_outputs(7861) <= a and not b;
    layer2_outputs(7862) <= not b;
    layer2_outputs(7863) <= not (a xor b);
    layer2_outputs(7864) <= a;
    layer2_outputs(7865) <= a xor b;
    layer2_outputs(7866) <= not (a xor b);
    layer2_outputs(7867) <= not a;
    layer2_outputs(7868) <= not b or a;
    layer2_outputs(7869) <= not (a xor b);
    layer2_outputs(7870) <= b;
    layer2_outputs(7871) <= a;
    layer2_outputs(7872) <= a and b;
    layer2_outputs(7873) <= not (a xor b);
    layer2_outputs(7874) <= not (a xor b);
    layer2_outputs(7875) <= a and b;
    layer2_outputs(7876) <= not b or a;
    layer2_outputs(7877) <= b;
    layer2_outputs(7878) <= b;
    layer2_outputs(7879) <= not a or b;
    layer2_outputs(7880) <= a;
    layer2_outputs(7881) <= b and not a;
    layer2_outputs(7882) <= b;
    layer2_outputs(7883) <= not b;
    layer2_outputs(7884) <= a or b;
    layer2_outputs(7885) <= not b or a;
    layer2_outputs(7886) <= b;
    layer2_outputs(7887) <= not b;
    layer2_outputs(7888) <= not b;
    layer2_outputs(7889) <= not a;
    layer2_outputs(7890) <= not (a and b);
    layer2_outputs(7891) <= b and not a;
    layer2_outputs(7892) <= a xor b;
    layer2_outputs(7893) <= not b;
    layer2_outputs(7894) <= a;
    layer2_outputs(7895) <= not a;
    layer2_outputs(7896) <= a or b;
    layer2_outputs(7897) <= not a or b;
    layer2_outputs(7898) <= a or b;
    layer2_outputs(7899) <= not (a and b);
    layer2_outputs(7900) <= b;
    layer2_outputs(7901) <= a xor b;
    layer2_outputs(7902) <= a or b;
    layer2_outputs(7903) <= a and b;
    layer2_outputs(7904) <= not b;
    layer2_outputs(7905) <= not a or b;
    layer2_outputs(7906) <= not a;
    layer2_outputs(7907) <= b and not a;
    layer2_outputs(7908) <= not (a or b);
    layer2_outputs(7909) <= a;
    layer2_outputs(7910) <= a and b;
    layer2_outputs(7911) <= b;
    layer2_outputs(7912) <= b;
    layer2_outputs(7913) <= a and b;
    layer2_outputs(7914) <= b and not a;
    layer2_outputs(7915) <= not (a xor b);
    layer2_outputs(7916) <= b;
    layer2_outputs(7917) <= a;
    layer2_outputs(7918) <= not a or b;
    layer2_outputs(7919) <= not a;
    layer2_outputs(7920) <= b and not a;
    layer2_outputs(7921) <= a or b;
    layer2_outputs(7922) <= not a;
    layer2_outputs(7923) <= a and b;
    layer2_outputs(7924) <= a and not b;
    layer2_outputs(7925) <= not a;
    layer2_outputs(7926) <= a or b;
    layer2_outputs(7927) <= not a or b;
    layer2_outputs(7928) <= not (a xor b);
    layer2_outputs(7929) <= b;
    layer2_outputs(7930) <= b;
    layer2_outputs(7931) <= b and not a;
    layer2_outputs(7932) <= not b;
    layer2_outputs(7933) <= not b;
    layer2_outputs(7934) <= not a or b;
    layer2_outputs(7935) <= not a;
    layer2_outputs(7936) <= not a or b;
    layer2_outputs(7937) <= a or b;
    layer2_outputs(7938) <= not (a or b);
    layer2_outputs(7939) <= not (a xor b);
    layer2_outputs(7940) <= not b;
    layer2_outputs(7941) <= not a or b;
    layer2_outputs(7942) <= '0';
    layer2_outputs(7943) <= not (a xor b);
    layer2_outputs(7944) <= a and b;
    layer2_outputs(7945) <= a and not b;
    layer2_outputs(7946) <= not a;
    layer2_outputs(7947) <= not b or a;
    layer2_outputs(7948) <= a and b;
    layer2_outputs(7949) <= b;
    layer2_outputs(7950) <= not a;
    layer2_outputs(7951) <= a and not b;
    layer2_outputs(7952) <= not (a or b);
    layer2_outputs(7953) <= b;
    layer2_outputs(7954) <= a;
    layer2_outputs(7955) <= not b or a;
    layer2_outputs(7956) <= a or b;
    layer2_outputs(7957) <= not (a xor b);
    layer2_outputs(7958) <= a or b;
    layer2_outputs(7959) <= '1';
    layer2_outputs(7960) <= a and b;
    layer2_outputs(7961) <= '1';
    layer2_outputs(7962) <= not (a xor b);
    layer2_outputs(7963) <= not (a and b);
    layer2_outputs(7964) <= not b;
    layer2_outputs(7965) <= not b or a;
    layer2_outputs(7966) <= not (a xor b);
    layer2_outputs(7967) <= not a;
    layer2_outputs(7968) <= a or b;
    layer2_outputs(7969) <= not b or a;
    layer2_outputs(7970) <= not a;
    layer2_outputs(7971) <= a or b;
    layer2_outputs(7972) <= a and b;
    layer2_outputs(7973) <= a;
    layer2_outputs(7974) <= not (a or b);
    layer2_outputs(7975) <= not b;
    layer2_outputs(7976) <= a or b;
    layer2_outputs(7977) <= not (a and b);
    layer2_outputs(7978) <= not (a xor b);
    layer2_outputs(7979) <= not a or b;
    layer2_outputs(7980) <= b and not a;
    layer2_outputs(7981) <= a or b;
    layer2_outputs(7982) <= a;
    layer2_outputs(7983) <= a xor b;
    layer2_outputs(7984) <= not a or b;
    layer2_outputs(7985) <= not (a xor b);
    layer2_outputs(7986) <= not (a and b);
    layer2_outputs(7987) <= not (a or b);
    layer2_outputs(7988) <= a xor b;
    layer2_outputs(7989) <= not a or b;
    layer2_outputs(7990) <= a or b;
    layer2_outputs(7991) <= not a;
    layer2_outputs(7992) <= not (a and b);
    layer2_outputs(7993) <= a;
    layer2_outputs(7994) <= not (a or b);
    layer2_outputs(7995) <= a xor b;
    layer2_outputs(7996) <= not a;
    layer2_outputs(7997) <= b and not a;
    layer2_outputs(7998) <= not b or a;
    layer2_outputs(7999) <= not (a xor b);
    layer2_outputs(8000) <= not (a xor b);
    layer2_outputs(8001) <= not b;
    layer2_outputs(8002) <= not (a and b);
    layer2_outputs(8003) <= not a;
    layer2_outputs(8004) <= b;
    layer2_outputs(8005) <= not b;
    layer2_outputs(8006) <= a or b;
    layer2_outputs(8007) <= not b or a;
    layer2_outputs(8008) <= a and not b;
    layer2_outputs(8009) <= not b;
    layer2_outputs(8010) <= a xor b;
    layer2_outputs(8011) <= a xor b;
    layer2_outputs(8012) <= not (a xor b);
    layer2_outputs(8013) <= not (a and b);
    layer2_outputs(8014) <= a;
    layer2_outputs(8015) <= not a or b;
    layer2_outputs(8016) <= not (a xor b);
    layer2_outputs(8017) <= not (a xor b);
    layer2_outputs(8018) <= not b;
    layer2_outputs(8019) <= a xor b;
    layer2_outputs(8020) <= b;
    layer2_outputs(8021) <= not (a xor b);
    layer2_outputs(8022) <= a xor b;
    layer2_outputs(8023) <= not (a or b);
    layer2_outputs(8024) <= a or b;
    layer2_outputs(8025) <= a xor b;
    layer2_outputs(8026) <= a or b;
    layer2_outputs(8027) <= not (a or b);
    layer2_outputs(8028) <= a and b;
    layer2_outputs(8029) <= '0';
    layer2_outputs(8030) <= not (a and b);
    layer2_outputs(8031) <= not a or b;
    layer2_outputs(8032) <= a xor b;
    layer2_outputs(8033) <= a or b;
    layer2_outputs(8034) <= b and not a;
    layer2_outputs(8035) <= not (a or b);
    layer2_outputs(8036) <= b;
    layer2_outputs(8037) <= not a;
    layer2_outputs(8038) <= not (a or b);
    layer2_outputs(8039) <= b;
    layer2_outputs(8040) <= a or b;
    layer2_outputs(8041) <= a and b;
    layer2_outputs(8042) <= not (a xor b);
    layer2_outputs(8043) <= not b;
    layer2_outputs(8044) <= not b;
    layer2_outputs(8045) <= not a;
    layer2_outputs(8046) <= b;
    layer2_outputs(8047) <= not a;
    layer2_outputs(8048) <= not (a xor b);
    layer2_outputs(8049) <= a and b;
    layer2_outputs(8050) <= not a;
    layer2_outputs(8051) <= not a;
    layer2_outputs(8052) <= b;
    layer2_outputs(8053) <= not (a xor b);
    layer2_outputs(8054) <= not a;
    layer2_outputs(8055) <= not a or b;
    layer2_outputs(8056) <= not b;
    layer2_outputs(8057) <= not (a and b);
    layer2_outputs(8058) <= not (a xor b);
    layer2_outputs(8059) <= not a or b;
    layer2_outputs(8060) <= a;
    layer2_outputs(8061) <= not b;
    layer2_outputs(8062) <= a or b;
    layer2_outputs(8063) <= not (a or b);
    layer2_outputs(8064) <= a;
    layer2_outputs(8065) <= not (a xor b);
    layer2_outputs(8066) <= not (a or b);
    layer2_outputs(8067) <= not (a xor b);
    layer2_outputs(8068) <= not b or a;
    layer2_outputs(8069) <= not b;
    layer2_outputs(8070) <= b;
    layer2_outputs(8071) <= a;
    layer2_outputs(8072) <= a or b;
    layer2_outputs(8073) <= '1';
    layer2_outputs(8074) <= b and not a;
    layer2_outputs(8075) <= a;
    layer2_outputs(8076) <= not a or b;
    layer2_outputs(8077) <= not (a xor b);
    layer2_outputs(8078) <= not (a xor b);
    layer2_outputs(8079) <= a;
    layer2_outputs(8080) <= a or b;
    layer2_outputs(8081) <= not a;
    layer2_outputs(8082) <= a and not b;
    layer2_outputs(8083) <= not b;
    layer2_outputs(8084) <= not (a or b);
    layer2_outputs(8085) <= b and not a;
    layer2_outputs(8086) <= b and not a;
    layer2_outputs(8087) <= b;
    layer2_outputs(8088) <= a xor b;
    layer2_outputs(8089) <= not b or a;
    layer2_outputs(8090) <= a xor b;
    layer2_outputs(8091) <= a;
    layer2_outputs(8092) <= not b;
    layer2_outputs(8093) <= a and b;
    layer2_outputs(8094) <= not b;
    layer2_outputs(8095) <= a and not b;
    layer2_outputs(8096) <= not a;
    layer2_outputs(8097) <= not a;
    layer2_outputs(8098) <= a or b;
    layer2_outputs(8099) <= b and not a;
    layer2_outputs(8100) <= b;
    layer2_outputs(8101) <= not b;
    layer2_outputs(8102) <= not a;
    layer2_outputs(8103) <= b and not a;
    layer2_outputs(8104) <= a and b;
    layer2_outputs(8105) <= b;
    layer2_outputs(8106) <= b;
    layer2_outputs(8107) <= a and not b;
    layer2_outputs(8108) <= a and not b;
    layer2_outputs(8109) <= a;
    layer2_outputs(8110) <= a and not b;
    layer2_outputs(8111) <= a and b;
    layer2_outputs(8112) <= a xor b;
    layer2_outputs(8113) <= a;
    layer2_outputs(8114) <= not (a or b);
    layer2_outputs(8115) <= b and not a;
    layer2_outputs(8116) <= not (a or b);
    layer2_outputs(8117) <= a;
    layer2_outputs(8118) <= b;
    layer2_outputs(8119) <= not (a or b);
    layer2_outputs(8120) <= not (a and b);
    layer2_outputs(8121) <= a and b;
    layer2_outputs(8122) <= not a;
    layer2_outputs(8123) <= a and not b;
    layer2_outputs(8124) <= a;
    layer2_outputs(8125) <= b;
    layer2_outputs(8126) <= b and not a;
    layer2_outputs(8127) <= not a;
    layer2_outputs(8128) <= b;
    layer2_outputs(8129) <= '1';
    layer2_outputs(8130) <= not a or b;
    layer2_outputs(8131) <= not b;
    layer2_outputs(8132) <= '1';
    layer2_outputs(8133) <= not (a and b);
    layer2_outputs(8134) <= b and not a;
    layer2_outputs(8135) <= not (a and b);
    layer2_outputs(8136) <= a and b;
    layer2_outputs(8137) <= not b;
    layer2_outputs(8138) <= not (a xor b);
    layer2_outputs(8139) <= not a or b;
    layer2_outputs(8140) <= a xor b;
    layer2_outputs(8141) <= a or b;
    layer2_outputs(8142) <= b;
    layer2_outputs(8143) <= b;
    layer2_outputs(8144) <= not (a xor b);
    layer2_outputs(8145) <= b;
    layer2_outputs(8146) <= a xor b;
    layer2_outputs(8147) <= b and not a;
    layer2_outputs(8148) <= a and b;
    layer2_outputs(8149) <= not (a xor b);
    layer2_outputs(8150) <= a and not b;
    layer2_outputs(8151) <= not (a or b);
    layer2_outputs(8152) <= not (a xor b);
    layer2_outputs(8153) <= not b;
    layer2_outputs(8154) <= not a;
    layer2_outputs(8155) <= not b or a;
    layer2_outputs(8156) <= not a;
    layer2_outputs(8157) <= not b or a;
    layer2_outputs(8158) <= a xor b;
    layer2_outputs(8159) <= not (a and b);
    layer2_outputs(8160) <= not (a xor b);
    layer2_outputs(8161) <= a xor b;
    layer2_outputs(8162) <= a;
    layer2_outputs(8163) <= not (a or b);
    layer2_outputs(8164) <= not b;
    layer2_outputs(8165) <= a xor b;
    layer2_outputs(8166) <= a;
    layer2_outputs(8167) <= a xor b;
    layer2_outputs(8168) <= not (a or b);
    layer2_outputs(8169) <= a or b;
    layer2_outputs(8170) <= not a;
    layer2_outputs(8171) <= a or b;
    layer2_outputs(8172) <= not a;
    layer2_outputs(8173) <= a;
    layer2_outputs(8174) <= a and not b;
    layer2_outputs(8175) <= b;
    layer2_outputs(8176) <= not a;
    layer2_outputs(8177) <= not a or b;
    layer2_outputs(8178) <= a or b;
    layer2_outputs(8179) <= not b;
    layer2_outputs(8180) <= not a;
    layer2_outputs(8181) <= not b or a;
    layer2_outputs(8182) <= a and not b;
    layer2_outputs(8183) <= not a;
    layer2_outputs(8184) <= not a or b;
    layer2_outputs(8185) <= b;
    layer2_outputs(8186) <= b;
    layer2_outputs(8187) <= a xor b;
    layer2_outputs(8188) <= not a;
    layer2_outputs(8189) <= a and b;
    layer2_outputs(8190) <= not b;
    layer2_outputs(8191) <= a and not b;
    layer2_outputs(8192) <= a xor b;
    layer2_outputs(8193) <= not (a xor b);
    layer2_outputs(8194) <= not a or b;
    layer2_outputs(8195) <= not (a xor b);
    layer2_outputs(8196) <= not (a xor b);
    layer2_outputs(8197) <= b;
    layer2_outputs(8198) <= a xor b;
    layer2_outputs(8199) <= not b;
    layer2_outputs(8200) <= not b or a;
    layer2_outputs(8201) <= not a;
    layer2_outputs(8202) <= b;
    layer2_outputs(8203) <= a xor b;
    layer2_outputs(8204) <= not b;
    layer2_outputs(8205) <= b;
    layer2_outputs(8206) <= not a or b;
    layer2_outputs(8207) <= not b or a;
    layer2_outputs(8208) <= b;
    layer2_outputs(8209) <= not a or b;
    layer2_outputs(8210) <= not b;
    layer2_outputs(8211) <= not (a xor b);
    layer2_outputs(8212) <= b;
    layer2_outputs(8213) <= not b;
    layer2_outputs(8214) <= a xor b;
    layer2_outputs(8215) <= a and not b;
    layer2_outputs(8216) <= a or b;
    layer2_outputs(8217) <= a and not b;
    layer2_outputs(8218) <= not (a xor b);
    layer2_outputs(8219) <= a;
    layer2_outputs(8220) <= b;
    layer2_outputs(8221) <= not a;
    layer2_outputs(8222) <= a xor b;
    layer2_outputs(8223) <= b;
    layer2_outputs(8224) <= a or b;
    layer2_outputs(8225) <= not (a and b);
    layer2_outputs(8226) <= a and not b;
    layer2_outputs(8227) <= b;
    layer2_outputs(8228) <= a;
    layer2_outputs(8229) <= not a;
    layer2_outputs(8230) <= a or b;
    layer2_outputs(8231) <= not a;
    layer2_outputs(8232) <= not a;
    layer2_outputs(8233) <= not (a xor b);
    layer2_outputs(8234) <= not a;
    layer2_outputs(8235) <= a;
    layer2_outputs(8236) <= '0';
    layer2_outputs(8237) <= b;
    layer2_outputs(8238) <= not a;
    layer2_outputs(8239) <= not (a xor b);
    layer2_outputs(8240) <= b;
    layer2_outputs(8241) <= not b;
    layer2_outputs(8242) <= a;
    layer2_outputs(8243) <= not (a or b);
    layer2_outputs(8244) <= a;
    layer2_outputs(8245) <= not a;
    layer2_outputs(8246) <= not (a xor b);
    layer2_outputs(8247) <= b;
    layer2_outputs(8248) <= a and not b;
    layer2_outputs(8249) <= not b;
    layer2_outputs(8250) <= a or b;
    layer2_outputs(8251) <= a and b;
    layer2_outputs(8252) <= not a;
    layer2_outputs(8253) <= b and not a;
    layer2_outputs(8254) <= not (a xor b);
    layer2_outputs(8255) <= not a or b;
    layer2_outputs(8256) <= not a;
    layer2_outputs(8257) <= not a or b;
    layer2_outputs(8258) <= not (a and b);
    layer2_outputs(8259) <= b and not a;
    layer2_outputs(8260) <= not (a and b);
    layer2_outputs(8261) <= a or b;
    layer2_outputs(8262) <= not a or b;
    layer2_outputs(8263) <= a and b;
    layer2_outputs(8264) <= not a;
    layer2_outputs(8265) <= not a;
    layer2_outputs(8266) <= a and not b;
    layer2_outputs(8267) <= not (a and b);
    layer2_outputs(8268) <= a and b;
    layer2_outputs(8269) <= a;
    layer2_outputs(8270) <= b;
    layer2_outputs(8271) <= not b;
    layer2_outputs(8272) <= a;
    layer2_outputs(8273) <= not a or b;
    layer2_outputs(8274) <= a;
    layer2_outputs(8275) <= not (a xor b);
    layer2_outputs(8276) <= b and not a;
    layer2_outputs(8277) <= not b;
    layer2_outputs(8278) <= a and not b;
    layer2_outputs(8279) <= a xor b;
    layer2_outputs(8280) <= not a;
    layer2_outputs(8281) <= b and not a;
    layer2_outputs(8282) <= a;
    layer2_outputs(8283) <= not b;
    layer2_outputs(8284) <= not b or a;
    layer2_outputs(8285) <= not b or a;
    layer2_outputs(8286) <= not (a and b);
    layer2_outputs(8287) <= a and b;
    layer2_outputs(8288) <= '0';
    layer2_outputs(8289) <= not b;
    layer2_outputs(8290) <= not (a xor b);
    layer2_outputs(8291) <= a and not b;
    layer2_outputs(8292) <= not (a or b);
    layer2_outputs(8293) <= not b;
    layer2_outputs(8294) <= a or b;
    layer2_outputs(8295) <= not b;
    layer2_outputs(8296) <= not a;
    layer2_outputs(8297) <= not b;
    layer2_outputs(8298) <= b and not a;
    layer2_outputs(8299) <= b;
    layer2_outputs(8300) <= not b;
    layer2_outputs(8301) <= a;
    layer2_outputs(8302) <= not (a or b);
    layer2_outputs(8303) <= not (a and b);
    layer2_outputs(8304) <= a and b;
    layer2_outputs(8305) <= not (a or b);
    layer2_outputs(8306) <= not b or a;
    layer2_outputs(8307) <= not b;
    layer2_outputs(8308) <= a;
    layer2_outputs(8309) <= a;
    layer2_outputs(8310) <= b;
    layer2_outputs(8311) <= not (a xor b);
    layer2_outputs(8312) <= not b;
    layer2_outputs(8313) <= a xor b;
    layer2_outputs(8314) <= b and not a;
    layer2_outputs(8315) <= not b or a;
    layer2_outputs(8316) <= a xor b;
    layer2_outputs(8317) <= b;
    layer2_outputs(8318) <= b;
    layer2_outputs(8319) <= not b;
    layer2_outputs(8320) <= not a;
    layer2_outputs(8321) <= a and not b;
    layer2_outputs(8322) <= a and b;
    layer2_outputs(8323) <= a or b;
    layer2_outputs(8324) <= b and not a;
    layer2_outputs(8325) <= a and not b;
    layer2_outputs(8326) <= a or b;
    layer2_outputs(8327) <= b;
    layer2_outputs(8328) <= not b;
    layer2_outputs(8329) <= not (a and b);
    layer2_outputs(8330) <= not (a or b);
    layer2_outputs(8331) <= not b or a;
    layer2_outputs(8332) <= b;
    layer2_outputs(8333) <= not b or a;
    layer2_outputs(8334) <= a or b;
    layer2_outputs(8335) <= a and not b;
    layer2_outputs(8336) <= not b;
    layer2_outputs(8337) <= not b;
    layer2_outputs(8338) <= a xor b;
    layer2_outputs(8339) <= b;
    layer2_outputs(8340) <= a xor b;
    layer2_outputs(8341) <= not (a xor b);
    layer2_outputs(8342) <= not a;
    layer2_outputs(8343) <= a and not b;
    layer2_outputs(8344) <= b;
    layer2_outputs(8345) <= a xor b;
    layer2_outputs(8346) <= a or b;
    layer2_outputs(8347) <= not a or b;
    layer2_outputs(8348) <= b and not a;
    layer2_outputs(8349) <= a;
    layer2_outputs(8350) <= a and not b;
    layer2_outputs(8351) <= b and not a;
    layer2_outputs(8352) <= a;
    layer2_outputs(8353) <= a and not b;
    layer2_outputs(8354) <= not b;
    layer2_outputs(8355) <= not b;
    layer2_outputs(8356) <= b and not a;
    layer2_outputs(8357) <= b and not a;
    layer2_outputs(8358) <= b and not a;
    layer2_outputs(8359) <= b and not a;
    layer2_outputs(8360) <= not a or b;
    layer2_outputs(8361) <= not (a and b);
    layer2_outputs(8362) <= a and not b;
    layer2_outputs(8363) <= b;
    layer2_outputs(8364) <= not a or b;
    layer2_outputs(8365) <= b and not a;
    layer2_outputs(8366) <= b;
    layer2_outputs(8367) <= a;
    layer2_outputs(8368) <= a;
    layer2_outputs(8369) <= not b or a;
    layer2_outputs(8370) <= not b;
    layer2_outputs(8371) <= a;
    layer2_outputs(8372) <= a xor b;
    layer2_outputs(8373) <= not a;
    layer2_outputs(8374) <= b and not a;
    layer2_outputs(8375) <= a xor b;
    layer2_outputs(8376) <= not b;
    layer2_outputs(8377) <= not a;
    layer2_outputs(8378) <= not b;
    layer2_outputs(8379) <= not b;
    layer2_outputs(8380) <= a and not b;
    layer2_outputs(8381) <= not (a and b);
    layer2_outputs(8382) <= '1';
    layer2_outputs(8383) <= b;
    layer2_outputs(8384) <= not (a and b);
    layer2_outputs(8385) <= not a;
    layer2_outputs(8386) <= not b;
    layer2_outputs(8387) <= not b;
    layer2_outputs(8388) <= b;
    layer2_outputs(8389) <= a and b;
    layer2_outputs(8390) <= not a;
    layer2_outputs(8391) <= not a or b;
    layer2_outputs(8392) <= a xor b;
    layer2_outputs(8393) <= not a;
    layer2_outputs(8394) <= a;
    layer2_outputs(8395) <= not (a and b);
    layer2_outputs(8396) <= not b;
    layer2_outputs(8397) <= not a or b;
    layer2_outputs(8398) <= b and not a;
    layer2_outputs(8399) <= a and b;
    layer2_outputs(8400) <= a;
    layer2_outputs(8401) <= not (a and b);
    layer2_outputs(8402) <= not b;
    layer2_outputs(8403) <= b;
    layer2_outputs(8404) <= not b or a;
    layer2_outputs(8405) <= a;
    layer2_outputs(8406) <= a xor b;
    layer2_outputs(8407) <= not a;
    layer2_outputs(8408) <= not a;
    layer2_outputs(8409) <= not a;
    layer2_outputs(8410) <= b and not a;
    layer2_outputs(8411) <= a;
    layer2_outputs(8412) <= not b;
    layer2_outputs(8413) <= a and not b;
    layer2_outputs(8414) <= b;
    layer2_outputs(8415) <= b;
    layer2_outputs(8416) <= a;
    layer2_outputs(8417) <= '1';
    layer2_outputs(8418) <= b;
    layer2_outputs(8419) <= not b;
    layer2_outputs(8420) <= a or b;
    layer2_outputs(8421) <= a or b;
    layer2_outputs(8422) <= not a;
    layer2_outputs(8423) <= not b;
    layer2_outputs(8424) <= b;
    layer2_outputs(8425) <= not a;
    layer2_outputs(8426) <= not b;
    layer2_outputs(8427) <= b and not a;
    layer2_outputs(8428) <= not b;
    layer2_outputs(8429) <= b and not a;
    layer2_outputs(8430) <= not (a or b);
    layer2_outputs(8431) <= not (a or b);
    layer2_outputs(8432) <= not a or b;
    layer2_outputs(8433) <= b;
    layer2_outputs(8434) <= not b or a;
    layer2_outputs(8435) <= a and b;
    layer2_outputs(8436) <= not (a and b);
    layer2_outputs(8437) <= not a;
    layer2_outputs(8438) <= a;
    layer2_outputs(8439) <= a;
    layer2_outputs(8440) <= a and not b;
    layer2_outputs(8441) <= b;
    layer2_outputs(8442) <= not a;
    layer2_outputs(8443) <= not a or b;
    layer2_outputs(8444) <= not a or b;
    layer2_outputs(8445) <= a and b;
    layer2_outputs(8446) <= a and b;
    layer2_outputs(8447) <= b;
    layer2_outputs(8448) <= a and b;
    layer2_outputs(8449) <= not (a or b);
    layer2_outputs(8450) <= not (a xor b);
    layer2_outputs(8451) <= a or b;
    layer2_outputs(8452) <= a;
    layer2_outputs(8453) <= a;
    layer2_outputs(8454) <= a;
    layer2_outputs(8455) <= a and b;
    layer2_outputs(8456) <= b;
    layer2_outputs(8457) <= a or b;
    layer2_outputs(8458) <= not b;
    layer2_outputs(8459) <= not b or a;
    layer2_outputs(8460) <= not a or b;
    layer2_outputs(8461) <= a and not b;
    layer2_outputs(8462) <= a xor b;
    layer2_outputs(8463) <= b and not a;
    layer2_outputs(8464) <= not (a xor b);
    layer2_outputs(8465) <= not (a xor b);
    layer2_outputs(8466) <= not b;
    layer2_outputs(8467) <= a xor b;
    layer2_outputs(8468) <= not b;
    layer2_outputs(8469) <= a;
    layer2_outputs(8470) <= a and b;
    layer2_outputs(8471) <= not (a or b);
    layer2_outputs(8472) <= a and not b;
    layer2_outputs(8473) <= a;
    layer2_outputs(8474) <= not b;
    layer2_outputs(8475) <= not a;
    layer2_outputs(8476) <= not b;
    layer2_outputs(8477) <= not b or a;
    layer2_outputs(8478) <= a;
    layer2_outputs(8479) <= '0';
    layer2_outputs(8480) <= not a;
    layer2_outputs(8481) <= a and b;
    layer2_outputs(8482) <= a or b;
    layer2_outputs(8483) <= not (a and b);
    layer2_outputs(8484) <= not a or b;
    layer2_outputs(8485) <= not b;
    layer2_outputs(8486) <= b;
    layer2_outputs(8487) <= a;
    layer2_outputs(8488) <= b;
    layer2_outputs(8489) <= a and b;
    layer2_outputs(8490) <= a xor b;
    layer2_outputs(8491) <= b;
    layer2_outputs(8492) <= not b;
    layer2_outputs(8493) <= not (a xor b);
    layer2_outputs(8494) <= a;
    layer2_outputs(8495) <= not (a and b);
    layer2_outputs(8496) <= not a;
    layer2_outputs(8497) <= not a;
    layer2_outputs(8498) <= a and not b;
    layer2_outputs(8499) <= not (a and b);
    layer2_outputs(8500) <= not b;
    layer2_outputs(8501) <= a and not b;
    layer2_outputs(8502) <= not a or b;
    layer2_outputs(8503) <= not b;
    layer2_outputs(8504) <= a;
    layer2_outputs(8505) <= b;
    layer2_outputs(8506) <= a;
    layer2_outputs(8507) <= not (a xor b);
    layer2_outputs(8508) <= a;
    layer2_outputs(8509) <= a xor b;
    layer2_outputs(8510) <= not b;
    layer2_outputs(8511) <= not b or a;
    layer2_outputs(8512) <= not b;
    layer2_outputs(8513) <= a and b;
    layer2_outputs(8514) <= not (a xor b);
    layer2_outputs(8515) <= a xor b;
    layer2_outputs(8516) <= a xor b;
    layer2_outputs(8517) <= not (a xor b);
    layer2_outputs(8518) <= a xor b;
    layer2_outputs(8519) <= not a or b;
    layer2_outputs(8520) <= not (a or b);
    layer2_outputs(8521) <= a or b;
    layer2_outputs(8522) <= not (a and b);
    layer2_outputs(8523) <= not (a xor b);
    layer2_outputs(8524) <= b;
    layer2_outputs(8525) <= not a;
    layer2_outputs(8526) <= not b;
    layer2_outputs(8527) <= not b or a;
    layer2_outputs(8528) <= a or b;
    layer2_outputs(8529) <= a and b;
    layer2_outputs(8530) <= not (a or b);
    layer2_outputs(8531) <= b;
    layer2_outputs(8532) <= a or b;
    layer2_outputs(8533) <= a;
    layer2_outputs(8534) <= a xor b;
    layer2_outputs(8535) <= not (a and b);
    layer2_outputs(8536) <= not b;
    layer2_outputs(8537) <= a and not b;
    layer2_outputs(8538) <= not (a and b);
    layer2_outputs(8539) <= a and b;
    layer2_outputs(8540) <= a and b;
    layer2_outputs(8541) <= a;
    layer2_outputs(8542) <= not a;
    layer2_outputs(8543) <= not (a xor b);
    layer2_outputs(8544) <= not b or a;
    layer2_outputs(8545) <= not (a or b);
    layer2_outputs(8546) <= not (a xor b);
    layer2_outputs(8547) <= not a or b;
    layer2_outputs(8548) <= not a or b;
    layer2_outputs(8549) <= not a or b;
    layer2_outputs(8550) <= a and b;
    layer2_outputs(8551) <= '0';
    layer2_outputs(8552) <= not a;
    layer2_outputs(8553) <= not b;
    layer2_outputs(8554) <= not b or a;
    layer2_outputs(8555) <= not (a xor b);
    layer2_outputs(8556) <= a or b;
    layer2_outputs(8557) <= a;
    layer2_outputs(8558) <= not (a or b);
    layer2_outputs(8559) <= b;
    layer2_outputs(8560) <= not a;
    layer2_outputs(8561) <= not (a and b);
    layer2_outputs(8562) <= a xor b;
    layer2_outputs(8563) <= b;
    layer2_outputs(8564) <= not b or a;
    layer2_outputs(8565) <= b;
    layer2_outputs(8566) <= a or b;
    layer2_outputs(8567) <= a and b;
    layer2_outputs(8568) <= not b;
    layer2_outputs(8569) <= not a;
    layer2_outputs(8570) <= a xor b;
    layer2_outputs(8571) <= not a;
    layer2_outputs(8572) <= not (a and b);
    layer2_outputs(8573) <= b;
    layer2_outputs(8574) <= not a;
    layer2_outputs(8575) <= a and b;
    layer2_outputs(8576) <= b and not a;
    layer2_outputs(8577) <= not a;
    layer2_outputs(8578) <= not a;
    layer2_outputs(8579) <= not a or b;
    layer2_outputs(8580) <= b;
    layer2_outputs(8581) <= not (a or b);
    layer2_outputs(8582) <= not b or a;
    layer2_outputs(8583) <= not (a xor b);
    layer2_outputs(8584) <= a xor b;
    layer2_outputs(8585) <= not (a xor b);
    layer2_outputs(8586) <= not a;
    layer2_outputs(8587) <= not (a or b);
    layer2_outputs(8588) <= a or b;
    layer2_outputs(8589) <= not b;
    layer2_outputs(8590) <= a;
    layer2_outputs(8591) <= not b or a;
    layer2_outputs(8592) <= not (a xor b);
    layer2_outputs(8593) <= b;
    layer2_outputs(8594) <= not b;
    layer2_outputs(8595) <= a;
    layer2_outputs(8596) <= not a or b;
    layer2_outputs(8597) <= not b;
    layer2_outputs(8598) <= a xor b;
    layer2_outputs(8599) <= a and not b;
    layer2_outputs(8600) <= a and b;
    layer2_outputs(8601) <= a;
    layer2_outputs(8602) <= b;
    layer2_outputs(8603) <= not a;
    layer2_outputs(8604) <= a;
    layer2_outputs(8605) <= not (a xor b);
    layer2_outputs(8606) <= not a or b;
    layer2_outputs(8607) <= b;
    layer2_outputs(8608) <= a or b;
    layer2_outputs(8609) <= b;
    layer2_outputs(8610) <= a or b;
    layer2_outputs(8611) <= not a;
    layer2_outputs(8612) <= a xor b;
    layer2_outputs(8613) <= a and b;
    layer2_outputs(8614) <= a xor b;
    layer2_outputs(8615) <= a;
    layer2_outputs(8616) <= not (a or b);
    layer2_outputs(8617) <= b and not a;
    layer2_outputs(8618) <= not a;
    layer2_outputs(8619) <= a or b;
    layer2_outputs(8620) <= b;
    layer2_outputs(8621) <= a and b;
    layer2_outputs(8622) <= a and not b;
    layer2_outputs(8623) <= not (a and b);
    layer2_outputs(8624) <= a and b;
    layer2_outputs(8625) <= a and not b;
    layer2_outputs(8626) <= not b;
    layer2_outputs(8627) <= not b or a;
    layer2_outputs(8628) <= a and b;
    layer2_outputs(8629) <= a;
    layer2_outputs(8630) <= not a;
    layer2_outputs(8631) <= not a;
    layer2_outputs(8632) <= b and not a;
    layer2_outputs(8633) <= a;
    layer2_outputs(8634) <= a;
    layer2_outputs(8635) <= not b;
    layer2_outputs(8636) <= a and not b;
    layer2_outputs(8637) <= not (a and b);
    layer2_outputs(8638) <= not (a xor b);
    layer2_outputs(8639) <= not b;
    layer2_outputs(8640) <= a xor b;
    layer2_outputs(8641) <= a or b;
    layer2_outputs(8642) <= not (a or b);
    layer2_outputs(8643) <= b and not a;
    layer2_outputs(8644) <= not (a xor b);
    layer2_outputs(8645) <= a or b;
    layer2_outputs(8646) <= a xor b;
    layer2_outputs(8647) <= a or b;
    layer2_outputs(8648) <= a or b;
    layer2_outputs(8649) <= a;
    layer2_outputs(8650) <= a and not b;
    layer2_outputs(8651) <= a;
    layer2_outputs(8652) <= not a;
    layer2_outputs(8653) <= not b or a;
    layer2_outputs(8654) <= a and not b;
    layer2_outputs(8655) <= not b;
    layer2_outputs(8656) <= a;
    layer2_outputs(8657) <= a;
    layer2_outputs(8658) <= not a or b;
    layer2_outputs(8659) <= a and not b;
    layer2_outputs(8660) <= a;
    layer2_outputs(8661) <= a;
    layer2_outputs(8662) <= '1';
    layer2_outputs(8663) <= not a;
    layer2_outputs(8664) <= not (a xor b);
    layer2_outputs(8665) <= not a;
    layer2_outputs(8666) <= a;
    layer2_outputs(8667) <= not b or a;
    layer2_outputs(8668) <= not (a xor b);
    layer2_outputs(8669) <= not b;
    layer2_outputs(8670) <= a;
    layer2_outputs(8671) <= not b or a;
    layer2_outputs(8672) <= not b;
    layer2_outputs(8673) <= a;
    layer2_outputs(8674) <= not (a or b);
    layer2_outputs(8675) <= not (a or b);
    layer2_outputs(8676) <= not (a and b);
    layer2_outputs(8677) <= a;
    layer2_outputs(8678) <= b;
    layer2_outputs(8679) <= not (a and b);
    layer2_outputs(8680) <= not b;
    layer2_outputs(8681) <= b;
    layer2_outputs(8682) <= not a;
    layer2_outputs(8683) <= b;
    layer2_outputs(8684) <= not a;
    layer2_outputs(8685) <= b;
    layer2_outputs(8686) <= not a or b;
    layer2_outputs(8687) <= not (a and b);
    layer2_outputs(8688) <= not (a or b);
    layer2_outputs(8689) <= b;
    layer2_outputs(8690) <= not b or a;
    layer2_outputs(8691) <= not a;
    layer2_outputs(8692) <= not a or b;
    layer2_outputs(8693) <= a and not b;
    layer2_outputs(8694) <= not b or a;
    layer2_outputs(8695) <= a xor b;
    layer2_outputs(8696) <= b and not a;
    layer2_outputs(8697) <= a and b;
    layer2_outputs(8698) <= not (a xor b);
    layer2_outputs(8699) <= a;
    layer2_outputs(8700) <= b and not a;
    layer2_outputs(8701) <= not b;
    layer2_outputs(8702) <= not a;
    layer2_outputs(8703) <= b;
    layer2_outputs(8704) <= not b or a;
    layer2_outputs(8705) <= not (a and b);
    layer2_outputs(8706) <= not a or b;
    layer2_outputs(8707) <= a;
    layer2_outputs(8708) <= not (a and b);
    layer2_outputs(8709) <= not (a xor b);
    layer2_outputs(8710) <= not a;
    layer2_outputs(8711) <= not a;
    layer2_outputs(8712) <= '1';
    layer2_outputs(8713) <= not (a and b);
    layer2_outputs(8714) <= b;
    layer2_outputs(8715) <= a and b;
    layer2_outputs(8716) <= not a;
    layer2_outputs(8717) <= not a or b;
    layer2_outputs(8718) <= b;
    layer2_outputs(8719) <= not (a xor b);
    layer2_outputs(8720) <= a xor b;
    layer2_outputs(8721) <= not (a and b);
    layer2_outputs(8722) <= a xor b;
    layer2_outputs(8723) <= a and b;
    layer2_outputs(8724) <= not b;
    layer2_outputs(8725) <= b;
    layer2_outputs(8726) <= not (a xor b);
    layer2_outputs(8727) <= b;
    layer2_outputs(8728) <= a;
    layer2_outputs(8729) <= a xor b;
    layer2_outputs(8730) <= not (a or b);
    layer2_outputs(8731) <= not b;
    layer2_outputs(8732) <= a;
    layer2_outputs(8733) <= not a or b;
    layer2_outputs(8734) <= a xor b;
    layer2_outputs(8735) <= a and b;
    layer2_outputs(8736) <= not a;
    layer2_outputs(8737) <= not a or b;
    layer2_outputs(8738) <= not (a xor b);
    layer2_outputs(8739) <= not a;
    layer2_outputs(8740) <= not (a xor b);
    layer2_outputs(8741) <= a and not b;
    layer2_outputs(8742) <= a or b;
    layer2_outputs(8743) <= a or b;
    layer2_outputs(8744) <= not a or b;
    layer2_outputs(8745) <= not (a xor b);
    layer2_outputs(8746) <= not a;
    layer2_outputs(8747) <= not b;
    layer2_outputs(8748) <= not (a xor b);
    layer2_outputs(8749) <= a xor b;
    layer2_outputs(8750) <= not b or a;
    layer2_outputs(8751) <= a;
    layer2_outputs(8752) <= b;
    layer2_outputs(8753) <= not a or b;
    layer2_outputs(8754) <= b;
    layer2_outputs(8755) <= not (a xor b);
    layer2_outputs(8756) <= a;
    layer2_outputs(8757) <= a xor b;
    layer2_outputs(8758) <= a xor b;
    layer2_outputs(8759) <= a and not b;
    layer2_outputs(8760) <= a or b;
    layer2_outputs(8761) <= a xor b;
    layer2_outputs(8762) <= not (a xor b);
    layer2_outputs(8763) <= a and not b;
    layer2_outputs(8764) <= a;
    layer2_outputs(8765) <= a or b;
    layer2_outputs(8766) <= a and not b;
    layer2_outputs(8767) <= not a or b;
    layer2_outputs(8768) <= a xor b;
    layer2_outputs(8769) <= b;
    layer2_outputs(8770) <= a;
    layer2_outputs(8771) <= not b;
    layer2_outputs(8772) <= a xor b;
    layer2_outputs(8773) <= not a;
    layer2_outputs(8774) <= not (a and b);
    layer2_outputs(8775) <= b and not a;
    layer2_outputs(8776) <= not (a xor b);
    layer2_outputs(8777) <= a;
    layer2_outputs(8778) <= a and b;
    layer2_outputs(8779) <= not b or a;
    layer2_outputs(8780) <= not b;
    layer2_outputs(8781) <= not (a and b);
    layer2_outputs(8782) <= not b or a;
    layer2_outputs(8783) <= not (a or b);
    layer2_outputs(8784) <= a and b;
    layer2_outputs(8785) <= not a;
    layer2_outputs(8786) <= not a;
    layer2_outputs(8787) <= b;
    layer2_outputs(8788) <= not b;
    layer2_outputs(8789) <= a and not b;
    layer2_outputs(8790) <= a or b;
    layer2_outputs(8791) <= not b;
    layer2_outputs(8792) <= not (a xor b);
    layer2_outputs(8793) <= not (a xor b);
    layer2_outputs(8794) <= not a;
    layer2_outputs(8795) <= not (a xor b);
    layer2_outputs(8796) <= a;
    layer2_outputs(8797) <= not a;
    layer2_outputs(8798) <= not a;
    layer2_outputs(8799) <= not b or a;
    layer2_outputs(8800) <= b and not a;
    layer2_outputs(8801) <= a and b;
    layer2_outputs(8802) <= not a or b;
    layer2_outputs(8803) <= a xor b;
    layer2_outputs(8804) <= a and b;
    layer2_outputs(8805) <= not (a or b);
    layer2_outputs(8806) <= not b;
    layer2_outputs(8807) <= a;
    layer2_outputs(8808) <= b;
    layer2_outputs(8809) <= not (a xor b);
    layer2_outputs(8810) <= not b or a;
    layer2_outputs(8811) <= not (a and b);
    layer2_outputs(8812) <= b;
    layer2_outputs(8813) <= b and not a;
    layer2_outputs(8814) <= not b;
    layer2_outputs(8815) <= a xor b;
    layer2_outputs(8816) <= a and b;
    layer2_outputs(8817) <= not b or a;
    layer2_outputs(8818) <= a xor b;
    layer2_outputs(8819) <= not (a and b);
    layer2_outputs(8820) <= a and not b;
    layer2_outputs(8821) <= not b;
    layer2_outputs(8822) <= b;
    layer2_outputs(8823) <= not a;
    layer2_outputs(8824) <= a or b;
    layer2_outputs(8825) <= b and not a;
    layer2_outputs(8826) <= b;
    layer2_outputs(8827) <= not b;
    layer2_outputs(8828) <= not (a or b);
    layer2_outputs(8829) <= a xor b;
    layer2_outputs(8830) <= a xor b;
    layer2_outputs(8831) <= b and not a;
    layer2_outputs(8832) <= not (a and b);
    layer2_outputs(8833) <= not b or a;
    layer2_outputs(8834) <= a;
    layer2_outputs(8835) <= not a;
    layer2_outputs(8836) <= a;
    layer2_outputs(8837) <= not b;
    layer2_outputs(8838) <= not a;
    layer2_outputs(8839) <= b;
    layer2_outputs(8840) <= a;
    layer2_outputs(8841) <= a and b;
    layer2_outputs(8842) <= not (a or b);
    layer2_outputs(8843) <= b;
    layer2_outputs(8844) <= a xor b;
    layer2_outputs(8845) <= not b;
    layer2_outputs(8846) <= not b;
    layer2_outputs(8847) <= not (a or b);
    layer2_outputs(8848) <= not (a or b);
    layer2_outputs(8849) <= a;
    layer2_outputs(8850) <= not b;
    layer2_outputs(8851) <= a;
    layer2_outputs(8852) <= b;
    layer2_outputs(8853) <= b and not a;
    layer2_outputs(8854) <= b;
    layer2_outputs(8855) <= a and not b;
    layer2_outputs(8856) <= a xor b;
    layer2_outputs(8857) <= not a or b;
    layer2_outputs(8858) <= not b or a;
    layer2_outputs(8859) <= not a or b;
    layer2_outputs(8860) <= not b;
    layer2_outputs(8861) <= a xor b;
    layer2_outputs(8862) <= not (a xor b);
    layer2_outputs(8863) <= not a;
    layer2_outputs(8864) <= a xor b;
    layer2_outputs(8865) <= not (a and b);
    layer2_outputs(8866) <= a and b;
    layer2_outputs(8867) <= not (a xor b);
    layer2_outputs(8868) <= a;
    layer2_outputs(8869) <= not (a and b);
    layer2_outputs(8870) <= b;
    layer2_outputs(8871) <= not (a or b);
    layer2_outputs(8872) <= '1';
    layer2_outputs(8873) <= a and not b;
    layer2_outputs(8874) <= b;
    layer2_outputs(8875) <= not (a xor b);
    layer2_outputs(8876) <= a;
    layer2_outputs(8877) <= b and not a;
    layer2_outputs(8878) <= b;
    layer2_outputs(8879) <= not a;
    layer2_outputs(8880) <= b;
    layer2_outputs(8881) <= a xor b;
    layer2_outputs(8882) <= not a;
    layer2_outputs(8883) <= not (a xor b);
    layer2_outputs(8884) <= a and b;
    layer2_outputs(8885) <= a xor b;
    layer2_outputs(8886) <= not (a and b);
    layer2_outputs(8887) <= a and b;
    layer2_outputs(8888) <= not a or b;
    layer2_outputs(8889) <= a;
    layer2_outputs(8890) <= a xor b;
    layer2_outputs(8891) <= a;
    layer2_outputs(8892) <= a xor b;
    layer2_outputs(8893) <= not a;
    layer2_outputs(8894) <= a;
    layer2_outputs(8895) <= not (a or b);
    layer2_outputs(8896) <= not b;
    layer2_outputs(8897) <= a;
    layer2_outputs(8898) <= a or b;
    layer2_outputs(8899) <= a or b;
    layer2_outputs(8900) <= not (a or b);
    layer2_outputs(8901) <= a and b;
    layer2_outputs(8902) <= b and not a;
    layer2_outputs(8903) <= b;
    layer2_outputs(8904) <= not a;
    layer2_outputs(8905) <= a;
    layer2_outputs(8906) <= not a;
    layer2_outputs(8907) <= not a;
    layer2_outputs(8908) <= not a;
    layer2_outputs(8909) <= b and not a;
    layer2_outputs(8910) <= not a;
    layer2_outputs(8911) <= not b or a;
    layer2_outputs(8912) <= not (a or b);
    layer2_outputs(8913) <= a xor b;
    layer2_outputs(8914) <= not (a and b);
    layer2_outputs(8915) <= not a;
    layer2_outputs(8916) <= not b;
    layer2_outputs(8917) <= a;
    layer2_outputs(8918) <= a and b;
    layer2_outputs(8919) <= not a or b;
    layer2_outputs(8920) <= not (a and b);
    layer2_outputs(8921) <= a and not b;
    layer2_outputs(8922) <= not b;
    layer2_outputs(8923) <= b;
    layer2_outputs(8924) <= not (a and b);
    layer2_outputs(8925) <= a xor b;
    layer2_outputs(8926) <= a and not b;
    layer2_outputs(8927) <= b and not a;
    layer2_outputs(8928) <= not a;
    layer2_outputs(8929) <= not a or b;
    layer2_outputs(8930) <= a and b;
    layer2_outputs(8931) <= not (a and b);
    layer2_outputs(8932) <= not (a and b);
    layer2_outputs(8933) <= not b;
    layer2_outputs(8934) <= not (a xor b);
    layer2_outputs(8935) <= not a;
    layer2_outputs(8936) <= not (a and b);
    layer2_outputs(8937) <= not a;
    layer2_outputs(8938) <= a or b;
    layer2_outputs(8939) <= not (a or b);
    layer2_outputs(8940) <= a;
    layer2_outputs(8941) <= not b or a;
    layer2_outputs(8942) <= not a;
    layer2_outputs(8943) <= not (a or b);
    layer2_outputs(8944) <= '0';
    layer2_outputs(8945) <= a xor b;
    layer2_outputs(8946) <= not a;
    layer2_outputs(8947) <= b;
    layer2_outputs(8948) <= a and b;
    layer2_outputs(8949) <= a and b;
    layer2_outputs(8950) <= a xor b;
    layer2_outputs(8951) <= b;
    layer2_outputs(8952) <= not b;
    layer2_outputs(8953) <= a xor b;
    layer2_outputs(8954) <= a and not b;
    layer2_outputs(8955) <= not b;
    layer2_outputs(8956) <= a xor b;
    layer2_outputs(8957) <= a;
    layer2_outputs(8958) <= not b or a;
    layer2_outputs(8959) <= a;
    layer2_outputs(8960) <= not a;
    layer2_outputs(8961) <= a and not b;
    layer2_outputs(8962) <= not b or a;
    layer2_outputs(8963) <= not b;
    layer2_outputs(8964) <= a;
    layer2_outputs(8965) <= a;
    layer2_outputs(8966) <= not b;
    layer2_outputs(8967) <= a xor b;
    layer2_outputs(8968) <= b;
    layer2_outputs(8969) <= not b or a;
    layer2_outputs(8970) <= not a or b;
    layer2_outputs(8971) <= not (a or b);
    layer2_outputs(8972) <= not (a or b);
    layer2_outputs(8973) <= a and b;
    layer2_outputs(8974) <= not a;
    layer2_outputs(8975) <= not b or a;
    layer2_outputs(8976) <= a xor b;
    layer2_outputs(8977) <= a xor b;
    layer2_outputs(8978) <= b;
    layer2_outputs(8979) <= not b;
    layer2_outputs(8980) <= not (a xor b);
    layer2_outputs(8981) <= not a;
    layer2_outputs(8982) <= a and not b;
    layer2_outputs(8983) <= not (a xor b);
    layer2_outputs(8984) <= b;
    layer2_outputs(8985) <= not a or b;
    layer2_outputs(8986) <= not a;
    layer2_outputs(8987) <= a and b;
    layer2_outputs(8988) <= not a;
    layer2_outputs(8989) <= not b or a;
    layer2_outputs(8990) <= a;
    layer2_outputs(8991) <= a or b;
    layer2_outputs(8992) <= b and not a;
    layer2_outputs(8993) <= not a;
    layer2_outputs(8994) <= b;
    layer2_outputs(8995) <= not a;
    layer2_outputs(8996) <= a xor b;
    layer2_outputs(8997) <= not (a xor b);
    layer2_outputs(8998) <= not b or a;
    layer2_outputs(8999) <= not (a and b);
    layer2_outputs(9000) <= not (a xor b);
    layer2_outputs(9001) <= not a or b;
    layer2_outputs(9002) <= a and not b;
    layer2_outputs(9003) <= not a;
    layer2_outputs(9004) <= not (a xor b);
    layer2_outputs(9005) <= not (a xor b);
    layer2_outputs(9006) <= a and not b;
    layer2_outputs(9007) <= a or b;
    layer2_outputs(9008) <= not (a xor b);
    layer2_outputs(9009) <= not (a xor b);
    layer2_outputs(9010) <= not (a and b);
    layer2_outputs(9011) <= a;
    layer2_outputs(9012) <= not (a xor b);
    layer2_outputs(9013) <= not (a and b);
    layer2_outputs(9014) <= not b;
    layer2_outputs(9015) <= not b or a;
    layer2_outputs(9016) <= not a or b;
    layer2_outputs(9017) <= not b or a;
    layer2_outputs(9018) <= not (a xor b);
    layer2_outputs(9019) <= not a;
    layer2_outputs(9020) <= not a;
    layer2_outputs(9021) <= b;
    layer2_outputs(9022) <= a;
    layer2_outputs(9023) <= b and not a;
    layer2_outputs(9024) <= a;
    layer2_outputs(9025) <= b;
    layer2_outputs(9026) <= a and b;
    layer2_outputs(9027) <= a xor b;
    layer2_outputs(9028) <= b;
    layer2_outputs(9029) <= not (a or b);
    layer2_outputs(9030) <= not (a xor b);
    layer2_outputs(9031) <= b;
    layer2_outputs(9032) <= a xor b;
    layer2_outputs(9033) <= not b;
    layer2_outputs(9034) <= a xor b;
    layer2_outputs(9035) <= a and b;
    layer2_outputs(9036) <= a or b;
    layer2_outputs(9037) <= not b;
    layer2_outputs(9038) <= a xor b;
    layer2_outputs(9039) <= b;
    layer2_outputs(9040) <= a xor b;
    layer2_outputs(9041) <= b and not a;
    layer2_outputs(9042) <= not (a xor b);
    layer2_outputs(9043) <= not (a xor b);
    layer2_outputs(9044) <= a;
    layer2_outputs(9045) <= b and not a;
    layer2_outputs(9046) <= not (a and b);
    layer2_outputs(9047) <= not (a and b);
    layer2_outputs(9048) <= a;
    layer2_outputs(9049) <= not b or a;
    layer2_outputs(9050) <= not a;
    layer2_outputs(9051) <= a;
    layer2_outputs(9052) <= b;
    layer2_outputs(9053) <= not a;
    layer2_outputs(9054) <= a or b;
    layer2_outputs(9055) <= a and b;
    layer2_outputs(9056) <= not a or b;
    layer2_outputs(9057) <= '0';
    layer2_outputs(9058) <= not a or b;
    layer2_outputs(9059) <= not (a xor b);
    layer2_outputs(9060) <= not b;
    layer2_outputs(9061) <= not a or b;
    layer2_outputs(9062) <= b;
    layer2_outputs(9063) <= a;
    layer2_outputs(9064) <= b and not a;
    layer2_outputs(9065) <= not (a and b);
    layer2_outputs(9066) <= a xor b;
    layer2_outputs(9067) <= a and not b;
    layer2_outputs(9068) <= a xor b;
    layer2_outputs(9069) <= a and b;
    layer2_outputs(9070) <= not a;
    layer2_outputs(9071) <= a and b;
    layer2_outputs(9072) <= b and not a;
    layer2_outputs(9073) <= not b;
    layer2_outputs(9074) <= a and not b;
    layer2_outputs(9075) <= not a;
    layer2_outputs(9076) <= '1';
    layer2_outputs(9077) <= not a or b;
    layer2_outputs(9078) <= a and b;
    layer2_outputs(9079) <= a;
    layer2_outputs(9080) <= b;
    layer2_outputs(9081) <= not (a or b);
    layer2_outputs(9082) <= b;
    layer2_outputs(9083) <= not a or b;
    layer2_outputs(9084) <= not a or b;
    layer2_outputs(9085) <= not (a xor b);
    layer2_outputs(9086) <= not (a xor b);
    layer2_outputs(9087) <= a xor b;
    layer2_outputs(9088) <= a;
    layer2_outputs(9089) <= b and not a;
    layer2_outputs(9090) <= not (a or b);
    layer2_outputs(9091) <= not (a and b);
    layer2_outputs(9092) <= not (a or b);
    layer2_outputs(9093) <= b;
    layer2_outputs(9094) <= not a;
    layer2_outputs(9095) <= b;
    layer2_outputs(9096) <= not (a and b);
    layer2_outputs(9097) <= not b or a;
    layer2_outputs(9098) <= a and not b;
    layer2_outputs(9099) <= not (a or b);
    layer2_outputs(9100) <= b and not a;
    layer2_outputs(9101) <= not a;
    layer2_outputs(9102) <= not b;
    layer2_outputs(9103) <= not (a and b);
    layer2_outputs(9104) <= not (a xor b);
    layer2_outputs(9105) <= a or b;
    layer2_outputs(9106) <= not b or a;
    layer2_outputs(9107) <= a;
    layer2_outputs(9108) <= not a;
    layer2_outputs(9109) <= not (a xor b);
    layer2_outputs(9110) <= a xor b;
    layer2_outputs(9111) <= not a;
    layer2_outputs(9112) <= not b;
    layer2_outputs(9113) <= a;
    layer2_outputs(9114) <= a and not b;
    layer2_outputs(9115) <= not a;
    layer2_outputs(9116) <= a and b;
    layer2_outputs(9117) <= a;
    layer2_outputs(9118) <= a;
    layer2_outputs(9119) <= b;
    layer2_outputs(9120) <= not (a or b);
    layer2_outputs(9121) <= not (a xor b);
    layer2_outputs(9122) <= not a;
    layer2_outputs(9123) <= a or b;
    layer2_outputs(9124) <= not (a and b);
    layer2_outputs(9125) <= a xor b;
    layer2_outputs(9126) <= not a or b;
    layer2_outputs(9127) <= not (a xor b);
    layer2_outputs(9128) <= not (a xor b);
    layer2_outputs(9129) <= b;
    layer2_outputs(9130) <= not b;
    layer2_outputs(9131) <= b and not a;
    layer2_outputs(9132) <= not a;
    layer2_outputs(9133) <= not b;
    layer2_outputs(9134) <= a and b;
    layer2_outputs(9135) <= not b;
    layer2_outputs(9136) <= b;
    layer2_outputs(9137) <= b;
    layer2_outputs(9138) <= a;
    layer2_outputs(9139) <= b;
    layer2_outputs(9140) <= a and b;
    layer2_outputs(9141) <= a;
    layer2_outputs(9142) <= b and not a;
    layer2_outputs(9143) <= a;
    layer2_outputs(9144) <= not a or b;
    layer2_outputs(9145) <= not b or a;
    layer2_outputs(9146) <= not b or a;
    layer2_outputs(9147) <= not (a xor b);
    layer2_outputs(9148) <= b;
    layer2_outputs(9149) <= a and b;
    layer2_outputs(9150) <= a;
    layer2_outputs(9151) <= not a;
    layer2_outputs(9152) <= b and not a;
    layer2_outputs(9153) <= a;
    layer2_outputs(9154) <= not (a xor b);
    layer2_outputs(9155) <= a xor b;
    layer2_outputs(9156) <= a;
    layer2_outputs(9157) <= not a;
    layer2_outputs(9158) <= not a;
    layer2_outputs(9159) <= a xor b;
    layer2_outputs(9160) <= b;
    layer2_outputs(9161) <= not (a xor b);
    layer2_outputs(9162) <= not b;
    layer2_outputs(9163) <= not a or b;
    layer2_outputs(9164) <= not a;
    layer2_outputs(9165) <= not b;
    layer2_outputs(9166) <= not (a and b);
    layer2_outputs(9167) <= not b or a;
    layer2_outputs(9168) <= not (a and b);
    layer2_outputs(9169) <= not b;
    layer2_outputs(9170) <= a;
    layer2_outputs(9171) <= a;
    layer2_outputs(9172) <= not (a xor b);
    layer2_outputs(9173) <= not (a or b);
    layer2_outputs(9174) <= not a;
    layer2_outputs(9175) <= not b;
    layer2_outputs(9176) <= not (a xor b);
    layer2_outputs(9177) <= not (a and b);
    layer2_outputs(9178) <= a xor b;
    layer2_outputs(9179) <= not b or a;
    layer2_outputs(9180) <= not (a or b);
    layer2_outputs(9181) <= not b;
    layer2_outputs(9182) <= a and not b;
    layer2_outputs(9183) <= not a;
    layer2_outputs(9184) <= not a or b;
    layer2_outputs(9185) <= a and b;
    layer2_outputs(9186) <= not b or a;
    layer2_outputs(9187) <= b;
    layer2_outputs(9188) <= not (a xor b);
    layer2_outputs(9189) <= b;
    layer2_outputs(9190) <= not b or a;
    layer2_outputs(9191) <= not a or b;
    layer2_outputs(9192) <= a and b;
    layer2_outputs(9193) <= not (a xor b);
    layer2_outputs(9194) <= not b;
    layer2_outputs(9195) <= b;
    layer2_outputs(9196) <= not a;
    layer2_outputs(9197) <= not (a and b);
    layer2_outputs(9198) <= a;
    layer2_outputs(9199) <= a xor b;
    layer2_outputs(9200) <= b and not a;
    layer2_outputs(9201) <= not b or a;
    layer2_outputs(9202) <= not (a xor b);
    layer2_outputs(9203) <= not b or a;
    layer2_outputs(9204) <= a and not b;
    layer2_outputs(9205) <= not a;
    layer2_outputs(9206) <= not a;
    layer2_outputs(9207) <= not (a or b);
    layer2_outputs(9208) <= not b;
    layer2_outputs(9209) <= not a;
    layer2_outputs(9210) <= not b;
    layer2_outputs(9211) <= b and not a;
    layer2_outputs(9212) <= not b;
    layer2_outputs(9213) <= not b;
    layer2_outputs(9214) <= a and not b;
    layer2_outputs(9215) <= not (a or b);
    layer2_outputs(9216) <= not (a or b);
    layer2_outputs(9217) <= a;
    layer2_outputs(9218) <= not b or a;
    layer2_outputs(9219) <= b and not a;
    layer2_outputs(9220) <= not (a xor b);
    layer2_outputs(9221) <= not a;
    layer2_outputs(9222) <= b;
    layer2_outputs(9223) <= not b;
    layer2_outputs(9224) <= not b;
    layer2_outputs(9225) <= b;
    layer2_outputs(9226) <= not (a xor b);
    layer2_outputs(9227) <= not (a xor b);
    layer2_outputs(9228) <= not a;
    layer2_outputs(9229) <= not b;
    layer2_outputs(9230) <= not (a and b);
    layer2_outputs(9231) <= b;
    layer2_outputs(9232) <= not a;
    layer2_outputs(9233) <= not (a xor b);
    layer2_outputs(9234) <= b;
    layer2_outputs(9235) <= not b or a;
    layer2_outputs(9236) <= not a;
    layer2_outputs(9237) <= a;
    layer2_outputs(9238) <= a and not b;
    layer2_outputs(9239) <= not (a and b);
    layer2_outputs(9240) <= b;
    layer2_outputs(9241) <= a and not b;
    layer2_outputs(9242) <= a and not b;
    layer2_outputs(9243) <= not b;
    layer2_outputs(9244) <= a;
    layer2_outputs(9245) <= not b;
    layer2_outputs(9246) <= not a;
    layer2_outputs(9247) <= a or b;
    layer2_outputs(9248) <= a;
    layer2_outputs(9249) <= a or b;
    layer2_outputs(9250) <= a;
    layer2_outputs(9251) <= a and not b;
    layer2_outputs(9252) <= a and b;
    layer2_outputs(9253) <= a and b;
    layer2_outputs(9254) <= not a or b;
    layer2_outputs(9255) <= a and b;
    layer2_outputs(9256) <= '1';
    layer2_outputs(9257) <= a and not b;
    layer2_outputs(9258) <= not b;
    layer2_outputs(9259) <= not b;
    layer2_outputs(9260) <= a and not b;
    layer2_outputs(9261) <= not (a xor b);
    layer2_outputs(9262) <= a and not b;
    layer2_outputs(9263) <= not (a and b);
    layer2_outputs(9264) <= a and b;
    layer2_outputs(9265) <= not b or a;
    layer2_outputs(9266) <= not b or a;
    layer2_outputs(9267) <= b;
    layer2_outputs(9268) <= a and b;
    layer2_outputs(9269) <= not (a or b);
    layer2_outputs(9270) <= a xor b;
    layer2_outputs(9271) <= a xor b;
    layer2_outputs(9272) <= not (a xor b);
    layer2_outputs(9273) <= not b;
    layer2_outputs(9274) <= not b;
    layer2_outputs(9275) <= not b;
    layer2_outputs(9276) <= not a or b;
    layer2_outputs(9277) <= a and not b;
    layer2_outputs(9278) <= not a;
    layer2_outputs(9279) <= not (a or b);
    layer2_outputs(9280) <= not b;
    layer2_outputs(9281) <= a;
    layer2_outputs(9282) <= not a;
    layer2_outputs(9283) <= b;
    layer2_outputs(9284) <= a and b;
    layer2_outputs(9285) <= b;
    layer2_outputs(9286) <= b and not a;
    layer2_outputs(9287) <= a;
    layer2_outputs(9288) <= a and b;
    layer2_outputs(9289) <= a or b;
    layer2_outputs(9290) <= not (a or b);
    layer2_outputs(9291) <= a and not b;
    layer2_outputs(9292) <= a and b;
    layer2_outputs(9293) <= not b;
    layer2_outputs(9294) <= not (a and b);
    layer2_outputs(9295) <= not (a or b);
    layer2_outputs(9296) <= b and not a;
    layer2_outputs(9297) <= not b or a;
    layer2_outputs(9298) <= a or b;
    layer2_outputs(9299) <= not b;
    layer2_outputs(9300) <= b and not a;
    layer2_outputs(9301) <= not a or b;
    layer2_outputs(9302) <= not (a or b);
    layer2_outputs(9303) <= a;
    layer2_outputs(9304) <= a and not b;
    layer2_outputs(9305) <= '1';
    layer2_outputs(9306) <= a and not b;
    layer2_outputs(9307) <= not b;
    layer2_outputs(9308) <= a and not b;
    layer2_outputs(9309) <= b;
    layer2_outputs(9310) <= not b;
    layer2_outputs(9311) <= not a or b;
    layer2_outputs(9312) <= not b;
    layer2_outputs(9313) <= a;
    layer2_outputs(9314) <= a xor b;
    layer2_outputs(9315) <= not (a and b);
    layer2_outputs(9316) <= a and not b;
    layer2_outputs(9317) <= not a;
    layer2_outputs(9318) <= a and b;
    layer2_outputs(9319) <= a or b;
    layer2_outputs(9320) <= a or b;
    layer2_outputs(9321) <= not b or a;
    layer2_outputs(9322) <= b and not a;
    layer2_outputs(9323) <= not b;
    layer2_outputs(9324) <= not b or a;
    layer2_outputs(9325) <= a;
    layer2_outputs(9326) <= b;
    layer2_outputs(9327) <= not b or a;
    layer2_outputs(9328) <= not b;
    layer2_outputs(9329) <= not b;
    layer2_outputs(9330) <= not (a xor b);
    layer2_outputs(9331) <= not (a and b);
    layer2_outputs(9332) <= a;
    layer2_outputs(9333) <= not b;
    layer2_outputs(9334) <= not (a xor b);
    layer2_outputs(9335) <= a and not b;
    layer2_outputs(9336) <= a xor b;
    layer2_outputs(9337) <= not b;
    layer2_outputs(9338) <= not (a and b);
    layer2_outputs(9339) <= a and not b;
    layer2_outputs(9340) <= not b or a;
    layer2_outputs(9341) <= a;
    layer2_outputs(9342) <= a;
    layer2_outputs(9343) <= not (a and b);
    layer2_outputs(9344) <= not b;
    layer2_outputs(9345) <= a and b;
    layer2_outputs(9346) <= not (a xor b);
    layer2_outputs(9347) <= not (a xor b);
    layer2_outputs(9348) <= b and not a;
    layer2_outputs(9349) <= b;
    layer2_outputs(9350) <= not a;
    layer2_outputs(9351) <= a xor b;
    layer2_outputs(9352) <= not (a and b);
    layer2_outputs(9353) <= a and b;
    layer2_outputs(9354) <= not b;
    layer2_outputs(9355) <= '1';
    layer2_outputs(9356) <= not a;
    layer2_outputs(9357) <= a;
    layer2_outputs(9358) <= b and not a;
    layer2_outputs(9359) <= b;
    layer2_outputs(9360) <= a;
    layer2_outputs(9361) <= not a or b;
    layer2_outputs(9362) <= not a;
    layer2_outputs(9363) <= not (a xor b);
    layer2_outputs(9364) <= not b or a;
    layer2_outputs(9365) <= not b;
    layer2_outputs(9366) <= a xor b;
    layer2_outputs(9367) <= not (a or b);
    layer2_outputs(9368) <= not a;
    layer2_outputs(9369) <= not b or a;
    layer2_outputs(9370) <= not a or b;
    layer2_outputs(9371) <= not b;
    layer2_outputs(9372) <= not (a or b);
    layer2_outputs(9373) <= not b or a;
    layer2_outputs(9374) <= a and b;
    layer2_outputs(9375) <= not a;
    layer2_outputs(9376) <= a and b;
    layer2_outputs(9377) <= not b;
    layer2_outputs(9378) <= not (a xor b);
    layer2_outputs(9379) <= a;
    layer2_outputs(9380) <= not b;
    layer2_outputs(9381) <= not (a and b);
    layer2_outputs(9382) <= a;
    layer2_outputs(9383) <= not (a and b);
    layer2_outputs(9384) <= a and b;
    layer2_outputs(9385) <= not (a xor b);
    layer2_outputs(9386) <= not a;
    layer2_outputs(9387) <= not a;
    layer2_outputs(9388) <= not a;
    layer2_outputs(9389) <= not (a and b);
    layer2_outputs(9390) <= not (a xor b);
    layer2_outputs(9391) <= not a;
    layer2_outputs(9392) <= a;
    layer2_outputs(9393) <= a;
    layer2_outputs(9394) <= not (a or b);
    layer2_outputs(9395) <= not a or b;
    layer2_outputs(9396) <= b;
    layer2_outputs(9397) <= b and not a;
    layer2_outputs(9398) <= a and not b;
    layer2_outputs(9399) <= not b;
    layer2_outputs(9400) <= b;
    layer2_outputs(9401) <= not a or b;
    layer2_outputs(9402) <= a;
    layer2_outputs(9403) <= a or b;
    layer2_outputs(9404) <= b;
    layer2_outputs(9405) <= a and b;
    layer2_outputs(9406) <= b and not a;
    layer2_outputs(9407) <= a or b;
    layer2_outputs(9408) <= a or b;
    layer2_outputs(9409) <= b;
    layer2_outputs(9410) <= b;
    layer2_outputs(9411) <= not (a xor b);
    layer2_outputs(9412) <= a or b;
    layer2_outputs(9413) <= a xor b;
    layer2_outputs(9414) <= a and b;
    layer2_outputs(9415) <= a;
    layer2_outputs(9416) <= b;
    layer2_outputs(9417) <= a and not b;
    layer2_outputs(9418) <= not b;
    layer2_outputs(9419) <= not b;
    layer2_outputs(9420) <= a xor b;
    layer2_outputs(9421) <= a and not b;
    layer2_outputs(9422) <= not a;
    layer2_outputs(9423) <= b;
    layer2_outputs(9424) <= not (a xor b);
    layer2_outputs(9425) <= not b or a;
    layer2_outputs(9426) <= a or b;
    layer2_outputs(9427) <= not a or b;
    layer2_outputs(9428) <= a or b;
    layer2_outputs(9429) <= not b;
    layer2_outputs(9430) <= not a;
    layer2_outputs(9431) <= a xor b;
    layer2_outputs(9432) <= a;
    layer2_outputs(9433) <= not a or b;
    layer2_outputs(9434) <= a and not b;
    layer2_outputs(9435) <= a;
    layer2_outputs(9436) <= not b;
    layer2_outputs(9437) <= not b or a;
    layer2_outputs(9438) <= a and b;
    layer2_outputs(9439) <= not (a xor b);
    layer2_outputs(9440) <= '1';
    layer2_outputs(9441) <= not a;
    layer2_outputs(9442) <= not b or a;
    layer2_outputs(9443) <= a;
    layer2_outputs(9444) <= a and b;
    layer2_outputs(9445) <= a xor b;
    layer2_outputs(9446) <= not b or a;
    layer2_outputs(9447) <= not b or a;
    layer2_outputs(9448) <= not a;
    layer2_outputs(9449) <= a xor b;
    layer2_outputs(9450) <= b;
    layer2_outputs(9451) <= a and not b;
    layer2_outputs(9452) <= not b;
    layer2_outputs(9453) <= a and not b;
    layer2_outputs(9454) <= not (a or b);
    layer2_outputs(9455) <= not a;
    layer2_outputs(9456) <= not b;
    layer2_outputs(9457) <= a;
    layer2_outputs(9458) <= not (a or b);
    layer2_outputs(9459) <= not a or b;
    layer2_outputs(9460) <= not a;
    layer2_outputs(9461) <= not b or a;
    layer2_outputs(9462) <= a and not b;
    layer2_outputs(9463) <= a and b;
    layer2_outputs(9464) <= not (a xor b);
    layer2_outputs(9465) <= b and not a;
    layer2_outputs(9466) <= a and not b;
    layer2_outputs(9467) <= not b;
    layer2_outputs(9468) <= a;
    layer2_outputs(9469) <= a or b;
    layer2_outputs(9470) <= a xor b;
    layer2_outputs(9471) <= a;
    layer2_outputs(9472) <= a;
    layer2_outputs(9473) <= a;
    layer2_outputs(9474) <= b;
    layer2_outputs(9475) <= a or b;
    layer2_outputs(9476) <= a or b;
    layer2_outputs(9477) <= b;
    layer2_outputs(9478) <= a and b;
    layer2_outputs(9479) <= b;
    layer2_outputs(9480) <= not a;
    layer2_outputs(9481) <= a;
    layer2_outputs(9482) <= not (a or b);
    layer2_outputs(9483) <= not (a or b);
    layer2_outputs(9484) <= not a;
    layer2_outputs(9485) <= b and not a;
    layer2_outputs(9486) <= not a;
    layer2_outputs(9487) <= a and not b;
    layer2_outputs(9488) <= not a or b;
    layer2_outputs(9489) <= not a;
    layer2_outputs(9490) <= not (a or b);
    layer2_outputs(9491) <= b;
    layer2_outputs(9492) <= not a;
    layer2_outputs(9493) <= a and b;
    layer2_outputs(9494) <= a or b;
    layer2_outputs(9495) <= a or b;
    layer2_outputs(9496) <= not b;
    layer2_outputs(9497) <= not (a and b);
    layer2_outputs(9498) <= a or b;
    layer2_outputs(9499) <= b and not a;
    layer2_outputs(9500) <= not (a or b);
    layer2_outputs(9501) <= not (a or b);
    layer2_outputs(9502) <= a;
    layer2_outputs(9503) <= not a;
    layer2_outputs(9504) <= not (a xor b);
    layer2_outputs(9505) <= not b;
    layer2_outputs(9506) <= not b;
    layer2_outputs(9507) <= not a;
    layer2_outputs(9508) <= a;
    layer2_outputs(9509) <= a xor b;
    layer2_outputs(9510) <= b and not a;
    layer2_outputs(9511) <= not a or b;
    layer2_outputs(9512) <= not (a and b);
    layer2_outputs(9513) <= not (a or b);
    layer2_outputs(9514) <= not (a and b);
    layer2_outputs(9515) <= a;
    layer2_outputs(9516) <= not (a and b);
    layer2_outputs(9517) <= b;
    layer2_outputs(9518) <= not b or a;
    layer2_outputs(9519) <= not a or b;
    layer2_outputs(9520) <= a xor b;
    layer2_outputs(9521) <= not (a xor b);
    layer2_outputs(9522) <= a or b;
    layer2_outputs(9523) <= a;
    layer2_outputs(9524) <= a;
    layer2_outputs(9525) <= a or b;
    layer2_outputs(9526) <= not (a xor b);
    layer2_outputs(9527) <= a or b;
    layer2_outputs(9528) <= not b;
    layer2_outputs(9529) <= a;
    layer2_outputs(9530) <= not b or a;
    layer2_outputs(9531) <= a and b;
    layer2_outputs(9532) <= a and b;
    layer2_outputs(9533) <= not (a or b);
    layer2_outputs(9534) <= not b or a;
    layer2_outputs(9535) <= a xor b;
    layer2_outputs(9536) <= a and not b;
    layer2_outputs(9537) <= a and not b;
    layer2_outputs(9538) <= a;
    layer2_outputs(9539) <= not a;
    layer2_outputs(9540) <= not a or b;
    layer2_outputs(9541) <= a;
    layer2_outputs(9542) <= a;
    layer2_outputs(9543) <= b and not a;
    layer2_outputs(9544) <= not (a or b);
    layer2_outputs(9545) <= b and not a;
    layer2_outputs(9546) <= not (a and b);
    layer2_outputs(9547) <= a;
    layer2_outputs(9548) <= not b;
    layer2_outputs(9549) <= not (a xor b);
    layer2_outputs(9550) <= not (a xor b);
    layer2_outputs(9551) <= a xor b;
    layer2_outputs(9552) <= a;
    layer2_outputs(9553) <= not b or a;
    layer2_outputs(9554) <= a xor b;
    layer2_outputs(9555) <= not a or b;
    layer2_outputs(9556) <= not a;
    layer2_outputs(9557) <= not a;
    layer2_outputs(9558) <= b;
    layer2_outputs(9559) <= a and b;
    layer2_outputs(9560) <= not a or b;
    layer2_outputs(9561) <= '0';
    layer2_outputs(9562) <= a;
    layer2_outputs(9563) <= a and not b;
    layer2_outputs(9564) <= not a;
    layer2_outputs(9565) <= not b;
    layer2_outputs(9566) <= b;
    layer2_outputs(9567) <= not (a xor b);
    layer2_outputs(9568) <= not b;
    layer2_outputs(9569) <= not a;
    layer2_outputs(9570) <= a and b;
    layer2_outputs(9571) <= b and not a;
    layer2_outputs(9572) <= not a;
    layer2_outputs(9573) <= b and not a;
    layer2_outputs(9574) <= not (a xor b);
    layer2_outputs(9575) <= b;
    layer2_outputs(9576) <= not (a and b);
    layer2_outputs(9577) <= not b or a;
    layer2_outputs(9578) <= not (a or b);
    layer2_outputs(9579) <= b;
    layer2_outputs(9580) <= not b;
    layer2_outputs(9581) <= a;
    layer2_outputs(9582) <= not (a xor b);
    layer2_outputs(9583) <= not b;
    layer2_outputs(9584) <= not (a xor b);
    layer2_outputs(9585) <= not b;
    layer2_outputs(9586) <= not b;
    layer2_outputs(9587) <= a and not b;
    layer2_outputs(9588) <= b and not a;
    layer2_outputs(9589) <= a xor b;
    layer2_outputs(9590) <= a and not b;
    layer2_outputs(9591) <= a xor b;
    layer2_outputs(9592) <= not b or a;
    layer2_outputs(9593) <= a xor b;
    layer2_outputs(9594) <= b;
    layer2_outputs(9595) <= a and not b;
    layer2_outputs(9596) <= not a;
    layer2_outputs(9597) <= a xor b;
    layer2_outputs(9598) <= b;
    layer2_outputs(9599) <= not (a and b);
    layer2_outputs(9600) <= not b;
    layer2_outputs(9601) <= not (a and b);
    layer2_outputs(9602) <= not (a or b);
    layer2_outputs(9603) <= a and b;
    layer2_outputs(9604) <= not b or a;
    layer2_outputs(9605) <= a;
    layer2_outputs(9606) <= not b;
    layer2_outputs(9607) <= a xor b;
    layer2_outputs(9608) <= a or b;
    layer2_outputs(9609) <= a or b;
    layer2_outputs(9610) <= b and not a;
    layer2_outputs(9611) <= a and b;
    layer2_outputs(9612) <= not (a or b);
    layer2_outputs(9613) <= b;
    layer2_outputs(9614) <= a;
    layer2_outputs(9615) <= not b;
    layer2_outputs(9616) <= b;
    layer2_outputs(9617) <= b;
    layer2_outputs(9618) <= not a or b;
    layer2_outputs(9619) <= a or b;
    layer2_outputs(9620) <= not a or b;
    layer2_outputs(9621) <= not b;
    layer2_outputs(9622) <= not a;
    layer2_outputs(9623) <= not b;
    layer2_outputs(9624) <= a or b;
    layer2_outputs(9625) <= not b;
    layer2_outputs(9626) <= a xor b;
    layer2_outputs(9627) <= a xor b;
    layer2_outputs(9628) <= not (a and b);
    layer2_outputs(9629) <= not b or a;
    layer2_outputs(9630) <= not a or b;
    layer2_outputs(9631) <= not a;
    layer2_outputs(9632) <= not a;
    layer2_outputs(9633) <= a xor b;
    layer2_outputs(9634) <= a and not b;
    layer2_outputs(9635) <= not a;
    layer2_outputs(9636) <= a;
    layer2_outputs(9637) <= b;
    layer2_outputs(9638) <= not (a xor b);
    layer2_outputs(9639) <= b and not a;
    layer2_outputs(9640) <= not (a or b);
    layer2_outputs(9641) <= a xor b;
    layer2_outputs(9642) <= not (a or b);
    layer2_outputs(9643) <= a and not b;
    layer2_outputs(9644) <= a;
    layer2_outputs(9645) <= not b or a;
    layer2_outputs(9646) <= b and not a;
    layer2_outputs(9647) <= not (a or b);
    layer2_outputs(9648) <= not b or a;
    layer2_outputs(9649) <= a xor b;
    layer2_outputs(9650) <= a;
    layer2_outputs(9651) <= b and not a;
    layer2_outputs(9652) <= '0';
    layer2_outputs(9653) <= b;
    layer2_outputs(9654) <= a xor b;
    layer2_outputs(9655) <= not (a and b);
    layer2_outputs(9656) <= not (a or b);
    layer2_outputs(9657) <= not a or b;
    layer2_outputs(9658) <= not a;
    layer2_outputs(9659) <= b;
    layer2_outputs(9660) <= not (a xor b);
    layer2_outputs(9661) <= a;
    layer2_outputs(9662) <= a and b;
    layer2_outputs(9663) <= not (a or b);
    layer2_outputs(9664) <= a xor b;
    layer2_outputs(9665) <= not b;
    layer2_outputs(9666) <= a;
    layer2_outputs(9667) <= not a;
    layer2_outputs(9668) <= b and not a;
    layer2_outputs(9669) <= a xor b;
    layer2_outputs(9670) <= a or b;
    layer2_outputs(9671) <= b;
    layer2_outputs(9672) <= not b;
    layer2_outputs(9673) <= a xor b;
    layer2_outputs(9674) <= a;
    layer2_outputs(9675) <= a xor b;
    layer2_outputs(9676) <= not (a and b);
    layer2_outputs(9677) <= not b;
    layer2_outputs(9678) <= a or b;
    layer2_outputs(9679) <= a xor b;
    layer2_outputs(9680) <= a and b;
    layer2_outputs(9681) <= not a or b;
    layer2_outputs(9682) <= b;
    layer2_outputs(9683) <= not (a xor b);
    layer2_outputs(9684) <= not a or b;
    layer2_outputs(9685) <= a or b;
    layer2_outputs(9686) <= b and not a;
    layer2_outputs(9687) <= not (a or b);
    layer2_outputs(9688) <= not a or b;
    layer2_outputs(9689) <= a and not b;
    layer2_outputs(9690) <= b and not a;
    layer2_outputs(9691) <= a;
    layer2_outputs(9692) <= not (a and b);
    layer2_outputs(9693) <= a or b;
    layer2_outputs(9694) <= not b;
    layer2_outputs(9695) <= not (a xor b);
    layer2_outputs(9696) <= not (a or b);
    layer2_outputs(9697) <= a xor b;
    layer2_outputs(9698) <= not (a xor b);
    layer2_outputs(9699) <= not (a or b);
    layer2_outputs(9700) <= a or b;
    layer2_outputs(9701) <= not a or b;
    layer2_outputs(9702) <= not a;
    layer2_outputs(9703) <= not (a xor b);
    layer2_outputs(9704) <= not b or a;
    layer2_outputs(9705) <= a;
    layer2_outputs(9706) <= a xor b;
    layer2_outputs(9707) <= not a;
    layer2_outputs(9708) <= a;
    layer2_outputs(9709) <= b and not a;
    layer2_outputs(9710) <= not b;
    layer2_outputs(9711) <= not (a and b);
    layer2_outputs(9712) <= b;
    layer2_outputs(9713) <= not b;
    layer2_outputs(9714) <= not a or b;
    layer2_outputs(9715) <= not a;
    layer2_outputs(9716) <= not (a or b);
    layer2_outputs(9717) <= not a;
    layer2_outputs(9718) <= a and b;
    layer2_outputs(9719) <= b;
    layer2_outputs(9720) <= not a;
    layer2_outputs(9721) <= b;
    layer2_outputs(9722) <= b;
    layer2_outputs(9723) <= not b or a;
    layer2_outputs(9724) <= not b;
    layer2_outputs(9725) <= not (a xor b);
    layer2_outputs(9726) <= not a or b;
    layer2_outputs(9727) <= a and b;
    layer2_outputs(9728) <= not b or a;
    layer2_outputs(9729) <= a or b;
    layer2_outputs(9730) <= not a;
    layer2_outputs(9731) <= not (a or b);
    layer2_outputs(9732) <= not a;
    layer2_outputs(9733) <= a or b;
    layer2_outputs(9734) <= b;
    layer2_outputs(9735) <= a and not b;
    layer2_outputs(9736) <= not a;
    layer2_outputs(9737) <= not b;
    layer2_outputs(9738) <= not (a xor b);
    layer2_outputs(9739) <= b and not a;
    layer2_outputs(9740) <= not (a or b);
    layer2_outputs(9741) <= not (a xor b);
    layer2_outputs(9742) <= not b or a;
    layer2_outputs(9743) <= a;
    layer2_outputs(9744) <= a and b;
    layer2_outputs(9745) <= not (a and b);
    layer2_outputs(9746) <= a xor b;
    layer2_outputs(9747) <= a;
    layer2_outputs(9748) <= not (a and b);
    layer2_outputs(9749) <= a and b;
    layer2_outputs(9750) <= a;
    layer2_outputs(9751) <= not (a or b);
    layer2_outputs(9752) <= b;
    layer2_outputs(9753) <= a xor b;
    layer2_outputs(9754) <= a and b;
    layer2_outputs(9755) <= a;
    layer2_outputs(9756) <= not (a and b);
    layer2_outputs(9757) <= a xor b;
    layer2_outputs(9758) <= a;
    layer2_outputs(9759) <= b;
    layer2_outputs(9760) <= not b;
    layer2_outputs(9761) <= a and b;
    layer2_outputs(9762) <= not a;
    layer2_outputs(9763) <= b;
    layer2_outputs(9764) <= a and b;
    layer2_outputs(9765) <= a;
    layer2_outputs(9766) <= not (a or b);
    layer2_outputs(9767) <= not (a or b);
    layer2_outputs(9768) <= not a;
    layer2_outputs(9769) <= not b;
    layer2_outputs(9770) <= not b;
    layer2_outputs(9771) <= a;
    layer2_outputs(9772) <= a and not b;
    layer2_outputs(9773) <= not (a xor b);
    layer2_outputs(9774) <= not b;
    layer2_outputs(9775) <= not (a or b);
    layer2_outputs(9776) <= a;
    layer2_outputs(9777) <= a;
    layer2_outputs(9778) <= not (a xor b);
    layer2_outputs(9779) <= a;
    layer2_outputs(9780) <= b;
    layer2_outputs(9781) <= not (a and b);
    layer2_outputs(9782) <= a and not b;
    layer2_outputs(9783) <= a;
    layer2_outputs(9784) <= a;
    layer2_outputs(9785) <= a;
    layer2_outputs(9786) <= a and b;
    layer2_outputs(9787) <= a;
    layer2_outputs(9788) <= a and not b;
    layer2_outputs(9789) <= not a or b;
    layer2_outputs(9790) <= a;
    layer2_outputs(9791) <= not a or b;
    layer2_outputs(9792) <= b and not a;
    layer2_outputs(9793) <= a;
    layer2_outputs(9794) <= b and not a;
    layer2_outputs(9795) <= a;
    layer2_outputs(9796) <= a and b;
    layer2_outputs(9797) <= a and b;
    layer2_outputs(9798) <= a xor b;
    layer2_outputs(9799) <= not (a xor b);
    layer2_outputs(9800) <= not b or a;
    layer2_outputs(9801) <= b;
    layer2_outputs(9802) <= a xor b;
    layer2_outputs(9803) <= a or b;
    layer2_outputs(9804) <= not (a xor b);
    layer2_outputs(9805) <= a xor b;
    layer2_outputs(9806) <= b and not a;
    layer2_outputs(9807) <= a or b;
    layer2_outputs(9808) <= a or b;
    layer2_outputs(9809) <= a or b;
    layer2_outputs(9810) <= a and b;
    layer2_outputs(9811) <= b;
    layer2_outputs(9812) <= a and b;
    layer2_outputs(9813) <= not a or b;
    layer2_outputs(9814) <= not b or a;
    layer2_outputs(9815) <= not (a and b);
    layer2_outputs(9816) <= a and b;
    layer2_outputs(9817) <= not b or a;
    layer2_outputs(9818) <= a and b;
    layer2_outputs(9819) <= b;
    layer2_outputs(9820) <= not a;
    layer2_outputs(9821) <= a;
    layer2_outputs(9822) <= a or b;
    layer2_outputs(9823) <= b;
    layer2_outputs(9824) <= b and not a;
    layer2_outputs(9825) <= a and not b;
    layer2_outputs(9826) <= not a;
    layer2_outputs(9827) <= not b;
    layer2_outputs(9828) <= not (a xor b);
    layer2_outputs(9829) <= b and not a;
    layer2_outputs(9830) <= a and not b;
    layer2_outputs(9831) <= not a;
    layer2_outputs(9832) <= not (a or b);
    layer2_outputs(9833) <= a;
    layer2_outputs(9834) <= a and not b;
    layer2_outputs(9835) <= not a;
    layer2_outputs(9836) <= not (a xor b);
    layer2_outputs(9837) <= a xor b;
    layer2_outputs(9838) <= a;
    layer2_outputs(9839) <= a xor b;
    layer2_outputs(9840) <= a or b;
    layer2_outputs(9841) <= not (a and b);
    layer2_outputs(9842) <= a;
    layer2_outputs(9843) <= a xor b;
    layer2_outputs(9844) <= a;
    layer2_outputs(9845) <= b;
    layer2_outputs(9846) <= not a;
    layer2_outputs(9847) <= a and b;
    layer2_outputs(9848) <= not (a xor b);
    layer2_outputs(9849) <= a;
    layer2_outputs(9850) <= not b or a;
    layer2_outputs(9851) <= not (a and b);
    layer2_outputs(9852) <= not b;
    layer2_outputs(9853) <= a;
    layer2_outputs(9854) <= not b;
    layer2_outputs(9855) <= a or b;
    layer2_outputs(9856) <= b;
    layer2_outputs(9857) <= a;
    layer2_outputs(9858) <= a;
    layer2_outputs(9859) <= b and not a;
    layer2_outputs(9860) <= a;
    layer2_outputs(9861) <= not (a and b);
    layer2_outputs(9862) <= b;
    layer2_outputs(9863) <= a;
    layer2_outputs(9864) <= not (a or b);
    layer2_outputs(9865) <= b;
    layer2_outputs(9866) <= not a;
    layer2_outputs(9867) <= not b or a;
    layer2_outputs(9868) <= not b or a;
    layer2_outputs(9869) <= b and not a;
    layer2_outputs(9870) <= not (a and b);
    layer2_outputs(9871) <= not a;
    layer2_outputs(9872) <= a;
    layer2_outputs(9873) <= a;
    layer2_outputs(9874) <= a xor b;
    layer2_outputs(9875) <= b;
    layer2_outputs(9876) <= a and not b;
    layer2_outputs(9877) <= not (a xor b);
    layer2_outputs(9878) <= not b or a;
    layer2_outputs(9879) <= not (a xor b);
    layer2_outputs(9880) <= a or b;
    layer2_outputs(9881) <= not a;
    layer2_outputs(9882) <= a or b;
    layer2_outputs(9883) <= not (a or b);
    layer2_outputs(9884) <= not (a xor b);
    layer2_outputs(9885) <= b;
    layer2_outputs(9886) <= not (a and b);
    layer2_outputs(9887) <= a or b;
    layer2_outputs(9888) <= b;
    layer2_outputs(9889) <= a or b;
    layer2_outputs(9890) <= not a;
    layer2_outputs(9891) <= a and b;
    layer2_outputs(9892) <= not (a xor b);
    layer2_outputs(9893) <= not a;
    layer2_outputs(9894) <= b;
    layer2_outputs(9895) <= b;
    layer2_outputs(9896) <= a xor b;
    layer2_outputs(9897) <= not a or b;
    layer2_outputs(9898) <= '1';
    layer2_outputs(9899) <= a and not b;
    layer2_outputs(9900) <= not (a or b);
    layer2_outputs(9901) <= a and not b;
    layer2_outputs(9902) <= not a;
    layer2_outputs(9903) <= not a or b;
    layer2_outputs(9904) <= a and b;
    layer2_outputs(9905) <= a xor b;
    layer2_outputs(9906) <= b and not a;
    layer2_outputs(9907) <= b;
    layer2_outputs(9908) <= not b;
    layer2_outputs(9909) <= a;
    layer2_outputs(9910) <= a;
    layer2_outputs(9911) <= not (a xor b);
    layer2_outputs(9912) <= not a or b;
    layer2_outputs(9913) <= not a;
    layer2_outputs(9914) <= not b;
    layer2_outputs(9915) <= a and b;
    layer2_outputs(9916) <= not (a xor b);
    layer2_outputs(9917) <= b;
    layer2_outputs(9918) <= a or b;
    layer2_outputs(9919) <= a;
    layer2_outputs(9920) <= not a or b;
    layer2_outputs(9921) <= not (a xor b);
    layer2_outputs(9922) <= b;
    layer2_outputs(9923) <= not (a and b);
    layer2_outputs(9924) <= a xor b;
    layer2_outputs(9925) <= not a;
    layer2_outputs(9926) <= a;
    layer2_outputs(9927) <= not (a or b);
    layer2_outputs(9928) <= a and not b;
    layer2_outputs(9929) <= a and b;
    layer2_outputs(9930) <= not (a and b);
    layer2_outputs(9931) <= not b;
    layer2_outputs(9932) <= not b;
    layer2_outputs(9933) <= b and not a;
    layer2_outputs(9934) <= a and not b;
    layer2_outputs(9935) <= not a or b;
    layer2_outputs(9936) <= a and b;
    layer2_outputs(9937) <= not (a or b);
    layer2_outputs(9938) <= not (a xor b);
    layer2_outputs(9939) <= a and b;
    layer2_outputs(9940) <= not (a xor b);
    layer2_outputs(9941) <= a and b;
    layer2_outputs(9942) <= not a or b;
    layer2_outputs(9943) <= not (a and b);
    layer2_outputs(9944) <= a and not b;
    layer2_outputs(9945) <= a xor b;
    layer2_outputs(9946) <= not (a xor b);
    layer2_outputs(9947) <= not (a xor b);
    layer2_outputs(9948) <= a xor b;
    layer2_outputs(9949) <= not a or b;
    layer2_outputs(9950) <= not (a or b);
    layer2_outputs(9951) <= a;
    layer2_outputs(9952) <= not a or b;
    layer2_outputs(9953) <= not a;
    layer2_outputs(9954) <= not (a and b);
    layer2_outputs(9955) <= b and not a;
    layer2_outputs(9956) <= not (a or b);
    layer2_outputs(9957) <= b;
    layer2_outputs(9958) <= '0';
    layer2_outputs(9959) <= not a;
    layer2_outputs(9960) <= b;
    layer2_outputs(9961) <= b;
    layer2_outputs(9962) <= not a;
    layer2_outputs(9963) <= not (a xor b);
    layer2_outputs(9964) <= not (a and b);
    layer2_outputs(9965) <= not a;
    layer2_outputs(9966) <= not a or b;
    layer2_outputs(9967) <= not b;
    layer2_outputs(9968) <= b;
    layer2_outputs(9969) <= a xor b;
    layer2_outputs(9970) <= '0';
    layer2_outputs(9971) <= a or b;
    layer2_outputs(9972) <= not b or a;
    layer2_outputs(9973) <= not (a xor b);
    layer2_outputs(9974) <= a and not b;
    layer2_outputs(9975) <= a xor b;
    layer2_outputs(9976) <= not a or b;
    layer2_outputs(9977) <= a and b;
    layer2_outputs(9978) <= a and not b;
    layer2_outputs(9979) <= not (a xor b);
    layer2_outputs(9980) <= not b;
    layer2_outputs(9981) <= a;
    layer2_outputs(9982) <= not (a xor b);
    layer2_outputs(9983) <= a;
    layer2_outputs(9984) <= not (a and b);
    layer2_outputs(9985) <= not (a xor b);
    layer2_outputs(9986) <= a xor b;
    layer2_outputs(9987) <= not a;
    layer2_outputs(9988) <= not (a xor b);
    layer2_outputs(9989) <= not a or b;
    layer2_outputs(9990) <= a;
    layer2_outputs(9991) <= not (a or b);
    layer2_outputs(9992) <= not (a xor b);
    layer2_outputs(9993) <= b;
    layer2_outputs(9994) <= not (a or b);
    layer2_outputs(9995) <= '0';
    layer2_outputs(9996) <= not b;
    layer2_outputs(9997) <= a and not b;
    layer2_outputs(9998) <= not (a xor b);
    layer2_outputs(9999) <= not a or b;
    layer2_outputs(10000) <= a;
    layer2_outputs(10001) <= not (a xor b);
    layer2_outputs(10002) <= a or b;
    layer2_outputs(10003) <= not a or b;
    layer2_outputs(10004) <= b and not a;
    layer2_outputs(10005) <= not a;
    layer2_outputs(10006) <= a or b;
    layer2_outputs(10007) <= a or b;
    layer2_outputs(10008) <= not (a xor b);
    layer2_outputs(10009) <= not (a xor b);
    layer2_outputs(10010) <= not (a xor b);
    layer2_outputs(10011) <= not (a xor b);
    layer2_outputs(10012) <= not a or b;
    layer2_outputs(10013) <= not a or b;
    layer2_outputs(10014) <= not a or b;
    layer2_outputs(10015) <= a and not b;
    layer2_outputs(10016) <= b;
    layer2_outputs(10017) <= not a;
    layer2_outputs(10018) <= not (a or b);
    layer2_outputs(10019) <= '0';
    layer2_outputs(10020) <= not a;
    layer2_outputs(10021) <= a or b;
    layer2_outputs(10022) <= not (a and b);
    layer2_outputs(10023) <= not a;
    layer2_outputs(10024) <= a;
    layer2_outputs(10025) <= b;
    layer2_outputs(10026) <= b;
    layer2_outputs(10027) <= not a;
    layer2_outputs(10028) <= a;
    layer2_outputs(10029) <= a and not b;
    layer2_outputs(10030) <= b;
    layer2_outputs(10031) <= not b;
    layer2_outputs(10032) <= not (a and b);
    layer2_outputs(10033) <= not a or b;
    layer2_outputs(10034) <= not (a xor b);
    layer2_outputs(10035) <= a;
    layer2_outputs(10036) <= b;
    layer2_outputs(10037) <= not (a xor b);
    layer2_outputs(10038) <= a;
    layer2_outputs(10039) <= b and not a;
    layer2_outputs(10040) <= not (a and b);
    layer2_outputs(10041) <= not (a xor b);
    layer2_outputs(10042) <= not a;
    layer2_outputs(10043) <= a xor b;
    layer2_outputs(10044) <= not (a xor b);
    layer2_outputs(10045) <= not b;
    layer2_outputs(10046) <= a;
    layer2_outputs(10047) <= b and not a;
    layer2_outputs(10048) <= a xor b;
    layer2_outputs(10049) <= a;
    layer2_outputs(10050) <= not a;
    layer2_outputs(10051) <= not b or a;
    layer2_outputs(10052) <= not b;
    layer2_outputs(10053) <= a xor b;
    layer2_outputs(10054) <= a;
    layer2_outputs(10055) <= a and not b;
    layer2_outputs(10056) <= a;
    layer2_outputs(10057) <= a and b;
    layer2_outputs(10058) <= not (a and b);
    layer2_outputs(10059) <= a;
    layer2_outputs(10060) <= not (a or b);
    layer2_outputs(10061) <= not a;
    layer2_outputs(10062) <= not a;
    layer2_outputs(10063) <= a or b;
    layer2_outputs(10064) <= not b;
    layer2_outputs(10065) <= not a;
    layer2_outputs(10066) <= not (a and b);
    layer2_outputs(10067) <= b;
    layer2_outputs(10068) <= not b;
    layer2_outputs(10069) <= a;
    layer2_outputs(10070) <= not (a xor b);
    layer2_outputs(10071) <= not b;
    layer2_outputs(10072) <= a xor b;
    layer2_outputs(10073) <= a xor b;
    layer2_outputs(10074) <= not b;
    layer2_outputs(10075) <= not a;
    layer2_outputs(10076) <= b and not a;
    layer2_outputs(10077) <= not (a and b);
    layer2_outputs(10078) <= a xor b;
    layer2_outputs(10079) <= a or b;
    layer2_outputs(10080) <= not b or a;
    layer2_outputs(10081) <= a xor b;
    layer2_outputs(10082) <= not b;
    layer2_outputs(10083) <= b;
    layer2_outputs(10084) <= not b;
    layer2_outputs(10085) <= a;
    layer2_outputs(10086) <= a;
    layer2_outputs(10087) <= a;
    layer2_outputs(10088) <= not a;
    layer2_outputs(10089) <= b and not a;
    layer2_outputs(10090) <= not (a xor b);
    layer2_outputs(10091) <= a and not b;
    layer2_outputs(10092) <= a or b;
    layer2_outputs(10093) <= not (a and b);
    layer2_outputs(10094) <= b and not a;
    layer2_outputs(10095) <= not (a xor b);
    layer2_outputs(10096) <= b;
    layer2_outputs(10097) <= not a or b;
    layer2_outputs(10098) <= not b;
    layer2_outputs(10099) <= not b;
    layer2_outputs(10100) <= not a;
    layer2_outputs(10101) <= not b or a;
    layer2_outputs(10102) <= not (a or b);
    layer2_outputs(10103) <= b and not a;
    layer2_outputs(10104) <= not (a or b);
    layer2_outputs(10105) <= a;
    layer2_outputs(10106) <= not (a xor b);
    layer2_outputs(10107) <= not a;
    layer2_outputs(10108) <= b;
    layer2_outputs(10109) <= b and not a;
    layer2_outputs(10110) <= a xor b;
    layer2_outputs(10111) <= b and not a;
    layer2_outputs(10112) <= not (a and b);
    layer2_outputs(10113) <= not a or b;
    layer2_outputs(10114) <= b and not a;
    layer2_outputs(10115) <= a xor b;
    layer2_outputs(10116) <= not (a xor b);
    layer2_outputs(10117) <= b;
    layer2_outputs(10118) <= not b or a;
    layer2_outputs(10119) <= a xor b;
    layer2_outputs(10120) <= a;
    layer2_outputs(10121) <= b;
    layer2_outputs(10122) <= a;
    layer2_outputs(10123) <= not b;
    layer2_outputs(10124) <= not (a and b);
    layer2_outputs(10125) <= b and not a;
    layer2_outputs(10126) <= a xor b;
    layer2_outputs(10127) <= not a;
    layer2_outputs(10128) <= not b or a;
    layer2_outputs(10129) <= not (a or b);
    layer2_outputs(10130) <= a xor b;
    layer2_outputs(10131) <= not a;
    layer2_outputs(10132) <= not a;
    layer2_outputs(10133) <= a or b;
    layer2_outputs(10134) <= '0';
    layer2_outputs(10135) <= a and b;
    layer2_outputs(10136) <= '0';
    layer2_outputs(10137) <= not (a xor b);
    layer2_outputs(10138) <= b;
    layer2_outputs(10139) <= not a;
    layer2_outputs(10140) <= not (a xor b);
    layer2_outputs(10141) <= a or b;
    layer2_outputs(10142) <= a and not b;
    layer2_outputs(10143) <= not (a xor b);
    layer2_outputs(10144) <= not (a xor b);
    layer2_outputs(10145) <= a and not b;
    layer2_outputs(10146) <= a and not b;
    layer2_outputs(10147) <= not b;
    layer2_outputs(10148) <= a and b;
    layer2_outputs(10149) <= a and not b;
    layer2_outputs(10150) <= not b or a;
    layer2_outputs(10151) <= b;
    layer2_outputs(10152) <= a and b;
    layer2_outputs(10153) <= a xor b;
    layer2_outputs(10154) <= not a or b;
    layer2_outputs(10155) <= not (a and b);
    layer2_outputs(10156) <= b and not a;
    layer2_outputs(10157) <= '0';
    layer2_outputs(10158) <= a;
    layer2_outputs(10159) <= b and not a;
    layer2_outputs(10160) <= b and not a;
    layer2_outputs(10161) <= a and b;
    layer2_outputs(10162) <= b and not a;
    layer2_outputs(10163) <= a xor b;
    layer2_outputs(10164) <= a;
    layer2_outputs(10165) <= a and not b;
    layer2_outputs(10166) <= not a;
    layer2_outputs(10167) <= a;
    layer2_outputs(10168) <= b;
    layer2_outputs(10169) <= b and not a;
    layer2_outputs(10170) <= not (a xor b);
    layer2_outputs(10171) <= not (a xor b);
    layer2_outputs(10172) <= a and b;
    layer2_outputs(10173) <= b and not a;
    layer2_outputs(10174) <= not b;
    layer2_outputs(10175) <= a and b;
    layer2_outputs(10176) <= not a;
    layer2_outputs(10177) <= b and not a;
    layer2_outputs(10178) <= not (a xor b);
    layer2_outputs(10179) <= b;
    layer2_outputs(10180) <= not b or a;
    layer2_outputs(10181) <= not (a or b);
    layer2_outputs(10182) <= not (a xor b);
    layer2_outputs(10183) <= a or b;
    layer2_outputs(10184) <= b and not a;
    layer2_outputs(10185) <= not b or a;
    layer2_outputs(10186) <= not b or a;
    layer2_outputs(10187) <= a;
    layer2_outputs(10188) <= not a;
    layer2_outputs(10189) <= b and not a;
    layer2_outputs(10190) <= not (a xor b);
    layer2_outputs(10191) <= b and not a;
    layer2_outputs(10192) <= a;
    layer2_outputs(10193) <= not (a xor b);
    layer2_outputs(10194) <= not b;
    layer2_outputs(10195) <= a xor b;
    layer2_outputs(10196) <= a and not b;
    layer2_outputs(10197) <= a xor b;
    layer2_outputs(10198) <= a;
    layer2_outputs(10199) <= a and b;
    layer2_outputs(10200) <= a xor b;
    layer2_outputs(10201) <= b;
    layer2_outputs(10202) <= not (a or b);
    layer2_outputs(10203) <= not b or a;
    layer2_outputs(10204) <= not a or b;
    layer2_outputs(10205) <= a;
    layer2_outputs(10206) <= b;
    layer2_outputs(10207) <= not (a and b);
    layer2_outputs(10208) <= b and not a;
    layer2_outputs(10209) <= a or b;
    layer2_outputs(10210) <= a and b;
    layer2_outputs(10211) <= not (a xor b);
    layer2_outputs(10212) <= b;
    layer2_outputs(10213) <= a and b;
    layer2_outputs(10214) <= b and not a;
    layer2_outputs(10215) <= not b;
    layer2_outputs(10216) <= a and b;
    layer2_outputs(10217) <= '1';
    layer2_outputs(10218) <= not (a xor b);
    layer2_outputs(10219) <= not b;
    layer2_outputs(10220) <= not b;
    layer2_outputs(10221) <= not b;
    layer2_outputs(10222) <= not b;
    layer2_outputs(10223) <= not (a xor b);
    layer2_outputs(10224) <= not a;
    layer2_outputs(10225) <= a;
    layer2_outputs(10226) <= b;
    layer2_outputs(10227) <= not b or a;
    layer2_outputs(10228) <= not (a xor b);
    layer2_outputs(10229) <= b;
    layer2_outputs(10230) <= a;
    layer2_outputs(10231) <= not (a or b);
    layer2_outputs(10232) <= a xor b;
    layer2_outputs(10233) <= b and not a;
    layer2_outputs(10234) <= b and not a;
    layer2_outputs(10235) <= not b or a;
    layer2_outputs(10236) <= not a or b;
    layer2_outputs(10237) <= a xor b;
    layer2_outputs(10238) <= a xor b;
    layer2_outputs(10239) <= b;
    outputs(0) <= b;
    outputs(1) <= b;
    outputs(2) <= b and not a;
    outputs(3) <= a xor b;
    outputs(4) <= not a;
    outputs(5) <= b;
    outputs(6) <= not b;
    outputs(7) <= not a or b;
    outputs(8) <= a;
    outputs(9) <= a and not b;
    outputs(10) <= not a;
    outputs(11) <= a;
    outputs(12) <= a xor b;
    outputs(13) <= not a;
    outputs(14) <= not a or b;
    outputs(15) <= a;
    outputs(16) <= not a;
    outputs(17) <= not (a xor b);
    outputs(18) <= not (a or b);
    outputs(19) <= not (a or b);
    outputs(20) <= not a;
    outputs(21) <= a and b;
    outputs(22) <= b;
    outputs(23) <= b;
    outputs(24) <= not a;
    outputs(25) <= a and b;
    outputs(26) <= not b;
    outputs(27) <= b;
    outputs(28) <= a xor b;
    outputs(29) <= not b;
    outputs(30) <= a;
    outputs(31) <= a;
    outputs(32) <= a xor b;
    outputs(33) <= a;
    outputs(34) <= not b;
    outputs(35) <= not (a xor b);
    outputs(36) <= not (a or b);
    outputs(37) <= a xor b;
    outputs(38) <= b;
    outputs(39) <= a;
    outputs(40) <= not b or a;
    outputs(41) <= b;
    outputs(42) <= not b or a;
    outputs(43) <= b;
    outputs(44) <= a;
    outputs(45) <= a and b;
    outputs(46) <= not a;
    outputs(47) <= a or b;
    outputs(48) <= not a;
    outputs(49) <= a or b;
    outputs(50) <= not (a or b);
    outputs(51) <= a and not b;
    outputs(52) <= a;
    outputs(53) <= a;
    outputs(54) <= a xor b;
    outputs(55) <= a;
    outputs(56) <= not b;
    outputs(57) <= b;
    outputs(58) <= not a;
    outputs(59) <= a and not b;
    outputs(60) <= not (a or b);
    outputs(61) <= not b;
    outputs(62) <= a;
    outputs(63) <= b;
    outputs(64) <= not (a or b);
    outputs(65) <= a xor b;
    outputs(66) <= a;
    outputs(67) <= not b;
    outputs(68) <= b;
    outputs(69) <= not a;
    outputs(70) <= not b;
    outputs(71) <= a xor b;
    outputs(72) <= not (a or b);
    outputs(73) <= a and b;
    outputs(74) <= not a;
    outputs(75) <= not b;
    outputs(76) <= not (a or b);
    outputs(77) <= not (a xor b);
    outputs(78) <= b;
    outputs(79) <= a or b;
    outputs(80) <= b;
    outputs(81) <= a;
    outputs(82) <= not b;
    outputs(83) <= a;
    outputs(84) <= not a;
    outputs(85) <= a and b;
    outputs(86) <= not a;
    outputs(87) <= not a;
    outputs(88) <= not a;
    outputs(89) <= a;
    outputs(90) <= b;
    outputs(91) <= not (a and b);
    outputs(92) <= a;
    outputs(93) <= not b;
    outputs(94) <= not b or a;
    outputs(95) <= a;
    outputs(96) <= not (a and b);
    outputs(97) <= not (a or b);
    outputs(98) <= not (a or b);
    outputs(99) <= not b;
    outputs(100) <= a xor b;
    outputs(101) <= a xor b;
    outputs(102) <= not (a xor b);
    outputs(103) <= b and not a;
    outputs(104) <= not (a xor b);
    outputs(105) <= not b or a;
    outputs(106) <= not b;
    outputs(107) <= not b;
    outputs(108) <= not b;
    outputs(109) <= not (a xor b);
    outputs(110) <= not b;
    outputs(111) <= not b;
    outputs(112) <= b;
    outputs(113) <= not a or b;
    outputs(114) <= not (a or b);
    outputs(115) <= not a;
    outputs(116) <= not b;
    outputs(117) <= b;
    outputs(118) <= b and not a;
    outputs(119) <= a xor b;
    outputs(120) <= a;
    outputs(121) <= a;
    outputs(122) <= not (a or b);
    outputs(123) <= b;
    outputs(124) <= a xor b;
    outputs(125) <= not a;
    outputs(126) <= a;
    outputs(127) <= not b;
    outputs(128) <= not a or b;
    outputs(129) <= not a;
    outputs(130) <= not b;
    outputs(131) <= a;
    outputs(132) <= a or b;
    outputs(133) <= b;
    outputs(134) <= b;
    outputs(135) <= a;
    outputs(136) <= a xor b;
    outputs(137) <= a and b;
    outputs(138) <= a xor b;
    outputs(139) <= b and not a;
    outputs(140) <= b;
    outputs(141) <= not (a and b);
    outputs(142) <= not a;
    outputs(143) <= a xor b;
    outputs(144) <= not a;
    outputs(145) <= a;
    outputs(146) <= a xor b;
    outputs(147) <= a;
    outputs(148) <= not (a xor b);
    outputs(149) <= b and not a;
    outputs(150) <= a and not b;
    outputs(151) <= not (a xor b);
    outputs(152) <= a xor b;
    outputs(153) <= not b;
    outputs(154) <= a and b;
    outputs(155) <= b and not a;
    outputs(156) <= not b;
    outputs(157) <= a;
    outputs(158) <= a;
    outputs(159) <= a and not b;
    outputs(160) <= not b;
    outputs(161) <= a and not b;
    outputs(162) <= not b;
    outputs(163) <= a xor b;
    outputs(164) <= not a or b;
    outputs(165) <= not b;
    outputs(166) <= not a or b;
    outputs(167) <= not a;
    outputs(168) <= not b;
    outputs(169) <= not (a xor b);
    outputs(170) <= not a;
    outputs(171) <= a and b;
    outputs(172) <= a or b;
    outputs(173) <= a;
    outputs(174) <= not a;
    outputs(175) <= not a;
    outputs(176) <= not b;
    outputs(177) <= a xor b;
    outputs(178) <= a;
    outputs(179) <= not (a xor b);
    outputs(180) <= b;
    outputs(181) <= a and b;
    outputs(182) <= not (a xor b);
    outputs(183) <= b;
    outputs(184) <= a or b;
    outputs(185) <= b;
    outputs(186) <= not (a xor b);
    outputs(187) <= not (a and b);
    outputs(188) <= not b;
    outputs(189) <= not (a xor b);
    outputs(190) <= b;
    outputs(191) <= b;
    outputs(192) <= not (a xor b);
    outputs(193) <= not b;
    outputs(194) <= a xor b;
    outputs(195) <= not b;
    outputs(196) <= not b;
    outputs(197) <= a;
    outputs(198) <= not (a xor b);
    outputs(199) <= not a;
    outputs(200) <= a and not b;
    outputs(201) <= not (a or b);
    outputs(202) <= not b;
    outputs(203) <= a and b;
    outputs(204) <= not a;
    outputs(205) <= b;
    outputs(206) <= a;
    outputs(207) <= a;
    outputs(208) <= a and not b;
    outputs(209) <= not a;
    outputs(210) <= a and b;
    outputs(211) <= b and not a;
    outputs(212) <= a;
    outputs(213) <= not (a xor b);
    outputs(214) <= a and b;
    outputs(215) <= not (a and b);
    outputs(216) <= not b;
    outputs(217) <= a xor b;
    outputs(218) <= a and b;
    outputs(219) <= b and not a;
    outputs(220) <= a;
    outputs(221) <= not a;
    outputs(222) <= not b or a;
    outputs(223) <= not a;
    outputs(224) <= not a or b;
    outputs(225) <= a xor b;
    outputs(226) <= not b;
    outputs(227) <= b;
    outputs(228) <= not (a and b);
    outputs(229) <= a;
    outputs(230) <= b and not a;
    outputs(231) <= a;
    outputs(232) <= a xor b;
    outputs(233) <= not (a xor b);
    outputs(234) <= a;
    outputs(235) <= not (a xor b);
    outputs(236) <= not (a xor b);
    outputs(237) <= a and not b;
    outputs(238) <= not (a xor b);
    outputs(239) <= not a;
    outputs(240) <= not (a xor b);
    outputs(241) <= not (a xor b);
    outputs(242) <= a xor b;
    outputs(243) <= a;
    outputs(244) <= not (a or b);
    outputs(245) <= a;
    outputs(246) <= not (a xor b);
    outputs(247) <= a xor b;
    outputs(248) <= a and not b;
    outputs(249) <= not b;
    outputs(250) <= not (a xor b);
    outputs(251) <= b;
    outputs(252) <= a;
    outputs(253) <= a and not b;
    outputs(254) <= not a or b;
    outputs(255) <= a and not b;
    outputs(256) <= a xor b;
    outputs(257) <= not b;
    outputs(258) <= b;
    outputs(259) <= a and not b;
    outputs(260) <= a;
    outputs(261) <= a xor b;
    outputs(262) <= a;
    outputs(263) <= not a;
    outputs(264) <= a and b;
    outputs(265) <= not a;
    outputs(266) <= not (a xor b);
    outputs(267) <= a xor b;
    outputs(268) <= not a;
    outputs(269) <= not a;
    outputs(270) <= not (a or b);
    outputs(271) <= not (a or b);
    outputs(272) <= a and b;
    outputs(273) <= not (a xor b);
    outputs(274) <= not a;
    outputs(275) <= a xor b;
    outputs(276) <= not (a xor b);
    outputs(277) <= a and not b;
    outputs(278) <= not b;
    outputs(279) <= not a or b;
    outputs(280) <= not a;
    outputs(281) <= not (a and b);
    outputs(282) <= a and b;
    outputs(283) <= a xor b;
    outputs(284) <= b;
    outputs(285) <= a xor b;
    outputs(286) <= not b;
    outputs(287) <= b;
    outputs(288) <= not a;
    outputs(289) <= b;
    outputs(290) <= b;
    outputs(291) <= not a;
    outputs(292) <= not b;
    outputs(293) <= a xor b;
    outputs(294) <= not (a xor b);
    outputs(295) <= b;
    outputs(296) <= not b;
    outputs(297) <= not a;
    outputs(298) <= a;
    outputs(299) <= not b or a;
    outputs(300) <= b;
    outputs(301) <= not (a or b);
    outputs(302) <= not b or a;
    outputs(303) <= not b;
    outputs(304) <= b;
    outputs(305) <= a and b;
    outputs(306) <= not (a or b);
    outputs(307) <= b;
    outputs(308) <= not a;
    outputs(309) <= not b;
    outputs(310) <= not a or b;
    outputs(311) <= a;
    outputs(312) <= a xor b;
    outputs(313) <= not a;
    outputs(314) <= b and not a;
    outputs(315) <= not a;
    outputs(316) <= a and b;
    outputs(317) <= not (a and b);
    outputs(318) <= not b;
    outputs(319) <= a;
    outputs(320) <= not (a or b);
    outputs(321) <= not (a xor b);
    outputs(322) <= not b;
    outputs(323) <= not (a or b);
    outputs(324) <= a;
    outputs(325) <= not b or a;
    outputs(326) <= not a;
    outputs(327) <= b;
    outputs(328) <= not (a or b);
    outputs(329) <= not (a or b);
    outputs(330) <= not b;
    outputs(331) <= a xor b;
    outputs(332) <= not a;
    outputs(333) <= not b or a;
    outputs(334) <= b;
    outputs(335) <= a;
    outputs(336) <= a and b;
    outputs(337) <= not (a xor b);
    outputs(338) <= not (a or b);
    outputs(339) <= not b or a;
    outputs(340) <= not a;
    outputs(341) <= not (a and b);
    outputs(342) <= not a;
    outputs(343) <= a and not b;
    outputs(344) <= not a;
    outputs(345) <= a and b;
    outputs(346) <= not b;
    outputs(347) <= not a;
    outputs(348) <= a;
    outputs(349) <= a xor b;
    outputs(350) <= not (a or b);
    outputs(351) <= not b;
    outputs(352) <= not a;
    outputs(353) <= b;
    outputs(354) <= not (a or b);
    outputs(355) <= not (a xor b);
    outputs(356) <= not a;
    outputs(357) <= a and b;
    outputs(358) <= not b;
    outputs(359) <= not (a xor b);
    outputs(360) <= not (a and b);
    outputs(361) <= a xor b;
    outputs(362) <= a and b;
    outputs(363) <= not (a xor b);
    outputs(364) <= a and not b;
    outputs(365) <= not b;
    outputs(366) <= a xor b;
    outputs(367) <= a or b;
    outputs(368) <= not a;
    outputs(369) <= not (a xor b);
    outputs(370) <= a;
    outputs(371) <= a xor b;
    outputs(372) <= a or b;
    outputs(373) <= b;
    outputs(374) <= a xor b;
    outputs(375) <= not (a xor b);
    outputs(376) <= b;
    outputs(377) <= a and not b;
    outputs(378) <= a or b;
    outputs(379) <= a xor b;
    outputs(380) <= not (a or b);
    outputs(381) <= a;
    outputs(382) <= b;
    outputs(383) <= not (a xor b);
    outputs(384) <= a;
    outputs(385) <= a;
    outputs(386) <= b and not a;
    outputs(387) <= a and not b;
    outputs(388) <= a;
    outputs(389) <= b;
    outputs(390) <= not (a xor b);
    outputs(391) <= a xor b;
    outputs(392) <= a and b;
    outputs(393) <= a and not b;
    outputs(394) <= not (a xor b);
    outputs(395) <= not (a xor b);
    outputs(396) <= not b or a;
    outputs(397) <= not (a xor b);
    outputs(398) <= a and not b;
    outputs(399) <= not b;
    outputs(400) <= not b;
    outputs(401) <= a and b;
    outputs(402) <= not a or b;
    outputs(403) <= not b or a;
    outputs(404) <= b;
    outputs(405) <= a;
    outputs(406) <= not b;
    outputs(407) <= not a;
    outputs(408) <= not a or b;
    outputs(409) <= not (a xor b);
    outputs(410) <= not (a xor b);
    outputs(411) <= not a;
    outputs(412) <= not b;
    outputs(413) <= not (a and b);
    outputs(414) <= not (a and b);
    outputs(415) <= b and not a;
    outputs(416) <= not a;
    outputs(417) <= not a;
    outputs(418) <= a xor b;
    outputs(419) <= a and not b;
    outputs(420) <= not (a xor b);
    outputs(421) <= not (a xor b);
    outputs(422) <= a and b;
    outputs(423) <= not b;
    outputs(424) <= not (a xor b);
    outputs(425) <= b;
    outputs(426) <= not b;
    outputs(427) <= a;
    outputs(428) <= not b;
    outputs(429) <= b and not a;
    outputs(430) <= a;
    outputs(431) <= b;
    outputs(432) <= not (a xor b);
    outputs(433) <= b;
    outputs(434) <= b;
    outputs(435) <= not a;
    outputs(436) <= a and b;
    outputs(437) <= a;
    outputs(438) <= a xor b;
    outputs(439) <= a;
    outputs(440) <= not a;
    outputs(441) <= not b;
    outputs(442) <= not (a and b);
    outputs(443) <= not (a xor b);
    outputs(444) <= not b;
    outputs(445) <= b and not a;
    outputs(446) <= b;
    outputs(447) <= a;
    outputs(448) <= not a;
    outputs(449) <= not (a xor b);
    outputs(450) <= not b;
    outputs(451) <= b;
    outputs(452) <= not a or b;
    outputs(453) <= not (a or b);
    outputs(454) <= a and b;
    outputs(455) <= a and not b;
    outputs(456) <= not (a or b);
    outputs(457) <= a xor b;
    outputs(458) <= a or b;
    outputs(459) <= not a;
    outputs(460) <= a;
    outputs(461) <= not a;
    outputs(462) <= not a or b;
    outputs(463) <= a xor b;
    outputs(464) <= not b;
    outputs(465) <= a xor b;
    outputs(466) <= a;
    outputs(467) <= not (a xor b);
    outputs(468) <= b;
    outputs(469) <= a;
    outputs(470) <= b;
    outputs(471) <= not (a or b);
    outputs(472) <= a and b;
    outputs(473) <= b and not a;
    outputs(474) <= not (a xor b);
    outputs(475) <= b;
    outputs(476) <= a xor b;
    outputs(477) <= a xor b;
    outputs(478) <= a or b;
    outputs(479) <= a xor b;
    outputs(480) <= not a;
    outputs(481) <= a;
    outputs(482) <= not a;
    outputs(483) <= a;
    outputs(484) <= not (a or b);
    outputs(485) <= a;
    outputs(486) <= not (a and b);
    outputs(487) <= a xor b;
    outputs(488) <= a xor b;
    outputs(489) <= not a;
    outputs(490) <= not a;
    outputs(491) <= a;
    outputs(492) <= a;
    outputs(493) <= a or b;
    outputs(494) <= a and b;
    outputs(495) <= a;
    outputs(496) <= a and b;
    outputs(497) <= a and b;
    outputs(498) <= not a or b;
    outputs(499) <= not (a xor b);
    outputs(500) <= b;
    outputs(501) <= a xor b;
    outputs(502) <= b;
    outputs(503) <= not (a and b);
    outputs(504) <= not (a or b);
    outputs(505) <= b;
    outputs(506) <= not a;
    outputs(507) <= not a or b;
    outputs(508) <= not (a xor b);
    outputs(509) <= a and not b;
    outputs(510) <= not (a and b);
    outputs(511) <= a;
    outputs(512) <= a;
    outputs(513) <= not (a and b);
    outputs(514) <= not (a xor b);
    outputs(515) <= a xor b;
    outputs(516) <= not (a or b);
    outputs(517) <= not b;
    outputs(518) <= not b;
    outputs(519) <= not a;
    outputs(520) <= a and b;
    outputs(521) <= not (a xor b);
    outputs(522) <= b;
    outputs(523) <= a and not b;
    outputs(524) <= not a;
    outputs(525) <= not (a xor b);
    outputs(526) <= a;
    outputs(527) <= not b;
    outputs(528) <= a;
    outputs(529) <= a xor b;
    outputs(530) <= b and not a;
    outputs(531) <= b and not a;
    outputs(532) <= not a;
    outputs(533) <= a;
    outputs(534) <= a xor b;
    outputs(535) <= not (a xor b);
    outputs(536) <= a;
    outputs(537) <= a and not b;
    outputs(538) <= not b or a;
    outputs(539) <= not (a xor b);
    outputs(540) <= b;
    outputs(541) <= b and not a;
    outputs(542) <= not (a xor b);
    outputs(543) <= a;
    outputs(544) <= not a;
    outputs(545) <= not a;
    outputs(546) <= not (a xor b);
    outputs(547) <= b;
    outputs(548) <= a xor b;
    outputs(549) <= not b or a;
    outputs(550) <= a;
    outputs(551) <= a;
    outputs(552) <= a;
    outputs(553) <= not (a xor b);
    outputs(554) <= b and not a;
    outputs(555) <= not b;
    outputs(556) <= not (a xor b);
    outputs(557) <= not b;
    outputs(558) <= not a;
    outputs(559) <= a xor b;
    outputs(560) <= a;
    outputs(561) <= not b;
    outputs(562) <= a xor b;
    outputs(563) <= not b;
    outputs(564) <= not a;
    outputs(565) <= a;
    outputs(566) <= a xor b;
    outputs(567) <= a;
    outputs(568) <= not a;
    outputs(569) <= a and not b;
    outputs(570) <= not (a xor b);
    outputs(571) <= not a or b;
    outputs(572) <= a;
    outputs(573) <= a and not b;
    outputs(574) <= a and not b;
    outputs(575) <= not a;
    outputs(576) <= not a;
    outputs(577) <= b;
    outputs(578) <= a and not b;
    outputs(579) <= b;
    outputs(580) <= not b or a;
    outputs(581) <= not (a xor b);
    outputs(582) <= a xor b;
    outputs(583) <= a xor b;
    outputs(584) <= a and b;
    outputs(585) <= a and not b;
    outputs(586) <= a;
    outputs(587) <= not (a or b);
    outputs(588) <= not b;
    outputs(589) <= not b;
    outputs(590) <= not (a xor b);
    outputs(591) <= a and b;
    outputs(592) <= a xor b;
    outputs(593) <= not b or a;
    outputs(594) <= a;
    outputs(595) <= not a;
    outputs(596) <= a or b;
    outputs(597) <= b;
    outputs(598) <= a;
    outputs(599) <= not (a xor b);
    outputs(600) <= a xor b;
    outputs(601) <= not a;
    outputs(602) <= not b;
    outputs(603) <= not b;
    outputs(604) <= b and not a;
    outputs(605) <= not b;
    outputs(606) <= a xor b;
    outputs(607) <= not (a xor b);
    outputs(608) <= a or b;
    outputs(609) <= not b;
    outputs(610) <= a and b;
    outputs(611) <= not a;
    outputs(612) <= not (a xor b);
    outputs(613) <= not a;
    outputs(614) <= a;
    outputs(615) <= b and not a;
    outputs(616) <= a and not b;
    outputs(617) <= not a;
    outputs(618) <= a and b;
    outputs(619) <= a or b;
    outputs(620) <= not b;
    outputs(621) <= not a;
    outputs(622) <= a xor b;
    outputs(623) <= not b or a;
    outputs(624) <= not (a xor b);
    outputs(625) <= not (a and b);
    outputs(626) <= not (a or b);
    outputs(627) <= b;
    outputs(628) <= a and b;
    outputs(629) <= not b;
    outputs(630) <= not (a xor b);
    outputs(631) <= not b;
    outputs(632) <= not (a or b);
    outputs(633) <= not b;
    outputs(634) <= a;
    outputs(635) <= a or b;
    outputs(636) <= a;
    outputs(637) <= b;
    outputs(638) <= not b;
    outputs(639) <= not (a or b);
    outputs(640) <= a and not b;
    outputs(641) <= not (a or b);
    outputs(642) <= b;
    outputs(643) <= not a;
    outputs(644) <= not b;
    outputs(645) <= b;
    outputs(646) <= a and not b;
    outputs(647) <= a xor b;
    outputs(648) <= not (a xor b);
    outputs(649) <= not b;
    outputs(650) <= a and not b;
    outputs(651) <= not b;
    outputs(652) <= a xor b;
    outputs(653) <= a;
    outputs(654) <= not a;
    outputs(655) <= a xor b;
    outputs(656) <= b and not a;
    outputs(657) <= not a;
    outputs(658) <= a;
    outputs(659) <= a;
    outputs(660) <= a and b;
    outputs(661) <= a;
    outputs(662) <= b and not a;
    outputs(663) <= a;
    outputs(664) <= not (a xor b);
    outputs(665) <= b;
    outputs(666) <= b;
    outputs(667) <= not (a or b);
    outputs(668) <= not (a xor b);
    outputs(669) <= not b;
    outputs(670) <= not (a xor b);
    outputs(671) <= not b or a;
    outputs(672) <= not (a or b);
    outputs(673) <= not (a and b);
    outputs(674) <= b;
    outputs(675) <= a and not b;
    outputs(676) <= not (a xor b);
    outputs(677) <= a;
    outputs(678) <= a xor b;
    outputs(679) <= not b;
    outputs(680) <= not b or a;
    outputs(681) <= b;
    outputs(682) <= not (a xor b);
    outputs(683) <= a xor b;
    outputs(684) <= a or b;
    outputs(685) <= a xor b;
    outputs(686) <= not b or a;
    outputs(687) <= not b or a;
    outputs(688) <= not (a or b);
    outputs(689) <= not b;
    outputs(690) <= b;
    outputs(691) <= not (a xor b);
    outputs(692) <= b and not a;
    outputs(693) <= not a;
    outputs(694) <= b;
    outputs(695) <= not a;
    outputs(696) <= b;
    outputs(697) <= a xor b;
    outputs(698) <= b;
    outputs(699) <= not a;
    outputs(700) <= not b;
    outputs(701) <= b and not a;
    outputs(702) <= a xor b;
    outputs(703) <= not (a xor b);
    outputs(704) <= b;
    outputs(705) <= a;
    outputs(706) <= not (a or b);
    outputs(707) <= not (a and b);
    outputs(708) <= not (a xor b);
    outputs(709) <= not b;
    outputs(710) <= not (a xor b);
    outputs(711) <= a and not b;
    outputs(712) <= a;
    outputs(713) <= not (a xor b);
    outputs(714) <= b and not a;
    outputs(715) <= not (a or b);
    outputs(716) <= not (a xor b);
    outputs(717) <= not (a xor b);
    outputs(718) <= b;
    outputs(719) <= a and not b;
    outputs(720) <= a and b;
    outputs(721) <= a and not b;
    outputs(722) <= b and not a;
    outputs(723) <= b;
    outputs(724) <= b;
    outputs(725) <= not (a xor b);
    outputs(726) <= not b or a;
    outputs(727) <= not a;
    outputs(728) <= not (a xor b);
    outputs(729) <= not b;
    outputs(730) <= not b or a;
    outputs(731) <= not a;
    outputs(732) <= a;
    outputs(733) <= not a;
    outputs(734) <= not b;
    outputs(735) <= not a;
    outputs(736) <= b and not a;
    outputs(737) <= b;
    outputs(738) <= not (a xor b);
    outputs(739) <= a and not b;
    outputs(740) <= a xor b;
    outputs(741) <= not (a xor b);
    outputs(742) <= not (a xor b);
    outputs(743) <= a xor b;
    outputs(744) <= not b;
    outputs(745) <= not a;
    outputs(746) <= a;
    outputs(747) <= not (a and b);
    outputs(748) <= a;
    outputs(749) <= a xor b;
    outputs(750) <= a xor b;
    outputs(751) <= not (a or b);
    outputs(752) <= b and not a;
    outputs(753) <= not (a or b);
    outputs(754) <= not b;
    outputs(755) <= not b;
    outputs(756) <= not (a or b);
    outputs(757) <= a;
    outputs(758) <= not (a and b);
    outputs(759) <= a;
    outputs(760) <= not b;
    outputs(761) <= a and not b;
    outputs(762) <= a and not b;
    outputs(763) <= not (a or b);
    outputs(764) <= a;
    outputs(765) <= a xor b;
    outputs(766) <= not b or a;
    outputs(767) <= a;
    outputs(768) <= a or b;
    outputs(769) <= a xor b;
    outputs(770) <= b;
    outputs(771) <= a;
    outputs(772) <= a;
    outputs(773) <= not a;
    outputs(774) <= a and not b;
    outputs(775) <= b and not a;
    outputs(776) <= not a;
    outputs(777) <= not b;
    outputs(778) <= not a;
    outputs(779) <= not (a xor b);
    outputs(780) <= not a or b;
    outputs(781) <= a and b;
    outputs(782) <= a xor b;
    outputs(783) <= not b;
    outputs(784) <= b and not a;
    outputs(785) <= b;
    outputs(786) <= not b;
    outputs(787) <= a xor b;
    outputs(788) <= not a or b;
    outputs(789) <= not a;
    outputs(790) <= not b;
    outputs(791) <= a;
    outputs(792) <= b and not a;
    outputs(793) <= a;
    outputs(794) <= a;
    outputs(795) <= not (a xor b);
    outputs(796) <= a xor b;
    outputs(797) <= a;
    outputs(798) <= not b;
    outputs(799) <= a xor b;
    outputs(800) <= not b;
    outputs(801) <= a;
    outputs(802) <= a and not b;
    outputs(803) <= not a;
    outputs(804) <= a;
    outputs(805) <= b;
    outputs(806) <= not a;
    outputs(807) <= a xor b;
    outputs(808) <= b and not a;
    outputs(809) <= not (a xor b);
    outputs(810) <= a and not b;
    outputs(811) <= not (a or b);
    outputs(812) <= a;
    outputs(813) <= not b or a;
    outputs(814) <= not b;
    outputs(815) <= not a;
    outputs(816) <= b and not a;
    outputs(817) <= not b;
    outputs(818) <= b;
    outputs(819) <= not (a xor b);
    outputs(820) <= not (a xor b);
    outputs(821) <= b;
    outputs(822) <= not b;
    outputs(823) <= not b;
    outputs(824) <= not (a xor b);
    outputs(825) <= not (a xor b);
    outputs(826) <= a;
    outputs(827) <= b;
    outputs(828) <= a xor b;
    outputs(829) <= a and b;
    outputs(830) <= not a;
    outputs(831) <= not (a and b);
    outputs(832) <= not (a xor b);
    outputs(833) <= not (a and b);
    outputs(834) <= b;
    outputs(835) <= not (a or b);
    outputs(836) <= b and not a;
    outputs(837) <= not a;
    outputs(838) <= a xor b;
    outputs(839) <= not b;
    outputs(840) <= a and b;
    outputs(841) <= a;
    outputs(842) <= a xor b;
    outputs(843) <= b;
    outputs(844) <= a and b;
    outputs(845) <= not (a xor b);
    outputs(846) <= not b;
    outputs(847) <= a xor b;
    outputs(848) <= a xor b;
    outputs(849) <= not a or b;
    outputs(850) <= not (a xor b);
    outputs(851) <= a;
    outputs(852) <= a xor b;
    outputs(853) <= a or b;
    outputs(854) <= b;
    outputs(855) <= a xor b;
    outputs(856) <= a and b;
    outputs(857) <= b;
    outputs(858) <= not (a or b);
    outputs(859) <= b;
    outputs(860) <= a;
    outputs(861) <= b;
    outputs(862) <= a;
    outputs(863) <= not (a xor b);
    outputs(864) <= a and not b;
    outputs(865) <= not (a or b);
    outputs(866) <= not a;
    outputs(867) <= not b;
    outputs(868) <= b;
    outputs(869) <= not a or b;
    outputs(870) <= b;
    outputs(871) <= b and not a;
    outputs(872) <= not a;
    outputs(873) <= not b;
    outputs(874) <= not a;
    outputs(875) <= a and b;
    outputs(876) <= not (a or b);
    outputs(877) <= not (a or b);
    outputs(878) <= not b;
    outputs(879) <= a xor b;
    outputs(880) <= not b;
    outputs(881) <= not (a xor b);
    outputs(882) <= b;
    outputs(883) <= not b;
    outputs(884) <= b;
    outputs(885) <= not a;
    outputs(886) <= b;
    outputs(887) <= a and b;
    outputs(888) <= b and not a;
    outputs(889) <= a;
    outputs(890) <= a;
    outputs(891) <= not (a xor b);
    outputs(892) <= a or b;
    outputs(893) <= a;
    outputs(894) <= not (a xor b);
    outputs(895) <= not (a xor b);
    outputs(896) <= not (a xor b);
    outputs(897) <= a and not b;
    outputs(898) <= a xor b;
    outputs(899) <= not (a xor b);
    outputs(900) <= a;
    outputs(901) <= not b;
    outputs(902) <= b;
    outputs(903) <= b;
    outputs(904) <= a xor b;
    outputs(905) <= not b;
    outputs(906) <= not a;
    outputs(907) <= a and not b;
    outputs(908) <= a and not b;
    outputs(909) <= not a or b;
    outputs(910) <= not a;
    outputs(911) <= b and not a;
    outputs(912) <= a;
    outputs(913) <= a and b;
    outputs(914) <= not a or b;
    outputs(915) <= a or b;
    outputs(916) <= not a;
    outputs(917) <= a and b;
    outputs(918) <= not (a or b);
    outputs(919) <= a xor b;
    outputs(920) <= a xor b;
    outputs(921) <= a and not b;
    outputs(922) <= b;
    outputs(923) <= a;
    outputs(924) <= a or b;
    outputs(925) <= not (a xor b);
    outputs(926) <= b;
    outputs(927) <= not a;
    outputs(928) <= not b;
    outputs(929) <= b;
    outputs(930) <= not a;
    outputs(931) <= a;
    outputs(932) <= a xor b;
    outputs(933) <= a and b;
    outputs(934) <= not b;
    outputs(935) <= not b;
    outputs(936) <= not a or b;
    outputs(937) <= not (a xor b);
    outputs(938) <= not a;
    outputs(939) <= a xor b;
    outputs(940) <= b;
    outputs(941) <= not (a xor b);
    outputs(942) <= a or b;
    outputs(943) <= not a;
    outputs(944) <= not a or b;
    outputs(945) <= a xor b;
    outputs(946) <= not (a and b);
    outputs(947) <= b;
    outputs(948) <= a and b;
    outputs(949) <= b and not a;
    outputs(950) <= not (a xor b);
    outputs(951) <= a;
    outputs(952) <= a and not b;
    outputs(953) <= a xor b;
    outputs(954) <= b and not a;
    outputs(955) <= not a;
    outputs(956) <= a;
    outputs(957) <= not b;
    outputs(958) <= b and not a;
    outputs(959) <= not (a xor b);
    outputs(960) <= a or b;
    outputs(961) <= not b;
    outputs(962) <= a xor b;
    outputs(963) <= not a;
    outputs(964) <= not a or b;
    outputs(965) <= not b or a;
    outputs(966) <= b;
    outputs(967) <= not b;
    outputs(968) <= b;
    outputs(969) <= not b;
    outputs(970) <= not b;
    outputs(971) <= not a;
    outputs(972) <= not a;
    outputs(973) <= a;
    outputs(974) <= b;
    outputs(975) <= a;
    outputs(976) <= not (a xor b);
    outputs(977) <= not b or a;
    outputs(978) <= not b or a;
    outputs(979) <= not b;
    outputs(980) <= not a;
    outputs(981) <= a and b;
    outputs(982) <= not a;
    outputs(983) <= b;
    outputs(984) <= a xor b;
    outputs(985) <= not (a xor b);
    outputs(986) <= not a;
    outputs(987) <= not b;
    outputs(988) <= b and not a;
    outputs(989) <= b;
    outputs(990) <= not (a xor b);
    outputs(991) <= not b;
    outputs(992) <= a and not b;
    outputs(993) <= not (a xor b);
    outputs(994) <= b;
    outputs(995) <= a or b;
    outputs(996) <= not (a and b);
    outputs(997) <= not (a and b);
    outputs(998) <= a and not b;
    outputs(999) <= not b;
    outputs(1000) <= b;
    outputs(1001) <= not b;
    outputs(1002) <= a xor b;
    outputs(1003) <= not (a xor b);
    outputs(1004) <= not a;
    outputs(1005) <= b;
    outputs(1006) <= b;
    outputs(1007) <= b;
    outputs(1008) <= not (a or b);
    outputs(1009) <= not (a xor b);
    outputs(1010) <= a;
    outputs(1011) <= not (a xor b);
    outputs(1012) <= not (a xor b);
    outputs(1013) <= not (a xor b);
    outputs(1014) <= not (a xor b);
    outputs(1015) <= b;
    outputs(1016) <= a or b;
    outputs(1017) <= not (a xor b);
    outputs(1018) <= b;
    outputs(1019) <= b;
    outputs(1020) <= not a;
    outputs(1021) <= not (a xor b);
    outputs(1022) <= a xor b;
    outputs(1023) <= not b;
    outputs(1024) <= a and b;
    outputs(1025) <= not (a xor b);
    outputs(1026) <= a xor b;
    outputs(1027) <= a and b;
    outputs(1028) <= a xor b;
    outputs(1029) <= b;
    outputs(1030) <= not (a or b);
    outputs(1031) <= not b;
    outputs(1032) <= a xor b;
    outputs(1033) <= not b;
    outputs(1034) <= a xor b;
    outputs(1035) <= b;
    outputs(1036) <= b;
    outputs(1037) <= b and not a;
    outputs(1038) <= a xor b;
    outputs(1039) <= a and b;
    outputs(1040) <= not b;
    outputs(1041) <= b;
    outputs(1042) <= a xor b;
    outputs(1043) <= not b;
    outputs(1044) <= b;
    outputs(1045) <= not (a or b);
    outputs(1046) <= not a;
    outputs(1047) <= a xor b;
    outputs(1048) <= b and not a;
    outputs(1049) <= a;
    outputs(1050) <= not (a or b);
    outputs(1051) <= not (a xor b);
    outputs(1052) <= a and not b;
    outputs(1053) <= not (a or b);
    outputs(1054) <= not (a xor b);
    outputs(1055) <= a xor b;
    outputs(1056) <= a xor b;
    outputs(1057) <= not (a or b);
    outputs(1058) <= not (a xor b);
    outputs(1059) <= a xor b;
    outputs(1060) <= not (a or b);
    outputs(1061) <= not b;
    outputs(1062) <= a and not b;
    outputs(1063) <= not (a or b);
    outputs(1064) <= not (a xor b);
    outputs(1065) <= not (a or b);
    outputs(1066) <= not (a xor b);
    outputs(1067) <= b and not a;
    outputs(1068) <= b and not a;
    outputs(1069) <= a and not b;
    outputs(1070) <= a xor b;
    outputs(1071) <= not a or b;
    outputs(1072) <= '0';
    outputs(1073) <= not (a or b);
    outputs(1074) <= b and not a;
    outputs(1075) <= not (a xor b);
    outputs(1076) <= a;
    outputs(1077) <= a xor b;
    outputs(1078) <= a xor b;
    outputs(1079) <= a xor b;
    outputs(1080) <= a and b;
    outputs(1081) <= a xor b;
    outputs(1082) <= a xor b;
    outputs(1083) <= a and not b;
    outputs(1084) <= not b;
    outputs(1085) <= '0';
    outputs(1086) <= not (a or b);
    outputs(1087) <= a and not b;
    outputs(1088) <= not (a xor b);
    outputs(1089) <= not (a xor b);
    outputs(1090) <= not (a xor b);
    outputs(1091) <= a and not b;
    outputs(1092) <= not b;
    outputs(1093) <= a xor b;
    outputs(1094) <= a xor b;
    outputs(1095) <= not a;
    outputs(1096) <= a;
    outputs(1097) <= a;
    outputs(1098) <= b;
    outputs(1099) <= a and not b;
    outputs(1100) <= a and not b;
    outputs(1101) <= a and b;
    outputs(1102) <= b and not a;
    outputs(1103) <= not (a or b);
    outputs(1104) <= not (a or b);
    outputs(1105) <= b;
    outputs(1106) <= not a;
    outputs(1107) <= a xor b;
    outputs(1108) <= a and not b;
    outputs(1109) <= b and not a;
    outputs(1110) <= b and not a;
    outputs(1111) <= a xor b;
    outputs(1112) <= b;
    outputs(1113) <= not (a xor b);
    outputs(1114) <= a xor b;
    outputs(1115) <= not (a or b);
    outputs(1116) <= a xor b;
    outputs(1117) <= a and not b;
    outputs(1118) <= b;
    outputs(1119) <= b;
    outputs(1120) <= not (a xor b);
    outputs(1121) <= a xor b;
    outputs(1122) <= '0';
    outputs(1123) <= a xor b;
    outputs(1124) <= not (a or b);
    outputs(1125) <= not a or b;
    outputs(1126) <= not b;
    outputs(1127) <= a xor b;
    outputs(1128) <= a xor b;
    outputs(1129) <= not b;
    outputs(1130) <= b;
    outputs(1131) <= a;
    outputs(1132) <= a and b;
    outputs(1133) <= not b;
    outputs(1134) <= b;
    outputs(1135) <= not (a or b);
    outputs(1136) <= a xor b;
    outputs(1137) <= not b or a;
    outputs(1138) <= not b;
    outputs(1139) <= not (a xor b);
    outputs(1140) <= a;
    outputs(1141) <= not b;
    outputs(1142) <= a xor b;
    outputs(1143) <= not (a or b);
    outputs(1144) <= a and b;
    outputs(1145) <= not a;
    outputs(1146) <= a and b;
    outputs(1147) <= a xor b;
    outputs(1148) <= a xor b;
    outputs(1149) <= b and not a;
    outputs(1150) <= a xor b;
    outputs(1151) <= not (a xor b);
    outputs(1152) <= a;
    outputs(1153) <= b;
    outputs(1154) <= not (a xor b);
    outputs(1155) <= not b;
    outputs(1156) <= b;
    outputs(1157) <= a and b;
    outputs(1158) <= a xor b;
    outputs(1159) <= not a;
    outputs(1160) <= b and not a;
    outputs(1161) <= a or b;
    outputs(1162) <= b;
    outputs(1163) <= b;
    outputs(1164) <= a and b;
    outputs(1165) <= not a;
    outputs(1166) <= not (a xor b);
    outputs(1167) <= a xor b;
    outputs(1168) <= a xor b;
    outputs(1169) <= a xor b;
    outputs(1170) <= not (a xor b);
    outputs(1171) <= a and b;
    outputs(1172) <= '0';
    outputs(1173) <= not b;
    outputs(1174) <= b;
    outputs(1175) <= not a;
    outputs(1176) <= a and not b;
    outputs(1177) <= a xor b;
    outputs(1178) <= not (a xor b);
    outputs(1179) <= a xor b;
    outputs(1180) <= not (a or b);
    outputs(1181) <= not (a xor b);
    outputs(1182) <= not a or b;
    outputs(1183) <= b and not a;
    outputs(1184) <= a and not b;
    outputs(1185) <= a xor b;
    outputs(1186) <= not b;
    outputs(1187) <= not b;
    outputs(1188) <= a;
    outputs(1189) <= a and not b;
    outputs(1190) <= '0';
    outputs(1191) <= not (a xor b);
    outputs(1192) <= not (a or b);
    outputs(1193) <= b and not a;
    outputs(1194) <= a xor b;
    outputs(1195) <= not a;
    outputs(1196) <= a and b;
    outputs(1197) <= b;
    outputs(1198) <= not b or a;
    outputs(1199) <= not (a xor b);
    outputs(1200) <= not b;
    outputs(1201) <= not (a or b);
    outputs(1202) <= not (a or b);
    outputs(1203) <= not (a xor b);
    outputs(1204) <= not (a xor b);
    outputs(1205) <= a and not b;
    outputs(1206) <= not (a xor b);
    outputs(1207) <= not b;
    outputs(1208) <= not (a xor b);
    outputs(1209) <= a xor b;
    outputs(1210) <= b;
    outputs(1211) <= not a;
    outputs(1212) <= not (a or b);
    outputs(1213) <= a and b;
    outputs(1214) <= not (a xor b);
    outputs(1215) <= a and b;
    outputs(1216) <= a;
    outputs(1217) <= a xor b;
    outputs(1218) <= a and not b;
    outputs(1219) <= a xor b;
    outputs(1220) <= a;
    outputs(1221) <= a and not b;
    outputs(1222) <= a and b;
    outputs(1223) <= b;
    outputs(1224) <= a and not b;
    outputs(1225) <= b and not a;
    outputs(1226) <= a and b;
    outputs(1227) <= not a;
    outputs(1228) <= a xor b;
    outputs(1229) <= not (a or b);
    outputs(1230) <= not (a xor b);
    outputs(1231) <= not (a or b);
    outputs(1232) <= a xor b;
    outputs(1233) <= b and not a;
    outputs(1234) <= b and not a;
    outputs(1235) <= a and b;
    outputs(1236) <= a and not b;
    outputs(1237) <= a and b;
    outputs(1238) <= not (a xor b);
    outputs(1239) <= not (a or b);
    outputs(1240) <= a xor b;
    outputs(1241) <= not a;
    outputs(1242) <= a;
    outputs(1243) <= a;
    outputs(1244) <= not b;
    outputs(1245) <= not a;
    outputs(1246) <= b;
    outputs(1247) <= a xor b;
    outputs(1248) <= a;
    outputs(1249) <= a and not b;
    outputs(1250) <= a xor b;
    outputs(1251) <= not a;
    outputs(1252) <= b;
    outputs(1253) <= a or b;
    outputs(1254) <= b;
    outputs(1255) <= a;
    outputs(1256) <= not (a xor b);
    outputs(1257) <= a;
    outputs(1258) <= a xor b;
    outputs(1259) <= not a;
    outputs(1260) <= b;
    outputs(1261) <= b;
    outputs(1262) <= not (a xor b);
    outputs(1263) <= not b;
    outputs(1264) <= not b or a;
    outputs(1265) <= not (a xor b);
    outputs(1266) <= not b;
    outputs(1267) <= not b;
    outputs(1268) <= not a;
    outputs(1269) <= not b;
    outputs(1270) <= a and not b;
    outputs(1271) <= b and not a;
    outputs(1272) <= not a;
    outputs(1273) <= a;
    outputs(1274) <= not a;
    outputs(1275) <= not b;
    outputs(1276) <= not b;
    outputs(1277) <= a;
    outputs(1278) <= not (a xor b);
    outputs(1279) <= '0';
    outputs(1280) <= b and not a;
    outputs(1281) <= b and not a;
    outputs(1282) <= a xor b;
    outputs(1283) <= not a;
    outputs(1284) <= not (a xor b);
    outputs(1285) <= not a;
    outputs(1286) <= not (a xor b);
    outputs(1287) <= not (a or b);
    outputs(1288) <= '0';
    outputs(1289) <= b and not a;
    outputs(1290) <= a xor b;
    outputs(1291) <= not a;
    outputs(1292) <= b;
    outputs(1293) <= a and b;
    outputs(1294) <= a and not b;
    outputs(1295) <= b;
    outputs(1296) <= not b;
    outputs(1297) <= a xor b;
    outputs(1298) <= not a;
    outputs(1299) <= not (a or b);
    outputs(1300) <= b and not a;
    outputs(1301) <= not (a xor b);
    outputs(1302) <= not (a xor b);
    outputs(1303) <= a xor b;
    outputs(1304) <= a and b;
    outputs(1305) <= not b;
    outputs(1306) <= a xor b;
    outputs(1307) <= a and not b;
    outputs(1308) <= not b;
    outputs(1309) <= not b;
    outputs(1310) <= a and b;
    outputs(1311) <= not (a xor b);
    outputs(1312) <= not (a xor b);
    outputs(1313) <= not (a xor b);
    outputs(1314) <= not (a or b);
    outputs(1315) <= b;
    outputs(1316) <= not (a xor b);
    outputs(1317) <= not (a xor b);
    outputs(1318) <= not (a or b);
    outputs(1319) <= a and b;
    outputs(1320) <= not (a xor b);
    outputs(1321) <= a;
    outputs(1322) <= a and not b;
    outputs(1323) <= a xor b;
    outputs(1324) <= a and b;
    outputs(1325) <= a xor b;
    outputs(1326) <= b and not a;
    outputs(1327) <= not (a xor b);
    outputs(1328) <= not (a xor b);
    outputs(1329) <= b and not a;
    outputs(1330) <= a and not b;
    outputs(1331) <= a;
    outputs(1332) <= not a;
    outputs(1333) <= a or b;
    outputs(1334) <= a xor b;
    outputs(1335) <= not b;
    outputs(1336) <= not b;
    outputs(1337) <= not (a xor b);
    outputs(1338) <= not a;
    outputs(1339) <= not b;
    outputs(1340) <= not b;
    outputs(1341) <= a and b;
    outputs(1342) <= not b;
    outputs(1343) <= not (a xor b);
    outputs(1344) <= not b;
    outputs(1345) <= a xor b;
    outputs(1346) <= not (a xor b);
    outputs(1347) <= a and not b;
    outputs(1348) <= a;
    outputs(1349) <= b and not a;
    outputs(1350) <= not a;
    outputs(1351) <= a xor b;
    outputs(1352) <= not (a or b);
    outputs(1353) <= not a;
    outputs(1354) <= not (a or b);
    outputs(1355) <= not (a xor b);
    outputs(1356) <= not (a xor b);
    outputs(1357) <= not (a xor b);
    outputs(1358) <= not b;
    outputs(1359) <= b;
    outputs(1360) <= b;
    outputs(1361) <= not (a xor b);
    outputs(1362) <= not (a or b);
    outputs(1363) <= not b;
    outputs(1364) <= a and not b;
    outputs(1365) <= not (a or b);
    outputs(1366) <= not (a xor b);
    outputs(1367) <= not a;
    outputs(1368) <= a xor b;
    outputs(1369) <= not (a xor b);
    outputs(1370) <= not (a xor b);
    outputs(1371) <= a;
    outputs(1372) <= not a;
    outputs(1373) <= not a;
    outputs(1374) <= not (a xor b);
    outputs(1375) <= not a;
    outputs(1376) <= not a;
    outputs(1377) <= not (a xor b);
    outputs(1378) <= a;
    outputs(1379) <= b;
    outputs(1380) <= a xor b;
    outputs(1381) <= not (a xor b);
    outputs(1382) <= not b;
    outputs(1383) <= a xor b;
    outputs(1384) <= a xor b;
    outputs(1385) <= not (a xor b);
    outputs(1386) <= not (a xor b);
    outputs(1387) <= not (a xor b);
    outputs(1388) <= b;
    outputs(1389) <= a;
    outputs(1390) <= not a;
    outputs(1391) <= a and b;
    outputs(1392) <= a and not b;
    outputs(1393) <= not (a xor b);
    outputs(1394) <= not (a xor b);
    outputs(1395) <= a;
    outputs(1396) <= not (a xor b);
    outputs(1397) <= b and not a;
    outputs(1398) <= not (a xor b);
    outputs(1399) <= a and b;
    outputs(1400) <= a xor b;
    outputs(1401) <= a and not b;
    outputs(1402) <= '0';
    outputs(1403) <= not a;
    outputs(1404) <= b;
    outputs(1405) <= a and b;
    outputs(1406) <= not (a xor b);
    outputs(1407) <= not b;
    outputs(1408) <= not (a xor b);
    outputs(1409) <= a and not b;
    outputs(1410) <= not (a xor b);
    outputs(1411) <= not (a xor b);
    outputs(1412) <= a xor b;
    outputs(1413) <= a and b;
    outputs(1414) <= a xor b;
    outputs(1415) <= a and b;
    outputs(1416) <= a and b;
    outputs(1417) <= b and not a;
    outputs(1418) <= a and b;
    outputs(1419) <= not (a xor b);
    outputs(1420) <= not a;
    outputs(1421) <= not (a xor b);
    outputs(1422) <= not (a xor b);
    outputs(1423) <= not b;
    outputs(1424) <= not (a or b);
    outputs(1425) <= not (a xor b);
    outputs(1426) <= b and not a;
    outputs(1427) <= not (a xor b);
    outputs(1428) <= a xor b;
    outputs(1429) <= not b;
    outputs(1430) <= a and b;
    outputs(1431) <= a xor b;
    outputs(1432) <= not (a or b);
    outputs(1433) <= not (a or b);
    outputs(1434) <= a xor b;
    outputs(1435) <= not (a xor b);
    outputs(1436) <= a xor b;
    outputs(1437) <= not (a xor b);
    outputs(1438) <= a xor b;
    outputs(1439) <= a and b;
    outputs(1440) <= not (a xor b);
    outputs(1441) <= a;
    outputs(1442) <= not (a xor b);
    outputs(1443) <= b and not a;
    outputs(1444) <= not (a or b);
    outputs(1445) <= a and b;
    outputs(1446) <= b;
    outputs(1447) <= a xor b;
    outputs(1448) <= not (a or b);
    outputs(1449) <= b and not a;
    outputs(1450) <= a xor b;
    outputs(1451) <= a xor b;
    outputs(1452) <= not a;
    outputs(1453) <= a xor b;
    outputs(1454) <= not (a xor b);
    outputs(1455) <= a;
    outputs(1456) <= not b;
    outputs(1457) <= a;
    outputs(1458) <= '0';
    outputs(1459) <= b and not a;
    outputs(1460) <= not (a or b);
    outputs(1461) <= not b;
    outputs(1462) <= a;
    outputs(1463) <= not a;
    outputs(1464) <= not b or a;
    outputs(1465) <= not (a or b);
    outputs(1466) <= a xor b;
    outputs(1467) <= a and b;
    outputs(1468) <= a and b;
    outputs(1469) <= a xor b;
    outputs(1470) <= a and not b;
    outputs(1471) <= b;
    outputs(1472) <= not (a xor b);
    outputs(1473) <= a and not b;
    outputs(1474) <= not (a or b);
    outputs(1475) <= a and not b;
    outputs(1476) <= not b;
    outputs(1477) <= a xor b;
    outputs(1478) <= not (a xor b);
    outputs(1479) <= b and not a;
    outputs(1480) <= a and b;
    outputs(1481) <= a and not b;
    outputs(1482) <= not (a xor b);
    outputs(1483) <= b and not a;
    outputs(1484) <= a and b;
    outputs(1485) <= b and not a;
    outputs(1486) <= a xor b;
    outputs(1487) <= b and not a;
    outputs(1488) <= a and b;
    outputs(1489) <= a and b;
    outputs(1490) <= b;
    outputs(1491) <= not a;
    outputs(1492) <= not (a xor b);
    outputs(1493) <= a and b;
    outputs(1494) <= b and not a;
    outputs(1495) <= not b;
    outputs(1496) <= a and b;
    outputs(1497) <= '0';
    outputs(1498) <= not b;
    outputs(1499) <= not (a and b);
    outputs(1500) <= b and not a;
    outputs(1501) <= not (a or b);
    outputs(1502) <= a;
    outputs(1503) <= a xor b;
    outputs(1504) <= not b or a;
    outputs(1505) <= a;
    outputs(1506) <= a and not b;
    outputs(1507) <= not a;
    outputs(1508) <= a;
    outputs(1509) <= not b;
    outputs(1510) <= a xor b;
    outputs(1511) <= a and not b;
    outputs(1512) <= not a;
    outputs(1513) <= b and not a;
    outputs(1514) <= not (a or b);
    outputs(1515) <= not (a xor b);
    outputs(1516) <= not (a or b);
    outputs(1517) <= a xor b;
    outputs(1518) <= a;
    outputs(1519) <= not b;
    outputs(1520) <= a xor b;
    outputs(1521) <= a;
    outputs(1522) <= a and not b;
    outputs(1523) <= a and b;
    outputs(1524) <= a xor b;
    outputs(1525) <= not (a xor b);
    outputs(1526) <= not b;
    outputs(1527) <= a;
    outputs(1528) <= not (a or b);
    outputs(1529) <= not (a or b);
    outputs(1530) <= a xor b;
    outputs(1531) <= a and not b;
    outputs(1532) <= b;
    outputs(1533) <= not b;
    outputs(1534) <= not a;
    outputs(1535) <= b;
    outputs(1536) <= a and not b;
    outputs(1537) <= not (a xor b);
    outputs(1538) <= a xor b;
    outputs(1539) <= not (a xor b);
    outputs(1540) <= b;
    outputs(1541) <= a and b;
    outputs(1542) <= '0';
    outputs(1543) <= b;
    outputs(1544) <= a and not b;
    outputs(1545) <= a and b;
    outputs(1546) <= a xor b;
    outputs(1547) <= not b;
    outputs(1548) <= not (a xor b);
    outputs(1549) <= a and b;
    outputs(1550) <= a xor b;
    outputs(1551) <= not b;
    outputs(1552) <= not (a xor b);
    outputs(1553) <= b and not a;
    outputs(1554) <= a xor b;
    outputs(1555) <= not b;
    outputs(1556) <= not b;
    outputs(1557) <= a xor b;
    outputs(1558) <= a and not b;
    outputs(1559) <= not b;
    outputs(1560) <= a xor b;
    outputs(1561) <= b;
    outputs(1562) <= b;
    outputs(1563) <= not b;
    outputs(1564) <= not (a xor b);
    outputs(1565) <= not b;
    outputs(1566) <= not b;
    outputs(1567) <= a xor b;
    outputs(1568) <= not (a xor b);
    outputs(1569) <= a and b;
    outputs(1570) <= not (a xor b);
    outputs(1571) <= b;
    outputs(1572) <= not (a or b);
    outputs(1573) <= a xor b;
    outputs(1574) <= a and b;
    outputs(1575) <= a;
    outputs(1576) <= a xor b;
    outputs(1577) <= a and not b;
    outputs(1578) <= b;
    outputs(1579) <= not a;
    outputs(1580) <= b;
    outputs(1581) <= not (a or b);
    outputs(1582) <= a;
    outputs(1583) <= a xor b;
    outputs(1584) <= a and b;
    outputs(1585) <= b;
    outputs(1586) <= b and not a;
    outputs(1587) <= not (a xor b);
    outputs(1588) <= not (a xor b);
    outputs(1589) <= a;
    outputs(1590) <= a and b;
    outputs(1591) <= not (a or b);
    outputs(1592) <= a;
    outputs(1593) <= not (a or b);
    outputs(1594) <= b and not a;
    outputs(1595) <= b;
    outputs(1596) <= not (a xor b);
    outputs(1597) <= a and b;
    outputs(1598) <= not (a xor b);
    outputs(1599) <= not (a xor b);
    outputs(1600) <= a and b;
    outputs(1601) <= b;
    outputs(1602) <= not b;
    outputs(1603) <= not (a xor b);
    outputs(1604) <= not (a xor b);
    outputs(1605) <= not (a xor b);
    outputs(1606) <= b;
    outputs(1607) <= a;
    outputs(1608) <= not b;
    outputs(1609) <= a and b;
    outputs(1610) <= a or b;
    outputs(1611) <= a and b;
    outputs(1612) <= not b;
    outputs(1613) <= not (a or b);
    outputs(1614) <= a xor b;
    outputs(1615) <= not b;
    outputs(1616) <= a and b;
    outputs(1617) <= a and not b;
    outputs(1618) <= a and not b;
    outputs(1619) <= a and not b;
    outputs(1620) <= not (a xor b);
    outputs(1621) <= '0';
    outputs(1622) <= not (a or b);
    outputs(1623) <= not a;
    outputs(1624) <= not b or a;
    outputs(1625) <= not b;
    outputs(1626) <= not a;
    outputs(1627) <= a and not b;
    outputs(1628) <= a xor b;
    outputs(1629) <= not (a or b);
    outputs(1630) <= not (a xor b);
    outputs(1631) <= not b;
    outputs(1632) <= a and not b;
    outputs(1633) <= not a;
    outputs(1634) <= not (a or b);
    outputs(1635) <= not (a xor b);
    outputs(1636) <= a;
    outputs(1637) <= b;
    outputs(1638) <= not (a or b);
    outputs(1639) <= not a;
    outputs(1640) <= not b;
    outputs(1641) <= not (a or b);
    outputs(1642) <= a;
    outputs(1643) <= a xor b;
    outputs(1644) <= b;
    outputs(1645) <= a;
    outputs(1646) <= not a;
    outputs(1647) <= a;
    outputs(1648) <= a and not b;
    outputs(1649) <= a and b;
    outputs(1650) <= not (a or b);
    outputs(1651) <= a;
    outputs(1652) <= a and b;
    outputs(1653) <= a;
    outputs(1654) <= b and not a;
    outputs(1655) <= not (a xor b);
    outputs(1656) <= '0';
    outputs(1657) <= a or b;
    outputs(1658) <= not (a or b);
    outputs(1659) <= not (a xor b);
    outputs(1660) <= a and not b;
    outputs(1661) <= not (a or b);
    outputs(1662) <= not a;
    outputs(1663) <= a xor b;
    outputs(1664) <= not a;
    outputs(1665) <= b;
    outputs(1666) <= not (a or b);
    outputs(1667) <= not (a xor b);
    outputs(1668) <= not (a or b);
    outputs(1669) <= not a;
    outputs(1670) <= b and not a;
    outputs(1671) <= b and not a;
    outputs(1672) <= not b;
    outputs(1673) <= not (a xor b);
    outputs(1674) <= a;
    outputs(1675) <= not a;
    outputs(1676) <= b;
    outputs(1677) <= not (a xor b);
    outputs(1678) <= a xor b;
    outputs(1679) <= not b;
    outputs(1680) <= not (a xor b);
    outputs(1681) <= b;
    outputs(1682) <= b and not a;
    outputs(1683) <= a xor b;
    outputs(1684) <= not (a xor b);
    outputs(1685) <= a and b;
    outputs(1686) <= a xor b;
    outputs(1687) <= not (a and b);
    outputs(1688) <= not (a xor b);
    outputs(1689) <= not a;
    outputs(1690) <= a;
    outputs(1691) <= b;
    outputs(1692) <= not (a or b);
    outputs(1693) <= a and b;
    outputs(1694) <= b;
    outputs(1695) <= not b;
    outputs(1696) <= not a;
    outputs(1697) <= not a;
    outputs(1698) <= b;
    outputs(1699) <= b and not a;
    outputs(1700) <= not (a or b);
    outputs(1701) <= a and b;
    outputs(1702) <= not (a xor b);
    outputs(1703) <= not (a xor b);
    outputs(1704) <= a;
    outputs(1705) <= a and b;
    outputs(1706) <= a and b;
    outputs(1707) <= a and not b;
    outputs(1708) <= not (a or b);
    outputs(1709) <= a xor b;
    outputs(1710) <= a xor b;
    outputs(1711) <= not b;
    outputs(1712) <= not (a xor b);
    outputs(1713) <= b;
    outputs(1714) <= a and b;
    outputs(1715) <= not (a xor b);
    outputs(1716) <= b and not a;
    outputs(1717) <= not b or a;
    outputs(1718) <= not b;
    outputs(1719) <= a xor b;
    outputs(1720) <= a and not b;
    outputs(1721) <= b;
    outputs(1722) <= not a;
    outputs(1723) <= not a;
    outputs(1724) <= a and not b;
    outputs(1725) <= b;
    outputs(1726) <= b and not a;
    outputs(1727) <= not (a xor b);
    outputs(1728) <= not (a xor b);
    outputs(1729) <= b;
    outputs(1730) <= not (a or b);
    outputs(1731) <= not (a xor b);
    outputs(1732) <= not a;
    outputs(1733) <= a and not b;
    outputs(1734) <= b and not a;
    outputs(1735) <= not (a or b);
    outputs(1736) <= not (a xor b);
    outputs(1737) <= not (a or b);
    outputs(1738) <= a xor b;
    outputs(1739) <= a and b;
    outputs(1740) <= not (a xor b);
    outputs(1741) <= not a;
    outputs(1742) <= a;
    outputs(1743) <= b and not a;
    outputs(1744) <= not a;
    outputs(1745) <= not (a or b);
    outputs(1746) <= a xor b;
    outputs(1747) <= not b;
    outputs(1748) <= a and b;
    outputs(1749) <= not (a xor b);
    outputs(1750) <= a xor b;
    outputs(1751) <= not a or b;
    outputs(1752) <= a xor b;
    outputs(1753) <= a xor b;
    outputs(1754) <= a and not b;
    outputs(1755) <= b;
    outputs(1756) <= b;
    outputs(1757) <= not (a xor b);
    outputs(1758) <= not b;
    outputs(1759) <= not a;
    outputs(1760) <= not a;
    outputs(1761) <= b and not a;
    outputs(1762) <= not (a xor b);
    outputs(1763) <= a xor b;
    outputs(1764) <= a;
    outputs(1765) <= b;
    outputs(1766) <= not b;
    outputs(1767) <= not (a or b);
    outputs(1768) <= a xor b;
    outputs(1769) <= not (a xor b);
    outputs(1770) <= a and not b;
    outputs(1771) <= a and not b;
    outputs(1772) <= not a;
    outputs(1773) <= a;
    outputs(1774) <= a and not b;
    outputs(1775) <= a and not b;
    outputs(1776) <= b and not a;
    outputs(1777) <= not a;
    outputs(1778) <= a xor b;
    outputs(1779) <= not (a or b);
    outputs(1780) <= a and not b;
    outputs(1781) <= b and not a;
    outputs(1782) <= not a;
    outputs(1783) <= not a;
    outputs(1784) <= a xor b;
    outputs(1785) <= not b;
    outputs(1786) <= a and not b;
    outputs(1787) <= not b;
    outputs(1788) <= b and not a;
    outputs(1789) <= b;
    outputs(1790) <= a and b;
    outputs(1791) <= not b;
    outputs(1792) <= a xor b;
    outputs(1793) <= not (a xor b);
    outputs(1794) <= not (a or b);
    outputs(1795) <= a xor b;
    outputs(1796) <= a and not b;
    outputs(1797) <= not (a xor b);
    outputs(1798) <= b and not a;
    outputs(1799) <= not (a xor b);
    outputs(1800) <= not a;
    outputs(1801) <= a xor b;
    outputs(1802) <= b and not a;
    outputs(1803) <= '0';
    outputs(1804) <= not a;
    outputs(1805) <= a and not b;
    outputs(1806) <= not (a xor b);
    outputs(1807) <= not (a xor b);
    outputs(1808) <= not (a or b);
    outputs(1809) <= not (a xor b);
    outputs(1810) <= b and not a;
    outputs(1811) <= not a;
    outputs(1812) <= a and not b;
    outputs(1813) <= not (a xor b);
    outputs(1814) <= not b;
    outputs(1815) <= not (a xor b);
    outputs(1816) <= b and not a;
    outputs(1817) <= a and b;
    outputs(1818) <= a and b;
    outputs(1819) <= not (a xor b);
    outputs(1820) <= a and not b;
    outputs(1821) <= a and b;
    outputs(1822) <= not (a xor b);
    outputs(1823) <= a xor b;
    outputs(1824) <= '0';
    outputs(1825) <= a and not b;
    outputs(1826) <= not (a xor b);
    outputs(1827) <= a and not b;
    outputs(1828) <= not (a xor b);
    outputs(1829) <= a;
    outputs(1830) <= not (a or b);
    outputs(1831) <= not a;
    outputs(1832) <= b;
    outputs(1833) <= b;
    outputs(1834) <= a xor b;
    outputs(1835) <= a;
    outputs(1836) <= not (a xor b);
    outputs(1837) <= not b;
    outputs(1838) <= b and not a;
    outputs(1839) <= not a;
    outputs(1840) <= b and not a;
    outputs(1841) <= a and b;
    outputs(1842) <= a and not b;
    outputs(1843) <= not (a or b);
    outputs(1844) <= not (a xor b);
    outputs(1845) <= a;
    outputs(1846) <= a and b;
    outputs(1847) <= not (a or b);
    outputs(1848) <= not (a xor b);
    outputs(1849) <= a xor b;
    outputs(1850) <= a and b;
    outputs(1851) <= not (a xor b);
    outputs(1852) <= a xor b;
    outputs(1853) <= not (a or b);
    outputs(1854) <= a and not b;
    outputs(1855) <= not b;
    outputs(1856) <= not (a xor b);
    outputs(1857) <= not (a xor b);
    outputs(1858) <= a and not b;
    outputs(1859) <= not (a xor b);
    outputs(1860) <= a xor b;
    outputs(1861) <= not b;
    outputs(1862) <= a and b;
    outputs(1863) <= not b;
    outputs(1864) <= not b;
    outputs(1865) <= b and not a;
    outputs(1866) <= not (a xor b);
    outputs(1867) <= b and not a;
    outputs(1868) <= a and not b;
    outputs(1869) <= a xor b;
    outputs(1870) <= not a;
    outputs(1871) <= not b;
    outputs(1872) <= a xor b;
    outputs(1873) <= not (a or b);
    outputs(1874) <= not (a or b);
    outputs(1875) <= b and not a;
    outputs(1876) <= not (a xor b);
    outputs(1877) <= not a;
    outputs(1878) <= not (a or b);
    outputs(1879) <= a;
    outputs(1880) <= not (a or b);
    outputs(1881) <= a xor b;
    outputs(1882) <= a xor b;
    outputs(1883) <= a;
    outputs(1884) <= not (a xor b);
    outputs(1885) <= not b;
    outputs(1886) <= not (a and b);
    outputs(1887) <= a and not b;
    outputs(1888) <= a xor b;
    outputs(1889) <= a and b;
    outputs(1890) <= a;
    outputs(1891) <= a;
    outputs(1892) <= a xor b;
    outputs(1893) <= b and not a;
    outputs(1894) <= not (a or b);
    outputs(1895) <= a and not b;
    outputs(1896) <= b;
    outputs(1897) <= not (a or b);
    outputs(1898) <= not (a xor b);
    outputs(1899) <= b;
    outputs(1900) <= not (a or b);
    outputs(1901) <= not a;
    outputs(1902) <= a xor b;
    outputs(1903) <= a and not b;
    outputs(1904) <= a and b;
    outputs(1905) <= b;
    outputs(1906) <= a xor b;
    outputs(1907) <= a and not b;
    outputs(1908) <= b and not a;
    outputs(1909) <= a and b;
    outputs(1910) <= a xor b;
    outputs(1911) <= not (a xor b);
    outputs(1912) <= a xor b;
    outputs(1913) <= a and b;
    outputs(1914) <= not b;
    outputs(1915) <= a xor b;
    outputs(1916) <= not (a xor b);
    outputs(1917) <= a xor b;
    outputs(1918) <= '0';
    outputs(1919) <= not (a xor b);
    outputs(1920) <= b;
    outputs(1921) <= not (a xor b);
    outputs(1922) <= a xor b;
    outputs(1923) <= not (a xor b);
    outputs(1924) <= not b;
    outputs(1925) <= a;
    outputs(1926) <= not a;
    outputs(1927) <= a and not b;
    outputs(1928) <= not (a xor b);
    outputs(1929) <= a and b;
    outputs(1930) <= not b;
    outputs(1931) <= b and not a;
    outputs(1932) <= not (a or b);
    outputs(1933) <= not b or a;
    outputs(1934) <= not b;
    outputs(1935) <= not b;
    outputs(1936) <= b and not a;
    outputs(1937) <= not a;
    outputs(1938) <= a;
    outputs(1939) <= not (a or b);
    outputs(1940) <= a and b;
    outputs(1941) <= b;
    outputs(1942) <= b;
    outputs(1943) <= a and not b;
    outputs(1944) <= not (a xor b);
    outputs(1945) <= b;
    outputs(1946) <= a and b;
    outputs(1947) <= not (a xor b);
    outputs(1948) <= not a;
    outputs(1949) <= b and not a;
    outputs(1950) <= not (a xor b);
    outputs(1951) <= b;
    outputs(1952) <= a and b;
    outputs(1953) <= a and b;
    outputs(1954) <= not a;
    outputs(1955) <= b and not a;
    outputs(1956) <= not (a xor b);
    outputs(1957) <= a xor b;
    outputs(1958) <= a and b;
    outputs(1959) <= a xor b;
    outputs(1960) <= a and not b;
    outputs(1961) <= not a;
    outputs(1962) <= a and b;
    outputs(1963) <= not (a or b);
    outputs(1964) <= a xor b;
    outputs(1965) <= not a;
    outputs(1966) <= not (a or b);
    outputs(1967) <= not b;
    outputs(1968) <= b and not a;
    outputs(1969) <= not a;
    outputs(1970) <= a xor b;
    outputs(1971) <= a and b;
    outputs(1972) <= a xor b;
    outputs(1973) <= b and not a;
    outputs(1974) <= a;
    outputs(1975) <= not (a xor b);
    outputs(1976) <= not (a or b);
    outputs(1977) <= not (a xor b);
    outputs(1978) <= not a or b;
    outputs(1979) <= b;
    outputs(1980) <= not (a or b);
    outputs(1981) <= not (a xor b);
    outputs(1982) <= '0';
    outputs(1983) <= not b;
    outputs(1984) <= a xor b;
    outputs(1985) <= b;
    outputs(1986) <= a;
    outputs(1987) <= a and not b;
    outputs(1988) <= not (a xor b);
    outputs(1989) <= not (a xor b);
    outputs(1990) <= b and not a;
    outputs(1991) <= not (a or b);
    outputs(1992) <= a xor b;
    outputs(1993) <= not (a xor b);
    outputs(1994) <= a and not b;
    outputs(1995) <= b;
    outputs(1996) <= not (a or b);
    outputs(1997) <= not b;
    outputs(1998) <= b and not a;
    outputs(1999) <= not a;
    outputs(2000) <= not (a or b);
    outputs(2001) <= not (a or b);
    outputs(2002) <= a or b;
    outputs(2003) <= a;
    outputs(2004) <= a xor b;
    outputs(2005) <= not (a xor b);
    outputs(2006) <= not (a xor b);
    outputs(2007) <= not a;
    outputs(2008) <= b and not a;
    outputs(2009) <= a xor b;
    outputs(2010) <= a and not b;
    outputs(2011) <= not a;
    outputs(2012) <= a;
    outputs(2013) <= a;
    outputs(2014) <= '0';
    outputs(2015) <= a and not b;
    outputs(2016) <= not (a xor b);
    outputs(2017) <= b and not a;
    outputs(2018) <= a and not b;
    outputs(2019) <= not (a or b);
    outputs(2020) <= b;
    outputs(2021) <= b;
    outputs(2022) <= a and b;
    outputs(2023) <= a and b;
    outputs(2024) <= a xor b;
    outputs(2025) <= not (a xor b);
    outputs(2026) <= a xor b;
    outputs(2027) <= a and not b;
    outputs(2028) <= not b;
    outputs(2029) <= a and not b;
    outputs(2030) <= not (a xor b);
    outputs(2031) <= not b;
    outputs(2032) <= b;
    outputs(2033) <= a and b;
    outputs(2034) <= a and not b;
    outputs(2035) <= b;
    outputs(2036) <= not (a xor b);
    outputs(2037) <= b;
    outputs(2038) <= not (a xor b);
    outputs(2039) <= b;
    outputs(2040) <= not b;
    outputs(2041) <= b;
    outputs(2042) <= a xor b;
    outputs(2043) <= not (a xor b);
    outputs(2044) <= not (a xor b);
    outputs(2045) <= a;
    outputs(2046) <= b and not a;
    outputs(2047) <= a;
    outputs(2048) <= b;
    outputs(2049) <= a or b;
    outputs(2050) <= not b;
    outputs(2051) <= b;
    outputs(2052) <= not a;
    outputs(2053) <= a xor b;
    outputs(2054) <= a xor b;
    outputs(2055) <= not (a xor b);
    outputs(2056) <= b and not a;
    outputs(2057) <= a and b;
    outputs(2058) <= not (a xor b);
    outputs(2059) <= not a or b;
    outputs(2060) <= not a or b;
    outputs(2061) <= not (a xor b);
    outputs(2062) <= a or b;
    outputs(2063) <= a xor b;
    outputs(2064) <= a xor b;
    outputs(2065) <= not b or a;
    outputs(2066) <= not b;
    outputs(2067) <= not a;
    outputs(2068) <= not (a xor b);
    outputs(2069) <= not (a and b);
    outputs(2070) <= not a;
    outputs(2071) <= a;
    outputs(2072) <= a xor b;
    outputs(2073) <= b;
    outputs(2074) <= a;
    outputs(2075) <= a xor b;
    outputs(2076) <= not b;
    outputs(2077) <= not a;
    outputs(2078) <= a;
    outputs(2079) <= not a;
    outputs(2080) <= not (a xor b);
    outputs(2081) <= not b;
    outputs(2082) <= not a;
    outputs(2083) <= not (a xor b);
    outputs(2084) <= b;
    outputs(2085) <= not b or a;
    outputs(2086) <= not (a or b);
    outputs(2087) <= b;
    outputs(2088) <= not a;
    outputs(2089) <= a;
    outputs(2090) <= not a;
    outputs(2091) <= a and not b;
    outputs(2092) <= a;
    outputs(2093) <= not b;
    outputs(2094) <= not b;
    outputs(2095) <= not (a xor b);
    outputs(2096) <= b;
    outputs(2097) <= not b;
    outputs(2098) <= a;
    outputs(2099) <= not a or b;
    outputs(2100) <= not b;
    outputs(2101) <= a xor b;
    outputs(2102) <= a and b;
    outputs(2103) <= b;
    outputs(2104) <= not a;
    outputs(2105) <= a and b;
    outputs(2106) <= not b;
    outputs(2107) <= a;
    outputs(2108) <= not a;
    outputs(2109) <= not a;
    outputs(2110) <= not (a or b);
    outputs(2111) <= not (a and b);
    outputs(2112) <= a;
    outputs(2113) <= not (a xor b);
    outputs(2114) <= b and not a;
    outputs(2115) <= not (a xor b);
    outputs(2116) <= b and not a;
    outputs(2117) <= b;
    outputs(2118) <= a xor b;
    outputs(2119) <= not b or a;
    outputs(2120) <= not (a xor b);
    outputs(2121) <= a;
    outputs(2122) <= a;
    outputs(2123) <= a xor b;
    outputs(2124) <= a;
    outputs(2125) <= not (a xor b);
    outputs(2126) <= not (a and b);
    outputs(2127) <= a xor b;
    outputs(2128) <= not a or b;
    outputs(2129) <= a xor b;
    outputs(2130) <= a and not b;
    outputs(2131) <= not a;
    outputs(2132) <= b and not a;
    outputs(2133) <= not (a xor b);
    outputs(2134) <= a xor b;
    outputs(2135) <= not a or b;
    outputs(2136) <= a;
    outputs(2137) <= a xor b;
    outputs(2138) <= not (a or b);
    outputs(2139) <= not (a xor b);
    outputs(2140) <= not (a xor b);
    outputs(2141) <= a xor b;
    outputs(2142) <= not a;
    outputs(2143) <= b;
    outputs(2144) <= b and not a;
    outputs(2145) <= b;
    outputs(2146) <= not (a xor b);
    outputs(2147) <= not a;
    outputs(2148) <= b;
    outputs(2149) <= a xor b;
    outputs(2150) <= a xor b;
    outputs(2151) <= not b;
    outputs(2152) <= not b;
    outputs(2153) <= not a or b;
    outputs(2154) <= not a;
    outputs(2155) <= a or b;
    outputs(2156) <= not (a xor b);
    outputs(2157) <= not (a xor b);
    outputs(2158) <= not b;
    outputs(2159) <= not (a xor b);
    outputs(2160) <= b;
    outputs(2161) <= a;
    outputs(2162) <= not (a xor b);
    outputs(2163) <= a xor b;
    outputs(2164) <= not (a or b);
    outputs(2165) <= not a or b;
    outputs(2166) <= not a;
    outputs(2167) <= a xor b;
    outputs(2168) <= not b or a;
    outputs(2169) <= a and not b;
    outputs(2170) <= a or b;
    outputs(2171) <= a xor b;
    outputs(2172) <= a;
    outputs(2173) <= not (a or b);
    outputs(2174) <= a;
    outputs(2175) <= a or b;
    outputs(2176) <= not b;
    outputs(2177) <= a and b;
    outputs(2178) <= a or b;
    outputs(2179) <= not (a or b);
    outputs(2180) <= a xor b;
    outputs(2181) <= a and b;
    outputs(2182) <= b;
    outputs(2183) <= not b;
    outputs(2184) <= not a;
    outputs(2185) <= not a;
    outputs(2186) <= a and b;
    outputs(2187) <= a;
    outputs(2188) <= a xor b;
    outputs(2189) <= not a;
    outputs(2190) <= b;
    outputs(2191) <= not a;
    outputs(2192) <= a;
    outputs(2193) <= not (a xor b);
    outputs(2194) <= not (a xor b);
    outputs(2195) <= a;
    outputs(2196) <= a xor b;
    outputs(2197) <= not a;
    outputs(2198) <= b and not a;
    outputs(2199) <= a and not b;
    outputs(2200) <= not b or a;
    outputs(2201) <= a xor b;
    outputs(2202) <= b;
    outputs(2203) <= b and not a;
    outputs(2204) <= a xor b;
    outputs(2205) <= not (a xor b);
    outputs(2206) <= not a or b;
    outputs(2207) <= not (a xor b);
    outputs(2208) <= not b or a;
    outputs(2209) <= not (a xor b);
    outputs(2210) <= b;
    outputs(2211) <= a or b;
    outputs(2212) <= not (a xor b);
    outputs(2213) <= a xor b;
    outputs(2214) <= a;
    outputs(2215) <= not a;
    outputs(2216) <= a or b;
    outputs(2217) <= a xor b;
    outputs(2218) <= a xor b;
    outputs(2219) <= b;
    outputs(2220) <= not (a xor b);
    outputs(2221) <= not a or b;
    outputs(2222) <= b;
    outputs(2223) <= b;
    outputs(2224) <= a xor b;
    outputs(2225) <= not (a xor b);
    outputs(2226) <= a xor b;
    outputs(2227) <= not a or b;
    outputs(2228) <= not (a and b);
    outputs(2229) <= not a or b;
    outputs(2230) <= b;
    outputs(2231) <= not a or b;
    outputs(2232) <= not a or b;
    outputs(2233) <= a xor b;
    outputs(2234) <= a xor b;
    outputs(2235) <= not (a xor b);
    outputs(2236) <= not b or a;
    outputs(2237) <= not (a and b);
    outputs(2238) <= not a or b;
    outputs(2239) <= b;
    outputs(2240) <= b and not a;
    outputs(2241) <= not (a xor b);
    outputs(2242) <= a;
    outputs(2243) <= not (a or b);
    outputs(2244) <= b;
    outputs(2245) <= not (a xor b);
    outputs(2246) <= not b;
    outputs(2247) <= not (a and b);
    outputs(2248) <= b;
    outputs(2249) <= a xor b;
    outputs(2250) <= a;
    outputs(2251) <= not a;
    outputs(2252) <= not (a xor b);
    outputs(2253) <= a xor b;
    outputs(2254) <= a xor b;
    outputs(2255) <= a;
    outputs(2256) <= not (a or b);
    outputs(2257) <= b;
    outputs(2258) <= not (a and b);
    outputs(2259) <= a;
    outputs(2260) <= a or b;
    outputs(2261) <= a xor b;
    outputs(2262) <= not a;
    outputs(2263) <= a xor b;
    outputs(2264) <= a xor b;
    outputs(2265) <= a and b;
    outputs(2266) <= b;
    outputs(2267) <= a xor b;
    outputs(2268) <= not (a xor b);
    outputs(2269) <= not a or b;
    outputs(2270) <= not (a xor b);
    outputs(2271) <= a xor b;
    outputs(2272) <= not a or b;
    outputs(2273) <= not (a and b);
    outputs(2274) <= a;
    outputs(2275) <= not (a xor b);
    outputs(2276) <= b;
    outputs(2277) <= not a;
    outputs(2278) <= b;
    outputs(2279) <= not a;
    outputs(2280) <= not a;
    outputs(2281) <= not b or a;
    outputs(2282) <= not a;
    outputs(2283) <= a xor b;
    outputs(2284) <= not a;
    outputs(2285) <= a;
    outputs(2286) <= not (a and b);
    outputs(2287) <= a xor b;
    outputs(2288) <= a and not b;
    outputs(2289) <= not (a xor b);
    outputs(2290) <= a xor b;
    outputs(2291) <= a;
    outputs(2292) <= not (a xor b);
    outputs(2293) <= not (a xor b);
    outputs(2294) <= not (a xor b);
    outputs(2295) <= a xor b;
    outputs(2296) <= a xor b;
    outputs(2297) <= a xor b;
    outputs(2298) <= not (a and b);
    outputs(2299) <= not b or a;
    outputs(2300) <= not a or b;
    outputs(2301) <= not (a xor b);
    outputs(2302) <= not (a xor b);
    outputs(2303) <= a xor b;
    outputs(2304) <= not a;
    outputs(2305) <= not a or b;
    outputs(2306) <= not a;
    outputs(2307) <= a or b;
    outputs(2308) <= not b;
    outputs(2309) <= b;
    outputs(2310) <= not (a xor b);
    outputs(2311) <= b;
    outputs(2312) <= a and not b;
    outputs(2313) <= not (a and b);
    outputs(2314) <= a;
    outputs(2315) <= not (a or b);
    outputs(2316) <= not b;
    outputs(2317) <= a xor b;
    outputs(2318) <= b and not a;
    outputs(2319) <= not b or a;
    outputs(2320) <= a xor b;
    outputs(2321) <= a and not b;
    outputs(2322) <= not a;
    outputs(2323) <= b;
    outputs(2324) <= not (a and b);
    outputs(2325) <= not b;
    outputs(2326) <= a;
    outputs(2327) <= not b;
    outputs(2328) <= a;
    outputs(2329) <= not a;
    outputs(2330) <= b;
    outputs(2331) <= not (a xor b);
    outputs(2332) <= not a;
    outputs(2333) <= a xor b;
    outputs(2334) <= b;
    outputs(2335) <= not b or a;
    outputs(2336) <= not b;
    outputs(2337) <= not b;
    outputs(2338) <= not a or b;
    outputs(2339) <= a xor b;
    outputs(2340) <= b;
    outputs(2341) <= not a;
    outputs(2342) <= not (a xor b);
    outputs(2343) <= a xor b;
    outputs(2344) <= not a;
    outputs(2345) <= a and not b;
    outputs(2346) <= a;
    outputs(2347) <= not (a and b);
    outputs(2348) <= b;
    outputs(2349) <= a or b;
    outputs(2350) <= not a;
    outputs(2351) <= not (a and b);
    outputs(2352) <= b;
    outputs(2353) <= not b;
    outputs(2354) <= not (a xor b);
    outputs(2355) <= not b;
    outputs(2356) <= b;
    outputs(2357) <= a and not b;
    outputs(2358) <= a or b;
    outputs(2359) <= a;
    outputs(2360) <= b;
    outputs(2361) <= a;
    outputs(2362) <= b;
    outputs(2363) <= a;
    outputs(2364) <= not b or a;
    outputs(2365) <= a xor b;
    outputs(2366) <= a xor b;
    outputs(2367) <= a or b;
    outputs(2368) <= a and not b;
    outputs(2369) <= b;
    outputs(2370) <= not (a and b);
    outputs(2371) <= not (a or b);
    outputs(2372) <= a;
    outputs(2373) <= not (a xor b);
    outputs(2374) <= a xor b;
    outputs(2375) <= not a;
    outputs(2376) <= a xor b;
    outputs(2377) <= b;
    outputs(2378) <= a;
    outputs(2379) <= a xor b;
    outputs(2380) <= not (a or b);
    outputs(2381) <= a or b;
    outputs(2382) <= not (a xor b);
    outputs(2383) <= a xor b;
    outputs(2384) <= a;
    outputs(2385) <= a xor b;
    outputs(2386) <= a xor b;
    outputs(2387) <= not (a xor b);
    outputs(2388) <= not (a xor b);
    outputs(2389) <= a or b;
    outputs(2390) <= not a;
    outputs(2391) <= a;
    outputs(2392) <= not (a xor b);
    outputs(2393) <= not (a and b);
    outputs(2394) <= not (a xor b);
    outputs(2395) <= a;
    outputs(2396) <= a;
    outputs(2397) <= not a;
    outputs(2398) <= b;
    outputs(2399) <= not a;
    outputs(2400) <= a xor b;
    outputs(2401) <= not b;
    outputs(2402) <= a or b;
    outputs(2403) <= a xor b;
    outputs(2404) <= b and not a;
    outputs(2405) <= not (a or b);
    outputs(2406) <= not b;
    outputs(2407) <= b;
    outputs(2408) <= a xor b;
    outputs(2409) <= b;
    outputs(2410) <= b;
    outputs(2411) <= a;
    outputs(2412) <= not b or a;
    outputs(2413) <= not a;
    outputs(2414) <= not a;
    outputs(2415) <= a and not b;
    outputs(2416) <= not b;
    outputs(2417) <= not b;
    outputs(2418) <= not b;
    outputs(2419) <= a xor b;
    outputs(2420) <= not (a and b);
    outputs(2421) <= a and not b;
    outputs(2422) <= a and b;
    outputs(2423) <= a;
    outputs(2424) <= not (a xor b);
    outputs(2425) <= b and not a;
    outputs(2426) <= b;
    outputs(2427) <= not (a xor b);
    outputs(2428) <= not a or b;
    outputs(2429) <= a and not b;
    outputs(2430) <= not a or b;
    outputs(2431) <= not a;
    outputs(2432) <= a or b;
    outputs(2433) <= not (a and b);
    outputs(2434) <= not b;
    outputs(2435) <= not a;
    outputs(2436) <= not a;
    outputs(2437) <= not (a xor b);
    outputs(2438) <= a xor b;
    outputs(2439) <= not (a xor b);
    outputs(2440) <= not b or a;
    outputs(2441) <= not a;
    outputs(2442) <= not b;
    outputs(2443) <= not a;
    outputs(2444) <= not (a or b);
    outputs(2445) <= not (a or b);
    outputs(2446) <= a xor b;
    outputs(2447) <= not a;
    outputs(2448) <= a;
    outputs(2449) <= a;
    outputs(2450) <= not (a xor b);
    outputs(2451) <= not b;
    outputs(2452) <= not (a xor b);
    outputs(2453) <= a;
    outputs(2454) <= b;
    outputs(2455) <= b;
    outputs(2456) <= b and not a;
    outputs(2457) <= a or b;
    outputs(2458) <= a;
    outputs(2459) <= not b or a;
    outputs(2460) <= not a;
    outputs(2461) <= not a or b;
    outputs(2462) <= not (a xor b);
    outputs(2463) <= a or b;
    outputs(2464) <= a xor b;
    outputs(2465) <= a;
    outputs(2466) <= not b or a;
    outputs(2467) <= a or b;
    outputs(2468) <= not (a xor b);
    outputs(2469) <= b and not a;
    outputs(2470) <= not (a xor b);
    outputs(2471) <= b;
    outputs(2472) <= not (a xor b);
    outputs(2473) <= not (a or b);
    outputs(2474) <= not (a and b);
    outputs(2475) <= a and not b;
    outputs(2476) <= not (a xor b);
    outputs(2477) <= not (a or b);
    outputs(2478) <= not a;
    outputs(2479) <= a and not b;
    outputs(2480) <= a xor b;
    outputs(2481) <= not b;
    outputs(2482) <= a xor b;
    outputs(2483) <= a xor b;
    outputs(2484) <= not b;
    outputs(2485) <= not (a xor b);
    outputs(2486) <= not b or a;
    outputs(2487) <= b;
    outputs(2488) <= b;
    outputs(2489) <= not b;
    outputs(2490) <= not a;
    outputs(2491) <= not a or b;
    outputs(2492) <= a xor b;
    outputs(2493) <= not (a xor b);
    outputs(2494) <= not b or a;
    outputs(2495) <= not (a and b);
    outputs(2496) <= not (a and b);
    outputs(2497) <= not (a xor b);
    outputs(2498) <= not (a or b);
    outputs(2499) <= a or b;
    outputs(2500) <= a or b;
    outputs(2501) <= not a;
    outputs(2502) <= a;
    outputs(2503) <= a xor b;
    outputs(2504) <= not a or b;
    outputs(2505) <= not (a xor b);
    outputs(2506) <= not (a or b);
    outputs(2507) <= not (a xor b);
    outputs(2508) <= not b;
    outputs(2509) <= a xor b;
    outputs(2510) <= not (a xor b);
    outputs(2511) <= a xor b;
    outputs(2512) <= a and not b;
    outputs(2513) <= not b;
    outputs(2514) <= a and not b;
    outputs(2515) <= a and b;
    outputs(2516) <= a xor b;
    outputs(2517) <= not (a xor b);
    outputs(2518) <= a xor b;
    outputs(2519) <= not (a xor b);
    outputs(2520) <= a;
    outputs(2521) <= not (a and b);
    outputs(2522) <= not b;
    outputs(2523) <= not (a xor b);
    outputs(2524) <= not a;
    outputs(2525) <= a;
    outputs(2526) <= b;
    outputs(2527) <= a;
    outputs(2528) <= a or b;
    outputs(2529) <= b;
    outputs(2530) <= a xor b;
    outputs(2531) <= a and not b;
    outputs(2532) <= a;
    outputs(2533) <= not b or a;
    outputs(2534) <= a and not b;
    outputs(2535) <= not b;
    outputs(2536) <= a and not b;
    outputs(2537) <= not (a or b);
    outputs(2538) <= b;
    outputs(2539) <= b;
    outputs(2540) <= not b;
    outputs(2541) <= a xor b;
    outputs(2542) <= not (a xor b);
    outputs(2543) <= not a;
    outputs(2544) <= b and not a;
    outputs(2545) <= a or b;
    outputs(2546) <= not a or b;
    outputs(2547) <= not b;
    outputs(2548) <= a and b;
    outputs(2549) <= not (a and b);
    outputs(2550) <= not b;
    outputs(2551) <= a xor b;
    outputs(2552) <= not a;
    outputs(2553) <= a xor b;
    outputs(2554) <= b;
    outputs(2555) <= not b;
    outputs(2556) <= not (a xor b);
    outputs(2557) <= b;
    outputs(2558) <= a and not b;
    outputs(2559) <= b;
    outputs(2560) <= a and not b;
    outputs(2561) <= not a or b;
    outputs(2562) <= not (a or b);
    outputs(2563) <= a;
    outputs(2564) <= not (a xor b);
    outputs(2565) <= not a;
    outputs(2566) <= not a;
    outputs(2567) <= not (a or b);
    outputs(2568) <= b;
    outputs(2569) <= b;
    outputs(2570) <= not a;
    outputs(2571) <= b and not a;
    outputs(2572) <= a xor b;
    outputs(2573) <= a xor b;
    outputs(2574) <= not (a or b);
    outputs(2575) <= not (a xor b);
    outputs(2576) <= a and not b;
    outputs(2577) <= a and b;
    outputs(2578) <= a xor b;
    outputs(2579) <= a;
    outputs(2580) <= not (a xor b);
    outputs(2581) <= a;
    outputs(2582) <= not (a xor b);
    outputs(2583) <= not (a xor b);
    outputs(2584) <= not (a xor b);
    outputs(2585) <= b;
    outputs(2586) <= a;
    outputs(2587) <= not b;
    outputs(2588) <= a xor b;
    outputs(2589) <= a;
    outputs(2590) <= a xor b;
    outputs(2591) <= not a;
    outputs(2592) <= not a;
    outputs(2593) <= not a;
    outputs(2594) <= not a;
    outputs(2595) <= not a;
    outputs(2596) <= a;
    outputs(2597) <= not (a or b);
    outputs(2598) <= not (a xor b);
    outputs(2599) <= not a or b;
    outputs(2600) <= not a;
    outputs(2601) <= not a;
    outputs(2602) <= not (a or b);
    outputs(2603) <= not b;
    outputs(2604) <= not b;
    outputs(2605) <= a;
    outputs(2606) <= a;
    outputs(2607) <= not (a and b);
    outputs(2608) <= a;
    outputs(2609) <= not a;
    outputs(2610) <= b;
    outputs(2611) <= not (a xor b);
    outputs(2612) <= a xor b;
    outputs(2613) <= not (a xor b);
    outputs(2614) <= a xor b;
    outputs(2615) <= not b;
    outputs(2616) <= a xor b;
    outputs(2617) <= a or b;
    outputs(2618) <= a;
    outputs(2619) <= not (a or b);
    outputs(2620) <= a and not b;
    outputs(2621) <= not b or a;
    outputs(2622) <= a;
    outputs(2623) <= not (a xor b);
    outputs(2624) <= not b;
    outputs(2625) <= b and not a;
    outputs(2626) <= not a or b;
    outputs(2627) <= not a;
    outputs(2628) <= a xor b;
    outputs(2629) <= a;
    outputs(2630) <= a xor b;
    outputs(2631) <= not a;
    outputs(2632) <= not (a xor b);
    outputs(2633) <= a;
    outputs(2634) <= not (a and b);
    outputs(2635) <= not a or b;
    outputs(2636) <= b;
    outputs(2637) <= not a or b;
    outputs(2638) <= not (a or b);
    outputs(2639) <= not a;
    outputs(2640) <= not (a or b);
    outputs(2641) <= not (a xor b);
    outputs(2642) <= b;
    outputs(2643) <= b;
    outputs(2644) <= a xor b;
    outputs(2645) <= b;
    outputs(2646) <= not b or a;
    outputs(2647) <= not b;
    outputs(2648) <= not b or a;
    outputs(2649) <= not a;
    outputs(2650) <= not (a xor b);
    outputs(2651) <= not a;
    outputs(2652) <= a and b;
    outputs(2653) <= a;
    outputs(2654) <= a xor b;
    outputs(2655) <= not a;
    outputs(2656) <= a xor b;
    outputs(2657) <= a xor b;
    outputs(2658) <= not a;
    outputs(2659) <= not (a or b);
    outputs(2660) <= not a;
    outputs(2661) <= not (a xor b);
    outputs(2662) <= not a;
    outputs(2663) <= not b;
    outputs(2664) <= b;
    outputs(2665) <= not (a and b);
    outputs(2666) <= b and not a;
    outputs(2667) <= not a or b;
    outputs(2668) <= not a;
    outputs(2669) <= not (a xor b);
    outputs(2670) <= not (a xor b);
    outputs(2671) <= a xor b;
    outputs(2672) <= b;
    outputs(2673) <= b;
    outputs(2674) <= a;
    outputs(2675) <= a xor b;
    outputs(2676) <= b;
    outputs(2677) <= not b;
    outputs(2678) <= a xor b;
    outputs(2679) <= a xor b;
    outputs(2680) <= a xor b;
    outputs(2681) <= a and b;
    outputs(2682) <= not (a xor b);
    outputs(2683) <= a;
    outputs(2684) <= not a or b;
    outputs(2685) <= not (a xor b);
    outputs(2686) <= b;
    outputs(2687) <= not (a or b);
    outputs(2688) <= not (a xor b);
    outputs(2689) <= not b;
    outputs(2690) <= not (a and b);
    outputs(2691) <= b and not a;
    outputs(2692) <= a xor b;
    outputs(2693) <= not a;
    outputs(2694) <= b;
    outputs(2695) <= not a;
    outputs(2696) <= not b or a;
    outputs(2697) <= not a;
    outputs(2698) <= b;
    outputs(2699) <= not b;
    outputs(2700) <= not b;
    outputs(2701) <= b;
    outputs(2702) <= a xor b;
    outputs(2703) <= not a or b;
    outputs(2704) <= a xor b;
    outputs(2705) <= not a or b;
    outputs(2706) <= not a or b;
    outputs(2707) <= a xor b;
    outputs(2708) <= b;
    outputs(2709) <= not (a and b);
    outputs(2710) <= not a;
    outputs(2711) <= not b;
    outputs(2712) <= not b;
    outputs(2713) <= not b;
    outputs(2714) <= not (a xor b);
    outputs(2715) <= not a or b;
    outputs(2716) <= a and not b;
    outputs(2717) <= a or b;
    outputs(2718) <= a and not b;
    outputs(2719) <= not b or a;
    outputs(2720) <= a and not b;
    outputs(2721) <= a;
    outputs(2722) <= a or b;
    outputs(2723) <= a;
    outputs(2724) <= not (a xor b);
    outputs(2725) <= b and not a;
    outputs(2726) <= b and not a;
    outputs(2727) <= not (a and b);
    outputs(2728) <= a xor b;
    outputs(2729) <= a xor b;
    outputs(2730) <= b;
    outputs(2731) <= b;
    outputs(2732) <= b;
    outputs(2733) <= not (a or b);
    outputs(2734) <= not (a xor b);
    outputs(2735) <= not a;
    outputs(2736) <= not a;
    outputs(2737) <= not a;
    outputs(2738) <= not a or b;
    outputs(2739) <= not b;
    outputs(2740) <= not (a or b);
    outputs(2741) <= not a;
    outputs(2742) <= not (a and b);
    outputs(2743) <= not b;
    outputs(2744) <= a xor b;
    outputs(2745) <= a or b;
    outputs(2746) <= a;
    outputs(2747) <= not (a xor b);
    outputs(2748) <= a xor b;
    outputs(2749) <= a xor b;
    outputs(2750) <= not b;
    outputs(2751) <= a and not b;
    outputs(2752) <= a and not b;
    outputs(2753) <= not a;
    outputs(2754) <= not b;
    outputs(2755) <= a or b;
    outputs(2756) <= not (a or b);
    outputs(2757) <= a xor b;
    outputs(2758) <= not b or a;
    outputs(2759) <= a;
    outputs(2760) <= not (a xor b);
    outputs(2761) <= not a or b;
    outputs(2762) <= a xor b;
    outputs(2763) <= a xor b;
    outputs(2764) <= a;
    outputs(2765) <= a;
    outputs(2766) <= not b;
    outputs(2767) <= not a;
    outputs(2768) <= not a or b;
    outputs(2769) <= a;
    outputs(2770) <= not b;
    outputs(2771) <= not (a xor b);
    outputs(2772) <= not b;
    outputs(2773) <= a;
    outputs(2774) <= a or b;
    outputs(2775) <= not a;
    outputs(2776) <= a;
    outputs(2777) <= b;
    outputs(2778) <= not (a and b);
    outputs(2779) <= b;
    outputs(2780) <= not b;
    outputs(2781) <= a or b;
    outputs(2782) <= b;
    outputs(2783) <= a and not b;
    outputs(2784) <= not a;
    outputs(2785) <= b;
    outputs(2786) <= not (a or b);
    outputs(2787) <= a;
    outputs(2788) <= a xor b;
    outputs(2789) <= not b or a;
    outputs(2790) <= a or b;
    outputs(2791) <= not (a xor b);
    outputs(2792) <= a;
    outputs(2793) <= b and not a;
    outputs(2794) <= b;
    outputs(2795) <= not a or b;
    outputs(2796) <= a or b;
    outputs(2797) <= not a or b;
    outputs(2798) <= a xor b;
    outputs(2799) <= a;
    outputs(2800) <= not (a xor b);
    outputs(2801) <= a;
    outputs(2802) <= a xor b;
    outputs(2803) <= not (a xor b);
    outputs(2804) <= b;
    outputs(2805) <= b and not a;
    outputs(2806) <= a;
    outputs(2807) <= not (a xor b);
    outputs(2808) <= a xor b;
    outputs(2809) <= a xor b;
    outputs(2810) <= not b;
    outputs(2811) <= not a or b;
    outputs(2812) <= not (a xor b);
    outputs(2813) <= a xor b;
    outputs(2814) <= a and b;
    outputs(2815) <= a xor b;
    outputs(2816) <= not b;
    outputs(2817) <= not b or a;
    outputs(2818) <= not a or b;
    outputs(2819) <= not (a xor b);
    outputs(2820) <= a xor b;
    outputs(2821) <= not b or a;
    outputs(2822) <= a;
    outputs(2823) <= not (a xor b);
    outputs(2824) <= b;
    outputs(2825) <= a and b;
    outputs(2826) <= not b;
    outputs(2827) <= not b or a;
    outputs(2828) <= a;
    outputs(2829) <= a xor b;
    outputs(2830) <= a and not b;
    outputs(2831) <= not a;
    outputs(2832) <= a and b;
    outputs(2833) <= a;
    outputs(2834) <= a;
    outputs(2835) <= a;
    outputs(2836) <= a xor b;
    outputs(2837) <= a xor b;
    outputs(2838) <= a xor b;
    outputs(2839) <= a xor b;
    outputs(2840) <= a and b;
    outputs(2841) <= not b;
    outputs(2842) <= a xor b;
    outputs(2843) <= not (a or b);
    outputs(2844) <= a and not b;
    outputs(2845) <= a xor b;
    outputs(2846) <= not (a xor b);
    outputs(2847) <= a;
    outputs(2848) <= a;
    outputs(2849) <= not (a and b);
    outputs(2850) <= not (a xor b);
    outputs(2851) <= b and not a;
    outputs(2852) <= a or b;
    outputs(2853) <= a xor b;
    outputs(2854) <= not (a xor b);
    outputs(2855) <= b;
    outputs(2856) <= not a;
    outputs(2857) <= not b;
    outputs(2858) <= a and not b;
    outputs(2859) <= not (a xor b);
    outputs(2860) <= not (a xor b);
    outputs(2861) <= a or b;
    outputs(2862) <= not a;
    outputs(2863) <= not (a xor b);
    outputs(2864) <= a;
    outputs(2865) <= a;
    outputs(2866) <= not (a and b);
    outputs(2867) <= not a;
    outputs(2868) <= not b;
    outputs(2869) <= a and b;
    outputs(2870) <= not a or b;
    outputs(2871) <= not a;
    outputs(2872) <= a xor b;
    outputs(2873) <= a and not b;
    outputs(2874) <= not (a xor b);
    outputs(2875) <= not a;
    outputs(2876) <= not a;
    outputs(2877) <= a xor b;
    outputs(2878) <= not (a xor b);
    outputs(2879) <= not b;
    outputs(2880) <= b;
    outputs(2881) <= not (a xor b);
    outputs(2882) <= b;
    outputs(2883) <= not (a or b);
    outputs(2884) <= a or b;
    outputs(2885) <= a xor b;
    outputs(2886) <= not (a xor b);
    outputs(2887) <= not b;
    outputs(2888) <= a;
    outputs(2889) <= not a;
    outputs(2890) <= not b;
    outputs(2891) <= b;
    outputs(2892) <= not b;
    outputs(2893) <= not (a xor b);
    outputs(2894) <= b;
    outputs(2895) <= a xor b;
    outputs(2896) <= b;
    outputs(2897) <= not (a xor b);
    outputs(2898) <= b;
    outputs(2899) <= not (a xor b);
    outputs(2900) <= not (a or b);
    outputs(2901) <= not b;
    outputs(2902) <= not (a xor b);
    outputs(2903) <= a or b;
    outputs(2904) <= not a;
    outputs(2905) <= a or b;
    outputs(2906) <= a xor b;
    outputs(2907) <= a xor b;
    outputs(2908) <= b;
    outputs(2909) <= not (a xor b);
    outputs(2910) <= not b;
    outputs(2911) <= b;
    outputs(2912) <= a;
    outputs(2913) <= not b;
    outputs(2914) <= not (a xor b);
    outputs(2915) <= a and b;
    outputs(2916) <= not (a or b);
    outputs(2917) <= a xor b;
    outputs(2918) <= b;
    outputs(2919) <= not (a xor b);
    outputs(2920) <= b;
    outputs(2921) <= b;
    outputs(2922) <= not a;
    outputs(2923) <= not b or a;
    outputs(2924) <= not b;
    outputs(2925) <= b;
    outputs(2926) <= not b;
    outputs(2927) <= not a;
    outputs(2928) <= a xor b;
    outputs(2929) <= a;
    outputs(2930) <= not a;
    outputs(2931) <= not (a xor b);
    outputs(2932) <= not (a or b);
    outputs(2933) <= a;
    outputs(2934) <= not b or a;
    outputs(2935) <= a xor b;
    outputs(2936) <= a;
    outputs(2937) <= not b or a;
    outputs(2938) <= b;
    outputs(2939) <= a;
    outputs(2940) <= not a;
    outputs(2941) <= a;
    outputs(2942) <= not (a xor b);
    outputs(2943) <= not a;
    outputs(2944) <= a or b;
    outputs(2945) <= not (a or b);
    outputs(2946) <= b;
    outputs(2947) <= a;
    outputs(2948) <= b and not a;
    outputs(2949) <= b;
    outputs(2950) <= not (a or b);
    outputs(2951) <= a xor b;
    outputs(2952) <= b;
    outputs(2953) <= not (a xor b);
    outputs(2954) <= not a;
    outputs(2955) <= not (a and b);
    outputs(2956) <= b and not a;
    outputs(2957) <= b;
    outputs(2958) <= a and b;
    outputs(2959) <= not (a xor b);
    outputs(2960) <= a;
    outputs(2961) <= not (a and b);
    outputs(2962) <= not (a xor b);
    outputs(2963) <= not (a xor b);
    outputs(2964) <= not b;
    outputs(2965) <= not b or a;
    outputs(2966) <= not (a or b);
    outputs(2967) <= b and not a;
    outputs(2968) <= b;
    outputs(2969) <= b;
    outputs(2970) <= not (a xor b);
    outputs(2971) <= not b;
    outputs(2972) <= b;
    outputs(2973) <= b;
    outputs(2974) <= not b or a;
    outputs(2975) <= a and not b;
    outputs(2976) <= not a;
    outputs(2977) <= b;
    outputs(2978) <= not (a xor b);
    outputs(2979) <= a xor b;
    outputs(2980) <= not (a xor b);
    outputs(2981) <= b;
    outputs(2982) <= a xor b;
    outputs(2983) <= not b;
    outputs(2984) <= a;
    outputs(2985) <= b;
    outputs(2986) <= b and not a;
    outputs(2987) <= not a;
    outputs(2988) <= not a;
    outputs(2989) <= not b or a;
    outputs(2990) <= b;
    outputs(2991) <= not (a and b);
    outputs(2992) <= a xor b;
    outputs(2993) <= not b;
    outputs(2994) <= a;
    outputs(2995) <= a xor b;
    outputs(2996) <= a xor b;
    outputs(2997) <= not b or a;
    outputs(2998) <= b;
    outputs(2999) <= not (a xor b);
    outputs(3000) <= b;
    outputs(3001) <= a or b;
    outputs(3002) <= a and not b;
    outputs(3003) <= b;
    outputs(3004) <= a xor b;
    outputs(3005) <= a or b;
    outputs(3006) <= b;
    outputs(3007) <= a and b;
    outputs(3008) <= not (a and b);
    outputs(3009) <= not a;
    outputs(3010) <= a xor b;
    outputs(3011) <= a or b;
    outputs(3012) <= a xor b;
    outputs(3013) <= not (a xor b);
    outputs(3014) <= not (a and b);
    outputs(3015) <= not a or b;
    outputs(3016) <= not (a xor b);
    outputs(3017) <= not (a xor b);
    outputs(3018) <= not a;
    outputs(3019) <= not (a xor b);
    outputs(3020) <= not a or b;
    outputs(3021) <= a and not b;
    outputs(3022) <= not (a and b);
    outputs(3023) <= not (a xor b);
    outputs(3024) <= b and not a;
    outputs(3025) <= not b or a;
    outputs(3026) <= b and not a;
    outputs(3027) <= a and not b;
    outputs(3028) <= a xor b;
    outputs(3029) <= a and b;
    outputs(3030) <= not a;
    outputs(3031) <= not (a or b);
    outputs(3032) <= not b or a;
    outputs(3033) <= a xor b;
    outputs(3034) <= not a or b;
    outputs(3035) <= b and not a;
    outputs(3036) <= not b;
    outputs(3037) <= not (a or b);
    outputs(3038) <= b and not a;
    outputs(3039) <= b;
    outputs(3040) <= a and b;
    outputs(3041) <= not (a or b);
    outputs(3042) <= a;
    outputs(3043) <= a xor b;
    outputs(3044) <= a or b;
    outputs(3045) <= not a;
    outputs(3046) <= a or b;
    outputs(3047) <= a xor b;
    outputs(3048) <= not b;
    outputs(3049) <= a xor b;
    outputs(3050) <= a xor b;
    outputs(3051) <= not b;
    outputs(3052) <= a and b;
    outputs(3053) <= a xor b;
    outputs(3054) <= not a;
    outputs(3055) <= a and b;
    outputs(3056) <= a and not b;
    outputs(3057) <= a and b;
    outputs(3058) <= not b;
    outputs(3059) <= a xor b;
    outputs(3060) <= not (a and b);
    outputs(3061) <= a xor b;
    outputs(3062) <= not b;
    outputs(3063) <= a xor b;
    outputs(3064) <= not (a and b);
    outputs(3065) <= not b;
    outputs(3066) <= a;
    outputs(3067) <= b and not a;
    outputs(3068) <= a;
    outputs(3069) <= not b;
    outputs(3070) <= not a;
    outputs(3071) <= not a;
    outputs(3072) <= a xor b;
    outputs(3073) <= a and not b;
    outputs(3074) <= not (a and b);
    outputs(3075) <= a xor b;
    outputs(3076) <= b;
    outputs(3077) <= not a or b;
    outputs(3078) <= not (a xor b);
    outputs(3079) <= not a;
    outputs(3080) <= a xor b;
    outputs(3081) <= a and not b;
    outputs(3082) <= b;
    outputs(3083) <= not (a xor b);
    outputs(3084) <= not (a xor b);
    outputs(3085) <= b;
    outputs(3086) <= not (a xor b);
    outputs(3087) <= not a;
    outputs(3088) <= b;
    outputs(3089) <= b and not a;
    outputs(3090) <= a xor b;
    outputs(3091) <= a and b;
    outputs(3092) <= b;
    outputs(3093) <= a xor b;
    outputs(3094) <= b;
    outputs(3095) <= b;
    outputs(3096) <= not (a xor b);
    outputs(3097) <= not a or b;
    outputs(3098) <= not b;
    outputs(3099) <= not b;
    outputs(3100) <= a xor b;
    outputs(3101) <= not a or b;
    outputs(3102) <= a or b;
    outputs(3103) <= a;
    outputs(3104) <= not (a xor b);
    outputs(3105) <= a or b;
    outputs(3106) <= not b;
    outputs(3107) <= not (a and b);
    outputs(3108) <= a xor b;
    outputs(3109) <= a xor b;
    outputs(3110) <= not (a and b);
    outputs(3111) <= not (a xor b);
    outputs(3112) <= not b;
    outputs(3113) <= not a or b;
    outputs(3114) <= a xor b;
    outputs(3115) <= a xor b;
    outputs(3116) <= not (a xor b);
    outputs(3117) <= not a or b;
    outputs(3118) <= not a;
    outputs(3119) <= not a or b;
    outputs(3120) <= not (a xor b);
    outputs(3121) <= not (a xor b);
    outputs(3122) <= not (a xor b);
    outputs(3123) <= a and not b;
    outputs(3124) <= not (a and b);
    outputs(3125) <= a or b;
    outputs(3126) <= a;
    outputs(3127) <= not b;
    outputs(3128) <= a xor b;
    outputs(3129) <= a;
    outputs(3130) <= a and not b;
    outputs(3131) <= a or b;
    outputs(3132) <= not b or a;
    outputs(3133) <= a xor b;
    outputs(3134) <= not b;
    outputs(3135) <= not a;
    outputs(3136) <= b;
    outputs(3137) <= not b;
    outputs(3138) <= not a;
    outputs(3139) <= a;
    outputs(3140) <= b and not a;
    outputs(3141) <= a or b;
    outputs(3142) <= not a or b;
    outputs(3143) <= b and not a;
    outputs(3144) <= not (a xor b);
    outputs(3145) <= not (a xor b);
    outputs(3146) <= a;
    outputs(3147) <= a;
    outputs(3148) <= a;
    outputs(3149) <= not b;
    outputs(3150) <= not a;
    outputs(3151) <= b;
    outputs(3152) <= not a;
    outputs(3153) <= a xor b;
    outputs(3154) <= not (a xor b);
    outputs(3155) <= not a;
    outputs(3156) <= not b;
    outputs(3157) <= a or b;
    outputs(3158) <= b;
    outputs(3159) <= a and not b;
    outputs(3160) <= not (a or b);
    outputs(3161) <= not b;
    outputs(3162) <= not b or a;
    outputs(3163) <= a and b;
    outputs(3164) <= not (a xor b);
    outputs(3165) <= not b or a;
    outputs(3166) <= b and not a;
    outputs(3167) <= a xor b;
    outputs(3168) <= a xor b;
    outputs(3169) <= not (a or b);
    outputs(3170) <= a xor b;
    outputs(3171) <= not (a or b);
    outputs(3172) <= not (a xor b);
    outputs(3173) <= a and not b;
    outputs(3174) <= not (a xor b);
    outputs(3175) <= b;
    outputs(3176) <= b and not a;
    outputs(3177) <= a and b;
    outputs(3178) <= a xor b;
    outputs(3179) <= not b;
    outputs(3180) <= not (a xor b);
    outputs(3181) <= a xor b;
    outputs(3182) <= a xor b;
    outputs(3183) <= b;
    outputs(3184) <= not (a xor b);
    outputs(3185) <= not a or b;
    outputs(3186) <= a;
    outputs(3187) <= not a;
    outputs(3188) <= a xor b;
    outputs(3189) <= b and not a;
    outputs(3190) <= not b;
    outputs(3191) <= not (a or b);
    outputs(3192) <= not a;
    outputs(3193) <= not (a xor b);
    outputs(3194) <= a and not b;
    outputs(3195) <= not b;
    outputs(3196) <= a xor b;
    outputs(3197) <= a;
    outputs(3198) <= not (a xor b);
    outputs(3199) <= a xor b;
    outputs(3200) <= a;
    outputs(3201) <= not (a xor b);
    outputs(3202) <= not (a or b);
    outputs(3203) <= b;
    outputs(3204) <= a xor b;
    outputs(3205) <= not (a xor b);
    outputs(3206) <= not a;
    outputs(3207) <= not b;
    outputs(3208) <= not (a or b);
    outputs(3209) <= not b;
    outputs(3210) <= not (a xor b);
    outputs(3211) <= not b or a;
    outputs(3212) <= b and not a;
    outputs(3213) <= a and not b;
    outputs(3214) <= not (a xor b);
    outputs(3215) <= a or b;
    outputs(3216) <= not b;
    outputs(3217) <= not (a xor b);
    outputs(3218) <= not (a xor b);
    outputs(3219) <= a;
    outputs(3220) <= a and not b;
    outputs(3221) <= a;
    outputs(3222) <= a xor b;
    outputs(3223) <= b;
    outputs(3224) <= a;
    outputs(3225) <= not (a xor b);
    outputs(3226) <= a xor b;
    outputs(3227) <= a xor b;
    outputs(3228) <= not a;
    outputs(3229) <= not (a xor b);
    outputs(3230) <= b;
    outputs(3231) <= not (a or b);
    outputs(3232) <= not (a xor b);
    outputs(3233) <= a or b;
    outputs(3234) <= b;
    outputs(3235) <= b and not a;
    outputs(3236) <= not (a xor b);
    outputs(3237) <= not b;
    outputs(3238) <= a and not b;
    outputs(3239) <= b;
    outputs(3240) <= not (a xor b);
    outputs(3241) <= a xor b;
    outputs(3242) <= a xor b;
    outputs(3243) <= not b;
    outputs(3244) <= a xor b;
    outputs(3245) <= not b or a;
    outputs(3246) <= not (a and b);
    outputs(3247) <= b;
    outputs(3248) <= not (a xor b);
    outputs(3249) <= b;
    outputs(3250) <= not (a xor b);
    outputs(3251) <= not (a xor b);
    outputs(3252) <= b and not a;
    outputs(3253) <= not b or a;
    outputs(3254) <= a xor b;
    outputs(3255) <= a;
    outputs(3256) <= b;
    outputs(3257) <= a xor b;
    outputs(3258) <= a xor b;
    outputs(3259) <= b;
    outputs(3260) <= a and not b;
    outputs(3261) <= a xor b;
    outputs(3262) <= a xor b;
    outputs(3263) <= a xor b;
    outputs(3264) <= a and not b;
    outputs(3265) <= b and not a;
    outputs(3266) <= a and b;
    outputs(3267) <= a xor b;
    outputs(3268) <= not a or b;
    outputs(3269) <= not a;
    outputs(3270) <= b;
    outputs(3271) <= not (a or b);
    outputs(3272) <= a;
    outputs(3273) <= not b;
    outputs(3274) <= not (a or b);
    outputs(3275) <= not b;
    outputs(3276) <= a;
    outputs(3277) <= a;
    outputs(3278) <= a xor b;
    outputs(3279) <= a and b;
    outputs(3280) <= not (a and b);
    outputs(3281) <= a;
    outputs(3282) <= not (a xor b);
    outputs(3283) <= not a or b;
    outputs(3284) <= not (a xor b);
    outputs(3285) <= not (a or b);
    outputs(3286) <= b;
    outputs(3287) <= not (a xor b);
    outputs(3288) <= not (a or b);
    outputs(3289) <= not b;
    outputs(3290) <= b;
    outputs(3291) <= a and b;
    outputs(3292) <= b and not a;
    outputs(3293) <= not a;
    outputs(3294) <= a;
    outputs(3295) <= b and not a;
    outputs(3296) <= not (a xor b);
    outputs(3297) <= a xor b;
    outputs(3298) <= not a or b;
    outputs(3299) <= not a;
    outputs(3300) <= a;
    outputs(3301) <= a xor b;
    outputs(3302) <= not a;
    outputs(3303) <= not b;
    outputs(3304) <= not a or b;
    outputs(3305) <= a xor b;
    outputs(3306) <= a;
    outputs(3307) <= not (a xor b);
    outputs(3308) <= a xor b;
    outputs(3309) <= not (a xor b);
    outputs(3310) <= a;
    outputs(3311) <= not a or b;
    outputs(3312) <= not a;
    outputs(3313) <= b;
    outputs(3314) <= a xor b;
    outputs(3315) <= not a or b;
    outputs(3316) <= a or b;
    outputs(3317) <= not a;
    outputs(3318) <= not b;
    outputs(3319) <= not (a xor b);
    outputs(3320) <= not b or a;
    outputs(3321) <= not a;
    outputs(3322) <= not (a and b);
    outputs(3323) <= b;
    outputs(3324) <= not a;
    outputs(3325) <= a xor b;
    outputs(3326) <= a and not b;
    outputs(3327) <= not (a xor b);
    outputs(3328) <= a xor b;
    outputs(3329) <= a;
    outputs(3330) <= a xor b;
    outputs(3331) <= a xor b;
    outputs(3332) <= not a or b;
    outputs(3333) <= not b or a;
    outputs(3334) <= not b;
    outputs(3335) <= not a or b;
    outputs(3336) <= a and not b;
    outputs(3337) <= not (a or b);
    outputs(3338) <= not (a xor b);
    outputs(3339) <= not a;
    outputs(3340) <= not b or a;
    outputs(3341) <= a xor b;
    outputs(3342) <= not (a and b);
    outputs(3343) <= a;
    outputs(3344) <= not (a or b);
    outputs(3345) <= not b;
    outputs(3346) <= not (a xor b);
    outputs(3347) <= a and not b;
    outputs(3348) <= not a;
    outputs(3349) <= not (a xor b);
    outputs(3350) <= not a;
    outputs(3351) <= not (a xor b);
    outputs(3352) <= b;
    outputs(3353) <= not b;
    outputs(3354) <= not (a and b);
    outputs(3355) <= not a or b;
    outputs(3356) <= b;
    outputs(3357) <= not (a xor b);
    outputs(3358) <= a xor b;
    outputs(3359) <= a;
    outputs(3360) <= a and b;
    outputs(3361) <= a;
    outputs(3362) <= a;
    outputs(3363) <= a xor b;
    outputs(3364) <= not b;
    outputs(3365) <= not b;
    outputs(3366) <= not b or a;
    outputs(3367) <= not (a or b);
    outputs(3368) <= not b;
    outputs(3369) <= not (a xor b);
    outputs(3370) <= a;
    outputs(3371) <= a and b;
    outputs(3372) <= not (a xor b);
    outputs(3373) <= not b;
    outputs(3374) <= not a;
    outputs(3375) <= a;
    outputs(3376) <= a xor b;
    outputs(3377) <= not b or a;
    outputs(3378) <= not (a or b);
    outputs(3379) <= not b or a;
    outputs(3380) <= a;
    outputs(3381) <= a xor b;
    outputs(3382) <= not (a xor b);
    outputs(3383) <= a and not b;
    outputs(3384) <= a and not b;
    outputs(3385) <= not (a or b);
    outputs(3386) <= a;
    outputs(3387) <= b;
    outputs(3388) <= not b;
    outputs(3389) <= a xor b;
    outputs(3390) <= b;
    outputs(3391) <= a xor b;
    outputs(3392) <= a;
    outputs(3393) <= a;
    outputs(3394) <= not b;
    outputs(3395) <= not b;
    outputs(3396) <= a;
    outputs(3397) <= a or b;
    outputs(3398) <= not b;
    outputs(3399) <= a and not b;
    outputs(3400) <= not b;
    outputs(3401) <= not b;
    outputs(3402) <= a xor b;
    outputs(3403) <= b;
    outputs(3404) <= a;
    outputs(3405) <= not a;
    outputs(3406) <= a and b;
    outputs(3407) <= a or b;
    outputs(3408) <= b and not a;
    outputs(3409) <= a;
    outputs(3410) <= not a or b;
    outputs(3411) <= a xor b;
    outputs(3412) <= not b;
    outputs(3413) <= a;
    outputs(3414) <= not a or b;
    outputs(3415) <= not a;
    outputs(3416) <= b and not a;
    outputs(3417) <= not (a or b);
    outputs(3418) <= not a;
    outputs(3419) <= a;
    outputs(3420) <= not (a xor b);
    outputs(3421) <= not b or a;
    outputs(3422) <= a xor b;
    outputs(3423) <= not a;
    outputs(3424) <= a;
    outputs(3425) <= not (a or b);
    outputs(3426) <= a and b;
    outputs(3427) <= b and not a;
    outputs(3428) <= not (a xor b);
    outputs(3429) <= not a;
    outputs(3430) <= not b;
    outputs(3431) <= a;
    outputs(3432) <= a;
    outputs(3433) <= a xor b;
    outputs(3434) <= b;
    outputs(3435) <= not b or a;
    outputs(3436) <= not b;
    outputs(3437) <= a or b;
    outputs(3438) <= b;
    outputs(3439) <= b;
    outputs(3440) <= b;
    outputs(3441) <= not b;
    outputs(3442) <= b;
    outputs(3443) <= not b;
    outputs(3444) <= not a;
    outputs(3445) <= not (a or b);
    outputs(3446) <= not (a or b);
    outputs(3447) <= not (a and b);
    outputs(3448) <= a and not b;
    outputs(3449) <= a and b;
    outputs(3450) <= b;
    outputs(3451) <= a;
    outputs(3452) <= a xor b;
    outputs(3453) <= not (a or b);
    outputs(3454) <= b and not a;
    outputs(3455) <= a;
    outputs(3456) <= not a or b;
    outputs(3457) <= a;
    outputs(3458) <= not b;
    outputs(3459) <= b;
    outputs(3460) <= a and not b;
    outputs(3461) <= not (a and b);
    outputs(3462) <= not b;
    outputs(3463) <= not (a or b);
    outputs(3464) <= a and b;
    outputs(3465) <= not (a and b);
    outputs(3466) <= b;
    outputs(3467) <= not (a or b);
    outputs(3468) <= a and not b;
    outputs(3469) <= a or b;
    outputs(3470) <= not (a and b);
    outputs(3471) <= not b;
    outputs(3472) <= not b or a;
    outputs(3473) <= a;
    outputs(3474) <= b and not a;
    outputs(3475) <= a and not b;
    outputs(3476) <= not b;
    outputs(3477) <= b and not a;
    outputs(3478) <= not b;
    outputs(3479) <= a xor b;
    outputs(3480) <= not b;
    outputs(3481) <= not b or a;
    outputs(3482) <= a;
    outputs(3483) <= a xor b;
    outputs(3484) <= a xor b;
    outputs(3485) <= not a;
    outputs(3486) <= not (a xor b);
    outputs(3487) <= not (a and b);
    outputs(3488) <= a;
    outputs(3489) <= not (a and b);
    outputs(3490) <= not (a or b);
    outputs(3491) <= not (a xor b);
    outputs(3492) <= not b or a;
    outputs(3493) <= a or b;
    outputs(3494) <= not a;
    outputs(3495) <= not b;
    outputs(3496) <= b;
    outputs(3497) <= not b;
    outputs(3498) <= not b or a;
    outputs(3499) <= a xor b;
    outputs(3500) <= b;
    outputs(3501) <= a or b;
    outputs(3502) <= not b;
    outputs(3503) <= not (a and b);
    outputs(3504) <= b and not a;
    outputs(3505) <= b;
    outputs(3506) <= not b;
    outputs(3507) <= not a;
    outputs(3508) <= not (a xor b);
    outputs(3509) <= a xor b;
    outputs(3510) <= b;
    outputs(3511) <= a xor b;
    outputs(3512) <= not b;
    outputs(3513) <= b;
    outputs(3514) <= a;
    outputs(3515) <= not b;
    outputs(3516) <= a and b;
    outputs(3517) <= not (a and b);
    outputs(3518) <= a xor b;
    outputs(3519) <= not a or b;
    outputs(3520) <= not (a and b);
    outputs(3521) <= not a or b;
    outputs(3522) <= not a or b;
    outputs(3523) <= a or b;
    outputs(3524) <= not b or a;
    outputs(3525) <= not b or a;
    outputs(3526) <= not a;
    outputs(3527) <= not b;
    outputs(3528) <= not a or b;
    outputs(3529) <= a xor b;
    outputs(3530) <= not (a xor b);
    outputs(3531) <= a xor b;
    outputs(3532) <= not b;
    outputs(3533) <= b;
    outputs(3534) <= b;
    outputs(3535) <= a xor b;
    outputs(3536) <= a xor b;
    outputs(3537) <= a;
    outputs(3538) <= b and not a;
    outputs(3539) <= a xor b;
    outputs(3540) <= not a;
    outputs(3541) <= a;
    outputs(3542) <= not b;
    outputs(3543) <= a xor b;
    outputs(3544) <= not a or b;
    outputs(3545) <= not b;
    outputs(3546) <= a;
    outputs(3547) <= not a or b;
    outputs(3548) <= not (a xor b);
    outputs(3549) <= not (a xor b);
    outputs(3550) <= a xor b;
    outputs(3551) <= not b;
    outputs(3552) <= not b or a;
    outputs(3553) <= not a;
    outputs(3554) <= b;
    outputs(3555) <= b and not a;
    outputs(3556) <= a and not b;
    outputs(3557) <= a or b;
    outputs(3558) <= a xor b;
    outputs(3559) <= b and not a;
    outputs(3560) <= a xor b;
    outputs(3561) <= not b;
    outputs(3562) <= not (a xor b);
    outputs(3563) <= not b;
    outputs(3564) <= a xor b;
    outputs(3565) <= b;
    outputs(3566) <= not (a xor b);
    outputs(3567) <= not (a xor b);
    outputs(3568) <= not b;
    outputs(3569) <= a;
    outputs(3570) <= a;
    outputs(3571) <= b;
    outputs(3572) <= a;
    outputs(3573) <= a;
    outputs(3574) <= not b;
    outputs(3575) <= not a;
    outputs(3576) <= not b;
    outputs(3577) <= not (a xor b);
    outputs(3578) <= not (a xor b);
    outputs(3579) <= a and not b;
    outputs(3580) <= not (a and b);
    outputs(3581) <= a or b;
    outputs(3582) <= not (a xor b);
    outputs(3583) <= not b or a;
    outputs(3584) <= a and b;
    outputs(3585) <= b;
    outputs(3586) <= not b;
    outputs(3587) <= a and not b;
    outputs(3588) <= a or b;
    outputs(3589) <= not b or a;
    outputs(3590) <= not a;
    outputs(3591) <= not a;
    outputs(3592) <= a xor b;
    outputs(3593) <= not a;
    outputs(3594) <= a and not b;
    outputs(3595) <= not a;
    outputs(3596) <= not a;
    outputs(3597) <= a;
    outputs(3598) <= a xor b;
    outputs(3599) <= not a or b;
    outputs(3600) <= not (a xor b);
    outputs(3601) <= not b or a;
    outputs(3602) <= b;
    outputs(3603) <= a and b;
    outputs(3604) <= a xor b;
    outputs(3605) <= a xor b;
    outputs(3606) <= not (a xor b);
    outputs(3607) <= a;
    outputs(3608) <= a xor b;
    outputs(3609) <= not b;
    outputs(3610) <= not a;
    outputs(3611) <= a;
    outputs(3612) <= a and b;
    outputs(3613) <= a xor b;
    outputs(3614) <= a xor b;
    outputs(3615) <= not (a xor b);
    outputs(3616) <= not (a and b);
    outputs(3617) <= a;
    outputs(3618) <= a xor b;
    outputs(3619) <= not b or a;
    outputs(3620) <= not (a xor b);
    outputs(3621) <= not a or b;
    outputs(3622) <= not a;
    outputs(3623) <= a xor b;
    outputs(3624) <= b;
    outputs(3625) <= not a;
    outputs(3626) <= not (a xor b);
    outputs(3627) <= not a or b;
    outputs(3628) <= a;
    outputs(3629) <= b;
    outputs(3630) <= not a;
    outputs(3631) <= not (a xor b);
    outputs(3632) <= not (a xor b);
    outputs(3633) <= a xor b;
    outputs(3634) <= a xor b;
    outputs(3635) <= b;
    outputs(3636) <= not a;
    outputs(3637) <= a or b;
    outputs(3638) <= b and not a;
    outputs(3639) <= not (a or b);
    outputs(3640) <= not a;
    outputs(3641) <= not b;
    outputs(3642) <= a xor b;
    outputs(3643) <= a;
    outputs(3644) <= not (a and b);
    outputs(3645) <= b and not a;
    outputs(3646) <= b and not a;
    outputs(3647) <= not b or a;
    outputs(3648) <= a and b;
    outputs(3649) <= not b;
    outputs(3650) <= a and b;
    outputs(3651) <= a xor b;
    outputs(3652) <= not a or b;
    outputs(3653) <= b;
    outputs(3654) <= a or b;
    outputs(3655) <= a xor b;
    outputs(3656) <= not a;
    outputs(3657) <= not a;
    outputs(3658) <= not b;
    outputs(3659) <= a;
    outputs(3660) <= not b;
    outputs(3661) <= not a;
    outputs(3662) <= b and not a;
    outputs(3663) <= a;
    outputs(3664) <= b;
    outputs(3665) <= a;
    outputs(3666) <= a xor b;
    outputs(3667) <= not (a xor b);
    outputs(3668) <= not a;
    outputs(3669) <= a xor b;
    outputs(3670) <= not (a xor b);
    outputs(3671) <= b;
    outputs(3672) <= a;
    outputs(3673) <= b;
    outputs(3674) <= b and not a;
    outputs(3675) <= not a;
    outputs(3676) <= a and b;
    outputs(3677) <= a or b;
    outputs(3678) <= a;
    outputs(3679) <= not a;
    outputs(3680) <= not a or b;
    outputs(3681) <= a and b;
    outputs(3682) <= a and not b;
    outputs(3683) <= not (a xor b);
    outputs(3684) <= not (a xor b);
    outputs(3685) <= a xor b;
    outputs(3686) <= b;
    outputs(3687) <= not (a xor b);
    outputs(3688) <= not a;
    outputs(3689) <= not b;
    outputs(3690) <= not a or b;
    outputs(3691) <= not b;
    outputs(3692) <= a xor b;
    outputs(3693) <= a and not b;
    outputs(3694) <= a or b;
    outputs(3695) <= not (a xor b);
    outputs(3696) <= not (a xor b);
    outputs(3697) <= a and b;
    outputs(3698) <= not (a or b);
    outputs(3699) <= b;
    outputs(3700) <= not (a xor b);
    outputs(3701) <= not (a xor b);
    outputs(3702) <= not (a and b);
    outputs(3703) <= b and not a;
    outputs(3704) <= not b;
    outputs(3705) <= b;
    outputs(3706) <= not (a and b);
    outputs(3707) <= not (a xor b);
    outputs(3708) <= a xor b;
    outputs(3709) <= b and not a;
    outputs(3710) <= not (a or b);
    outputs(3711) <= not a;
    outputs(3712) <= not (a or b);
    outputs(3713) <= b and not a;
    outputs(3714) <= b and not a;
    outputs(3715) <= a and b;
    outputs(3716) <= not (a or b);
    outputs(3717) <= a;
    outputs(3718) <= a and not b;
    outputs(3719) <= not (a or b);
    outputs(3720) <= not a;
    outputs(3721) <= b and not a;
    outputs(3722) <= not b;
    outputs(3723) <= b;
    outputs(3724) <= a xor b;
    outputs(3725) <= a and b;
    outputs(3726) <= not (a and b);
    outputs(3727) <= b;
    outputs(3728) <= not a;
    outputs(3729) <= a xor b;
    outputs(3730) <= a and b;
    outputs(3731) <= b and not a;
    outputs(3732) <= not a;
    outputs(3733) <= not b;
    outputs(3734) <= a;
    outputs(3735) <= b;
    outputs(3736) <= b;
    outputs(3737) <= a xor b;
    outputs(3738) <= not (a xor b);
    outputs(3739) <= a and b;
    outputs(3740) <= a or b;
    outputs(3741) <= not b or a;
    outputs(3742) <= a;
    outputs(3743) <= a and not b;
    outputs(3744) <= a xor b;
    outputs(3745) <= a;
    outputs(3746) <= not b;
    outputs(3747) <= not a;
    outputs(3748) <= a;
    outputs(3749) <= not (a xor b);
    outputs(3750) <= not (a or b);
    outputs(3751) <= a and b;
    outputs(3752) <= a;
    outputs(3753) <= a and b;
    outputs(3754) <= not (a xor b);
    outputs(3755) <= not (a or b);
    outputs(3756) <= not b;
    outputs(3757) <= not b or a;
    outputs(3758) <= not b;
    outputs(3759) <= a xor b;
    outputs(3760) <= not (a xor b);
    outputs(3761) <= b and not a;
    outputs(3762) <= a xor b;
    outputs(3763) <= b and not a;
    outputs(3764) <= not (a xor b);
    outputs(3765) <= a and b;
    outputs(3766) <= a;
    outputs(3767) <= not b;
    outputs(3768) <= b;
    outputs(3769) <= a and not b;
    outputs(3770) <= not b or a;
    outputs(3771) <= not (a and b);
    outputs(3772) <= not (a and b);
    outputs(3773) <= a and b;
    outputs(3774) <= not (a xor b);
    outputs(3775) <= not a or b;
    outputs(3776) <= not (a xor b);
    outputs(3777) <= b and not a;
    outputs(3778) <= a;
    outputs(3779) <= not b;
    outputs(3780) <= not (a xor b);
    outputs(3781) <= a;
    outputs(3782) <= a and b;
    outputs(3783) <= not b or a;
    outputs(3784) <= b;
    outputs(3785) <= not b;
    outputs(3786) <= not a;
    outputs(3787) <= a;
    outputs(3788) <= not b;
    outputs(3789) <= not b or a;
    outputs(3790) <= not (a or b);
    outputs(3791) <= a;
    outputs(3792) <= not a;
    outputs(3793) <= not b or a;
    outputs(3794) <= b;
    outputs(3795) <= a;
    outputs(3796) <= a xor b;
    outputs(3797) <= not b;
    outputs(3798) <= not (a xor b);
    outputs(3799) <= b and not a;
    outputs(3800) <= not (a xor b);
    outputs(3801) <= not (a xor b);
    outputs(3802) <= not (a xor b);
    outputs(3803) <= not (a or b);
    outputs(3804) <= b and not a;
    outputs(3805) <= not b;
    outputs(3806) <= a xor b;
    outputs(3807) <= a;
    outputs(3808) <= a xor b;
    outputs(3809) <= not a or b;
    outputs(3810) <= not (a xor b);
    outputs(3811) <= a;
    outputs(3812) <= a xor b;
    outputs(3813) <= a xor b;
    outputs(3814) <= a or b;
    outputs(3815) <= a and b;
    outputs(3816) <= a and b;
    outputs(3817) <= not (a xor b);
    outputs(3818) <= a xor b;
    outputs(3819) <= a and not b;
    outputs(3820) <= a;
    outputs(3821) <= a or b;
    outputs(3822) <= not b or a;
    outputs(3823) <= not (a xor b);
    outputs(3824) <= not a;
    outputs(3825) <= a xor b;
    outputs(3826) <= not (a xor b);
    outputs(3827) <= not a;
    outputs(3828) <= a xor b;
    outputs(3829) <= not (a and b);
    outputs(3830) <= a and b;
    outputs(3831) <= a;
    outputs(3832) <= not b;
    outputs(3833) <= b;
    outputs(3834) <= not (a xor b);
    outputs(3835) <= a xor b;
    outputs(3836) <= not (a xor b);
    outputs(3837) <= not (a xor b);
    outputs(3838) <= a xor b;
    outputs(3839) <= not b or a;
    outputs(3840) <= b and not a;
    outputs(3841) <= a or b;
    outputs(3842) <= not a;
    outputs(3843) <= not b;
    outputs(3844) <= not (a and b);
    outputs(3845) <= b;
    outputs(3846) <= a xor b;
    outputs(3847) <= not b;
    outputs(3848) <= not b;
    outputs(3849) <= a xor b;
    outputs(3850) <= not (a xor b);
    outputs(3851) <= not b;
    outputs(3852) <= a and b;
    outputs(3853) <= not (a and b);
    outputs(3854) <= a;
    outputs(3855) <= a xor b;
    outputs(3856) <= a;
    outputs(3857) <= b;
    outputs(3858) <= b;
    outputs(3859) <= not (a xor b);
    outputs(3860) <= a or b;
    outputs(3861) <= a xor b;
    outputs(3862) <= not b;
    outputs(3863) <= not b;
    outputs(3864) <= not a;
    outputs(3865) <= a xor b;
    outputs(3866) <= not b;
    outputs(3867) <= not (a or b);
    outputs(3868) <= a and not b;
    outputs(3869) <= a;
    outputs(3870) <= a xor b;
    outputs(3871) <= not b or a;
    outputs(3872) <= a;
    outputs(3873) <= not (a or b);
    outputs(3874) <= not (a or b);
    outputs(3875) <= not (a xor b);
    outputs(3876) <= a xor b;
    outputs(3877) <= not b or a;
    outputs(3878) <= a;
    outputs(3879) <= a and not b;
    outputs(3880) <= not (a or b);
    outputs(3881) <= not a;
    outputs(3882) <= a xor b;
    outputs(3883) <= a or b;
    outputs(3884) <= a xor b;
    outputs(3885) <= not (a xor b);
    outputs(3886) <= b and not a;
    outputs(3887) <= b;
    outputs(3888) <= a xor b;
    outputs(3889) <= not a or b;
    outputs(3890) <= not (a xor b);
    outputs(3891) <= a xor b;
    outputs(3892) <= not b;
    outputs(3893) <= b and not a;
    outputs(3894) <= not a;
    outputs(3895) <= a xor b;
    outputs(3896) <= not a;
    outputs(3897) <= a;
    outputs(3898) <= b and not a;
    outputs(3899) <= a;
    outputs(3900) <= not b;
    outputs(3901) <= b and not a;
    outputs(3902) <= a;
    outputs(3903) <= not (a and b);
    outputs(3904) <= a xor b;
    outputs(3905) <= a xor b;
    outputs(3906) <= b and not a;
    outputs(3907) <= not b;
    outputs(3908) <= b;
    outputs(3909) <= not (a or b);
    outputs(3910) <= not b or a;
    outputs(3911) <= not b;
    outputs(3912) <= a;
    outputs(3913) <= not b;
    outputs(3914) <= not (a xor b);
    outputs(3915) <= a;
    outputs(3916) <= not (a and b);
    outputs(3917) <= not (a xor b);
    outputs(3918) <= a and not b;
    outputs(3919) <= a;
    outputs(3920) <= not a;
    outputs(3921) <= a and b;
    outputs(3922) <= not a or b;
    outputs(3923) <= not b or a;
    outputs(3924) <= a or b;
    outputs(3925) <= a or b;
    outputs(3926) <= not (a xor b);
    outputs(3927) <= b;
    outputs(3928) <= not b;
    outputs(3929) <= b and not a;
    outputs(3930) <= not a;
    outputs(3931) <= b;
    outputs(3932) <= not a;
    outputs(3933) <= not b or a;
    outputs(3934) <= a;
    outputs(3935) <= a xor b;
    outputs(3936) <= not b or a;
    outputs(3937) <= a;
    outputs(3938) <= not (a xor b);
    outputs(3939) <= a xor b;
    outputs(3940) <= not (a and b);
    outputs(3941) <= not a;
    outputs(3942) <= a xor b;
    outputs(3943) <= a;
    outputs(3944) <= a xor b;
    outputs(3945) <= a;
    outputs(3946) <= not a;
    outputs(3947) <= not b;
    outputs(3948) <= not (a or b);
    outputs(3949) <= a and not b;
    outputs(3950) <= not (a or b);
    outputs(3951) <= a and not b;
    outputs(3952) <= not (a xor b);
    outputs(3953) <= b;
    outputs(3954) <= not (a xor b);
    outputs(3955) <= not (a and b);
    outputs(3956) <= a xor b;
    outputs(3957) <= not (a or b);
    outputs(3958) <= not b;
    outputs(3959) <= not (a or b);
    outputs(3960) <= not b;
    outputs(3961) <= not (a xor b);
    outputs(3962) <= b;
    outputs(3963) <= a or b;
    outputs(3964) <= a and not b;
    outputs(3965) <= not (a or b);
    outputs(3966) <= a and b;
    outputs(3967) <= not (a xor b);
    outputs(3968) <= a and b;
    outputs(3969) <= b;
    outputs(3970) <= b and not a;
    outputs(3971) <= not (a or b);
    outputs(3972) <= b and not a;
    outputs(3973) <= not b;
    outputs(3974) <= a;
    outputs(3975) <= a and not b;
    outputs(3976) <= not a;
    outputs(3977) <= a xor b;
    outputs(3978) <= not (a xor b);
    outputs(3979) <= a;
    outputs(3980) <= a xor b;
    outputs(3981) <= a;
    outputs(3982) <= not b;
    outputs(3983) <= not (a xor b);
    outputs(3984) <= not (a or b);
    outputs(3985) <= a xor b;
    outputs(3986) <= a;
    outputs(3987) <= a;
    outputs(3988) <= not (a and b);
    outputs(3989) <= b and not a;
    outputs(3990) <= a and not b;
    outputs(3991) <= not b;
    outputs(3992) <= a;
    outputs(3993) <= a and b;
    outputs(3994) <= a;
    outputs(3995) <= b;
    outputs(3996) <= a xor b;
    outputs(3997) <= a;
    outputs(3998) <= not (a or b);
    outputs(3999) <= not (a or b);
    outputs(4000) <= not (a xor b);
    outputs(4001) <= not a;
    outputs(4002) <= not (a xor b);
    outputs(4003) <= not a;
    outputs(4004) <= a xor b;
    outputs(4005) <= a xor b;
    outputs(4006) <= not (a or b);
    outputs(4007) <= b;
    outputs(4008) <= not (a and b);
    outputs(4009) <= a xor b;
    outputs(4010) <= a xor b;
    outputs(4011) <= not (a or b);
    outputs(4012) <= not b;
    outputs(4013) <= b;
    outputs(4014) <= not b;
    outputs(4015) <= not a or b;
    outputs(4016) <= a and b;
    outputs(4017) <= not (a xor b);
    outputs(4018) <= a xor b;
    outputs(4019) <= b and not a;
    outputs(4020) <= a xor b;
    outputs(4021) <= a xor b;
    outputs(4022) <= not (a xor b);
    outputs(4023) <= not (a xor b);
    outputs(4024) <= not a or b;
    outputs(4025) <= not a;
    outputs(4026) <= not (a and b);
    outputs(4027) <= a;
    outputs(4028) <= b;
    outputs(4029) <= not (a xor b);
    outputs(4030) <= a and not b;
    outputs(4031) <= not (a xor b);
    outputs(4032) <= not a;
    outputs(4033) <= a;
    outputs(4034) <= a;
    outputs(4035) <= not (a or b);
    outputs(4036) <= a xor b;
    outputs(4037) <= b;
    outputs(4038) <= not b or a;
    outputs(4039) <= not (a xor b);
    outputs(4040) <= a and not b;
    outputs(4041) <= not b;
    outputs(4042) <= not b;
    outputs(4043) <= not b;
    outputs(4044) <= a;
    outputs(4045) <= not (a xor b);
    outputs(4046) <= a and b;
    outputs(4047) <= a xor b;
    outputs(4048) <= a xor b;
    outputs(4049) <= not (a xor b);
    outputs(4050) <= a and b;
    outputs(4051) <= not b;
    outputs(4052) <= b;
    outputs(4053) <= a and b;
    outputs(4054) <= a xor b;
    outputs(4055) <= not a;
    outputs(4056) <= not (a xor b);
    outputs(4057) <= not b or a;
    outputs(4058) <= not (a and b);
    outputs(4059) <= a and not b;
    outputs(4060) <= b;
    outputs(4061) <= not (a or b);
    outputs(4062) <= not a;
    outputs(4063) <= a;
    outputs(4064) <= not (a xor b);
    outputs(4065) <= b;
    outputs(4066) <= not b;
    outputs(4067) <= not (a xor b);
    outputs(4068) <= a;
    outputs(4069) <= b;
    outputs(4070) <= not a;
    outputs(4071) <= a and b;
    outputs(4072) <= a xor b;
    outputs(4073) <= not b or a;
    outputs(4074) <= not b;
    outputs(4075) <= a and b;
    outputs(4076) <= b;
    outputs(4077) <= b;
    outputs(4078) <= a or b;
    outputs(4079) <= a;
    outputs(4080) <= b;
    outputs(4081) <= not (a or b);
    outputs(4082) <= not (a or b);
    outputs(4083) <= b;
    outputs(4084) <= a;
    outputs(4085) <= not (a or b);
    outputs(4086) <= not b;
    outputs(4087) <= not b;
    outputs(4088) <= a xor b;
    outputs(4089) <= not b;
    outputs(4090) <= a;
    outputs(4091) <= not b or a;
    outputs(4092) <= not (a xor b);
    outputs(4093) <= not a;
    outputs(4094) <= a and not b;
    outputs(4095) <= not a;
    outputs(4096) <= a;
    outputs(4097) <= not (a and b);
    outputs(4098) <= a xor b;
    outputs(4099) <= a xor b;
    outputs(4100) <= a;
    outputs(4101) <= not a;
    outputs(4102) <= not a or b;
    outputs(4103) <= not a;
    outputs(4104) <= not (a xor b);
    outputs(4105) <= not (a or b);
    outputs(4106) <= not (a xor b);
    outputs(4107) <= not a;
    outputs(4108) <= a and b;
    outputs(4109) <= b;
    outputs(4110) <= not (a xor b);
    outputs(4111) <= a;
    outputs(4112) <= b;
    outputs(4113) <= not a or b;
    outputs(4114) <= not a or b;
    outputs(4115) <= not (a xor b);
    outputs(4116) <= a and not b;
    outputs(4117) <= not (a or b);
    outputs(4118) <= not (a and b);
    outputs(4119) <= a;
    outputs(4120) <= not a;
    outputs(4121) <= a and b;
    outputs(4122) <= b and not a;
    outputs(4123) <= not b;
    outputs(4124) <= a xor b;
    outputs(4125) <= not b;
    outputs(4126) <= not (a or b);
    outputs(4127) <= not (a xor b);
    outputs(4128) <= a and not b;
    outputs(4129) <= not a;
    outputs(4130) <= a xor b;
    outputs(4131) <= b and not a;
    outputs(4132) <= b;
    outputs(4133) <= a xor b;
    outputs(4134) <= a xor b;
    outputs(4135) <= a and not b;
    outputs(4136) <= not b;
    outputs(4137) <= b and not a;
    outputs(4138) <= a xor b;
    outputs(4139) <= a xor b;
    outputs(4140) <= a xor b;
    outputs(4141) <= not (a xor b);
    outputs(4142) <= not b or a;
    outputs(4143) <= not b;
    outputs(4144) <= a and not b;
    outputs(4145) <= not (a xor b);
    outputs(4146) <= a and not b;
    outputs(4147) <= a;
    outputs(4148) <= not (a xor b);
    outputs(4149) <= not b;
    outputs(4150) <= not b;
    outputs(4151) <= not a;
    outputs(4152) <= not b;
    outputs(4153) <= not a;
    outputs(4154) <= not a;
    outputs(4155) <= not b;
    outputs(4156) <= not (a xor b);
    outputs(4157) <= a and not b;
    outputs(4158) <= not b;
    outputs(4159) <= a or b;
    outputs(4160) <= not (a xor b);
    outputs(4161) <= not b;
    outputs(4162) <= a or b;
    outputs(4163) <= a xor b;
    outputs(4164) <= a xor b;
    outputs(4165) <= b and not a;
    outputs(4166) <= not (a xor b);
    outputs(4167) <= a;
    outputs(4168) <= a;
    outputs(4169) <= not b;
    outputs(4170) <= not b;
    outputs(4171) <= not (a xor b);
    outputs(4172) <= not b;
    outputs(4173) <= a xor b;
    outputs(4174) <= not (a xor b);
    outputs(4175) <= not a or b;
    outputs(4176) <= b and not a;
    outputs(4177) <= b;
    outputs(4178) <= a xor b;
    outputs(4179) <= a and b;
    outputs(4180) <= not a;
    outputs(4181) <= a and not b;
    outputs(4182) <= not (a xor b);
    outputs(4183) <= a xor b;
    outputs(4184) <= not b or a;
    outputs(4185) <= not (a xor b);
    outputs(4186) <= not a;
    outputs(4187) <= not a;
    outputs(4188) <= not a;
    outputs(4189) <= not (a and b);
    outputs(4190) <= not (a xor b);
    outputs(4191) <= a and b;
    outputs(4192) <= b and not a;
    outputs(4193) <= a;
    outputs(4194) <= a;
    outputs(4195) <= not (a xor b);
    outputs(4196) <= a xor b;
    outputs(4197) <= a and not b;
    outputs(4198) <= not b;
    outputs(4199) <= not b;
    outputs(4200) <= a;
    outputs(4201) <= b and not a;
    outputs(4202) <= a xor b;
    outputs(4203) <= not (a and b);
    outputs(4204) <= a xor b;
    outputs(4205) <= not a;
    outputs(4206) <= not (a or b);
    outputs(4207) <= a and not b;
    outputs(4208) <= not b;
    outputs(4209) <= a xor b;
    outputs(4210) <= not b;
    outputs(4211) <= a;
    outputs(4212) <= b;
    outputs(4213) <= b;
    outputs(4214) <= a;
    outputs(4215) <= a;
    outputs(4216) <= a xor b;
    outputs(4217) <= a;
    outputs(4218) <= a xor b;
    outputs(4219) <= not b;
    outputs(4220) <= not (a xor b);
    outputs(4221) <= a xor b;
    outputs(4222) <= a;
    outputs(4223) <= not b or a;
    outputs(4224) <= b;
    outputs(4225) <= not (a or b);
    outputs(4226) <= b;
    outputs(4227) <= not (a xor b);
    outputs(4228) <= a;
    outputs(4229) <= a and not b;
    outputs(4230) <= not (a or b);
    outputs(4231) <= a xor b;
    outputs(4232) <= not b;
    outputs(4233) <= not a;
    outputs(4234) <= not b;
    outputs(4235) <= a xor b;
    outputs(4236) <= not (a xor b);
    outputs(4237) <= b and not a;
    outputs(4238) <= b;
    outputs(4239) <= not (a xor b);
    outputs(4240) <= not (a xor b);
    outputs(4241) <= a;
    outputs(4242) <= a;
    outputs(4243) <= not a;
    outputs(4244) <= not (a xor b);
    outputs(4245) <= a xor b;
    outputs(4246) <= not (a xor b);
    outputs(4247) <= a and b;
    outputs(4248) <= not b;
    outputs(4249) <= not (a xor b);
    outputs(4250) <= not b;
    outputs(4251) <= a xor b;
    outputs(4252) <= a;
    outputs(4253) <= not b;
    outputs(4254) <= not (a xor b);
    outputs(4255) <= not (a or b);
    outputs(4256) <= not (a xor b);
    outputs(4257) <= not (a and b);
    outputs(4258) <= not a;
    outputs(4259) <= b and not a;
    outputs(4260) <= a;
    outputs(4261) <= a xor b;
    outputs(4262) <= a;
    outputs(4263) <= a;
    outputs(4264) <= a or b;
    outputs(4265) <= not a;
    outputs(4266) <= not b;
    outputs(4267) <= b and not a;
    outputs(4268) <= a or b;
    outputs(4269) <= not a;
    outputs(4270) <= b;
    outputs(4271) <= a and not b;
    outputs(4272) <= not a or b;
    outputs(4273) <= a;
    outputs(4274) <= a xor b;
    outputs(4275) <= a xor b;
    outputs(4276) <= a or b;
    outputs(4277) <= not (a xor b);
    outputs(4278) <= a xor b;
    outputs(4279) <= not a;
    outputs(4280) <= not a;
    outputs(4281) <= a;
    outputs(4282) <= not b;
    outputs(4283) <= not b;
    outputs(4284) <= a xor b;
    outputs(4285) <= a;
    outputs(4286) <= b;
    outputs(4287) <= not (a or b);
    outputs(4288) <= not b;
    outputs(4289) <= not (a xor b);
    outputs(4290) <= a;
    outputs(4291) <= a and not b;
    outputs(4292) <= not (a xor b);
    outputs(4293) <= not a;
    outputs(4294) <= not b;
    outputs(4295) <= b;
    outputs(4296) <= b and not a;
    outputs(4297) <= not a;
    outputs(4298) <= b;
    outputs(4299) <= not (a and b);
    outputs(4300) <= not (a xor b);
    outputs(4301) <= not b;
    outputs(4302) <= a and b;
    outputs(4303) <= not (a xor b);
    outputs(4304) <= a;
    outputs(4305) <= a and not b;
    outputs(4306) <= not (a xor b);
    outputs(4307) <= not (a xor b);
    outputs(4308) <= b and not a;
    outputs(4309) <= not (a xor b);
    outputs(4310) <= a;
    outputs(4311) <= a and b;
    outputs(4312) <= b and not a;
    outputs(4313) <= not a;
    outputs(4314) <= a xor b;
    outputs(4315) <= not (a and b);
    outputs(4316) <= a or b;
    outputs(4317) <= not a;
    outputs(4318) <= not a;
    outputs(4319) <= not (a xor b);
    outputs(4320) <= a;
    outputs(4321) <= a;
    outputs(4322) <= a or b;
    outputs(4323) <= not b or a;
    outputs(4324) <= not (a or b);
    outputs(4325) <= a;
    outputs(4326) <= b;
    outputs(4327) <= a and not b;
    outputs(4328) <= a and b;
    outputs(4329) <= a;
    outputs(4330) <= a;
    outputs(4331) <= a and not b;
    outputs(4332) <= not (a or b);
    outputs(4333) <= not (a or b);
    outputs(4334) <= not (a xor b);
    outputs(4335) <= a and b;
    outputs(4336) <= not (a xor b);
    outputs(4337) <= a and b;
    outputs(4338) <= not a;
    outputs(4339) <= a xor b;
    outputs(4340) <= a and b;
    outputs(4341) <= b and not a;
    outputs(4342) <= not (a xor b);
    outputs(4343) <= not (a and b);
    outputs(4344) <= not (a xor b);
    outputs(4345) <= a and not b;
    outputs(4346) <= not b;
    outputs(4347) <= a xor b;
    outputs(4348) <= not b;
    outputs(4349) <= not (a xor b);
    outputs(4350) <= b;
    outputs(4351) <= not (a or b);
    outputs(4352) <= not (a xor b);
    outputs(4353) <= not (a xor b);
    outputs(4354) <= a and not b;
    outputs(4355) <= a xor b;
    outputs(4356) <= not a;
    outputs(4357) <= a xor b;
    outputs(4358) <= not (a xor b);
    outputs(4359) <= not (a and b);
    outputs(4360) <= not b;
    outputs(4361) <= b;
    outputs(4362) <= not b;
    outputs(4363) <= b;
    outputs(4364) <= a and b;
    outputs(4365) <= a;
    outputs(4366) <= a and b;
    outputs(4367) <= a;
    outputs(4368) <= not (a xor b);
    outputs(4369) <= not (a xor b);
    outputs(4370) <= a xor b;
    outputs(4371) <= a xor b;
    outputs(4372) <= a and not b;
    outputs(4373) <= a xor b;
    outputs(4374) <= not (a or b);
    outputs(4375) <= not (a xor b);
    outputs(4376) <= a;
    outputs(4377) <= b;
    outputs(4378) <= a xor b;
    outputs(4379) <= not (a xor b);
    outputs(4380) <= not (a xor b);
    outputs(4381) <= b and not a;
    outputs(4382) <= b;
    outputs(4383) <= b and not a;
    outputs(4384) <= not (a or b);
    outputs(4385) <= a;
    outputs(4386) <= a or b;
    outputs(4387) <= a;
    outputs(4388) <= not (a xor b);
    outputs(4389) <= not a;
    outputs(4390) <= b;
    outputs(4391) <= b and not a;
    outputs(4392) <= not a;
    outputs(4393) <= a and not b;
    outputs(4394) <= not a or b;
    outputs(4395) <= not a;
    outputs(4396) <= a;
    outputs(4397) <= a and not b;
    outputs(4398) <= a and b;
    outputs(4399) <= b;
    outputs(4400) <= not (a xor b);
    outputs(4401) <= a xor b;
    outputs(4402) <= b;
    outputs(4403) <= not (a xor b);
    outputs(4404) <= not (a xor b);
    outputs(4405) <= not (a xor b);
    outputs(4406) <= not (a or b);
    outputs(4407) <= not a;
    outputs(4408) <= a xor b;
    outputs(4409) <= not (a xor b);
    outputs(4410) <= not b or a;
    outputs(4411) <= a and not b;
    outputs(4412) <= a or b;
    outputs(4413) <= a;
    outputs(4414) <= a and not b;
    outputs(4415) <= not a;
    outputs(4416) <= b;
    outputs(4417) <= not b;
    outputs(4418) <= not a;
    outputs(4419) <= not a;
    outputs(4420) <= b;
    outputs(4421) <= b;
    outputs(4422) <= not (a xor b);
    outputs(4423) <= '0';
    outputs(4424) <= a or b;
    outputs(4425) <= b and not a;
    outputs(4426) <= a xor b;
    outputs(4427) <= not (a xor b);
    outputs(4428) <= not b;
    outputs(4429) <= a or b;
    outputs(4430) <= not (a or b);
    outputs(4431) <= not b;
    outputs(4432) <= a xor b;
    outputs(4433) <= not b;
    outputs(4434) <= b and not a;
    outputs(4435) <= a and not b;
    outputs(4436) <= not a;
    outputs(4437) <= a;
    outputs(4438) <= b and not a;
    outputs(4439) <= not b;
    outputs(4440) <= b;
    outputs(4441) <= not a;
    outputs(4442) <= not a;
    outputs(4443) <= not b;
    outputs(4444) <= a and b;
    outputs(4445) <= b and not a;
    outputs(4446) <= a xor b;
    outputs(4447) <= not (a xor b);
    outputs(4448) <= a and not b;
    outputs(4449) <= b;
    outputs(4450) <= not (a xor b);
    outputs(4451) <= not a;
    outputs(4452) <= not (a or b);
    outputs(4453) <= not (a xor b);
    outputs(4454) <= a xor b;
    outputs(4455) <= not a;
    outputs(4456) <= a xor b;
    outputs(4457) <= b and not a;
    outputs(4458) <= not b or a;
    outputs(4459) <= b;
    outputs(4460) <= a xor b;
    outputs(4461) <= a xor b;
    outputs(4462) <= not b or a;
    outputs(4463) <= not b or a;
    outputs(4464) <= a;
    outputs(4465) <= not b;
    outputs(4466) <= a and not b;
    outputs(4467) <= a;
    outputs(4468) <= b and not a;
    outputs(4469) <= b;
    outputs(4470) <= a;
    outputs(4471) <= not a;
    outputs(4472) <= a xor b;
    outputs(4473) <= not a;
    outputs(4474) <= b and not a;
    outputs(4475) <= not b;
    outputs(4476) <= not (a xor b);
    outputs(4477) <= not a;
    outputs(4478) <= b and not a;
    outputs(4479) <= b;
    outputs(4480) <= b;
    outputs(4481) <= not (a xor b);
    outputs(4482) <= a xor b;
    outputs(4483) <= not b;
    outputs(4484) <= not b;
    outputs(4485) <= not a;
    outputs(4486) <= not a;
    outputs(4487) <= not a;
    outputs(4488) <= a xor b;
    outputs(4489) <= not (a xor b);
    outputs(4490) <= a xor b;
    outputs(4491) <= not (a or b);
    outputs(4492) <= a xor b;
    outputs(4493) <= not a;
    outputs(4494) <= not a;
    outputs(4495) <= not (a or b);
    outputs(4496) <= a xor b;
    outputs(4497) <= a and not b;
    outputs(4498) <= a xor b;
    outputs(4499) <= a and not b;
    outputs(4500) <= not b;
    outputs(4501) <= not (a xor b);
    outputs(4502) <= a and b;
    outputs(4503) <= b;
    outputs(4504) <= a and b;
    outputs(4505) <= not (a and b);
    outputs(4506) <= not (a xor b);
    outputs(4507) <= a and not b;
    outputs(4508) <= not b;
    outputs(4509) <= not a;
    outputs(4510) <= not b;
    outputs(4511) <= not (a and b);
    outputs(4512) <= not b;
    outputs(4513) <= not (a xor b);
    outputs(4514) <= a;
    outputs(4515) <= a and b;
    outputs(4516) <= a and b;
    outputs(4517) <= a xor b;
    outputs(4518) <= a;
    outputs(4519) <= not (a or b);
    outputs(4520) <= a;
    outputs(4521) <= a and not b;
    outputs(4522) <= not (a and b);
    outputs(4523) <= not (a xor b);
    outputs(4524) <= not (a xor b);
    outputs(4525) <= not a;
    outputs(4526) <= a and not b;
    outputs(4527) <= a;
    outputs(4528) <= b;
    outputs(4529) <= a;
    outputs(4530) <= not a;
    outputs(4531) <= a;
    outputs(4532) <= not (a and b);
    outputs(4533) <= not a;
    outputs(4534) <= a;
    outputs(4535) <= not b;
    outputs(4536) <= not (a xor b);
    outputs(4537) <= a xor b;
    outputs(4538) <= not (a xor b);
    outputs(4539) <= not b;
    outputs(4540) <= not (a xor b);
    outputs(4541) <= a and b;
    outputs(4542) <= a xor b;
    outputs(4543) <= a xor b;
    outputs(4544) <= a;
    outputs(4545) <= a xor b;
    outputs(4546) <= b;
    outputs(4547) <= b;
    outputs(4548) <= not a;
    outputs(4549) <= b;
    outputs(4550) <= a xor b;
    outputs(4551) <= not b;
    outputs(4552) <= not b;
    outputs(4553) <= b;
    outputs(4554) <= b;
    outputs(4555) <= a and b;
    outputs(4556) <= a and b;
    outputs(4557) <= not (a and b);
    outputs(4558) <= a xor b;
    outputs(4559) <= not b;
    outputs(4560) <= not a or b;
    outputs(4561) <= a;
    outputs(4562) <= not b;
    outputs(4563) <= a and b;
    outputs(4564) <= not b or a;
    outputs(4565) <= not (a or b);
    outputs(4566) <= a xor b;
    outputs(4567) <= a and b;
    outputs(4568) <= a;
    outputs(4569) <= a;
    outputs(4570) <= a;
    outputs(4571) <= not a or b;
    outputs(4572) <= not b;
    outputs(4573) <= a xor b;
    outputs(4574) <= not (a xor b);
    outputs(4575) <= not (a xor b);
    outputs(4576) <= a xor b;
    outputs(4577) <= not a;
    outputs(4578) <= a xor b;
    outputs(4579) <= not b;
    outputs(4580) <= b;
    outputs(4581) <= b and not a;
    outputs(4582) <= not (a xor b);
    outputs(4583) <= a xor b;
    outputs(4584) <= not (a xor b);
    outputs(4585) <= not (a xor b);
    outputs(4586) <= not b;
    outputs(4587) <= b;
    outputs(4588) <= a and b;
    outputs(4589) <= a xor b;
    outputs(4590) <= b and not a;
    outputs(4591) <= not a;
    outputs(4592) <= b;
    outputs(4593) <= a;
    outputs(4594) <= b and not a;
    outputs(4595) <= not b or a;
    outputs(4596) <= a;
    outputs(4597) <= a xor b;
    outputs(4598) <= not a;
    outputs(4599) <= not (a xor b);
    outputs(4600) <= a;
    outputs(4601) <= a and b;
    outputs(4602) <= not a;
    outputs(4603) <= not b;
    outputs(4604) <= not (a xor b);
    outputs(4605) <= not b;
    outputs(4606) <= not a;
    outputs(4607) <= a xor b;
    outputs(4608) <= not (a xor b);
    outputs(4609) <= not b;
    outputs(4610) <= a xor b;
    outputs(4611) <= not (a or b);
    outputs(4612) <= b;
    outputs(4613) <= a and not b;
    outputs(4614) <= a and not b;
    outputs(4615) <= not (a xor b);
    outputs(4616) <= a and not b;
    outputs(4617) <= b;
    outputs(4618) <= not b;
    outputs(4619) <= a and b;
    outputs(4620) <= b and not a;
    outputs(4621) <= a and b;
    outputs(4622) <= b;
    outputs(4623) <= a xor b;
    outputs(4624) <= a and b;
    outputs(4625) <= a and b;
    outputs(4626) <= a;
    outputs(4627) <= a;
    outputs(4628) <= b and not a;
    outputs(4629) <= not a;
    outputs(4630) <= not (a xor b);
    outputs(4631) <= a and not b;
    outputs(4632) <= not (a or b);
    outputs(4633) <= not b;
    outputs(4634) <= not (a xor b);
    outputs(4635) <= a or b;
    outputs(4636) <= a and not b;
    outputs(4637) <= a and not b;
    outputs(4638) <= not (a or b);
    outputs(4639) <= not b;
    outputs(4640) <= not a;
    outputs(4641) <= b and not a;
    outputs(4642) <= not a;
    outputs(4643) <= not (a xor b);
    outputs(4644) <= a or b;
    outputs(4645) <= not b;
    outputs(4646) <= not (a or b);
    outputs(4647) <= a;
    outputs(4648) <= not (a or b);
    outputs(4649) <= not a;
    outputs(4650) <= not a;
    outputs(4651) <= b;
    outputs(4652) <= a and b;
    outputs(4653) <= not (a xor b);
    outputs(4654) <= not b;
    outputs(4655) <= a and not b;
    outputs(4656) <= a and b;
    outputs(4657) <= not (a xor b);
    outputs(4658) <= b;
    outputs(4659) <= not a;
    outputs(4660) <= not (a and b);
    outputs(4661) <= a and b;
    outputs(4662) <= a;
    outputs(4663) <= not b or a;
    outputs(4664) <= not b;
    outputs(4665) <= a;
    outputs(4666) <= not b;
    outputs(4667) <= a and not b;
    outputs(4668) <= not a;
    outputs(4669) <= not (a and b);
    outputs(4670) <= not b;
    outputs(4671) <= not (a or b);
    outputs(4672) <= not (a xor b);
    outputs(4673) <= a xor b;
    outputs(4674) <= not a;
    outputs(4675) <= not a;
    outputs(4676) <= a;
    outputs(4677) <= not a;
    outputs(4678) <= not (a xor b);
    outputs(4679) <= a xor b;
    outputs(4680) <= b;
    outputs(4681) <= a xor b;
    outputs(4682) <= a xor b;
    outputs(4683) <= not (a xor b);
    outputs(4684) <= not a;
    outputs(4685) <= not (a and b);
    outputs(4686) <= a;
    outputs(4687) <= not (a or b);
    outputs(4688) <= not a or b;
    outputs(4689) <= a and not b;
    outputs(4690) <= not b;
    outputs(4691) <= b and not a;
    outputs(4692) <= not a or b;
    outputs(4693) <= not (a or b);
    outputs(4694) <= not a;
    outputs(4695) <= not (a xor b);
    outputs(4696) <= not (a xor b);
    outputs(4697) <= not a;
    outputs(4698) <= a and not b;
    outputs(4699) <= not a;
    outputs(4700) <= not (a or b);
    outputs(4701) <= not b;
    outputs(4702) <= a and b;
    outputs(4703) <= b and not a;
    outputs(4704) <= not b;
    outputs(4705) <= not (a xor b);
    outputs(4706) <= a and not b;
    outputs(4707) <= not (a or b);
    outputs(4708) <= b;
    outputs(4709) <= not (a or b);
    outputs(4710) <= b;
    outputs(4711) <= not a;
    outputs(4712) <= not b;
    outputs(4713) <= a xor b;
    outputs(4714) <= b;
    outputs(4715) <= a and not b;
    outputs(4716) <= not a;
    outputs(4717) <= a xor b;
    outputs(4718) <= not (a xor b);
    outputs(4719) <= a;
    outputs(4720) <= a xor b;
    outputs(4721) <= a xor b;
    outputs(4722) <= a xor b;
    outputs(4723) <= a xor b;
    outputs(4724) <= not (a xor b);
    outputs(4725) <= not a;
    outputs(4726) <= b;
    outputs(4727) <= not (a or b);
    outputs(4728) <= not (a xor b);
    outputs(4729) <= not a;
    outputs(4730) <= not b;
    outputs(4731) <= a xor b;
    outputs(4732) <= not (a xor b);
    outputs(4733) <= a xor b;
    outputs(4734) <= not (a xor b);
    outputs(4735) <= not a;
    outputs(4736) <= a and not b;
    outputs(4737) <= b;
    outputs(4738) <= not b;
    outputs(4739) <= a;
    outputs(4740) <= b;
    outputs(4741) <= not (a or b);
    outputs(4742) <= not (a xor b);
    outputs(4743) <= a and b;
    outputs(4744) <= b and not a;
    outputs(4745) <= not a;
    outputs(4746) <= not (a xor b);
    outputs(4747) <= a and not b;
    outputs(4748) <= not a;
    outputs(4749) <= a and not b;
    outputs(4750) <= not a or b;
    outputs(4751) <= not a;
    outputs(4752) <= not (a or b);
    outputs(4753) <= not (a xor b);
    outputs(4754) <= a or b;
    outputs(4755) <= not (a or b);
    outputs(4756) <= not a;
    outputs(4757) <= not b or a;
    outputs(4758) <= not b;
    outputs(4759) <= not a;
    outputs(4760) <= b;
    outputs(4761) <= b;
    outputs(4762) <= not (a xor b);
    outputs(4763) <= not (a xor b);
    outputs(4764) <= a xor b;
    outputs(4765) <= a xor b;
    outputs(4766) <= not b;
    outputs(4767) <= not a;
    outputs(4768) <= b;
    outputs(4769) <= not (a or b);
    outputs(4770) <= not a;
    outputs(4771) <= a;
    outputs(4772) <= not (a xor b);
    outputs(4773) <= not b;
    outputs(4774) <= a;
    outputs(4775) <= not (a and b);
    outputs(4776) <= not (a xor b);
    outputs(4777) <= not b;
    outputs(4778) <= a;
    outputs(4779) <= not b;
    outputs(4780) <= not a;
    outputs(4781) <= b and not a;
    outputs(4782) <= a and not b;
    outputs(4783) <= not a;
    outputs(4784) <= a and b;
    outputs(4785) <= b and not a;
    outputs(4786) <= not (a or b);
    outputs(4787) <= not (a or b);
    outputs(4788) <= a and b;
    outputs(4789) <= a;
    outputs(4790) <= b and not a;
    outputs(4791) <= a and not b;
    outputs(4792) <= a and not b;
    outputs(4793) <= not (a xor b);
    outputs(4794) <= a;
    outputs(4795) <= b;
    outputs(4796) <= not a;
    outputs(4797) <= not a;
    outputs(4798) <= b;
    outputs(4799) <= not (a and b);
    outputs(4800) <= a or b;
    outputs(4801) <= a xor b;
    outputs(4802) <= not a;
    outputs(4803) <= not a;
    outputs(4804) <= b;
    outputs(4805) <= a xor b;
    outputs(4806) <= not (a or b);
    outputs(4807) <= a and b;
    outputs(4808) <= b;
    outputs(4809) <= b and not a;
    outputs(4810) <= a xor b;
    outputs(4811) <= not a;
    outputs(4812) <= not (a or b);
    outputs(4813) <= not b;
    outputs(4814) <= a or b;
    outputs(4815) <= a xor b;
    outputs(4816) <= not (a xor b);
    outputs(4817) <= not b;
    outputs(4818) <= not (a xor b);
    outputs(4819) <= a xor b;
    outputs(4820) <= a;
    outputs(4821) <= b and not a;
    outputs(4822) <= b;
    outputs(4823) <= a xor b;
    outputs(4824) <= not b;
    outputs(4825) <= not (a xor b);
    outputs(4826) <= not (a xor b);
    outputs(4827) <= a xor b;
    outputs(4828) <= a xor b;
    outputs(4829) <= a and not b;
    outputs(4830) <= b;
    outputs(4831) <= a and not b;
    outputs(4832) <= a xor b;
    outputs(4833) <= b;
    outputs(4834) <= a;
    outputs(4835) <= not (a xor b);
    outputs(4836) <= not b or a;
    outputs(4837) <= not (a or b);
    outputs(4838) <= not (a or b);
    outputs(4839) <= a;
    outputs(4840) <= not b;
    outputs(4841) <= a;
    outputs(4842) <= b;
    outputs(4843) <= not (a or b);
    outputs(4844) <= not (a xor b);
    outputs(4845) <= a or b;
    outputs(4846) <= not a;
    outputs(4847) <= b and not a;
    outputs(4848) <= b;
    outputs(4849) <= not (a and b);
    outputs(4850) <= a xor b;
    outputs(4851) <= not a;
    outputs(4852) <= a;
    outputs(4853) <= a;
    outputs(4854) <= a and b;
    outputs(4855) <= a and not b;
    outputs(4856) <= not (a or b);
    outputs(4857) <= a;
    outputs(4858) <= not a;
    outputs(4859) <= b;
    outputs(4860) <= a xor b;
    outputs(4861) <= a;
    outputs(4862) <= a and not b;
    outputs(4863) <= not a;
    outputs(4864) <= not b;
    outputs(4865) <= b;
    outputs(4866) <= not a;
    outputs(4867) <= not (a or b);
    outputs(4868) <= b;
    outputs(4869) <= a xor b;
    outputs(4870) <= a;
    outputs(4871) <= not a;
    outputs(4872) <= b;
    outputs(4873) <= a and not b;
    outputs(4874) <= not (a or b);
    outputs(4875) <= not a;
    outputs(4876) <= not a;
    outputs(4877) <= not b;
    outputs(4878) <= not b;
    outputs(4879) <= not b;
    outputs(4880) <= a;
    outputs(4881) <= not (a xor b);
    outputs(4882) <= a and not b;
    outputs(4883) <= a xor b;
    outputs(4884) <= not b;
    outputs(4885) <= not b;
    outputs(4886) <= a and not b;
    outputs(4887) <= not (a xor b);
    outputs(4888) <= b;
    outputs(4889) <= b;
    outputs(4890) <= not b;
    outputs(4891) <= not (a xor b);
    outputs(4892) <= not a;
    outputs(4893) <= not b;
    outputs(4894) <= a and b;
    outputs(4895) <= not (a xor b);
    outputs(4896) <= not a;
    outputs(4897) <= not (a xor b);
    outputs(4898) <= not (a xor b);
    outputs(4899) <= b;
    outputs(4900) <= not a;
    outputs(4901) <= a and b;
    outputs(4902) <= not b or a;
    outputs(4903) <= a;
    outputs(4904) <= not (a xor b);
    outputs(4905) <= a or b;
    outputs(4906) <= a or b;
    outputs(4907) <= a xor b;
    outputs(4908) <= a and b;
    outputs(4909) <= not (a or b);
    outputs(4910) <= not (a or b);
    outputs(4911) <= not b or a;
    outputs(4912) <= not a or b;
    outputs(4913) <= a and b;
    outputs(4914) <= a xor b;
    outputs(4915) <= a xor b;
    outputs(4916) <= a;
    outputs(4917) <= b and not a;
    outputs(4918) <= a xor b;
    outputs(4919) <= a;
    outputs(4920) <= not b;
    outputs(4921) <= b;
    outputs(4922) <= a xor b;
    outputs(4923) <= a xor b;
    outputs(4924) <= not (a or b);
    outputs(4925) <= a xor b;
    outputs(4926) <= not b;
    outputs(4927) <= b;
    outputs(4928) <= a or b;
    outputs(4929) <= b;
    outputs(4930) <= a xor b;
    outputs(4931) <= not (a or b);
    outputs(4932) <= a;
    outputs(4933) <= not b;
    outputs(4934) <= not (a xor b);
    outputs(4935) <= b;
    outputs(4936) <= not b;
    outputs(4937) <= a xor b;
    outputs(4938) <= not (a xor b);
    outputs(4939) <= a;
    outputs(4940) <= a xor b;
    outputs(4941) <= not b;
    outputs(4942) <= not (a or b);
    outputs(4943) <= not b;
    outputs(4944) <= not a;
    outputs(4945) <= a;
    outputs(4946) <= not b or a;
    outputs(4947) <= a;
    outputs(4948) <= not b;
    outputs(4949) <= not b;
    outputs(4950) <= a xor b;
    outputs(4951) <= a;
    outputs(4952) <= a;
    outputs(4953) <= a;
    outputs(4954) <= not (a xor b);
    outputs(4955) <= a xor b;
    outputs(4956) <= a and not b;
    outputs(4957) <= not (a or b);
    outputs(4958) <= a xor b;
    outputs(4959) <= a;
    outputs(4960) <= b and not a;
    outputs(4961) <= a;
    outputs(4962) <= not b;
    outputs(4963) <= a xor b;
    outputs(4964) <= b and not a;
    outputs(4965) <= b;
    outputs(4966) <= b and not a;
    outputs(4967) <= a;
    outputs(4968) <= a xor b;
    outputs(4969) <= a;
    outputs(4970) <= b;
    outputs(4971) <= a and not b;
    outputs(4972) <= a and not b;
    outputs(4973) <= b and not a;
    outputs(4974) <= not (a xor b);
    outputs(4975) <= b;
    outputs(4976) <= a;
    outputs(4977) <= not (a xor b);
    outputs(4978) <= a and not b;
    outputs(4979) <= not (a xor b);
    outputs(4980) <= not a;
    outputs(4981) <= not b;
    outputs(4982) <= not a or b;
    outputs(4983) <= not b;
    outputs(4984) <= not b or a;
    outputs(4985) <= b;
    outputs(4986) <= b;
    outputs(4987) <= not a;
    outputs(4988) <= a and b;
    outputs(4989) <= b and not a;
    outputs(4990) <= not a;
    outputs(4991) <= a;
    outputs(4992) <= a and not b;
    outputs(4993) <= not (a xor b);
    outputs(4994) <= not (a xor b);
    outputs(4995) <= b;
    outputs(4996) <= not a;
    outputs(4997) <= not (a xor b);
    outputs(4998) <= not a;
    outputs(4999) <= b;
    outputs(5000) <= a and not b;
    outputs(5001) <= not a;
    outputs(5002) <= a xor b;
    outputs(5003) <= a or b;
    outputs(5004) <= b;
    outputs(5005) <= a and b;
    outputs(5006) <= a xor b;
    outputs(5007) <= not (a xor b);
    outputs(5008) <= a xor b;
    outputs(5009) <= not (a xor b);
    outputs(5010) <= not b;
    outputs(5011) <= not (a or b);
    outputs(5012) <= b and not a;
    outputs(5013) <= not (a xor b);
    outputs(5014) <= a and not b;
    outputs(5015) <= not (a or b);
    outputs(5016) <= not a;
    outputs(5017) <= not (a xor b);
    outputs(5018) <= a xor b;
    outputs(5019) <= a or b;
    outputs(5020) <= not a;
    outputs(5021) <= b and not a;
    outputs(5022) <= a;
    outputs(5023) <= not b;
    outputs(5024) <= not a;
    outputs(5025) <= b and not a;
    outputs(5026) <= b;
    outputs(5027) <= not b or a;
    outputs(5028) <= not (a xor b);
    outputs(5029) <= a xor b;
    outputs(5030) <= not b;
    outputs(5031) <= a;
    outputs(5032) <= not (a xor b);
    outputs(5033) <= a;
    outputs(5034) <= not (a xor b);
    outputs(5035) <= a;
    outputs(5036) <= not b;
    outputs(5037) <= not a;
    outputs(5038) <= not (a and b);
    outputs(5039) <= a;
    outputs(5040) <= b;
    outputs(5041) <= not a;
    outputs(5042) <= b;
    outputs(5043) <= a;
    outputs(5044) <= not a;
    outputs(5045) <= a xor b;
    outputs(5046) <= a;
    outputs(5047) <= not (a or b);
    outputs(5048) <= a and b;
    outputs(5049) <= a;
    outputs(5050) <= a;
    outputs(5051) <= a;
    outputs(5052) <= not (a xor b);
    outputs(5053) <= a and not b;
    outputs(5054) <= not a;
    outputs(5055) <= a;
    outputs(5056) <= not b;
    outputs(5057) <= not (a xor b);
    outputs(5058) <= not (a or b);
    outputs(5059) <= a or b;
    outputs(5060) <= b;
    outputs(5061) <= a xor b;
    outputs(5062) <= a;
    outputs(5063) <= b;
    outputs(5064) <= a xor b;
    outputs(5065) <= a xor b;
    outputs(5066) <= not (a xor b);
    outputs(5067) <= b;
    outputs(5068) <= not b;
    outputs(5069) <= not b or a;
    outputs(5070) <= not b;
    outputs(5071) <= not (a xor b);
    outputs(5072) <= a;
    outputs(5073) <= b;
    outputs(5074) <= a;
    outputs(5075) <= a xor b;
    outputs(5076) <= a and not b;
    outputs(5077) <= not (a xor b);
    outputs(5078) <= not a;
    outputs(5079) <= not a or b;
    outputs(5080) <= not (a xor b);
    outputs(5081) <= a and not b;
    outputs(5082) <= b and not a;
    outputs(5083) <= b;
    outputs(5084) <= not (a and b);
    outputs(5085) <= not a;
    outputs(5086) <= a xor b;
    outputs(5087) <= a xor b;
    outputs(5088) <= not a;
    outputs(5089) <= not b;
    outputs(5090) <= a and b;
    outputs(5091) <= not (a xor b);
    outputs(5092) <= not a;
    outputs(5093) <= not (a xor b);
    outputs(5094) <= b;
    outputs(5095) <= b and not a;
    outputs(5096) <= not (a xor b);
    outputs(5097) <= a xor b;
    outputs(5098) <= b;
    outputs(5099) <= a;
    outputs(5100) <= not (a xor b);
    outputs(5101) <= a xor b;
    outputs(5102) <= a xor b;
    outputs(5103) <= not a;
    outputs(5104) <= b;
    outputs(5105) <= b and not a;
    outputs(5106) <= a;
    outputs(5107) <= a xor b;
    outputs(5108) <= not a;
    outputs(5109) <= a or b;
    outputs(5110) <= a;
    outputs(5111) <= a;
    outputs(5112) <= a;
    outputs(5113) <= b and not a;
    outputs(5114) <= a or b;
    outputs(5115) <= not (a and b);
    outputs(5116) <= b;
    outputs(5117) <= not b;
    outputs(5118) <= not (a xor b);
    outputs(5119) <= not a;
    outputs(5120) <= b and not a;
    outputs(5121) <= not a or b;
    outputs(5122) <= a xor b;
    outputs(5123) <= not (a or b);
    outputs(5124) <= a xor b;
    outputs(5125) <= a xor b;
    outputs(5126) <= not b or a;
    outputs(5127) <= b and not a;
    outputs(5128) <= not b or a;
    outputs(5129) <= a xor b;
    outputs(5130) <= not (a and b);
    outputs(5131) <= b;
    outputs(5132) <= a xor b;
    outputs(5133) <= not a or b;
    outputs(5134) <= a;
    outputs(5135) <= a;
    outputs(5136) <= a and not b;
    outputs(5137) <= not (a xor b);
    outputs(5138) <= a xor b;
    outputs(5139) <= not (a and b);
    outputs(5140) <= a;
    outputs(5141) <= not b;
    outputs(5142) <= a;
    outputs(5143) <= not b;
    outputs(5144) <= not (a xor b);
    outputs(5145) <= a and b;
    outputs(5146) <= not (a or b);
    outputs(5147) <= not b;
    outputs(5148) <= a xor b;
    outputs(5149) <= not (a xor b);
    outputs(5150) <= a;
    outputs(5151) <= a xor b;
    outputs(5152) <= not a or b;
    outputs(5153) <= b and not a;
    outputs(5154) <= not a;
    outputs(5155) <= not b;
    outputs(5156) <= not a;
    outputs(5157) <= not a;
    outputs(5158) <= not a;
    outputs(5159) <= a and not b;
    outputs(5160) <= a and b;
    outputs(5161) <= b;
    outputs(5162) <= b and not a;
    outputs(5163) <= not (a xor b);
    outputs(5164) <= not (a and b);
    outputs(5165) <= a xor b;
    outputs(5166) <= not (a xor b);
    outputs(5167) <= not a;
    outputs(5168) <= a xor b;
    outputs(5169) <= a or b;
    outputs(5170) <= a;
    outputs(5171) <= not b or a;
    outputs(5172) <= not (a and b);
    outputs(5173) <= not (a xor b);
    outputs(5174) <= a xor b;
    outputs(5175) <= not (a or b);
    outputs(5176) <= not b;
    outputs(5177) <= not a;
    outputs(5178) <= not a;
    outputs(5179) <= not b;
    outputs(5180) <= not a;
    outputs(5181) <= a and not b;
    outputs(5182) <= not (a and b);
    outputs(5183) <= not b;
    outputs(5184) <= not a;
    outputs(5185) <= a xor b;
    outputs(5186) <= not (a and b);
    outputs(5187) <= a or b;
    outputs(5188) <= not (a xor b);
    outputs(5189) <= a xor b;
    outputs(5190) <= a;
    outputs(5191) <= not a;
    outputs(5192) <= not b;
    outputs(5193) <= b;
    outputs(5194) <= not (a or b);
    outputs(5195) <= a and b;
    outputs(5196) <= a or b;
    outputs(5197) <= a;
    outputs(5198) <= a or b;
    outputs(5199) <= not (a xor b);
    outputs(5200) <= a xor b;
    outputs(5201) <= a xor b;
    outputs(5202) <= a xor b;
    outputs(5203) <= not a;
    outputs(5204) <= not a or b;
    outputs(5205) <= not a;
    outputs(5206) <= not (a xor b);
    outputs(5207) <= not (a xor b);
    outputs(5208) <= not (a xor b);
    outputs(5209) <= not (a xor b);
    outputs(5210) <= not (a xor b);
    outputs(5211) <= a and not b;
    outputs(5212) <= b;
    outputs(5213) <= not (a xor b);
    outputs(5214) <= not (a xor b);
    outputs(5215) <= not (a xor b);
    outputs(5216) <= a;
    outputs(5217) <= not a;
    outputs(5218) <= not b;
    outputs(5219) <= a xor b;
    outputs(5220) <= a xor b;
    outputs(5221) <= not a;
    outputs(5222) <= a;
    outputs(5223) <= not (a xor b);
    outputs(5224) <= not a;
    outputs(5225) <= not b;
    outputs(5226) <= a xor b;
    outputs(5227) <= not a;
    outputs(5228) <= not b;
    outputs(5229) <= b;
    outputs(5230) <= not a;
    outputs(5231) <= b;
    outputs(5232) <= not (a xor b);
    outputs(5233) <= a xor b;
    outputs(5234) <= a and b;
    outputs(5235) <= not a;
    outputs(5236) <= b and not a;
    outputs(5237) <= not b;
    outputs(5238) <= not (a and b);
    outputs(5239) <= not (a or b);
    outputs(5240) <= not a;
    outputs(5241) <= b;
    outputs(5242) <= not a;
    outputs(5243) <= a xor b;
    outputs(5244) <= not b;
    outputs(5245) <= not (a xor b);
    outputs(5246) <= not (a xor b);
    outputs(5247) <= b;
    outputs(5248) <= not b or a;
    outputs(5249) <= b;
    outputs(5250) <= b;
    outputs(5251) <= a xor b;
    outputs(5252) <= not a or b;
    outputs(5253) <= b;
    outputs(5254) <= b;
    outputs(5255) <= not a;
    outputs(5256) <= a;
    outputs(5257) <= not a;
    outputs(5258) <= a xor b;
    outputs(5259) <= a xor b;
    outputs(5260) <= b;
    outputs(5261) <= a and b;
    outputs(5262) <= not (a xor b);
    outputs(5263) <= a xor b;
    outputs(5264) <= a xor b;
    outputs(5265) <= not a;
    outputs(5266) <= not b;
    outputs(5267) <= not a;
    outputs(5268) <= not a;
    outputs(5269) <= not a or b;
    outputs(5270) <= a or b;
    outputs(5271) <= a xor b;
    outputs(5272) <= a;
    outputs(5273) <= b;
    outputs(5274) <= b;
    outputs(5275) <= not (a or b);
    outputs(5276) <= not (a xor b);
    outputs(5277) <= not (a xor b);
    outputs(5278) <= a xor b;
    outputs(5279) <= not a or b;
    outputs(5280) <= not a;
    outputs(5281) <= b and not a;
    outputs(5282) <= not b;
    outputs(5283) <= a xor b;
    outputs(5284) <= a xor b;
    outputs(5285) <= a xor b;
    outputs(5286) <= a xor b;
    outputs(5287) <= b;
    outputs(5288) <= a xor b;
    outputs(5289) <= a and not b;
    outputs(5290) <= a xor b;
    outputs(5291) <= a or b;
    outputs(5292) <= a xor b;
    outputs(5293) <= not b;
    outputs(5294) <= a xor b;
    outputs(5295) <= not a;
    outputs(5296) <= not (a or b);
    outputs(5297) <= a and not b;
    outputs(5298) <= not (a xor b);
    outputs(5299) <= b and not a;
    outputs(5300) <= a xor b;
    outputs(5301) <= not b or a;
    outputs(5302) <= a xor b;
    outputs(5303) <= a xor b;
    outputs(5304) <= b;
    outputs(5305) <= not (a or b);
    outputs(5306) <= a xor b;
    outputs(5307) <= a xor b;
    outputs(5308) <= not (a xor b);
    outputs(5309) <= not (a and b);
    outputs(5310) <= not (a xor b);
    outputs(5311) <= b and not a;
    outputs(5312) <= not b;
    outputs(5313) <= not (a xor b);
    outputs(5314) <= not b;
    outputs(5315) <= not (a xor b);
    outputs(5316) <= not (a xor b);
    outputs(5317) <= not a;
    outputs(5318) <= b and not a;
    outputs(5319) <= a xor b;
    outputs(5320) <= not a;
    outputs(5321) <= not a or b;
    outputs(5322) <= a;
    outputs(5323) <= not (a xor b);
    outputs(5324) <= a xor b;
    outputs(5325) <= a and b;
    outputs(5326) <= not (a and b);
    outputs(5327) <= not a or b;
    outputs(5328) <= b and not a;
    outputs(5329) <= a xor b;
    outputs(5330) <= b and not a;
    outputs(5331) <= a xor b;
    outputs(5332) <= a;
    outputs(5333) <= not a or b;
    outputs(5334) <= not a;
    outputs(5335) <= a xor b;
    outputs(5336) <= not a;
    outputs(5337) <= not (a and b);
    outputs(5338) <= a xor b;
    outputs(5339) <= not b;
    outputs(5340) <= not b or a;
    outputs(5341) <= not (a xor b);
    outputs(5342) <= b;
    outputs(5343) <= a xor b;
    outputs(5344) <= b;
    outputs(5345) <= a xor b;
    outputs(5346) <= not (a xor b);
    outputs(5347) <= not b;
    outputs(5348) <= a xor b;
    outputs(5349) <= a xor b;
    outputs(5350) <= a or b;
    outputs(5351) <= not (a xor b);
    outputs(5352) <= not a;
    outputs(5353) <= not b;
    outputs(5354) <= not (a xor b);
    outputs(5355) <= not (a xor b);
    outputs(5356) <= not (a and b);
    outputs(5357) <= b;
    outputs(5358) <= not (a xor b);
    outputs(5359) <= a xor b;
    outputs(5360) <= not b;
    outputs(5361) <= a xor b;
    outputs(5362) <= a;
    outputs(5363) <= not b;
    outputs(5364) <= a xor b;
    outputs(5365) <= not b;
    outputs(5366) <= not b;
    outputs(5367) <= not a;
    outputs(5368) <= a;
    outputs(5369) <= b and not a;
    outputs(5370) <= a xor b;
    outputs(5371) <= not b;
    outputs(5372) <= a or b;
    outputs(5373) <= not a;
    outputs(5374) <= b and not a;
    outputs(5375) <= not (a xor b);
    outputs(5376) <= not (a or b);
    outputs(5377) <= not b;
    outputs(5378) <= a xor b;
    outputs(5379) <= b and not a;
    outputs(5380) <= not (a xor b);
    outputs(5381) <= not (a xor b);
    outputs(5382) <= not (a or b);
    outputs(5383) <= not b;
    outputs(5384) <= not a;
    outputs(5385) <= not (a xor b);
    outputs(5386) <= not a;
    outputs(5387) <= not a;
    outputs(5388) <= not (a xor b);
    outputs(5389) <= b and not a;
    outputs(5390) <= not a or b;
    outputs(5391) <= not (a and b);
    outputs(5392) <= a and b;
    outputs(5393) <= b;
    outputs(5394) <= b and not a;
    outputs(5395) <= a xor b;
    outputs(5396) <= a;
    outputs(5397) <= not (a or b);
    outputs(5398) <= a xor b;
    outputs(5399) <= a;
    outputs(5400) <= a;
    outputs(5401) <= a xor b;
    outputs(5402) <= not (a or b);
    outputs(5403) <= a xor b;
    outputs(5404) <= not (a xor b);
    outputs(5405) <= not (a and b);
    outputs(5406) <= not b or a;
    outputs(5407) <= not (a xor b);
    outputs(5408) <= a xor b;
    outputs(5409) <= not (a or b);
    outputs(5410) <= b;
    outputs(5411) <= not a;
    outputs(5412) <= not (a xor b);
    outputs(5413) <= not a;
    outputs(5414) <= not (a xor b);
    outputs(5415) <= a xor b;
    outputs(5416) <= a xor b;
    outputs(5417) <= b and not a;
    outputs(5418) <= not b or a;
    outputs(5419) <= a;
    outputs(5420) <= not a;
    outputs(5421) <= a xor b;
    outputs(5422) <= not (a xor b);
    outputs(5423) <= a xor b;
    outputs(5424) <= not a;
    outputs(5425) <= not (a xor b);
    outputs(5426) <= not (a xor b);
    outputs(5427) <= not b;
    outputs(5428) <= a xor b;
    outputs(5429) <= b;
    outputs(5430) <= b;
    outputs(5431) <= b;
    outputs(5432) <= b and not a;
    outputs(5433) <= not b;
    outputs(5434) <= a and b;
    outputs(5435) <= a xor b;
    outputs(5436) <= a xor b;
    outputs(5437) <= not b;
    outputs(5438) <= not (a or b);
    outputs(5439) <= not (a and b);
    outputs(5440) <= not (a xor b);
    outputs(5441) <= a xor b;
    outputs(5442) <= not (a xor b);
    outputs(5443) <= not a;
    outputs(5444) <= not (a xor b);
    outputs(5445) <= a;
    outputs(5446) <= a and b;
    outputs(5447) <= not (a xor b);
    outputs(5448) <= not (a xor b);
    outputs(5449) <= a;
    outputs(5450) <= a;
    outputs(5451) <= not (a xor b);
    outputs(5452) <= a;
    outputs(5453) <= not b;
    outputs(5454) <= not a;
    outputs(5455) <= b;
    outputs(5456) <= not (a xor b);
    outputs(5457) <= not (a and b);
    outputs(5458) <= a and b;
    outputs(5459) <= not a or b;
    outputs(5460) <= a and not b;
    outputs(5461) <= b;
    outputs(5462) <= a xor b;
    outputs(5463) <= a or b;
    outputs(5464) <= a;
    outputs(5465) <= not (a or b);
    outputs(5466) <= not (a xor b);
    outputs(5467) <= not (a xor b);
    outputs(5468) <= b;
    outputs(5469) <= b;
    outputs(5470) <= not a;
    outputs(5471) <= not (a and b);
    outputs(5472) <= a xor b;
    outputs(5473) <= a;
    outputs(5474) <= a xor b;
    outputs(5475) <= a xor b;
    outputs(5476) <= a and b;
    outputs(5477) <= b;
    outputs(5478) <= not (a xor b);
    outputs(5479) <= a and not b;
    outputs(5480) <= a xor b;
    outputs(5481) <= not (a xor b);
    outputs(5482) <= b;
    outputs(5483) <= a;
    outputs(5484) <= b and not a;
    outputs(5485) <= not (a xor b);
    outputs(5486) <= not (a xor b);
    outputs(5487) <= not b;
    outputs(5488) <= a;
    outputs(5489) <= a xor b;
    outputs(5490) <= b;
    outputs(5491) <= not a;
    outputs(5492) <= not b or a;
    outputs(5493) <= a;
    outputs(5494) <= not a or b;
    outputs(5495) <= not b or a;
    outputs(5496) <= a and b;
    outputs(5497) <= not (a xor b);
    outputs(5498) <= a;
    outputs(5499) <= a xor b;
    outputs(5500) <= b and not a;
    outputs(5501) <= not b or a;
    outputs(5502) <= not (a and b);
    outputs(5503) <= b;
    outputs(5504) <= a xor b;
    outputs(5505) <= not (a or b);
    outputs(5506) <= a xor b;
    outputs(5507) <= a;
    outputs(5508) <= not b;
    outputs(5509) <= not a or b;
    outputs(5510) <= not b;
    outputs(5511) <= not b;
    outputs(5512) <= not (a xor b);
    outputs(5513) <= not a;
    outputs(5514) <= a and not b;
    outputs(5515) <= b;
    outputs(5516) <= not (a or b);
    outputs(5517) <= a;
    outputs(5518) <= not a;
    outputs(5519) <= b;
    outputs(5520) <= not (a xor b);
    outputs(5521) <= b and not a;
    outputs(5522) <= a and b;
    outputs(5523) <= a or b;
    outputs(5524) <= not (a and b);
    outputs(5525) <= a xor b;
    outputs(5526) <= not (a or b);
    outputs(5527) <= not b;
    outputs(5528) <= not (a xor b);
    outputs(5529) <= b and not a;
    outputs(5530) <= b;
    outputs(5531) <= not b;
    outputs(5532) <= b;
    outputs(5533) <= a and b;
    outputs(5534) <= b;
    outputs(5535) <= not b;
    outputs(5536) <= a and b;
    outputs(5537) <= a xor b;
    outputs(5538) <= b and not a;
    outputs(5539) <= b;
    outputs(5540) <= not b;
    outputs(5541) <= a and not b;
    outputs(5542) <= not (a xor b);
    outputs(5543) <= a;
    outputs(5544) <= a xor b;
    outputs(5545) <= not a;
    outputs(5546) <= not a;
    outputs(5547) <= not (a and b);
    outputs(5548) <= a xor b;
    outputs(5549) <= a xor b;
    outputs(5550) <= b;
    outputs(5551) <= not a;
    outputs(5552) <= a;
    outputs(5553) <= not (a xor b);
    outputs(5554) <= not b;
    outputs(5555) <= a xor b;
    outputs(5556) <= not a;
    outputs(5557) <= not b;
    outputs(5558) <= b;
    outputs(5559) <= not b;
    outputs(5560) <= a xor b;
    outputs(5561) <= not a or b;
    outputs(5562) <= not (a and b);
    outputs(5563) <= not (a xor b);
    outputs(5564) <= not a;
    outputs(5565) <= a and not b;
    outputs(5566) <= a xor b;
    outputs(5567) <= b;
    outputs(5568) <= not (a or b);
    outputs(5569) <= not b;
    outputs(5570) <= not (a or b);
    outputs(5571) <= not a;
    outputs(5572) <= a;
    outputs(5573) <= not a;
    outputs(5574) <= not (a xor b);
    outputs(5575) <= a xor b;
    outputs(5576) <= a;
    outputs(5577) <= not (a xor b);
    outputs(5578) <= b;
    outputs(5579) <= not a;
    outputs(5580) <= not a;
    outputs(5581) <= not a;
    outputs(5582) <= not b;
    outputs(5583) <= not a;
    outputs(5584) <= not b;
    outputs(5585) <= not b or a;
    outputs(5586) <= a;
    outputs(5587) <= a and not b;
    outputs(5588) <= not b;
    outputs(5589) <= not a;
    outputs(5590) <= b;
    outputs(5591) <= a and b;
    outputs(5592) <= not (a xor b);
    outputs(5593) <= not b;
    outputs(5594) <= not (a xor b);
    outputs(5595) <= b;
    outputs(5596) <= b;
    outputs(5597) <= a xor b;
    outputs(5598) <= a xor b;
    outputs(5599) <= not (a xor b);
    outputs(5600) <= not b or a;
    outputs(5601) <= not b;
    outputs(5602) <= not a or b;
    outputs(5603) <= b and not a;
    outputs(5604) <= a xor b;
    outputs(5605) <= a xor b;
    outputs(5606) <= not a or b;
    outputs(5607) <= a and b;
    outputs(5608) <= a xor b;
    outputs(5609) <= a xor b;
    outputs(5610) <= not b or a;
    outputs(5611) <= not (a xor b);
    outputs(5612) <= b;
    outputs(5613) <= a and b;
    outputs(5614) <= b;
    outputs(5615) <= a xor b;
    outputs(5616) <= not b;
    outputs(5617) <= b;
    outputs(5618) <= a or b;
    outputs(5619) <= b;
    outputs(5620) <= not (a or b);
    outputs(5621) <= a xor b;
    outputs(5622) <= a xor b;
    outputs(5623) <= not a;
    outputs(5624) <= not a;
    outputs(5625) <= b;
    outputs(5626) <= b;
    outputs(5627) <= a xor b;
    outputs(5628) <= a xor b;
    outputs(5629) <= not (a xor b);
    outputs(5630) <= not a;
    outputs(5631) <= b and not a;
    outputs(5632) <= not b;
    outputs(5633) <= not (a or b);
    outputs(5634) <= a and not b;
    outputs(5635) <= a;
    outputs(5636) <= a and not b;
    outputs(5637) <= a and not b;
    outputs(5638) <= not (a xor b);
    outputs(5639) <= not a;
    outputs(5640) <= not b;
    outputs(5641) <= a;
    outputs(5642) <= not a;
    outputs(5643) <= not (a xor b);
    outputs(5644) <= b;
    outputs(5645) <= not a;
    outputs(5646) <= not b;
    outputs(5647) <= not a;
    outputs(5648) <= not (a xor b);
    outputs(5649) <= b;
    outputs(5650) <= not b;
    outputs(5651) <= not (a xor b);
    outputs(5652) <= a;
    outputs(5653) <= not (a xor b);
    outputs(5654) <= not (a or b);
    outputs(5655) <= not (a xor b);
    outputs(5656) <= not (a xor b);
    outputs(5657) <= not b;
    outputs(5658) <= a xor b;
    outputs(5659) <= not (a or b);
    outputs(5660) <= not b;
    outputs(5661) <= not b;
    outputs(5662) <= not (a xor b);
    outputs(5663) <= not (a or b);
    outputs(5664) <= a and not b;
    outputs(5665) <= a and not b;
    outputs(5666) <= b and not a;
    outputs(5667) <= b;
    outputs(5668) <= a xor b;
    outputs(5669) <= not b;
    outputs(5670) <= b;
    outputs(5671) <= b and not a;
    outputs(5672) <= a xor b;
    outputs(5673) <= not (a or b);
    outputs(5674) <= not a or b;
    outputs(5675) <= not a;
    outputs(5676) <= a xor b;
    outputs(5677) <= not b;
    outputs(5678) <= not (a or b);
    outputs(5679) <= not (a xor b);
    outputs(5680) <= a xor b;
    outputs(5681) <= not b;
    outputs(5682) <= a and not b;
    outputs(5683) <= a xor b;
    outputs(5684) <= not b;
    outputs(5685) <= not (a or b);
    outputs(5686) <= a xor b;
    outputs(5687) <= not b;
    outputs(5688) <= not b;
    outputs(5689) <= a;
    outputs(5690) <= a xor b;
    outputs(5691) <= not (a xor b);
    outputs(5692) <= a;
    outputs(5693) <= not a;
    outputs(5694) <= a xor b;
    outputs(5695) <= not (a and b);
    outputs(5696) <= not (a and b);
    outputs(5697) <= a and not b;
    outputs(5698) <= a;
    outputs(5699) <= b;
    outputs(5700) <= not b;
    outputs(5701) <= not (a or b);
    outputs(5702) <= not (a xor b);
    outputs(5703) <= not b;
    outputs(5704) <= a xor b;
    outputs(5705) <= not (a xor b);
    outputs(5706) <= b;
    outputs(5707) <= a or b;
    outputs(5708) <= a xor b;
    outputs(5709) <= a xor b;
    outputs(5710) <= not b;
    outputs(5711) <= not a;
    outputs(5712) <= b;
    outputs(5713) <= a xor b;
    outputs(5714) <= not a;
    outputs(5715) <= a xor b;
    outputs(5716) <= a;
    outputs(5717) <= not a or b;
    outputs(5718) <= b;
    outputs(5719) <= a and b;
    outputs(5720) <= a;
    outputs(5721) <= a xor b;
    outputs(5722) <= a;
    outputs(5723) <= a and b;
    outputs(5724) <= not (a xor b);
    outputs(5725) <= a or b;
    outputs(5726) <= not a;
    outputs(5727) <= not a;
    outputs(5728) <= not b;
    outputs(5729) <= not (a or b);
    outputs(5730) <= a xor b;
    outputs(5731) <= not (a xor b);
    outputs(5732) <= not (a and b);
    outputs(5733) <= not (a xor b);
    outputs(5734) <= b;
    outputs(5735) <= not (a and b);
    outputs(5736) <= a;
    outputs(5737) <= not a;
    outputs(5738) <= a and not b;
    outputs(5739) <= b;
    outputs(5740) <= not (a xor b);
    outputs(5741) <= a;
    outputs(5742) <= a and not b;
    outputs(5743) <= b and not a;
    outputs(5744) <= not (a xor b);
    outputs(5745) <= not (a xor b);
    outputs(5746) <= not b;
    outputs(5747) <= b;
    outputs(5748) <= a xor b;
    outputs(5749) <= not (a or b);
    outputs(5750) <= not b;
    outputs(5751) <= a or b;
    outputs(5752) <= a xor b;
    outputs(5753) <= a;
    outputs(5754) <= not (a and b);
    outputs(5755) <= not (a or b);
    outputs(5756) <= a xor b;
    outputs(5757) <= b;
    outputs(5758) <= not a;
    outputs(5759) <= a;
    outputs(5760) <= b;
    outputs(5761) <= not a;
    outputs(5762) <= not (a xor b);
    outputs(5763) <= b and not a;
    outputs(5764) <= not (a xor b);
    outputs(5765) <= not a;
    outputs(5766) <= not a;
    outputs(5767) <= not a or b;
    outputs(5768) <= a or b;
    outputs(5769) <= a xor b;
    outputs(5770) <= a xor b;
    outputs(5771) <= b and not a;
    outputs(5772) <= not (a xor b);
    outputs(5773) <= not (a xor b);
    outputs(5774) <= not b;
    outputs(5775) <= not b or a;
    outputs(5776) <= not a or b;
    outputs(5777) <= a or b;
    outputs(5778) <= not (a xor b);
    outputs(5779) <= not (a xor b);
    outputs(5780) <= a xor b;
    outputs(5781) <= a xor b;
    outputs(5782) <= a;
    outputs(5783) <= not (a or b);
    outputs(5784) <= not (a xor b);
    outputs(5785) <= a and b;
    outputs(5786) <= not b;
    outputs(5787) <= not (a xor b);
    outputs(5788) <= a and b;
    outputs(5789) <= a or b;
    outputs(5790) <= a xor b;
    outputs(5791) <= b and not a;
    outputs(5792) <= a and b;
    outputs(5793) <= a xor b;
    outputs(5794) <= not b;
    outputs(5795) <= not b;
    outputs(5796) <= a xor b;
    outputs(5797) <= not (a xor b);
    outputs(5798) <= not (a and b);
    outputs(5799) <= not (a xor b);
    outputs(5800) <= not b or a;
    outputs(5801) <= not (a xor b);
    outputs(5802) <= not (a xor b);
    outputs(5803) <= b;
    outputs(5804) <= not (a xor b);
    outputs(5805) <= not b;
    outputs(5806) <= not a;
    outputs(5807) <= not b or a;
    outputs(5808) <= not (a and b);
    outputs(5809) <= a;
    outputs(5810) <= a or b;
    outputs(5811) <= b;
    outputs(5812) <= a and not b;
    outputs(5813) <= b;
    outputs(5814) <= a and b;
    outputs(5815) <= not (a or b);
    outputs(5816) <= not b or a;
    outputs(5817) <= b;
    outputs(5818) <= a xor b;
    outputs(5819) <= not (a or b);
    outputs(5820) <= a xor b;
    outputs(5821) <= not (a xor b);
    outputs(5822) <= a and not b;
    outputs(5823) <= not a;
    outputs(5824) <= not a;
    outputs(5825) <= b;
    outputs(5826) <= not (a or b);
    outputs(5827) <= not b;
    outputs(5828) <= a and not b;
    outputs(5829) <= not (a xor b);
    outputs(5830) <= not a or b;
    outputs(5831) <= not b;
    outputs(5832) <= not b;
    outputs(5833) <= a xor b;
    outputs(5834) <= a xor b;
    outputs(5835) <= a and not b;
    outputs(5836) <= not a or b;
    outputs(5837) <= not b or a;
    outputs(5838) <= not b;
    outputs(5839) <= not (a xor b);
    outputs(5840) <= a and b;
    outputs(5841) <= b;
    outputs(5842) <= a xor b;
    outputs(5843) <= a;
    outputs(5844) <= not b or a;
    outputs(5845) <= a xor b;
    outputs(5846) <= not (a and b);
    outputs(5847) <= b;
    outputs(5848) <= not b;
    outputs(5849) <= a and not b;
    outputs(5850) <= a xor b;
    outputs(5851) <= a;
    outputs(5852) <= a and not b;
    outputs(5853) <= a xor b;
    outputs(5854) <= not (a xor b);
    outputs(5855) <= a xor b;
    outputs(5856) <= not (a and b);
    outputs(5857) <= b;
    outputs(5858) <= a and not b;
    outputs(5859) <= not b;
    outputs(5860) <= not a;
    outputs(5861) <= a xor b;
    outputs(5862) <= a;
    outputs(5863) <= not b;
    outputs(5864) <= not (a or b);
    outputs(5865) <= not b;
    outputs(5866) <= b and not a;
    outputs(5867) <= not a;
    outputs(5868) <= not b;
    outputs(5869) <= a xor b;
    outputs(5870) <= a xor b;
    outputs(5871) <= a xor b;
    outputs(5872) <= b;
    outputs(5873) <= not (a or b);
    outputs(5874) <= b;
    outputs(5875) <= not a;
    outputs(5876) <= b;
    outputs(5877) <= a;
    outputs(5878) <= not a;
    outputs(5879) <= not a;
    outputs(5880) <= a;
    outputs(5881) <= not b;
    outputs(5882) <= not a or b;
    outputs(5883) <= not a or b;
    outputs(5884) <= not a;
    outputs(5885) <= a and b;
    outputs(5886) <= not (a or b);
    outputs(5887) <= a;
    outputs(5888) <= b;
    outputs(5889) <= not a;
    outputs(5890) <= b;
    outputs(5891) <= a xor b;
    outputs(5892) <= not b;
    outputs(5893) <= a xor b;
    outputs(5894) <= not a;
    outputs(5895) <= a;
    outputs(5896) <= a;
    outputs(5897) <= a or b;
    outputs(5898) <= a and b;
    outputs(5899) <= a and b;
    outputs(5900) <= not a;
    outputs(5901) <= a and not b;
    outputs(5902) <= a xor b;
    outputs(5903) <= not b;
    outputs(5904) <= not (a xor b);
    outputs(5905) <= a;
    outputs(5906) <= not (a xor b);
    outputs(5907) <= not (a xor b);
    outputs(5908) <= not (a xor b);
    outputs(5909) <= not (a xor b);
    outputs(5910) <= not (a or b);
    outputs(5911) <= b and not a;
    outputs(5912) <= b;
    outputs(5913) <= not b;
    outputs(5914) <= b and not a;
    outputs(5915) <= not (a xor b);
    outputs(5916) <= not a;
    outputs(5917) <= a xor b;
    outputs(5918) <= not a;
    outputs(5919) <= a;
    outputs(5920) <= not (a xor b);
    outputs(5921) <= a;
    outputs(5922) <= not (a xor b);
    outputs(5923) <= a xor b;
    outputs(5924) <= a;
    outputs(5925) <= not a;
    outputs(5926) <= not a;
    outputs(5927) <= not a;
    outputs(5928) <= a xor b;
    outputs(5929) <= not (a xor b);
    outputs(5930) <= a xor b;
    outputs(5931) <= not b;
    outputs(5932) <= not (a and b);
    outputs(5933) <= not (a xor b);
    outputs(5934) <= not (a xor b);
    outputs(5935) <= not (a xor b);
    outputs(5936) <= a xor b;
    outputs(5937) <= a;
    outputs(5938) <= not b or a;
    outputs(5939) <= a;
    outputs(5940) <= a;
    outputs(5941) <= a xor b;
    outputs(5942) <= a xor b;
    outputs(5943) <= a xor b;
    outputs(5944) <= not b;
    outputs(5945) <= not a or b;
    outputs(5946) <= a xor b;
    outputs(5947) <= not (a xor b);
    outputs(5948) <= not a;
    outputs(5949) <= b;
    outputs(5950) <= a or b;
    outputs(5951) <= a and b;
    outputs(5952) <= a xor b;
    outputs(5953) <= not a;
    outputs(5954) <= not (a xor b);
    outputs(5955) <= b;
    outputs(5956) <= b;
    outputs(5957) <= b;
    outputs(5958) <= not (a and b);
    outputs(5959) <= a or b;
    outputs(5960) <= a xor b;
    outputs(5961) <= not b;
    outputs(5962) <= a xor b;
    outputs(5963) <= a;
    outputs(5964) <= not (a xor b);
    outputs(5965) <= not (a xor b);
    outputs(5966) <= b;
    outputs(5967) <= a or b;
    outputs(5968) <= not b;
    outputs(5969) <= not (a xor b);
    outputs(5970) <= b;
    outputs(5971) <= a;
    outputs(5972) <= not a;
    outputs(5973) <= a;
    outputs(5974) <= not (a xor b);
    outputs(5975) <= not b;
    outputs(5976) <= not (a xor b);
    outputs(5977) <= not b or a;
    outputs(5978) <= a;
    outputs(5979) <= not a;
    outputs(5980) <= a xor b;
    outputs(5981) <= a xor b;
    outputs(5982) <= a;
    outputs(5983) <= a or b;
    outputs(5984) <= not a;
    outputs(5985) <= not (a xor b);
    outputs(5986) <= a xor b;
    outputs(5987) <= a xor b;
    outputs(5988) <= a xor b;
    outputs(5989) <= not (a or b);
    outputs(5990) <= a;
    outputs(5991) <= b;
    outputs(5992) <= b and not a;
    outputs(5993) <= a xor b;
    outputs(5994) <= not a or b;
    outputs(5995) <= a;
    outputs(5996) <= b;
    outputs(5997) <= a and b;
    outputs(5998) <= b;
    outputs(5999) <= a and not b;
    outputs(6000) <= a xor b;
    outputs(6001) <= not (a xor b);
    outputs(6002) <= not (a xor b);
    outputs(6003) <= a or b;
    outputs(6004) <= a;
    outputs(6005) <= a xor b;
    outputs(6006) <= not (a xor b);
    outputs(6007) <= not b;
    outputs(6008) <= not (a or b);
    outputs(6009) <= not (a and b);
    outputs(6010) <= not a;
    outputs(6011) <= not (a xor b);
    outputs(6012) <= b and not a;
    outputs(6013) <= not b;
    outputs(6014) <= not (a xor b);
    outputs(6015) <= a;
    outputs(6016) <= not (a or b);
    outputs(6017) <= not (a xor b);
    outputs(6018) <= not a;
    outputs(6019) <= a;
    outputs(6020) <= a xor b;
    outputs(6021) <= not a;
    outputs(6022) <= not b or a;
    outputs(6023) <= not (a xor b);
    outputs(6024) <= not b or a;
    outputs(6025) <= not a;
    outputs(6026) <= not a;
    outputs(6027) <= a xor b;
    outputs(6028) <= b;
    outputs(6029) <= b;
    outputs(6030) <= a or b;
    outputs(6031) <= not (a xor b);
    outputs(6032) <= a xor b;
    outputs(6033) <= not (a xor b);
    outputs(6034) <= not (a or b);
    outputs(6035) <= not b;
    outputs(6036) <= a and not b;
    outputs(6037) <= a xor b;
    outputs(6038) <= not a;
    outputs(6039) <= a or b;
    outputs(6040) <= a xor b;
    outputs(6041) <= a xor b;
    outputs(6042) <= not (a xor b);
    outputs(6043) <= not a;
    outputs(6044) <= a;
    outputs(6045) <= b and not a;
    outputs(6046) <= not b;
    outputs(6047) <= a xor b;
    outputs(6048) <= not (a xor b);
    outputs(6049) <= not b;
    outputs(6050) <= b;
    outputs(6051) <= a and b;
    outputs(6052) <= not (a or b);
    outputs(6053) <= not a;
    outputs(6054) <= not b or a;
    outputs(6055) <= a;
    outputs(6056) <= not (a xor b);
    outputs(6057) <= b;
    outputs(6058) <= a and not b;
    outputs(6059) <= a or b;
    outputs(6060) <= not (a or b);
    outputs(6061) <= not a;
    outputs(6062) <= a xor b;
    outputs(6063) <= a and not b;
    outputs(6064) <= a or b;
    outputs(6065) <= not a;
    outputs(6066) <= a and not b;
    outputs(6067) <= not (a or b);
    outputs(6068) <= not a;
    outputs(6069) <= a xor b;
    outputs(6070) <= a xor b;
    outputs(6071) <= not a;
    outputs(6072) <= not a;
    outputs(6073) <= not b;
    outputs(6074) <= not (a or b);
    outputs(6075) <= not a or b;
    outputs(6076) <= a xor b;
    outputs(6077) <= b;
    outputs(6078) <= b;
    outputs(6079) <= a;
    outputs(6080) <= not b;
    outputs(6081) <= not b;
    outputs(6082) <= not a;
    outputs(6083) <= not a;
    outputs(6084) <= not a;
    outputs(6085) <= a and not b;
    outputs(6086) <= not b;
    outputs(6087) <= a and b;
    outputs(6088) <= a;
    outputs(6089) <= a xor b;
    outputs(6090) <= a or b;
    outputs(6091) <= not (a xor b);
    outputs(6092) <= not b or a;
    outputs(6093) <= a;
    outputs(6094) <= a or b;
    outputs(6095) <= b;
    outputs(6096) <= a xor b;
    outputs(6097) <= not a;
    outputs(6098) <= not (a xor b);
    outputs(6099) <= not a;
    outputs(6100) <= not (a xor b);
    outputs(6101) <= a xor b;
    outputs(6102) <= a xor b;
    outputs(6103) <= a;
    outputs(6104) <= a;
    outputs(6105) <= not (a or b);
    outputs(6106) <= b;
    outputs(6107) <= not (a xor b);
    outputs(6108) <= not (a or b);
    outputs(6109) <= not (a xor b);
    outputs(6110) <= not b;
    outputs(6111) <= a xor b;
    outputs(6112) <= not (a xor b);
    outputs(6113) <= a;
    outputs(6114) <= a;
    outputs(6115) <= a;
    outputs(6116) <= not (a xor b);
    outputs(6117) <= a;
    outputs(6118) <= not a;
    outputs(6119) <= not a or b;
    outputs(6120) <= not (a xor b);
    outputs(6121) <= not (a xor b);
    outputs(6122) <= not a or b;
    outputs(6123) <= not (a xor b);
    outputs(6124) <= a xor b;
    outputs(6125) <= a xor b;
    outputs(6126) <= not (a xor b);
    outputs(6127) <= not b;
    outputs(6128) <= not (a xor b);
    outputs(6129) <= b;
    outputs(6130) <= not (a or b);
    outputs(6131) <= not a;
    outputs(6132) <= b;
    outputs(6133) <= a xor b;
    outputs(6134) <= not (a xor b);
    outputs(6135) <= a;
    outputs(6136) <= not b;
    outputs(6137) <= not (a xor b);
    outputs(6138) <= a or b;
    outputs(6139) <= a;
    outputs(6140) <= not a;
    outputs(6141) <= a xor b;
    outputs(6142) <= a;
    outputs(6143) <= not (a or b);
    outputs(6144) <= a or b;
    outputs(6145) <= a xor b;
    outputs(6146) <= a;
    outputs(6147) <= b;
    outputs(6148) <= not b;
    outputs(6149) <= a xor b;
    outputs(6150) <= a;
    outputs(6151) <= a;
    outputs(6152) <= a;
    outputs(6153) <= b and not a;
    outputs(6154) <= not b;
    outputs(6155) <= not b;
    outputs(6156) <= b;
    outputs(6157) <= not (a or b);
    outputs(6158) <= b and not a;
    outputs(6159) <= not (a or b);
    outputs(6160) <= not (a xor b);
    outputs(6161) <= not (a or b);
    outputs(6162) <= not a;
    outputs(6163) <= b;
    outputs(6164) <= not a;
    outputs(6165) <= not (a xor b);
    outputs(6166) <= a and b;
    outputs(6167) <= a or b;
    outputs(6168) <= a xor b;
    outputs(6169) <= a xor b;
    outputs(6170) <= not (a and b);
    outputs(6171) <= not (a xor b);
    outputs(6172) <= not a or b;
    outputs(6173) <= not (a xor b);
    outputs(6174) <= not a;
    outputs(6175) <= a and b;
    outputs(6176) <= not b;
    outputs(6177) <= not a;
    outputs(6178) <= a;
    outputs(6179) <= a xor b;
    outputs(6180) <= a and b;
    outputs(6181) <= a xor b;
    outputs(6182) <= not (a and b);
    outputs(6183) <= not a;
    outputs(6184) <= b;
    outputs(6185) <= not b;
    outputs(6186) <= not b or a;
    outputs(6187) <= a and b;
    outputs(6188) <= a and not b;
    outputs(6189) <= b;
    outputs(6190) <= not a;
    outputs(6191) <= a and b;
    outputs(6192) <= a;
    outputs(6193) <= a;
    outputs(6194) <= not b;
    outputs(6195) <= not a;
    outputs(6196) <= not (a xor b);
    outputs(6197) <= not b;
    outputs(6198) <= not a;
    outputs(6199) <= not (a or b);
    outputs(6200) <= a xor b;
    outputs(6201) <= a xor b;
    outputs(6202) <= a xor b;
    outputs(6203) <= not (a xor b);
    outputs(6204) <= not a or b;
    outputs(6205) <= not a;
    outputs(6206) <= a;
    outputs(6207) <= not (a or b);
    outputs(6208) <= a;
    outputs(6209) <= a and b;
    outputs(6210) <= a xor b;
    outputs(6211) <= not a;
    outputs(6212) <= not b or a;
    outputs(6213) <= a xor b;
    outputs(6214) <= not a;
    outputs(6215) <= a xor b;
    outputs(6216) <= not (a xor b);
    outputs(6217) <= a;
    outputs(6218) <= a and b;
    outputs(6219) <= b;
    outputs(6220) <= not b;
    outputs(6221) <= b and not a;
    outputs(6222) <= not (a or b);
    outputs(6223) <= not a;
    outputs(6224) <= not (a or b);
    outputs(6225) <= not b;
    outputs(6226) <= b and not a;
    outputs(6227) <= b;
    outputs(6228) <= not a or b;
    outputs(6229) <= a;
    outputs(6230) <= not a;
    outputs(6231) <= a xor b;
    outputs(6232) <= not b or a;
    outputs(6233) <= a xor b;
    outputs(6234) <= a or b;
    outputs(6235) <= not a or b;
    outputs(6236) <= not a;
    outputs(6237) <= not b;
    outputs(6238) <= not a or b;
    outputs(6239) <= a xor b;
    outputs(6240) <= not (a or b);
    outputs(6241) <= not a;
    outputs(6242) <= not a or b;
    outputs(6243) <= not (a xor b);
    outputs(6244) <= a xor b;
    outputs(6245) <= a xor b;
    outputs(6246) <= not (a or b);
    outputs(6247) <= b;
    outputs(6248) <= not (a xor b);
    outputs(6249) <= not b;
    outputs(6250) <= not (a xor b);
    outputs(6251) <= a;
    outputs(6252) <= not b;
    outputs(6253) <= not (a xor b);
    outputs(6254) <= not b;
    outputs(6255) <= not b;
    outputs(6256) <= b;
    outputs(6257) <= a xor b;
    outputs(6258) <= a;
    outputs(6259) <= a;
    outputs(6260) <= a or b;
    outputs(6261) <= not a;
    outputs(6262) <= not (a xor b);
    outputs(6263) <= not (a xor b);
    outputs(6264) <= b;
    outputs(6265) <= a xor b;
    outputs(6266) <= a xor b;
    outputs(6267) <= not a;
    outputs(6268) <= not a;
    outputs(6269) <= not (a xor b);
    outputs(6270) <= a;
    outputs(6271) <= not b;
    outputs(6272) <= not (a xor b);
    outputs(6273) <= a and b;
    outputs(6274) <= not b;
    outputs(6275) <= b;
    outputs(6276) <= not b;
    outputs(6277) <= b and not a;
    outputs(6278) <= a xor b;
    outputs(6279) <= b;
    outputs(6280) <= a and b;
    outputs(6281) <= a and b;
    outputs(6282) <= not (a xor b);
    outputs(6283) <= b;
    outputs(6284) <= not (a xor b);
    outputs(6285) <= a;
    outputs(6286) <= a xor b;
    outputs(6287) <= a;
    outputs(6288) <= not a;
    outputs(6289) <= a xor b;
    outputs(6290) <= a xor b;
    outputs(6291) <= not b;
    outputs(6292) <= not (a xor b);
    outputs(6293) <= b and not a;
    outputs(6294) <= a xor b;
    outputs(6295) <= a and not b;
    outputs(6296) <= not b or a;
    outputs(6297) <= not a;
    outputs(6298) <= a or b;
    outputs(6299) <= not b;
    outputs(6300) <= a;
    outputs(6301) <= a and not b;
    outputs(6302) <= not (a xor b);
    outputs(6303) <= a;
    outputs(6304) <= b and not a;
    outputs(6305) <= b and not a;
    outputs(6306) <= not a;
    outputs(6307) <= a;
    outputs(6308) <= not b;
    outputs(6309) <= a and b;
    outputs(6310) <= not a;
    outputs(6311) <= not a or b;
    outputs(6312) <= a xor b;
    outputs(6313) <= a xor b;
    outputs(6314) <= a;
    outputs(6315) <= not b;
    outputs(6316) <= not b or a;
    outputs(6317) <= a xor b;
    outputs(6318) <= a and b;
    outputs(6319) <= b and not a;
    outputs(6320) <= not (a xor b);
    outputs(6321) <= not (a xor b);
    outputs(6322) <= a;
    outputs(6323) <= not (a xor b);
    outputs(6324) <= b;
    outputs(6325) <= not (a or b);
    outputs(6326) <= not (a xor b);
    outputs(6327) <= a xor b;
    outputs(6328) <= not b;
    outputs(6329) <= not (a xor b);
    outputs(6330) <= not b;
    outputs(6331) <= not (a xor b);
    outputs(6332) <= a and b;
    outputs(6333) <= not a or b;
    outputs(6334) <= not (a and b);
    outputs(6335) <= not a;
    outputs(6336) <= not a;
    outputs(6337) <= a xor b;
    outputs(6338) <= a and b;
    outputs(6339) <= not (a or b);
    outputs(6340) <= a xor b;
    outputs(6341) <= a and not b;
    outputs(6342) <= b;
    outputs(6343) <= not (a xor b);
    outputs(6344) <= not b;
    outputs(6345) <= not a;
    outputs(6346) <= a;
    outputs(6347) <= not a;
    outputs(6348) <= a and not b;
    outputs(6349) <= not a;
    outputs(6350) <= b;
    outputs(6351) <= not a;
    outputs(6352) <= not (a xor b);
    outputs(6353) <= a xor b;
    outputs(6354) <= not (a xor b);
    outputs(6355) <= a and not b;
    outputs(6356) <= a xor b;
    outputs(6357) <= b;
    outputs(6358) <= not b;
    outputs(6359) <= a;
    outputs(6360) <= b;
    outputs(6361) <= b and not a;
    outputs(6362) <= b;
    outputs(6363) <= not a or b;
    outputs(6364) <= a and b;
    outputs(6365) <= not a;
    outputs(6366) <= not b;
    outputs(6367) <= not (a and b);
    outputs(6368) <= not a or b;
    outputs(6369) <= not a;
    outputs(6370) <= a and b;
    outputs(6371) <= a;
    outputs(6372) <= not a;
    outputs(6373) <= not a;
    outputs(6374) <= not a;
    outputs(6375) <= not (a xor b);
    outputs(6376) <= not (a or b);
    outputs(6377) <= a;
    outputs(6378) <= a or b;
    outputs(6379) <= not b;
    outputs(6380) <= a xor b;
    outputs(6381) <= a or b;
    outputs(6382) <= not a;
    outputs(6383) <= b;
    outputs(6384) <= not (a xor b);
    outputs(6385) <= not b;
    outputs(6386) <= a xor b;
    outputs(6387) <= not (a xor b);
    outputs(6388) <= a xor b;
    outputs(6389) <= not (a xor b);
    outputs(6390) <= a;
    outputs(6391) <= not (a xor b);
    outputs(6392) <= a xor b;
    outputs(6393) <= a and not b;
    outputs(6394) <= b;
    outputs(6395) <= a;
    outputs(6396) <= b and not a;
    outputs(6397) <= not b;
    outputs(6398) <= a;
    outputs(6399) <= not (a xor b);
    outputs(6400) <= not b;
    outputs(6401) <= not (a xor b);
    outputs(6402) <= not (a xor b);
    outputs(6403) <= not (a xor b);
    outputs(6404) <= a and b;
    outputs(6405) <= not (a or b);
    outputs(6406) <= not a;
    outputs(6407) <= not (a and b);
    outputs(6408) <= a and b;
    outputs(6409) <= a xor b;
    outputs(6410) <= a xor b;
    outputs(6411) <= a and b;
    outputs(6412) <= not (a xor b);
    outputs(6413) <= a and not b;
    outputs(6414) <= a;
    outputs(6415) <= b and not a;
    outputs(6416) <= b and not a;
    outputs(6417) <= not b;
    outputs(6418) <= not (a xor b);
    outputs(6419) <= not a or b;
    outputs(6420) <= a xor b;
    outputs(6421) <= not a;
    outputs(6422) <= not (a or b);
    outputs(6423) <= not a;
    outputs(6424) <= not b;
    outputs(6425) <= not a or b;
    outputs(6426) <= b;
    outputs(6427) <= a;
    outputs(6428) <= b;
    outputs(6429) <= not a;
    outputs(6430) <= not (a or b);
    outputs(6431) <= not b;
    outputs(6432) <= not a;
    outputs(6433) <= a xor b;
    outputs(6434) <= a;
    outputs(6435) <= not b or a;
    outputs(6436) <= not (a xor b);
    outputs(6437) <= not (a or b);
    outputs(6438) <= a xor b;
    outputs(6439) <= a xor b;
    outputs(6440) <= not (a or b);
    outputs(6441) <= not (a xor b);
    outputs(6442) <= not b;
    outputs(6443) <= not b;
    outputs(6444) <= not b;
    outputs(6445) <= a xor b;
    outputs(6446) <= not a;
    outputs(6447) <= a xor b;
    outputs(6448) <= not a or b;
    outputs(6449) <= not (a or b);
    outputs(6450) <= b;
    outputs(6451) <= not a;
    outputs(6452) <= not b;
    outputs(6453) <= not b;
    outputs(6454) <= not (a xor b);
    outputs(6455) <= not (a xor b);
    outputs(6456) <= b;
    outputs(6457) <= a and not b;
    outputs(6458) <= not a;
    outputs(6459) <= not (a xor b);
    outputs(6460) <= not a;
    outputs(6461) <= a xor b;
    outputs(6462) <= not b;
    outputs(6463) <= a and not b;
    outputs(6464) <= b;
    outputs(6465) <= a xor b;
    outputs(6466) <= not b;
    outputs(6467) <= not a or b;
    outputs(6468) <= not a or b;
    outputs(6469) <= a;
    outputs(6470) <= not a;
    outputs(6471) <= not (a and b);
    outputs(6472) <= b;
    outputs(6473) <= not a or b;
    outputs(6474) <= a and not b;
    outputs(6475) <= b;
    outputs(6476) <= b;
    outputs(6477) <= a and b;
    outputs(6478) <= not (a or b);
    outputs(6479) <= a or b;
    outputs(6480) <= a and not b;
    outputs(6481) <= not b;
    outputs(6482) <= not a;
    outputs(6483) <= a and b;
    outputs(6484) <= not b;
    outputs(6485) <= not (a xor b);
    outputs(6486) <= not (a xor b);
    outputs(6487) <= a xor b;
    outputs(6488) <= a and b;
    outputs(6489) <= not (a xor b);
    outputs(6490) <= not (a xor b);
    outputs(6491) <= not b;
    outputs(6492) <= not b;
    outputs(6493) <= not (a or b);
    outputs(6494) <= not (a or b);
    outputs(6495) <= a xor b;
    outputs(6496) <= a;
    outputs(6497) <= b and not a;
    outputs(6498) <= a;
    outputs(6499) <= a xor b;
    outputs(6500) <= not (a or b);
    outputs(6501) <= not (a xor b);
    outputs(6502) <= a xor b;
    outputs(6503) <= not b;
    outputs(6504) <= a;
    outputs(6505) <= not b;
    outputs(6506) <= a;
    outputs(6507) <= not (a or b);
    outputs(6508) <= a;
    outputs(6509) <= not b;
    outputs(6510) <= a xor b;
    outputs(6511) <= not b;
    outputs(6512) <= not b or a;
    outputs(6513) <= a xor b;
    outputs(6514) <= not (a xor b);
    outputs(6515) <= a xor b;
    outputs(6516) <= not (a and b);
    outputs(6517) <= b;
    outputs(6518) <= b;
    outputs(6519) <= b;
    outputs(6520) <= not b;
    outputs(6521) <= a;
    outputs(6522) <= a and not b;
    outputs(6523) <= a;
    outputs(6524) <= not a;
    outputs(6525) <= not (a xor b);
    outputs(6526) <= b and not a;
    outputs(6527) <= not (a xor b);
    outputs(6528) <= not b;
    outputs(6529) <= b and not a;
    outputs(6530) <= a and not b;
    outputs(6531) <= not (a xor b);
    outputs(6532) <= not b;
    outputs(6533) <= not b or a;
    outputs(6534) <= a;
    outputs(6535) <= a xor b;
    outputs(6536) <= b and not a;
    outputs(6537) <= a;
    outputs(6538) <= a;
    outputs(6539) <= a and b;
    outputs(6540) <= a;
    outputs(6541) <= b;
    outputs(6542) <= not b;
    outputs(6543) <= not a;
    outputs(6544) <= not a;
    outputs(6545) <= not a;
    outputs(6546) <= not a;
    outputs(6547) <= a and b;
    outputs(6548) <= not (a xor b);
    outputs(6549) <= a xor b;
    outputs(6550) <= not a;
    outputs(6551) <= a;
    outputs(6552) <= a;
    outputs(6553) <= not a;
    outputs(6554) <= not b or a;
    outputs(6555) <= b;
    outputs(6556) <= a;
    outputs(6557) <= not a;
    outputs(6558) <= a xor b;
    outputs(6559) <= not (a xor b);
    outputs(6560) <= a;
    outputs(6561) <= a and not b;
    outputs(6562) <= not (a xor b);
    outputs(6563) <= not a or b;
    outputs(6564) <= b and not a;
    outputs(6565) <= not (a and b);
    outputs(6566) <= a;
    outputs(6567) <= not (a xor b);
    outputs(6568) <= a xor b;
    outputs(6569) <= b;
    outputs(6570) <= a;
    outputs(6571) <= a and b;
    outputs(6572) <= a and b;
    outputs(6573) <= a xor b;
    outputs(6574) <= not (a xor b);
    outputs(6575) <= a xor b;
    outputs(6576) <= not a;
    outputs(6577) <= not b;
    outputs(6578) <= a;
    outputs(6579) <= not b or a;
    outputs(6580) <= not a;
    outputs(6581) <= a;
    outputs(6582) <= not (a xor b);
    outputs(6583) <= not b;
    outputs(6584) <= not b;
    outputs(6585) <= not a;
    outputs(6586) <= not a;
    outputs(6587) <= not a;
    outputs(6588) <= not (a xor b);
    outputs(6589) <= not a;
    outputs(6590) <= a and not b;
    outputs(6591) <= not b or a;
    outputs(6592) <= a and b;
    outputs(6593) <= a xor b;
    outputs(6594) <= not b;
    outputs(6595) <= b;
    outputs(6596) <= a and not b;
    outputs(6597) <= not (a or b);
    outputs(6598) <= b and not a;
    outputs(6599) <= not a;
    outputs(6600) <= not (a xor b);
    outputs(6601) <= not b;
    outputs(6602) <= not (a or b);
    outputs(6603) <= a;
    outputs(6604) <= a xor b;
    outputs(6605) <= not a;
    outputs(6606) <= b and not a;
    outputs(6607) <= a or b;
    outputs(6608) <= not (a xor b);
    outputs(6609) <= a xor b;
    outputs(6610) <= not (a xor b);
    outputs(6611) <= not (a xor b);
    outputs(6612) <= a;
    outputs(6613) <= b and not a;
    outputs(6614) <= a xor b;
    outputs(6615) <= not (a xor b);
    outputs(6616) <= not a;
    outputs(6617) <= a;
    outputs(6618) <= b and not a;
    outputs(6619) <= b;
    outputs(6620) <= a;
    outputs(6621) <= b and not a;
    outputs(6622) <= a xor b;
    outputs(6623) <= a or b;
    outputs(6624) <= a;
    outputs(6625) <= b;
    outputs(6626) <= a;
    outputs(6627) <= not (a or b);
    outputs(6628) <= not b;
    outputs(6629) <= not (a xor b);
    outputs(6630) <= not a;
    outputs(6631) <= not b;
    outputs(6632) <= a;
    outputs(6633) <= b and not a;
    outputs(6634) <= a and not b;
    outputs(6635) <= a and b;
    outputs(6636) <= a xor b;
    outputs(6637) <= not (a xor b);
    outputs(6638) <= a and b;
    outputs(6639) <= not a;
    outputs(6640) <= not (a xor b);
    outputs(6641) <= not b;
    outputs(6642) <= not (a or b);
    outputs(6643) <= not a;
    outputs(6644) <= not (a xor b);
    outputs(6645) <= b;
    outputs(6646) <= a and not b;
    outputs(6647) <= not a or b;
    outputs(6648) <= not b;
    outputs(6649) <= a xor b;
    outputs(6650) <= a xor b;
    outputs(6651) <= not b or a;
    outputs(6652) <= a xor b;
    outputs(6653) <= not b;
    outputs(6654) <= a and b;
    outputs(6655) <= not a;
    outputs(6656) <= not a;
    outputs(6657) <= a;
    outputs(6658) <= a xor b;
    outputs(6659) <= b and not a;
    outputs(6660) <= not a or b;
    outputs(6661) <= not (a xor b);
    outputs(6662) <= not a;
    outputs(6663) <= a;
    outputs(6664) <= not (a or b);
    outputs(6665) <= not a;
    outputs(6666) <= not a;
    outputs(6667) <= b and not a;
    outputs(6668) <= a or b;
    outputs(6669) <= a xor b;
    outputs(6670) <= not b;
    outputs(6671) <= not (a xor b);
    outputs(6672) <= not b;
    outputs(6673) <= a and not b;
    outputs(6674) <= a and b;
    outputs(6675) <= a and b;
    outputs(6676) <= not (a xor b);
    outputs(6677) <= b;
    outputs(6678) <= a xor b;
    outputs(6679) <= not (a xor b);
    outputs(6680) <= not (a xor b);
    outputs(6681) <= not (a xor b);
    outputs(6682) <= not b;
    outputs(6683) <= not a;
    outputs(6684) <= not (a xor b);
    outputs(6685) <= not a;
    outputs(6686) <= a;
    outputs(6687) <= b and not a;
    outputs(6688) <= a and not b;
    outputs(6689) <= b;
    outputs(6690) <= not b;
    outputs(6691) <= b;
    outputs(6692) <= not a;
    outputs(6693) <= not b;
    outputs(6694) <= a;
    outputs(6695) <= a xor b;
    outputs(6696) <= not (a and b);
    outputs(6697) <= a;
    outputs(6698) <= a;
    outputs(6699) <= not (a xor b);
    outputs(6700) <= not b;
    outputs(6701) <= a;
    outputs(6702) <= b;
    outputs(6703) <= a xor b;
    outputs(6704) <= not (a xor b);
    outputs(6705) <= not (a xor b);
    outputs(6706) <= not (a xor b);
    outputs(6707) <= not (a xor b);
    outputs(6708) <= b;
    outputs(6709) <= a xor b;
    outputs(6710) <= a xor b;
    outputs(6711) <= a;
    outputs(6712) <= not b;
    outputs(6713) <= a;
    outputs(6714) <= not a;
    outputs(6715) <= a and not b;
    outputs(6716) <= not (a xor b);
    outputs(6717) <= not b or a;
    outputs(6718) <= not a or b;
    outputs(6719) <= b;
    outputs(6720) <= a xor b;
    outputs(6721) <= not b or a;
    outputs(6722) <= not a;
    outputs(6723) <= b and not a;
    outputs(6724) <= a and b;
    outputs(6725) <= b and not a;
    outputs(6726) <= not b;
    outputs(6727) <= not a;
    outputs(6728) <= not (a xor b);
    outputs(6729) <= a and b;
    outputs(6730) <= b;
    outputs(6731) <= a;
    outputs(6732) <= not a or b;
    outputs(6733) <= b and not a;
    outputs(6734) <= not a;
    outputs(6735) <= not (a or b);
    outputs(6736) <= a xor b;
    outputs(6737) <= not (a xor b);
    outputs(6738) <= not b;
    outputs(6739) <= a or b;
    outputs(6740) <= a or b;
    outputs(6741) <= b;
    outputs(6742) <= b;
    outputs(6743) <= not (a or b);
    outputs(6744) <= b and not a;
    outputs(6745) <= not a;
    outputs(6746) <= a xor b;
    outputs(6747) <= b and not a;
    outputs(6748) <= a and not b;
    outputs(6749) <= b;
    outputs(6750) <= not a or b;
    outputs(6751) <= a;
    outputs(6752) <= a xor b;
    outputs(6753) <= a or b;
    outputs(6754) <= not (a xor b);
    outputs(6755) <= a;
    outputs(6756) <= b;
    outputs(6757) <= b;
    outputs(6758) <= a;
    outputs(6759) <= b and not a;
    outputs(6760) <= a and b;
    outputs(6761) <= b and not a;
    outputs(6762) <= not b;
    outputs(6763) <= not b;
    outputs(6764) <= a or b;
    outputs(6765) <= a;
    outputs(6766) <= a and not b;
    outputs(6767) <= a and not b;
    outputs(6768) <= not a;
    outputs(6769) <= a xor b;
    outputs(6770) <= a;
    outputs(6771) <= not (a and b);
    outputs(6772) <= a;
    outputs(6773) <= a;
    outputs(6774) <= not a or b;
    outputs(6775) <= a and not b;
    outputs(6776) <= not b;
    outputs(6777) <= not (a and b);
    outputs(6778) <= not (a or b);
    outputs(6779) <= not (a xor b);
    outputs(6780) <= not (a xor b);
    outputs(6781) <= not b or a;
    outputs(6782) <= b and not a;
    outputs(6783) <= a;
    outputs(6784) <= not (a xor b);
    outputs(6785) <= a and not b;
    outputs(6786) <= a or b;
    outputs(6787) <= not (a and b);
    outputs(6788) <= not b or a;
    outputs(6789) <= not a;
    outputs(6790) <= b;
    outputs(6791) <= not (a or b);
    outputs(6792) <= a and not b;
    outputs(6793) <= a xor b;
    outputs(6794) <= a;
    outputs(6795) <= not a;
    outputs(6796) <= not b or a;
    outputs(6797) <= not a;
    outputs(6798) <= not b;
    outputs(6799) <= a and b;
    outputs(6800) <= not b;
    outputs(6801) <= a xor b;
    outputs(6802) <= a xor b;
    outputs(6803) <= a xor b;
    outputs(6804) <= a xor b;
    outputs(6805) <= b and not a;
    outputs(6806) <= a and not b;
    outputs(6807) <= a and not b;
    outputs(6808) <= a or b;
    outputs(6809) <= not (a xor b);
    outputs(6810) <= not (a xor b);
    outputs(6811) <= b;
    outputs(6812) <= not (a or b);
    outputs(6813) <= not b;
    outputs(6814) <= not (a or b);
    outputs(6815) <= not b;
    outputs(6816) <= a;
    outputs(6817) <= not a;
    outputs(6818) <= not (a xor b);
    outputs(6819) <= b and not a;
    outputs(6820) <= a xor b;
    outputs(6821) <= not a;
    outputs(6822) <= not b;
    outputs(6823) <= b;
    outputs(6824) <= not b;
    outputs(6825) <= not b;
    outputs(6826) <= a and not b;
    outputs(6827) <= b and not a;
    outputs(6828) <= a and b;
    outputs(6829) <= not a;
    outputs(6830) <= b;
    outputs(6831) <= not b;
    outputs(6832) <= a xor b;
    outputs(6833) <= not b;
    outputs(6834) <= b and not a;
    outputs(6835) <= a and b;
    outputs(6836) <= a xor b;
    outputs(6837) <= not a;
    outputs(6838) <= a;
    outputs(6839) <= a;
    outputs(6840) <= not b or a;
    outputs(6841) <= a and b;
    outputs(6842) <= b;
    outputs(6843) <= a xor b;
    outputs(6844) <= not b;
    outputs(6845) <= not (a and b);
    outputs(6846) <= not (a xor b);
    outputs(6847) <= not a;
    outputs(6848) <= not (a xor b);
    outputs(6849) <= not a or b;
    outputs(6850) <= a;
    outputs(6851) <= a xor b;
    outputs(6852) <= not b;
    outputs(6853) <= b;
    outputs(6854) <= b and not a;
    outputs(6855) <= b;
    outputs(6856) <= not a;
    outputs(6857) <= not a;
    outputs(6858) <= b and not a;
    outputs(6859) <= a and not b;
    outputs(6860) <= a xor b;
    outputs(6861) <= not b;
    outputs(6862) <= not (a xor b);
    outputs(6863) <= not (a and b);
    outputs(6864) <= a and not b;
    outputs(6865) <= a xor b;
    outputs(6866) <= not b;
    outputs(6867) <= b;
    outputs(6868) <= a xor b;
    outputs(6869) <= a and b;
    outputs(6870) <= a;
    outputs(6871) <= not (a xor b);
    outputs(6872) <= not b;
    outputs(6873) <= not (a xor b);
    outputs(6874) <= a or b;
    outputs(6875) <= b and not a;
    outputs(6876) <= not (a xor b);
    outputs(6877) <= b;
    outputs(6878) <= not b;
    outputs(6879) <= a xor b;
    outputs(6880) <= not a;
    outputs(6881) <= b and not a;
    outputs(6882) <= not a;
    outputs(6883) <= a;
    outputs(6884) <= not b;
    outputs(6885) <= a xor b;
    outputs(6886) <= a;
    outputs(6887) <= a;
    outputs(6888) <= not a;
    outputs(6889) <= b;
    outputs(6890) <= a xor b;
    outputs(6891) <= a xor b;
    outputs(6892) <= a and b;
    outputs(6893) <= not b;
    outputs(6894) <= not b;
    outputs(6895) <= not (a xor b);
    outputs(6896) <= a and not b;
    outputs(6897) <= a xor b;
    outputs(6898) <= not a;
    outputs(6899) <= a and b;
    outputs(6900) <= not b;
    outputs(6901) <= b;
    outputs(6902) <= not a;
    outputs(6903) <= a;
    outputs(6904) <= a xor b;
    outputs(6905) <= a and not b;
    outputs(6906) <= a or b;
    outputs(6907) <= not a;
    outputs(6908) <= not a;
    outputs(6909) <= a;
    outputs(6910) <= b and not a;
    outputs(6911) <= not b;
    outputs(6912) <= a xor b;
    outputs(6913) <= a and not b;
    outputs(6914) <= a;
    outputs(6915) <= a xor b;
    outputs(6916) <= a;
    outputs(6917) <= a and not b;
    outputs(6918) <= not b;
    outputs(6919) <= a and b;
    outputs(6920) <= not (a or b);
    outputs(6921) <= not (a and b);
    outputs(6922) <= not a;
    outputs(6923) <= a xor b;
    outputs(6924) <= a;
    outputs(6925) <= not a;
    outputs(6926) <= not a;
    outputs(6927) <= a and not b;
    outputs(6928) <= not (a or b);
    outputs(6929) <= not (a xor b);
    outputs(6930) <= a xor b;
    outputs(6931) <= a xor b;
    outputs(6932) <= a and b;
    outputs(6933) <= not (a and b);
    outputs(6934) <= not b;
    outputs(6935) <= a;
    outputs(6936) <= not b;
    outputs(6937) <= not (a or b);
    outputs(6938) <= a and not b;
    outputs(6939) <= not (a and b);
    outputs(6940) <= b;
    outputs(6941) <= not a;
    outputs(6942) <= not b;
    outputs(6943) <= not (a and b);
    outputs(6944) <= a xor b;
    outputs(6945) <= not b;
    outputs(6946) <= b;
    outputs(6947) <= b and not a;
    outputs(6948) <= not (a and b);
    outputs(6949) <= not b;
    outputs(6950) <= a and not b;
    outputs(6951) <= a or b;
    outputs(6952) <= not (a xor b);
    outputs(6953) <= not a;
    outputs(6954) <= b and not a;
    outputs(6955) <= not a or b;
    outputs(6956) <= a;
    outputs(6957) <= b and not a;
    outputs(6958) <= b;
    outputs(6959) <= not b or a;
    outputs(6960) <= not a;
    outputs(6961) <= not b;
    outputs(6962) <= not (a xor b);
    outputs(6963) <= a or b;
    outputs(6964) <= not (a xor b);
    outputs(6965) <= a or b;
    outputs(6966) <= a or b;
    outputs(6967) <= a and not b;
    outputs(6968) <= a;
    outputs(6969) <= a;
    outputs(6970) <= a and not b;
    outputs(6971) <= a xor b;
    outputs(6972) <= b;
    outputs(6973) <= a and not b;
    outputs(6974) <= not a;
    outputs(6975) <= a xor b;
    outputs(6976) <= a and not b;
    outputs(6977) <= not b;
    outputs(6978) <= a xor b;
    outputs(6979) <= not (a xor b);
    outputs(6980) <= a;
    outputs(6981) <= not (a xor b);
    outputs(6982) <= b;
    outputs(6983) <= not a;
    outputs(6984) <= not a;
    outputs(6985) <= not (a or b);
    outputs(6986) <= b and not a;
    outputs(6987) <= a;
    outputs(6988) <= a;
    outputs(6989) <= not a;
    outputs(6990) <= a xor b;
    outputs(6991) <= not b;
    outputs(6992) <= not a;
    outputs(6993) <= b;
    outputs(6994) <= not a;
    outputs(6995) <= not (a xor b);
    outputs(6996) <= b;
    outputs(6997) <= not a;
    outputs(6998) <= a xor b;
    outputs(6999) <= not b;
    outputs(7000) <= a;
    outputs(7001) <= a;
    outputs(7002) <= a xor b;
    outputs(7003) <= not (a xor b);
    outputs(7004) <= a xor b;
    outputs(7005) <= a and b;
    outputs(7006) <= not b;
    outputs(7007) <= not a;
    outputs(7008) <= not b;
    outputs(7009) <= b and not a;
    outputs(7010) <= a and not b;
    outputs(7011) <= not (a xor b);
    outputs(7012) <= not a or b;
    outputs(7013) <= not a;
    outputs(7014) <= not b;
    outputs(7015) <= not b;
    outputs(7016) <= a and b;
    outputs(7017) <= b and not a;
    outputs(7018) <= a xor b;
    outputs(7019) <= b and not a;
    outputs(7020) <= b;
    outputs(7021) <= not (a xor b);
    outputs(7022) <= not b;
    outputs(7023) <= not (a or b);
    outputs(7024) <= not b or a;
    outputs(7025) <= b and not a;
    outputs(7026) <= a;
    outputs(7027) <= a xor b;
    outputs(7028) <= b and not a;
    outputs(7029) <= b;
    outputs(7030) <= a;
    outputs(7031) <= a xor b;
    outputs(7032) <= a xor b;
    outputs(7033) <= not b;
    outputs(7034) <= not (a xor b);
    outputs(7035) <= b and not a;
    outputs(7036) <= not a;
    outputs(7037) <= a;
    outputs(7038) <= a or b;
    outputs(7039) <= a and b;
    outputs(7040) <= a xor b;
    outputs(7041) <= a xor b;
    outputs(7042) <= b and not a;
    outputs(7043) <= a;
    outputs(7044) <= not a;
    outputs(7045) <= not a;
    outputs(7046) <= a;
    outputs(7047) <= b;
    outputs(7048) <= b;
    outputs(7049) <= a xor b;
    outputs(7050) <= a and not b;
    outputs(7051) <= a xor b;
    outputs(7052) <= b and not a;
    outputs(7053) <= not (a or b);
    outputs(7054) <= not a or b;
    outputs(7055) <= b;
    outputs(7056) <= not b;
    outputs(7057) <= not (a or b);
    outputs(7058) <= not b;
    outputs(7059) <= not (a xor b);
    outputs(7060) <= a xor b;
    outputs(7061) <= b;
    outputs(7062) <= b and not a;
    outputs(7063) <= a xor b;
    outputs(7064) <= b;
    outputs(7065) <= a xor b;
    outputs(7066) <= not (a and b);
    outputs(7067) <= b;
    outputs(7068) <= not (a xor b);
    outputs(7069) <= b and not a;
    outputs(7070) <= a and not b;
    outputs(7071) <= a or b;
    outputs(7072) <= not b or a;
    outputs(7073) <= not (a and b);
    outputs(7074) <= not (a xor b);
    outputs(7075) <= a and not b;
    outputs(7076) <= b and not a;
    outputs(7077) <= a xor b;
    outputs(7078) <= not (a xor b);
    outputs(7079) <= not b;
    outputs(7080) <= not a;
    outputs(7081) <= a;
    outputs(7082) <= b;
    outputs(7083) <= a xor b;
    outputs(7084) <= not b or a;
    outputs(7085) <= not a;
    outputs(7086) <= not b or a;
    outputs(7087) <= not a;
    outputs(7088) <= a;
    outputs(7089) <= a and not b;
    outputs(7090) <= not (a xor b);
    outputs(7091) <= a;
    outputs(7092) <= a xor b;
    outputs(7093) <= not a;
    outputs(7094) <= b;
    outputs(7095) <= not a;
    outputs(7096) <= not a or b;
    outputs(7097) <= b;
    outputs(7098) <= b and not a;
    outputs(7099) <= b;
    outputs(7100) <= b;
    outputs(7101) <= b;
    outputs(7102) <= a xor b;
    outputs(7103) <= not a;
    outputs(7104) <= not (a xor b);
    outputs(7105) <= a xor b;
    outputs(7106) <= a;
    outputs(7107) <= not b;
    outputs(7108) <= b;
    outputs(7109) <= a xor b;
    outputs(7110) <= not (a xor b);
    outputs(7111) <= a or b;
    outputs(7112) <= not b or a;
    outputs(7113) <= a xor b;
    outputs(7114) <= b;
    outputs(7115) <= b;
    outputs(7116) <= not a;
    outputs(7117) <= not a or b;
    outputs(7118) <= a and not b;
    outputs(7119) <= a xor b;
    outputs(7120) <= not (a xor b);
    outputs(7121) <= a xor b;
    outputs(7122) <= a;
    outputs(7123) <= a xor b;
    outputs(7124) <= a xor b;
    outputs(7125) <= b;
    outputs(7126) <= not a;
    outputs(7127) <= not a or b;
    outputs(7128) <= not b;
    outputs(7129) <= a;
    outputs(7130) <= not b;
    outputs(7131) <= a;
    outputs(7132) <= a;
    outputs(7133) <= not b;
    outputs(7134) <= not b;
    outputs(7135) <= not a;
    outputs(7136) <= a and b;
    outputs(7137) <= a xor b;
    outputs(7138) <= not b;
    outputs(7139) <= not a;
    outputs(7140) <= a xor b;
    outputs(7141) <= not a or b;
    outputs(7142) <= not (a xor b);
    outputs(7143) <= not (a xor b);
    outputs(7144) <= a xor b;
    outputs(7145) <= b and not a;
    outputs(7146) <= not a;
    outputs(7147) <= b and not a;
    outputs(7148) <= a xor b;
    outputs(7149) <= not (a or b);
    outputs(7150) <= a and b;
    outputs(7151) <= not (a xor b);
    outputs(7152) <= not a;
    outputs(7153) <= a xor b;
    outputs(7154) <= a and not b;
    outputs(7155) <= a;
    outputs(7156) <= b;
    outputs(7157) <= not b;
    outputs(7158) <= not (a or b);
    outputs(7159) <= b;
    outputs(7160) <= not b;
    outputs(7161) <= not b;
    outputs(7162) <= not (a xor b);
    outputs(7163) <= not b;
    outputs(7164) <= a;
    outputs(7165) <= a xor b;
    outputs(7166) <= a;
    outputs(7167) <= not (a xor b);
    outputs(7168) <= not (a xor b);
    outputs(7169) <= b;
    outputs(7170) <= b and not a;
    outputs(7171) <= not a or b;
    outputs(7172) <= not b;
    outputs(7173) <= not (a xor b);
    outputs(7174) <= not b;
    outputs(7175) <= not (a xor b);
    outputs(7176) <= a xor b;
    outputs(7177) <= not a;
    outputs(7178) <= a;
    outputs(7179) <= b;
    outputs(7180) <= b;
    outputs(7181) <= not (a xor b);
    outputs(7182) <= not (a xor b);
    outputs(7183) <= a and b;
    outputs(7184) <= not a or b;
    outputs(7185) <= a;
    outputs(7186) <= not a;
    outputs(7187) <= b;
    outputs(7188) <= not (a or b);
    outputs(7189) <= a;
    outputs(7190) <= a;
    outputs(7191) <= a and not b;
    outputs(7192) <= not b;
    outputs(7193) <= b and not a;
    outputs(7194) <= not b or a;
    outputs(7195) <= b;
    outputs(7196) <= a and not b;
    outputs(7197) <= not (a or b);
    outputs(7198) <= a or b;
    outputs(7199) <= b;
    outputs(7200) <= a and not b;
    outputs(7201) <= not a or b;
    outputs(7202) <= not a;
    outputs(7203) <= a;
    outputs(7204) <= a and b;
    outputs(7205) <= not (a xor b);
    outputs(7206) <= not b;
    outputs(7207) <= not (a xor b);
    outputs(7208) <= a and b;
    outputs(7209) <= not (a or b);
    outputs(7210) <= b;
    outputs(7211) <= a and not b;
    outputs(7212) <= a xor b;
    outputs(7213) <= not a;
    outputs(7214) <= b and not a;
    outputs(7215) <= a xor b;
    outputs(7216) <= not (a and b);
    outputs(7217) <= not (a xor b);
    outputs(7218) <= b and not a;
    outputs(7219) <= a and not b;
    outputs(7220) <= b;
    outputs(7221) <= a and b;
    outputs(7222) <= a xor b;
    outputs(7223) <= b and not a;
    outputs(7224) <= a;
    outputs(7225) <= a and b;
    outputs(7226) <= b;
    outputs(7227) <= b and not a;
    outputs(7228) <= a;
    outputs(7229) <= not (a or b);
    outputs(7230) <= a or b;
    outputs(7231) <= a xor b;
    outputs(7232) <= a xor b;
    outputs(7233) <= not (a xor b);
    outputs(7234) <= not b or a;
    outputs(7235) <= not b;
    outputs(7236) <= a xor b;
    outputs(7237) <= b and not a;
    outputs(7238) <= not a or b;
    outputs(7239) <= b and not a;
    outputs(7240) <= b;
    outputs(7241) <= not a;
    outputs(7242) <= b and not a;
    outputs(7243) <= a;
    outputs(7244) <= '0';
    outputs(7245) <= not (a xor b);
    outputs(7246) <= not (a and b);
    outputs(7247) <= a xor b;
    outputs(7248) <= not (a and b);
    outputs(7249) <= not b;
    outputs(7250) <= not b;
    outputs(7251) <= not a;
    outputs(7252) <= a;
    outputs(7253) <= not a or b;
    outputs(7254) <= not (a xor b);
    outputs(7255) <= not (a or b);
    outputs(7256) <= not b or a;
    outputs(7257) <= a xor b;
    outputs(7258) <= a and b;
    outputs(7259) <= a;
    outputs(7260) <= b;
    outputs(7261) <= a;
    outputs(7262) <= not a;
    outputs(7263) <= not a;
    outputs(7264) <= a or b;
    outputs(7265) <= a;
    outputs(7266) <= b;
    outputs(7267) <= not (a xor b);
    outputs(7268) <= not a;
    outputs(7269) <= not a;
    outputs(7270) <= a xor b;
    outputs(7271) <= not (a or b);
    outputs(7272) <= a or b;
    outputs(7273) <= not b;
    outputs(7274) <= not a;
    outputs(7275) <= not (a and b);
    outputs(7276) <= b and not a;
    outputs(7277) <= a;
    outputs(7278) <= a;
    outputs(7279) <= not (a or b);
    outputs(7280) <= b;
    outputs(7281) <= not a;
    outputs(7282) <= a;
    outputs(7283) <= not b;
    outputs(7284) <= not (a xor b);
    outputs(7285) <= not b;
    outputs(7286) <= b;
    outputs(7287) <= a xor b;
    outputs(7288) <= b and not a;
    outputs(7289) <= a or b;
    outputs(7290) <= not (a and b);
    outputs(7291) <= a xor b;
    outputs(7292) <= not (a xor b);
    outputs(7293) <= a xor b;
    outputs(7294) <= a xor b;
    outputs(7295) <= b;
    outputs(7296) <= a xor b;
    outputs(7297) <= not a;
    outputs(7298) <= b;
    outputs(7299) <= not (a or b);
    outputs(7300) <= a or b;
    outputs(7301) <= not (a xor b);
    outputs(7302) <= b and not a;
    outputs(7303) <= a or b;
    outputs(7304) <= not b;
    outputs(7305) <= b and not a;
    outputs(7306) <= a;
    outputs(7307) <= a and b;
    outputs(7308) <= b;
    outputs(7309) <= a xor b;
    outputs(7310) <= b;
    outputs(7311) <= not b or a;
    outputs(7312) <= a;
    outputs(7313) <= not (a or b);
    outputs(7314) <= not (a or b);
    outputs(7315) <= a and b;
    outputs(7316) <= b and not a;
    outputs(7317) <= a or b;
    outputs(7318) <= a;
    outputs(7319) <= not (a xor b);
    outputs(7320) <= a;
    outputs(7321) <= not (a or b);
    outputs(7322) <= b and not a;
    outputs(7323) <= a;
    outputs(7324) <= b and not a;
    outputs(7325) <= a;
    outputs(7326) <= not a;
    outputs(7327) <= a and b;
    outputs(7328) <= a xor b;
    outputs(7329) <= not (a and b);
    outputs(7330) <= a xor b;
    outputs(7331) <= a;
    outputs(7332) <= not b or a;
    outputs(7333) <= not b or a;
    outputs(7334) <= not b;
    outputs(7335) <= not b;
    outputs(7336) <= not a;
    outputs(7337) <= a and not b;
    outputs(7338) <= not (a or b);
    outputs(7339) <= a xor b;
    outputs(7340) <= b and not a;
    outputs(7341) <= b;
    outputs(7342) <= a and b;
    outputs(7343) <= not b;
    outputs(7344) <= a and b;
    outputs(7345) <= not (a or b);
    outputs(7346) <= b;
    outputs(7347) <= b and not a;
    outputs(7348) <= a and not b;
    outputs(7349) <= a and not b;
    outputs(7350) <= not a;
    outputs(7351) <= b;
    outputs(7352) <= not b or a;
    outputs(7353) <= not a;
    outputs(7354) <= a and not b;
    outputs(7355) <= a;
    outputs(7356) <= b and not a;
    outputs(7357) <= a xor b;
    outputs(7358) <= a xor b;
    outputs(7359) <= not b;
    outputs(7360) <= a and not b;
    outputs(7361) <= b;
    outputs(7362) <= b;
    outputs(7363) <= a and b;
    outputs(7364) <= not b;
    outputs(7365) <= not a;
    outputs(7366) <= a and not b;
    outputs(7367) <= not b;
    outputs(7368) <= not (a xor b);
    outputs(7369) <= a xor b;
    outputs(7370) <= b;
    outputs(7371) <= not (a or b);
    outputs(7372) <= a xor b;
    outputs(7373) <= a or b;
    outputs(7374) <= not b;
    outputs(7375) <= a and not b;
    outputs(7376) <= a and not b;
    outputs(7377) <= a xor b;
    outputs(7378) <= b;
    outputs(7379) <= b;
    outputs(7380) <= a;
    outputs(7381) <= not b;
    outputs(7382) <= not b;
    outputs(7383) <= b;
    outputs(7384) <= not b;
    outputs(7385) <= a;
    outputs(7386) <= a;
    outputs(7387) <= not b;
    outputs(7388) <= a;
    outputs(7389) <= a;
    outputs(7390) <= b and not a;
    outputs(7391) <= not a;
    outputs(7392) <= a;
    outputs(7393) <= a and not b;
    outputs(7394) <= a;
    outputs(7395) <= not a;
    outputs(7396) <= a and not b;
    outputs(7397) <= not (a and b);
    outputs(7398) <= b;
    outputs(7399) <= a xor b;
    outputs(7400) <= a and not b;
    outputs(7401) <= not (a xor b);
    outputs(7402) <= b;
    outputs(7403) <= a;
    outputs(7404) <= b;
    outputs(7405) <= a xor b;
    outputs(7406) <= a;
    outputs(7407) <= a xor b;
    outputs(7408) <= a and b;
    outputs(7409) <= not (a or b);
    outputs(7410) <= not (a xor b);
    outputs(7411) <= b and not a;
    outputs(7412) <= not a;
    outputs(7413) <= b;
    outputs(7414) <= a xor b;
    outputs(7415) <= b;
    outputs(7416) <= b and not a;
    outputs(7417) <= b;
    outputs(7418) <= not b or a;
    outputs(7419) <= a and not b;
    outputs(7420) <= not a;
    outputs(7421) <= not a or b;
    outputs(7422) <= b;
    outputs(7423) <= not b;
    outputs(7424) <= not b;
    outputs(7425) <= not b;
    outputs(7426) <= not b;
    outputs(7427) <= a xor b;
    outputs(7428) <= not (a or b);
    outputs(7429) <= a;
    outputs(7430) <= b;
    outputs(7431) <= b;
    outputs(7432) <= b;
    outputs(7433) <= not (a xor b);
    outputs(7434) <= a;
    outputs(7435) <= not (a xor b);
    outputs(7436) <= not b or a;
    outputs(7437) <= a xor b;
    outputs(7438) <= not (a xor b);
    outputs(7439) <= a xor b;
    outputs(7440) <= b;
    outputs(7441) <= a and not b;
    outputs(7442) <= b;
    outputs(7443) <= b;
    outputs(7444) <= b;
    outputs(7445) <= not (a or b);
    outputs(7446) <= not (a xor b);
    outputs(7447) <= a and not b;
    outputs(7448) <= a xor b;
    outputs(7449) <= b;
    outputs(7450) <= a;
    outputs(7451) <= a;
    outputs(7452) <= a;
    outputs(7453) <= not a;
    outputs(7454) <= a and not b;
    outputs(7455) <= a xor b;
    outputs(7456) <= b;
    outputs(7457) <= b;
    outputs(7458) <= not a;
    outputs(7459) <= not (a or b);
    outputs(7460) <= not (a and b);
    outputs(7461) <= not a;
    outputs(7462) <= a and not b;
    outputs(7463) <= not (a and b);
    outputs(7464) <= a xor b;
    outputs(7465) <= b;
    outputs(7466) <= a or b;
    outputs(7467) <= b and not a;
    outputs(7468) <= not (a xor b);
    outputs(7469) <= not b;
    outputs(7470) <= not (a xor b);
    outputs(7471) <= b;
    outputs(7472) <= not (a or b);
    outputs(7473) <= a xor b;
    outputs(7474) <= a and not b;
    outputs(7475) <= not (a xor b);
    outputs(7476) <= a;
    outputs(7477) <= b and not a;
    outputs(7478) <= a xor b;
    outputs(7479) <= not b;
    outputs(7480) <= not (a xor b);
    outputs(7481) <= a xor b;
    outputs(7482) <= not b or a;
    outputs(7483) <= not a;
    outputs(7484) <= not b;
    outputs(7485) <= a xor b;
    outputs(7486) <= a and b;
    outputs(7487) <= b;
    outputs(7488) <= not (a xor b);
    outputs(7489) <= not (a or b);
    outputs(7490) <= not (a and b);
    outputs(7491) <= not (a xor b);
    outputs(7492) <= a and b;
    outputs(7493) <= b;
    outputs(7494) <= not a;
    outputs(7495) <= b;
    outputs(7496) <= a;
    outputs(7497) <= a and not b;
    outputs(7498) <= b;
    outputs(7499) <= a and b;
    outputs(7500) <= b and not a;
    outputs(7501) <= a;
    outputs(7502) <= a xor b;
    outputs(7503) <= a;
    outputs(7504) <= not (a or b);
    outputs(7505) <= b;
    outputs(7506) <= a;
    outputs(7507) <= not a or b;
    outputs(7508) <= b;
    outputs(7509) <= not a;
    outputs(7510) <= not (a xor b);
    outputs(7511) <= not (a xor b);
    outputs(7512) <= a and b;
    outputs(7513) <= b;
    outputs(7514) <= not (a or b);
    outputs(7515) <= a;
    outputs(7516) <= not (a xor b);
    outputs(7517) <= a xor b;
    outputs(7518) <= a and b;
    outputs(7519) <= not (a and b);
    outputs(7520) <= b and not a;
    outputs(7521) <= not b;
    outputs(7522) <= not b;
    outputs(7523) <= b and not a;
    outputs(7524) <= a xor b;
    outputs(7525) <= not (a xor b);
    outputs(7526) <= a;
    outputs(7527) <= a xor b;
    outputs(7528) <= b;
    outputs(7529) <= a;
    outputs(7530) <= not b;
    outputs(7531) <= a xor b;
    outputs(7532) <= not (a xor b);
    outputs(7533) <= a;
    outputs(7534) <= b;
    outputs(7535) <= not (a xor b);
    outputs(7536) <= not (a xor b);
    outputs(7537) <= a;
    outputs(7538) <= a;
    outputs(7539) <= a;
    outputs(7540) <= not (a xor b);
    outputs(7541) <= not b;
    outputs(7542) <= a;
    outputs(7543) <= a;
    outputs(7544) <= a and not b;
    outputs(7545) <= b and not a;
    outputs(7546) <= a;
    outputs(7547) <= b;
    outputs(7548) <= not a;
    outputs(7549) <= a xor b;
    outputs(7550) <= not b;
    outputs(7551) <= a and b;
    outputs(7552) <= b;
    outputs(7553) <= not (a xor b);
    outputs(7554) <= a and not b;
    outputs(7555) <= not b;
    outputs(7556) <= not a;
    outputs(7557) <= not (a or b);
    outputs(7558) <= b;
    outputs(7559) <= not b;
    outputs(7560) <= a xor b;
    outputs(7561) <= a and not b;
    outputs(7562) <= a or b;
    outputs(7563) <= not a;
    outputs(7564) <= not b;
    outputs(7565) <= not b;
    outputs(7566) <= a and b;
    outputs(7567) <= not b or a;
    outputs(7568) <= a and b;
    outputs(7569) <= a xor b;
    outputs(7570) <= not b;
    outputs(7571) <= b and not a;
    outputs(7572) <= not (a xor b);
    outputs(7573) <= b and not a;
    outputs(7574) <= not a;
    outputs(7575) <= a and b;
    outputs(7576) <= b and not a;
    outputs(7577) <= b and not a;
    outputs(7578) <= a and b;
    outputs(7579) <= b and not a;
    outputs(7580) <= not a;
    outputs(7581) <= a and not b;
    outputs(7582) <= not b;
    outputs(7583) <= a and not b;
    outputs(7584) <= b and not a;
    outputs(7585) <= a and not b;
    outputs(7586) <= not a;
    outputs(7587) <= not a;
    outputs(7588) <= not b;
    outputs(7589) <= a;
    outputs(7590) <= a and b;
    outputs(7591) <= a xor b;
    outputs(7592) <= a xor b;
    outputs(7593) <= a xor b;
    outputs(7594) <= not (a or b);
    outputs(7595) <= a xor b;
    outputs(7596) <= not (a xor b);
    outputs(7597) <= a xor b;
    outputs(7598) <= a and not b;
    outputs(7599) <= b;
    outputs(7600) <= not (a xor b);
    outputs(7601) <= not (a xor b);
    outputs(7602) <= a;
    outputs(7603) <= not (a and b);
    outputs(7604) <= not (a xor b);
    outputs(7605) <= b and not a;
    outputs(7606) <= not (a or b);
    outputs(7607) <= not (a xor b);
    outputs(7608) <= not (a or b);
    outputs(7609) <= b and not a;
    outputs(7610) <= a xor b;
    outputs(7611) <= a;
    outputs(7612) <= b;
    outputs(7613) <= a;
    outputs(7614) <= a;
    outputs(7615) <= a and b;
    outputs(7616) <= a xor b;
    outputs(7617) <= a or b;
    outputs(7618) <= not b or a;
    outputs(7619) <= a xor b;
    outputs(7620) <= not (a xor b);
    outputs(7621) <= b and not a;
    outputs(7622) <= a xor b;
    outputs(7623) <= a xor b;
    outputs(7624) <= b and not a;
    outputs(7625) <= b;
    outputs(7626) <= a;
    outputs(7627) <= a;
    outputs(7628) <= b;
    outputs(7629) <= not (a xor b);
    outputs(7630) <= a and not b;
    outputs(7631) <= b;
    outputs(7632) <= not (a xor b);
    outputs(7633) <= a and b;
    outputs(7634) <= a and b;
    outputs(7635) <= b and not a;
    outputs(7636) <= b and not a;
    outputs(7637) <= not a;
    outputs(7638) <= b and not a;
    outputs(7639) <= b and not a;
    outputs(7640) <= a or b;
    outputs(7641) <= a xor b;
    outputs(7642) <= b;
    outputs(7643) <= a;
    outputs(7644) <= a xor b;
    outputs(7645) <= a xor b;
    outputs(7646) <= not b or a;
    outputs(7647) <= a and b;
    outputs(7648) <= not a or b;
    outputs(7649) <= a xor b;
    outputs(7650) <= not a;
    outputs(7651) <= not b;
    outputs(7652) <= b;
    outputs(7653) <= b;
    outputs(7654) <= not (a xor b);
    outputs(7655) <= a xor b;
    outputs(7656) <= not a;
    outputs(7657) <= b and not a;
    outputs(7658) <= a and b;
    outputs(7659) <= not a;
    outputs(7660) <= not (a xor b);
    outputs(7661) <= not b or a;
    outputs(7662) <= not (a or b);
    outputs(7663) <= not (a xor b);
    outputs(7664) <= a;
    outputs(7665) <= a xor b;
    outputs(7666) <= b;
    outputs(7667) <= a xor b;
    outputs(7668) <= a xor b;
    outputs(7669) <= a and b;
    outputs(7670) <= a;
    outputs(7671) <= not a;
    outputs(7672) <= a xor b;
    outputs(7673) <= not (a and b);
    outputs(7674) <= a;
    outputs(7675) <= a;
    outputs(7676) <= a and b;
    outputs(7677) <= a and not b;
    outputs(7678) <= not a;
    outputs(7679) <= a and b;
    outputs(7680) <= a xor b;
    outputs(7681) <= b and not a;
    outputs(7682) <= not b;
    outputs(7683) <= not a;
    outputs(7684) <= b;
    outputs(7685) <= not (a and b);
    outputs(7686) <= not (a and b);
    outputs(7687) <= a xor b;
    outputs(7688) <= a and b;
    outputs(7689) <= not (a and b);
    outputs(7690) <= a;
    outputs(7691) <= a;
    outputs(7692) <= a xor b;
    outputs(7693) <= a xor b;
    outputs(7694) <= not (a or b);
    outputs(7695) <= not b;
    outputs(7696) <= not (a and b);
    outputs(7697) <= not a;
    outputs(7698) <= not a;
    outputs(7699) <= not (a xor b);
    outputs(7700) <= a xor b;
    outputs(7701) <= b;
    outputs(7702) <= a xor b;
    outputs(7703) <= a and b;
    outputs(7704) <= b;
    outputs(7705) <= not b;
    outputs(7706) <= b;
    outputs(7707) <= not b;
    outputs(7708) <= a and not b;
    outputs(7709) <= a;
    outputs(7710) <= not (a or b);
    outputs(7711) <= a and b;
    outputs(7712) <= not b or a;
    outputs(7713) <= a and b;
    outputs(7714) <= b;
    outputs(7715) <= a xor b;
    outputs(7716) <= a xor b;
    outputs(7717) <= a and b;
    outputs(7718) <= not a or b;
    outputs(7719) <= a and not b;
    outputs(7720) <= not b;
    outputs(7721) <= not (a xor b);
    outputs(7722) <= not (a xor b);
    outputs(7723) <= b;
    outputs(7724) <= not (a or b);
    outputs(7725) <= b and not a;
    outputs(7726) <= a;
    outputs(7727) <= not b or a;
    outputs(7728) <= not b;
    outputs(7729) <= b;
    outputs(7730) <= not a or b;
    outputs(7731) <= not b;
    outputs(7732) <= not a;
    outputs(7733) <= a and b;
    outputs(7734) <= a;
    outputs(7735) <= a xor b;
    outputs(7736) <= not b or a;
    outputs(7737) <= a xor b;
    outputs(7738) <= not a or b;
    outputs(7739) <= not a;
    outputs(7740) <= a xor b;
    outputs(7741) <= not (a or b);
    outputs(7742) <= a;
    outputs(7743) <= a;
    outputs(7744) <= b;
    outputs(7745) <= not a;
    outputs(7746) <= not b;
    outputs(7747) <= a;
    outputs(7748) <= b and not a;
    outputs(7749) <= not (a xor b);
    outputs(7750) <= not b or a;
    outputs(7751) <= b and not a;
    outputs(7752) <= a and not b;
    outputs(7753) <= not a;
    outputs(7754) <= b and not a;
    outputs(7755) <= not b or a;
    outputs(7756) <= not a or b;
    outputs(7757) <= a and b;
    outputs(7758) <= not b;
    outputs(7759) <= a and b;
    outputs(7760) <= a and b;
    outputs(7761) <= a or b;
    outputs(7762) <= a xor b;
    outputs(7763) <= not a;
    outputs(7764) <= not a or b;
    outputs(7765) <= not b;
    outputs(7766) <= b;
    outputs(7767) <= not (a xor b);
    outputs(7768) <= b and not a;
    outputs(7769) <= not (a xor b);
    outputs(7770) <= b;
    outputs(7771) <= a;
    outputs(7772) <= a and not b;
    outputs(7773) <= not (a and b);
    outputs(7774) <= a;
    outputs(7775) <= a xor b;
    outputs(7776) <= a xor b;
    outputs(7777) <= not a or b;
    outputs(7778) <= b and not a;
    outputs(7779) <= a;
    outputs(7780) <= b and not a;
    outputs(7781) <= not (a xor b);
    outputs(7782) <= not a;
    outputs(7783) <= a and b;
    outputs(7784) <= not (a or b);
    outputs(7785) <= a;
    outputs(7786) <= a;
    outputs(7787) <= b;
    outputs(7788) <= not (a xor b);
    outputs(7789) <= not (a xor b);
    outputs(7790) <= a;
    outputs(7791) <= a and not b;
    outputs(7792) <= a;
    outputs(7793) <= not a;
    outputs(7794) <= not (a xor b);
    outputs(7795) <= not (a xor b);
    outputs(7796) <= not b;
    outputs(7797) <= b;
    outputs(7798) <= a and b;
    outputs(7799) <= not a;
    outputs(7800) <= a xor b;
    outputs(7801) <= a or b;
    outputs(7802) <= b;
    outputs(7803) <= a and b;
    outputs(7804) <= a and b;
    outputs(7805) <= not b;
    outputs(7806) <= not (a xor b);
    outputs(7807) <= not (a xor b);
    outputs(7808) <= not b;
    outputs(7809) <= b and not a;
    outputs(7810) <= a xor b;
    outputs(7811) <= a and b;
    outputs(7812) <= not a or b;
    outputs(7813) <= not (a or b);
    outputs(7814) <= not (a or b);
    outputs(7815) <= not a;
    outputs(7816) <= not (a or b);
    outputs(7817) <= a;
    outputs(7818) <= a and not b;
    outputs(7819) <= not a;
    outputs(7820) <= a xor b;
    outputs(7821) <= b;
    outputs(7822) <= b and not a;
    outputs(7823) <= a and not b;
    outputs(7824) <= not (a xor b);
    outputs(7825) <= not (a xor b);
    outputs(7826) <= a and b;
    outputs(7827) <= not a or b;
    outputs(7828) <= not a or b;
    outputs(7829) <= b;
    outputs(7830) <= a and not b;
    outputs(7831) <= a xor b;
    outputs(7832) <= not b;
    outputs(7833) <= not b;
    outputs(7834) <= a;
    outputs(7835) <= a and b;
    outputs(7836) <= not (a xor b);
    outputs(7837) <= not a;
    outputs(7838) <= a xor b;
    outputs(7839) <= b;
    outputs(7840) <= not b;
    outputs(7841) <= a xor b;
    outputs(7842) <= not b or a;
    outputs(7843) <= not (a or b);
    outputs(7844) <= not b;
    outputs(7845) <= not b;
    outputs(7846) <= a;
    outputs(7847) <= not b;
    outputs(7848) <= not b;
    outputs(7849) <= not (a xor b);
    outputs(7850) <= a or b;
    outputs(7851) <= b;
    outputs(7852) <= a;
    outputs(7853) <= b and not a;
    outputs(7854) <= not a or b;
    outputs(7855) <= b and not a;
    outputs(7856) <= a;
    outputs(7857) <= not a;
    outputs(7858) <= a and b;
    outputs(7859) <= not a or b;
    outputs(7860) <= not a;
    outputs(7861) <= not b;
    outputs(7862) <= not (a or b);
    outputs(7863) <= a and not b;
    outputs(7864) <= not b;
    outputs(7865) <= not (a xor b);
    outputs(7866) <= a or b;
    outputs(7867) <= not a;
    outputs(7868) <= a and b;
    outputs(7869) <= a or b;
    outputs(7870) <= not (a and b);
    outputs(7871) <= not a or b;
    outputs(7872) <= not b;
    outputs(7873) <= not (a xor b);
    outputs(7874) <= b;
    outputs(7875) <= not (a xor b);
    outputs(7876) <= not b;
    outputs(7877) <= a;
    outputs(7878) <= not b or a;
    outputs(7879) <= a and not b;
    outputs(7880) <= not (a or b);
    outputs(7881) <= not b;
    outputs(7882) <= not (a or b);
    outputs(7883) <= not a;
    outputs(7884) <= a;
    outputs(7885) <= not b;
    outputs(7886) <= not b;
    outputs(7887) <= a;
    outputs(7888) <= a and not b;
    outputs(7889) <= not (a xor b);
    outputs(7890) <= not a;
    outputs(7891) <= a and not b;
    outputs(7892) <= a and b;
    outputs(7893) <= not b;
    outputs(7894) <= a;
    outputs(7895) <= not (a xor b);
    outputs(7896) <= b;
    outputs(7897) <= b;
    outputs(7898) <= a xor b;
    outputs(7899) <= a or b;
    outputs(7900) <= not a;
    outputs(7901) <= not (a xor b);
    outputs(7902) <= not (a xor b);
    outputs(7903) <= not (a or b);
    outputs(7904) <= not b or a;
    outputs(7905) <= not a;
    outputs(7906) <= not a;
    outputs(7907) <= b;
    outputs(7908) <= not a;
    outputs(7909) <= not b;
    outputs(7910) <= a xor b;
    outputs(7911) <= not (a xor b);
    outputs(7912) <= a and b;
    outputs(7913) <= not (a and b);
    outputs(7914) <= a;
    outputs(7915) <= a;
    outputs(7916) <= b;
    outputs(7917) <= b;
    outputs(7918) <= a;
    outputs(7919) <= not (a xor b);
    outputs(7920) <= not a;
    outputs(7921) <= not a;
    outputs(7922) <= not (a and b);
    outputs(7923) <= a xor b;
    outputs(7924) <= a;
    outputs(7925) <= a and not b;
    outputs(7926) <= a;
    outputs(7927) <= not (a xor b);
    outputs(7928) <= a xor b;
    outputs(7929) <= b;
    outputs(7930) <= not a;
    outputs(7931) <= b and not a;
    outputs(7932) <= b;
    outputs(7933) <= b and not a;
    outputs(7934) <= b and not a;
    outputs(7935) <= b;
    outputs(7936) <= not a;
    outputs(7937) <= not b;
    outputs(7938) <= a;
    outputs(7939) <= not b;
    outputs(7940) <= not b;
    outputs(7941) <= a xor b;
    outputs(7942) <= a xor b;
    outputs(7943) <= not (a and b);
    outputs(7944) <= not (a or b);
    outputs(7945) <= not b;
    outputs(7946) <= a xor b;
    outputs(7947) <= a and b;
    outputs(7948) <= b;
    outputs(7949) <= not b;
    outputs(7950) <= a and b;
    outputs(7951) <= a and b;
    outputs(7952) <= a and not b;
    outputs(7953) <= not (a or b);
    outputs(7954) <= b;
    outputs(7955) <= b and not a;
    outputs(7956) <= a and not b;
    outputs(7957) <= not a or b;
    outputs(7958) <= a xor b;
    outputs(7959) <= a;
    outputs(7960) <= a or b;
    outputs(7961) <= a and not b;
    outputs(7962) <= not b;
    outputs(7963) <= a and b;
    outputs(7964) <= b;
    outputs(7965) <= not b or a;
    outputs(7966) <= not (a xor b);
    outputs(7967) <= a xor b;
    outputs(7968) <= b;
    outputs(7969) <= a;
    outputs(7970) <= a;
    outputs(7971) <= a and b;
    outputs(7972) <= not a;
    outputs(7973) <= not b;
    outputs(7974) <= b;
    outputs(7975) <= not a or b;
    outputs(7976) <= not a;
    outputs(7977) <= a and b;
    outputs(7978) <= a xor b;
    outputs(7979) <= a;
    outputs(7980) <= a and b;
    outputs(7981) <= a and not b;
    outputs(7982) <= not b;
    outputs(7983) <= a;
    outputs(7984) <= a;
    outputs(7985) <= b and not a;
    outputs(7986) <= a xor b;
    outputs(7987) <= not (a or b);
    outputs(7988) <= a;
    outputs(7989) <= not b;
    outputs(7990) <= not (a xor b);
    outputs(7991) <= not a;
    outputs(7992) <= b;
    outputs(7993) <= not b;
    outputs(7994) <= a and b;
    outputs(7995) <= not a;
    outputs(7996) <= not b;
    outputs(7997) <= not a;
    outputs(7998) <= not b;
    outputs(7999) <= not b;
    outputs(8000) <= not (a or b);
    outputs(8001) <= not (a xor b);
    outputs(8002) <= a and not b;
    outputs(8003) <= not (a xor b);
    outputs(8004) <= not a;
    outputs(8005) <= a and b;
    outputs(8006) <= a and b;
    outputs(8007) <= b;
    outputs(8008) <= not (a or b);
    outputs(8009) <= a or b;
    outputs(8010) <= a;
    outputs(8011) <= not a;
    outputs(8012) <= a and not b;
    outputs(8013) <= a xor b;
    outputs(8014) <= not a;
    outputs(8015) <= a xor b;
    outputs(8016) <= a and not b;
    outputs(8017) <= not (a and b);
    outputs(8018) <= not a;
    outputs(8019) <= a;
    outputs(8020) <= a;
    outputs(8021) <= not b;
    outputs(8022) <= a xor b;
    outputs(8023) <= a;
    outputs(8024) <= a and b;
    outputs(8025) <= a and not b;
    outputs(8026) <= b;
    outputs(8027) <= not b;
    outputs(8028) <= b;
    outputs(8029) <= not a;
    outputs(8030) <= a and b;
    outputs(8031) <= not (a and b);
    outputs(8032) <= a xor b;
    outputs(8033) <= not a;
    outputs(8034) <= a xor b;
    outputs(8035) <= a;
    outputs(8036) <= a;
    outputs(8037) <= not b or a;
    outputs(8038) <= not (a xor b);
    outputs(8039) <= a xor b;
    outputs(8040) <= a xor b;
    outputs(8041) <= not (a xor b);
    outputs(8042) <= not a or b;
    outputs(8043) <= a xor b;
    outputs(8044) <= b;
    outputs(8045) <= b;
    outputs(8046) <= a or b;
    outputs(8047) <= a;
    outputs(8048) <= not a;
    outputs(8049) <= a xor b;
    outputs(8050) <= a;
    outputs(8051) <= not b;
    outputs(8052) <= not (a xor b);
    outputs(8053) <= a or b;
    outputs(8054) <= not (a and b);
    outputs(8055) <= a;
    outputs(8056) <= not a;
    outputs(8057) <= a or b;
    outputs(8058) <= not (a or b);
    outputs(8059) <= a or b;
    outputs(8060) <= not a;
    outputs(8061) <= not (a and b);
    outputs(8062) <= not (a xor b);
    outputs(8063) <= not (a or b);
    outputs(8064) <= not (a or b);
    outputs(8065) <= not a;
    outputs(8066) <= a xor b;
    outputs(8067) <= a or b;
    outputs(8068) <= a and not b;
    outputs(8069) <= a;
    outputs(8070) <= not b or a;
    outputs(8071) <= not a;
    outputs(8072) <= b;
    outputs(8073) <= a;
    outputs(8074) <= a;
    outputs(8075) <= not b;
    outputs(8076) <= a xor b;
    outputs(8077) <= b;
    outputs(8078) <= a xor b;
    outputs(8079) <= not (a or b);
    outputs(8080) <= a and b;
    outputs(8081) <= a;
    outputs(8082) <= not a;
    outputs(8083) <= not a;
    outputs(8084) <= b;
    outputs(8085) <= not (a or b);
    outputs(8086) <= a;
    outputs(8087) <= not (a xor b);
    outputs(8088) <= b;
    outputs(8089) <= b;
    outputs(8090) <= not (a xor b);
    outputs(8091) <= not b;
    outputs(8092) <= b;
    outputs(8093) <= a and b;
    outputs(8094) <= not a or b;
    outputs(8095) <= a xor b;
    outputs(8096) <= not (a xor b);
    outputs(8097) <= not a;
    outputs(8098) <= not b;
    outputs(8099) <= a xor b;
    outputs(8100) <= a xor b;
    outputs(8101) <= b;
    outputs(8102) <= a xor b;
    outputs(8103) <= a;
    outputs(8104) <= a and b;
    outputs(8105) <= not (a xor b);
    outputs(8106) <= b;
    outputs(8107) <= a and b;
    outputs(8108) <= a;
    outputs(8109) <= not b;
    outputs(8110) <= not a;
    outputs(8111) <= not a or b;
    outputs(8112) <= b and not a;
    outputs(8113) <= not (a or b);
    outputs(8114) <= b and not a;
    outputs(8115) <= not b;
    outputs(8116) <= a and b;
    outputs(8117) <= a xor b;
    outputs(8118) <= not (a or b);
    outputs(8119) <= b and not a;
    outputs(8120) <= b;
    outputs(8121) <= not (a xor b);
    outputs(8122) <= not b;
    outputs(8123) <= not (a xor b);
    outputs(8124) <= not a;
    outputs(8125) <= a and not b;
    outputs(8126) <= not (a xor b);
    outputs(8127) <= a;
    outputs(8128) <= not b;
    outputs(8129) <= a xor b;
    outputs(8130) <= a xor b;
    outputs(8131) <= a xor b;
    outputs(8132) <= not (a or b);
    outputs(8133) <= not (a or b);
    outputs(8134) <= a;
    outputs(8135) <= a xor b;
    outputs(8136) <= a or b;
    outputs(8137) <= a xor b;
    outputs(8138) <= not (a and b);
    outputs(8139) <= not (a and b);
    outputs(8140) <= not (a or b);
    outputs(8141) <= a and not b;
    outputs(8142) <= a and not b;
    outputs(8143) <= not b;
    outputs(8144) <= not (a and b);
    outputs(8145) <= not a;
    outputs(8146) <= not a;
    outputs(8147) <= not a;
    outputs(8148) <= a and not b;
    outputs(8149) <= not a;
    outputs(8150) <= a xor b;
    outputs(8151) <= not a;
    outputs(8152) <= b;
    outputs(8153) <= not (a xor b);
    outputs(8154) <= not (a or b);
    outputs(8155) <= a xor b;
    outputs(8156) <= b;
    outputs(8157) <= a xor b;
    outputs(8158) <= b and not a;
    outputs(8159) <= not a;
    outputs(8160) <= a or b;
    outputs(8161) <= b;
    outputs(8162) <= a;
    outputs(8163) <= not a or b;
    outputs(8164) <= not a;
    outputs(8165) <= b and not a;
    outputs(8166) <= b and not a;
    outputs(8167) <= a and b;
    outputs(8168) <= a;
    outputs(8169) <= a xor b;
    outputs(8170) <= a;
    outputs(8171) <= a and b;
    outputs(8172) <= a;
    outputs(8173) <= a;
    outputs(8174) <= a and b;
    outputs(8175) <= a and b;
    outputs(8176) <= not a;
    outputs(8177) <= a xor b;
    outputs(8178) <= a xor b;
    outputs(8179) <= b and not a;
    outputs(8180) <= a and not b;
    outputs(8181) <= b and not a;
    outputs(8182) <= not (a and b);
    outputs(8183) <= a or b;
    outputs(8184) <= a and b;
    outputs(8185) <= not (a or b);
    outputs(8186) <= not b or a;
    outputs(8187) <= not b;
    outputs(8188) <= b;
    outputs(8189) <= not (a xor b);
    outputs(8190) <= not (a xor b);
    outputs(8191) <= not a;
    outputs(8192) <= not (a xor b);
    outputs(8193) <= not b;
    outputs(8194) <= b;
    outputs(8195) <= a xor b;
    outputs(8196) <= a xor b;
    outputs(8197) <= not (a or b);
    outputs(8198) <= not b;
    outputs(8199) <= a xor b;
    outputs(8200) <= a xor b;
    outputs(8201) <= not b;
    outputs(8202) <= not b;
    outputs(8203) <= not b or a;
    outputs(8204) <= not b or a;
    outputs(8205) <= a xor b;
    outputs(8206) <= b;
    outputs(8207) <= b and not a;
    outputs(8208) <= a xor b;
    outputs(8209) <= not b;
    outputs(8210) <= a or b;
    outputs(8211) <= b;
    outputs(8212) <= a or b;
    outputs(8213) <= not a or b;
    outputs(8214) <= b and not a;
    outputs(8215) <= a or b;
    outputs(8216) <= not (a xor b);
    outputs(8217) <= a;
    outputs(8218) <= a xor b;
    outputs(8219) <= not (a or b);
    outputs(8220) <= not (a xor b);
    outputs(8221) <= a;
    outputs(8222) <= not b or a;
    outputs(8223) <= not (a xor b);
    outputs(8224) <= not a;
    outputs(8225) <= b and not a;
    outputs(8226) <= not (a xor b);
    outputs(8227) <= not (a xor b);
    outputs(8228) <= not (a xor b);
    outputs(8229) <= b;
    outputs(8230) <= a or b;
    outputs(8231) <= not a;
    outputs(8232) <= a or b;
    outputs(8233) <= not (a xor b);
    outputs(8234) <= a;
    outputs(8235) <= not a or b;
    outputs(8236) <= a or b;
    outputs(8237) <= a xor b;
    outputs(8238) <= b;
    outputs(8239) <= not (a xor b);
    outputs(8240) <= a and not b;
    outputs(8241) <= a;
    outputs(8242) <= a xor b;
    outputs(8243) <= a xor b;
    outputs(8244) <= not (a xor b);
    outputs(8245) <= b;
    outputs(8246) <= a xor b;
    outputs(8247) <= a xor b;
    outputs(8248) <= b;
    outputs(8249) <= a;
    outputs(8250) <= not (a or b);
    outputs(8251) <= b and not a;
    outputs(8252) <= not b;
    outputs(8253) <= not a;
    outputs(8254) <= not (a and b);
    outputs(8255) <= a xor b;
    outputs(8256) <= not (a and b);
    outputs(8257) <= not b or a;
    outputs(8258) <= a;
    outputs(8259) <= a xor b;
    outputs(8260) <= not a or b;
    outputs(8261) <= not a;
    outputs(8262) <= b and not a;
    outputs(8263) <= a and not b;
    outputs(8264) <= not (a and b);
    outputs(8265) <= a;
    outputs(8266) <= not b or a;
    outputs(8267) <= not (a xor b);
    outputs(8268) <= not a;
    outputs(8269) <= a xor b;
    outputs(8270) <= not (a xor b);
    outputs(8271) <= a;
    outputs(8272) <= b and not a;
    outputs(8273) <= not b or a;
    outputs(8274) <= b;
    outputs(8275) <= a or b;
    outputs(8276) <= not a or b;
    outputs(8277) <= not (a xor b);
    outputs(8278) <= b;
    outputs(8279) <= a and not b;
    outputs(8280) <= a xor b;
    outputs(8281) <= not a;
    outputs(8282) <= not a;
    outputs(8283) <= not (a and b);
    outputs(8284) <= not a;
    outputs(8285) <= a or b;
    outputs(8286) <= b;
    outputs(8287) <= a;
    outputs(8288) <= not a;
    outputs(8289) <= a or b;
    outputs(8290) <= a;
    outputs(8291) <= a xor b;
    outputs(8292) <= a xor b;
    outputs(8293) <= b;
    outputs(8294) <= not b or a;
    outputs(8295) <= not b;
    outputs(8296) <= not (a xor b);
    outputs(8297) <= not b;
    outputs(8298) <= a or b;
    outputs(8299) <= b;
    outputs(8300) <= not a;
    outputs(8301) <= a xor b;
    outputs(8302) <= not (a xor b);
    outputs(8303) <= a and b;
    outputs(8304) <= not (a xor b);
    outputs(8305) <= b;
    outputs(8306) <= a xor b;
    outputs(8307) <= not (a or b);
    outputs(8308) <= a or b;
    outputs(8309) <= not a or b;
    outputs(8310) <= a xor b;
    outputs(8311) <= a xor b;
    outputs(8312) <= a;
    outputs(8313) <= not (a or b);
    outputs(8314) <= a xor b;
    outputs(8315) <= not a;
    outputs(8316) <= b;
    outputs(8317) <= b and not a;
    outputs(8318) <= not (a xor b);
    outputs(8319) <= a;
    outputs(8320) <= not (a xor b);
    outputs(8321) <= b;
    outputs(8322) <= a xor b;
    outputs(8323) <= a;
    outputs(8324) <= not a;
    outputs(8325) <= b;
    outputs(8326) <= a;
    outputs(8327) <= not (a xor b);
    outputs(8328) <= b and not a;
    outputs(8329) <= not (a and b);
    outputs(8330) <= not a or b;
    outputs(8331) <= not (a or b);
    outputs(8332) <= a;
    outputs(8333) <= not (a xor b);
    outputs(8334) <= b;
    outputs(8335) <= not (a xor b);
    outputs(8336) <= not (a xor b);
    outputs(8337) <= not a;
    outputs(8338) <= not b;
    outputs(8339) <= not b or a;
    outputs(8340) <= a xor b;
    outputs(8341) <= not a;
    outputs(8342) <= a xor b;
    outputs(8343) <= not (a xor b);
    outputs(8344) <= a xor b;
    outputs(8345) <= a xor b;
    outputs(8346) <= not (a xor b);
    outputs(8347) <= a xor b;
    outputs(8348) <= a xor b;
    outputs(8349) <= not b;
    outputs(8350) <= a xor b;
    outputs(8351) <= not a;
    outputs(8352) <= not (a xor b);
    outputs(8353) <= not (a xor b);
    outputs(8354) <= a;
    outputs(8355) <= a and b;
    outputs(8356) <= not (a xor b);
    outputs(8357) <= not (a xor b);
    outputs(8358) <= not b;
    outputs(8359) <= b;
    outputs(8360) <= a xor b;
    outputs(8361) <= not a or b;
    outputs(8362) <= not a;
    outputs(8363) <= not (a or b);
    outputs(8364) <= a xor b;
    outputs(8365) <= b;
    outputs(8366) <= not (a or b);
    outputs(8367) <= a xor b;
    outputs(8368) <= a xor b;
    outputs(8369) <= a;
    outputs(8370) <= not b;
    outputs(8371) <= a xor b;
    outputs(8372) <= not a;
    outputs(8373) <= a and not b;
    outputs(8374) <= not a;
    outputs(8375) <= b;
    outputs(8376) <= b;
    outputs(8377) <= not (a xor b);
    outputs(8378) <= a xor b;
    outputs(8379) <= a;
    outputs(8380) <= a;
    outputs(8381) <= not (a xor b);
    outputs(8382) <= not (a xor b);
    outputs(8383) <= a;
    outputs(8384) <= a;
    outputs(8385) <= a xor b;
    outputs(8386) <= b;
    outputs(8387) <= not (a xor b);
    outputs(8388) <= not b;
    outputs(8389) <= not (a and b);
    outputs(8390) <= not b or a;
    outputs(8391) <= b;
    outputs(8392) <= not a or b;
    outputs(8393) <= not a;
    outputs(8394) <= not a;
    outputs(8395) <= not a;
    outputs(8396) <= a;
    outputs(8397) <= a xor b;
    outputs(8398) <= not (a xor b);
    outputs(8399) <= not b;
    outputs(8400) <= b;
    outputs(8401) <= a xor b;
    outputs(8402) <= not (a xor b);
    outputs(8403) <= not a or b;
    outputs(8404) <= b;
    outputs(8405) <= a and b;
    outputs(8406) <= a or b;
    outputs(8407) <= not (a xor b);
    outputs(8408) <= not a or b;
    outputs(8409) <= b;
    outputs(8410) <= a xor b;
    outputs(8411) <= not a or b;
    outputs(8412) <= not (a or b);
    outputs(8413) <= a;
    outputs(8414) <= not (a or b);
    outputs(8415) <= not (a and b);
    outputs(8416) <= a xor b;
    outputs(8417) <= not (a xor b);
    outputs(8418) <= not (a and b);
    outputs(8419) <= not a;
    outputs(8420) <= a or b;
    outputs(8421) <= a xor b;
    outputs(8422) <= a and b;
    outputs(8423) <= a;
    outputs(8424) <= b;
    outputs(8425) <= not a;
    outputs(8426) <= not (a and b);
    outputs(8427) <= not b or a;
    outputs(8428) <= b;
    outputs(8429) <= not (a and b);
    outputs(8430) <= a and b;
    outputs(8431) <= not a;
    outputs(8432) <= not a or b;
    outputs(8433) <= not (a xor b);
    outputs(8434) <= a xor b;
    outputs(8435) <= b;
    outputs(8436) <= b and not a;
    outputs(8437) <= not (a xor b);
    outputs(8438) <= not a or b;
    outputs(8439) <= b and not a;
    outputs(8440) <= not (a xor b);
    outputs(8441) <= not a;
    outputs(8442) <= not b;
    outputs(8443) <= not (a xor b);
    outputs(8444) <= not (a xor b);
    outputs(8445) <= a;
    outputs(8446) <= a;
    outputs(8447) <= b and not a;
    outputs(8448) <= not (a and b);
    outputs(8449) <= not (a xor b);
    outputs(8450) <= not (a and b);
    outputs(8451) <= not (a or b);
    outputs(8452) <= not a;
    outputs(8453) <= a xor b;
    outputs(8454) <= not a or b;
    outputs(8455) <= b and not a;
    outputs(8456) <= not a;
    outputs(8457) <= not (a xor b);
    outputs(8458) <= a xor b;
    outputs(8459) <= not (a xor b);
    outputs(8460) <= b;
    outputs(8461) <= not b;
    outputs(8462) <= not (a and b);
    outputs(8463) <= a xor b;
    outputs(8464) <= not (a xor b);
    outputs(8465) <= not (a xor b);
    outputs(8466) <= not (a xor b);
    outputs(8467) <= not (a or b);
    outputs(8468) <= not a;
    outputs(8469) <= not b;
    outputs(8470) <= not (a or b);
    outputs(8471) <= not b;
    outputs(8472) <= not b;
    outputs(8473) <= not (a and b);
    outputs(8474) <= a and not b;
    outputs(8475) <= a xor b;
    outputs(8476) <= a;
    outputs(8477) <= not (a or b);
    outputs(8478) <= not (a and b);
    outputs(8479) <= not a or b;
    outputs(8480) <= not (a or b);
    outputs(8481) <= not (a and b);
    outputs(8482) <= not a;
    outputs(8483) <= a;
    outputs(8484) <= not a or b;
    outputs(8485) <= not (a and b);
    outputs(8486) <= not (a or b);
    outputs(8487) <= b;
    outputs(8488) <= not (a xor b);
    outputs(8489) <= a;
    outputs(8490) <= not b;
    outputs(8491) <= a;
    outputs(8492) <= b and not a;
    outputs(8493) <= b;
    outputs(8494) <= not (a xor b);
    outputs(8495) <= not b;
    outputs(8496) <= b and not a;
    outputs(8497) <= not a or b;
    outputs(8498) <= a xor b;
    outputs(8499) <= not (a xor b);
    outputs(8500) <= a xor b;
    outputs(8501) <= not (a xor b);
    outputs(8502) <= a and b;
    outputs(8503) <= b and not a;
    outputs(8504) <= a;
    outputs(8505) <= a and not b;
    outputs(8506) <= b;
    outputs(8507) <= not b;
    outputs(8508) <= not (a xor b);
    outputs(8509) <= a and b;
    outputs(8510) <= a or b;
    outputs(8511) <= b;
    outputs(8512) <= b;
    outputs(8513) <= a xor b;
    outputs(8514) <= not a;
    outputs(8515) <= not (a and b);
    outputs(8516) <= a;
    outputs(8517) <= a;
    outputs(8518) <= a xor b;
    outputs(8519) <= not (a xor b);
    outputs(8520) <= not (a and b);
    outputs(8521) <= not b or a;
    outputs(8522) <= not (a xor b);
    outputs(8523) <= not a;
    outputs(8524) <= not b;
    outputs(8525) <= a and not b;
    outputs(8526) <= not a;
    outputs(8527) <= a xor b;
    outputs(8528) <= b;
    outputs(8529) <= not a or b;
    outputs(8530) <= b;
    outputs(8531) <= not (a and b);
    outputs(8532) <= b;
    outputs(8533) <= a or b;
    outputs(8534) <= not b or a;
    outputs(8535) <= not a;
    outputs(8536) <= not (a xor b);
    outputs(8537) <= b and not a;
    outputs(8538) <= a xor b;
    outputs(8539) <= a xor b;
    outputs(8540) <= not b;
    outputs(8541) <= not a or b;
    outputs(8542) <= b;
    outputs(8543) <= a;
    outputs(8544) <= a xor b;
    outputs(8545) <= not a or b;
    outputs(8546) <= not b or a;
    outputs(8547) <= not b;
    outputs(8548) <= not b or a;
    outputs(8549) <= a;
    outputs(8550) <= a and b;
    outputs(8551) <= b;
    outputs(8552) <= not (a and b);
    outputs(8553) <= not a or b;
    outputs(8554) <= b;
    outputs(8555) <= a xor b;
    outputs(8556) <= a and b;
    outputs(8557) <= not (a xor b);
    outputs(8558) <= not (a xor b);
    outputs(8559) <= not a or b;
    outputs(8560) <= a or b;
    outputs(8561) <= not a;
    outputs(8562) <= b and not a;
    outputs(8563) <= a xor b;
    outputs(8564) <= b;
    outputs(8565) <= b and not a;
    outputs(8566) <= b;
    outputs(8567) <= not b;
    outputs(8568) <= a xor b;
    outputs(8569) <= not (a xor b);
    outputs(8570) <= a or b;
    outputs(8571) <= b;
    outputs(8572) <= not (a and b);
    outputs(8573) <= not a;
    outputs(8574) <= not (a xor b);
    outputs(8575) <= a or b;
    outputs(8576) <= not a;
    outputs(8577) <= a;
    outputs(8578) <= a;
    outputs(8579) <= a;
    outputs(8580) <= not b;
    outputs(8581) <= not a or b;
    outputs(8582) <= not a;
    outputs(8583) <= not (a and b);
    outputs(8584) <= not a;
    outputs(8585) <= b and not a;
    outputs(8586) <= a;
    outputs(8587) <= a;
    outputs(8588) <= not a;
    outputs(8589) <= a xor b;
    outputs(8590) <= not (a xor b);
    outputs(8591) <= not a or b;
    outputs(8592) <= a;
    outputs(8593) <= a;
    outputs(8594) <= not b;
    outputs(8595) <= not (a and b);
    outputs(8596) <= not (a and b);
    outputs(8597) <= b;
    outputs(8598) <= a xor b;
    outputs(8599) <= not b or a;
    outputs(8600) <= not (a and b);
    outputs(8601) <= a xor b;
    outputs(8602) <= not a or b;
    outputs(8603) <= a;
    outputs(8604) <= b;
    outputs(8605) <= not b or a;
    outputs(8606) <= not (a and b);
    outputs(8607) <= not (a xor b);
    outputs(8608) <= not b;
    outputs(8609) <= not (a xor b);
    outputs(8610) <= not a;
    outputs(8611) <= not (a xor b);
    outputs(8612) <= not a or b;
    outputs(8613) <= not b;
    outputs(8614) <= a;
    outputs(8615) <= a;
    outputs(8616) <= a;
    outputs(8617) <= not b or a;
    outputs(8618) <= a;
    outputs(8619) <= a xor b;
    outputs(8620) <= a xor b;
    outputs(8621) <= a;
    outputs(8622) <= not b;
    outputs(8623) <= a;
    outputs(8624) <= not a;
    outputs(8625) <= not b or a;
    outputs(8626) <= a and not b;
    outputs(8627) <= not (a and b);
    outputs(8628) <= not (a xor b);
    outputs(8629) <= not a or b;
    outputs(8630) <= not b or a;
    outputs(8631) <= not (a xor b);
    outputs(8632) <= not (a xor b);
    outputs(8633) <= a xor b;
    outputs(8634) <= not a;
    outputs(8635) <= a;
    outputs(8636) <= b and not a;
    outputs(8637) <= a xor b;
    outputs(8638) <= not a;
    outputs(8639) <= a xor b;
    outputs(8640) <= not (a xor b);
    outputs(8641) <= not (a or b);
    outputs(8642) <= a xor b;
    outputs(8643) <= not (a and b);
    outputs(8644) <= a xor b;
    outputs(8645) <= a xor b;
    outputs(8646) <= not (a and b);
    outputs(8647) <= not b;
    outputs(8648) <= a and not b;
    outputs(8649) <= not (a xor b);
    outputs(8650) <= not b;
    outputs(8651) <= not (a or b);
    outputs(8652) <= a and not b;
    outputs(8653) <= b;
    outputs(8654) <= a xor b;
    outputs(8655) <= a and not b;
    outputs(8656) <= not (a and b);
    outputs(8657) <= not b;
    outputs(8658) <= a xor b;
    outputs(8659) <= a xor b;
    outputs(8660) <= not a;
    outputs(8661) <= not b;
    outputs(8662) <= not b or a;
    outputs(8663) <= a;
    outputs(8664) <= not b;
    outputs(8665) <= not (a xor b);
    outputs(8666) <= not b;
    outputs(8667) <= not b;
    outputs(8668) <= a;
    outputs(8669) <= not a or b;
    outputs(8670) <= b;
    outputs(8671) <= a and b;
    outputs(8672) <= b;
    outputs(8673) <= not (a and b);
    outputs(8674) <= a;
    outputs(8675) <= not b;
    outputs(8676) <= not (a or b);
    outputs(8677) <= not (a and b);
    outputs(8678) <= not (a and b);
    outputs(8679) <= a xor b;
    outputs(8680) <= a or b;
    outputs(8681) <= b;
    outputs(8682) <= not (a and b);
    outputs(8683) <= not (a xor b);
    outputs(8684) <= b;
    outputs(8685) <= a or b;
    outputs(8686) <= a and not b;
    outputs(8687) <= a xor b;
    outputs(8688) <= not (a xor b);
    outputs(8689) <= a xor b;
    outputs(8690) <= not a;
    outputs(8691) <= not (a and b);
    outputs(8692) <= not b;
    outputs(8693) <= not b or a;
    outputs(8694) <= a xor b;
    outputs(8695) <= a xor b;
    outputs(8696) <= a and not b;
    outputs(8697) <= a xor b;
    outputs(8698) <= not (a xor b);
    outputs(8699) <= not (a xor b);
    outputs(8700) <= b and not a;
    outputs(8701) <= a xor b;
    outputs(8702) <= a xor b;
    outputs(8703) <= not (a xor b);
    outputs(8704) <= not (a xor b);
    outputs(8705) <= not a;
    outputs(8706) <= not b;
    outputs(8707) <= not a;
    outputs(8708) <= b;
    outputs(8709) <= b;
    outputs(8710) <= not a;
    outputs(8711) <= not (a and b);
    outputs(8712) <= not (a xor b);
    outputs(8713) <= a or b;
    outputs(8714) <= not (a xor b);
    outputs(8715) <= a xor b;
    outputs(8716) <= not a;
    outputs(8717) <= not a or b;
    outputs(8718) <= a and not b;
    outputs(8719) <= not a or b;
    outputs(8720) <= not (a or b);
    outputs(8721) <= not a;
    outputs(8722) <= not a;
    outputs(8723) <= b;
    outputs(8724) <= b;
    outputs(8725) <= a xor b;
    outputs(8726) <= not (a xor b);
    outputs(8727) <= not (a or b);
    outputs(8728) <= a xor b;
    outputs(8729) <= not a or b;
    outputs(8730) <= not b or a;
    outputs(8731) <= a xor b;
    outputs(8732) <= not b;
    outputs(8733) <= not a;
    outputs(8734) <= not (a xor b);
    outputs(8735) <= b;
    outputs(8736) <= not (a and b);
    outputs(8737) <= not (a and b);
    outputs(8738) <= a;
    outputs(8739) <= not b;
    outputs(8740) <= a xor b;
    outputs(8741) <= b;
    outputs(8742) <= not b;
    outputs(8743) <= not (a xor b);
    outputs(8744) <= not (a xor b);
    outputs(8745) <= not a or b;
    outputs(8746) <= a xor b;
    outputs(8747) <= not b;
    outputs(8748) <= a and not b;
    outputs(8749) <= a;
    outputs(8750) <= a and not b;
    outputs(8751) <= a xor b;
    outputs(8752) <= a and b;
    outputs(8753) <= not (a or b);
    outputs(8754) <= not b or a;
    outputs(8755) <= not a;
    outputs(8756) <= not (a and b);
    outputs(8757) <= not a;
    outputs(8758) <= not (a xor b);
    outputs(8759) <= not (a and b);
    outputs(8760) <= not (a xor b);
    outputs(8761) <= not (a xor b);
    outputs(8762) <= b;
    outputs(8763) <= not (a xor b);
    outputs(8764) <= not a;
    outputs(8765) <= a;
    outputs(8766) <= a and b;
    outputs(8767) <= not (a xor b);
    outputs(8768) <= a;
    outputs(8769) <= not a;
    outputs(8770) <= not b or a;
    outputs(8771) <= not a;
    outputs(8772) <= not (a or b);
    outputs(8773) <= not a;
    outputs(8774) <= not a;
    outputs(8775) <= not b;
    outputs(8776) <= a;
    outputs(8777) <= not (a xor b);
    outputs(8778) <= not b;
    outputs(8779) <= not a or b;
    outputs(8780) <= not (a xor b);
    outputs(8781) <= b;
    outputs(8782) <= a xor b;
    outputs(8783) <= not (a xor b);
    outputs(8784) <= a;
    outputs(8785) <= not (a xor b);
    outputs(8786) <= a xor b;
    outputs(8787) <= not (a and b);
    outputs(8788) <= not a or b;
    outputs(8789) <= not a or b;
    outputs(8790) <= a xor b;
    outputs(8791) <= a and not b;
    outputs(8792) <= a xor b;
    outputs(8793) <= b;
    outputs(8794) <= not (a xor b);
    outputs(8795) <= not a;
    outputs(8796) <= b and not a;
    outputs(8797) <= a xor b;
    outputs(8798) <= not (a xor b);
    outputs(8799) <= a or b;
    outputs(8800) <= not a;
    outputs(8801) <= not a or b;
    outputs(8802) <= a or b;
    outputs(8803) <= a;
    outputs(8804) <= a xor b;
    outputs(8805) <= not a or b;
    outputs(8806) <= not (a or b);
    outputs(8807) <= a;
    outputs(8808) <= not a or b;
    outputs(8809) <= not a;
    outputs(8810) <= a xor b;
    outputs(8811) <= a;
    outputs(8812) <= not b;
    outputs(8813) <= not (a xor b);
    outputs(8814) <= not b;
    outputs(8815) <= not a;
    outputs(8816) <= a and not b;
    outputs(8817) <= a and not b;
    outputs(8818) <= a xor b;
    outputs(8819) <= not a;
    outputs(8820) <= not a;
    outputs(8821) <= a xor b;
    outputs(8822) <= b;
    outputs(8823) <= b;
    outputs(8824) <= a xor b;
    outputs(8825) <= b;
    outputs(8826) <= a and b;
    outputs(8827) <= not a;
    outputs(8828) <= a or b;
    outputs(8829) <= a xor b;
    outputs(8830) <= a xor b;
    outputs(8831) <= a;
    outputs(8832) <= not (a and b);
    outputs(8833) <= a xor b;
    outputs(8834) <= a or b;
    outputs(8835) <= not (a xor b);
    outputs(8836) <= not (a xor b);
    outputs(8837) <= not a;
    outputs(8838) <= not b or a;
    outputs(8839) <= not (a xor b);
    outputs(8840) <= not a or b;
    outputs(8841) <= a xor b;
    outputs(8842) <= a xor b;
    outputs(8843) <= b and not a;
    outputs(8844) <= not (a and b);
    outputs(8845) <= a xor b;
    outputs(8846) <= a xor b;
    outputs(8847) <= not (a xor b);
    outputs(8848) <= not (a xor b);
    outputs(8849) <= a and b;
    outputs(8850) <= a and b;
    outputs(8851) <= a or b;
    outputs(8852) <= a or b;
    outputs(8853) <= not (a xor b);
    outputs(8854) <= a xor b;
    outputs(8855) <= not a;
    outputs(8856) <= not (a xor b);
    outputs(8857) <= not a or b;
    outputs(8858) <= a;
    outputs(8859) <= b and not a;
    outputs(8860) <= b and not a;
    outputs(8861) <= a xor b;
    outputs(8862) <= b;
    outputs(8863) <= a xor b;
    outputs(8864) <= b and not a;
    outputs(8865) <= not a or b;
    outputs(8866) <= b and not a;
    outputs(8867) <= a;
    outputs(8868) <= not b;
    outputs(8869) <= not b;
    outputs(8870) <= a;
    outputs(8871) <= b;
    outputs(8872) <= not (a xor b);
    outputs(8873) <= not (a xor b);
    outputs(8874) <= b;
    outputs(8875) <= not b or a;
    outputs(8876) <= a;
    outputs(8877) <= not (a xor b);
    outputs(8878) <= not (a or b);
    outputs(8879) <= not (a xor b);
    outputs(8880) <= not (a xor b);
    outputs(8881) <= b and not a;
    outputs(8882) <= a and not b;
    outputs(8883) <= b;
    outputs(8884) <= not b;
    outputs(8885) <= b;
    outputs(8886) <= b;
    outputs(8887) <= not (a xor b);
    outputs(8888) <= not (a xor b);
    outputs(8889) <= not a;
    outputs(8890) <= a;
    outputs(8891) <= a xor b;
    outputs(8892) <= not b;
    outputs(8893) <= a xor b;
    outputs(8894) <= not (a xor b);
    outputs(8895) <= a;
    outputs(8896) <= a xor b;
    outputs(8897) <= a;
    outputs(8898) <= a or b;
    outputs(8899) <= not (a xor b);
    outputs(8900) <= not b or a;
    outputs(8901) <= a and not b;
    outputs(8902) <= a xor b;
    outputs(8903) <= a;
    outputs(8904) <= a xor b;
    outputs(8905) <= not a;
    outputs(8906) <= not (a xor b);
    outputs(8907) <= a xor b;
    outputs(8908) <= a and not b;
    outputs(8909) <= not a or b;
    outputs(8910) <= not (a and b);
    outputs(8911) <= a xor b;
    outputs(8912) <= not (a xor b);
    outputs(8913) <= not b;
    outputs(8914) <= not b or a;
    outputs(8915) <= a xor b;
    outputs(8916) <= a and b;
    outputs(8917) <= not a or b;
    outputs(8918) <= b;
    outputs(8919) <= not a;
    outputs(8920) <= b and not a;
    outputs(8921) <= a;
    outputs(8922) <= not a;
    outputs(8923) <= not (a xor b);
    outputs(8924) <= not (a xor b);
    outputs(8925) <= a xor b;
    outputs(8926) <= not (a xor b);
    outputs(8927) <= not b;
    outputs(8928) <= a xor b;
    outputs(8929) <= not (a xor b);
    outputs(8930) <= not a or b;
    outputs(8931) <= a xor b;
    outputs(8932) <= not (a xor b);
    outputs(8933) <= not (a xor b);
    outputs(8934) <= not b or a;
    outputs(8935) <= not (a or b);
    outputs(8936) <= not (a xor b);
    outputs(8937) <= a;
    outputs(8938) <= not a;
    outputs(8939) <= b;
    outputs(8940) <= not (a xor b);
    outputs(8941) <= not (a and b);
    outputs(8942) <= not a;
    outputs(8943) <= not (a xor b);
    outputs(8944) <= not b or a;
    outputs(8945) <= not b;
    outputs(8946) <= not (a xor b);
    outputs(8947) <= not b;
    outputs(8948) <= not a or b;
    outputs(8949) <= not (a xor b);
    outputs(8950) <= a;
    outputs(8951) <= not (a and b);
    outputs(8952) <= not a or b;
    outputs(8953) <= not (a or b);
    outputs(8954) <= not (a xor b);
    outputs(8955) <= a or b;
    outputs(8956) <= b and not a;
    outputs(8957) <= b;
    outputs(8958) <= not b or a;
    outputs(8959) <= not b or a;
    outputs(8960) <= not (a and b);
    outputs(8961) <= not (a xor b);
    outputs(8962) <= a and b;
    outputs(8963) <= a xor b;
    outputs(8964) <= not (a and b);
    outputs(8965) <= not b;
    outputs(8966) <= not b;
    outputs(8967) <= not b;
    outputs(8968) <= a;
    outputs(8969) <= not b;
    outputs(8970) <= a;
    outputs(8971) <= not a;
    outputs(8972) <= not (a and b);
    outputs(8973) <= a;
    outputs(8974) <= not a;
    outputs(8975) <= a xor b;
    outputs(8976) <= not (a xor b);
    outputs(8977) <= a xor b;
    outputs(8978) <= a xor b;
    outputs(8979) <= a xor b;
    outputs(8980) <= not (a xor b);
    outputs(8981) <= a xor b;
    outputs(8982) <= b;
    outputs(8983) <= a;
    outputs(8984) <= b and not a;
    outputs(8985) <= not b;
    outputs(8986) <= not a;
    outputs(8987) <= not a;
    outputs(8988) <= not (a xor b);
    outputs(8989) <= a xor b;
    outputs(8990) <= not (a xor b);
    outputs(8991) <= not b;
    outputs(8992) <= not (a xor b);
    outputs(8993) <= b;
    outputs(8994) <= a or b;
    outputs(8995) <= not b;
    outputs(8996) <= b;
    outputs(8997) <= not (a xor b);
    outputs(8998) <= not (a xor b);
    outputs(8999) <= not (a or b);
    outputs(9000) <= not (a xor b);
    outputs(9001) <= not b;
    outputs(9002) <= not b;
    outputs(9003) <= a or b;
    outputs(9004) <= not (a and b);
    outputs(9005) <= a or b;
    outputs(9006) <= a and b;
    outputs(9007) <= not (a xor b);
    outputs(9008) <= b;
    outputs(9009) <= not a;
    outputs(9010) <= a xor b;
    outputs(9011) <= not b;
    outputs(9012) <= not a or b;
    outputs(9013) <= b;
    outputs(9014) <= not a;
    outputs(9015) <= b;
    outputs(9016) <= a or b;
    outputs(9017) <= not b or a;
    outputs(9018) <= a and not b;
    outputs(9019) <= a;
    outputs(9020) <= not (a and b);
    outputs(9021) <= a or b;
    outputs(9022) <= not (a and b);
    outputs(9023) <= a and not b;
    outputs(9024) <= a xor b;
    outputs(9025) <= a or b;
    outputs(9026) <= not b;
    outputs(9027) <= not (a xor b);
    outputs(9028) <= a and not b;
    outputs(9029) <= a xor b;
    outputs(9030) <= not (a xor b);
    outputs(9031) <= a;
    outputs(9032) <= not a;
    outputs(9033) <= a xor b;
    outputs(9034) <= a xor b;
    outputs(9035) <= not b;
    outputs(9036) <= a and b;
    outputs(9037) <= b and not a;
    outputs(9038) <= a;
    outputs(9039) <= a xor b;
    outputs(9040) <= not (a xor b);
    outputs(9041) <= not (a and b);
    outputs(9042) <= not (a xor b);
    outputs(9043) <= not b or a;
    outputs(9044) <= not a or b;
    outputs(9045) <= not b;
    outputs(9046) <= not b;
    outputs(9047) <= a xor b;
    outputs(9048) <= not (a xor b);
    outputs(9049) <= not b or a;
    outputs(9050) <= a and not b;
    outputs(9051) <= a xor b;
    outputs(9052) <= not (a xor b);
    outputs(9053) <= not b;
    outputs(9054) <= b;
    outputs(9055) <= b and not a;
    outputs(9056) <= a;
    outputs(9057) <= a;
    outputs(9058) <= a and not b;
    outputs(9059) <= a or b;
    outputs(9060) <= a xor b;
    outputs(9061) <= not (a and b);
    outputs(9062) <= a xor b;
    outputs(9063) <= b;
    outputs(9064) <= not (a or b);
    outputs(9065) <= not b;
    outputs(9066) <= b;
    outputs(9067) <= b and not a;
    outputs(9068) <= not (a and b);
    outputs(9069) <= a;
    outputs(9070) <= not a;
    outputs(9071) <= not (a xor b);
    outputs(9072) <= not (a xor b);
    outputs(9073) <= not (a or b);
    outputs(9074) <= a xor b;
    outputs(9075) <= not (a and b);
    outputs(9076) <= b and not a;
    outputs(9077) <= b;
    outputs(9078) <= a or b;
    outputs(9079) <= not (a or b);
    outputs(9080) <= a xor b;
    outputs(9081) <= a xor b;
    outputs(9082) <= a xor b;
    outputs(9083) <= a xor b;
    outputs(9084) <= b and not a;
    outputs(9085) <= not (a and b);
    outputs(9086) <= a and not b;
    outputs(9087) <= a;
    outputs(9088) <= a and b;
    outputs(9089) <= b;
    outputs(9090) <= a xor b;
    outputs(9091) <= a xor b;
    outputs(9092) <= not (a xor b);
    outputs(9093) <= not (a xor b);
    outputs(9094) <= a xor b;
    outputs(9095) <= a and b;
    outputs(9096) <= a and not b;
    outputs(9097) <= not b;
    outputs(9098) <= not (a or b);
    outputs(9099) <= a or b;
    outputs(9100) <= not (a xor b);
    outputs(9101) <= not b or a;
    outputs(9102) <= a or b;
    outputs(9103) <= not (a xor b);
    outputs(9104) <= a or b;
    outputs(9105) <= not b;
    outputs(9106) <= b;
    outputs(9107) <= not (a xor b);
    outputs(9108) <= not b;
    outputs(9109) <= not (a xor b);
    outputs(9110) <= b;
    outputs(9111) <= b and not a;
    outputs(9112) <= not a;
    outputs(9113) <= not (a xor b);
    outputs(9114) <= a and b;
    outputs(9115) <= not a;
    outputs(9116) <= b;
    outputs(9117) <= b;
    outputs(9118) <= a;
    outputs(9119) <= b and not a;
    outputs(9120) <= not b or a;
    outputs(9121) <= b and not a;
    outputs(9122) <= b;
    outputs(9123) <= a xor b;
    outputs(9124) <= a;
    outputs(9125) <= a and b;
    outputs(9126) <= a and b;
    outputs(9127) <= not (a xor b);
    outputs(9128) <= b;
    outputs(9129) <= a xor b;
    outputs(9130) <= b;
    outputs(9131) <= b;
    outputs(9132) <= a xor b;
    outputs(9133) <= a xor b;
    outputs(9134) <= not a;
    outputs(9135) <= not a;
    outputs(9136) <= not (a xor b);
    outputs(9137) <= a and b;
    outputs(9138) <= b;
    outputs(9139) <= a xor b;
    outputs(9140) <= not a;
    outputs(9141) <= a and not b;
    outputs(9142) <= a xor b;
    outputs(9143) <= not b;
    outputs(9144) <= not a;
    outputs(9145) <= not (a xor b);
    outputs(9146) <= b;
    outputs(9147) <= not b;
    outputs(9148) <= a or b;
    outputs(9149) <= not (a or b);
    outputs(9150) <= a;
    outputs(9151) <= a or b;
    outputs(9152) <= not (a and b);
    outputs(9153) <= not (a xor b);
    outputs(9154) <= not (a or b);
    outputs(9155) <= a;
    outputs(9156) <= a xor b;
    outputs(9157) <= not a;
    outputs(9158) <= not b or a;
    outputs(9159) <= not b or a;
    outputs(9160) <= a xor b;
    outputs(9161) <= not a;
    outputs(9162) <= a;
    outputs(9163) <= a or b;
    outputs(9164) <= not (a xor b);
    outputs(9165) <= a xor b;
    outputs(9166) <= not (a and b);
    outputs(9167) <= not (a xor b);
    outputs(9168) <= not a;
    outputs(9169) <= a;
    outputs(9170) <= not b;
    outputs(9171) <= a;
    outputs(9172) <= not b;
    outputs(9173) <= a or b;
    outputs(9174) <= b;
    outputs(9175) <= not a or b;
    outputs(9176) <= a and b;
    outputs(9177) <= a or b;
    outputs(9178) <= not (a xor b);
    outputs(9179) <= a;
    outputs(9180) <= not (a and b);
    outputs(9181) <= not a;
    outputs(9182) <= not a;
    outputs(9183) <= a xor b;
    outputs(9184) <= a or b;
    outputs(9185) <= a xor b;
    outputs(9186) <= not a or b;
    outputs(9187) <= b and not a;
    outputs(9188) <= not b or a;
    outputs(9189) <= a xor b;
    outputs(9190) <= a;
    outputs(9191) <= b and not a;
    outputs(9192) <= a xor b;
    outputs(9193) <= a or b;
    outputs(9194) <= not (a xor b);
    outputs(9195) <= b;
    outputs(9196) <= a;
    outputs(9197) <= b and not a;
    outputs(9198) <= a xor b;
    outputs(9199) <= a;
    outputs(9200) <= a and not b;
    outputs(9201) <= not b;
    outputs(9202) <= not a;
    outputs(9203) <= not b or a;
    outputs(9204) <= not (a xor b);
    outputs(9205) <= b and not a;
    outputs(9206) <= a and b;
    outputs(9207) <= a xor b;
    outputs(9208) <= a xor b;
    outputs(9209) <= not (a xor b);
    outputs(9210) <= b;
    outputs(9211) <= b;
    outputs(9212) <= b;
    outputs(9213) <= not a or b;
    outputs(9214) <= a xor b;
    outputs(9215) <= not (a and b);
    outputs(9216) <= b;
    outputs(9217) <= not b;
    outputs(9218) <= not (a or b);
    outputs(9219) <= not (a and b);
    outputs(9220) <= a;
    outputs(9221) <= a xor b;
    outputs(9222) <= not (a or b);
    outputs(9223) <= a and not b;
    outputs(9224) <= a xor b;
    outputs(9225) <= b;
    outputs(9226) <= a xor b;
    outputs(9227) <= not b;
    outputs(9228) <= not (a or b);
    outputs(9229) <= a xor b;
    outputs(9230) <= b and not a;
    outputs(9231) <= not (a and b);
    outputs(9232) <= a xor b;
    outputs(9233) <= not (a xor b);
    outputs(9234) <= a and b;
    outputs(9235) <= a and b;
    outputs(9236) <= not (a xor b);
    outputs(9237) <= a and not b;
    outputs(9238) <= not (a or b);
    outputs(9239) <= a or b;
    outputs(9240) <= not a;
    outputs(9241) <= a xor b;
    outputs(9242) <= b;
    outputs(9243) <= not a;
    outputs(9244) <= a xor b;
    outputs(9245) <= a and b;
    outputs(9246) <= not (a xor b);
    outputs(9247) <= not b;
    outputs(9248) <= a xor b;
    outputs(9249) <= a;
    outputs(9250) <= a;
    outputs(9251) <= a or b;
    outputs(9252) <= b;
    outputs(9253) <= not a;
    outputs(9254) <= not (a xor b);
    outputs(9255) <= a;
    outputs(9256) <= not b;
    outputs(9257) <= a xor b;
    outputs(9258) <= not a;
    outputs(9259) <= not a;
    outputs(9260) <= not (a or b);
    outputs(9261) <= b and not a;
    outputs(9262) <= a xor b;
    outputs(9263) <= a;
    outputs(9264) <= a xor b;
    outputs(9265) <= not b or a;
    outputs(9266) <= a and b;
    outputs(9267) <= b;
    outputs(9268) <= a or b;
    outputs(9269) <= a xor b;
    outputs(9270) <= a xor b;
    outputs(9271) <= b;
    outputs(9272) <= a xor b;
    outputs(9273) <= a;
    outputs(9274) <= not a;
    outputs(9275) <= b;
    outputs(9276) <= b;
    outputs(9277) <= a xor b;
    outputs(9278) <= not (a xor b);
    outputs(9279) <= not (a xor b);
    outputs(9280) <= a and b;
    outputs(9281) <= not b;
    outputs(9282) <= a;
    outputs(9283) <= a xor b;
    outputs(9284) <= a xor b;
    outputs(9285) <= not a;
    outputs(9286) <= not (a and b);
    outputs(9287) <= a xor b;
    outputs(9288) <= not (a xor b);
    outputs(9289) <= a xor b;
    outputs(9290) <= not b;
    outputs(9291) <= a xor b;
    outputs(9292) <= not a or b;
    outputs(9293) <= b;
    outputs(9294) <= not (a xor b);
    outputs(9295) <= not (a or b);
    outputs(9296) <= a xor b;
    outputs(9297) <= a or b;
    outputs(9298) <= a and b;
    outputs(9299) <= a and b;
    outputs(9300) <= b and not a;
    outputs(9301) <= not (a xor b);
    outputs(9302) <= b and not a;
    outputs(9303) <= b and not a;
    outputs(9304) <= a;
    outputs(9305) <= not a;
    outputs(9306) <= a xor b;
    outputs(9307) <= not (a xor b);
    outputs(9308) <= a and not b;
    outputs(9309) <= a xor b;
    outputs(9310) <= b;
    outputs(9311) <= a;
    outputs(9312) <= a;
    outputs(9313) <= a xor b;
    outputs(9314) <= not b;
    outputs(9315) <= a and b;
    outputs(9316) <= a or b;
    outputs(9317) <= b;
    outputs(9318) <= not (a xor b);
    outputs(9319) <= a and b;
    outputs(9320) <= a xor b;
    outputs(9321) <= b;
    outputs(9322) <= b;
    outputs(9323) <= a or b;
    outputs(9324) <= not a;
    outputs(9325) <= b and not a;
    outputs(9326) <= b and not a;
    outputs(9327) <= b and not a;
    outputs(9328) <= not (a xor b);
    outputs(9329) <= b and not a;
    outputs(9330) <= a and not b;
    outputs(9331) <= a and not b;
    outputs(9332) <= not (a xor b);
    outputs(9333) <= b;
    outputs(9334) <= not a or b;
    outputs(9335) <= b;
    outputs(9336) <= a xor b;
    outputs(9337) <= a xor b;
    outputs(9338) <= a and b;
    outputs(9339) <= not a;
    outputs(9340) <= a xor b;
    outputs(9341) <= not b;
    outputs(9342) <= not a;
    outputs(9343) <= not (a and b);
    outputs(9344) <= a or b;
    outputs(9345) <= not a;
    outputs(9346) <= b;
    outputs(9347) <= not (a xor b);
    outputs(9348) <= a and not b;
    outputs(9349) <= a xor b;
    outputs(9350) <= a;
    outputs(9351) <= not b;
    outputs(9352) <= b and not a;
    outputs(9353) <= not b;
    outputs(9354) <= not b or a;
    outputs(9355) <= not (a xor b);
    outputs(9356) <= not a;
    outputs(9357) <= not a or b;
    outputs(9358) <= b;
    outputs(9359) <= a and not b;
    outputs(9360) <= b;
    outputs(9361) <= not a;
    outputs(9362) <= b and not a;
    outputs(9363) <= not (a xor b);
    outputs(9364) <= not a;
    outputs(9365) <= a xor b;
    outputs(9366) <= not a;
    outputs(9367) <= b;
    outputs(9368) <= not a;
    outputs(9369) <= not b;
    outputs(9370) <= a;
    outputs(9371) <= a and b;
    outputs(9372) <= a and b;
    outputs(9373) <= a xor b;
    outputs(9374) <= not b;
    outputs(9375) <= not a;
    outputs(9376) <= b;
    outputs(9377) <= a xor b;
    outputs(9378) <= not a;
    outputs(9379) <= not b;
    outputs(9380) <= a;
    outputs(9381) <= b and not a;
    outputs(9382) <= a;
    outputs(9383) <= not b;
    outputs(9384) <= not (a xor b);
    outputs(9385) <= b;
    outputs(9386) <= a xor b;
    outputs(9387) <= a and b;
    outputs(9388) <= a xor b;
    outputs(9389) <= a xor b;
    outputs(9390) <= not b;
    outputs(9391) <= b;
    outputs(9392) <= not (a xor b);
    outputs(9393) <= not (a xor b);
    outputs(9394) <= not (a or b);
    outputs(9395) <= not b;
    outputs(9396) <= not a;
    outputs(9397) <= a and b;
    outputs(9398) <= a;
    outputs(9399) <= not (a or b);
    outputs(9400) <= a and not b;
    outputs(9401) <= not (a xor b);
    outputs(9402) <= b and not a;
    outputs(9403) <= a xor b;
    outputs(9404) <= not b or a;
    outputs(9405) <= b;
    outputs(9406) <= not (a xor b);
    outputs(9407) <= not (a xor b);
    outputs(9408) <= a;
    outputs(9409) <= a or b;
    outputs(9410) <= a xor b;
    outputs(9411) <= not a;
    outputs(9412) <= not b;
    outputs(9413) <= a xor b;
    outputs(9414) <= not b;
    outputs(9415) <= not a;
    outputs(9416) <= b and not a;
    outputs(9417) <= a or b;
    outputs(9418) <= b;
    outputs(9419) <= not a;
    outputs(9420) <= a;
    outputs(9421) <= not (a xor b);
    outputs(9422) <= a;
    outputs(9423) <= a xor b;
    outputs(9424) <= a and b;
    outputs(9425) <= not b;
    outputs(9426) <= not (a xor b);
    outputs(9427) <= a;
    outputs(9428) <= not b;
    outputs(9429) <= a and not b;
    outputs(9430) <= not (a and b);
    outputs(9431) <= not (a and b);
    outputs(9432) <= a;
    outputs(9433) <= a xor b;
    outputs(9434) <= a xor b;
    outputs(9435) <= a and b;
    outputs(9436) <= not (a xor b);
    outputs(9437) <= not a;
    outputs(9438) <= a xor b;
    outputs(9439) <= not (a xor b);
    outputs(9440) <= a xor b;
    outputs(9441) <= a;
    outputs(9442) <= not (a or b);
    outputs(9443) <= not a;
    outputs(9444) <= not (a xor b);
    outputs(9445) <= not b;
    outputs(9446) <= not (a xor b);
    outputs(9447) <= b;
    outputs(9448) <= not a;
    outputs(9449) <= b;
    outputs(9450) <= b;
    outputs(9451) <= not (a xor b);
    outputs(9452) <= a and not b;
    outputs(9453) <= not a;
    outputs(9454) <= b and not a;
    outputs(9455) <= a and not b;
    outputs(9456) <= a xor b;
    outputs(9457) <= not (a xor b);
    outputs(9458) <= b;
    outputs(9459) <= not (a or b);
    outputs(9460) <= not b;
    outputs(9461) <= a and b;
    outputs(9462) <= not (a xor b);
    outputs(9463) <= a;
    outputs(9464) <= a and not b;
    outputs(9465) <= not a;
    outputs(9466) <= b;
    outputs(9467) <= b;
    outputs(9468) <= not a;
    outputs(9469) <= not a;
    outputs(9470) <= not (a or b);
    outputs(9471) <= not b or a;
    outputs(9472) <= not a;
    outputs(9473) <= b;
    outputs(9474) <= not a or b;
    outputs(9475) <= a;
    outputs(9476) <= not b;
    outputs(9477) <= a or b;
    outputs(9478) <= a xor b;
    outputs(9479) <= a;
    outputs(9480) <= not a;
    outputs(9481) <= a xor b;
    outputs(9482) <= a xor b;
    outputs(9483) <= not (a and b);
    outputs(9484) <= not a;
    outputs(9485) <= a and b;
    outputs(9486) <= a;
    outputs(9487) <= not (a xor b);
    outputs(9488) <= not (a xor b);
    outputs(9489) <= a xor b;
    outputs(9490) <= not a;
    outputs(9491) <= not (a xor b);
    outputs(9492) <= a and not b;
    outputs(9493) <= b;
    outputs(9494) <= not (a xor b);
    outputs(9495) <= b and not a;
    outputs(9496) <= a xor b;
    outputs(9497) <= a and b;
    outputs(9498) <= not a;
    outputs(9499) <= not a;
    outputs(9500) <= a xor b;
    outputs(9501) <= b;
    outputs(9502) <= a;
    outputs(9503) <= not a;
    outputs(9504) <= not a or b;
    outputs(9505) <= not (a xor b);
    outputs(9506) <= b;
    outputs(9507) <= b;
    outputs(9508) <= a or b;
    outputs(9509) <= a and not b;
    outputs(9510) <= a xor b;
    outputs(9511) <= a xor b;
    outputs(9512) <= not a;
    outputs(9513) <= not b or a;
    outputs(9514) <= not (a xor b);
    outputs(9515) <= a;
    outputs(9516) <= b;
    outputs(9517) <= not (a xor b);
    outputs(9518) <= not a or b;
    outputs(9519) <= not a;
    outputs(9520) <= a or b;
    outputs(9521) <= not (a xor b);
    outputs(9522) <= a;
    outputs(9523) <= not (a xor b);
    outputs(9524) <= not (a xor b);
    outputs(9525) <= b and not a;
    outputs(9526) <= not b or a;
    outputs(9527) <= b and not a;
    outputs(9528) <= not (a and b);
    outputs(9529) <= not b;
    outputs(9530) <= b;
    outputs(9531) <= not (a or b);
    outputs(9532) <= b and not a;
    outputs(9533) <= a xor b;
    outputs(9534) <= not b or a;
    outputs(9535) <= not (a xor b);
    outputs(9536) <= b;
    outputs(9537) <= not a;
    outputs(9538) <= a;
    outputs(9539) <= not (a xor b);
    outputs(9540) <= not (a xor b);
    outputs(9541) <= not (a or b);
    outputs(9542) <= not (a xor b);
    outputs(9543) <= not (a or b);
    outputs(9544) <= b and not a;
    outputs(9545) <= a xor b;
    outputs(9546) <= not (a xor b);
    outputs(9547) <= a;
    outputs(9548) <= b and not a;
    outputs(9549) <= not b;
    outputs(9550) <= not (a or b);
    outputs(9551) <= a xor b;
    outputs(9552) <= b;
    outputs(9553) <= a and b;
    outputs(9554) <= b;
    outputs(9555) <= not b;
    outputs(9556) <= a and not b;
    outputs(9557) <= not b;
    outputs(9558) <= a and b;
    outputs(9559) <= b;
    outputs(9560) <= not a;
    outputs(9561) <= not b;
    outputs(9562) <= a or b;
    outputs(9563) <= not (a xor b);
    outputs(9564) <= not b;
    outputs(9565) <= a;
    outputs(9566) <= a xor b;
    outputs(9567) <= a xor b;
    outputs(9568) <= not (a xor b);
    outputs(9569) <= a and not b;
    outputs(9570) <= b and not a;
    outputs(9571) <= a and b;
    outputs(9572) <= a xor b;
    outputs(9573) <= b;
    outputs(9574) <= not (a and b);
    outputs(9575) <= b;
    outputs(9576) <= not b;
    outputs(9577) <= not a;
    outputs(9578) <= b and not a;
    outputs(9579) <= not (a xor b);
    outputs(9580) <= not a;
    outputs(9581) <= not (a xor b);
    outputs(9582) <= b;
    outputs(9583) <= not (a xor b);
    outputs(9584) <= not (a xor b);
    outputs(9585) <= a xor b;
    outputs(9586) <= b;
    outputs(9587) <= a;
    outputs(9588) <= not (a xor b);
    outputs(9589) <= not (a xor b);
    outputs(9590) <= not (a xor b);
    outputs(9591) <= a and not b;
    outputs(9592) <= a;
    outputs(9593) <= not b or a;
    outputs(9594) <= a;
    outputs(9595) <= b and not a;
    outputs(9596) <= not (a xor b);
    outputs(9597) <= not a;
    outputs(9598) <= not a or b;
    outputs(9599) <= not (a xor b);
    outputs(9600) <= not b;
    outputs(9601) <= not (a or b);
    outputs(9602) <= not b;
    outputs(9603) <= a;
    outputs(9604) <= not (a xor b);
    outputs(9605) <= a;
    outputs(9606) <= a and b;
    outputs(9607) <= a or b;
    outputs(9608) <= not (a xor b);
    outputs(9609) <= a and b;
    outputs(9610) <= not (a xor b);
    outputs(9611) <= a and b;
    outputs(9612) <= a xor b;
    outputs(9613) <= a xor b;
    outputs(9614) <= a xor b;
    outputs(9615) <= not b;
    outputs(9616) <= a xor b;
    outputs(9617) <= b;
    outputs(9618) <= b;
    outputs(9619) <= a;
    outputs(9620) <= not b;
    outputs(9621) <= not a or b;
    outputs(9622) <= not a;
    outputs(9623) <= b and not a;
    outputs(9624) <= b and not a;
    outputs(9625) <= not (a xor b);
    outputs(9626) <= not b;
    outputs(9627) <= a and b;
    outputs(9628) <= not b;
    outputs(9629) <= not a;
    outputs(9630) <= b and not a;
    outputs(9631) <= not (a or b);
    outputs(9632) <= a xor b;
    outputs(9633) <= a;
    outputs(9634) <= not (a xor b);
    outputs(9635) <= b and not a;
    outputs(9636) <= not (a xor b);
    outputs(9637) <= not (a xor b);
    outputs(9638) <= not (a xor b);
    outputs(9639) <= a xor b;
    outputs(9640) <= not (a xor b);
    outputs(9641) <= b and not a;
    outputs(9642) <= b;
    outputs(9643) <= b and not a;
    outputs(9644) <= not a;
    outputs(9645) <= a;
    outputs(9646) <= not b;
    outputs(9647) <= a;
    outputs(9648) <= a;
    outputs(9649) <= a and b;
    outputs(9650) <= a;
    outputs(9651) <= a xor b;
    outputs(9652) <= b;
    outputs(9653) <= not (a xor b);
    outputs(9654) <= b;
    outputs(9655) <= not b or a;
    outputs(9656) <= not a;
    outputs(9657) <= not (a xor b);
    outputs(9658) <= a;
    outputs(9659) <= not (a xor b);
    outputs(9660) <= a;
    outputs(9661) <= not b;
    outputs(9662) <= not a;
    outputs(9663) <= b;
    outputs(9664) <= not b;
    outputs(9665) <= a xor b;
    outputs(9666) <= b;
    outputs(9667) <= a and not b;
    outputs(9668) <= a;
    outputs(9669) <= not (a xor b);
    outputs(9670) <= b;
    outputs(9671) <= a and not b;
    outputs(9672) <= not (a or b);
    outputs(9673) <= not (a or b);
    outputs(9674) <= a;
    outputs(9675) <= b;
    outputs(9676) <= a and b;
    outputs(9677) <= b and not a;
    outputs(9678) <= a xor b;
    outputs(9679) <= b and not a;
    outputs(9680) <= not (a xor b);
    outputs(9681) <= not (a xor b);
    outputs(9682) <= a;
    outputs(9683) <= a and b;
    outputs(9684) <= not a;
    outputs(9685) <= a;
    outputs(9686) <= not a or b;
    outputs(9687) <= a and not b;
    outputs(9688) <= a xor b;
    outputs(9689) <= not (a xor b);
    outputs(9690) <= not b;
    outputs(9691) <= not (a xor b);
    outputs(9692) <= b and not a;
    outputs(9693) <= b and not a;
    outputs(9694) <= a and b;
    outputs(9695) <= not (a xor b);
    outputs(9696) <= not a;
    outputs(9697) <= b;
    outputs(9698) <= b and not a;
    outputs(9699) <= a and b;
    outputs(9700) <= a and b;
    outputs(9701) <= not (a xor b);
    outputs(9702) <= a xor b;
    outputs(9703) <= a and not b;
    outputs(9704) <= not (a xor b);
    outputs(9705) <= not a;
    outputs(9706) <= a and not b;
    outputs(9707) <= not b;
    outputs(9708) <= a xor b;
    outputs(9709) <= b;
    outputs(9710) <= not (a or b);
    outputs(9711) <= b;
    outputs(9712) <= b;
    outputs(9713) <= a xor b;
    outputs(9714) <= not b;
    outputs(9715) <= not b;
    outputs(9716) <= a and b;
    outputs(9717) <= b and not a;
    outputs(9718) <= b;
    outputs(9719) <= a xor b;
    outputs(9720) <= b;
    outputs(9721) <= not (a and b);
    outputs(9722) <= b and not a;
    outputs(9723) <= a xor b;
    outputs(9724) <= a or b;
    outputs(9725) <= b and not a;
    outputs(9726) <= a and not b;
    outputs(9727) <= not (a xor b);
    outputs(9728) <= a;
    outputs(9729) <= not a;
    outputs(9730) <= not (a or b);
    outputs(9731) <= a xor b;
    outputs(9732) <= not (a xor b);
    outputs(9733) <= a and not b;
    outputs(9734) <= not (a xor b);
    outputs(9735) <= not (a or b);
    outputs(9736) <= a xor b;
    outputs(9737) <= a or b;
    outputs(9738) <= not b;
    outputs(9739) <= not (a or b);
    outputs(9740) <= a or b;
    outputs(9741) <= a xor b;
    outputs(9742) <= a and b;
    outputs(9743) <= not (a xor b);
    outputs(9744) <= b and not a;
    outputs(9745) <= b and not a;
    outputs(9746) <= not (a or b);
    outputs(9747) <= not a;
    outputs(9748) <= not (a xor b);
    outputs(9749) <= b;
    outputs(9750) <= not a;
    outputs(9751) <= not a;
    outputs(9752) <= not (a and b);
    outputs(9753) <= not b or a;
    outputs(9754) <= not a;
    outputs(9755) <= a xor b;
    outputs(9756) <= a xor b;
    outputs(9757) <= not b;
    outputs(9758) <= a xor b;
    outputs(9759) <= not (a and b);
    outputs(9760) <= not a or b;
    outputs(9761) <= a;
    outputs(9762) <= not (a xor b);
    outputs(9763) <= a and not b;
    outputs(9764) <= a and not b;
    outputs(9765) <= a;
    outputs(9766) <= b and not a;
    outputs(9767) <= a and not b;
    outputs(9768) <= not (a xor b);
    outputs(9769) <= not a;
    outputs(9770) <= not a or b;
    outputs(9771) <= not (a xor b);
    outputs(9772) <= b and not a;
    outputs(9773) <= a xor b;
    outputs(9774) <= not (a xor b);
    outputs(9775) <= a and b;
    outputs(9776) <= b;
    outputs(9777) <= a xor b;
    outputs(9778) <= not a;
    outputs(9779) <= not a or b;
    outputs(9780) <= not b or a;
    outputs(9781) <= a;
    outputs(9782) <= not (a and b);
    outputs(9783) <= a xor b;
    outputs(9784) <= a xor b;
    outputs(9785) <= not (a or b);
    outputs(9786) <= a xor b;
    outputs(9787) <= not (a xor b);
    outputs(9788) <= not (a or b);
    outputs(9789) <= a and not b;
    outputs(9790) <= not (a xor b);
    outputs(9791) <= not (a xor b);
    outputs(9792) <= b and not a;
    outputs(9793) <= a xor b;
    outputs(9794) <= not b;
    outputs(9795) <= not (a or b);
    outputs(9796) <= b;
    outputs(9797) <= not b;
    outputs(9798) <= a and b;
    outputs(9799) <= not b;
    outputs(9800) <= a;
    outputs(9801) <= a xor b;
    outputs(9802) <= not a;
    outputs(9803) <= not a or b;
    outputs(9804) <= a;
    outputs(9805) <= b and not a;
    outputs(9806) <= a xor b;
    outputs(9807) <= a xor b;
    outputs(9808) <= a and b;
    outputs(9809) <= b and not a;
    outputs(9810) <= not (a or b);
    outputs(9811) <= not (a xor b);
    outputs(9812) <= a xor b;
    outputs(9813) <= not (a xor b);
    outputs(9814) <= not (a or b);
    outputs(9815) <= not (a xor b);
    outputs(9816) <= not a;
    outputs(9817) <= a and b;
    outputs(9818) <= b;
    outputs(9819) <= not (a or b);
    outputs(9820) <= b;
    outputs(9821) <= not a;
    outputs(9822) <= not (a xor b);
    outputs(9823) <= not b;
    outputs(9824) <= not (a xor b);
    outputs(9825) <= not a;
    outputs(9826) <= not (a xor b);
    outputs(9827) <= a xor b;
    outputs(9828) <= b;
    outputs(9829) <= not a;
    outputs(9830) <= a and not b;
    outputs(9831) <= a;
    outputs(9832) <= a or b;
    outputs(9833) <= not (a xor b);
    outputs(9834) <= not a;
    outputs(9835) <= b;
    outputs(9836) <= b;
    outputs(9837) <= a or b;
    outputs(9838) <= not (a xor b);
    outputs(9839) <= not a;
    outputs(9840) <= not (a xor b);
    outputs(9841) <= not (a or b);
    outputs(9842) <= b;
    outputs(9843) <= a and not b;
    outputs(9844) <= not (a and b);
    outputs(9845) <= not a;
    outputs(9846) <= a and b;
    outputs(9847) <= b;
    outputs(9848) <= b and not a;
    outputs(9849) <= not b;
    outputs(9850) <= a xor b;
    outputs(9851) <= a and b;
    outputs(9852) <= not a or b;
    outputs(9853) <= not (a xor b);
    outputs(9854) <= a;
    outputs(9855) <= not a;
    outputs(9856) <= not a;
    outputs(9857) <= a;
    outputs(9858) <= a;
    outputs(9859) <= a and b;
    outputs(9860) <= a;
    outputs(9861) <= a xor b;
    outputs(9862) <= b;
    outputs(9863) <= not (a or b);
    outputs(9864) <= not b or a;
    outputs(9865) <= a or b;
    outputs(9866) <= not a;
    outputs(9867) <= not (a or b);
    outputs(9868) <= b;
    outputs(9869) <= not (a and b);
    outputs(9870) <= not a;
    outputs(9871) <= a and not b;
    outputs(9872) <= not a or b;
    outputs(9873) <= not (a xor b);
    outputs(9874) <= a and not b;
    outputs(9875) <= a;
    outputs(9876) <= not (a xor b);
    outputs(9877) <= not b;
    outputs(9878) <= not a or b;
    outputs(9879) <= not b;
    outputs(9880) <= a and b;
    outputs(9881) <= a and b;
    outputs(9882) <= a xor b;
    outputs(9883) <= not (a or b);
    outputs(9884) <= not (a or b);
    outputs(9885) <= not b;
    outputs(9886) <= not b;
    outputs(9887) <= b and not a;
    outputs(9888) <= b and not a;
    outputs(9889) <= b and not a;
    outputs(9890) <= a;
    outputs(9891) <= not a;
    outputs(9892) <= not (a or b);
    outputs(9893) <= a xor b;
    outputs(9894) <= b;
    outputs(9895) <= a;
    outputs(9896) <= not a;
    outputs(9897) <= not b;
    outputs(9898) <= not b;
    outputs(9899) <= not a;
    outputs(9900) <= not a;
    outputs(9901) <= not a;
    outputs(9902) <= a and b;
    outputs(9903) <= not b or a;
    outputs(9904) <= not b;
    outputs(9905) <= not (a or b);
    outputs(9906) <= b and not a;
    outputs(9907) <= a xor b;
    outputs(9908) <= not a;
    outputs(9909) <= a and b;
    outputs(9910) <= not b or a;
    outputs(9911) <= a;
    outputs(9912) <= a xor b;
    outputs(9913) <= not b;
    outputs(9914) <= not (a and b);
    outputs(9915) <= a;
    outputs(9916) <= a xor b;
    outputs(9917) <= a;
    outputs(9918) <= not a;
    outputs(9919) <= a and b;
    outputs(9920) <= a and b;
    outputs(9921) <= not (a xor b);
    outputs(9922) <= not (a xor b);
    outputs(9923) <= not b;
    outputs(9924) <= a xor b;
    outputs(9925) <= a and b;
    outputs(9926) <= not (a or b);
    outputs(9927) <= not b;
    outputs(9928) <= a xor b;
    outputs(9929) <= a xor b;
    outputs(9930) <= b;
    outputs(9931) <= a;
    outputs(9932) <= not (a or b);
    outputs(9933) <= a;
    outputs(9934) <= not (a xor b);
    outputs(9935) <= b;
    outputs(9936) <= b and not a;
    outputs(9937) <= not a;
    outputs(9938) <= not (a xor b);
    outputs(9939) <= a;
    outputs(9940) <= a;
    outputs(9941) <= a;
    outputs(9942) <= not (a xor b);
    outputs(9943) <= not b;
    outputs(9944) <= not (a xor b);
    outputs(9945) <= a and not b;
    outputs(9946) <= a;
    outputs(9947) <= not (a and b);
    outputs(9948) <= b and not a;
    outputs(9949) <= not (a xor b);
    outputs(9950) <= b;
    outputs(9951) <= a and b;
    outputs(9952) <= not (a xor b);
    outputs(9953) <= not (a or b);
    outputs(9954) <= a;
    outputs(9955) <= not a;
    outputs(9956) <= not (a and b);
    outputs(9957) <= b and not a;
    outputs(9958) <= a;
    outputs(9959) <= not (a xor b);
    outputs(9960) <= not a or b;
    outputs(9961) <= not a or b;
    outputs(9962) <= not a;
    outputs(9963) <= not b;
    outputs(9964) <= a;
    outputs(9965) <= not b;
    outputs(9966) <= not (a xor b);
    outputs(9967) <= a;
    outputs(9968) <= not (a xor b);
    outputs(9969) <= not b;
    outputs(9970) <= not (a xor b);
    outputs(9971) <= not b;
    outputs(9972) <= a;
    outputs(9973) <= a xor b;
    outputs(9974) <= a;
    outputs(9975) <= a and b;
    outputs(9976) <= a and b;
    outputs(9977) <= a xor b;
    outputs(9978) <= a xor b;
    outputs(9979) <= a or b;
    outputs(9980) <= a xor b;
    outputs(9981) <= a xor b;
    outputs(9982) <= not (a xor b);
    outputs(9983) <= not (a xor b);
    outputs(9984) <= not a;
    outputs(9985) <= a and not b;
    outputs(9986) <= not a;
    outputs(9987) <= b;
    outputs(9988) <= a and not b;
    outputs(9989) <= a xor b;
    outputs(9990) <= a xor b;
    outputs(9991) <= not a;
    outputs(9992) <= not a;
    outputs(9993) <= not (a and b);
    outputs(9994) <= a and not b;
    outputs(9995) <= not b or a;
    outputs(9996) <= not (a xor b);
    outputs(9997) <= a xor b;
    outputs(9998) <= not (a xor b);
    outputs(9999) <= not (a xor b);
    outputs(10000) <= not b;
    outputs(10001) <= not (a xor b);
    outputs(10002) <= a xor b;
    outputs(10003) <= not a;
    outputs(10004) <= a;
    outputs(10005) <= not a;
    outputs(10006) <= a xor b;
    outputs(10007) <= a;
    outputs(10008) <= not (a or b);
    outputs(10009) <= not b;
    outputs(10010) <= not (a or b);
    outputs(10011) <= not b;
    outputs(10012) <= not (a or b);
    outputs(10013) <= not (a and b);
    outputs(10014) <= not (a xor b);
    outputs(10015) <= a and not b;
    outputs(10016) <= not (a xor b);
    outputs(10017) <= a xor b;
    outputs(10018) <= not a;
    outputs(10019) <= a xor b;
    outputs(10020) <= not a;
    outputs(10021) <= a or b;
    outputs(10022) <= a xor b;
    outputs(10023) <= not a;
    outputs(10024) <= not b;
    outputs(10025) <= not a or b;
    outputs(10026) <= not b;
    outputs(10027) <= not a or b;
    outputs(10028) <= not a;
    outputs(10029) <= not (a xor b);
    outputs(10030) <= a and not b;
    outputs(10031) <= b and not a;
    outputs(10032) <= a xor b;
    outputs(10033) <= b;
    outputs(10034) <= not (a and b);
    outputs(10035) <= not a;
    outputs(10036) <= not (a xor b);
    outputs(10037) <= not b;
    outputs(10038) <= a and b;
    outputs(10039) <= not a;
    outputs(10040) <= a and b;
    outputs(10041) <= '0';
    outputs(10042) <= not a;
    outputs(10043) <= not (a xor b);
    outputs(10044) <= a and not b;
    outputs(10045) <= b and not a;
    outputs(10046) <= a;
    outputs(10047) <= b;
    outputs(10048) <= a xor b;
    outputs(10049) <= b;
    outputs(10050) <= a or b;
    outputs(10051) <= not (a or b);
    outputs(10052) <= a xor b;
    outputs(10053) <= not (a xor b);
    outputs(10054) <= a xor b;
    outputs(10055) <= not (a xor b);
    outputs(10056) <= not b;
    outputs(10057) <= a;
    outputs(10058) <= b;
    outputs(10059) <= a;
    outputs(10060) <= a xor b;
    outputs(10061) <= a and b;
    outputs(10062) <= not (a or b);
    outputs(10063) <= not a;
    outputs(10064) <= a xor b;
    outputs(10065) <= b and not a;
    outputs(10066) <= a and b;
    outputs(10067) <= a xor b;
    outputs(10068) <= b and not a;
    outputs(10069) <= not a;
    outputs(10070) <= b and not a;
    outputs(10071) <= a or b;
    outputs(10072) <= b and not a;
    outputs(10073) <= not b;
    outputs(10074) <= not a;
    outputs(10075) <= not b or a;
    outputs(10076) <= not (a or b);
    outputs(10077) <= not a;
    outputs(10078) <= a xor b;
    outputs(10079) <= a xor b;
    outputs(10080) <= not (a xor b);
    outputs(10081) <= not a;
    outputs(10082) <= a xor b;
    outputs(10083) <= a xor b;
    outputs(10084) <= not (a xor b);
    outputs(10085) <= b;
    outputs(10086) <= not b;
    outputs(10087) <= b;
    outputs(10088) <= b;
    outputs(10089) <= a and b;
    outputs(10090) <= a and not b;
    outputs(10091) <= not a;
    outputs(10092) <= b;
    outputs(10093) <= a;
    outputs(10094) <= a xor b;
    outputs(10095) <= a xor b;
    outputs(10096) <= a and not b;
    outputs(10097) <= a xor b;
    outputs(10098) <= b;
    outputs(10099) <= not b;
    outputs(10100) <= a xor b;
    outputs(10101) <= a xor b;
    outputs(10102) <= a xor b;
    outputs(10103) <= a xor b;
    outputs(10104) <= a xor b;
    outputs(10105) <= a;
    outputs(10106) <= not b;
    outputs(10107) <= not b or a;
    outputs(10108) <= not (a xor b);
    outputs(10109) <= b;
    outputs(10110) <= not (a or b);
    outputs(10111) <= '1';
    outputs(10112) <= not (a xor b);
    outputs(10113) <= a xor b;
    outputs(10114) <= b;
    outputs(10115) <= not b;
    outputs(10116) <= a;
    outputs(10117) <= a;
    outputs(10118) <= a and not b;
    outputs(10119) <= not a;
    outputs(10120) <= a;
    outputs(10121) <= not a;
    outputs(10122) <= a or b;
    outputs(10123) <= not (a xor b);
    outputs(10124) <= a xor b;
    outputs(10125) <= not b;
    outputs(10126) <= a xor b;
    outputs(10127) <= a and b;
    outputs(10128) <= a xor b;
    outputs(10129) <= not (a and b);
    outputs(10130) <= not (a xor b);
    outputs(10131) <= a xor b;
    outputs(10132) <= not b;
    outputs(10133) <= a and b;
    outputs(10134) <= not (a or b);
    outputs(10135) <= not (a xor b);
    outputs(10136) <= a;
    outputs(10137) <= b and not a;
    outputs(10138) <= a xor b;
    outputs(10139) <= a and not b;
    outputs(10140) <= a and not b;
    outputs(10141) <= not (a xor b);
    outputs(10142) <= a;
    outputs(10143) <= a xor b;
    outputs(10144) <= not (a xor b);
    outputs(10145) <= b;
    outputs(10146) <= not a;
    outputs(10147) <= a and not b;
    outputs(10148) <= not (a xor b);
    outputs(10149) <= a;
    outputs(10150) <= not (a or b);
    outputs(10151) <= a and not b;
    outputs(10152) <= a;
    outputs(10153) <= not (a xor b);
    outputs(10154) <= a;
    outputs(10155) <= a xor b;
    outputs(10156) <= a;
    outputs(10157) <= b and not a;
    outputs(10158) <= a and not b;
    outputs(10159) <= b and not a;
    outputs(10160) <= a xor b;
    outputs(10161) <= b;
    outputs(10162) <= not (a xor b);
    outputs(10163) <= a xor b;
    outputs(10164) <= not (a xor b);
    outputs(10165) <= not a;
    outputs(10166) <= not (a xor b);
    outputs(10167) <= b and not a;
    outputs(10168) <= not b;
    outputs(10169) <= a or b;
    outputs(10170) <= not (a and b);
    outputs(10171) <= not (a xor b);
    outputs(10172) <= b;
    outputs(10173) <= a;
    outputs(10174) <= a and not b;
    outputs(10175) <= not b;
    outputs(10176) <= not (a xor b);
    outputs(10177) <= not b;
    outputs(10178) <= not b;
    outputs(10179) <= not a;
    outputs(10180) <= a and not b;
    outputs(10181) <= a;
    outputs(10182) <= not a;
    outputs(10183) <= not (a xor b);
    outputs(10184) <= b;
    outputs(10185) <= not b;
    outputs(10186) <= not (a xor b);
    outputs(10187) <= b;
    outputs(10188) <= not (a xor b);
    outputs(10189) <= not b;
    outputs(10190) <= not a or b;
    outputs(10191) <= not (a xor b);
    outputs(10192) <= a and not b;
    outputs(10193) <= not a;
    outputs(10194) <= not b;
    outputs(10195) <= a xor b;
    outputs(10196) <= a and not b;
    outputs(10197) <= a and b;
    outputs(10198) <= not (a xor b);
    outputs(10199) <= a and b;
    outputs(10200) <= a;
    outputs(10201) <= a xor b;
    outputs(10202) <= not a;
    outputs(10203) <= not b or a;
    outputs(10204) <= a and not b;
    outputs(10205) <= b;
    outputs(10206) <= not (a xor b);
    outputs(10207) <= a xor b;
    outputs(10208) <= a and b;
    outputs(10209) <= a xor b;
    outputs(10210) <= a xor b;
    outputs(10211) <= not (a xor b);
    outputs(10212) <= a;
    outputs(10213) <= not a;
    outputs(10214) <= b and not a;
    outputs(10215) <= not b;
    outputs(10216) <= a xor b;
    outputs(10217) <= a;
    outputs(10218) <= a and b;
    outputs(10219) <= not b;
    outputs(10220) <= not (a xor b);
    outputs(10221) <= not a;
    outputs(10222) <= a xor b;
    outputs(10223) <= not (a xor b);
    outputs(10224) <= not (a xor b);
    outputs(10225) <= a and not b;
    outputs(10226) <= not (a xor b);
    outputs(10227) <= not a;
    outputs(10228) <= a and b;
    outputs(10229) <= not a;
    outputs(10230) <= not (a and b);
    outputs(10231) <= not a;
    outputs(10232) <= a xor b;
    outputs(10233) <= a xor b;
    outputs(10234) <= not b;
    outputs(10235) <= a xor b;
    outputs(10236) <= not a;
    outputs(10237) <= a xor b;
    outputs(10238) <= a and b;
    outputs(10239) <= a;
end Behavioral;
