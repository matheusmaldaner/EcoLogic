library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs: in std_logic_vector(1023 downto 0);
        outputs: out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs: std_logic_vector(5119 downto 0);
    signal layer1_outputs: std_logic_vector(5119 downto 0);
    signal layer2_outputs: std_logic_vector(5119 downto 0);
    signal layer3_outputs: std_logic_vector(5119 downto 0);
    signal layer4_outputs: std_logic_vector(5119 downto 0);
    signal layer5_outputs: std_logic_vector(5119 downto 0);
    signal layer6_outputs: std_logic_vector(5119 downto 0);
    signal layer7_outputs: std_logic_vector(5119 downto 0);
    signal layer8_outputs: std_logic_vector(5119 downto 0);

begin
    layer0_outputs(0) <= '1';
    layer0_outputs(1) <= a and b;
    layer0_outputs(2) <= not b;
    layer0_outputs(3) <= a and b;
    layer0_outputs(4) <= b;
    layer0_outputs(5) <= '0';
    layer0_outputs(6) <= not a;
    layer0_outputs(7) <= a xor b;
    layer0_outputs(8) <= not (a or b);
    layer0_outputs(9) <= not a or b;
    layer0_outputs(10) <= a xor b;
    layer0_outputs(11) <= '0';
    layer0_outputs(12) <= not (a or b);
    layer0_outputs(13) <= '0';
    layer0_outputs(14) <= not (a or b);
    layer0_outputs(15) <= a and b;
    layer0_outputs(16) <= b;
    layer0_outputs(17) <= not a;
    layer0_outputs(18) <= a or b;
    layer0_outputs(19) <= a and b;
    layer0_outputs(20) <= a;
    layer0_outputs(21) <= b;
    layer0_outputs(22) <= a;
    layer0_outputs(23) <= not a;
    layer0_outputs(24) <= a and b;
    layer0_outputs(25) <= a and not b;
    layer0_outputs(26) <= '1';
    layer0_outputs(27) <= not b or a;
    layer0_outputs(28) <= not (a and b);
    layer0_outputs(29) <= not b;
    layer0_outputs(30) <= not a;
    layer0_outputs(31) <= a xor b;
    layer0_outputs(32) <= a xor b;
    layer0_outputs(33) <= not a;
    layer0_outputs(34) <= '1';
    layer0_outputs(35) <= not (a and b);
    layer0_outputs(36) <= a and not b;
    layer0_outputs(37) <= not a;
    layer0_outputs(38) <= not a or b;
    layer0_outputs(39) <= a or b;
    layer0_outputs(40) <= a and b;
    layer0_outputs(41) <= b;
    layer0_outputs(42) <= b and not a;
    layer0_outputs(43) <= a or b;
    layer0_outputs(44) <= not a or b;
    layer0_outputs(45) <= not (a xor b);
    layer0_outputs(46) <= '0';
    layer0_outputs(47) <= not a or b;
    layer0_outputs(48) <= not (a or b);
    layer0_outputs(49) <= not b or a;
    layer0_outputs(50) <= not a;
    layer0_outputs(51) <= a and b;
    layer0_outputs(52) <= not (a and b);
    layer0_outputs(53) <= not a;
    layer0_outputs(54) <= '1';
    layer0_outputs(55) <= b and not a;
    layer0_outputs(56) <= not (a and b);
    layer0_outputs(57) <= '0';
    layer0_outputs(58) <= not (a and b);
    layer0_outputs(59) <= not b;
    layer0_outputs(60) <= a or b;
    layer0_outputs(61) <= a and b;
    layer0_outputs(62) <= a and not b;
    layer0_outputs(63) <= a xor b;
    layer0_outputs(64) <= not (a xor b);
    layer0_outputs(65) <= not (a or b);
    layer0_outputs(66) <= not b or a;
    layer0_outputs(67) <= not (a or b);
    layer0_outputs(68) <= '0';
    layer0_outputs(69) <= a or b;
    layer0_outputs(70) <= a;
    layer0_outputs(71) <= b and not a;
    layer0_outputs(72) <= not b or a;
    layer0_outputs(73) <= not a;
    layer0_outputs(74) <= not a;
    layer0_outputs(75) <= a or b;
    layer0_outputs(76) <= b;
    layer0_outputs(77) <= not b or a;
    layer0_outputs(78) <= a;
    layer0_outputs(79) <= a;
    layer0_outputs(80) <= not (a or b);
    layer0_outputs(81) <= not a;
    layer0_outputs(82) <= b;
    layer0_outputs(83) <= not b;
    layer0_outputs(84) <= not b;
    layer0_outputs(85) <= not (a and b);
    layer0_outputs(86) <= a or b;
    layer0_outputs(87) <= '0';
    layer0_outputs(88) <= not (a or b);
    layer0_outputs(89) <= a and not b;
    layer0_outputs(90) <= not b;
    layer0_outputs(91) <= not (a or b);
    layer0_outputs(92) <= not b or a;
    layer0_outputs(93) <= a xor b;
    layer0_outputs(94) <= a and b;
    layer0_outputs(95) <= b;
    layer0_outputs(96) <= a;
    layer0_outputs(97) <= '0';
    layer0_outputs(98) <= a and b;
    layer0_outputs(99) <= b;
    layer0_outputs(100) <= not b;
    layer0_outputs(101) <= '1';
    layer0_outputs(102) <= a or b;
    layer0_outputs(103) <= b and not a;
    layer0_outputs(104) <= not b or a;
    layer0_outputs(105) <= a xor b;
    layer0_outputs(106) <= a;
    layer0_outputs(107) <= not (a or b);
    layer0_outputs(108) <= a or b;
    layer0_outputs(109) <= a or b;
    layer0_outputs(110) <= not a or b;
    layer0_outputs(111) <= b;
    layer0_outputs(112) <= not b or a;
    layer0_outputs(113) <= a and b;
    layer0_outputs(114) <= '0';
    layer0_outputs(115) <= not a;
    layer0_outputs(116) <= b and not a;
    layer0_outputs(117) <= not b or a;
    layer0_outputs(118) <= '1';
    layer0_outputs(119) <= a xor b;
    layer0_outputs(120) <= a;
    layer0_outputs(121) <= not b or a;
    layer0_outputs(122) <= '0';
    layer0_outputs(123) <= not a or b;
    layer0_outputs(124) <= '0';
    layer0_outputs(125) <= a;
    layer0_outputs(126) <= not b or a;
    layer0_outputs(127) <= not a or b;
    layer0_outputs(128) <= a xor b;
    layer0_outputs(129) <= a and not b;
    layer0_outputs(130) <= a and not b;
    layer0_outputs(131) <= b and not a;
    layer0_outputs(132) <= a and b;
    layer0_outputs(133) <= not b;
    layer0_outputs(134) <= not a;
    layer0_outputs(135) <= not (a or b);
    layer0_outputs(136) <= not (a xor b);
    layer0_outputs(137) <= a and not b;
    layer0_outputs(138) <= not (a or b);
    layer0_outputs(139) <= not a or b;
    layer0_outputs(140) <= b;
    layer0_outputs(141) <= '1';
    layer0_outputs(142) <= a xor b;
    layer0_outputs(143) <= not a;
    layer0_outputs(144) <= '0';
    layer0_outputs(145) <= a xor b;
    layer0_outputs(146) <= not (a and b);
    layer0_outputs(147) <= '0';
    layer0_outputs(148) <= a xor b;
    layer0_outputs(149) <= not (a xor b);
    layer0_outputs(150) <= not (a xor b);
    layer0_outputs(151) <= a or b;
    layer0_outputs(152) <= '0';
    layer0_outputs(153) <= b;
    layer0_outputs(154) <= not a;
    layer0_outputs(155) <= not (a and b);
    layer0_outputs(156) <= a and not b;
    layer0_outputs(157) <= not a;
    layer0_outputs(158) <= b and not a;
    layer0_outputs(159) <= not a or b;
    layer0_outputs(160) <= not a;
    layer0_outputs(161) <= b;
    layer0_outputs(162) <= a or b;
    layer0_outputs(163) <= not (a and b);
    layer0_outputs(164) <= not (a or b);
    layer0_outputs(165) <= not (a xor b);
    layer0_outputs(166) <= not b or a;
    layer0_outputs(167) <= '0';
    layer0_outputs(168) <= a xor b;
    layer0_outputs(169) <= b and not a;
    layer0_outputs(170) <= not b or a;
    layer0_outputs(171) <= a;
    layer0_outputs(172) <= a;
    layer0_outputs(173) <= '0';
    layer0_outputs(174) <= not (a xor b);
    layer0_outputs(175) <= b;
    layer0_outputs(176) <= a and b;
    layer0_outputs(177) <= not b;
    layer0_outputs(178) <= not (a or b);
    layer0_outputs(179) <= not a;
    layer0_outputs(180) <= not b;
    layer0_outputs(181) <= b and not a;
    layer0_outputs(182) <= not a or b;
    layer0_outputs(183) <= not a or b;
    layer0_outputs(184) <= not b;
    layer0_outputs(185) <= b and not a;
    layer0_outputs(186) <= '1';
    layer0_outputs(187) <= b;
    layer0_outputs(188) <= '0';
    layer0_outputs(189) <= a and b;
    layer0_outputs(190) <= a and b;
    layer0_outputs(191) <= a xor b;
    layer0_outputs(192) <= not b;
    layer0_outputs(193) <= b and not a;
    layer0_outputs(194) <= a;
    layer0_outputs(195) <= a xor b;
    layer0_outputs(196) <= '0';
    layer0_outputs(197) <= not b or a;
    layer0_outputs(198) <= not b;
    layer0_outputs(199) <= not (a xor b);
    layer0_outputs(200) <= a;
    layer0_outputs(201) <= not (a or b);
    layer0_outputs(202) <= not a or b;
    layer0_outputs(203) <= '0';
    layer0_outputs(204) <= b;
    layer0_outputs(205) <= not b;
    layer0_outputs(206) <= not (a or b);
    layer0_outputs(207) <= not (a or b);
    layer0_outputs(208) <= a xor b;
    layer0_outputs(209) <= '1';
    layer0_outputs(210) <= not (a xor b);
    layer0_outputs(211) <= not a;
    layer0_outputs(212) <= '1';
    layer0_outputs(213) <= '0';
    layer0_outputs(214) <= '0';
    layer0_outputs(215) <= not b;
    layer0_outputs(216) <= not (a and b);
    layer0_outputs(217) <= b and not a;
    layer0_outputs(218) <= a and not b;
    layer0_outputs(219) <= '0';
    layer0_outputs(220) <= b and not a;
    layer0_outputs(221) <= not (a xor b);
    layer0_outputs(222) <= '0';
    layer0_outputs(223) <= b and not a;
    layer0_outputs(224) <= '1';
    layer0_outputs(225) <= not b;
    layer0_outputs(226) <= not b or a;
    layer0_outputs(227) <= b and not a;
    layer0_outputs(228) <= b;
    layer0_outputs(229) <= a and b;
    layer0_outputs(230) <= b;
    layer0_outputs(231) <= not a;
    layer0_outputs(232) <= b and not a;
    layer0_outputs(233) <= b and not a;
    layer0_outputs(234) <= not (a xor b);
    layer0_outputs(235) <= a and not b;
    layer0_outputs(236) <= not (a and b);
    layer0_outputs(237) <= b and not a;
    layer0_outputs(238) <= not b or a;
    layer0_outputs(239) <= not (a or b);
    layer0_outputs(240) <= not (a or b);
    layer0_outputs(241) <= b;
    layer0_outputs(242) <= not a;
    layer0_outputs(243) <= not b or a;
    layer0_outputs(244) <= a and b;
    layer0_outputs(245) <= b;
    layer0_outputs(246) <= a and b;
    layer0_outputs(247) <= not a;
    layer0_outputs(248) <= not (a or b);
    layer0_outputs(249) <= a xor b;
    layer0_outputs(250) <= a and not b;
    layer0_outputs(251) <= b and not a;
    layer0_outputs(252) <= not (a xor b);
    layer0_outputs(253) <= b and not a;
    layer0_outputs(254) <= not (a xor b);
    layer0_outputs(255) <= '0';
    layer0_outputs(256) <= not (a or b);
    layer0_outputs(257) <= not (a xor b);
    layer0_outputs(258) <= a xor b;
    layer0_outputs(259) <= not b or a;
    layer0_outputs(260) <= not a or b;
    layer0_outputs(261) <= not b or a;
    layer0_outputs(262) <= not b;
    layer0_outputs(263) <= a or b;
    layer0_outputs(264) <= a;
    layer0_outputs(265) <= '1';
    layer0_outputs(266) <= a;
    layer0_outputs(267) <= '1';
    layer0_outputs(268) <= not (a or b);
    layer0_outputs(269) <= a and b;
    layer0_outputs(270) <= '1';
    layer0_outputs(271) <= a;
    layer0_outputs(272) <= b and not a;
    layer0_outputs(273) <= '1';
    layer0_outputs(274) <= a and b;
    layer0_outputs(275) <= not (a and b);
    layer0_outputs(276) <= a and b;
    layer0_outputs(277) <= not a;
    layer0_outputs(278) <= '1';
    layer0_outputs(279) <= not (a xor b);
    layer0_outputs(280) <= '0';
    layer0_outputs(281) <= not (a xor b);
    layer0_outputs(282) <= not a or b;
    layer0_outputs(283) <= '1';
    layer0_outputs(284) <= a and b;
    layer0_outputs(285) <= a xor b;
    layer0_outputs(286) <= a or b;
    layer0_outputs(287) <= not b;
    layer0_outputs(288) <= a and not b;
    layer0_outputs(289) <= '1';
    layer0_outputs(290) <= not a or b;
    layer0_outputs(291) <= not b;
    layer0_outputs(292) <= not a;
    layer0_outputs(293) <= b and not a;
    layer0_outputs(294) <= a;
    layer0_outputs(295) <= not b or a;
    layer0_outputs(296) <= '0';
    layer0_outputs(297) <= '0';
    layer0_outputs(298) <= not b;
    layer0_outputs(299) <= not a or b;
    layer0_outputs(300) <= not a or b;
    layer0_outputs(301) <= '1';
    layer0_outputs(302) <= a and not b;
    layer0_outputs(303) <= '0';
    layer0_outputs(304) <= a;
    layer0_outputs(305) <= '1';
    layer0_outputs(306) <= a and b;
    layer0_outputs(307) <= a and b;
    layer0_outputs(308) <= a xor b;
    layer0_outputs(309) <= '0';
    layer0_outputs(310) <= a and not b;
    layer0_outputs(311) <= a;
    layer0_outputs(312) <= a or b;
    layer0_outputs(313) <= '1';
    layer0_outputs(314) <= not (a and b);
    layer0_outputs(315) <= a and not b;
    layer0_outputs(316) <= not b or a;
    layer0_outputs(317) <= a or b;
    layer0_outputs(318) <= not (a and b);
    layer0_outputs(319) <= not b;
    layer0_outputs(320) <= a xor b;
    layer0_outputs(321) <= not (a xor b);
    layer0_outputs(322) <= not b;
    layer0_outputs(323) <= not b;
    layer0_outputs(324) <= b;
    layer0_outputs(325) <= a xor b;
    layer0_outputs(326) <= a xor b;
    layer0_outputs(327) <= not a;
    layer0_outputs(328) <= a and not b;
    layer0_outputs(329) <= a and not b;
    layer0_outputs(330) <= not (a xor b);
    layer0_outputs(331) <= '1';
    layer0_outputs(332) <= not b;
    layer0_outputs(333) <= b and not a;
    layer0_outputs(334) <= a and b;
    layer0_outputs(335) <= not a;
    layer0_outputs(336) <= not a or b;
    layer0_outputs(337) <= not a or b;
    layer0_outputs(338) <= a and b;
    layer0_outputs(339) <= not a or b;
    layer0_outputs(340) <= a;
    layer0_outputs(341) <= not (a xor b);
    layer0_outputs(342) <= '1';
    layer0_outputs(343) <= b;
    layer0_outputs(344) <= a and not b;
    layer0_outputs(345) <= not (a xor b);
    layer0_outputs(346) <= a and not b;
    layer0_outputs(347) <= b;
    layer0_outputs(348) <= a or b;
    layer0_outputs(349) <= not a;
    layer0_outputs(350) <= b and not a;
    layer0_outputs(351) <= '1';
    layer0_outputs(352) <= a and b;
    layer0_outputs(353) <= not b or a;
    layer0_outputs(354) <= a and b;
    layer0_outputs(355) <= not b or a;
    layer0_outputs(356) <= '1';
    layer0_outputs(357) <= not a;
    layer0_outputs(358) <= not a;
    layer0_outputs(359) <= not (a or b);
    layer0_outputs(360) <= '1';
    layer0_outputs(361) <= not a;
    layer0_outputs(362) <= a;
    layer0_outputs(363) <= a and b;
    layer0_outputs(364) <= a xor b;
    layer0_outputs(365) <= not (a xor b);
    layer0_outputs(366) <= not b or a;
    layer0_outputs(367) <= '1';
    layer0_outputs(368) <= a or b;
    layer0_outputs(369) <= not b;
    layer0_outputs(370) <= not a;
    layer0_outputs(371) <= a;
    layer0_outputs(372) <= b;
    layer0_outputs(373) <= a and not b;
    layer0_outputs(374) <= b;
    layer0_outputs(375) <= not b or a;
    layer0_outputs(376) <= not (a or b);
    layer0_outputs(377) <= a xor b;
    layer0_outputs(378) <= not (a or b);
    layer0_outputs(379) <= not b or a;
    layer0_outputs(380) <= a and not b;
    layer0_outputs(381) <= a and b;
    layer0_outputs(382) <= '1';
    layer0_outputs(383) <= not b;
    layer0_outputs(384) <= '0';
    layer0_outputs(385) <= a;
    layer0_outputs(386) <= b and not a;
    layer0_outputs(387) <= not b;
    layer0_outputs(388) <= a;
    layer0_outputs(389) <= a and b;
    layer0_outputs(390) <= not b;
    layer0_outputs(391) <= '0';
    layer0_outputs(392) <= not b;
    layer0_outputs(393) <= b and not a;
    layer0_outputs(394) <= not (a and b);
    layer0_outputs(395) <= a xor b;
    layer0_outputs(396) <= not (a and b);
    layer0_outputs(397) <= a and not b;
    layer0_outputs(398) <= b;
    layer0_outputs(399) <= not a;
    layer0_outputs(400) <= b;
    layer0_outputs(401) <= a and not b;
    layer0_outputs(402) <= a or b;
    layer0_outputs(403) <= not a or b;
    layer0_outputs(404) <= b;
    layer0_outputs(405) <= a and b;
    layer0_outputs(406) <= a;
    layer0_outputs(407) <= a;
    layer0_outputs(408) <= a and not b;
    layer0_outputs(409) <= not a or b;
    layer0_outputs(410) <= '1';
    layer0_outputs(411) <= not a;
    layer0_outputs(412) <= a or b;
    layer0_outputs(413) <= not (a and b);
    layer0_outputs(414) <= not (a and b);
    layer0_outputs(415) <= not (a xor b);
    layer0_outputs(416) <= a and b;
    layer0_outputs(417) <= '0';
    layer0_outputs(418) <= not (a and b);
    layer0_outputs(419) <= not a or b;
    layer0_outputs(420) <= '0';
    layer0_outputs(421) <= not (a and b);
    layer0_outputs(422) <= not (a xor b);
    layer0_outputs(423) <= a;
    layer0_outputs(424) <= not (a or b);
    layer0_outputs(425) <= '0';
    layer0_outputs(426) <= a;
    layer0_outputs(427) <= not b or a;
    layer0_outputs(428) <= a and b;
    layer0_outputs(429) <= a and not b;
    layer0_outputs(430) <= a or b;
    layer0_outputs(431) <= '0';
    layer0_outputs(432) <= '0';
    layer0_outputs(433) <= '0';
    layer0_outputs(434) <= not (a and b);
    layer0_outputs(435) <= not (a xor b);
    layer0_outputs(436) <= a and b;
    layer0_outputs(437) <= not (a or b);
    layer0_outputs(438) <= a or b;
    layer0_outputs(439) <= not (a xor b);
    layer0_outputs(440) <= not (a and b);
    layer0_outputs(441) <= '0';
    layer0_outputs(442) <= not (a xor b);
    layer0_outputs(443) <= not b or a;
    layer0_outputs(444) <= not a;
    layer0_outputs(445) <= a;
    layer0_outputs(446) <= not b or a;
    layer0_outputs(447) <= a xor b;
    layer0_outputs(448) <= not b;
    layer0_outputs(449) <= a xor b;
    layer0_outputs(450) <= a;
    layer0_outputs(451) <= a and not b;
    layer0_outputs(452) <= not a;
    layer0_outputs(453) <= not b or a;
    layer0_outputs(454) <= b;
    layer0_outputs(455) <= not b;
    layer0_outputs(456) <= '0';
    layer0_outputs(457) <= not (a and b);
    layer0_outputs(458) <= a or b;
    layer0_outputs(459) <= a and b;
    layer0_outputs(460) <= a and b;
    layer0_outputs(461) <= a or b;
    layer0_outputs(462) <= not b;
    layer0_outputs(463) <= a;
    layer0_outputs(464) <= not b;
    layer0_outputs(465) <= a and b;
    layer0_outputs(466) <= '1';
    layer0_outputs(467) <= not a or b;
    layer0_outputs(468) <= b;
    layer0_outputs(469) <= not a or b;
    layer0_outputs(470) <= '1';
    layer0_outputs(471) <= a and b;
    layer0_outputs(472) <= '0';
    layer0_outputs(473) <= not b or a;
    layer0_outputs(474) <= b and not a;
    layer0_outputs(475) <= not b or a;
    layer0_outputs(476) <= not a;
    layer0_outputs(477) <= '1';
    layer0_outputs(478) <= not b;
    layer0_outputs(479) <= not (a or b);
    layer0_outputs(480) <= '0';
    layer0_outputs(481) <= not (a xor b);
    layer0_outputs(482) <= '1';
    layer0_outputs(483) <= b;
    layer0_outputs(484) <= '0';
    layer0_outputs(485) <= not (a or b);
    layer0_outputs(486) <= a and not b;
    layer0_outputs(487) <= not a or b;
    layer0_outputs(488) <= not (a xor b);
    layer0_outputs(489) <= not a;
    layer0_outputs(490) <= not a or b;
    layer0_outputs(491) <= '0';
    layer0_outputs(492) <= '1';
    layer0_outputs(493) <= not b;
    layer0_outputs(494) <= not a or b;
    layer0_outputs(495) <= not a or b;
    layer0_outputs(496) <= not b;
    layer0_outputs(497) <= b and not a;
    layer0_outputs(498) <= a and b;
    layer0_outputs(499) <= not a;
    layer0_outputs(500) <= a;
    layer0_outputs(501) <= a or b;
    layer0_outputs(502) <= not (a and b);
    layer0_outputs(503) <= b;
    layer0_outputs(504) <= not a;
    layer0_outputs(505) <= b and not a;
    layer0_outputs(506) <= not b or a;
    layer0_outputs(507) <= not a or b;
    layer0_outputs(508) <= not (a and b);
    layer0_outputs(509) <= a;
    layer0_outputs(510) <= b;
    layer0_outputs(511) <= not a;
    layer0_outputs(512) <= not (a xor b);
    layer0_outputs(513) <= b and not a;
    layer0_outputs(514) <= not (a and b);
    layer0_outputs(515) <= b and not a;
    layer0_outputs(516) <= not (a or b);
    layer0_outputs(517) <= not (a and b);
    layer0_outputs(518) <= not b;
    layer0_outputs(519) <= not (a or b);
    layer0_outputs(520) <= b and not a;
    layer0_outputs(521) <= not (a and b);
    layer0_outputs(522) <= '1';
    layer0_outputs(523) <= not a;
    layer0_outputs(524) <= '1';
    layer0_outputs(525) <= not b;
    layer0_outputs(526) <= a;
    layer0_outputs(527) <= a xor b;
    layer0_outputs(528) <= a or b;
    layer0_outputs(529) <= not b or a;
    layer0_outputs(530) <= b;
    layer0_outputs(531) <= not a or b;
    layer0_outputs(532) <= b and not a;
    layer0_outputs(533) <= a or b;
    layer0_outputs(534) <= a xor b;
    layer0_outputs(535) <= a;
    layer0_outputs(536) <= '0';
    layer0_outputs(537) <= a and not b;
    layer0_outputs(538) <= a and b;
    layer0_outputs(539) <= not b;
    layer0_outputs(540) <= a;
    layer0_outputs(541) <= a and b;
    layer0_outputs(542) <= not a;
    layer0_outputs(543) <= a or b;
    layer0_outputs(544) <= not (a xor b);
    layer0_outputs(545) <= '1';
    layer0_outputs(546) <= a;
    layer0_outputs(547) <= not a or b;
    layer0_outputs(548) <= a;
    layer0_outputs(549) <= '0';
    layer0_outputs(550) <= b;
    layer0_outputs(551) <= '1';
    layer0_outputs(552) <= '1';
    layer0_outputs(553) <= a and not b;
    layer0_outputs(554) <= not b or a;
    layer0_outputs(555) <= not a or b;
    layer0_outputs(556) <= not (a xor b);
    layer0_outputs(557) <= not a or b;
    layer0_outputs(558) <= '1';
    layer0_outputs(559) <= not b or a;
    layer0_outputs(560) <= '1';
    layer0_outputs(561) <= a and not b;
    layer0_outputs(562) <= b;
    layer0_outputs(563) <= not (a and b);
    layer0_outputs(564) <= a and not b;
    layer0_outputs(565) <= not (a and b);
    layer0_outputs(566) <= not a;
    layer0_outputs(567) <= not a;
    layer0_outputs(568) <= not (a or b);
    layer0_outputs(569) <= not a or b;
    layer0_outputs(570) <= not b or a;
    layer0_outputs(571) <= a xor b;
    layer0_outputs(572) <= a;
    layer0_outputs(573) <= not (a and b);
    layer0_outputs(574) <= not a;
    layer0_outputs(575) <= not (a or b);
    layer0_outputs(576) <= a xor b;
    layer0_outputs(577) <= a;
    layer0_outputs(578) <= '0';
    layer0_outputs(579) <= a xor b;
    layer0_outputs(580) <= b and not a;
    layer0_outputs(581) <= not b or a;
    layer0_outputs(582) <= '0';
    layer0_outputs(583) <= not a or b;
    layer0_outputs(584) <= a;
    layer0_outputs(585) <= not a;
    layer0_outputs(586) <= a and not b;
    layer0_outputs(587) <= not b;
    layer0_outputs(588) <= not a or b;
    layer0_outputs(589) <= a or b;
    layer0_outputs(590) <= '0';
    layer0_outputs(591) <= a;
    layer0_outputs(592) <= not (a or b);
    layer0_outputs(593) <= not (a xor b);
    layer0_outputs(594) <= not (a xor b);
    layer0_outputs(595) <= a and b;
    layer0_outputs(596) <= a or b;
    layer0_outputs(597) <= not a or b;
    layer0_outputs(598) <= not a or b;
    layer0_outputs(599) <= not b or a;
    layer0_outputs(600) <= a or b;
    layer0_outputs(601) <= not a;
    layer0_outputs(602) <= b and not a;
    layer0_outputs(603) <= b;
    layer0_outputs(604) <= a and b;
    layer0_outputs(605) <= b and not a;
    layer0_outputs(606) <= not a;
    layer0_outputs(607) <= b;
    layer0_outputs(608) <= b and not a;
    layer0_outputs(609) <= not a;
    layer0_outputs(610) <= '1';
    layer0_outputs(611) <= a xor b;
    layer0_outputs(612) <= b and not a;
    layer0_outputs(613) <= a and b;
    layer0_outputs(614) <= not a or b;
    layer0_outputs(615) <= not a or b;
    layer0_outputs(616) <= a;
    layer0_outputs(617) <= a xor b;
    layer0_outputs(618) <= a and not b;
    layer0_outputs(619) <= a and b;
    layer0_outputs(620) <= not (a and b);
    layer0_outputs(621) <= b;
    layer0_outputs(622) <= not a or b;
    layer0_outputs(623) <= not b or a;
    layer0_outputs(624) <= '1';
    layer0_outputs(625) <= '1';
    layer0_outputs(626) <= a and b;
    layer0_outputs(627) <= '0';
    layer0_outputs(628) <= a and b;
    layer0_outputs(629) <= '1';
    layer0_outputs(630) <= not b or a;
    layer0_outputs(631) <= a xor b;
    layer0_outputs(632) <= a xor b;
    layer0_outputs(633) <= not a or b;
    layer0_outputs(634) <= not b;
    layer0_outputs(635) <= not a;
    layer0_outputs(636) <= '0';
    layer0_outputs(637) <= not (a or b);
    layer0_outputs(638) <= not b or a;
    layer0_outputs(639) <= a and not b;
    layer0_outputs(640) <= '0';
    layer0_outputs(641) <= not (a and b);
    layer0_outputs(642) <= not (a or b);
    layer0_outputs(643) <= b and not a;
    layer0_outputs(644) <= not (a and b);
    layer0_outputs(645) <= b and not a;
    layer0_outputs(646) <= a or b;
    layer0_outputs(647) <= not b or a;
    layer0_outputs(648) <= not b or a;
    layer0_outputs(649) <= '0';
    layer0_outputs(650) <= '0';
    layer0_outputs(651) <= a and b;
    layer0_outputs(652) <= '0';
    layer0_outputs(653) <= not (a or b);
    layer0_outputs(654) <= a;
    layer0_outputs(655) <= a;
    layer0_outputs(656) <= not (a or b);
    layer0_outputs(657) <= b and not a;
    layer0_outputs(658) <= b and not a;
    layer0_outputs(659) <= a and b;
    layer0_outputs(660) <= '0';
    layer0_outputs(661) <= not (a and b);
    layer0_outputs(662) <= '1';
    layer0_outputs(663) <= not (a xor b);
    layer0_outputs(664) <= not (a and b);
    layer0_outputs(665) <= b and not a;
    layer0_outputs(666) <= not (a xor b);
    layer0_outputs(667) <= not (a xor b);
    layer0_outputs(668) <= not (a and b);
    layer0_outputs(669) <= not b or a;
    layer0_outputs(670) <= a xor b;
    layer0_outputs(671) <= a;
    layer0_outputs(672) <= '1';
    layer0_outputs(673) <= a;
    layer0_outputs(674) <= not (a and b);
    layer0_outputs(675) <= not a;
    layer0_outputs(676) <= '0';
    layer0_outputs(677) <= a;
    layer0_outputs(678) <= a and b;
    layer0_outputs(679) <= a;
    layer0_outputs(680) <= '0';
    layer0_outputs(681) <= not (a or b);
    layer0_outputs(682) <= a and b;
    layer0_outputs(683) <= not (a xor b);
    layer0_outputs(684) <= a and not b;
    layer0_outputs(685) <= a and not b;
    layer0_outputs(686) <= a or b;
    layer0_outputs(687) <= not (a xor b);
    layer0_outputs(688) <= a xor b;
    layer0_outputs(689) <= a;
    layer0_outputs(690) <= '1';
    layer0_outputs(691) <= a;
    layer0_outputs(692) <= a xor b;
    layer0_outputs(693) <= not a;
    layer0_outputs(694) <= a;
    layer0_outputs(695) <= a and not b;
    layer0_outputs(696) <= a and not b;
    layer0_outputs(697) <= '1';
    layer0_outputs(698) <= not b;
    layer0_outputs(699) <= a and not b;
    layer0_outputs(700) <= b;
    layer0_outputs(701) <= b;
    layer0_outputs(702) <= a or b;
    layer0_outputs(703) <= a xor b;
    layer0_outputs(704) <= '1';
    layer0_outputs(705) <= a and b;
    layer0_outputs(706) <= not b or a;
    layer0_outputs(707) <= b and not a;
    layer0_outputs(708) <= '1';
    layer0_outputs(709) <= not a;
    layer0_outputs(710) <= a and b;
    layer0_outputs(711) <= a;
    layer0_outputs(712) <= b;
    layer0_outputs(713) <= a;
    layer0_outputs(714) <= not a or b;
    layer0_outputs(715) <= not (a xor b);
    layer0_outputs(716) <= not (a or b);
    layer0_outputs(717) <= a;
    layer0_outputs(718) <= not b;
    layer0_outputs(719) <= not a or b;
    layer0_outputs(720) <= not a or b;
    layer0_outputs(721) <= b;
    layer0_outputs(722) <= a or b;
    layer0_outputs(723) <= b;
    layer0_outputs(724) <= not a;
    layer0_outputs(725) <= b and not a;
    layer0_outputs(726) <= b;
    layer0_outputs(727) <= not (a and b);
    layer0_outputs(728) <= not (a and b);
    layer0_outputs(729) <= not b or a;
    layer0_outputs(730) <= b and not a;
    layer0_outputs(731) <= not a or b;
    layer0_outputs(732) <= a and b;
    layer0_outputs(733) <= '1';
    layer0_outputs(734) <= not (a xor b);
    layer0_outputs(735) <= a;
    layer0_outputs(736) <= not a;
    layer0_outputs(737) <= b;
    layer0_outputs(738) <= not (a or b);
    layer0_outputs(739) <= a or b;
    layer0_outputs(740) <= not (a or b);
    layer0_outputs(741) <= not (a and b);
    layer0_outputs(742) <= b;
    layer0_outputs(743) <= b and not a;
    layer0_outputs(744) <= not (a or b);
    layer0_outputs(745) <= not (a xor b);
    layer0_outputs(746) <= b;
    layer0_outputs(747) <= a;
    layer0_outputs(748) <= not a or b;
    layer0_outputs(749) <= not b or a;
    layer0_outputs(750) <= '1';
    layer0_outputs(751) <= a xor b;
    layer0_outputs(752) <= a or b;
    layer0_outputs(753) <= not b;
    layer0_outputs(754) <= b and not a;
    layer0_outputs(755) <= a and b;
    layer0_outputs(756) <= not b or a;
    layer0_outputs(757) <= '1';
    layer0_outputs(758) <= b and not a;
    layer0_outputs(759) <= a and not b;
    layer0_outputs(760) <= not b;
    layer0_outputs(761) <= not a;
    layer0_outputs(762) <= not (a and b);
    layer0_outputs(763) <= a xor b;
    layer0_outputs(764) <= not b or a;
    layer0_outputs(765) <= a or b;
    layer0_outputs(766) <= not (a or b);
    layer0_outputs(767) <= a and b;
    layer0_outputs(768) <= not (a and b);
    layer0_outputs(769) <= not (a or b);
    layer0_outputs(770) <= b;
    layer0_outputs(771) <= '1';
    layer0_outputs(772) <= not b;
    layer0_outputs(773) <= a xor b;
    layer0_outputs(774) <= not (a xor b);
    layer0_outputs(775) <= '0';
    layer0_outputs(776) <= a and b;
    layer0_outputs(777) <= b;
    layer0_outputs(778) <= a and b;
    layer0_outputs(779) <= not b;
    layer0_outputs(780) <= b;
    layer0_outputs(781) <= not (a or b);
    layer0_outputs(782) <= a or b;
    layer0_outputs(783) <= a and b;
    layer0_outputs(784) <= a;
    layer0_outputs(785) <= a;
    layer0_outputs(786) <= '0';
    layer0_outputs(787) <= '0';
    layer0_outputs(788) <= a;
    layer0_outputs(789) <= a xor b;
    layer0_outputs(790) <= a or b;
    layer0_outputs(791) <= '0';
    layer0_outputs(792) <= not (a and b);
    layer0_outputs(793) <= a or b;
    layer0_outputs(794) <= not b or a;
    layer0_outputs(795) <= '1';
    layer0_outputs(796) <= not a;
    layer0_outputs(797) <= a and b;
    layer0_outputs(798) <= a and not b;
    layer0_outputs(799) <= a;
    layer0_outputs(800) <= not (a and b);
    layer0_outputs(801) <= b and not a;
    layer0_outputs(802) <= a and not b;
    layer0_outputs(803) <= not (a or b);
    layer0_outputs(804) <= b and not a;
    layer0_outputs(805) <= b;
    layer0_outputs(806) <= a and not b;
    layer0_outputs(807) <= not (a and b);
    layer0_outputs(808) <= a;
    layer0_outputs(809) <= not b or a;
    layer0_outputs(810) <= not b;
    layer0_outputs(811) <= not a or b;
    layer0_outputs(812) <= not (a and b);
    layer0_outputs(813) <= b and not a;
    layer0_outputs(814) <= not a or b;
    layer0_outputs(815) <= a and not b;
    layer0_outputs(816) <= '1';
    layer0_outputs(817) <= a and b;
    layer0_outputs(818) <= not (a or b);
    layer0_outputs(819) <= not (a or b);
    layer0_outputs(820) <= a;
    layer0_outputs(821) <= b;
    layer0_outputs(822) <= not (a xor b);
    layer0_outputs(823) <= a and b;
    layer0_outputs(824) <= not a or b;
    layer0_outputs(825) <= not a or b;
    layer0_outputs(826) <= not b;
    layer0_outputs(827) <= b;
    layer0_outputs(828) <= not a or b;
    layer0_outputs(829) <= a and not b;
    layer0_outputs(830) <= not b;
    layer0_outputs(831) <= a;
    layer0_outputs(832) <= a or b;
    layer0_outputs(833) <= '1';
    layer0_outputs(834) <= not (a or b);
    layer0_outputs(835) <= b;
    layer0_outputs(836) <= not (a or b);
    layer0_outputs(837) <= '0';
    layer0_outputs(838) <= a xor b;
    layer0_outputs(839) <= a and b;
    layer0_outputs(840) <= not b;
    layer0_outputs(841) <= not b or a;
    layer0_outputs(842) <= not b;
    layer0_outputs(843) <= not (a or b);
    layer0_outputs(844) <= a;
    layer0_outputs(845) <= not b or a;
    layer0_outputs(846) <= not (a or b);
    layer0_outputs(847) <= a;
    layer0_outputs(848) <= '1';
    layer0_outputs(849) <= a or b;
    layer0_outputs(850) <= a xor b;
    layer0_outputs(851) <= b;
    layer0_outputs(852) <= not b;
    layer0_outputs(853) <= a xor b;
    layer0_outputs(854) <= a xor b;
    layer0_outputs(855) <= '1';
    layer0_outputs(856) <= not (a and b);
    layer0_outputs(857) <= b and not a;
    layer0_outputs(858) <= not (a and b);
    layer0_outputs(859) <= '0';
    layer0_outputs(860) <= '0';
    layer0_outputs(861) <= not b;
    layer0_outputs(862) <= '0';
    layer0_outputs(863) <= not (a and b);
    layer0_outputs(864) <= '1';
    layer0_outputs(865) <= not (a and b);
    layer0_outputs(866) <= not b;
    layer0_outputs(867) <= not (a or b);
    layer0_outputs(868) <= b and not a;
    layer0_outputs(869) <= '1';
    layer0_outputs(870) <= not a;
    layer0_outputs(871) <= not a or b;
    layer0_outputs(872) <= not (a or b);
    layer0_outputs(873) <= not (a xor b);
    layer0_outputs(874) <= b and not a;
    layer0_outputs(875) <= not (a or b);
    layer0_outputs(876) <= b and not a;
    layer0_outputs(877) <= not (a and b);
    layer0_outputs(878) <= a or b;
    layer0_outputs(879) <= a and not b;
    layer0_outputs(880) <= not a;
    layer0_outputs(881) <= a;
    layer0_outputs(882) <= not a;
    layer0_outputs(883) <= not a;
    layer0_outputs(884) <= not b;
    layer0_outputs(885) <= not a;
    layer0_outputs(886) <= not (a and b);
    layer0_outputs(887) <= b;
    layer0_outputs(888) <= not (a or b);
    layer0_outputs(889) <= a or b;
    layer0_outputs(890) <= '1';
    layer0_outputs(891) <= not b;
    layer0_outputs(892) <= not b or a;
    layer0_outputs(893) <= not b or a;
    layer0_outputs(894) <= not (a and b);
    layer0_outputs(895) <= not (a or b);
    layer0_outputs(896) <= not (a and b);
    layer0_outputs(897) <= not b;
    layer0_outputs(898) <= b and not a;
    layer0_outputs(899) <= '1';
    layer0_outputs(900) <= not b;
    layer0_outputs(901) <= a xor b;
    layer0_outputs(902) <= not (a or b);
    layer0_outputs(903) <= a or b;
    layer0_outputs(904) <= not a or b;
    layer0_outputs(905) <= a and b;
    layer0_outputs(906) <= b;
    layer0_outputs(907) <= a or b;
    layer0_outputs(908) <= not a;
    layer0_outputs(909) <= not (a xor b);
    layer0_outputs(910) <= not (a and b);
    layer0_outputs(911) <= not b or a;
    layer0_outputs(912) <= not (a or b);
    layer0_outputs(913) <= not b;
    layer0_outputs(914) <= a xor b;
    layer0_outputs(915) <= a;
    layer0_outputs(916) <= a and b;
    layer0_outputs(917) <= not (a and b);
    layer0_outputs(918) <= a;
    layer0_outputs(919) <= '1';
    layer0_outputs(920) <= a or b;
    layer0_outputs(921) <= not a or b;
    layer0_outputs(922) <= not (a or b);
    layer0_outputs(923) <= not a;
    layer0_outputs(924) <= '0';
    layer0_outputs(925) <= not a;
    layer0_outputs(926) <= b;
    layer0_outputs(927) <= not a or b;
    layer0_outputs(928) <= a and b;
    layer0_outputs(929) <= b and not a;
    layer0_outputs(930) <= b and not a;
    layer0_outputs(931) <= a and not b;
    layer0_outputs(932) <= not a or b;
    layer0_outputs(933) <= a or b;
    layer0_outputs(934) <= b and not a;
    layer0_outputs(935) <= not (a and b);
    layer0_outputs(936) <= '1';
    layer0_outputs(937) <= not (a or b);
    layer0_outputs(938) <= '1';
    layer0_outputs(939) <= not (a and b);
    layer0_outputs(940) <= a and not b;
    layer0_outputs(941) <= not (a xor b);
    layer0_outputs(942) <= b;
    layer0_outputs(943) <= b;
    layer0_outputs(944) <= a or b;
    layer0_outputs(945) <= b;
    layer0_outputs(946) <= a and not b;
    layer0_outputs(947) <= b and not a;
    layer0_outputs(948) <= not b or a;
    layer0_outputs(949) <= not a or b;
    layer0_outputs(950) <= a or b;
    layer0_outputs(951) <= not (a and b);
    layer0_outputs(952) <= not b or a;
    layer0_outputs(953) <= b and not a;
    layer0_outputs(954) <= a or b;
    layer0_outputs(955) <= a xor b;
    layer0_outputs(956) <= '0';
    layer0_outputs(957) <= b and not a;
    layer0_outputs(958) <= b and not a;
    layer0_outputs(959) <= not a;
    layer0_outputs(960) <= a and b;
    layer0_outputs(961) <= '1';
    layer0_outputs(962) <= a;
    layer0_outputs(963) <= a xor b;
    layer0_outputs(964) <= a and not b;
    layer0_outputs(965) <= a and b;
    layer0_outputs(966) <= b and not a;
    layer0_outputs(967) <= a and not b;
    layer0_outputs(968) <= b;
    layer0_outputs(969) <= not a or b;
    layer0_outputs(970) <= a xor b;
    layer0_outputs(971) <= b;
    layer0_outputs(972) <= not (a or b);
    layer0_outputs(973) <= not a;
    layer0_outputs(974) <= a and b;
    layer0_outputs(975) <= not a or b;
    layer0_outputs(976) <= not (a and b);
    layer0_outputs(977) <= b and not a;
    layer0_outputs(978) <= b and not a;
    layer0_outputs(979) <= a xor b;
    layer0_outputs(980) <= not (a or b);
    layer0_outputs(981) <= not (a or b);
    layer0_outputs(982) <= a and b;
    layer0_outputs(983) <= a and b;
    layer0_outputs(984) <= '0';
    layer0_outputs(985) <= a or b;
    layer0_outputs(986) <= not a;
    layer0_outputs(987) <= not (a xor b);
    layer0_outputs(988) <= not (a and b);
    layer0_outputs(989) <= a or b;
    layer0_outputs(990) <= '0';
    layer0_outputs(991) <= a or b;
    layer0_outputs(992) <= not a;
    layer0_outputs(993) <= not (a or b);
    layer0_outputs(994) <= not a;
    layer0_outputs(995) <= a and b;
    layer0_outputs(996) <= not b;
    layer0_outputs(997) <= not a or b;
    layer0_outputs(998) <= b;
    layer0_outputs(999) <= not (a and b);
    layer0_outputs(1000) <= '0';
    layer0_outputs(1001) <= not b or a;
    layer0_outputs(1002) <= not (a xor b);
    layer0_outputs(1003) <= a and not b;
    layer0_outputs(1004) <= a and b;
    layer0_outputs(1005) <= not b;
    layer0_outputs(1006) <= not b or a;
    layer0_outputs(1007) <= '1';
    layer0_outputs(1008) <= a;
    layer0_outputs(1009) <= '1';
    layer0_outputs(1010) <= b;
    layer0_outputs(1011) <= not b or a;
    layer0_outputs(1012) <= not (a and b);
    layer0_outputs(1013) <= not (a or b);
    layer0_outputs(1014) <= b;
    layer0_outputs(1015) <= a and not b;
    layer0_outputs(1016) <= b and not a;
    layer0_outputs(1017) <= not a or b;
    layer0_outputs(1018) <= a and b;
    layer0_outputs(1019) <= '0';
    layer0_outputs(1020) <= '0';
    layer0_outputs(1021) <= '1';
    layer0_outputs(1022) <= not (a or b);
    layer0_outputs(1023) <= b and not a;
    layer0_outputs(1024) <= not a or b;
    layer0_outputs(1025) <= b and not a;
    layer0_outputs(1026) <= a;
    layer0_outputs(1027) <= a and b;
    layer0_outputs(1028) <= not (a or b);
    layer0_outputs(1029) <= not b;
    layer0_outputs(1030) <= not (a or b);
    layer0_outputs(1031) <= '0';
    layer0_outputs(1032) <= a or b;
    layer0_outputs(1033) <= '0';
    layer0_outputs(1034) <= a or b;
    layer0_outputs(1035) <= not (a and b);
    layer0_outputs(1036) <= '1';
    layer0_outputs(1037) <= a and b;
    layer0_outputs(1038) <= a;
    layer0_outputs(1039) <= not a;
    layer0_outputs(1040) <= not (a xor b);
    layer0_outputs(1041) <= not (a xor b);
    layer0_outputs(1042) <= a and not b;
    layer0_outputs(1043) <= b and not a;
    layer0_outputs(1044) <= a;
    layer0_outputs(1045) <= b;
    layer0_outputs(1046) <= not (a xor b);
    layer0_outputs(1047) <= a and b;
    layer0_outputs(1048) <= not (a xor b);
    layer0_outputs(1049) <= not (a or b);
    layer0_outputs(1050) <= not a or b;
    layer0_outputs(1051) <= a and not b;
    layer0_outputs(1052) <= a;
    layer0_outputs(1053) <= not (a xor b);
    layer0_outputs(1054) <= not (a and b);
    layer0_outputs(1055) <= '1';
    layer0_outputs(1056) <= a or b;
    layer0_outputs(1057) <= not a or b;
    layer0_outputs(1058) <= a and b;
    layer0_outputs(1059) <= not b;
    layer0_outputs(1060) <= b;
    layer0_outputs(1061) <= not (a or b);
    layer0_outputs(1062) <= not (a or b);
    layer0_outputs(1063) <= b;
    layer0_outputs(1064) <= b and not a;
    layer0_outputs(1065) <= '1';
    layer0_outputs(1066) <= a xor b;
    layer0_outputs(1067) <= not (a xor b);
    layer0_outputs(1068) <= '0';
    layer0_outputs(1069) <= '0';
    layer0_outputs(1070) <= a;
    layer0_outputs(1071) <= not b;
    layer0_outputs(1072) <= not (a or b);
    layer0_outputs(1073) <= not (a or b);
    layer0_outputs(1074) <= not b;
    layer0_outputs(1075) <= not a or b;
    layer0_outputs(1076) <= b and not a;
    layer0_outputs(1077) <= not (a and b);
    layer0_outputs(1078) <= '1';
    layer0_outputs(1079) <= a and b;
    layer0_outputs(1080) <= not b;
    layer0_outputs(1081) <= not (a or b);
    layer0_outputs(1082) <= a;
    layer0_outputs(1083) <= not (a xor b);
    layer0_outputs(1084) <= b;
    layer0_outputs(1085) <= '0';
    layer0_outputs(1086) <= not b or a;
    layer0_outputs(1087) <= a and b;
    layer0_outputs(1088) <= not a;
    layer0_outputs(1089) <= b;
    layer0_outputs(1090) <= '0';
    layer0_outputs(1091) <= '0';
    layer0_outputs(1092) <= not (a or b);
    layer0_outputs(1093) <= a or b;
    layer0_outputs(1094) <= not b;
    layer0_outputs(1095) <= not a or b;
    layer0_outputs(1096) <= a or b;
    layer0_outputs(1097) <= '0';
    layer0_outputs(1098) <= a or b;
    layer0_outputs(1099) <= a or b;
    layer0_outputs(1100) <= '1';
    layer0_outputs(1101) <= not b or a;
    layer0_outputs(1102) <= not b or a;
    layer0_outputs(1103) <= '0';
    layer0_outputs(1104) <= a and b;
    layer0_outputs(1105) <= not (a or b);
    layer0_outputs(1106) <= not b or a;
    layer0_outputs(1107) <= a and not b;
    layer0_outputs(1108) <= a xor b;
    layer0_outputs(1109) <= a and not b;
    layer0_outputs(1110) <= not b;
    layer0_outputs(1111) <= not (a or b);
    layer0_outputs(1112) <= '1';
    layer0_outputs(1113) <= not b;
    layer0_outputs(1114) <= not b or a;
    layer0_outputs(1115) <= not b or a;
    layer0_outputs(1116) <= a;
    layer0_outputs(1117) <= not a or b;
    layer0_outputs(1118) <= not a or b;
    layer0_outputs(1119) <= b and not a;
    layer0_outputs(1120) <= b;
    layer0_outputs(1121) <= not b;
    layer0_outputs(1122) <= a xor b;
    layer0_outputs(1123) <= not b;
    layer0_outputs(1124) <= not b;
    layer0_outputs(1125) <= a and not b;
    layer0_outputs(1126) <= b and not a;
    layer0_outputs(1127) <= a;
    layer0_outputs(1128) <= a and not b;
    layer0_outputs(1129) <= b;
    layer0_outputs(1130) <= not b;
    layer0_outputs(1131) <= not b;
    layer0_outputs(1132) <= '1';
    layer0_outputs(1133) <= b and not a;
    layer0_outputs(1134) <= not a or b;
    layer0_outputs(1135) <= '1';
    layer0_outputs(1136) <= b and not a;
    layer0_outputs(1137) <= a and b;
    layer0_outputs(1138) <= not (a and b);
    layer0_outputs(1139) <= not b or a;
    layer0_outputs(1140) <= not a or b;
    layer0_outputs(1141) <= not a or b;
    layer0_outputs(1142) <= not (a and b);
    layer0_outputs(1143) <= not (a xor b);
    layer0_outputs(1144) <= a and not b;
    layer0_outputs(1145) <= not b;
    layer0_outputs(1146) <= b and not a;
    layer0_outputs(1147) <= '0';
    layer0_outputs(1148) <= b and not a;
    layer0_outputs(1149) <= '1';
    layer0_outputs(1150) <= a and b;
    layer0_outputs(1151) <= b;
    layer0_outputs(1152) <= not (a or b);
    layer0_outputs(1153) <= '1';
    layer0_outputs(1154) <= not b or a;
    layer0_outputs(1155) <= b;
    layer0_outputs(1156) <= not a or b;
    layer0_outputs(1157) <= not (a and b);
    layer0_outputs(1158) <= not (a or b);
    layer0_outputs(1159) <= a;
    layer0_outputs(1160) <= b and not a;
    layer0_outputs(1161) <= not (a xor b);
    layer0_outputs(1162) <= not b;
    layer0_outputs(1163) <= a;
    layer0_outputs(1164) <= '0';
    layer0_outputs(1165) <= not b or a;
    layer0_outputs(1166) <= not (a or b);
    layer0_outputs(1167) <= b;
    layer0_outputs(1168) <= a;
    layer0_outputs(1169) <= not a;
    layer0_outputs(1170) <= not (a or b);
    layer0_outputs(1171) <= b and not a;
    layer0_outputs(1172) <= not a;
    layer0_outputs(1173) <= a;
    layer0_outputs(1174) <= a;
    layer0_outputs(1175) <= a and not b;
    layer0_outputs(1176) <= not b or a;
    layer0_outputs(1177) <= not b or a;
    layer0_outputs(1178) <= a;
    layer0_outputs(1179) <= a and not b;
    layer0_outputs(1180) <= a xor b;
    layer0_outputs(1181) <= not b or a;
    layer0_outputs(1182) <= '1';
    layer0_outputs(1183) <= a and b;
    layer0_outputs(1184) <= b and not a;
    layer0_outputs(1185) <= a or b;
    layer0_outputs(1186) <= a and b;
    layer0_outputs(1187) <= not b;
    layer0_outputs(1188) <= a and not b;
    layer0_outputs(1189) <= a;
    layer0_outputs(1190) <= '0';
    layer0_outputs(1191) <= not a;
    layer0_outputs(1192) <= b;
    layer0_outputs(1193) <= not b;
    layer0_outputs(1194) <= not a or b;
    layer0_outputs(1195) <= not a or b;
    layer0_outputs(1196) <= a or b;
    layer0_outputs(1197) <= b;
    layer0_outputs(1198) <= '0';
    layer0_outputs(1199) <= '0';
    layer0_outputs(1200) <= a;
    layer0_outputs(1201) <= not b;
    layer0_outputs(1202) <= b;
    layer0_outputs(1203) <= b;
    layer0_outputs(1204) <= a xor b;
    layer0_outputs(1205) <= not (a and b);
    layer0_outputs(1206) <= '1';
    layer0_outputs(1207) <= b;
    layer0_outputs(1208) <= not (a and b);
    layer0_outputs(1209) <= '0';
    layer0_outputs(1210) <= not a or b;
    layer0_outputs(1211) <= a and not b;
    layer0_outputs(1212) <= not (a xor b);
    layer0_outputs(1213) <= a or b;
    layer0_outputs(1214) <= not (a and b);
    layer0_outputs(1215) <= not (a and b);
    layer0_outputs(1216) <= a;
    layer0_outputs(1217) <= '0';
    layer0_outputs(1218) <= not b;
    layer0_outputs(1219) <= a and not b;
    layer0_outputs(1220) <= not b or a;
    layer0_outputs(1221) <= a and b;
    layer0_outputs(1222) <= not (a and b);
    layer0_outputs(1223) <= not (a and b);
    layer0_outputs(1224) <= not a;
    layer0_outputs(1225) <= a or b;
    layer0_outputs(1226) <= not a or b;
    layer0_outputs(1227) <= not (a or b);
    layer0_outputs(1228) <= '0';
    layer0_outputs(1229) <= b;
    layer0_outputs(1230) <= a or b;
    layer0_outputs(1231) <= a and b;
    layer0_outputs(1232) <= b;
    layer0_outputs(1233) <= not b;
    layer0_outputs(1234) <= a and b;
    layer0_outputs(1235) <= not (a or b);
    layer0_outputs(1236) <= a;
    layer0_outputs(1237) <= not b or a;
    layer0_outputs(1238) <= not (a xor b);
    layer0_outputs(1239) <= not b;
    layer0_outputs(1240) <= '0';
    layer0_outputs(1241) <= not b or a;
    layer0_outputs(1242) <= not b or a;
    layer0_outputs(1243) <= a;
    layer0_outputs(1244) <= a;
    layer0_outputs(1245) <= a and not b;
    layer0_outputs(1246) <= '0';
    layer0_outputs(1247) <= a or b;
    layer0_outputs(1248) <= a or b;
    layer0_outputs(1249) <= a and not b;
    layer0_outputs(1250) <= a;
    layer0_outputs(1251) <= a or b;
    layer0_outputs(1252) <= not b;
    layer0_outputs(1253) <= not b;
    layer0_outputs(1254) <= not (a and b);
    layer0_outputs(1255) <= not b;
    layer0_outputs(1256) <= '1';
    layer0_outputs(1257) <= '0';
    layer0_outputs(1258) <= '1';
    layer0_outputs(1259) <= a and b;
    layer0_outputs(1260) <= not b or a;
    layer0_outputs(1261) <= a and b;
    layer0_outputs(1262) <= not b;
    layer0_outputs(1263) <= not (a and b);
    layer0_outputs(1264) <= not a or b;
    layer0_outputs(1265) <= not (a xor b);
    layer0_outputs(1266) <= not b;
    layer0_outputs(1267) <= a and b;
    layer0_outputs(1268) <= not b or a;
    layer0_outputs(1269) <= a and not b;
    layer0_outputs(1270) <= not (a and b);
    layer0_outputs(1271) <= a and b;
    layer0_outputs(1272) <= '1';
    layer0_outputs(1273) <= not b;
    layer0_outputs(1274) <= '0';
    layer0_outputs(1275) <= b;
    layer0_outputs(1276) <= a and not b;
    layer0_outputs(1277) <= not b or a;
    layer0_outputs(1278) <= not a;
    layer0_outputs(1279) <= b;
    layer0_outputs(1280) <= a;
    layer0_outputs(1281) <= not b;
    layer0_outputs(1282) <= '1';
    layer0_outputs(1283) <= not a;
    layer0_outputs(1284) <= b;
    layer0_outputs(1285) <= '1';
    layer0_outputs(1286) <= a and not b;
    layer0_outputs(1287) <= a and b;
    layer0_outputs(1288) <= not a;
    layer0_outputs(1289) <= not b;
    layer0_outputs(1290) <= a and not b;
    layer0_outputs(1291) <= not a or b;
    layer0_outputs(1292) <= a or b;
    layer0_outputs(1293) <= b;
    layer0_outputs(1294) <= a;
    layer0_outputs(1295) <= a;
    layer0_outputs(1296) <= not a;
    layer0_outputs(1297) <= '0';
    layer0_outputs(1298) <= a xor b;
    layer0_outputs(1299) <= a and not b;
    layer0_outputs(1300) <= not a or b;
    layer0_outputs(1301) <= b and not a;
    layer0_outputs(1302) <= b;
    layer0_outputs(1303) <= a xor b;
    layer0_outputs(1304) <= not (a or b);
    layer0_outputs(1305) <= b and not a;
    layer0_outputs(1306) <= not (a and b);
    layer0_outputs(1307) <= a and b;
    layer0_outputs(1308) <= b;
    layer0_outputs(1309) <= a and not b;
    layer0_outputs(1310) <= not b;
    layer0_outputs(1311) <= not (a and b);
    layer0_outputs(1312) <= b;
    layer0_outputs(1313) <= '0';
    layer0_outputs(1314) <= a xor b;
    layer0_outputs(1315) <= not b or a;
    layer0_outputs(1316) <= not a or b;
    layer0_outputs(1317) <= not (a xor b);
    layer0_outputs(1318) <= a;
    layer0_outputs(1319) <= not a or b;
    layer0_outputs(1320) <= not (a or b);
    layer0_outputs(1321) <= not b or a;
    layer0_outputs(1322) <= b;
    layer0_outputs(1323) <= '1';
    layer0_outputs(1324) <= a and b;
    layer0_outputs(1325) <= b;
    layer0_outputs(1326) <= a and b;
    layer0_outputs(1327) <= a and not b;
    layer0_outputs(1328) <= not (a xor b);
    layer0_outputs(1329) <= a and not b;
    layer0_outputs(1330) <= not b;
    layer0_outputs(1331) <= not a;
    layer0_outputs(1332) <= not b;
    layer0_outputs(1333) <= '1';
    layer0_outputs(1334) <= '1';
    layer0_outputs(1335) <= a xor b;
    layer0_outputs(1336) <= a and not b;
    layer0_outputs(1337) <= '0';
    layer0_outputs(1338) <= not (a xor b);
    layer0_outputs(1339) <= b;
    layer0_outputs(1340) <= a xor b;
    layer0_outputs(1341) <= not b or a;
    layer0_outputs(1342) <= '0';
    layer0_outputs(1343) <= not (a or b);
    layer0_outputs(1344) <= a;
    layer0_outputs(1345) <= not (a and b);
    layer0_outputs(1346) <= '0';
    layer0_outputs(1347) <= not (a xor b);
    layer0_outputs(1348) <= not a;
    layer0_outputs(1349) <= a xor b;
    layer0_outputs(1350) <= a;
    layer0_outputs(1351) <= not b;
    layer0_outputs(1352) <= a and b;
    layer0_outputs(1353) <= not b;
    layer0_outputs(1354) <= '0';
    layer0_outputs(1355) <= not (a xor b);
    layer0_outputs(1356) <= a and b;
    layer0_outputs(1357) <= not b or a;
    layer0_outputs(1358) <= not b or a;
    layer0_outputs(1359) <= '0';
    layer0_outputs(1360) <= not (a or b);
    layer0_outputs(1361) <= a xor b;
    layer0_outputs(1362) <= not b;
    layer0_outputs(1363) <= not (a or b);
    layer0_outputs(1364) <= not (a and b);
    layer0_outputs(1365) <= a and b;
    layer0_outputs(1366) <= a or b;
    layer0_outputs(1367) <= not (a xor b);
    layer0_outputs(1368) <= a or b;
    layer0_outputs(1369) <= b and not a;
    layer0_outputs(1370) <= a xor b;
    layer0_outputs(1371) <= '1';
    layer0_outputs(1372) <= '0';
    layer0_outputs(1373) <= a or b;
    layer0_outputs(1374) <= b and not a;
    layer0_outputs(1375) <= '1';
    layer0_outputs(1376) <= a;
    layer0_outputs(1377) <= not (a xor b);
    layer0_outputs(1378) <= '1';
    layer0_outputs(1379) <= a and b;
    layer0_outputs(1380) <= a;
    layer0_outputs(1381) <= not (a and b);
    layer0_outputs(1382) <= not b;
    layer0_outputs(1383) <= a;
    layer0_outputs(1384) <= '0';
    layer0_outputs(1385) <= not (a or b);
    layer0_outputs(1386) <= not (a xor b);
    layer0_outputs(1387) <= a;
    layer0_outputs(1388) <= '0';
    layer0_outputs(1389) <= not b;
    layer0_outputs(1390) <= not a;
    layer0_outputs(1391) <= not (a and b);
    layer0_outputs(1392) <= not b;
    layer0_outputs(1393) <= not (a xor b);
    layer0_outputs(1394) <= '0';
    layer0_outputs(1395) <= '0';
    layer0_outputs(1396) <= '1';
    layer0_outputs(1397) <= b and not a;
    layer0_outputs(1398) <= not a or b;
    layer0_outputs(1399) <= not a;
    layer0_outputs(1400) <= not (a or b);
    layer0_outputs(1401) <= a xor b;
    layer0_outputs(1402) <= not (a or b);
    layer0_outputs(1403) <= not b;
    layer0_outputs(1404) <= not b or a;
    layer0_outputs(1405) <= not a or b;
    layer0_outputs(1406) <= '0';
    layer0_outputs(1407) <= not (a or b);
    layer0_outputs(1408) <= not a or b;
    layer0_outputs(1409) <= not b or a;
    layer0_outputs(1410) <= '1';
    layer0_outputs(1411) <= a or b;
    layer0_outputs(1412) <= not (a and b);
    layer0_outputs(1413) <= a or b;
    layer0_outputs(1414) <= not a or b;
    layer0_outputs(1415) <= '0';
    layer0_outputs(1416) <= '1';
    layer0_outputs(1417) <= a;
    layer0_outputs(1418) <= not b or a;
    layer0_outputs(1419) <= '0';
    layer0_outputs(1420) <= not a or b;
    layer0_outputs(1421) <= a and not b;
    layer0_outputs(1422) <= a or b;
    layer0_outputs(1423) <= '1';
    layer0_outputs(1424) <= b;
    layer0_outputs(1425) <= b and not a;
    layer0_outputs(1426) <= not b;
    layer0_outputs(1427) <= a;
    layer0_outputs(1428) <= b;
    layer0_outputs(1429) <= not (a and b);
    layer0_outputs(1430) <= not (a xor b);
    layer0_outputs(1431) <= not (a xor b);
    layer0_outputs(1432) <= not a or b;
    layer0_outputs(1433) <= not b;
    layer0_outputs(1434) <= not a;
    layer0_outputs(1435) <= not (a xor b);
    layer0_outputs(1436) <= '0';
    layer0_outputs(1437) <= not a;
    layer0_outputs(1438) <= not b or a;
    layer0_outputs(1439) <= not b or a;
    layer0_outputs(1440) <= '1';
    layer0_outputs(1441) <= not a;
    layer0_outputs(1442) <= not b or a;
    layer0_outputs(1443) <= not b;
    layer0_outputs(1444) <= not b;
    layer0_outputs(1445) <= not (a xor b);
    layer0_outputs(1446) <= b;
    layer0_outputs(1447) <= '0';
    layer0_outputs(1448) <= not a;
    layer0_outputs(1449) <= not b;
    layer0_outputs(1450) <= not a or b;
    layer0_outputs(1451) <= a;
    layer0_outputs(1452) <= not (a and b);
    layer0_outputs(1453) <= b;
    layer0_outputs(1454) <= a or b;
    layer0_outputs(1455) <= b;
    layer0_outputs(1456) <= '0';
    layer0_outputs(1457) <= not (a xor b);
    layer0_outputs(1458) <= not (a or b);
    layer0_outputs(1459) <= b;
    layer0_outputs(1460) <= not (a or b);
    layer0_outputs(1461) <= not a;
    layer0_outputs(1462) <= not a;
    layer0_outputs(1463) <= not b or a;
    layer0_outputs(1464) <= not a or b;
    layer0_outputs(1465) <= a or b;
    layer0_outputs(1466) <= not b;
    layer0_outputs(1467) <= not a;
    layer0_outputs(1468) <= '1';
    layer0_outputs(1469) <= b;
    layer0_outputs(1470) <= not (a and b);
    layer0_outputs(1471) <= '1';
    layer0_outputs(1472) <= not (a and b);
    layer0_outputs(1473) <= '1';
    layer0_outputs(1474) <= '0';
    layer0_outputs(1475) <= not b or a;
    layer0_outputs(1476) <= not b;
    layer0_outputs(1477) <= a or b;
    layer0_outputs(1478) <= a xor b;
    layer0_outputs(1479) <= not (a and b);
    layer0_outputs(1480) <= b and not a;
    layer0_outputs(1481) <= not b or a;
    layer0_outputs(1482) <= b and not a;
    layer0_outputs(1483) <= not a;
    layer0_outputs(1484) <= '0';
    layer0_outputs(1485) <= not (a or b);
    layer0_outputs(1486) <= not b;
    layer0_outputs(1487) <= not b or a;
    layer0_outputs(1488) <= a;
    layer0_outputs(1489) <= a and b;
    layer0_outputs(1490) <= b and not a;
    layer0_outputs(1491) <= not a or b;
    layer0_outputs(1492) <= a and not b;
    layer0_outputs(1493) <= a and not b;
    layer0_outputs(1494) <= '1';
    layer0_outputs(1495) <= '1';
    layer0_outputs(1496) <= not (a and b);
    layer0_outputs(1497) <= '1';
    layer0_outputs(1498) <= not (a and b);
    layer0_outputs(1499) <= a xor b;
    layer0_outputs(1500) <= a;
    layer0_outputs(1501) <= a or b;
    layer0_outputs(1502) <= a xor b;
    layer0_outputs(1503) <= '1';
    layer0_outputs(1504) <= '0';
    layer0_outputs(1505) <= not (a or b);
    layer0_outputs(1506) <= not b;
    layer0_outputs(1507) <= not b;
    layer0_outputs(1508) <= a and not b;
    layer0_outputs(1509) <= a;
    layer0_outputs(1510) <= not (a xor b);
    layer0_outputs(1511) <= not (a or b);
    layer0_outputs(1512) <= not b or a;
    layer0_outputs(1513) <= a and not b;
    layer0_outputs(1514) <= not b or a;
    layer0_outputs(1515) <= not (a or b);
    layer0_outputs(1516) <= not a;
    layer0_outputs(1517) <= b and not a;
    layer0_outputs(1518) <= a and b;
    layer0_outputs(1519) <= '1';
    layer0_outputs(1520) <= not b or a;
    layer0_outputs(1521) <= a and b;
    layer0_outputs(1522) <= '0';
    layer0_outputs(1523) <= not b or a;
    layer0_outputs(1524) <= b and not a;
    layer0_outputs(1525) <= '0';
    layer0_outputs(1526) <= '0';
    layer0_outputs(1527) <= b and not a;
    layer0_outputs(1528) <= not (a xor b);
    layer0_outputs(1529) <= '0';
    layer0_outputs(1530) <= b;
    layer0_outputs(1531) <= '1';
    layer0_outputs(1532) <= not a or b;
    layer0_outputs(1533) <= not (a and b);
    layer0_outputs(1534) <= a and b;
    layer0_outputs(1535) <= not (a or b);
    layer0_outputs(1536) <= a;
    layer0_outputs(1537) <= not b;
    layer0_outputs(1538) <= not (a xor b);
    layer0_outputs(1539) <= '0';
    layer0_outputs(1540) <= '0';
    layer0_outputs(1541) <= not a;
    layer0_outputs(1542) <= not b;
    layer0_outputs(1543) <= b;
    layer0_outputs(1544) <= not a;
    layer0_outputs(1545) <= b and not a;
    layer0_outputs(1546) <= '1';
    layer0_outputs(1547) <= a and b;
    layer0_outputs(1548) <= a xor b;
    layer0_outputs(1549) <= a xor b;
    layer0_outputs(1550) <= not (a xor b);
    layer0_outputs(1551) <= not b or a;
    layer0_outputs(1552) <= '0';
    layer0_outputs(1553) <= b;
    layer0_outputs(1554) <= a and not b;
    layer0_outputs(1555) <= not (a xor b);
    layer0_outputs(1556) <= a and not b;
    layer0_outputs(1557) <= a xor b;
    layer0_outputs(1558) <= not (a or b);
    layer0_outputs(1559) <= a and b;
    layer0_outputs(1560) <= not a;
    layer0_outputs(1561) <= '0';
    layer0_outputs(1562) <= b;
    layer0_outputs(1563) <= '0';
    layer0_outputs(1564) <= b and not a;
    layer0_outputs(1565) <= a;
    layer0_outputs(1566) <= a and not b;
    layer0_outputs(1567) <= '0';
    layer0_outputs(1568) <= b;
    layer0_outputs(1569) <= '0';
    layer0_outputs(1570) <= not b or a;
    layer0_outputs(1571) <= not a or b;
    layer0_outputs(1572) <= a or b;
    layer0_outputs(1573) <= b;
    layer0_outputs(1574) <= not (a or b);
    layer0_outputs(1575) <= b;
    layer0_outputs(1576) <= '1';
    layer0_outputs(1577) <= '0';
    layer0_outputs(1578) <= not (a xor b);
    layer0_outputs(1579) <= a and not b;
    layer0_outputs(1580) <= not (a and b);
    layer0_outputs(1581) <= not (a xor b);
    layer0_outputs(1582) <= not a;
    layer0_outputs(1583) <= not (a xor b);
    layer0_outputs(1584) <= not (a and b);
    layer0_outputs(1585) <= a;
    layer0_outputs(1586) <= a and b;
    layer0_outputs(1587) <= not (a and b);
    layer0_outputs(1588) <= not (a or b);
    layer0_outputs(1589) <= b;
    layer0_outputs(1590) <= not (a or b);
    layer0_outputs(1591) <= a or b;
    layer0_outputs(1592) <= not (a and b);
    layer0_outputs(1593) <= not b;
    layer0_outputs(1594) <= not a;
    layer0_outputs(1595) <= not (a or b);
    layer0_outputs(1596) <= b;
    layer0_outputs(1597) <= b and not a;
    layer0_outputs(1598) <= a;
    layer0_outputs(1599) <= '1';
    layer0_outputs(1600) <= not a;
    layer0_outputs(1601) <= a xor b;
    layer0_outputs(1602) <= not (a and b);
    layer0_outputs(1603) <= not (a or b);
    layer0_outputs(1604) <= a or b;
    layer0_outputs(1605) <= '0';
    layer0_outputs(1606) <= '1';
    layer0_outputs(1607) <= not a;
    layer0_outputs(1608) <= a or b;
    layer0_outputs(1609) <= not a or b;
    layer0_outputs(1610) <= a and b;
    layer0_outputs(1611) <= a;
    layer0_outputs(1612) <= a xor b;
    layer0_outputs(1613) <= a xor b;
    layer0_outputs(1614) <= not (a and b);
    layer0_outputs(1615) <= not b or a;
    layer0_outputs(1616) <= '1';
    layer0_outputs(1617) <= not b or a;
    layer0_outputs(1618) <= b and not a;
    layer0_outputs(1619) <= not a;
    layer0_outputs(1620) <= b and not a;
    layer0_outputs(1621) <= a xor b;
    layer0_outputs(1622) <= not b or a;
    layer0_outputs(1623) <= a or b;
    layer0_outputs(1624) <= '0';
    layer0_outputs(1625) <= not b or a;
    layer0_outputs(1626) <= '0';
    layer0_outputs(1627) <= '1';
    layer0_outputs(1628) <= not a;
    layer0_outputs(1629) <= not b or a;
    layer0_outputs(1630) <= b and not a;
    layer0_outputs(1631) <= '1';
    layer0_outputs(1632) <= '1';
    layer0_outputs(1633) <= not b;
    layer0_outputs(1634) <= not b;
    layer0_outputs(1635) <= not (a or b);
    layer0_outputs(1636) <= a and b;
    layer0_outputs(1637) <= '1';
    layer0_outputs(1638) <= not (a and b);
    layer0_outputs(1639) <= a and b;
    layer0_outputs(1640) <= not b or a;
    layer0_outputs(1641) <= a;
    layer0_outputs(1642) <= not (a and b);
    layer0_outputs(1643) <= not b;
    layer0_outputs(1644) <= a xor b;
    layer0_outputs(1645) <= not (a or b);
    layer0_outputs(1646) <= a;
    layer0_outputs(1647) <= '0';
    layer0_outputs(1648) <= not b;
    layer0_outputs(1649) <= b and not a;
    layer0_outputs(1650) <= b and not a;
    layer0_outputs(1651) <= a or b;
    layer0_outputs(1652) <= b;
    layer0_outputs(1653) <= '1';
    layer0_outputs(1654) <= '1';
    layer0_outputs(1655) <= a;
    layer0_outputs(1656) <= a and not b;
    layer0_outputs(1657) <= a;
    layer0_outputs(1658) <= a and b;
    layer0_outputs(1659) <= not (a and b);
    layer0_outputs(1660) <= not (a and b);
    layer0_outputs(1661) <= not (a or b);
    layer0_outputs(1662) <= a xor b;
    layer0_outputs(1663) <= b;
    layer0_outputs(1664) <= not a or b;
    layer0_outputs(1665) <= '1';
    layer0_outputs(1666) <= a and not b;
    layer0_outputs(1667) <= '0';
    layer0_outputs(1668) <= not b or a;
    layer0_outputs(1669) <= '1';
    layer0_outputs(1670) <= not b or a;
    layer0_outputs(1671) <= '1';
    layer0_outputs(1672) <= not b;
    layer0_outputs(1673) <= a or b;
    layer0_outputs(1674) <= a and b;
    layer0_outputs(1675) <= '1';
    layer0_outputs(1676) <= '1';
    layer0_outputs(1677) <= not b or a;
    layer0_outputs(1678) <= not (a and b);
    layer0_outputs(1679) <= not a;
    layer0_outputs(1680) <= not (a and b);
    layer0_outputs(1681) <= b;
    layer0_outputs(1682) <= a;
    layer0_outputs(1683) <= a or b;
    layer0_outputs(1684) <= not (a xor b);
    layer0_outputs(1685) <= not (a and b);
    layer0_outputs(1686) <= a and not b;
    layer0_outputs(1687) <= not b;
    layer0_outputs(1688) <= not (a xor b);
    layer0_outputs(1689) <= not a or b;
    layer0_outputs(1690) <= a and b;
    layer0_outputs(1691) <= a and not b;
    layer0_outputs(1692) <= not b or a;
    layer0_outputs(1693) <= a;
    layer0_outputs(1694) <= not (a and b);
    layer0_outputs(1695) <= not (a or b);
    layer0_outputs(1696) <= '1';
    layer0_outputs(1697) <= a and b;
    layer0_outputs(1698) <= b;
    layer0_outputs(1699) <= a;
    layer0_outputs(1700) <= not b;
    layer0_outputs(1701) <= not b;
    layer0_outputs(1702) <= b and not a;
    layer0_outputs(1703) <= '1';
    layer0_outputs(1704) <= a;
    layer0_outputs(1705) <= not (a or b);
    layer0_outputs(1706) <= a and not b;
    layer0_outputs(1707) <= '0';
    layer0_outputs(1708) <= b;
    layer0_outputs(1709) <= not (a and b);
    layer0_outputs(1710) <= not (a or b);
    layer0_outputs(1711) <= not a;
    layer0_outputs(1712) <= b;
    layer0_outputs(1713) <= not a;
    layer0_outputs(1714) <= a and not b;
    layer0_outputs(1715) <= a;
    layer0_outputs(1716) <= a;
    layer0_outputs(1717) <= not a or b;
    layer0_outputs(1718) <= not b;
    layer0_outputs(1719) <= a xor b;
    layer0_outputs(1720) <= a;
    layer0_outputs(1721) <= b and not a;
    layer0_outputs(1722) <= not b or a;
    layer0_outputs(1723) <= not b;
    layer0_outputs(1724) <= b;
    layer0_outputs(1725) <= not a;
    layer0_outputs(1726) <= '0';
    layer0_outputs(1727) <= a and not b;
    layer0_outputs(1728) <= a or b;
    layer0_outputs(1729) <= a and not b;
    layer0_outputs(1730) <= not (a and b);
    layer0_outputs(1731) <= '0';
    layer0_outputs(1732) <= not (a or b);
    layer0_outputs(1733) <= b and not a;
    layer0_outputs(1734) <= not a or b;
    layer0_outputs(1735) <= not a;
    layer0_outputs(1736) <= a and not b;
    layer0_outputs(1737) <= not b;
    layer0_outputs(1738) <= '0';
    layer0_outputs(1739) <= not b or a;
    layer0_outputs(1740) <= not b or a;
    layer0_outputs(1741) <= a xor b;
    layer0_outputs(1742) <= a;
    layer0_outputs(1743) <= not (a and b);
    layer0_outputs(1744) <= not (a or b);
    layer0_outputs(1745) <= a xor b;
    layer0_outputs(1746) <= not a or b;
    layer0_outputs(1747) <= '1';
    layer0_outputs(1748) <= not b;
    layer0_outputs(1749) <= not (a and b);
    layer0_outputs(1750) <= b;
    layer0_outputs(1751) <= b and not a;
    layer0_outputs(1752) <= not (a or b);
    layer0_outputs(1753) <= '0';
    layer0_outputs(1754) <= a;
    layer0_outputs(1755) <= not b;
    layer0_outputs(1756) <= not (a and b);
    layer0_outputs(1757) <= not b or a;
    layer0_outputs(1758) <= not (a or b);
    layer0_outputs(1759) <= not (a and b);
    layer0_outputs(1760) <= '0';
    layer0_outputs(1761) <= not a or b;
    layer0_outputs(1762) <= not (a and b);
    layer0_outputs(1763) <= not (a xor b);
    layer0_outputs(1764) <= '1';
    layer0_outputs(1765) <= b and not a;
    layer0_outputs(1766) <= not b;
    layer0_outputs(1767) <= a and not b;
    layer0_outputs(1768) <= not (a and b);
    layer0_outputs(1769) <= b;
    layer0_outputs(1770) <= b and not a;
    layer0_outputs(1771) <= not b;
    layer0_outputs(1772) <= a or b;
    layer0_outputs(1773) <= not a or b;
    layer0_outputs(1774) <= not (a and b);
    layer0_outputs(1775) <= a and not b;
    layer0_outputs(1776) <= not (a or b);
    layer0_outputs(1777) <= not (a and b);
    layer0_outputs(1778) <= not (a and b);
    layer0_outputs(1779) <= not b or a;
    layer0_outputs(1780) <= a;
    layer0_outputs(1781) <= not b;
    layer0_outputs(1782) <= a;
    layer0_outputs(1783) <= not (a xor b);
    layer0_outputs(1784) <= not a;
    layer0_outputs(1785) <= not b;
    layer0_outputs(1786) <= '1';
    layer0_outputs(1787) <= not (a and b);
    layer0_outputs(1788) <= not b;
    layer0_outputs(1789) <= not a;
    layer0_outputs(1790) <= a and b;
    layer0_outputs(1791) <= a;
    layer0_outputs(1792) <= a and b;
    layer0_outputs(1793) <= not (a and b);
    layer0_outputs(1794) <= '1';
    layer0_outputs(1795) <= a xor b;
    layer0_outputs(1796) <= a and b;
    layer0_outputs(1797) <= not (a xor b);
    layer0_outputs(1798) <= a xor b;
    layer0_outputs(1799) <= not b or a;
    layer0_outputs(1800) <= not a or b;
    layer0_outputs(1801) <= b and not a;
    layer0_outputs(1802) <= a and b;
    layer0_outputs(1803) <= '0';
    layer0_outputs(1804) <= not a;
    layer0_outputs(1805) <= '1';
    layer0_outputs(1806) <= '1';
    layer0_outputs(1807) <= a xor b;
    layer0_outputs(1808) <= '0';
    layer0_outputs(1809) <= not (a and b);
    layer0_outputs(1810) <= a xor b;
    layer0_outputs(1811) <= b and not a;
    layer0_outputs(1812) <= not (a and b);
    layer0_outputs(1813) <= not a or b;
    layer0_outputs(1814) <= a or b;
    layer0_outputs(1815) <= b;
    layer0_outputs(1816) <= '1';
    layer0_outputs(1817) <= a or b;
    layer0_outputs(1818) <= a;
    layer0_outputs(1819) <= not a;
    layer0_outputs(1820) <= not (a and b);
    layer0_outputs(1821) <= a or b;
    layer0_outputs(1822) <= b;
    layer0_outputs(1823) <= not a;
    layer0_outputs(1824) <= '0';
    layer0_outputs(1825) <= a;
    layer0_outputs(1826) <= '1';
    layer0_outputs(1827) <= not (a and b);
    layer0_outputs(1828) <= a and not b;
    layer0_outputs(1829) <= a or b;
    layer0_outputs(1830) <= a and not b;
    layer0_outputs(1831) <= '1';
    layer0_outputs(1832) <= not a;
    layer0_outputs(1833) <= a and not b;
    layer0_outputs(1834) <= b and not a;
    layer0_outputs(1835) <= not (a and b);
    layer0_outputs(1836) <= a or b;
    layer0_outputs(1837) <= not (a and b);
    layer0_outputs(1838) <= '0';
    layer0_outputs(1839) <= a and not b;
    layer0_outputs(1840) <= not b or a;
    layer0_outputs(1841) <= a or b;
    layer0_outputs(1842) <= a;
    layer0_outputs(1843) <= not a;
    layer0_outputs(1844) <= not a or b;
    layer0_outputs(1845) <= b and not a;
    layer0_outputs(1846) <= a and b;
    layer0_outputs(1847) <= not b or a;
    layer0_outputs(1848) <= not (a and b);
    layer0_outputs(1849) <= not (a or b);
    layer0_outputs(1850) <= not a or b;
    layer0_outputs(1851) <= a xor b;
    layer0_outputs(1852) <= not (a and b);
    layer0_outputs(1853) <= a and b;
    layer0_outputs(1854) <= '0';
    layer0_outputs(1855) <= not a or b;
    layer0_outputs(1856) <= b;
    layer0_outputs(1857) <= a or b;
    layer0_outputs(1858) <= not a or b;
    layer0_outputs(1859) <= '0';
    layer0_outputs(1860) <= a and not b;
    layer0_outputs(1861) <= not a;
    layer0_outputs(1862) <= b;
    layer0_outputs(1863) <= '1';
    layer0_outputs(1864) <= a or b;
    layer0_outputs(1865) <= a and not b;
    layer0_outputs(1866) <= a and b;
    layer0_outputs(1867) <= b;
    layer0_outputs(1868) <= not a;
    layer0_outputs(1869) <= a;
    layer0_outputs(1870) <= not (a xor b);
    layer0_outputs(1871) <= '1';
    layer0_outputs(1872) <= '1';
    layer0_outputs(1873) <= a;
    layer0_outputs(1874) <= not a;
    layer0_outputs(1875) <= a and b;
    layer0_outputs(1876) <= a or b;
    layer0_outputs(1877) <= '1';
    layer0_outputs(1878) <= not b or a;
    layer0_outputs(1879) <= b;
    layer0_outputs(1880) <= not (a xor b);
    layer0_outputs(1881) <= not b or a;
    layer0_outputs(1882) <= b and not a;
    layer0_outputs(1883) <= a;
    layer0_outputs(1884) <= a and not b;
    layer0_outputs(1885) <= not b or a;
    layer0_outputs(1886) <= not (a xor b);
    layer0_outputs(1887) <= a or b;
    layer0_outputs(1888) <= b and not a;
    layer0_outputs(1889) <= not (a and b);
    layer0_outputs(1890) <= not b or a;
    layer0_outputs(1891) <= not (a xor b);
    layer0_outputs(1892) <= not a;
    layer0_outputs(1893) <= not (a or b);
    layer0_outputs(1894) <= not a or b;
    layer0_outputs(1895) <= '1';
    layer0_outputs(1896) <= '1';
    layer0_outputs(1897) <= '1';
    layer0_outputs(1898) <= a xor b;
    layer0_outputs(1899) <= a and b;
    layer0_outputs(1900) <= not b;
    layer0_outputs(1901) <= '0';
    layer0_outputs(1902) <= '1';
    layer0_outputs(1903) <= a xor b;
    layer0_outputs(1904) <= '0';
    layer0_outputs(1905) <= not (a and b);
    layer0_outputs(1906) <= '1';
    layer0_outputs(1907) <= a xor b;
    layer0_outputs(1908) <= not a;
    layer0_outputs(1909) <= a and b;
    layer0_outputs(1910) <= not b;
    layer0_outputs(1911) <= not a;
    layer0_outputs(1912) <= a and not b;
    layer0_outputs(1913) <= '0';
    layer0_outputs(1914) <= not (a xor b);
    layer0_outputs(1915) <= not (a and b);
    layer0_outputs(1916) <= not (a or b);
    layer0_outputs(1917) <= not a or b;
    layer0_outputs(1918) <= not (a or b);
    layer0_outputs(1919) <= not b;
    layer0_outputs(1920) <= a;
    layer0_outputs(1921) <= a and b;
    layer0_outputs(1922) <= not a;
    layer0_outputs(1923) <= '1';
    layer0_outputs(1924) <= b;
    layer0_outputs(1925) <= not (a or b);
    layer0_outputs(1926) <= a and not b;
    layer0_outputs(1927) <= not a;
    layer0_outputs(1928) <= '0';
    layer0_outputs(1929) <= not a or b;
    layer0_outputs(1930) <= a or b;
    layer0_outputs(1931) <= b;
    layer0_outputs(1932) <= b;
    layer0_outputs(1933) <= '0';
    layer0_outputs(1934) <= '1';
    layer0_outputs(1935) <= a or b;
    layer0_outputs(1936) <= a or b;
    layer0_outputs(1937) <= a and b;
    layer0_outputs(1938) <= not (a or b);
    layer0_outputs(1939) <= not (a or b);
    layer0_outputs(1940) <= a;
    layer0_outputs(1941) <= a and b;
    layer0_outputs(1942) <= b;
    layer0_outputs(1943) <= not b;
    layer0_outputs(1944) <= a;
    layer0_outputs(1945) <= a and not b;
    layer0_outputs(1946) <= '1';
    layer0_outputs(1947) <= a and not b;
    layer0_outputs(1948) <= a or b;
    layer0_outputs(1949) <= not a or b;
    layer0_outputs(1950) <= a;
    layer0_outputs(1951) <= '0';
    layer0_outputs(1952) <= a and b;
    layer0_outputs(1953) <= not a or b;
    layer0_outputs(1954) <= a or b;
    layer0_outputs(1955) <= '1';
    layer0_outputs(1956) <= a and b;
    layer0_outputs(1957) <= '1';
    layer0_outputs(1958) <= not a or b;
    layer0_outputs(1959) <= not (a or b);
    layer0_outputs(1960) <= not a or b;
    layer0_outputs(1961) <= not (a or b);
    layer0_outputs(1962) <= not a;
    layer0_outputs(1963) <= not (a and b);
    layer0_outputs(1964) <= a xor b;
    layer0_outputs(1965) <= a;
    layer0_outputs(1966) <= a or b;
    layer0_outputs(1967) <= '0';
    layer0_outputs(1968) <= '0';
    layer0_outputs(1969) <= not (a or b);
    layer0_outputs(1970) <= not a;
    layer0_outputs(1971) <= a;
    layer0_outputs(1972) <= not (a or b);
    layer0_outputs(1973) <= '0';
    layer0_outputs(1974) <= not (a xor b);
    layer0_outputs(1975) <= a;
    layer0_outputs(1976) <= b and not a;
    layer0_outputs(1977) <= '1';
    layer0_outputs(1978) <= a;
    layer0_outputs(1979) <= a and b;
    layer0_outputs(1980) <= a or b;
    layer0_outputs(1981) <= not b or a;
    layer0_outputs(1982) <= a xor b;
    layer0_outputs(1983) <= a;
    layer0_outputs(1984) <= a or b;
    layer0_outputs(1985) <= a or b;
    layer0_outputs(1986) <= not b or a;
    layer0_outputs(1987) <= not (a or b);
    layer0_outputs(1988) <= b and not a;
    layer0_outputs(1989) <= not (a and b);
    layer0_outputs(1990) <= b;
    layer0_outputs(1991) <= '0';
    layer0_outputs(1992) <= '0';
    layer0_outputs(1993) <= not (a or b);
    layer0_outputs(1994) <= b and not a;
    layer0_outputs(1995) <= a and b;
    layer0_outputs(1996) <= '1';
    layer0_outputs(1997) <= a xor b;
    layer0_outputs(1998) <= b;
    layer0_outputs(1999) <= not a;
    layer0_outputs(2000) <= '1';
    layer0_outputs(2001) <= not a or b;
    layer0_outputs(2002) <= not b or a;
    layer0_outputs(2003) <= b and not a;
    layer0_outputs(2004) <= a and b;
    layer0_outputs(2005) <= '0';
    layer0_outputs(2006) <= a and b;
    layer0_outputs(2007) <= '1';
    layer0_outputs(2008) <= not a;
    layer0_outputs(2009) <= not (a or b);
    layer0_outputs(2010) <= not (a xor b);
    layer0_outputs(2011) <= a and not b;
    layer0_outputs(2012) <= not (a and b);
    layer0_outputs(2013) <= not (a xor b);
    layer0_outputs(2014) <= a xor b;
    layer0_outputs(2015) <= '0';
    layer0_outputs(2016) <= not b;
    layer0_outputs(2017) <= a;
    layer0_outputs(2018) <= b;
    layer0_outputs(2019) <= not b or a;
    layer0_outputs(2020) <= b and not a;
    layer0_outputs(2021) <= a or b;
    layer0_outputs(2022) <= a xor b;
    layer0_outputs(2023) <= not (a xor b);
    layer0_outputs(2024) <= a and not b;
    layer0_outputs(2025) <= a;
    layer0_outputs(2026) <= a or b;
    layer0_outputs(2027) <= a or b;
    layer0_outputs(2028) <= not (a or b);
    layer0_outputs(2029) <= b;
    layer0_outputs(2030) <= a or b;
    layer0_outputs(2031) <= a xor b;
    layer0_outputs(2032) <= '1';
    layer0_outputs(2033) <= a;
    layer0_outputs(2034) <= a and not b;
    layer0_outputs(2035) <= a;
    layer0_outputs(2036) <= a;
    layer0_outputs(2037) <= '0';
    layer0_outputs(2038) <= not b;
    layer0_outputs(2039) <= '0';
    layer0_outputs(2040) <= a;
    layer0_outputs(2041) <= not a;
    layer0_outputs(2042) <= not a;
    layer0_outputs(2043) <= '1';
    layer0_outputs(2044) <= not b;
    layer0_outputs(2045) <= not (a or b);
    layer0_outputs(2046) <= not (a xor b);
    layer0_outputs(2047) <= not (a and b);
    layer0_outputs(2048) <= '1';
    layer0_outputs(2049) <= b and not a;
    layer0_outputs(2050) <= a;
    layer0_outputs(2051) <= a xor b;
    layer0_outputs(2052) <= a or b;
    layer0_outputs(2053) <= not b;
    layer0_outputs(2054) <= not a or b;
    layer0_outputs(2055) <= not b;
    layer0_outputs(2056) <= not b;
    layer0_outputs(2057) <= not (a xor b);
    layer0_outputs(2058) <= a or b;
    layer0_outputs(2059) <= a or b;
    layer0_outputs(2060) <= not (a and b);
    layer0_outputs(2061) <= not b;
    layer0_outputs(2062) <= a xor b;
    layer0_outputs(2063) <= not a;
    layer0_outputs(2064) <= a and b;
    layer0_outputs(2065) <= '1';
    layer0_outputs(2066) <= b;
    layer0_outputs(2067) <= not (a or b);
    layer0_outputs(2068) <= not a;
    layer0_outputs(2069) <= not a;
    layer0_outputs(2070) <= not (a or b);
    layer0_outputs(2071) <= a;
    layer0_outputs(2072) <= '1';
    layer0_outputs(2073) <= a and b;
    layer0_outputs(2074) <= '1';
    layer0_outputs(2075) <= a and b;
    layer0_outputs(2076) <= a xor b;
    layer0_outputs(2077) <= not a;
    layer0_outputs(2078) <= not a or b;
    layer0_outputs(2079) <= a;
    layer0_outputs(2080) <= a or b;
    layer0_outputs(2081) <= not b;
    layer0_outputs(2082) <= not (a or b);
    layer0_outputs(2083) <= not (a or b);
    layer0_outputs(2084) <= not a or b;
    layer0_outputs(2085) <= not (a and b);
    layer0_outputs(2086) <= not (a and b);
    layer0_outputs(2087) <= a or b;
    layer0_outputs(2088) <= '1';
    layer0_outputs(2089) <= not (a or b);
    layer0_outputs(2090) <= not a;
    layer0_outputs(2091) <= a xor b;
    layer0_outputs(2092) <= b;
    layer0_outputs(2093) <= '0';
    layer0_outputs(2094) <= a and b;
    layer0_outputs(2095) <= not b or a;
    layer0_outputs(2096) <= '0';
    layer0_outputs(2097) <= '0';
    layer0_outputs(2098) <= not b;
    layer0_outputs(2099) <= b;
    layer0_outputs(2100) <= a xor b;
    layer0_outputs(2101) <= not a;
    layer0_outputs(2102) <= a and b;
    layer0_outputs(2103) <= b and not a;
    layer0_outputs(2104) <= '1';
    layer0_outputs(2105) <= a and not b;
    layer0_outputs(2106) <= not a or b;
    layer0_outputs(2107) <= a;
    layer0_outputs(2108) <= '1';
    layer0_outputs(2109) <= not (a and b);
    layer0_outputs(2110) <= not b or a;
    layer0_outputs(2111) <= '1';
    layer0_outputs(2112) <= not (a and b);
    layer0_outputs(2113) <= not b;
    layer0_outputs(2114) <= '0';
    layer0_outputs(2115) <= a or b;
    layer0_outputs(2116) <= not a;
    layer0_outputs(2117) <= not (a and b);
    layer0_outputs(2118) <= b;
    layer0_outputs(2119) <= a or b;
    layer0_outputs(2120) <= a;
    layer0_outputs(2121) <= a;
    layer0_outputs(2122) <= not (a xor b);
    layer0_outputs(2123) <= '1';
    layer0_outputs(2124) <= a and b;
    layer0_outputs(2125) <= not b;
    layer0_outputs(2126) <= a or b;
    layer0_outputs(2127) <= not b;
    layer0_outputs(2128) <= not (a xor b);
    layer0_outputs(2129) <= not b;
    layer0_outputs(2130) <= '0';
    layer0_outputs(2131) <= b;
    layer0_outputs(2132) <= not (a xor b);
    layer0_outputs(2133) <= a;
    layer0_outputs(2134) <= not a;
    layer0_outputs(2135) <= a and b;
    layer0_outputs(2136) <= not b;
    layer0_outputs(2137) <= b and not a;
    layer0_outputs(2138) <= not b;
    layer0_outputs(2139) <= a and not b;
    layer0_outputs(2140) <= a;
    layer0_outputs(2141) <= b and not a;
    layer0_outputs(2142) <= a and b;
    layer0_outputs(2143) <= not b or a;
    layer0_outputs(2144) <= a or b;
    layer0_outputs(2145) <= a;
    layer0_outputs(2146) <= a and b;
    layer0_outputs(2147) <= '0';
    layer0_outputs(2148) <= '1';
    layer0_outputs(2149) <= a or b;
    layer0_outputs(2150) <= not a;
    layer0_outputs(2151) <= not a;
    layer0_outputs(2152) <= b and not a;
    layer0_outputs(2153) <= not b or a;
    layer0_outputs(2154) <= a and b;
    layer0_outputs(2155) <= not (a or b);
    layer0_outputs(2156) <= '1';
    layer0_outputs(2157) <= not (a xor b);
    layer0_outputs(2158) <= b;
    layer0_outputs(2159) <= not a or b;
    layer0_outputs(2160) <= '1';
    layer0_outputs(2161) <= not a;
    layer0_outputs(2162) <= b;
    layer0_outputs(2163) <= b;
    layer0_outputs(2164) <= a and b;
    layer0_outputs(2165) <= not (a or b);
    layer0_outputs(2166) <= not a;
    layer0_outputs(2167) <= not a;
    layer0_outputs(2168) <= '0';
    layer0_outputs(2169) <= a xor b;
    layer0_outputs(2170) <= '0';
    layer0_outputs(2171) <= a or b;
    layer0_outputs(2172) <= a and not b;
    layer0_outputs(2173) <= not a;
    layer0_outputs(2174) <= b;
    layer0_outputs(2175) <= a and not b;
    layer0_outputs(2176) <= b;
    layer0_outputs(2177) <= b and not a;
    layer0_outputs(2178) <= not b;
    layer0_outputs(2179) <= a xor b;
    layer0_outputs(2180) <= '1';
    layer0_outputs(2181) <= a;
    layer0_outputs(2182) <= not (a or b);
    layer0_outputs(2183) <= not a;
    layer0_outputs(2184) <= b and not a;
    layer0_outputs(2185) <= not b;
    layer0_outputs(2186) <= not b;
    layer0_outputs(2187) <= a and b;
    layer0_outputs(2188) <= not b;
    layer0_outputs(2189) <= a and b;
    layer0_outputs(2190) <= a and not b;
    layer0_outputs(2191) <= not (a xor b);
    layer0_outputs(2192) <= not b;
    layer0_outputs(2193) <= a and b;
    layer0_outputs(2194) <= b and not a;
    layer0_outputs(2195) <= '0';
    layer0_outputs(2196) <= not a;
    layer0_outputs(2197) <= a or b;
    layer0_outputs(2198) <= a and not b;
    layer0_outputs(2199) <= not a or b;
    layer0_outputs(2200) <= a and b;
    layer0_outputs(2201) <= not (a or b);
    layer0_outputs(2202) <= a;
    layer0_outputs(2203) <= a and not b;
    layer0_outputs(2204) <= '0';
    layer0_outputs(2205) <= '0';
    layer0_outputs(2206) <= not (a or b);
    layer0_outputs(2207) <= not (a and b);
    layer0_outputs(2208) <= a and b;
    layer0_outputs(2209) <= not a or b;
    layer0_outputs(2210) <= not a or b;
    layer0_outputs(2211) <= a;
    layer0_outputs(2212) <= a or b;
    layer0_outputs(2213) <= '0';
    layer0_outputs(2214) <= not b;
    layer0_outputs(2215) <= b and not a;
    layer0_outputs(2216) <= a;
    layer0_outputs(2217) <= not (a or b);
    layer0_outputs(2218) <= not b or a;
    layer0_outputs(2219) <= not (a and b);
    layer0_outputs(2220) <= '1';
    layer0_outputs(2221) <= not b;
    layer0_outputs(2222) <= '1';
    layer0_outputs(2223) <= a and b;
    layer0_outputs(2224) <= a and not b;
    layer0_outputs(2225) <= b;
    layer0_outputs(2226) <= not (a or b);
    layer0_outputs(2227) <= a and not b;
    layer0_outputs(2228) <= not a;
    layer0_outputs(2229) <= '1';
    layer0_outputs(2230) <= not b;
    layer0_outputs(2231) <= a and b;
    layer0_outputs(2232) <= not (a xor b);
    layer0_outputs(2233) <= '1';
    layer0_outputs(2234) <= not a;
    layer0_outputs(2235) <= a and b;
    layer0_outputs(2236) <= b;
    layer0_outputs(2237) <= not (a and b);
    layer0_outputs(2238) <= a or b;
    layer0_outputs(2239) <= not (a and b);
    layer0_outputs(2240) <= a or b;
    layer0_outputs(2241) <= not (a and b);
    layer0_outputs(2242) <= not (a or b);
    layer0_outputs(2243) <= '0';
    layer0_outputs(2244) <= a or b;
    layer0_outputs(2245) <= b and not a;
    layer0_outputs(2246) <= not a or b;
    layer0_outputs(2247) <= '1';
    layer0_outputs(2248) <= a;
    layer0_outputs(2249) <= '1';
    layer0_outputs(2250) <= b and not a;
    layer0_outputs(2251) <= not b or a;
    layer0_outputs(2252) <= not b;
    layer0_outputs(2253) <= b;
    layer0_outputs(2254) <= a and b;
    layer0_outputs(2255) <= a and not b;
    layer0_outputs(2256) <= b;
    layer0_outputs(2257) <= '1';
    layer0_outputs(2258) <= '1';
    layer0_outputs(2259) <= a and b;
    layer0_outputs(2260) <= '1';
    layer0_outputs(2261) <= b and not a;
    layer0_outputs(2262) <= b;
    layer0_outputs(2263) <= not b or a;
    layer0_outputs(2264) <= a and not b;
    layer0_outputs(2265) <= not b or a;
    layer0_outputs(2266) <= a xor b;
    layer0_outputs(2267) <= not a;
    layer0_outputs(2268) <= a;
    layer0_outputs(2269) <= a or b;
    layer0_outputs(2270) <= not a;
    layer0_outputs(2271) <= '1';
    layer0_outputs(2272) <= a xor b;
    layer0_outputs(2273) <= b;
    layer0_outputs(2274) <= '1';
    layer0_outputs(2275) <= '0';
    layer0_outputs(2276) <= '1';
    layer0_outputs(2277) <= not (a and b);
    layer0_outputs(2278) <= not (a or b);
    layer0_outputs(2279) <= a;
    layer0_outputs(2280) <= a xor b;
    layer0_outputs(2281) <= not (a xor b);
    layer0_outputs(2282) <= not b;
    layer0_outputs(2283) <= b;
    layer0_outputs(2284) <= not b or a;
    layer0_outputs(2285) <= b;
    layer0_outputs(2286) <= not a;
    layer0_outputs(2287) <= a and b;
    layer0_outputs(2288) <= b;
    layer0_outputs(2289) <= a or b;
    layer0_outputs(2290) <= b and not a;
    layer0_outputs(2291) <= b and not a;
    layer0_outputs(2292) <= not a or b;
    layer0_outputs(2293) <= a xor b;
    layer0_outputs(2294) <= '0';
    layer0_outputs(2295) <= not (a or b);
    layer0_outputs(2296) <= a or b;
    layer0_outputs(2297) <= a and not b;
    layer0_outputs(2298) <= a or b;
    layer0_outputs(2299) <= a and not b;
    layer0_outputs(2300) <= not a or b;
    layer0_outputs(2301) <= b;
    layer0_outputs(2302) <= '0';
    layer0_outputs(2303) <= a;
    layer0_outputs(2304) <= b and not a;
    layer0_outputs(2305) <= not b or a;
    layer0_outputs(2306) <= not a or b;
    layer0_outputs(2307) <= a and not b;
    layer0_outputs(2308) <= not b;
    layer0_outputs(2309) <= not a or b;
    layer0_outputs(2310) <= not (a and b);
    layer0_outputs(2311) <= a and b;
    layer0_outputs(2312) <= not (a or b);
    layer0_outputs(2313) <= not a or b;
    layer0_outputs(2314) <= a;
    layer0_outputs(2315) <= '1';
    layer0_outputs(2316) <= a;
    layer0_outputs(2317) <= '0';
    layer0_outputs(2318) <= a;
    layer0_outputs(2319) <= a and not b;
    layer0_outputs(2320) <= a and b;
    layer0_outputs(2321) <= not (a xor b);
    layer0_outputs(2322) <= b and not a;
    layer0_outputs(2323) <= a;
    layer0_outputs(2324) <= not (a or b);
    layer0_outputs(2325) <= '0';
    layer0_outputs(2326) <= a and not b;
    layer0_outputs(2327) <= not a;
    layer0_outputs(2328) <= a and not b;
    layer0_outputs(2329) <= not a or b;
    layer0_outputs(2330) <= a and not b;
    layer0_outputs(2331) <= a or b;
    layer0_outputs(2332) <= '0';
    layer0_outputs(2333) <= not b or a;
    layer0_outputs(2334) <= a or b;
    layer0_outputs(2335) <= not (a or b);
    layer0_outputs(2336) <= not (a and b);
    layer0_outputs(2337) <= '1';
    layer0_outputs(2338) <= a;
    layer0_outputs(2339) <= '0';
    layer0_outputs(2340) <= '0';
    layer0_outputs(2341) <= '0';
    layer0_outputs(2342) <= not b;
    layer0_outputs(2343) <= a and b;
    layer0_outputs(2344) <= a or b;
    layer0_outputs(2345) <= b;
    layer0_outputs(2346) <= a or b;
    layer0_outputs(2347) <= b;
    layer0_outputs(2348) <= not (a and b);
    layer0_outputs(2349) <= b;
    layer0_outputs(2350) <= not (a and b);
    layer0_outputs(2351) <= a or b;
    layer0_outputs(2352) <= not b;
    layer0_outputs(2353) <= not a or b;
    layer0_outputs(2354) <= '0';
    layer0_outputs(2355) <= '1';
    layer0_outputs(2356) <= not b;
    layer0_outputs(2357) <= not b or a;
    layer0_outputs(2358) <= not a or b;
    layer0_outputs(2359) <= a;
    layer0_outputs(2360) <= a;
    layer0_outputs(2361) <= a or b;
    layer0_outputs(2362) <= not b or a;
    layer0_outputs(2363) <= '1';
    layer0_outputs(2364) <= a xor b;
    layer0_outputs(2365) <= '0';
    layer0_outputs(2366) <= not a;
    layer0_outputs(2367) <= a and b;
    layer0_outputs(2368) <= '1';
    layer0_outputs(2369) <= b and not a;
    layer0_outputs(2370) <= not a or b;
    layer0_outputs(2371) <= not (a xor b);
    layer0_outputs(2372) <= a xor b;
    layer0_outputs(2373) <= not b or a;
    layer0_outputs(2374) <= '1';
    layer0_outputs(2375) <= '1';
    layer0_outputs(2376) <= not (a or b);
    layer0_outputs(2377) <= a and b;
    layer0_outputs(2378) <= a and b;
    layer0_outputs(2379) <= not a;
    layer0_outputs(2380) <= not b;
    layer0_outputs(2381) <= not (a or b);
    layer0_outputs(2382) <= '0';
    layer0_outputs(2383) <= '1';
    layer0_outputs(2384) <= not a;
    layer0_outputs(2385) <= a and b;
    layer0_outputs(2386) <= not (a xor b);
    layer0_outputs(2387) <= a and b;
    layer0_outputs(2388) <= '1';
    layer0_outputs(2389) <= '0';
    layer0_outputs(2390) <= a and b;
    layer0_outputs(2391) <= not a;
    layer0_outputs(2392) <= not (a or b);
    layer0_outputs(2393) <= not a;
    layer0_outputs(2394) <= b and not a;
    layer0_outputs(2395) <= '1';
    layer0_outputs(2396) <= not b or a;
    layer0_outputs(2397) <= not (a or b);
    layer0_outputs(2398) <= not b or a;
    layer0_outputs(2399) <= not a;
    layer0_outputs(2400) <= b;
    layer0_outputs(2401) <= '1';
    layer0_outputs(2402) <= not b;
    layer0_outputs(2403) <= a and not b;
    layer0_outputs(2404) <= a and b;
    layer0_outputs(2405) <= not a or b;
    layer0_outputs(2406) <= not b;
    layer0_outputs(2407) <= a or b;
    layer0_outputs(2408) <= a xor b;
    layer0_outputs(2409) <= a or b;
    layer0_outputs(2410) <= not b;
    layer0_outputs(2411) <= a;
    layer0_outputs(2412) <= b and not a;
    layer0_outputs(2413) <= a or b;
    layer0_outputs(2414) <= a and b;
    layer0_outputs(2415) <= not a;
    layer0_outputs(2416) <= '0';
    layer0_outputs(2417) <= a;
    layer0_outputs(2418) <= not b or a;
    layer0_outputs(2419) <= a or b;
    layer0_outputs(2420) <= a and b;
    layer0_outputs(2421) <= a or b;
    layer0_outputs(2422) <= a and b;
    layer0_outputs(2423) <= not (a or b);
    layer0_outputs(2424) <= b and not a;
    layer0_outputs(2425) <= not b;
    layer0_outputs(2426) <= b;
    layer0_outputs(2427) <= not a or b;
    layer0_outputs(2428) <= not (a or b);
    layer0_outputs(2429) <= a and not b;
    layer0_outputs(2430) <= not a;
    layer0_outputs(2431) <= not (a and b);
    layer0_outputs(2432) <= not (a xor b);
    layer0_outputs(2433) <= b;
    layer0_outputs(2434) <= not a or b;
    layer0_outputs(2435) <= '1';
    layer0_outputs(2436) <= a or b;
    layer0_outputs(2437) <= '1';
    layer0_outputs(2438) <= not (a xor b);
    layer0_outputs(2439) <= a and b;
    layer0_outputs(2440) <= '1';
    layer0_outputs(2441) <= a or b;
    layer0_outputs(2442) <= a and not b;
    layer0_outputs(2443) <= a or b;
    layer0_outputs(2444) <= b and not a;
    layer0_outputs(2445) <= not (a and b);
    layer0_outputs(2446) <= not (a xor b);
    layer0_outputs(2447) <= not (a and b);
    layer0_outputs(2448) <= not a or b;
    layer0_outputs(2449) <= a;
    layer0_outputs(2450) <= '1';
    layer0_outputs(2451) <= a and not b;
    layer0_outputs(2452) <= not a or b;
    layer0_outputs(2453) <= not (a or b);
    layer0_outputs(2454) <= not b;
    layer0_outputs(2455) <= not (a and b);
    layer0_outputs(2456) <= a and b;
    layer0_outputs(2457) <= not b;
    layer0_outputs(2458) <= b;
    layer0_outputs(2459) <= a;
    layer0_outputs(2460) <= not (a and b);
    layer0_outputs(2461) <= not b or a;
    layer0_outputs(2462) <= not a;
    layer0_outputs(2463) <= a;
    layer0_outputs(2464) <= a and b;
    layer0_outputs(2465) <= not (a or b);
    layer0_outputs(2466) <= not (a and b);
    layer0_outputs(2467) <= not (a or b);
    layer0_outputs(2468) <= '0';
    layer0_outputs(2469) <= '0';
    layer0_outputs(2470) <= a and b;
    layer0_outputs(2471) <= '1';
    layer0_outputs(2472) <= b and not a;
    layer0_outputs(2473) <= a;
    layer0_outputs(2474) <= a and not b;
    layer0_outputs(2475) <= not (a or b);
    layer0_outputs(2476) <= not (a and b);
    layer0_outputs(2477) <= a;
    layer0_outputs(2478) <= b;
    layer0_outputs(2479) <= not (a and b);
    layer0_outputs(2480) <= not (a or b);
    layer0_outputs(2481) <= not a or b;
    layer0_outputs(2482) <= not (a or b);
    layer0_outputs(2483) <= '1';
    layer0_outputs(2484) <= a or b;
    layer0_outputs(2485) <= '1';
    layer0_outputs(2486) <= '1';
    layer0_outputs(2487) <= '0';
    layer0_outputs(2488) <= not (a or b);
    layer0_outputs(2489) <= not a or b;
    layer0_outputs(2490) <= a xor b;
    layer0_outputs(2491) <= a and not b;
    layer0_outputs(2492) <= not a or b;
    layer0_outputs(2493) <= not b;
    layer0_outputs(2494) <= a xor b;
    layer0_outputs(2495) <= b and not a;
    layer0_outputs(2496) <= not (a and b);
    layer0_outputs(2497) <= b;
    layer0_outputs(2498) <= a;
    layer0_outputs(2499) <= a or b;
    layer0_outputs(2500) <= not a;
    layer0_outputs(2501) <= '1';
    layer0_outputs(2502) <= not a;
    layer0_outputs(2503) <= '1';
    layer0_outputs(2504) <= a and not b;
    layer0_outputs(2505) <= b;
    layer0_outputs(2506) <= b and not a;
    layer0_outputs(2507) <= not a or b;
    layer0_outputs(2508) <= not (a and b);
    layer0_outputs(2509) <= a;
    layer0_outputs(2510) <= '1';
    layer0_outputs(2511) <= not a or b;
    layer0_outputs(2512) <= '0';
    layer0_outputs(2513) <= a and not b;
    layer0_outputs(2514) <= not (a and b);
    layer0_outputs(2515) <= not (a xor b);
    layer0_outputs(2516) <= a;
    layer0_outputs(2517) <= a or b;
    layer0_outputs(2518) <= a;
    layer0_outputs(2519) <= not b or a;
    layer0_outputs(2520) <= not (a xor b);
    layer0_outputs(2521) <= not (a and b);
    layer0_outputs(2522) <= not b or a;
    layer0_outputs(2523) <= not a or b;
    layer0_outputs(2524) <= '0';
    layer0_outputs(2525) <= '0';
    layer0_outputs(2526) <= b;
    layer0_outputs(2527) <= not b;
    layer0_outputs(2528) <= b and not a;
    layer0_outputs(2529) <= not (a and b);
    layer0_outputs(2530) <= '0';
    layer0_outputs(2531) <= '0';
    layer0_outputs(2532) <= not (a or b);
    layer0_outputs(2533) <= a;
    layer0_outputs(2534) <= b and not a;
    layer0_outputs(2535) <= a xor b;
    layer0_outputs(2536) <= not b;
    layer0_outputs(2537) <= not (a and b);
    layer0_outputs(2538) <= '1';
    layer0_outputs(2539) <= not a;
    layer0_outputs(2540) <= not b or a;
    layer0_outputs(2541) <= not (a xor b);
    layer0_outputs(2542) <= not (a xor b);
    layer0_outputs(2543) <= not a or b;
    layer0_outputs(2544) <= b;
    layer0_outputs(2545) <= not b;
    layer0_outputs(2546) <= not b or a;
    layer0_outputs(2547) <= '1';
    layer0_outputs(2548) <= not b;
    layer0_outputs(2549) <= not b or a;
    layer0_outputs(2550) <= a or b;
    layer0_outputs(2551) <= not (a or b);
    layer0_outputs(2552) <= not b or a;
    layer0_outputs(2553) <= not (a and b);
    layer0_outputs(2554) <= not (a and b);
    layer0_outputs(2555) <= '0';
    layer0_outputs(2556) <= not b or a;
    layer0_outputs(2557) <= not a;
    layer0_outputs(2558) <= not a;
    layer0_outputs(2559) <= a and b;
    layer0_outputs(2560) <= not (a and b);
    layer0_outputs(2561) <= a and b;
    layer0_outputs(2562) <= a and not b;
    layer0_outputs(2563) <= a and not b;
    layer0_outputs(2564) <= not (a and b);
    layer0_outputs(2565) <= a and b;
    layer0_outputs(2566) <= not (a and b);
    layer0_outputs(2567) <= a;
    layer0_outputs(2568) <= a;
    layer0_outputs(2569) <= not b;
    layer0_outputs(2570) <= b and not a;
    layer0_outputs(2571) <= not b or a;
    layer0_outputs(2572) <= a or b;
    layer0_outputs(2573) <= not (a and b);
    layer0_outputs(2574) <= not b;
    layer0_outputs(2575) <= '0';
    layer0_outputs(2576) <= b and not a;
    layer0_outputs(2577) <= a;
    layer0_outputs(2578) <= not a or b;
    layer0_outputs(2579) <= b;
    layer0_outputs(2580) <= not b or a;
    layer0_outputs(2581) <= a and not b;
    layer0_outputs(2582) <= not b;
    layer0_outputs(2583) <= a or b;
    layer0_outputs(2584) <= a;
    layer0_outputs(2585) <= a;
    layer0_outputs(2586) <= a and b;
    layer0_outputs(2587) <= a and b;
    layer0_outputs(2588) <= not (a or b);
    layer0_outputs(2589) <= not (a and b);
    layer0_outputs(2590) <= not a;
    layer0_outputs(2591) <= not b or a;
    layer0_outputs(2592) <= a or b;
    layer0_outputs(2593) <= not (a and b);
    layer0_outputs(2594) <= not a;
    layer0_outputs(2595) <= '0';
    layer0_outputs(2596) <= '0';
    layer0_outputs(2597) <= not (a or b);
    layer0_outputs(2598) <= not a;
    layer0_outputs(2599) <= not a;
    layer0_outputs(2600) <= a and b;
    layer0_outputs(2601) <= a or b;
    layer0_outputs(2602) <= not b;
    layer0_outputs(2603) <= '1';
    layer0_outputs(2604) <= not (a xor b);
    layer0_outputs(2605) <= not a;
    layer0_outputs(2606) <= a or b;
    layer0_outputs(2607) <= not (a and b);
    layer0_outputs(2608) <= not b or a;
    layer0_outputs(2609) <= not a or b;
    layer0_outputs(2610) <= not (a and b);
    layer0_outputs(2611) <= a and b;
    layer0_outputs(2612) <= '0';
    layer0_outputs(2613) <= not b or a;
    layer0_outputs(2614) <= a;
    layer0_outputs(2615) <= a;
    layer0_outputs(2616) <= not a or b;
    layer0_outputs(2617) <= not b or a;
    layer0_outputs(2618) <= not (a or b);
    layer0_outputs(2619) <= not (a and b);
    layer0_outputs(2620) <= '0';
    layer0_outputs(2621) <= '1';
    layer0_outputs(2622) <= a and not b;
    layer0_outputs(2623) <= not a;
    layer0_outputs(2624) <= a and b;
    layer0_outputs(2625) <= b;
    layer0_outputs(2626) <= not a;
    layer0_outputs(2627) <= '1';
    layer0_outputs(2628) <= not a or b;
    layer0_outputs(2629) <= '1';
    layer0_outputs(2630) <= a;
    layer0_outputs(2631) <= '1';
    layer0_outputs(2632) <= a and b;
    layer0_outputs(2633) <= not (a or b);
    layer0_outputs(2634) <= '0';
    layer0_outputs(2635) <= '1';
    layer0_outputs(2636) <= a and b;
    layer0_outputs(2637) <= '1';
    layer0_outputs(2638) <= not (a or b);
    layer0_outputs(2639) <= a or b;
    layer0_outputs(2640) <= a or b;
    layer0_outputs(2641) <= not b or a;
    layer0_outputs(2642) <= not (a or b);
    layer0_outputs(2643) <= not b;
    layer0_outputs(2644) <= a;
    layer0_outputs(2645) <= not b;
    layer0_outputs(2646) <= not (a and b);
    layer0_outputs(2647) <= '1';
    layer0_outputs(2648) <= not b;
    layer0_outputs(2649) <= not (a and b);
    layer0_outputs(2650) <= a xor b;
    layer0_outputs(2651) <= a and b;
    layer0_outputs(2652) <= not b;
    layer0_outputs(2653) <= not a or b;
    layer0_outputs(2654) <= not a;
    layer0_outputs(2655) <= not (a or b);
    layer0_outputs(2656) <= b;
    layer0_outputs(2657) <= not a or b;
    layer0_outputs(2658) <= a or b;
    layer0_outputs(2659) <= not b;
    layer0_outputs(2660) <= '1';
    layer0_outputs(2661) <= a or b;
    layer0_outputs(2662) <= not (a xor b);
    layer0_outputs(2663) <= not b;
    layer0_outputs(2664) <= a or b;
    layer0_outputs(2665) <= not a or b;
    layer0_outputs(2666) <= a;
    layer0_outputs(2667) <= not a;
    layer0_outputs(2668) <= not a;
    layer0_outputs(2669) <= '1';
    layer0_outputs(2670) <= '0';
    layer0_outputs(2671) <= not b;
    layer0_outputs(2672) <= a or b;
    layer0_outputs(2673) <= b;
    layer0_outputs(2674) <= b;
    layer0_outputs(2675) <= b;
    layer0_outputs(2676) <= not b or a;
    layer0_outputs(2677) <= '0';
    layer0_outputs(2678) <= not (a or b);
    layer0_outputs(2679) <= not a;
    layer0_outputs(2680) <= not b;
    layer0_outputs(2681) <= '0';
    layer0_outputs(2682) <= not (a xor b);
    layer0_outputs(2683) <= b;
    layer0_outputs(2684) <= not b or a;
    layer0_outputs(2685) <= not b or a;
    layer0_outputs(2686) <= not a;
    layer0_outputs(2687) <= b;
    layer0_outputs(2688) <= not (a or b);
    layer0_outputs(2689) <= not a;
    layer0_outputs(2690) <= not a or b;
    layer0_outputs(2691) <= not a;
    layer0_outputs(2692) <= not b;
    layer0_outputs(2693) <= a xor b;
    layer0_outputs(2694) <= '1';
    layer0_outputs(2695) <= a and b;
    layer0_outputs(2696) <= b;
    layer0_outputs(2697) <= b;
    layer0_outputs(2698) <= '0';
    layer0_outputs(2699) <= '1';
    layer0_outputs(2700) <= a;
    layer0_outputs(2701) <= not b;
    layer0_outputs(2702) <= not a;
    layer0_outputs(2703) <= b;
    layer0_outputs(2704) <= not (a or b);
    layer0_outputs(2705) <= a;
    layer0_outputs(2706) <= a and not b;
    layer0_outputs(2707) <= a or b;
    layer0_outputs(2708) <= a xor b;
    layer0_outputs(2709) <= not (a and b);
    layer0_outputs(2710) <= '1';
    layer0_outputs(2711) <= a or b;
    layer0_outputs(2712) <= '1';
    layer0_outputs(2713) <= a xor b;
    layer0_outputs(2714) <= not (a and b);
    layer0_outputs(2715) <= '1';
    layer0_outputs(2716) <= not b or a;
    layer0_outputs(2717) <= '0';
    layer0_outputs(2718) <= a;
    layer0_outputs(2719) <= a xor b;
    layer0_outputs(2720) <= '0';
    layer0_outputs(2721) <= a;
    layer0_outputs(2722) <= not a;
    layer0_outputs(2723) <= not b;
    layer0_outputs(2724) <= not b or a;
    layer0_outputs(2725) <= not a;
    layer0_outputs(2726) <= not a;
    layer0_outputs(2727) <= not (a or b);
    layer0_outputs(2728) <= not b or a;
    layer0_outputs(2729) <= a xor b;
    layer0_outputs(2730) <= not a;
    layer0_outputs(2731) <= a;
    layer0_outputs(2732) <= not a or b;
    layer0_outputs(2733) <= '0';
    layer0_outputs(2734) <= not (a and b);
    layer0_outputs(2735) <= not (a xor b);
    layer0_outputs(2736) <= not a;
    layer0_outputs(2737) <= not b or a;
    layer0_outputs(2738) <= not (a xor b);
    layer0_outputs(2739) <= a and not b;
    layer0_outputs(2740) <= not (a or b);
    layer0_outputs(2741) <= a or b;
    layer0_outputs(2742) <= b;
    layer0_outputs(2743) <= a and b;
    layer0_outputs(2744) <= not b;
    layer0_outputs(2745) <= not b;
    layer0_outputs(2746) <= a;
    layer0_outputs(2747) <= b and not a;
    layer0_outputs(2748) <= a and b;
    layer0_outputs(2749) <= b;
    layer0_outputs(2750) <= not a;
    layer0_outputs(2751) <= b;
    layer0_outputs(2752) <= not (a or b);
    layer0_outputs(2753) <= a;
    layer0_outputs(2754) <= a;
    layer0_outputs(2755) <= b and not a;
    layer0_outputs(2756) <= b;
    layer0_outputs(2757) <= not a or b;
    layer0_outputs(2758) <= not (a and b);
    layer0_outputs(2759) <= not a;
    layer0_outputs(2760) <= not b;
    layer0_outputs(2761) <= not (a or b);
    layer0_outputs(2762) <= a or b;
    layer0_outputs(2763) <= a xor b;
    layer0_outputs(2764) <= not (a or b);
    layer0_outputs(2765) <= a;
    layer0_outputs(2766) <= a or b;
    layer0_outputs(2767) <= not (a and b);
    layer0_outputs(2768) <= not b or a;
    layer0_outputs(2769) <= a xor b;
    layer0_outputs(2770) <= not (a and b);
    layer0_outputs(2771) <= not (a and b);
    layer0_outputs(2772) <= b;
    layer0_outputs(2773) <= a or b;
    layer0_outputs(2774) <= '0';
    layer0_outputs(2775) <= not b or a;
    layer0_outputs(2776) <= b and not a;
    layer0_outputs(2777) <= '1';
    layer0_outputs(2778) <= not (a and b);
    layer0_outputs(2779) <= a xor b;
    layer0_outputs(2780) <= not b or a;
    layer0_outputs(2781) <= '1';
    layer0_outputs(2782) <= a;
    layer0_outputs(2783) <= b and not a;
    layer0_outputs(2784) <= not (a and b);
    layer0_outputs(2785) <= a and not b;
    layer0_outputs(2786) <= not (a and b);
    layer0_outputs(2787) <= not (a and b);
    layer0_outputs(2788) <= '1';
    layer0_outputs(2789) <= '0';
    layer0_outputs(2790) <= not b or a;
    layer0_outputs(2791) <= not a;
    layer0_outputs(2792) <= a and b;
    layer0_outputs(2793) <= a and not b;
    layer0_outputs(2794) <= '1';
    layer0_outputs(2795) <= not a;
    layer0_outputs(2796) <= not (a or b);
    layer0_outputs(2797) <= '1';
    layer0_outputs(2798) <= b and not a;
    layer0_outputs(2799) <= '1';
    layer0_outputs(2800) <= not b;
    layer0_outputs(2801) <= a and not b;
    layer0_outputs(2802) <= not b or a;
    layer0_outputs(2803) <= not (a or b);
    layer0_outputs(2804) <= not a;
    layer0_outputs(2805) <= not b;
    layer0_outputs(2806) <= not b or a;
    layer0_outputs(2807) <= not (a xor b);
    layer0_outputs(2808) <= not b or a;
    layer0_outputs(2809) <= a;
    layer0_outputs(2810) <= b;
    layer0_outputs(2811) <= a and b;
    layer0_outputs(2812) <= not a or b;
    layer0_outputs(2813) <= b and not a;
    layer0_outputs(2814) <= '0';
    layer0_outputs(2815) <= not a;
    layer0_outputs(2816) <= a and not b;
    layer0_outputs(2817) <= not b;
    layer0_outputs(2818) <= not (a xor b);
    layer0_outputs(2819) <= b and not a;
    layer0_outputs(2820) <= not b;
    layer0_outputs(2821) <= a;
    layer0_outputs(2822) <= a;
    layer0_outputs(2823) <= b;
    layer0_outputs(2824) <= not a;
    layer0_outputs(2825) <= not (a or b);
    layer0_outputs(2826) <= not (a or b);
    layer0_outputs(2827) <= a and not b;
    layer0_outputs(2828) <= b;
    layer0_outputs(2829) <= not (a and b);
    layer0_outputs(2830) <= not b or a;
    layer0_outputs(2831) <= '0';
    layer0_outputs(2832) <= a;
    layer0_outputs(2833) <= not a or b;
    layer0_outputs(2834) <= '0';
    layer0_outputs(2835) <= a and b;
    layer0_outputs(2836) <= b;
    layer0_outputs(2837) <= not a;
    layer0_outputs(2838) <= not (a and b);
    layer0_outputs(2839) <= not b or a;
    layer0_outputs(2840) <= '0';
    layer0_outputs(2841) <= b;
    layer0_outputs(2842) <= '1';
    layer0_outputs(2843) <= a or b;
    layer0_outputs(2844) <= not (a or b);
    layer0_outputs(2845) <= not b or a;
    layer0_outputs(2846) <= a or b;
    layer0_outputs(2847) <= not (a and b);
    layer0_outputs(2848) <= not (a or b);
    layer0_outputs(2849) <= not a or b;
    layer0_outputs(2850) <= not (a and b);
    layer0_outputs(2851) <= b;
    layer0_outputs(2852) <= not a or b;
    layer0_outputs(2853) <= not (a or b);
    layer0_outputs(2854) <= not a or b;
    layer0_outputs(2855) <= not b;
    layer0_outputs(2856) <= not a;
    layer0_outputs(2857) <= a and b;
    layer0_outputs(2858) <= not b or a;
    layer0_outputs(2859) <= not (a xor b);
    layer0_outputs(2860) <= b and not a;
    layer0_outputs(2861) <= a;
    layer0_outputs(2862) <= b and not a;
    layer0_outputs(2863) <= b;
    layer0_outputs(2864) <= not b;
    layer0_outputs(2865) <= b;
    layer0_outputs(2866) <= not (a and b);
    layer0_outputs(2867) <= not b or a;
    layer0_outputs(2868) <= not a or b;
    layer0_outputs(2869) <= a xor b;
    layer0_outputs(2870) <= not (a xor b);
    layer0_outputs(2871) <= not b;
    layer0_outputs(2872) <= '0';
    layer0_outputs(2873) <= not a;
    layer0_outputs(2874) <= a;
    layer0_outputs(2875) <= not a;
    layer0_outputs(2876) <= not b or a;
    layer0_outputs(2877) <= a and b;
    layer0_outputs(2878) <= a;
    layer0_outputs(2879) <= not a or b;
    layer0_outputs(2880) <= a xor b;
    layer0_outputs(2881) <= a or b;
    layer0_outputs(2882) <= b;
    layer0_outputs(2883) <= a xor b;
    layer0_outputs(2884) <= a or b;
    layer0_outputs(2885) <= a or b;
    layer0_outputs(2886) <= b and not a;
    layer0_outputs(2887) <= a or b;
    layer0_outputs(2888) <= a or b;
    layer0_outputs(2889) <= '1';
    layer0_outputs(2890) <= a;
    layer0_outputs(2891) <= not (a and b);
    layer0_outputs(2892) <= not (a xor b);
    layer0_outputs(2893) <= a or b;
    layer0_outputs(2894) <= a or b;
    layer0_outputs(2895) <= '0';
    layer0_outputs(2896) <= not b or a;
    layer0_outputs(2897) <= '0';
    layer0_outputs(2898) <= not a or b;
    layer0_outputs(2899) <= a;
    layer0_outputs(2900) <= a and b;
    layer0_outputs(2901) <= not (a xor b);
    layer0_outputs(2902) <= a and b;
    layer0_outputs(2903) <= not (a xor b);
    layer0_outputs(2904) <= '0';
    layer0_outputs(2905) <= '0';
    layer0_outputs(2906) <= b and not a;
    layer0_outputs(2907) <= b and not a;
    layer0_outputs(2908) <= not (a or b);
    layer0_outputs(2909) <= not b;
    layer0_outputs(2910) <= a or b;
    layer0_outputs(2911) <= a;
    layer0_outputs(2912) <= '0';
    layer0_outputs(2913) <= not a;
    layer0_outputs(2914) <= a and not b;
    layer0_outputs(2915) <= a or b;
    layer0_outputs(2916) <= not b;
    layer0_outputs(2917) <= not a or b;
    layer0_outputs(2918) <= '1';
    layer0_outputs(2919) <= a and b;
    layer0_outputs(2920) <= not (a and b);
    layer0_outputs(2921) <= not a;
    layer0_outputs(2922) <= not (a and b);
    layer0_outputs(2923) <= '0';
    layer0_outputs(2924) <= not b;
    layer0_outputs(2925) <= not (a xor b);
    layer0_outputs(2926) <= a;
    layer0_outputs(2927) <= a and b;
    layer0_outputs(2928) <= a;
    layer0_outputs(2929) <= a or b;
    layer0_outputs(2930) <= not (a or b);
    layer0_outputs(2931) <= '0';
    layer0_outputs(2932) <= not a;
    layer0_outputs(2933) <= a;
    layer0_outputs(2934) <= '1';
    layer0_outputs(2935) <= not (a or b);
    layer0_outputs(2936) <= a and b;
    layer0_outputs(2937) <= not a;
    layer0_outputs(2938) <= not b or a;
    layer0_outputs(2939) <= not b or a;
    layer0_outputs(2940) <= '0';
    layer0_outputs(2941) <= '0';
    layer0_outputs(2942) <= a and b;
    layer0_outputs(2943) <= not (a or b);
    layer0_outputs(2944) <= b;
    layer0_outputs(2945) <= a xor b;
    layer0_outputs(2946) <= b;
    layer0_outputs(2947) <= '1';
    layer0_outputs(2948) <= b;
    layer0_outputs(2949) <= a;
    layer0_outputs(2950) <= '0';
    layer0_outputs(2951) <= not a or b;
    layer0_outputs(2952) <= a;
    layer0_outputs(2953) <= not a;
    layer0_outputs(2954) <= '0';
    layer0_outputs(2955) <= b and not a;
    layer0_outputs(2956) <= not b or a;
    layer0_outputs(2957) <= not (a or b);
    layer0_outputs(2958) <= b and not a;
    layer0_outputs(2959) <= b and not a;
    layer0_outputs(2960) <= not (a and b);
    layer0_outputs(2961) <= b and not a;
    layer0_outputs(2962) <= not b;
    layer0_outputs(2963) <= not a;
    layer0_outputs(2964) <= a and b;
    layer0_outputs(2965) <= b and not a;
    layer0_outputs(2966) <= not (a or b);
    layer0_outputs(2967) <= not a;
    layer0_outputs(2968) <= not a;
    layer0_outputs(2969) <= '1';
    layer0_outputs(2970) <= not (a or b);
    layer0_outputs(2971) <= '0';
    layer0_outputs(2972) <= b;
    layer0_outputs(2973) <= '0';
    layer0_outputs(2974) <= a and b;
    layer0_outputs(2975) <= b;
    layer0_outputs(2976) <= a xor b;
    layer0_outputs(2977) <= not b or a;
    layer0_outputs(2978) <= a xor b;
    layer0_outputs(2979) <= a;
    layer0_outputs(2980) <= '1';
    layer0_outputs(2981) <= not (a or b);
    layer0_outputs(2982) <= b;
    layer0_outputs(2983) <= a or b;
    layer0_outputs(2984) <= not b or a;
    layer0_outputs(2985) <= not (a and b);
    layer0_outputs(2986) <= not b or a;
    layer0_outputs(2987) <= '1';
    layer0_outputs(2988) <= b;
    layer0_outputs(2989) <= '0';
    layer0_outputs(2990) <= not a or b;
    layer0_outputs(2991) <= '0';
    layer0_outputs(2992) <= '0';
    layer0_outputs(2993) <= '1';
    layer0_outputs(2994) <= not b;
    layer0_outputs(2995) <= '1';
    layer0_outputs(2996) <= a or b;
    layer0_outputs(2997) <= b;
    layer0_outputs(2998) <= not (a xor b);
    layer0_outputs(2999) <= a;
    layer0_outputs(3000) <= a and not b;
    layer0_outputs(3001) <= a and b;
    layer0_outputs(3002) <= not a;
    layer0_outputs(3003) <= not (a and b);
    layer0_outputs(3004) <= not (a and b);
    layer0_outputs(3005) <= '0';
    layer0_outputs(3006) <= a;
    layer0_outputs(3007) <= '0';
    layer0_outputs(3008) <= '1';
    layer0_outputs(3009) <= not b or a;
    layer0_outputs(3010) <= a and b;
    layer0_outputs(3011) <= a and not b;
    layer0_outputs(3012) <= '1';
    layer0_outputs(3013) <= not b;
    layer0_outputs(3014) <= not (a xor b);
    layer0_outputs(3015) <= not (a or b);
    layer0_outputs(3016) <= '0';
    layer0_outputs(3017) <= not a or b;
    layer0_outputs(3018) <= not b;
    layer0_outputs(3019) <= not a;
    layer0_outputs(3020) <= not (a xor b);
    layer0_outputs(3021) <= a and not b;
    layer0_outputs(3022) <= not b;
    layer0_outputs(3023) <= not b;
    layer0_outputs(3024) <= not b or a;
    layer0_outputs(3025) <= '1';
    layer0_outputs(3026) <= a xor b;
    layer0_outputs(3027) <= a;
    layer0_outputs(3028) <= '1';
    layer0_outputs(3029) <= b and not a;
    layer0_outputs(3030) <= a and not b;
    layer0_outputs(3031) <= not a;
    layer0_outputs(3032) <= not (a and b);
    layer0_outputs(3033) <= '1';
    layer0_outputs(3034) <= not a;
    layer0_outputs(3035) <= b and not a;
    layer0_outputs(3036) <= b;
    layer0_outputs(3037) <= not (a or b);
    layer0_outputs(3038) <= not b or a;
    layer0_outputs(3039) <= b and not a;
    layer0_outputs(3040) <= a and not b;
    layer0_outputs(3041) <= a xor b;
    layer0_outputs(3042) <= not b or a;
    layer0_outputs(3043) <= a and not b;
    layer0_outputs(3044) <= b and not a;
    layer0_outputs(3045) <= b and not a;
    layer0_outputs(3046) <= a xor b;
    layer0_outputs(3047) <= not a or b;
    layer0_outputs(3048) <= not a;
    layer0_outputs(3049) <= not a;
    layer0_outputs(3050) <= '1';
    layer0_outputs(3051) <= not b;
    layer0_outputs(3052) <= a and not b;
    layer0_outputs(3053) <= '1';
    layer0_outputs(3054) <= a;
    layer0_outputs(3055) <= a;
    layer0_outputs(3056) <= '0';
    layer0_outputs(3057) <= b and not a;
    layer0_outputs(3058) <= not b;
    layer0_outputs(3059) <= not a;
    layer0_outputs(3060) <= a and not b;
    layer0_outputs(3061) <= a;
    layer0_outputs(3062) <= a or b;
    layer0_outputs(3063) <= '1';
    layer0_outputs(3064) <= not b;
    layer0_outputs(3065) <= b;
    layer0_outputs(3066) <= a or b;
    layer0_outputs(3067) <= '1';
    layer0_outputs(3068) <= not a;
    layer0_outputs(3069) <= '0';
    layer0_outputs(3070) <= '0';
    layer0_outputs(3071) <= a;
    layer0_outputs(3072) <= '0';
    layer0_outputs(3073) <= a and not b;
    layer0_outputs(3074) <= a;
    layer0_outputs(3075) <= not a or b;
    layer0_outputs(3076) <= not a;
    layer0_outputs(3077) <= a;
    layer0_outputs(3078) <= not (a xor b);
    layer0_outputs(3079) <= a and not b;
    layer0_outputs(3080) <= a;
    layer0_outputs(3081) <= a;
    layer0_outputs(3082) <= a and b;
    layer0_outputs(3083) <= '0';
    layer0_outputs(3084) <= not a or b;
    layer0_outputs(3085) <= a and b;
    layer0_outputs(3086) <= '1';
    layer0_outputs(3087) <= '1';
    layer0_outputs(3088) <= a and not b;
    layer0_outputs(3089) <= a and b;
    layer0_outputs(3090) <= a and not b;
    layer0_outputs(3091) <= not b;
    layer0_outputs(3092) <= not (a and b);
    layer0_outputs(3093) <= not a;
    layer0_outputs(3094) <= a xor b;
    layer0_outputs(3095) <= not b;
    layer0_outputs(3096) <= '0';
    layer0_outputs(3097) <= not a or b;
    layer0_outputs(3098) <= not (a or b);
    layer0_outputs(3099) <= not b;
    layer0_outputs(3100) <= a or b;
    layer0_outputs(3101) <= a xor b;
    layer0_outputs(3102) <= not (a and b);
    layer0_outputs(3103) <= '0';
    layer0_outputs(3104) <= not (a or b);
    layer0_outputs(3105) <= not a;
    layer0_outputs(3106) <= b;
    layer0_outputs(3107) <= '0';
    layer0_outputs(3108) <= '1';
    layer0_outputs(3109) <= a and not b;
    layer0_outputs(3110) <= not a or b;
    layer0_outputs(3111) <= a and not b;
    layer0_outputs(3112) <= a;
    layer0_outputs(3113) <= not a or b;
    layer0_outputs(3114) <= '1';
    layer0_outputs(3115) <= a and not b;
    layer0_outputs(3116) <= not (a and b);
    layer0_outputs(3117) <= a and not b;
    layer0_outputs(3118) <= b;
    layer0_outputs(3119) <= not a;
    layer0_outputs(3120) <= not (a or b);
    layer0_outputs(3121) <= not b;
    layer0_outputs(3122) <= not b or a;
    layer0_outputs(3123) <= a and not b;
    layer0_outputs(3124) <= a and b;
    layer0_outputs(3125) <= not b or a;
    layer0_outputs(3126) <= not (a xor b);
    layer0_outputs(3127) <= not a;
    layer0_outputs(3128) <= not (a or b);
    layer0_outputs(3129) <= '0';
    layer0_outputs(3130) <= a xor b;
    layer0_outputs(3131) <= not a;
    layer0_outputs(3132) <= '0';
    layer0_outputs(3133) <= not a;
    layer0_outputs(3134) <= b and not a;
    layer0_outputs(3135) <= not a or b;
    layer0_outputs(3136) <= a or b;
    layer0_outputs(3137) <= '1';
    layer0_outputs(3138) <= b;
    layer0_outputs(3139) <= a or b;
    layer0_outputs(3140) <= a and b;
    layer0_outputs(3141) <= not b or a;
    layer0_outputs(3142) <= not b or a;
    layer0_outputs(3143) <= a xor b;
    layer0_outputs(3144) <= not b;
    layer0_outputs(3145) <= not (a xor b);
    layer0_outputs(3146) <= a;
    layer0_outputs(3147) <= a and b;
    layer0_outputs(3148) <= not (a xor b);
    layer0_outputs(3149) <= '1';
    layer0_outputs(3150) <= not b or a;
    layer0_outputs(3151) <= not b or a;
    layer0_outputs(3152) <= not a;
    layer0_outputs(3153) <= not b;
    layer0_outputs(3154) <= not (a or b);
    layer0_outputs(3155) <= '0';
    layer0_outputs(3156) <= not (a and b);
    layer0_outputs(3157) <= not (a or b);
    layer0_outputs(3158) <= not (a xor b);
    layer0_outputs(3159) <= not b;
    layer0_outputs(3160) <= b and not a;
    layer0_outputs(3161) <= b and not a;
    layer0_outputs(3162) <= '0';
    layer0_outputs(3163) <= b and not a;
    layer0_outputs(3164) <= a and not b;
    layer0_outputs(3165) <= a;
    layer0_outputs(3166) <= not b;
    layer0_outputs(3167) <= '1';
    layer0_outputs(3168) <= b;
    layer0_outputs(3169) <= not b;
    layer0_outputs(3170) <= b and not a;
    layer0_outputs(3171) <= not b;
    layer0_outputs(3172) <= '1';
    layer0_outputs(3173) <= not (a and b);
    layer0_outputs(3174) <= a and not b;
    layer0_outputs(3175) <= a and b;
    layer0_outputs(3176) <= a or b;
    layer0_outputs(3177) <= not (a or b);
    layer0_outputs(3178) <= not a or b;
    layer0_outputs(3179) <= '1';
    layer0_outputs(3180) <= a and b;
    layer0_outputs(3181) <= '1';
    layer0_outputs(3182) <= a;
    layer0_outputs(3183) <= a and b;
    layer0_outputs(3184) <= not (a and b);
    layer0_outputs(3185) <= a and not b;
    layer0_outputs(3186) <= not a;
    layer0_outputs(3187) <= not (a or b);
    layer0_outputs(3188) <= a and not b;
    layer0_outputs(3189) <= b and not a;
    layer0_outputs(3190) <= a xor b;
    layer0_outputs(3191) <= not a;
    layer0_outputs(3192) <= not b or a;
    layer0_outputs(3193) <= '0';
    layer0_outputs(3194) <= '1';
    layer0_outputs(3195) <= b;
    layer0_outputs(3196) <= a;
    layer0_outputs(3197) <= '1';
    layer0_outputs(3198) <= '0';
    layer0_outputs(3199) <= not (a or b);
    layer0_outputs(3200) <= not a or b;
    layer0_outputs(3201) <= a or b;
    layer0_outputs(3202) <= '1';
    layer0_outputs(3203) <= not b or a;
    layer0_outputs(3204) <= not a;
    layer0_outputs(3205) <= a and b;
    layer0_outputs(3206) <= a and not b;
    layer0_outputs(3207) <= '1';
    layer0_outputs(3208) <= not (a xor b);
    layer0_outputs(3209) <= not b;
    layer0_outputs(3210) <= '0';
    layer0_outputs(3211) <= not b;
    layer0_outputs(3212) <= a;
    layer0_outputs(3213) <= '1';
    layer0_outputs(3214) <= a and not b;
    layer0_outputs(3215) <= a and not b;
    layer0_outputs(3216) <= b and not a;
    layer0_outputs(3217) <= not b or a;
    layer0_outputs(3218) <= not (a xor b);
    layer0_outputs(3219) <= not b;
    layer0_outputs(3220) <= a and b;
    layer0_outputs(3221) <= not a or b;
    layer0_outputs(3222) <= a and not b;
    layer0_outputs(3223) <= '1';
    layer0_outputs(3224) <= '0';
    layer0_outputs(3225) <= a or b;
    layer0_outputs(3226) <= a and not b;
    layer0_outputs(3227) <= b;
    layer0_outputs(3228) <= not b;
    layer0_outputs(3229) <= not (a or b);
    layer0_outputs(3230) <= '1';
    layer0_outputs(3231) <= not (a or b);
    layer0_outputs(3232) <= not (a or b);
    layer0_outputs(3233) <= a and b;
    layer0_outputs(3234) <= b and not a;
    layer0_outputs(3235) <= b and not a;
    layer0_outputs(3236) <= a or b;
    layer0_outputs(3237) <= b and not a;
    layer0_outputs(3238) <= not a or b;
    layer0_outputs(3239) <= a;
    layer0_outputs(3240) <= '1';
    layer0_outputs(3241) <= not b or a;
    layer0_outputs(3242) <= a and b;
    layer0_outputs(3243) <= not (a and b);
    layer0_outputs(3244) <= not (a and b);
    layer0_outputs(3245) <= not a;
    layer0_outputs(3246) <= not a or b;
    layer0_outputs(3247) <= '0';
    layer0_outputs(3248) <= not a or b;
    layer0_outputs(3249) <= a or b;
    layer0_outputs(3250) <= not (a and b);
    layer0_outputs(3251) <= a;
    layer0_outputs(3252) <= b and not a;
    layer0_outputs(3253) <= not (a or b);
    layer0_outputs(3254) <= a xor b;
    layer0_outputs(3255) <= '1';
    layer0_outputs(3256) <= b;
    layer0_outputs(3257) <= '0';
    layer0_outputs(3258) <= not (a or b);
    layer0_outputs(3259) <= b and not a;
    layer0_outputs(3260) <= b;
    layer0_outputs(3261) <= b;
    layer0_outputs(3262) <= not (a and b);
    layer0_outputs(3263) <= '0';
    layer0_outputs(3264) <= a and not b;
    layer0_outputs(3265) <= a and not b;
    layer0_outputs(3266) <= not a;
    layer0_outputs(3267) <= not a or b;
    layer0_outputs(3268) <= b;
    layer0_outputs(3269) <= a and not b;
    layer0_outputs(3270) <= b;
    layer0_outputs(3271) <= '1';
    layer0_outputs(3272) <= not b;
    layer0_outputs(3273) <= not (a or b);
    layer0_outputs(3274) <= not a or b;
    layer0_outputs(3275) <= a and not b;
    layer0_outputs(3276) <= '0';
    layer0_outputs(3277) <= not a or b;
    layer0_outputs(3278) <= b and not a;
    layer0_outputs(3279) <= a and not b;
    layer0_outputs(3280) <= b;
    layer0_outputs(3281) <= a xor b;
    layer0_outputs(3282) <= b and not a;
    layer0_outputs(3283) <= not (a or b);
    layer0_outputs(3284) <= b;
    layer0_outputs(3285) <= a xor b;
    layer0_outputs(3286) <= a and b;
    layer0_outputs(3287) <= not b or a;
    layer0_outputs(3288) <= a;
    layer0_outputs(3289) <= not (a or b);
    layer0_outputs(3290) <= a and not b;
    layer0_outputs(3291) <= a or b;
    layer0_outputs(3292) <= b;
    layer0_outputs(3293) <= a;
    layer0_outputs(3294) <= a;
    layer0_outputs(3295) <= not b or a;
    layer0_outputs(3296) <= a xor b;
    layer0_outputs(3297) <= not a;
    layer0_outputs(3298) <= b and not a;
    layer0_outputs(3299) <= not a or b;
    layer0_outputs(3300) <= a or b;
    layer0_outputs(3301) <= '0';
    layer0_outputs(3302) <= not a;
    layer0_outputs(3303) <= not a;
    layer0_outputs(3304) <= b;
    layer0_outputs(3305) <= not (a or b);
    layer0_outputs(3306) <= b and not a;
    layer0_outputs(3307) <= not b or a;
    layer0_outputs(3308) <= a;
    layer0_outputs(3309) <= a and b;
    layer0_outputs(3310) <= not a;
    layer0_outputs(3311) <= not (a xor b);
    layer0_outputs(3312) <= b;
    layer0_outputs(3313) <= b and not a;
    layer0_outputs(3314) <= a;
    layer0_outputs(3315) <= '1';
    layer0_outputs(3316) <= '1';
    layer0_outputs(3317) <= not b;
    layer0_outputs(3318) <= not (a and b);
    layer0_outputs(3319) <= '0';
    layer0_outputs(3320) <= '0';
    layer0_outputs(3321) <= a and b;
    layer0_outputs(3322) <= not (a and b);
    layer0_outputs(3323) <= not (a or b);
    layer0_outputs(3324) <= a xor b;
    layer0_outputs(3325) <= not b;
    layer0_outputs(3326) <= b and not a;
    layer0_outputs(3327) <= b;
    layer0_outputs(3328) <= not b or a;
    layer0_outputs(3329) <= not a or b;
    layer0_outputs(3330) <= '0';
    layer0_outputs(3331) <= not a;
    layer0_outputs(3332) <= '1';
    layer0_outputs(3333) <= '1';
    layer0_outputs(3334) <= not b;
    layer0_outputs(3335) <= '0';
    layer0_outputs(3336) <= not (a or b);
    layer0_outputs(3337) <= not a or b;
    layer0_outputs(3338) <= a or b;
    layer0_outputs(3339) <= b;
    layer0_outputs(3340) <= not a;
    layer0_outputs(3341) <= a and not b;
    layer0_outputs(3342) <= '1';
    layer0_outputs(3343) <= b;
    layer0_outputs(3344) <= '0';
    layer0_outputs(3345) <= not a or b;
    layer0_outputs(3346) <= a and not b;
    layer0_outputs(3347) <= a;
    layer0_outputs(3348) <= not b or a;
    layer0_outputs(3349) <= '0';
    layer0_outputs(3350) <= not a;
    layer0_outputs(3351) <= not b or a;
    layer0_outputs(3352) <= '1';
    layer0_outputs(3353) <= '1';
    layer0_outputs(3354) <= a and not b;
    layer0_outputs(3355) <= not a;
    layer0_outputs(3356) <= not b;
    layer0_outputs(3357) <= a and b;
    layer0_outputs(3358) <= not b;
    layer0_outputs(3359) <= b and not a;
    layer0_outputs(3360) <= not b or a;
    layer0_outputs(3361) <= '0';
    layer0_outputs(3362) <= not (a or b);
    layer0_outputs(3363) <= not a;
    layer0_outputs(3364) <= not (a and b);
    layer0_outputs(3365) <= a and not b;
    layer0_outputs(3366) <= not b or a;
    layer0_outputs(3367) <= b;
    layer0_outputs(3368) <= not (a or b);
    layer0_outputs(3369) <= a and not b;
    layer0_outputs(3370) <= '0';
    layer0_outputs(3371) <= not (a and b);
    layer0_outputs(3372) <= a and not b;
    layer0_outputs(3373) <= not (a or b);
    layer0_outputs(3374) <= not b or a;
    layer0_outputs(3375) <= not a or b;
    layer0_outputs(3376) <= not (a and b);
    layer0_outputs(3377) <= b and not a;
    layer0_outputs(3378) <= a or b;
    layer0_outputs(3379) <= '1';
    layer0_outputs(3380) <= b;
    layer0_outputs(3381) <= not a or b;
    layer0_outputs(3382) <= not a;
    layer0_outputs(3383) <= not (a xor b);
    layer0_outputs(3384) <= a or b;
    layer0_outputs(3385) <= not a or b;
    layer0_outputs(3386) <= '1';
    layer0_outputs(3387) <= '1';
    layer0_outputs(3388) <= not (a and b);
    layer0_outputs(3389) <= a;
    layer0_outputs(3390) <= not (a and b);
    layer0_outputs(3391) <= a xor b;
    layer0_outputs(3392) <= not a;
    layer0_outputs(3393) <= not a;
    layer0_outputs(3394) <= '0';
    layer0_outputs(3395) <= a and not b;
    layer0_outputs(3396) <= '1';
    layer0_outputs(3397) <= '0';
    layer0_outputs(3398) <= '0';
    layer0_outputs(3399) <= a and not b;
    layer0_outputs(3400) <= not a or b;
    layer0_outputs(3401) <= '0';
    layer0_outputs(3402) <= b;
    layer0_outputs(3403) <= b;
    layer0_outputs(3404) <= not b;
    layer0_outputs(3405) <= '1';
    layer0_outputs(3406) <= b;
    layer0_outputs(3407) <= a and not b;
    layer0_outputs(3408) <= not b or a;
    layer0_outputs(3409) <= not (a xor b);
    layer0_outputs(3410) <= not b or a;
    layer0_outputs(3411) <= a or b;
    layer0_outputs(3412) <= not b or a;
    layer0_outputs(3413) <= b;
    layer0_outputs(3414) <= not b;
    layer0_outputs(3415) <= '1';
    layer0_outputs(3416) <= not b or a;
    layer0_outputs(3417) <= a;
    layer0_outputs(3418) <= a;
    layer0_outputs(3419) <= b and not a;
    layer0_outputs(3420) <= not (a and b);
    layer0_outputs(3421) <= not b or a;
    layer0_outputs(3422) <= b and not a;
    layer0_outputs(3423) <= b and not a;
    layer0_outputs(3424) <= not (a and b);
    layer0_outputs(3425) <= a;
    layer0_outputs(3426) <= '0';
    layer0_outputs(3427) <= a;
    layer0_outputs(3428) <= '1';
    layer0_outputs(3429) <= a and b;
    layer0_outputs(3430) <= not b;
    layer0_outputs(3431) <= not b;
    layer0_outputs(3432) <= not a or b;
    layer0_outputs(3433) <= '1';
    layer0_outputs(3434) <= a and not b;
    layer0_outputs(3435) <= b and not a;
    layer0_outputs(3436) <= a and b;
    layer0_outputs(3437) <= not (a or b);
    layer0_outputs(3438) <= not (a xor b);
    layer0_outputs(3439) <= '0';
    layer0_outputs(3440) <= a and not b;
    layer0_outputs(3441) <= not (a or b);
    layer0_outputs(3442) <= not b or a;
    layer0_outputs(3443) <= b;
    layer0_outputs(3444) <= '1';
    layer0_outputs(3445) <= not (a or b);
    layer0_outputs(3446) <= not (a or b);
    layer0_outputs(3447) <= not a or b;
    layer0_outputs(3448) <= '0';
    layer0_outputs(3449) <= not b;
    layer0_outputs(3450) <= b;
    layer0_outputs(3451) <= a or b;
    layer0_outputs(3452) <= not (a xor b);
    layer0_outputs(3453) <= a and b;
    layer0_outputs(3454) <= a or b;
    layer0_outputs(3455) <= '0';
    layer0_outputs(3456) <= b;
    layer0_outputs(3457) <= a and not b;
    layer0_outputs(3458) <= not b or a;
    layer0_outputs(3459) <= a and b;
    layer0_outputs(3460) <= b;
    layer0_outputs(3461) <= not (a or b);
    layer0_outputs(3462) <= not (a xor b);
    layer0_outputs(3463) <= not (a and b);
    layer0_outputs(3464) <= a or b;
    layer0_outputs(3465) <= not b or a;
    layer0_outputs(3466) <= '0';
    layer0_outputs(3467) <= not (a and b);
    layer0_outputs(3468) <= not b;
    layer0_outputs(3469) <= not a;
    layer0_outputs(3470) <= not b;
    layer0_outputs(3471) <= not a or b;
    layer0_outputs(3472) <= not (a or b);
    layer0_outputs(3473) <= a;
    layer0_outputs(3474) <= a xor b;
    layer0_outputs(3475) <= '1';
    layer0_outputs(3476) <= not (a xor b);
    layer0_outputs(3477) <= not a or b;
    layer0_outputs(3478) <= a xor b;
    layer0_outputs(3479) <= '1';
    layer0_outputs(3480) <= not b or a;
    layer0_outputs(3481) <= a and b;
    layer0_outputs(3482) <= not a;
    layer0_outputs(3483) <= b;
    layer0_outputs(3484) <= not (a xor b);
    layer0_outputs(3485) <= not b;
    layer0_outputs(3486) <= a and not b;
    layer0_outputs(3487) <= '0';
    layer0_outputs(3488) <= '0';
    layer0_outputs(3489) <= b;
    layer0_outputs(3490) <= a or b;
    layer0_outputs(3491) <= b and not a;
    layer0_outputs(3492) <= not b;
    layer0_outputs(3493) <= not a;
    layer0_outputs(3494) <= a or b;
    layer0_outputs(3495) <= a;
    layer0_outputs(3496) <= not a or b;
    layer0_outputs(3497) <= b and not a;
    layer0_outputs(3498) <= a or b;
    layer0_outputs(3499) <= '0';
    layer0_outputs(3500) <= not a or b;
    layer0_outputs(3501) <= '0';
    layer0_outputs(3502) <= '0';
    layer0_outputs(3503) <= a and not b;
    layer0_outputs(3504) <= b;
    layer0_outputs(3505) <= b;
    layer0_outputs(3506) <= a;
    layer0_outputs(3507) <= a and not b;
    layer0_outputs(3508) <= not b or a;
    layer0_outputs(3509) <= b;
    layer0_outputs(3510) <= a or b;
    layer0_outputs(3511) <= a or b;
    layer0_outputs(3512) <= '1';
    layer0_outputs(3513) <= a or b;
    layer0_outputs(3514) <= b;
    layer0_outputs(3515) <= '0';
    layer0_outputs(3516) <= '1';
    layer0_outputs(3517) <= '1';
    layer0_outputs(3518) <= '0';
    layer0_outputs(3519) <= b and not a;
    layer0_outputs(3520) <= '1';
    layer0_outputs(3521) <= a and not b;
    layer0_outputs(3522) <= not a;
    layer0_outputs(3523) <= '0';
    layer0_outputs(3524) <= a;
    layer0_outputs(3525) <= a;
    layer0_outputs(3526) <= a and not b;
    layer0_outputs(3527) <= a and not b;
    layer0_outputs(3528) <= '1';
    layer0_outputs(3529) <= a;
    layer0_outputs(3530) <= not b or a;
    layer0_outputs(3531) <= a and not b;
    layer0_outputs(3532) <= not a or b;
    layer0_outputs(3533) <= not (a and b);
    layer0_outputs(3534) <= not b;
    layer0_outputs(3535) <= not (a or b);
    layer0_outputs(3536) <= not (a xor b);
    layer0_outputs(3537) <= a and not b;
    layer0_outputs(3538) <= a xor b;
    layer0_outputs(3539) <= '1';
    layer0_outputs(3540) <= b;
    layer0_outputs(3541) <= not b;
    layer0_outputs(3542) <= not (a or b);
    layer0_outputs(3543) <= '0';
    layer0_outputs(3544) <= not a or b;
    layer0_outputs(3545) <= '1';
    layer0_outputs(3546) <= not a or b;
    layer0_outputs(3547) <= not (a or b);
    layer0_outputs(3548) <= b;
    layer0_outputs(3549) <= not (a and b);
    layer0_outputs(3550) <= a;
    layer0_outputs(3551) <= not a;
    layer0_outputs(3552) <= '0';
    layer0_outputs(3553) <= a and not b;
    layer0_outputs(3554) <= not (a and b);
    layer0_outputs(3555) <= not a or b;
    layer0_outputs(3556) <= a;
    layer0_outputs(3557) <= a and not b;
    layer0_outputs(3558) <= a and b;
    layer0_outputs(3559) <= a and b;
    layer0_outputs(3560) <= not (a and b);
    layer0_outputs(3561) <= '0';
    layer0_outputs(3562) <= a;
    layer0_outputs(3563) <= not (a and b);
    layer0_outputs(3564) <= not (a or b);
    layer0_outputs(3565) <= b and not a;
    layer0_outputs(3566) <= b;
    layer0_outputs(3567) <= a and b;
    layer0_outputs(3568) <= '1';
    layer0_outputs(3569) <= not (a or b);
    layer0_outputs(3570) <= not (a or b);
    layer0_outputs(3571) <= not b or a;
    layer0_outputs(3572) <= a xor b;
    layer0_outputs(3573) <= '1';
    layer0_outputs(3574) <= not (a xor b);
    layer0_outputs(3575) <= b and not a;
    layer0_outputs(3576) <= not b or a;
    layer0_outputs(3577) <= not b or a;
    layer0_outputs(3578) <= a and b;
    layer0_outputs(3579) <= not (a and b);
    layer0_outputs(3580) <= a and b;
    layer0_outputs(3581) <= b and not a;
    layer0_outputs(3582) <= '1';
    layer0_outputs(3583) <= '0';
    layer0_outputs(3584) <= a;
    layer0_outputs(3585) <= not a;
    layer0_outputs(3586) <= not (a xor b);
    layer0_outputs(3587) <= not b;
    layer0_outputs(3588) <= b and not a;
    layer0_outputs(3589) <= b;
    layer0_outputs(3590) <= not (a and b);
    layer0_outputs(3591) <= a and b;
    layer0_outputs(3592) <= not (a and b);
    layer0_outputs(3593) <= a and not b;
    layer0_outputs(3594) <= b and not a;
    layer0_outputs(3595) <= '1';
    layer0_outputs(3596) <= '0';
    layer0_outputs(3597) <= '1';
    layer0_outputs(3598) <= a and not b;
    layer0_outputs(3599) <= not b;
    layer0_outputs(3600) <= not b or a;
    layer0_outputs(3601) <= a;
    layer0_outputs(3602) <= not b;
    layer0_outputs(3603) <= b;
    layer0_outputs(3604) <= '1';
    layer0_outputs(3605) <= not (a xor b);
    layer0_outputs(3606) <= '1';
    layer0_outputs(3607) <= not (a or b);
    layer0_outputs(3608) <= a or b;
    layer0_outputs(3609) <= b and not a;
    layer0_outputs(3610) <= b and not a;
    layer0_outputs(3611) <= not (a or b);
    layer0_outputs(3612) <= a and b;
    layer0_outputs(3613) <= not (a xor b);
    layer0_outputs(3614) <= '0';
    layer0_outputs(3615) <= not (a or b);
    layer0_outputs(3616) <= not (a xor b);
    layer0_outputs(3617) <= '1';
    layer0_outputs(3618) <= '0';
    layer0_outputs(3619) <= not (a xor b);
    layer0_outputs(3620) <= a and b;
    layer0_outputs(3621) <= not (a or b);
    layer0_outputs(3622) <= a or b;
    layer0_outputs(3623) <= a;
    layer0_outputs(3624) <= '1';
    layer0_outputs(3625) <= a;
    layer0_outputs(3626) <= b and not a;
    layer0_outputs(3627) <= b;
    layer0_outputs(3628) <= not (a and b);
    layer0_outputs(3629) <= b and not a;
    layer0_outputs(3630) <= not a or b;
    layer0_outputs(3631) <= not a;
    layer0_outputs(3632) <= not b;
    layer0_outputs(3633) <= a;
    layer0_outputs(3634) <= not a;
    layer0_outputs(3635) <= not b or a;
    layer0_outputs(3636) <= not b or a;
    layer0_outputs(3637) <= not b or a;
    layer0_outputs(3638) <= not b or a;
    layer0_outputs(3639) <= a or b;
    layer0_outputs(3640) <= a and b;
    layer0_outputs(3641) <= a;
    layer0_outputs(3642) <= a;
    layer0_outputs(3643) <= a and not b;
    layer0_outputs(3644) <= b;
    layer0_outputs(3645) <= '0';
    layer0_outputs(3646) <= b;
    layer0_outputs(3647) <= b and not a;
    layer0_outputs(3648) <= a xor b;
    layer0_outputs(3649) <= a and not b;
    layer0_outputs(3650) <= b;
    layer0_outputs(3651) <= a or b;
    layer0_outputs(3652) <= '1';
    layer0_outputs(3653) <= '0';
    layer0_outputs(3654) <= '1';
    layer0_outputs(3655) <= a and not b;
    layer0_outputs(3656) <= not b;
    layer0_outputs(3657) <= not (a or b);
    layer0_outputs(3658) <= not (a xor b);
    layer0_outputs(3659) <= '0';
    layer0_outputs(3660) <= a and not b;
    layer0_outputs(3661) <= a and not b;
    layer0_outputs(3662) <= not b or a;
    layer0_outputs(3663) <= '1';
    layer0_outputs(3664) <= not (a and b);
    layer0_outputs(3665) <= not (a and b);
    layer0_outputs(3666) <= a and b;
    layer0_outputs(3667) <= not (a xor b);
    layer0_outputs(3668) <= a;
    layer0_outputs(3669) <= not (a and b);
    layer0_outputs(3670) <= not a or b;
    layer0_outputs(3671) <= '1';
    layer0_outputs(3672) <= a;
    layer0_outputs(3673) <= not a or b;
    layer0_outputs(3674) <= not a or b;
    layer0_outputs(3675) <= a;
    layer0_outputs(3676) <= a and b;
    layer0_outputs(3677) <= not a;
    layer0_outputs(3678) <= '1';
    layer0_outputs(3679) <= a and not b;
    layer0_outputs(3680) <= not b;
    layer0_outputs(3681) <= not (a xor b);
    layer0_outputs(3682) <= not (a xor b);
    layer0_outputs(3683) <= not b;
    layer0_outputs(3684) <= a xor b;
    layer0_outputs(3685) <= not (a and b);
    layer0_outputs(3686) <= not b;
    layer0_outputs(3687) <= a xor b;
    layer0_outputs(3688) <= a xor b;
    layer0_outputs(3689) <= a or b;
    layer0_outputs(3690) <= a;
    layer0_outputs(3691) <= a and not b;
    layer0_outputs(3692) <= a or b;
    layer0_outputs(3693) <= not (a or b);
    layer0_outputs(3694) <= not (a or b);
    layer0_outputs(3695) <= b;
    layer0_outputs(3696) <= a;
    layer0_outputs(3697) <= b and not a;
    layer0_outputs(3698) <= '0';
    layer0_outputs(3699) <= a xor b;
    layer0_outputs(3700) <= b;
    layer0_outputs(3701) <= not b;
    layer0_outputs(3702) <= not a;
    layer0_outputs(3703) <= not (a or b);
    layer0_outputs(3704) <= not (a and b);
    layer0_outputs(3705) <= a or b;
    layer0_outputs(3706) <= a xor b;
    layer0_outputs(3707) <= '0';
    layer0_outputs(3708) <= '0';
    layer0_outputs(3709) <= '0';
    layer0_outputs(3710) <= b;
    layer0_outputs(3711) <= not (a xor b);
    layer0_outputs(3712) <= a or b;
    layer0_outputs(3713) <= not b or a;
    layer0_outputs(3714) <= a;
    layer0_outputs(3715) <= not (a and b);
    layer0_outputs(3716) <= not a;
    layer0_outputs(3717) <= b;
    layer0_outputs(3718) <= '0';
    layer0_outputs(3719) <= a or b;
    layer0_outputs(3720) <= a;
    layer0_outputs(3721) <= not b;
    layer0_outputs(3722) <= a and not b;
    layer0_outputs(3723) <= not b or a;
    layer0_outputs(3724) <= a and b;
    layer0_outputs(3725) <= a xor b;
    layer0_outputs(3726) <= a and b;
    layer0_outputs(3727) <= a and b;
    layer0_outputs(3728) <= a and b;
    layer0_outputs(3729) <= b and not a;
    layer0_outputs(3730) <= b and not a;
    layer0_outputs(3731) <= a and b;
    layer0_outputs(3732) <= not (a or b);
    layer0_outputs(3733) <= not b or a;
    layer0_outputs(3734) <= '0';
    layer0_outputs(3735) <= '1';
    layer0_outputs(3736) <= not (a or b);
    layer0_outputs(3737) <= '0';
    layer0_outputs(3738) <= '0';
    layer0_outputs(3739) <= '1';
    layer0_outputs(3740) <= a xor b;
    layer0_outputs(3741) <= not b or a;
    layer0_outputs(3742) <= not b;
    layer0_outputs(3743) <= a and b;
    layer0_outputs(3744) <= a;
    layer0_outputs(3745) <= '1';
    layer0_outputs(3746) <= a and not b;
    layer0_outputs(3747) <= not b;
    layer0_outputs(3748) <= not b or a;
    layer0_outputs(3749) <= a or b;
    layer0_outputs(3750) <= not b or a;
    layer0_outputs(3751) <= '1';
    layer0_outputs(3752) <= a and b;
    layer0_outputs(3753) <= not (a and b);
    layer0_outputs(3754) <= b and not a;
    layer0_outputs(3755) <= not b or a;
    layer0_outputs(3756) <= not a;
    layer0_outputs(3757) <= a xor b;
    layer0_outputs(3758) <= not (a or b);
    layer0_outputs(3759) <= '1';
    layer0_outputs(3760) <= not b or a;
    layer0_outputs(3761) <= b and not a;
    layer0_outputs(3762) <= b;
    layer0_outputs(3763) <= a and b;
    layer0_outputs(3764) <= not b or a;
    layer0_outputs(3765) <= not (a or b);
    layer0_outputs(3766) <= not a;
    layer0_outputs(3767) <= a or b;
    layer0_outputs(3768) <= not b or a;
    layer0_outputs(3769) <= not (a and b);
    layer0_outputs(3770) <= a;
    layer0_outputs(3771) <= not b;
    layer0_outputs(3772) <= a xor b;
    layer0_outputs(3773) <= a;
    layer0_outputs(3774) <= a or b;
    layer0_outputs(3775) <= not b;
    layer0_outputs(3776) <= a and not b;
    layer0_outputs(3777) <= not a or b;
    layer0_outputs(3778) <= '1';
    layer0_outputs(3779) <= a and not b;
    layer0_outputs(3780) <= not b or a;
    layer0_outputs(3781) <= not (a or b);
    layer0_outputs(3782) <= a or b;
    layer0_outputs(3783) <= a and not b;
    layer0_outputs(3784) <= '0';
    layer0_outputs(3785) <= not (a or b);
    layer0_outputs(3786) <= not (a and b);
    layer0_outputs(3787) <= a;
    layer0_outputs(3788) <= not (a or b);
    layer0_outputs(3789) <= a and b;
    layer0_outputs(3790) <= b;
    layer0_outputs(3791) <= '1';
    layer0_outputs(3792) <= b;
    layer0_outputs(3793) <= a xor b;
    layer0_outputs(3794) <= a xor b;
    layer0_outputs(3795) <= not a or b;
    layer0_outputs(3796) <= not a or b;
    layer0_outputs(3797) <= b;
    layer0_outputs(3798) <= a and b;
    layer0_outputs(3799) <= a and b;
    layer0_outputs(3800) <= not b;
    layer0_outputs(3801) <= a or b;
    layer0_outputs(3802) <= not b;
    layer0_outputs(3803) <= a xor b;
    layer0_outputs(3804) <= b and not a;
    layer0_outputs(3805) <= not b;
    layer0_outputs(3806) <= not b;
    layer0_outputs(3807) <= a and b;
    layer0_outputs(3808) <= '0';
    layer0_outputs(3809) <= a xor b;
    layer0_outputs(3810) <= b and not a;
    layer0_outputs(3811) <= not (a or b);
    layer0_outputs(3812) <= a or b;
    layer0_outputs(3813) <= b and not a;
    layer0_outputs(3814) <= a or b;
    layer0_outputs(3815) <= a or b;
    layer0_outputs(3816) <= not b;
    layer0_outputs(3817) <= '0';
    layer0_outputs(3818) <= b and not a;
    layer0_outputs(3819) <= b;
    layer0_outputs(3820) <= not b;
    layer0_outputs(3821) <= not (a or b);
    layer0_outputs(3822) <= not (a and b);
    layer0_outputs(3823) <= '1';
    layer0_outputs(3824) <= '0';
    layer0_outputs(3825) <= '1';
    layer0_outputs(3826) <= b;
    layer0_outputs(3827) <= a or b;
    layer0_outputs(3828) <= b;
    layer0_outputs(3829) <= '0';
    layer0_outputs(3830) <= '1';
    layer0_outputs(3831) <= a and not b;
    layer0_outputs(3832) <= not (a or b);
    layer0_outputs(3833) <= '1';
    layer0_outputs(3834) <= '1';
    layer0_outputs(3835) <= a;
    layer0_outputs(3836) <= not b;
    layer0_outputs(3837) <= a and b;
    layer0_outputs(3838) <= a;
    layer0_outputs(3839) <= a and not b;
    layer0_outputs(3840) <= not (a xor b);
    layer0_outputs(3841) <= not (a and b);
    layer0_outputs(3842) <= not (a or b);
    layer0_outputs(3843) <= not a or b;
    layer0_outputs(3844) <= not (a and b);
    layer0_outputs(3845) <= a;
    layer0_outputs(3846) <= not b;
    layer0_outputs(3847) <= not (a or b);
    layer0_outputs(3848) <= '1';
    layer0_outputs(3849) <= a;
    layer0_outputs(3850) <= not b;
    layer0_outputs(3851) <= a and b;
    layer0_outputs(3852) <= not b or a;
    layer0_outputs(3853) <= '1';
    layer0_outputs(3854) <= b;
    layer0_outputs(3855) <= a and not b;
    layer0_outputs(3856) <= '1';
    layer0_outputs(3857) <= not (a and b);
    layer0_outputs(3858) <= not a or b;
    layer0_outputs(3859) <= not (a and b);
    layer0_outputs(3860) <= a;
    layer0_outputs(3861) <= not (a xor b);
    layer0_outputs(3862) <= '0';
    layer0_outputs(3863) <= not a or b;
    layer0_outputs(3864) <= '0';
    layer0_outputs(3865) <= not b or a;
    layer0_outputs(3866) <= not b or a;
    layer0_outputs(3867) <= a;
    layer0_outputs(3868) <= not a or b;
    layer0_outputs(3869) <= b;
    layer0_outputs(3870) <= a;
    layer0_outputs(3871) <= not (a or b);
    layer0_outputs(3872) <= a or b;
    layer0_outputs(3873) <= not (a and b);
    layer0_outputs(3874) <= not (a xor b);
    layer0_outputs(3875) <= a or b;
    layer0_outputs(3876) <= not a;
    layer0_outputs(3877) <= a xor b;
    layer0_outputs(3878) <= not (a or b);
    layer0_outputs(3879) <= not b or a;
    layer0_outputs(3880) <= b and not a;
    layer0_outputs(3881) <= not a;
    layer0_outputs(3882) <= a and b;
    layer0_outputs(3883) <= '1';
    layer0_outputs(3884) <= not b or a;
    layer0_outputs(3885) <= a and not b;
    layer0_outputs(3886) <= not b;
    layer0_outputs(3887) <= not (a or b);
    layer0_outputs(3888) <= not b or a;
    layer0_outputs(3889) <= a or b;
    layer0_outputs(3890) <= not b or a;
    layer0_outputs(3891) <= not (a or b);
    layer0_outputs(3892) <= not b or a;
    layer0_outputs(3893) <= a;
    layer0_outputs(3894) <= a xor b;
    layer0_outputs(3895) <= a;
    layer0_outputs(3896) <= b and not a;
    layer0_outputs(3897) <= '1';
    layer0_outputs(3898) <= not b;
    layer0_outputs(3899) <= not a or b;
    layer0_outputs(3900) <= a or b;
    layer0_outputs(3901) <= a;
    layer0_outputs(3902) <= not a;
    layer0_outputs(3903) <= a or b;
    layer0_outputs(3904) <= not (a or b);
    layer0_outputs(3905) <= b;
    layer0_outputs(3906) <= not (a or b);
    layer0_outputs(3907) <= a;
    layer0_outputs(3908) <= not b;
    layer0_outputs(3909) <= '1';
    layer0_outputs(3910) <= a and b;
    layer0_outputs(3911) <= not a;
    layer0_outputs(3912) <= not a;
    layer0_outputs(3913) <= not (a and b);
    layer0_outputs(3914) <= a and b;
    layer0_outputs(3915) <= '1';
    layer0_outputs(3916) <= '1';
    layer0_outputs(3917) <= not a or b;
    layer0_outputs(3918) <= a;
    layer0_outputs(3919) <= not (a xor b);
    layer0_outputs(3920) <= '1';
    layer0_outputs(3921) <= not a;
    layer0_outputs(3922) <= b;
    layer0_outputs(3923) <= a and not b;
    layer0_outputs(3924) <= not (a or b);
    layer0_outputs(3925) <= a and b;
    layer0_outputs(3926) <= '0';
    layer0_outputs(3927) <= b and not a;
    layer0_outputs(3928) <= b and not a;
    layer0_outputs(3929) <= b;
    layer0_outputs(3930) <= not b;
    layer0_outputs(3931) <= '1';
    layer0_outputs(3932) <= not b;
    layer0_outputs(3933) <= not (a or b);
    layer0_outputs(3934) <= '1';
    layer0_outputs(3935) <= '0';
    layer0_outputs(3936) <= a and not b;
    layer0_outputs(3937) <= not a;
    layer0_outputs(3938) <= not b;
    layer0_outputs(3939) <= not b;
    layer0_outputs(3940) <= not a or b;
    layer0_outputs(3941) <= not a or b;
    layer0_outputs(3942) <= '1';
    layer0_outputs(3943) <= not (a or b);
    layer0_outputs(3944) <= a;
    layer0_outputs(3945) <= a;
    layer0_outputs(3946) <= not (a or b);
    layer0_outputs(3947) <= not b or a;
    layer0_outputs(3948) <= not (a or b);
    layer0_outputs(3949) <= a and b;
    layer0_outputs(3950) <= a and not b;
    layer0_outputs(3951) <= not (a xor b);
    layer0_outputs(3952) <= not b or a;
    layer0_outputs(3953) <= not (a or b);
    layer0_outputs(3954) <= not (a or b);
    layer0_outputs(3955) <= a and not b;
    layer0_outputs(3956) <= not a or b;
    layer0_outputs(3957) <= a or b;
    layer0_outputs(3958) <= a;
    layer0_outputs(3959) <= '0';
    layer0_outputs(3960) <= not b;
    layer0_outputs(3961) <= not b or a;
    layer0_outputs(3962) <= not a or b;
    layer0_outputs(3963) <= b and not a;
    layer0_outputs(3964) <= not a;
    layer0_outputs(3965) <= a and b;
    layer0_outputs(3966) <= '0';
    layer0_outputs(3967) <= not (a xor b);
    layer0_outputs(3968) <= not b;
    layer0_outputs(3969) <= '1';
    layer0_outputs(3970) <= not a or b;
    layer0_outputs(3971) <= not a or b;
    layer0_outputs(3972) <= a xor b;
    layer0_outputs(3973) <= a or b;
    layer0_outputs(3974) <= not (a or b);
    layer0_outputs(3975) <= a;
    layer0_outputs(3976) <= not (a and b);
    layer0_outputs(3977) <= not b or a;
    layer0_outputs(3978) <= b and not a;
    layer0_outputs(3979) <= not (a or b);
    layer0_outputs(3980) <= a;
    layer0_outputs(3981) <= not (a xor b);
    layer0_outputs(3982) <= not (a and b);
    layer0_outputs(3983) <= a;
    layer0_outputs(3984) <= '0';
    layer0_outputs(3985) <= not (a and b);
    layer0_outputs(3986) <= not a;
    layer0_outputs(3987) <= a;
    layer0_outputs(3988) <= b and not a;
    layer0_outputs(3989) <= not a or b;
    layer0_outputs(3990) <= b;
    layer0_outputs(3991) <= not (a and b);
    layer0_outputs(3992) <= a and b;
    layer0_outputs(3993) <= a;
    layer0_outputs(3994) <= not b;
    layer0_outputs(3995) <= not (a xor b);
    layer0_outputs(3996) <= b and not a;
    layer0_outputs(3997) <= not a or b;
    layer0_outputs(3998) <= not a or b;
    layer0_outputs(3999) <= not a;
    layer0_outputs(4000) <= a and not b;
    layer0_outputs(4001) <= not (a and b);
    layer0_outputs(4002) <= not a;
    layer0_outputs(4003) <= a;
    layer0_outputs(4004) <= a;
    layer0_outputs(4005) <= not (a or b);
    layer0_outputs(4006) <= '0';
    layer0_outputs(4007) <= not b or a;
    layer0_outputs(4008) <= b;
    layer0_outputs(4009) <= not (a and b);
    layer0_outputs(4010) <= a;
    layer0_outputs(4011) <= b and not a;
    layer0_outputs(4012) <= a or b;
    layer0_outputs(4013) <= a or b;
    layer0_outputs(4014) <= not a or b;
    layer0_outputs(4015) <= a and not b;
    layer0_outputs(4016) <= not (a and b);
    layer0_outputs(4017) <= '1';
    layer0_outputs(4018) <= a or b;
    layer0_outputs(4019) <= a and not b;
    layer0_outputs(4020) <= a or b;
    layer0_outputs(4021) <= not (a and b);
    layer0_outputs(4022) <= not b;
    layer0_outputs(4023) <= not b;
    layer0_outputs(4024) <= not b or a;
    layer0_outputs(4025) <= a xor b;
    layer0_outputs(4026) <= not b or a;
    layer0_outputs(4027) <= b;
    layer0_outputs(4028) <= not (a or b);
    layer0_outputs(4029) <= not (a or b);
    layer0_outputs(4030) <= a or b;
    layer0_outputs(4031) <= not a or b;
    layer0_outputs(4032) <= a xor b;
    layer0_outputs(4033) <= not a;
    layer0_outputs(4034) <= b;
    layer0_outputs(4035) <= a or b;
    layer0_outputs(4036) <= not a or b;
    layer0_outputs(4037) <= not (a or b);
    layer0_outputs(4038) <= not (a and b);
    layer0_outputs(4039) <= b and not a;
    layer0_outputs(4040) <= '1';
    layer0_outputs(4041) <= not a;
    layer0_outputs(4042) <= not b;
    layer0_outputs(4043) <= not (a or b);
    layer0_outputs(4044) <= not a;
    layer0_outputs(4045) <= a xor b;
    layer0_outputs(4046) <= a and b;
    layer0_outputs(4047) <= not b or a;
    layer0_outputs(4048) <= a;
    layer0_outputs(4049) <= not a;
    layer0_outputs(4050) <= not a;
    layer0_outputs(4051) <= '0';
    layer0_outputs(4052) <= not (a or b);
    layer0_outputs(4053) <= a;
    layer0_outputs(4054) <= b and not a;
    layer0_outputs(4055) <= not a or b;
    layer0_outputs(4056) <= '1';
    layer0_outputs(4057) <= '0';
    layer0_outputs(4058) <= not a;
    layer0_outputs(4059) <= not b or a;
    layer0_outputs(4060) <= not (a and b);
    layer0_outputs(4061) <= not b or a;
    layer0_outputs(4062) <= a;
    layer0_outputs(4063) <= '1';
    layer0_outputs(4064) <= not a;
    layer0_outputs(4065) <= a or b;
    layer0_outputs(4066) <= not (a and b);
    layer0_outputs(4067) <= a or b;
    layer0_outputs(4068) <= '0';
    layer0_outputs(4069) <= a;
    layer0_outputs(4070) <= not b or a;
    layer0_outputs(4071) <= a;
    layer0_outputs(4072) <= '1';
    layer0_outputs(4073) <= a and b;
    layer0_outputs(4074) <= a and b;
    layer0_outputs(4075) <= '1';
    layer0_outputs(4076) <= not (a or b);
    layer0_outputs(4077) <= a and not b;
    layer0_outputs(4078) <= not (a and b);
    layer0_outputs(4079) <= not a or b;
    layer0_outputs(4080) <= b;
    layer0_outputs(4081) <= a;
    layer0_outputs(4082) <= not (a xor b);
    layer0_outputs(4083) <= not (a xor b);
    layer0_outputs(4084) <= a;
    layer0_outputs(4085) <= a and not b;
    layer0_outputs(4086) <= not a;
    layer0_outputs(4087) <= a;
    layer0_outputs(4088) <= not b;
    layer0_outputs(4089) <= a and not b;
    layer0_outputs(4090) <= a;
    layer0_outputs(4091) <= b and not a;
    layer0_outputs(4092) <= not b;
    layer0_outputs(4093) <= not a;
    layer0_outputs(4094) <= a;
    layer0_outputs(4095) <= not b or a;
    layer0_outputs(4096) <= a and not b;
    layer0_outputs(4097) <= a or b;
    layer0_outputs(4098) <= a xor b;
    layer0_outputs(4099) <= not a;
    layer0_outputs(4100) <= not b or a;
    layer0_outputs(4101) <= '1';
    layer0_outputs(4102) <= '0';
    layer0_outputs(4103) <= '0';
    layer0_outputs(4104) <= '1';
    layer0_outputs(4105) <= '1';
    layer0_outputs(4106) <= not (a and b);
    layer0_outputs(4107) <= a and b;
    layer0_outputs(4108) <= not (a xor b);
    layer0_outputs(4109) <= not (a or b);
    layer0_outputs(4110) <= '1';
    layer0_outputs(4111) <= '0';
    layer0_outputs(4112) <= b;
    layer0_outputs(4113) <= a or b;
    layer0_outputs(4114) <= not b;
    layer0_outputs(4115) <= a and b;
    layer0_outputs(4116) <= a;
    layer0_outputs(4117) <= not b or a;
    layer0_outputs(4118) <= not (a and b);
    layer0_outputs(4119) <= a;
    layer0_outputs(4120) <= not a;
    layer0_outputs(4121) <= a or b;
    layer0_outputs(4122) <= a or b;
    layer0_outputs(4123) <= not (a or b);
    layer0_outputs(4124) <= not a or b;
    layer0_outputs(4125) <= not b or a;
    layer0_outputs(4126) <= not (a xor b);
    layer0_outputs(4127) <= b and not a;
    layer0_outputs(4128) <= not a;
    layer0_outputs(4129) <= not a;
    layer0_outputs(4130) <= '1';
    layer0_outputs(4131) <= a or b;
    layer0_outputs(4132) <= '1';
    layer0_outputs(4133) <= a and b;
    layer0_outputs(4134) <= a;
    layer0_outputs(4135) <= a;
    layer0_outputs(4136) <= a;
    layer0_outputs(4137) <= not a;
    layer0_outputs(4138) <= a xor b;
    layer0_outputs(4139) <= not a;
    layer0_outputs(4140) <= not a or b;
    layer0_outputs(4141) <= a and not b;
    layer0_outputs(4142) <= a;
    layer0_outputs(4143) <= '1';
    layer0_outputs(4144) <= a and not b;
    layer0_outputs(4145) <= not a or b;
    layer0_outputs(4146) <= b;
    layer0_outputs(4147) <= b;
    layer0_outputs(4148) <= not (a and b);
    layer0_outputs(4149) <= not (a or b);
    layer0_outputs(4150) <= b and not a;
    layer0_outputs(4151) <= not a;
    layer0_outputs(4152) <= not b;
    layer0_outputs(4153) <= not (a xor b);
    layer0_outputs(4154) <= a and b;
    layer0_outputs(4155) <= not (a xor b);
    layer0_outputs(4156) <= a xor b;
    layer0_outputs(4157) <= not a or b;
    layer0_outputs(4158) <= not b;
    layer0_outputs(4159) <= not (a or b);
    layer0_outputs(4160) <= not a or b;
    layer0_outputs(4161) <= b and not a;
    layer0_outputs(4162) <= '1';
    layer0_outputs(4163) <= not a;
    layer0_outputs(4164) <= a;
    layer0_outputs(4165) <= not (a and b);
    layer0_outputs(4166) <= not b;
    layer0_outputs(4167) <= not b or a;
    layer0_outputs(4168) <= a and not b;
    layer0_outputs(4169) <= b and not a;
    layer0_outputs(4170) <= '1';
    layer0_outputs(4171) <= '1';
    layer0_outputs(4172) <= not (a xor b);
    layer0_outputs(4173) <= '1';
    layer0_outputs(4174) <= b;
    layer0_outputs(4175) <= b;
    layer0_outputs(4176) <= not a;
    layer0_outputs(4177) <= '1';
    layer0_outputs(4178) <= a;
    layer0_outputs(4179) <= not (a or b);
    layer0_outputs(4180) <= a or b;
    layer0_outputs(4181) <= a and not b;
    layer0_outputs(4182) <= a or b;
    layer0_outputs(4183) <= not b or a;
    layer0_outputs(4184) <= not (a and b);
    layer0_outputs(4185) <= b;
    layer0_outputs(4186) <= b;
    layer0_outputs(4187) <= not (a and b);
    layer0_outputs(4188) <= not (a or b);
    layer0_outputs(4189) <= b and not a;
    layer0_outputs(4190) <= '1';
    layer0_outputs(4191) <= b;
    layer0_outputs(4192) <= not b or a;
    layer0_outputs(4193) <= b;
    layer0_outputs(4194) <= a;
    layer0_outputs(4195) <= not a;
    layer0_outputs(4196) <= not a;
    layer0_outputs(4197) <= a or b;
    layer0_outputs(4198) <= b and not a;
    layer0_outputs(4199) <= not (a and b);
    layer0_outputs(4200) <= a;
    layer0_outputs(4201) <= b and not a;
    layer0_outputs(4202) <= b and not a;
    layer0_outputs(4203) <= a;
    layer0_outputs(4204) <= not (a xor b);
    layer0_outputs(4205) <= not a;
    layer0_outputs(4206) <= '1';
    layer0_outputs(4207) <= b and not a;
    layer0_outputs(4208) <= b and not a;
    layer0_outputs(4209) <= '1';
    layer0_outputs(4210) <= not a or b;
    layer0_outputs(4211) <= b and not a;
    layer0_outputs(4212) <= b;
    layer0_outputs(4213) <= '0';
    layer0_outputs(4214) <= a xor b;
    layer0_outputs(4215) <= not a;
    layer0_outputs(4216) <= a;
    layer0_outputs(4217) <= not b or a;
    layer0_outputs(4218) <= a;
    layer0_outputs(4219) <= a;
    layer0_outputs(4220) <= not a or b;
    layer0_outputs(4221) <= a xor b;
    layer0_outputs(4222) <= b;
    layer0_outputs(4223) <= not b or a;
    layer0_outputs(4224) <= a;
    layer0_outputs(4225) <= not (a or b);
    layer0_outputs(4226) <= b;
    layer0_outputs(4227) <= not a;
    layer0_outputs(4228) <= not a or b;
    layer0_outputs(4229) <= '0';
    layer0_outputs(4230) <= '0';
    layer0_outputs(4231) <= b;
    layer0_outputs(4232) <= a;
    layer0_outputs(4233) <= b;
    layer0_outputs(4234) <= not b or a;
    layer0_outputs(4235) <= not a;
    layer0_outputs(4236) <= not a or b;
    layer0_outputs(4237) <= b;
    layer0_outputs(4238) <= a;
    layer0_outputs(4239) <= a and not b;
    layer0_outputs(4240) <= not (a or b);
    layer0_outputs(4241) <= b;
    layer0_outputs(4242) <= not (a or b);
    layer0_outputs(4243) <= a and not b;
    layer0_outputs(4244) <= not b or a;
    layer0_outputs(4245) <= b and not a;
    layer0_outputs(4246) <= a xor b;
    layer0_outputs(4247) <= not a or b;
    layer0_outputs(4248) <= not a;
    layer0_outputs(4249) <= a;
    layer0_outputs(4250) <= not a or b;
    layer0_outputs(4251) <= not (a and b);
    layer0_outputs(4252) <= b;
    layer0_outputs(4253) <= not b;
    layer0_outputs(4254) <= b and not a;
    layer0_outputs(4255) <= a and b;
    layer0_outputs(4256) <= not a or b;
    layer0_outputs(4257) <= not (a or b);
    layer0_outputs(4258) <= a and not b;
    layer0_outputs(4259) <= not (a or b);
    layer0_outputs(4260) <= not a;
    layer0_outputs(4261) <= not (a or b);
    layer0_outputs(4262) <= a and not b;
    layer0_outputs(4263) <= not (a or b);
    layer0_outputs(4264) <= b and not a;
    layer0_outputs(4265) <= not a or b;
    layer0_outputs(4266) <= b;
    layer0_outputs(4267) <= '1';
    layer0_outputs(4268) <= not b or a;
    layer0_outputs(4269) <= a;
    layer0_outputs(4270) <= b and not a;
    layer0_outputs(4271) <= not b or a;
    layer0_outputs(4272) <= b;
    layer0_outputs(4273) <= a;
    layer0_outputs(4274) <= not (a or b);
    layer0_outputs(4275) <= '1';
    layer0_outputs(4276) <= '1';
    layer0_outputs(4277) <= b and not a;
    layer0_outputs(4278) <= a and not b;
    layer0_outputs(4279) <= a and b;
    layer0_outputs(4280) <= a and b;
    layer0_outputs(4281) <= not a or b;
    layer0_outputs(4282) <= a;
    layer0_outputs(4283) <= not (a and b);
    layer0_outputs(4284) <= a and b;
    layer0_outputs(4285) <= a or b;
    layer0_outputs(4286) <= b;
    layer0_outputs(4287) <= '0';
    layer0_outputs(4288) <= b and not a;
    layer0_outputs(4289) <= a xor b;
    layer0_outputs(4290) <= a xor b;
    layer0_outputs(4291) <= b;
    layer0_outputs(4292) <= a xor b;
    layer0_outputs(4293) <= '1';
    layer0_outputs(4294) <= not (a or b);
    layer0_outputs(4295) <= not b or a;
    layer0_outputs(4296) <= not a or b;
    layer0_outputs(4297) <= '1';
    layer0_outputs(4298) <= a and not b;
    layer0_outputs(4299) <= b;
    layer0_outputs(4300) <= not (a xor b);
    layer0_outputs(4301) <= a or b;
    layer0_outputs(4302) <= not (a and b);
    layer0_outputs(4303) <= not (a or b);
    layer0_outputs(4304) <= a and not b;
    layer0_outputs(4305) <= a;
    layer0_outputs(4306) <= a or b;
    layer0_outputs(4307) <= not (a xor b);
    layer0_outputs(4308) <= not (a xor b);
    layer0_outputs(4309) <= not (a or b);
    layer0_outputs(4310) <= b and not a;
    layer0_outputs(4311) <= a xor b;
    layer0_outputs(4312) <= a xor b;
    layer0_outputs(4313) <= not (a or b);
    layer0_outputs(4314) <= not a or b;
    layer0_outputs(4315) <= a and not b;
    layer0_outputs(4316) <= not b;
    layer0_outputs(4317) <= a;
    layer0_outputs(4318) <= a;
    layer0_outputs(4319) <= a or b;
    layer0_outputs(4320) <= '1';
    layer0_outputs(4321) <= not a;
    layer0_outputs(4322) <= not (a and b);
    layer0_outputs(4323) <= not a;
    layer0_outputs(4324) <= not (a xor b);
    layer0_outputs(4325) <= a or b;
    layer0_outputs(4326) <= b;
    layer0_outputs(4327) <= not b or a;
    layer0_outputs(4328) <= b;
    layer0_outputs(4329) <= not b;
    layer0_outputs(4330) <= b and not a;
    layer0_outputs(4331) <= not a or b;
    layer0_outputs(4332) <= not a or b;
    layer0_outputs(4333) <= a and not b;
    layer0_outputs(4334) <= a or b;
    layer0_outputs(4335) <= b and not a;
    layer0_outputs(4336) <= not b;
    layer0_outputs(4337) <= '0';
    layer0_outputs(4338) <= not b or a;
    layer0_outputs(4339) <= not (a or b);
    layer0_outputs(4340) <= a xor b;
    layer0_outputs(4341) <= '0';
    layer0_outputs(4342) <= not (a or b);
    layer0_outputs(4343) <= not a or b;
    layer0_outputs(4344) <= '0';
    layer0_outputs(4345) <= a and b;
    layer0_outputs(4346) <= b and not a;
    layer0_outputs(4347) <= a or b;
    layer0_outputs(4348) <= '1';
    layer0_outputs(4349) <= '0';
    layer0_outputs(4350) <= '1';
    layer0_outputs(4351) <= not (a or b);
    layer0_outputs(4352) <= a or b;
    layer0_outputs(4353) <= a;
    layer0_outputs(4354) <= not (a or b);
    layer0_outputs(4355) <= not a;
    layer0_outputs(4356) <= a or b;
    layer0_outputs(4357) <= not (a and b);
    layer0_outputs(4358) <= b;
    layer0_outputs(4359) <= '0';
    layer0_outputs(4360) <= '1';
    layer0_outputs(4361) <= '0';
    layer0_outputs(4362) <= '0';
    layer0_outputs(4363) <= not (a xor b);
    layer0_outputs(4364) <= not (a or b);
    layer0_outputs(4365) <= a or b;
    layer0_outputs(4366) <= '1';
    layer0_outputs(4367) <= a;
    layer0_outputs(4368) <= not (a or b);
    layer0_outputs(4369) <= not (a and b);
    layer0_outputs(4370) <= a and b;
    layer0_outputs(4371) <= '1';
    layer0_outputs(4372) <= b and not a;
    layer0_outputs(4373) <= '0';
    layer0_outputs(4374) <= b;
    layer0_outputs(4375) <= not b;
    layer0_outputs(4376) <= not a or b;
    layer0_outputs(4377) <= not a or b;
    layer0_outputs(4378) <= '0';
    layer0_outputs(4379) <= not (a or b);
    layer0_outputs(4380) <= not (a xor b);
    layer0_outputs(4381) <= not (a xor b);
    layer0_outputs(4382) <= a;
    layer0_outputs(4383) <= not (a xor b);
    layer0_outputs(4384) <= '0';
    layer0_outputs(4385) <= not a or b;
    layer0_outputs(4386) <= not (a and b);
    layer0_outputs(4387) <= not (a xor b);
    layer0_outputs(4388) <= a and not b;
    layer0_outputs(4389) <= a or b;
    layer0_outputs(4390) <= '0';
    layer0_outputs(4391) <= b;
    layer0_outputs(4392) <= a and b;
    layer0_outputs(4393) <= b;
    layer0_outputs(4394) <= not (a or b);
    layer0_outputs(4395) <= '0';
    layer0_outputs(4396) <= not a;
    layer0_outputs(4397) <= a;
    layer0_outputs(4398) <= a xor b;
    layer0_outputs(4399) <= a;
    layer0_outputs(4400) <= not b or a;
    layer0_outputs(4401) <= not a or b;
    layer0_outputs(4402) <= '0';
    layer0_outputs(4403) <= not (a xor b);
    layer0_outputs(4404) <= not a;
    layer0_outputs(4405) <= '1';
    layer0_outputs(4406) <= a and not b;
    layer0_outputs(4407) <= not (a or b);
    layer0_outputs(4408) <= b;
    layer0_outputs(4409) <= not (a and b);
    layer0_outputs(4410) <= '0';
    layer0_outputs(4411) <= a;
    layer0_outputs(4412) <= b;
    layer0_outputs(4413) <= '1';
    layer0_outputs(4414) <= a;
    layer0_outputs(4415) <= '0';
    layer0_outputs(4416) <= b and not a;
    layer0_outputs(4417) <= not a;
    layer0_outputs(4418) <= b and not a;
    layer0_outputs(4419) <= '0';
    layer0_outputs(4420) <= not b or a;
    layer0_outputs(4421) <= a and not b;
    layer0_outputs(4422) <= a and b;
    layer0_outputs(4423) <= not (a and b);
    layer0_outputs(4424) <= a and b;
    layer0_outputs(4425) <= not (a xor b);
    layer0_outputs(4426) <= a xor b;
    layer0_outputs(4427) <= b;
    layer0_outputs(4428) <= not b;
    layer0_outputs(4429) <= b and not a;
    layer0_outputs(4430) <= '1';
    layer0_outputs(4431) <= a and not b;
    layer0_outputs(4432) <= not a;
    layer0_outputs(4433) <= b;
    layer0_outputs(4434) <= b;
    layer0_outputs(4435) <= a;
    layer0_outputs(4436) <= a and b;
    layer0_outputs(4437) <= not b or a;
    layer0_outputs(4438) <= not b or a;
    layer0_outputs(4439) <= not a;
    layer0_outputs(4440) <= a xor b;
    layer0_outputs(4441) <= not a;
    layer0_outputs(4442) <= not a or b;
    layer0_outputs(4443) <= not (a or b);
    layer0_outputs(4444) <= not (a or b);
    layer0_outputs(4445) <= b and not a;
    layer0_outputs(4446) <= not b;
    layer0_outputs(4447) <= not (a or b);
    layer0_outputs(4448) <= not (a and b);
    layer0_outputs(4449) <= '0';
    layer0_outputs(4450) <= a and not b;
    layer0_outputs(4451) <= a and b;
    layer0_outputs(4452) <= not b or a;
    layer0_outputs(4453) <= not (a and b);
    layer0_outputs(4454) <= a and b;
    layer0_outputs(4455) <= a xor b;
    layer0_outputs(4456) <= b and not a;
    layer0_outputs(4457) <= b;
    layer0_outputs(4458) <= '0';
    layer0_outputs(4459) <= not b or a;
    layer0_outputs(4460) <= '0';
    layer0_outputs(4461) <= not a or b;
    layer0_outputs(4462) <= a and b;
    layer0_outputs(4463) <= not b;
    layer0_outputs(4464) <= '0';
    layer0_outputs(4465) <= b;
    layer0_outputs(4466) <= not a or b;
    layer0_outputs(4467) <= a and not b;
    layer0_outputs(4468) <= a and not b;
    layer0_outputs(4469) <= not a;
    layer0_outputs(4470) <= not (a xor b);
    layer0_outputs(4471) <= a and not b;
    layer0_outputs(4472) <= not b;
    layer0_outputs(4473) <= '0';
    layer0_outputs(4474) <= a;
    layer0_outputs(4475) <= '0';
    layer0_outputs(4476) <= not a;
    layer0_outputs(4477) <= not b or a;
    layer0_outputs(4478) <= b and not a;
    layer0_outputs(4479) <= a and b;
    layer0_outputs(4480) <= not (a or b);
    layer0_outputs(4481) <= '1';
    layer0_outputs(4482) <= not a;
    layer0_outputs(4483) <= not a or b;
    layer0_outputs(4484) <= not b;
    layer0_outputs(4485) <= a;
    layer0_outputs(4486) <= a;
    layer0_outputs(4487) <= '1';
    layer0_outputs(4488) <= not (a xor b);
    layer0_outputs(4489) <= a and not b;
    layer0_outputs(4490) <= '1';
    layer0_outputs(4491) <= a or b;
    layer0_outputs(4492) <= a xor b;
    layer0_outputs(4493) <= a or b;
    layer0_outputs(4494) <= b;
    layer0_outputs(4495) <= not (a and b);
    layer0_outputs(4496) <= not a;
    layer0_outputs(4497) <= a xor b;
    layer0_outputs(4498) <= b;
    layer0_outputs(4499) <= not a or b;
    layer0_outputs(4500) <= not a;
    layer0_outputs(4501) <= not a or b;
    layer0_outputs(4502) <= not b;
    layer0_outputs(4503) <= '0';
    layer0_outputs(4504) <= not a or b;
    layer0_outputs(4505) <= '0';
    layer0_outputs(4506) <= not a;
    layer0_outputs(4507) <= a or b;
    layer0_outputs(4508) <= not (a and b);
    layer0_outputs(4509) <= not b or a;
    layer0_outputs(4510) <= '1';
    layer0_outputs(4511) <= '1';
    layer0_outputs(4512) <= not a or b;
    layer0_outputs(4513) <= not (a and b);
    layer0_outputs(4514) <= '0';
    layer0_outputs(4515) <= '0';
    layer0_outputs(4516) <= not (a and b);
    layer0_outputs(4517) <= not a;
    layer0_outputs(4518) <= b;
    layer0_outputs(4519) <= not (a and b);
    layer0_outputs(4520) <= a;
    layer0_outputs(4521) <= not b;
    layer0_outputs(4522) <= not (a or b);
    layer0_outputs(4523) <= '0';
    layer0_outputs(4524) <= a xor b;
    layer0_outputs(4525) <= a or b;
    layer0_outputs(4526) <= '1';
    layer0_outputs(4527) <= not (a xor b);
    layer0_outputs(4528) <= not b;
    layer0_outputs(4529) <= a or b;
    layer0_outputs(4530) <= not b;
    layer0_outputs(4531) <= a or b;
    layer0_outputs(4532) <= not (a xor b);
    layer0_outputs(4533) <= not (a and b);
    layer0_outputs(4534) <= not (a or b);
    layer0_outputs(4535) <= not a;
    layer0_outputs(4536) <= a or b;
    layer0_outputs(4537) <= not a or b;
    layer0_outputs(4538) <= not b or a;
    layer0_outputs(4539) <= b;
    layer0_outputs(4540) <= '0';
    layer0_outputs(4541) <= a and b;
    layer0_outputs(4542) <= a and not b;
    layer0_outputs(4543) <= b and not a;
    layer0_outputs(4544) <= a and b;
    layer0_outputs(4545) <= not (a xor b);
    layer0_outputs(4546) <= a and b;
    layer0_outputs(4547) <= '0';
    layer0_outputs(4548) <= a or b;
    layer0_outputs(4549) <= '0';
    layer0_outputs(4550) <= not b or a;
    layer0_outputs(4551) <= b;
    layer0_outputs(4552) <= not a;
    layer0_outputs(4553) <= not (a xor b);
    layer0_outputs(4554) <= '0';
    layer0_outputs(4555) <= a;
    layer0_outputs(4556) <= not a;
    layer0_outputs(4557) <= a and not b;
    layer0_outputs(4558) <= b and not a;
    layer0_outputs(4559) <= not (a or b);
    layer0_outputs(4560) <= not a or b;
    layer0_outputs(4561) <= b;
    layer0_outputs(4562) <= not b;
    layer0_outputs(4563) <= not b or a;
    layer0_outputs(4564) <= not a;
    layer0_outputs(4565) <= a or b;
    layer0_outputs(4566) <= b and not a;
    layer0_outputs(4567) <= '0';
    layer0_outputs(4568) <= a and b;
    layer0_outputs(4569) <= a and not b;
    layer0_outputs(4570) <= a;
    layer0_outputs(4571) <= not a or b;
    layer0_outputs(4572) <= not (a or b);
    layer0_outputs(4573) <= not a or b;
    layer0_outputs(4574) <= not b or a;
    layer0_outputs(4575) <= not b or a;
    layer0_outputs(4576) <= a and b;
    layer0_outputs(4577) <= not (a and b);
    layer0_outputs(4578) <= a or b;
    layer0_outputs(4579) <= not b;
    layer0_outputs(4580) <= a and b;
    layer0_outputs(4581) <= '1';
    layer0_outputs(4582) <= not a or b;
    layer0_outputs(4583) <= a and not b;
    layer0_outputs(4584) <= not a;
    layer0_outputs(4585) <= a;
    layer0_outputs(4586) <= '0';
    layer0_outputs(4587) <= '1';
    layer0_outputs(4588) <= a and not b;
    layer0_outputs(4589) <= b;
    layer0_outputs(4590) <= a and b;
    layer0_outputs(4591) <= '1';
    layer0_outputs(4592) <= '1';
    layer0_outputs(4593) <= not a;
    layer0_outputs(4594) <= not (a xor b);
    layer0_outputs(4595) <= not (a or b);
    layer0_outputs(4596) <= '0';
    layer0_outputs(4597) <= not (a and b);
    layer0_outputs(4598) <= not (a or b);
    layer0_outputs(4599) <= not a or b;
    layer0_outputs(4600) <= '1';
    layer0_outputs(4601) <= a and not b;
    layer0_outputs(4602) <= '1';
    layer0_outputs(4603) <= a and not b;
    layer0_outputs(4604) <= not b or a;
    layer0_outputs(4605) <= a and b;
    layer0_outputs(4606) <= b and not a;
    layer0_outputs(4607) <= '1';
    layer0_outputs(4608) <= not a;
    layer0_outputs(4609) <= a;
    layer0_outputs(4610) <= '0';
    layer0_outputs(4611) <= b and not a;
    layer0_outputs(4612) <= a and not b;
    layer0_outputs(4613) <= '1';
    layer0_outputs(4614) <= not b;
    layer0_outputs(4615) <= not (a or b);
    layer0_outputs(4616) <= not (a or b);
    layer0_outputs(4617) <= not (a or b);
    layer0_outputs(4618) <= not a;
    layer0_outputs(4619) <= b and not a;
    layer0_outputs(4620) <= not b or a;
    layer0_outputs(4621) <= not a or b;
    layer0_outputs(4622) <= b and not a;
    layer0_outputs(4623) <= b;
    layer0_outputs(4624) <= not b or a;
    layer0_outputs(4625) <= a xor b;
    layer0_outputs(4626) <= not (a and b);
    layer0_outputs(4627) <= not b;
    layer0_outputs(4628) <= not a or b;
    layer0_outputs(4629) <= b;
    layer0_outputs(4630) <= a xor b;
    layer0_outputs(4631) <= '1';
    layer0_outputs(4632) <= a and not b;
    layer0_outputs(4633) <= '1';
    layer0_outputs(4634) <= b;
    layer0_outputs(4635) <= not b or a;
    layer0_outputs(4636) <= not (a and b);
    layer0_outputs(4637) <= not a;
    layer0_outputs(4638) <= not b;
    layer0_outputs(4639) <= '0';
    layer0_outputs(4640) <= not (a or b);
    layer0_outputs(4641) <= not b or a;
    layer0_outputs(4642) <= '0';
    layer0_outputs(4643) <= not (a and b);
    layer0_outputs(4644) <= a;
    layer0_outputs(4645) <= b and not a;
    layer0_outputs(4646) <= '1';
    layer0_outputs(4647) <= b and not a;
    layer0_outputs(4648) <= '1';
    layer0_outputs(4649) <= '0';
    layer0_outputs(4650) <= not (a or b);
    layer0_outputs(4651) <= '0';
    layer0_outputs(4652) <= not a;
    layer0_outputs(4653) <= a and not b;
    layer0_outputs(4654) <= not b or a;
    layer0_outputs(4655) <= '1';
    layer0_outputs(4656) <= not (a and b);
    layer0_outputs(4657) <= '1';
    layer0_outputs(4658) <= a;
    layer0_outputs(4659) <= not a;
    layer0_outputs(4660) <= a and not b;
    layer0_outputs(4661) <= not a;
    layer0_outputs(4662) <= not b;
    layer0_outputs(4663) <= '1';
    layer0_outputs(4664) <= a xor b;
    layer0_outputs(4665) <= not a;
    layer0_outputs(4666) <= a and not b;
    layer0_outputs(4667) <= a;
    layer0_outputs(4668) <= a xor b;
    layer0_outputs(4669) <= a and not b;
    layer0_outputs(4670) <= a and b;
    layer0_outputs(4671) <= not (a xor b);
    layer0_outputs(4672) <= not b or a;
    layer0_outputs(4673) <= b;
    layer0_outputs(4674) <= a;
    layer0_outputs(4675) <= not (a xor b);
    layer0_outputs(4676) <= '0';
    layer0_outputs(4677) <= not (a and b);
    layer0_outputs(4678) <= a or b;
    layer0_outputs(4679) <= not a;
    layer0_outputs(4680) <= '0';
    layer0_outputs(4681) <= a and b;
    layer0_outputs(4682) <= not b or a;
    layer0_outputs(4683) <= not a or b;
    layer0_outputs(4684) <= not a;
    layer0_outputs(4685) <= a and b;
    layer0_outputs(4686) <= not (a and b);
    layer0_outputs(4687) <= not b or a;
    layer0_outputs(4688) <= a;
    layer0_outputs(4689) <= a and not b;
    layer0_outputs(4690) <= b;
    layer0_outputs(4691) <= not b or a;
    layer0_outputs(4692) <= '1';
    layer0_outputs(4693) <= b;
    layer0_outputs(4694) <= not b or a;
    layer0_outputs(4695) <= '0';
    layer0_outputs(4696) <= b;
    layer0_outputs(4697) <= '1';
    layer0_outputs(4698) <= not (a or b);
    layer0_outputs(4699) <= not (a or b);
    layer0_outputs(4700) <= not a;
    layer0_outputs(4701) <= '1';
    layer0_outputs(4702) <= not a or b;
    layer0_outputs(4703) <= not a;
    layer0_outputs(4704) <= '1';
    layer0_outputs(4705) <= not b or a;
    layer0_outputs(4706) <= not b;
    layer0_outputs(4707) <= b and not a;
    layer0_outputs(4708) <= not b or a;
    layer0_outputs(4709) <= not (a or b);
    layer0_outputs(4710) <= not (a and b);
    layer0_outputs(4711) <= '1';
    layer0_outputs(4712) <= a or b;
    layer0_outputs(4713) <= a xor b;
    layer0_outputs(4714) <= a;
    layer0_outputs(4715) <= not b;
    layer0_outputs(4716) <= '1';
    layer0_outputs(4717) <= not a or b;
    layer0_outputs(4718) <= a and not b;
    layer0_outputs(4719) <= not (a and b);
    layer0_outputs(4720) <= not (a and b);
    layer0_outputs(4721) <= '0';
    layer0_outputs(4722) <= a;
    layer0_outputs(4723) <= '1';
    layer0_outputs(4724) <= '1';
    layer0_outputs(4725) <= not b;
    layer0_outputs(4726) <= '0';
    layer0_outputs(4727) <= a;
    layer0_outputs(4728) <= not a or b;
    layer0_outputs(4729) <= not (a xor b);
    layer0_outputs(4730) <= '0';
    layer0_outputs(4731) <= a or b;
    layer0_outputs(4732) <= a or b;
    layer0_outputs(4733) <= a xor b;
    layer0_outputs(4734) <= '0';
    layer0_outputs(4735) <= a or b;
    layer0_outputs(4736) <= a and not b;
    layer0_outputs(4737) <= not a;
    layer0_outputs(4738) <= not (a xor b);
    layer0_outputs(4739) <= a;
    layer0_outputs(4740) <= a and not b;
    layer0_outputs(4741) <= not (a or b);
    layer0_outputs(4742) <= not (a or b);
    layer0_outputs(4743) <= '0';
    layer0_outputs(4744) <= '1';
    layer0_outputs(4745) <= b and not a;
    layer0_outputs(4746) <= a;
    layer0_outputs(4747) <= '1';
    layer0_outputs(4748) <= '1';
    layer0_outputs(4749) <= a or b;
    layer0_outputs(4750) <= a;
    layer0_outputs(4751) <= not (a or b);
    layer0_outputs(4752) <= a;
    layer0_outputs(4753) <= b;
    layer0_outputs(4754) <= '0';
    layer0_outputs(4755) <= a and not b;
    layer0_outputs(4756) <= not b or a;
    layer0_outputs(4757) <= not (a xor b);
    layer0_outputs(4758) <= a or b;
    layer0_outputs(4759) <= not b;
    layer0_outputs(4760) <= b;
    layer0_outputs(4761) <= not (a and b);
    layer0_outputs(4762) <= not a;
    layer0_outputs(4763) <= not a;
    layer0_outputs(4764) <= not a;
    layer0_outputs(4765) <= not (a xor b);
    layer0_outputs(4766) <= a and b;
    layer0_outputs(4767) <= b;
    layer0_outputs(4768) <= not (a or b);
    layer0_outputs(4769) <= a or b;
    layer0_outputs(4770) <= not (a and b);
    layer0_outputs(4771) <= '1';
    layer0_outputs(4772) <= not (a xor b);
    layer0_outputs(4773) <= not (a xor b);
    layer0_outputs(4774) <= a and b;
    layer0_outputs(4775) <= not (a and b);
    layer0_outputs(4776) <= not a;
    layer0_outputs(4777) <= b and not a;
    layer0_outputs(4778) <= b;
    layer0_outputs(4779) <= b and not a;
    layer0_outputs(4780) <= b;
    layer0_outputs(4781) <= a;
    layer0_outputs(4782) <= a;
    layer0_outputs(4783) <= a and b;
    layer0_outputs(4784) <= not (a or b);
    layer0_outputs(4785) <= not a or b;
    layer0_outputs(4786) <= b;
    layer0_outputs(4787) <= '0';
    layer0_outputs(4788) <= '1';
    layer0_outputs(4789) <= not b;
    layer0_outputs(4790) <= a and not b;
    layer0_outputs(4791) <= b and not a;
    layer0_outputs(4792) <= not (a or b);
    layer0_outputs(4793) <= not b or a;
    layer0_outputs(4794) <= not (a xor b);
    layer0_outputs(4795) <= not (a and b);
    layer0_outputs(4796) <= not b;
    layer0_outputs(4797) <= not b;
    layer0_outputs(4798) <= '1';
    layer0_outputs(4799) <= not (a xor b);
    layer0_outputs(4800) <= a;
    layer0_outputs(4801) <= a;
    layer0_outputs(4802) <= b;
    layer0_outputs(4803) <= not (a xor b);
    layer0_outputs(4804) <= a;
    layer0_outputs(4805) <= '1';
    layer0_outputs(4806) <= not b or a;
    layer0_outputs(4807) <= a;
    layer0_outputs(4808) <= a and b;
    layer0_outputs(4809) <= a xor b;
    layer0_outputs(4810) <= not a;
    layer0_outputs(4811) <= not a;
    layer0_outputs(4812) <= '0';
    layer0_outputs(4813) <= not (a or b);
    layer0_outputs(4814) <= not (a or b);
    layer0_outputs(4815) <= a and not b;
    layer0_outputs(4816) <= not (a xor b);
    layer0_outputs(4817) <= not a;
    layer0_outputs(4818) <= b and not a;
    layer0_outputs(4819) <= b;
    layer0_outputs(4820) <= a or b;
    layer0_outputs(4821) <= not a or b;
    layer0_outputs(4822) <= not (a xor b);
    layer0_outputs(4823) <= '0';
    layer0_outputs(4824) <= a;
    layer0_outputs(4825) <= b and not a;
    layer0_outputs(4826) <= not b or a;
    layer0_outputs(4827) <= not b;
    layer0_outputs(4828) <= b;
    layer0_outputs(4829) <= not (a or b);
    layer0_outputs(4830) <= '1';
    layer0_outputs(4831) <= not a or b;
    layer0_outputs(4832) <= a;
    layer0_outputs(4833) <= not (a and b);
    layer0_outputs(4834) <= a and not b;
    layer0_outputs(4835) <= a xor b;
    layer0_outputs(4836) <= '0';
    layer0_outputs(4837) <= '0';
    layer0_outputs(4838) <= b and not a;
    layer0_outputs(4839) <= a and not b;
    layer0_outputs(4840) <= not (a and b);
    layer0_outputs(4841) <= not (a or b);
    layer0_outputs(4842) <= b;
    layer0_outputs(4843) <= '0';
    layer0_outputs(4844) <= a xor b;
    layer0_outputs(4845) <= not (a or b);
    layer0_outputs(4846) <= not (a and b);
    layer0_outputs(4847) <= not (a xor b);
    layer0_outputs(4848) <= '0';
    layer0_outputs(4849) <= b;
    layer0_outputs(4850) <= '0';
    layer0_outputs(4851) <= not b;
    layer0_outputs(4852) <= not b or a;
    layer0_outputs(4853) <= not (a or b);
    layer0_outputs(4854) <= not (a and b);
    layer0_outputs(4855) <= not a;
    layer0_outputs(4856) <= a or b;
    layer0_outputs(4857) <= not a;
    layer0_outputs(4858) <= a and b;
    layer0_outputs(4859) <= not (a xor b);
    layer0_outputs(4860) <= b;
    layer0_outputs(4861) <= a xor b;
    layer0_outputs(4862) <= not a or b;
    layer0_outputs(4863) <= b and not a;
    layer0_outputs(4864) <= not b or a;
    layer0_outputs(4865) <= b and not a;
    layer0_outputs(4866) <= a and not b;
    layer0_outputs(4867) <= a;
    layer0_outputs(4868) <= '0';
    layer0_outputs(4869) <= a and b;
    layer0_outputs(4870) <= '0';
    layer0_outputs(4871) <= not (a xor b);
    layer0_outputs(4872) <= not a or b;
    layer0_outputs(4873) <= not b or a;
    layer0_outputs(4874) <= b and not a;
    layer0_outputs(4875) <= not a;
    layer0_outputs(4876) <= a or b;
    layer0_outputs(4877) <= not a;
    layer0_outputs(4878) <= a and not b;
    layer0_outputs(4879) <= a;
    layer0_outputs(4880) <= not (a or b);
    layer0_outputs(4881) <= a and not b;
    layer0_outputs(4882) <= b and not a;
    layer0_outputs(4883) <= b;
    layer0_outputs(4884) <= a or b;
    layer0_outputs(4885) <= not b;
    layer0_outputs(4886) <= '1';
    layer0_outputs(4887) <= not b or a;
    layer0_outputs(4888) <= a and b;
    layer0_outputs(4889) <= a or b;
    layer0_outputs(4890) <= a xor b;
    layer0_outputs(4891) <= b;
    layer0_outputs(4892) <= a xor b;
    layer0_outputs(4893) <= not a;
    layer0_outputs(4894) <= a or b;
    layer0_outputs(4895) <= not a or b;
    layer0_outputs(4896) <= a and not b;
    layer0_outputs(4897) <= '0';
    layer0_outputs(4898) <= '0';
    layer0_outputs(4899) <= not a or b;
    layer0_outputs(4900) <= a xor b;
    layer0_outputs(4901) <= not (a or b);
    layer0_outputs(4902) <= a;
    layer0_outputs(4903) <= not b or a;
    layer0_outputs(4904) <= b and not a;
    layer0_outputs(4905) <= a;
    layer0_outputs(4906) <= b and not a;
    layer0_outputs(4907) <= '1';
    layer0_outputs(4908) <= a xor b;
    layer0_outputs(4909) <= b and not a;
    layer0_outputs(4910) <= not (a and b);
    layer0_outputs(4911) <= a xor b;
    layer0_outputs(4912) <= a and b;
    layer0_outputs(4913) <= not b or a;
    layer0_outputs(4914) <= not (a or b);
    layer0_outputs(4915) <= not b or a;
    layer0_outputs(4916) <= not (a xor b);
    layer0_outputs(4917) <= not (a and b);
    layer0_outputs(4918) <= a;
    layer0_outputs(4919) <= a xor b;
    layer0_outputs(4920) <= a and b;
    layer0_outputs(4921) <= '1';
    layer0_outputs(4922) <= not a;
    layer0_outputs(4923) <= not (a or b);
    layer0_outputs(4924) <= not b or a;
    layer0_outputs(4925) <= a or b;
    layer0_outputs(4926) <= not b;
    layer0_outputs(4927) <= a;
    layer0_outputs(4928) <= not a or b;
    layer0_outputs(4929) <= a;
    layer0_outputs(4930) <= not (a or b);
    layer0_outputs(4931) <= not b or a;
    layer0_outputs(4932) <= not a;
    layer0_outputs(4933) <= not a or b;
    layer0_outputs(4934) <= a and b;
    layer0_outputs(4935) <= not (a xor b);
    layer0_outputs(4936) <= '0';
    layer0_outputs(4937) <= a;
    layer0_outputs(4938) <= '1';
    layer0_outputs(4939) <= not b or a;
    layer0_outputs(4940) <= not (a or b);
    layer0_outputs(4941) <= a and not b;
    layer0_outputs(4942) <= not a or b;
    layer0_outputs(4943) <= a and b;
    layer0_outputs(4944) <= not (a xor b);
    layer0_outputs(4945) <= a xor b;
    layer0_outputs(4946) <= a xor b;
    layer0_outputs(4947) <= not (a and b);
    layer0_outputs(4948) <= b and not a;
    layer0_outputs(4949) <= not b;
    layer0_outputs(4950) <= '0';
    layer0_outputs(4951) <= b;
    layer0_outputs(4952) <= a and not b;
    layer0_outputs(4953) <= b and not a;
    layer0_outputs(4954) <= b;
    layer0_outputs(4955) <= '1';
    layer0_outputs(4956) <= a or b;
    layer0_outputs(4957) <= a or b;
    layer0_outputs(4958) <= not b or a;
    layer0_outputs(4959) <= '1';
    layer0_outputs(4960) <= '1';
    layer0_outputs(4961) <= a xor b;
    layer0_outputs(4962) <= not b or a;
    layer0_outputs(4963) <= a or b;
    layer0_outputs(4964) <= a and not b;
    layer0_outputs(4965) <= b;
    layer0_outputs(4966) <= '1';
    layer0_outputs(4967) <= '0';
    layer0_outputs(4968) <= a and not b;
    layer0_outputs(4969) <= a and b;
    layer0_outputs(4970) <= a;
    layer0_outputs(4971) <= not (a xor b);
    layer0_outputs(4972) <= a xor b;
    layer0_outputs(4973) <= not a;
    layer0_outputs(4974) <= not (a and b);
    layer0_outputs(4975) <= not a or b;
    layer0_outputs(4976) <= not (a or b);
    layer0_outputs(4977) <= '1';
    layer0_outputs(4978) <= b and not a;
    layer0_outputs(4979) <= b and not a;
    layer0_outputs(4980) <= a;
    layer0_outputs(4981) <= not (a and b);
    layer0_outputs(4982) <= b and not a;
    layer0_outputs(4983) <= b;
    layer0_outputs(4984) <= '1';
    layer0_outputs(4985) <= not b or a;
    layer0_outputs(4986) <= not (a xor b);
    layer0_outputs(4987) <= not (a xor b);
    layer0_outputs(4988) <= not a or b;
    layer0_outputs(4989) <= a and b;
    layer0_outputs(4990) <= a and not b;
    layer0_outputs(4991) <= a or b;
    layer0_outputs(4992) <= a and b;
    layer0_outputs(4993) <= not b;
    layer0_outputs(4994) <= a and b;
    layer0_outputs(4995) <= not (a or b);
    layer0_outputs(4996) <= b;
    layer0_outputs(4997) <= b;
    layer0_outputs(4998) <= a;
    layer0_outputs(4999) <= '1';
    layer0_outputs(5000) <= not a;
    layer0_outputs(5001) <= not a;
    layer0_outputs(5002) <= '0';
    layer0_outputs(5003) <= a xor b;
    layer0_outputs(5004) <= a;
    layer0_outputs(5005) <= not b or a;
    layer0_outputs(5006) <= a and not b;
    layer0_outputs(5007) <= not b;
    layer0_outputs(5008) <= a;
    layer0_outputs(5009) <= not a or b;
    layer0_outputs(5010) <= b and not a;
    layer0_outputs(5011) <= '0';
    layer0_outputs(5012) <= not (a or b);
    layer0_outputs(5013) <= not b;
    layer0_outputs(5014) <= not a;
    layer0_outputs(5015) <= b and not a;
    layer0_outputs(5016) <= not (a and b);
    layer0_outputs(5017) <= '1';
    layer0_outputs(5018) <= a;
    layer0_outputs(5019) <= not b;
    layer0_outputs(5020) <= '1';
    layer0_outputs(5021) <= '1';
    layer0_outputs(5022) <= not a;
    layer0_outputs(5023) <= b;
    layer0_outputs(5024) <= not b;
    layer0_outputs(5025) <= not (a xor b);
    layer0_outputs(5026) <= a and not b;
    layer0_outputs(5027) <= not a or b;
    layer0_outputs(5028) <= not (a and b);
    layer0_outputs(5029) <= '0';
    layer0_outputs(5030) <= '1';
    layer0_outputs(5031) <= b;
    layer0_outputs(5032) <= a and not b;
    layer0_outputs(5033) <= not (a xor b);
    layer0_outputs(5034) <= '1';
    layer0_outputs(5035) <= a and not b;
    layer0_outputs(5036) <= a xor b;
    layer0_outputs(5037) <= not a or b;
    layer0_outputs(5038) <= a or b;
    layer0_outputs(5039) <= not b or a;
    layer0_outputs(5040) <= a;
    layer0_outputs(5041) <= '1';
    layer0_outputs(5042) <= not (a and b);
    layer0_outputs(5043) <= not a;
    layer0_outputs(5044) <= a;
    layer0_outputs(5045) <= a and b;
    layer0_outputs(5046) <= a or b;
    layer0_outputs(5047) <= not a or b;
    layer0_outputs(5048) <= not (a and b);
    layer0_outputs(5049) <= '1';
    layer0_outputs(5050) <= not (a or b);
    layer0_outputs(5051) <= not (a and b);
    layer0_outputs(5052) <= not a;
    layer0_outputs(5053) <= b;
    layer0_outputs(5054) <= not (a or b);
    layer0_outputs(5055) <= not (a or b);
    layer0_outputs(5056) <= '1';
    layer0_outputs(5057) <= '0';
    layer0_outputs(5058) <= not a or b;
    layer0_outputs(5059) <= '0';
    layer0_outputs(5060) <= b;
    layer0_outputs(5061) <= b and not a;
    layer0_outputs(5062) <= not b;
    layer0_outputs(5063) <= not b or a;
    layer0_outputs(5064) <= not a;
    layer0_outputs(5065) <= b;
    layer0_outputs(5066) <= b;
    layer0_outputs(5067) <= '0';
    layer0_outputs(5068) <= not a;
    layer0_outputs(5069) <= '0';
    layer0_outputs(5070) <= not (a xor b);
    layer0_outputs(5071) <= not a;
    layer0_outputs(5072) <= a and not b;
    layer0_outputs(5073) <= '0';
    layer0_outputs(5074) <= b;
    layer0_outputs(5075) <= a and b;
    layer0_outputs(5076) <= not (a or b);
    layer0_outputs(5077) <= b and not a;
    layer0_outputs(5078) <= not b or a;
    layer0_outputs(5079) <= '0';
    layer0_outputs(5080) <= '1';
    layer0_outputs(5081) <= '0';
    layer0_outputs(5082) <= not (a xor b);
    layer0_outputs(5083) <= '0';
    layer0_outputs(5084) <= not a or b;
    layer0_outputs(5085) <= a xor b;
    layer0_outputs(5086) <= a xor b;
    layer0_outputs(5087) <= b;
    layer0_outputs(5088) <= not (a and b);
    layer0_outputs(5089) <= not b;
    layer0_outputs(5090) <= not (a xor b);
    layer0_outputs(5091) <= a;
    layer0_outputs(5092) <= not a or b;
    layer0_outputs(5093) <= '1';
    layer0_outputs(5094) <= not a or b;
    layer0_outputs(5095) <= a;
    layer0_outputs(5096) <= a;
    layer0_outputs(5097) <= not b or a;
    layer0_outputs(5098) <= not (a and b);
    layer0_outputs(5099) <= b;
    layer0_outputs(5100) <= a and not b;
    layer0_outputs(5101) <= '1';
    layer0_outputs(5102) <= a or b;
    layer0_outputs(5103) <= b;
    layer0_outputs(5104) <= a and not b;
    layer0_outputs(5105) <= not (a xor b);
    layer0_outputs(5106) <= not b or a;
    layer0_outputs(5107) <= '1';
    layer0_outputs(5108) <= a and b;
    layer0_outputs(5109) <= not (a or b);
    layer0_outputs(5110) <= '0';
    layer0_outputs(5111) <= a;
    layer0_outputs(5112) <= b;
    layer0_outputs(5113) <= '1';
    layer0_outputs(5114) <= '0';
    layer0_outputs(5115) <= not b;
    layer0_outputs(5116) <= '0';
    layer0_outputs(5117) <= not b or a;
    layer0_outputs(5118) <= b;
    layer0_outputs(5119) <= not (a and b);
    layer1_outputs(0) <= a and b;
    layer1_outputs(1) <= not a;
    layer1_outputs(2) <= b and not a;
    layer1_outputs(3) <= '1';
    layer1_outputs(4) <= b;
    layer1_outputs(5) <= b and not a;
    layer1_outputs(6) <= not a or b;
    layer1_outputs(7) <= '1';
    layer1_outputs(8) <= b;
    layer1_outputs(9) <= not (a and b);
    layer1_outputs(10) <= not a;
    layer1_outputs(11) <= not a or b;
    layer1_outputs(12) <= b;
    layer1_outputs(13) <= '0';
    layer1_outputs(14) <= not (a and b);
    layer1_outputs(15) <= '0';
    layer1_outputs(16) <= a and not b;
    layer1_outputs(17) <= not a or b;
    layer1_outputs(18) <= not (a and b);
    layer1_outputs(19) <= b and not a;
    layer1_outputs(20) <= b and not a;
    layer1_outputs(21) <= a;
    layer1_outputs(22) <= not b;
    layer1_outputs(23) <= a and not b;
    layer1_outputs(24) <= '0';
    layer1_outputs(25) <= not (a and b);
    layer1_outputs(26) <= a or b;
    layer1_outputs(27) <= '1';
    layer1_outputs(28) <= b;
    layer1_outputs(29) <= not b or a;
    layer1_outputs(30) <= not b or a;
    layer1_outputs(31) <= not a or b;
    layer1_outputs(32) <= a or b;
    layer1_outputs(33) <= b and not a;
    layer1_outputs(34) <= not b or a;
    layer1_outputs(35) <= not (a or b);
    layer1_outputs(36) <= '0';
    layer1_outputs(37) <= not (a or b);
    layer1_outputs(38) <= not b or a;
    layer1_outputs(39) <= not b;
    layer1_outputs(40) <= '1';
    layer1_outputs(41) <= '0';
    layer1_outputs(42) <= a or b;
    layer1_outputs(43) <= '1';
    layer1_outputs(44) <= a and not b;
    layer1_outputs(45) <= b and not a;
    layer1_outputs(46) <= '0';
    layer1_outputs(47) <= '1';
    layer1_outputs(48) <= a or b;
    layer1_outputs(49) <= not (a or b);
    layer1_outputs(50) <= '1';
    layer1_outputs(51) <= b;
    layer1_outputs(52) <= a and b;
    layer1_outputs(53) <= b and not a;
    layer1_outputs(54) <= b;
    layer1_outputs(55) <= not (a and b);
    layer1_outputs(56) <= not b;
    layer1_outputs(57) <= a;
    layer1_outputs(58) <= a or b;
    layer1_outputs(59) <= not a;
    layer1_outputs(60) <= not b;
    layer1_outputs(61) <= '1';
    layer1_outputs(62) <= '0';
    layer1_outputs(63) <= not (a or b);
    layer1_outputs(64) <= not (a or b);
    layer1_outputs(65) <= '0';
    layer1_outputs(66) <= not (a and b);
    layer1_outputs(67) <= a and b;
    layer1_outputs(68) <= a and not b;
    layer1_outputs(69) <= '0';
    layer1_outputs(70) <= not (a or b);
    layer1_outputs(71) <= not a or b;
    layer1_outputs(72) <= a or b;
    layer1_outputs(73) <= not b;
    layer1_outputs(74) <= a and b;
    layer1_outputs(75) <= '0';
    layer1_outputs(76) <= a and not b;
    layer1_outputs(77) <= not (a or b);
    layer1_outputs(78) <= not a or b;
    layer1_outputs(79) <= not b;
    layer1_outputs(80) <= not (a or b);
    layer1_outputs(81) <= not (a and b);
    layer1_outputs(82) <= b;
    layer1_outputs(83) <= a or b;
    layer1_outputs(84) <= a and b;
    layer1_outputs(85) <= not (a and b);
    layer1_outputs(86) <= b;
    layer1_outputs(87) <= a;
    layer1_outputs(88) <= not (a xor b);
    layer1_outputs(89) <= a and b;
    layer1_outputs(90) <= not (a or b);
    layer1_outputs(91) <= not a;
    layer1_outputs(92) <= not b;
    layer1_outputs(93) <= '0';
    layer1_outputs(94) <= '0';
    layer1_outputs(95) <= not (a or b);
    layer1_outputs(96) <= b and not a;
    layer1_outputs(97) <= '1';
    layer1_outputs(98) <= not (a and b);
    layer1_outputs(99) <= not b or a;
    layer1_outputs(100) <= '0';
    layer1_outputs(101) <= '1';
    layer1_outputs(102) <= a;
    layer1_outputs(103) <= a xor b;
    layer1_outputs(104) <= a;
    layer1_outputs(105) <= not (a or b);
    layer1_outputs(106) <= a xor b;
    layer1_outputs(107) <= '1';
    layer1_outputs(108) <= '1';
    layer1_outputs(109) <= a;
    layer1_outputs(110) <= b and not a;
    layer1_outputs(111) <= not (a or b);
    layer1_outputs(112) <= b;
    layer1_outputs(113) <= '0';
    layer1_outputs(114) <= b;
    layer1_outputs(115) <= a and not b;
    layer1_outputs(116) <= a and not b;
    layer1_outputs(117) <= a and b;
    layer1_outputs(118) <= a xor b;
    layer1_outputs(119) <= b and not a;
    layer1_outputs(120) <= '0';
    layer1_outputs(121) <= b and not a;
    layer1_outputs(122) <= a;
    layer1_outputs(123) <= not (a or b);
    layer1_outputs(124) <= not (a xor b);
    layer1_outputs(125) <= not (a and b);
    layer1_outputs(126) <= not b or a;
    layer1_outputs(127) <= a and b;
    layer1_outputs(128) <= a xor b;
    layer1_outputs(129) <= not b;
    layer1_outputs(130) <= b and not a;
    layer1_outputs(131) <= b and not a;
    layer1_outputs(132) <= a and b;
    layer1_outputs(133) <= not a;
    layer1_outputs(134) <= a and b;
    layer1_outputs(135) <= '0';
    layer1_outputs(136) <= '0';
    layer1_outputs(137) <= a and not b;
    layer1_outputs(138) <= not (a or b);
    layer1_outputs(139) <= a and not b;
    layer1_outputs(140) <= b and not a;
    layer1_outputs(141) <= a and not b;
    layer1_outputs(142) <= not (a or b);
    layer1_outputs(143) <= b and not a;
    layer1_outputs(144) <= not a or b;
    layer1_outputs(145) <= not a;
    layer1_outputs(146) <= not (a xor b);
    layer1_outputs(147) <= b and not a;
    layer1_outputs(148) <= '0';
    layer1_outputs(149) <= a and b;
    layer1_outputs(150) <= not a or b;
    layer1_outputs(151) <= a and b;
    layer1_outputs(152) <= a and b;
    layer1_outputs(153) <= not (a or b);
    layer1_outputs(154) <= not (a or b);
    layer1_outputs(155) <= '1';
    layer1_outputs(156) <= a;
    layer1_outputs(157) <= a and b;
    layer1_outputs(158) <= not (a or b);
    layer1_outputs(159) <= '1';
    layer1_outputs(160) <= '1';
    layer1_outputs(161) <= not (a or b);
    layer1_outputs(162) <= not b or a;
    layer1_outputs(163) <= not a or b;
    layer1_outputs(164) <= not a or b;
    layer1_outputs(165) <= not a or b;
    layer1_outputs(166) <= b;
    layer1_outputs(167) <= '1';
    layer1_outputs(168) <= b;
    layer1_outputs(169) <= b;
    layer1_outputs(170) <= '1';
    layer1_outputs(171) <= a;
    layer1_outputs(172) <= a and b;
    layer1_outputs(173) <= a and not b;
    layer1_outputs(174) <= b;
    layer1_outputs(175) <= not b or a;
    layer1_outputs(176) <= not (a or b);
    layer1_outputs(177) <= b;
    layer1_outputs(178) <= a xor b;
    layer1_outputs(179) <= a or b;
    layer1_outputs(180) <= not (a or b);
    layer1_outputs(181) <= a and not b;
    layer1_outputs(182) <= a and not b;
    layer1_outputs(183) <= '0';
    layer1_outputs(184) <= b;
    layer1_outputs(185) <= not a;
    layer1_outputs(186) <= not (a xor b);
    layer1_outputs(187) <= not a or b;
    layer1_outputs(188) <= b and not a;
    layer1_outputs(189) <= not (a xor b);
    layer1_outputs(190) <= '1';
    layer1_outputs(191) <= not b or a;
    layer1_outputs(192) <= b and not a;
    layer1_outputs(193) <= b;
    layer1_outputs(194) <= a and not b;
    layer1_outputs(195) <= b;
    layer1_outputs(196) <= not a;
    layer1_outputs(197) <= a and not b;
    layer1_outputs(198) <= a;
    layer1_outputs(199) <= not (a or b);
    layer1_outputs(200) <= '1';
    layer1_outputs(201) <= a and b;
    layer1_outputs(202) <= not b or a;
    layer1_outputs(203) <= a and b;
    layer1_outputs(204) <= b;
    layer1_outputs(205) <= not a;
    layer1_outputs(206) <= not b or a;
    layer1_outputs(207) <= not (a and b);
    layer1_outputs(208) <= '1';
    layer1_outputs(209) <= b and not a;
    layer1_outputs(210) <= '1';
    layer1_outputs(211) <= b;
    layer1_outputs(212) <= not a;
    layer1_outputs(213) <= b and not a;
    layer1_outputs(214) <= '1';
    layer1_outputs(215) <= a and b;
    layer1_outputs(216) <= b and not a;
    layer1_outputs(217) <= a;
    layer1_outputs(218) <= not a or b;
    layer1_outputs(219) <= not b or a;
    layer1_outputs(220) <= not (a and b);
    layer1_outputs(221) <= '1';
    layer1_outputs(222) <= a or b;
    layer1_outputs(223) <= not a or b;
    layer1_outputs(224) <= not a;
    layer1_outputs(225) <= a or b;
    layer1_outputs(226) <= '1';
    layer1_outputs(227) <= not b or a;
    layer1_outputs(228) <= not b;
    layer1_outputs(229) <= not b or a;
    layer1_outputs(230) <= a and not b;
    layer1_outputs(231) <= not a or b;
    layer1_outputs(232) <= '1';
    layer1_outputs(233) <= not b;
    layer1_outputs(234) <= a and not b;
    layer1_outputs(235) <= b and not a;
    layer1_outputs(236) <= '0';
    layer1_outputs(237) <= not a;
    layer1_outputs(238) <= a and not b;
    layer1_outputs(239) <= a;
    layer1_outputs(240) <= not a or b;
    layer1_outputs(241) <= not (a or b);
    layer1_outputs(242) <= a or b;
    layer1_outputs(243) <= a and b;
    layer1_outputs(244) <= not a;
    layer1_outputs(245) <= '0';
    layer1_outputs(246) <= not a;
    layer1_outputs(247) <= not (a or b);
    layer1_outputs(248) <= b;
    layer1_outputs(249) <= b and not a;
    layer1_outputs(250) <= '0';
    layer1_outputs(251) <= not (a and b);
    layer1_outputs(252) <= not (a and b);
    layer1_outputs(253) <= a and b;
    layer1_outputs(254) <= a and b;
    layer1_outputs(255) <= a xor b;
    layer1_outputs(256) <= '0';
    layer1_outputs(257) <= '0';
    layer1_outputs(258) <= not (a or b);
    layer1_outputs(259) <= not b;
    layer1_outputs(260) <= '0';
    layer1_outputs(261) <= not b or a;
    layer1_outputs(262) <= not b;
    layer1_outputs(263) <= not (a and b);
    layer1_outputs(264) <= '1';
    layer1_outputs(265) <= a or b;
    layer1_outputs(266) <= '1';
    layer1_outputs(267) <= b and not a;
    layer1_outputs(268) <= a xor b;
    layer1_outputs(269) <= '0';
    layer1_outputs(270) <= not b;
    layer1_outputs(271) <= a;
    layer1_outputs(272) <= a;
    layer1_outputs(273) <= '1';
    layer1_outputs(274) <= '0';
    layer1_outputs(275) <= '1';
    layer1_outputs(276) <= a and not b;
    layer1_outputs(277) <= '1';
    layer1_outputs(278) <= not b;
    layer1_outputs(279) <= not a;
    layer1_outputs(280) <= not a or b;
    layer1_outputs(281) <= not b or a;
    layer1_outputs(282) <= not (a or b);
    layer1_outputs(283) <= not (a or b);
    layer1_outputs(284) <= a and not b;
    layer1_outputs(285) <= not a or b;
    layer1_outputs(286) <= a or b;
    layer1_outputs(287) <= a and b;
    layer1_outputs(288) <= a or b;
    layer1_outputs(289) <= '0';
    layer1_outputs(290) <= not a or b;
    layer1_outputs(291) <= not b;
    layer1_outputs(292) <= b;
    layer1_outputs(293) <= not b;
    layer1_outputs(294) <= b;
    layer1_outputs(295) <= not (a and b);
    layer1_outputs(296) <= not a or b;
    layer1_outputs(297) <= a;
    layer1_outputs(298) <= not (a and b);
    layer1_outputs(299) <= not (a or b);
    layer1_outputs(300) <= a;
    layer1_outputs(301) <= a;
    layer1_outputs(302) <= not a;
    layer1_outputs(303) <= not (a and b);
    layer1_outputs(304) <= not (a and b);
    layer1_outputs(305) <= a;
    layer1_outputs(306) <= a and b;
    layer1_outputs(307) <= '0';
    layer1_outputs(308) <= a and not b;
    layer1_outputs(309) <= not (a and b);
    layer1_outputs(310) <= b;
    layer1_outputs(311) <= b and not a;
    layer1_outputs(312) <= a and b;
    layer1_outputs(313) <= not b;
    layer1_outputs(314) <= a;
    layer1_outputs(315) <= not a or b;
    layer1_outputs(316) <= a and not b;
    layer1_outputs(317) <= a and b;
    layer1_outputs(318) <= not b or a;
    layer1_outputs(319) <= a or b;
    layer1_outputs(320) <= b;
    layer1_outputs(321) <= a;
    layer1_outputs(322) <= a and not b;
    layer1_outputs(323) <= not (a and b);
    layer1_outputs(324) <= not (a or b);
    layer1_outputs(325) <= not b;
    layer1_outputs(326) <= a and b;
    layer1_outputs(327) <= '1';
    layer1_outputs(328) <= a and b;
    layer1_outputs(329) <= not b;
    layer1_outputs(330) <= b and not a;
    layer1_outputs(331) <= not b;
    layer1_outputs(332) <= '0';
    layer1_outputs(333) <= not (a xor b);
    layer1_outputs(334) <= a and not b;
    layer1_outputs(335) <= a and not b;
    layer1_outputs(336) <= '0';
    layer1_outputs(337) <= not b;
    layer1_outputs(338) <= a and not b;
    layer1_outputs(339) <= not b;
    layer1_outputs(340) <= not b;
    layer1_outputs(341) <= a and b;
    layer1_outputs(342) <= not b;
    layer1_outputs(343) <= not a;
    layer1_outputs(344) <= a;
    layer1_outputs(345) <= a or b;
    layer1_outputs(346) <= b and not a;
    layer1_outputs(347) <= b and not a;
    layer1_outputs(348) <= '1';
    layer1_outputs(349) <= not (a or b);
    layer1_outputs(350) <= b and not a;
    layer1_outputs(351) <= '0';
    layer1_outputs(352) <= not b or a;
    layer1_outputs(353) <= not (a or b);
    layer1_outputs(354) <= not b;
    layer1_outputs(355) <= '1';
    layer1_outputs(356) <= not (a xor b);
    layer1_outputs(357) <= not b;
    layer1_outputs(358) <= not (a or b);
    layer1_outputs(359) <= a or b;
    layer1_outputs(360) <= '1';
    layer1_outputs(361) <= a or b;
    layer1_outputs(362) <= not b;
    layer1_outputs(363) <= '0';
    layer1_outputs(364) <= not a;
    layer1_outputs(365) <= a and b;
    layer1_outputs(366) <= not (a and b);
    layer1_outputs(367) <= not (a or b);
    layer1_outputs(368) <= '1';
    layer1_outputs(369) <= a;
    layer1_outputs(370) <= not (a or b);
    layer1_outputs(371) <= not (a and b);
    layer1_outputs(372) <= '0';
    layer1_outputs(373) <= not b or a;
    layer1_outputs(374) <= not (a or b);
    layer1_outputs(375) <= '0';
    layer1_outputs(376) <= not a or b;
    layer1_outputs(377) <= not b or a;
    layer1_outputs(378) <= '1';
    layer1_outputs(379) <= '0';
    layer1_outputs(380) <= a or b;
    layer1_outputs(381) <= not (a and b);
    layer1_outputs(382) <= a and not b;
    layer1_outputs(383) <= not (a xor b);
    layer1_outputs(384) <= b and not a;
    layer1_outputs(385) <= b and not a;
    layer1_outputs(386) <= b;
    layer1_outputs(387) <= a and not b;
    layer1_outputs(388) <= '0';
    layer1_outputs(389) <= a or b;
    layer1_outputs(390) <= a or b;
    layer1_outputs(391) <= not b;
    layer1_outputs(392) <= a and not b;
    layer1_outputs(393) <= '0';
    layer1_outputs(394) <= not (a or b);
    layer1_outputs(395) <= not b;
    layer1_outputs(396) <= not (a or b);
    layer1_outputs(397) <= '0';
    layer1_outputs(398) <= '0';
    layer1_outputs(399) <= not b or a;
    layer1_outputs(400) <= a and b;
    layer1_outputs(401) <= a or b;
    layer1_outputs(402) <= not (a and b);
    layer1_outputs(403) <= b;
    layer1_outputs(404) <= not b;
    layer1_outputs(405) <= a and not b;
    layer1_outputs(406) <= not (a or b);
    layer1_outputs(407) <= not a;
    layer1_outputs(408) <= not b or a;
    layer1_outputs(409) <= a;
    layer1_outputs(410) <= not a;
    layer1_outputs(411) <= a and not b;
    layer1_outputs(412) <= not a;
    layer1_outputs(413) <= not b or a;
    layer1_outputs(414) <= not a or b;
    layer1_outputs(415) <= not b;
    layer1_outputs(416) <= not a or b;
    layer1_outputs(417) <= not (a or b);
    layer1_outputs(418) <= a and b;
    layer1_outputs(419) <= not (a or b);
    layer1_outputs(420) <= a and not b;
    layer1_outputs(421) <= not b or a;
    layer1_outputs(422) <= not b or a;
    layer1_outputs(423) <= a and not b;
    layer1_outputs(424) <= not b;
    layer1_outputs(425) <= a and not b;
    layer1_outputs(426) <= not (a and b);
    layer1_outputs(427) <= a or b;
    layer1_outputs(428) <= b;
    layer1_outputs(429) <= a or b;
    layer1_outputs(430) <= b;
    layer1_outputs(431) <= a or b;
    layer1_outputs(432) <= not a or b;
    layer1_outputs(433) <= b and not a;
    layer1_outputs(434) <= not b or a;
    layer1_outputs(435) <= b;
    layer1_outputs(436) <= a and b;
    layer1_outputs(437) <= not (a and b);
    layer1_outputs(438) <= '0';
    layer1_outputs(439) <= not (a or b);
    layer1_outputs(440) <= b and not a;
    layer1_outputs(441) <= not (a xor b);
    layer1_outputs(442) <= not a or b;
    layer1_outputs(443) <= a and not b;
    layer1_outputs(444) <= not a;
    layer1_outputs(445) <= a and b;
    layer1_outputs(446) <= not (a or b);
    layer1_outputs(447) <= a and b;
    layer1_outputs(448) <= b;
    layer1_outputs(449) <= b;
    layer1_outputs(450) <= a or b;
    layer1_outputs(451) <= a and not b;
    layer1_outputs(452) <= '0';
    layer1_outputs(453) <= not a or b;
    layer1_outputs(454) <= b and not a;
    layer1_outputs(455) <= not b;
    layer1_outputs(456) <= b and not a;
    layer1_outputs(457) <= not b;
    layer1_outputs(458) <= b;
    layer1_outputs(459) <= '0';
    layer1_outputs(460) <= a or b;
    layer1_outputs(461) <= not a;
    layer1_outputs(462) <= b;
    layer1_outputs(463) <= '1';
    layer1_outputs(464) <= not (a or b);
    layer1_outputs(465) <= b and not a;
    layer1_outputs(466) <= a and not b;
    layer1_outputs(467) <= '0';
    layer1_outputs(468) <= a;
    layer1_outputs(469) <= a or b;
    layer1_outputs(470) <= '1';
    layer1_outputs(471) <= not a;
    layer1_outputs(472) <= a and not b;
    layer1_outputs(473) <= '1';
    layer1_outputs(474) <= not a;
    layer1_outputs(475) <= b and not a;
    layer1_outputs(476) <= b and not a;
    layer1_outputs(477) <= '1';
    layer1_outputs(478) <= not a or b;
    layer1_outputs(479) <= '0';
    layer1_outputs(480) <= a and b;
    layer1_outputs(481) <= not (a and b);
    layer1_outputs(482) <= a or b;
    layer1_outputs(483) <= '0';
    layer1_outputs(484) <= not (a or b);
    layer1_outputs(485) <= a or b;
    layer1_outputs(486) <= b;
    layer1_outputs(487) <= a and not b;
    layer1_outputs(488) <= not b;
    layer1_outputs(489) <= not b or a;
    layer1_outputs(490) <= not b or a;
    layer1_outputs(491) <= '0';
    layer1_outputs(492) <= not b or a;
    layer1_outputs(493) <= not a;
    layer1_outputs(494) <= a and not b;
    layer1_outputs(495) <= a and b;
    layer1_outputs(496) <= not b or a;
    layer1_outputs(497) <= '0';
    layer1_outputs(498) <= not (a and b);
    layer1_outputs(499) <= not a;
    layer1_outputs(500) <= not b or a;
    layer1_outputs(501) <= a and b;
    layer1_outputs(502) <= not b or a;
    layer1_outputs(503) <= not a;
    layer1_outputs(504) <= a or b;
    layer1_outputs(505) <= not b or a;
    layer1_outputs(506) <= not b;
    layer1_outputs(507) <= not (a or b);
    layer1_outputs(508) <= not a;
    layer1_outputs(509) <= not b or a;
    layer1_outputs(510) <= a and b;
    layer1_outputs(511) <= a and b;
    layer1_outputs(512) <= '0';
    layer1_outputs(513) <= b and not a;
    layer1_outputs(514) <= not b or a;
    layer1_outputs(515) <= b;
    layer1_outputs(516) <= not a or b;
    layer1_outputs(517) <= b and not a;
    layer1_outputs(518) <= a and b;
    layer1_outputs(519) <= a or b;
    layer1_outputs(520) <= not a or b;
    layer1_outputs(521) <= not b or a;
    layer1_outputs(522) <= not a;
    layer1_outputs(523) <= not b or a;
    layer1_outputs(524) <= not a;
    layer1_outputs(525) <= not b or a;
    layer1_outputs(526) <= not (a or b);
    layer1_outputs(527) <= not a or b;
    layer1_outputs(528) <= not a or b;
    layer1_outputs(529) <= not a or b;
    layer1_outputs(530) <= a;
    layer1_outputs(531) <= not (a or b);
    layer1_outputs(532) <= not (a or b);
    layer1_outputs(533) <= a and b;
    layer1_outputs(534) <= not b;
    layer1_outputs(535) <= not (a or b);
    layer1_outputs(536) <= a and not b;
    layer1_outputs(537) <= not a or b;
    layer1_outputs(538) <= a or b;
    layer1_outputs(539) <= a or b;
    layer1_outputs(540) <= not (a or b);
    layer1_outputs(541) <= not (a or b);
    layer1_outputs(542) <= '1';
    layer1_outputs(543) <= '1';
    layer1_outputs(544) <= not b or a;
    layer1_outputs(545) <= not b or a;
    layer1_outputs(546) <= not (a and b);
    layer1_outputs(547) <= not (a or b);
    layer1_outputs(548) <= not (a or b);
    layer1_outputs(549) <= '1';
    layer1_outputs(550) <= not (a and b);
    layer1_outputs(551) <= a;
    layer1_outputs(552) <= not (a and b);
    layer1_outputs(553) <= a and not b;
    layer1_outputs(554) <= b and not a;
    layer1_outputs(555) <= not b;
    layer1_outputs(556) <= not b or a;
    layer1_outputs(557) <= not b or a;
    layer1_outputs(558) <= a and b;
    layer1_outputs(559) <= a and not b;
    layer1_outputs(560) <= a or b;
    layer1_outputs(561) <= '0';
    layer1_outputs(562) <= '0';
    layer1_outputs(563) <= b;
    layer1_outputs(564) <= b;
    layer1_outputs(565) <= not (a and b);
    layer1_outputs(566) <= not a or b;
    layer1_outputs(567) <= not a or b;
    layer1_outputs(568) <= b and not a;
    layer1_outputs(569) <= not (a or b);
    layer1_outputs(570) <= not a or b;
    layer1_outputs(571) <= a and b;
    layer1_outputs(572) <= not b or a;
    layer1_outputs(573) <= not (a xor b);
    layer1_outputs(574) <= a and b;
    layer1_outputs(575) <= not a;
    layer1_outputs(576) <= a;
    layer1_outputs(577) <= a or b;
    layer1_outputs(578) <= '0';
    layer1_outputs(579) <= not b or a;
    layer1_outputs(580) <= a and not b;
    layer1_outputs(581) <= not a or b;
    layer1_outputs(582) <= a and b;
    layer1_outputs(583) <= '0';
    layer1_outputs(584) <= '0';
    layer1_outputs(585) <= '1';
    layer1_outputs(586) <= not a;
    layer1_outputs(587) <= not b or a;
    layer1_outputs(588) <= not b or a;
    layer1_outputs(589) <= not b;
    layer1_outputs(590) <= a or b;
    layer1_outputs(591) <= not a;
    layer1_outputs(592) <= '0';
    layer1_outputs(593) <= not a;
    layer1_outputs(594) <= not (a and b);
    layer1_outputs(595) <= not b;
    layer1_outputs(596) <= a and b;
    layer1_outputs(597) <= not b or a;
    layer1_outputs(598) <= a and b;
    layer1_outputs(599) <= a or b;
    layer1_outputs(600) <= not (a or b);
    layer1_outputs(601) <= not a or b;
    layer1_outputs(602) <= not a or b;
    layer1_outputs(603) <= '0';
    layer1_outputs(604) <= '1';
    layer1_outputs(605) <= not (a and b);
    layer1_outputs(606) <= b and not a;
    layer1_outputs(607) <= not b;
    layer1_outputs(608) <= not a;
    layer1_outputs(609) <= '1';
    layer1_outputs(610) <= not a;
    layer1_outputs(611) <= not (a or b);
    layer1_outputs(612) <= b;
    layer1_outputs(613) <= not (a and b);
    layer1_outputs(614) <= not a or b;
    layer1_outputs(615) <= not (a or b);
    layer1_outputs(616) <= a xor b;
    layer1_outputs(617) <= a and not b;
    layer1_outputs(618) <= not b or a;
    layer1_outputs(619) <= '1';
    layer1_outputs(620) <= not b;
    layer1_outputs(621) <= a or b;
    layer1_outputs(622) <= not a or b;
    layer1_outputs(623) <= a or b;
    layer1_outputs(624) <= not a;
    layer1_outputs(625) <= a and not b;
    layer1_outputs(626) <= not (a and b);
    layer1_outputs(627) <= a and b;
    layer1_outputs(628) <= not b;
    layer1_outputs(629) <= '1';
    layer1_outputs(630) <= '0';
    layer1_outputs(631) <= b and not a;
    layer1_outputs(632) <= '0';
    layer1_outputs(633) <= not (a and b);
    layer1_outputs(634) <= a xor b;
    layer1_outputs(635) <= not b or a;
    layer1_outputs(636) <= a and not b;
    layer1_outputs(637) <= a and not b;
    layer1_outputs(638) <= not (a and b);
    layer1_outputs(639) <= a and b;
    layer1_outputs(640) <= '0';
    layer1_outputs(641) <= not (a or b);
    layer1_outputs(642) <= b;
    layer1_outputs(643) <= '1';
    layer1_outputs(644) <= not (a or b);
    layer1_outputs(645) <= a and not b;
    layer1_outputs(646) <= not b or a;
    layer1_outputs(647) <= not a or b;
    layer1_outputs(648) <= not b or a;
    layer1_outputs(649) <= a and not b;
    layer1_outputs(650) <= a or b;
    layer1_outputs(651) <= not a;
    layer1_outputs(652) <= a or b;
    layer1_outputs(653) <= a and b;
    layer1_outputs(654) <= not (a or b);
    layer1_outputs(655) <= not a or b;
    layer1_outputs(656) <= a and not b;
    layer1_outputs(657) <= not (a or b);
    layer1_outputs(658) <= a;
    layer1_outputs(659) <= a and not b;
    layer1_outputs(660) <= not (a and b);
    layer1_outputs(661) <= a and not b;
    layer1_outputs(662) <= a and not b;
    layer1_outputs(663) <= a;
    layer1_outputs(664) <= not (a and b);
    layer1_outputs(665) <= '0';
    layer1_outputs(666) <= a xor b;
    layer1_outputs(667) <= not (a and b);
    layer1_outputs(668) <= not b or a;
    layer1_outputs(669) <= a;
    layer1_outputs(670) <= not a;
    layer1_outputs(671) <= a and not b;
    layer1_outputs(672) <= a or b;
    layer1_outputs(673) <= '1';
    layer1_outputs(674) <= '0';
    layer1_outputs(675) <= b and not a;
    layer1_outputs(676) <= a and not b;
    layer1_outputs(677) <= b;
    layer1_outputs(678) <= not b;
    layer1_outputs(679) <= b and not a;
    layer1_outputs(680) <= a;
    layer1_outputs(681) <= a or b;
    layer1_outputs(682) <= '0';
    layer1_outputs(683) <= '0';
    layer1_outputs(684) <= not a or b;
    layer1_outputs(685) <= b;
    layer1_outputs(686) <= not b;
    layer1_outputs(687) <= a and b;
    layer1_outputs(688) <= a and b;
    layer1_outputs(689) <= a and b;
    layer1_outputs(690) <= not a;
    layer1_outputs(691) <= a and not b;
    layer1_outputs(692) <= not (a and b);
    layer1_outputs(693) <= a and b;
    layer1_outputs(694) <= a and b;
    layer1_outputs(695) <= a or b;
    layer1_outputs(696) <= a;
    layer1_outputs(697) <= a and not b;
    layer1_outputs(698) <= b and not a;
    layer1_outputs(699) <= '0';
    layer1_outputs(700) <= not (a and b);
    layer1_outputs(701) <= '1';
    layer1_outputs(702) <= '0';
    layer1_outputs(703) <= not (a and b);
    layer1_outputs(704) <= a;
    layer1_outputs(705) <= a;
    layer1_outputs(706) <= not b or a;
    layer1_outputs(707) <= a and not b;
    layer1_outputs(708) <= not a or b;
    layer1_outputs(709) <= not b;
    layer1_outputs(710) <= '1';
    layer1_outputs(711) <= a or b;
    layer1_outputs(712) <= a;
    layer1_outputs(713) <= not a;
    layer1_outputs(714) <= b and not a;
    layer1_outputs(715) <= '0';
    layer1_outputs(716) <= a;
    layer1_outputs(717) <= not a;
    layer1_outputs(718) <= b;
    layer1_outputs(719) <= not a;
    layer1_outputs(720) <= b;
    layer1_outputs(721) <= not (a and b);
    layer1_outputs(722) <= a xor b;
    layer1_outputs(723) <= not (a xor b);
    layer1_outputs(724) <= a;
    layer1_outputs(725) <= a and not b;
    layer1_outputs(726) <= '0';
    layer1_outputs(727) <= '0';
    layer1_outputs(728) <= b and not a;
    layer1_outputs(729) <= not b;
    layer1_outputs(730) <= '1';
    layer1_outputs(731) <= not (a or b);
    layer1_outputs(732) <= b and not a;
    layer1_outputs(733) <= a and b;
    layer1_outputs(734) <= not a;
    layer1_outputs(735) <= a and not b;
    layer1_outputs(736) <= not (a or b);
    layer1_outputs(737) <= '0';
    layer1_outputs(738) <= '0';
    layer1_outputs(739) <= not b;
    layer1_outputs(740) <= not b;
    layer1_outputs(741) <= a and b;
    layer1_outputs(742) <= a xor b;
    layer1_outputs(743) <= not b or a;
    layer1_outputs(744) <= '0';
    layer1_outputs(745) <= not b;
    layer1_outputs(746) <= not b or a;
    layer1_outputs(747) <= '0';
    layer1_outputs(748) <= a and not b;
    layer1_outputs(749) <= not (a or b);
    layer1_outputs(750) <= b;
    layer1_outputs(751) <= not (a and b);
    layer1_outputs(752) <= a and b;
    layer1_outputs(753) <= not a or b;
    layer1_outputs(754) <= not a;
    layer1_outputs(755) <= a;
    layer1_outputs(756) <= '1';
    layer1_outputs(757) <= a or b;
    layer1_outputs(758) <= a or b;
    layer1_outputs(759) <= '1';
    layer1_outputs(760) <= not b;
    layer1_outputs(761) <= a xor b;
    layer1_outputs(762) <= a and not b;
    layer1_outputs(763) <= not a;
    layer1_outputs(764) <= b and not a;
    layer1_outputs(765) <= b and not a;
    layer1_outputs(766) <= not a or b;
    layer1_outputs(767) <= b;
    layer1_outputs(768) <= a and not b;
    layer1_outputs(769) <= not b;
    layer1_outputs(770) <= '1';
    layer1_outputs(771) <= a and not b;
    layer1_outputs(772) <= not (a and b);
    layer1_outputs(773) <= not b;
    layer1_outputs(774) <= '0';
    layer1_outputs(775) <= not (a and b);
    layer1_outputs(776) <= b and not a;
    layer1_outputs(777) <= not b or a;
    layer1_outputs(778) <= a;
    layer1_outputs(779) <= not b;
    layer1_outputs(780) <= '1';
    layer1_outputs(781) <= not a or b;
    layer1_outputs(782) <= a and not b;
    layer1_outputs(783) <= '0';
    layer1_outputs(784) <= b;
    layer1_outputs(785) <= a;
    layer1_outputs(786) <= a and not b;
    layer1_outputs(787) <= '1';
    layer1_outputs(788) <= not a or b;
    layer1_outputs(789) <= a or b;
    layer1_outputs(790) <= '1';
    layer1_outputs(791) <= a and b;
    layer1_outputs(792) <= not a or b;
    layer1_outputs(793) <= a xor b;
    layer1_outputs(794) <= b and not a;
    layer1_outputs(795) <= not b;
    layer1_outputs(796) <= not a or b;
    layer1_outputs(797) <= a and not b;
    layer1_outputs(798) <= a;
    layer1_outputs(799) <= not b;
    layer1_outputs(800) <= a or b;
    layer1_outputs(801) <= a and not b;
    layer1_outputs(802) <= b and not a;
    layer1_outputs(803) <= '0';
    layer1_outputs(804) <= a and b;
    layer1_outputs(805) <= not a or b;
    layer1_outputs(806) <= '0';
    layer1_outputs(807) <= not a or b;
    layer1_outputs(808) <= not b;
    layer1_outputs(809) <= not (a and b);
    layer1_outputs(810) <= a or b;
    layer1_outputs(811) <= not a or b;
    layer1_outputs(812) <= '1';
    layer1_outputs(813) <= a or b;
    layer1_outputs(814) <= a and not b;
    layer1_outputs(815) <= not a;
    layer1_outputs(816) <= not (a or b);
    layer1_outputs(817) <= b and not a;
    layer1_outputs(818) <= a;
    layer1_outputs(819) <= a;
    layer1_outputs(820) <= not b or a;
    layer1_outputs(821) <= a;
    layer1_outputs(822) <= b;
    layer1_outputs(823) <= not (a xor b);
    layer1_outputs(824) <= not a or b;
    layer1_outputs(825) <= not b;
    layer1_outputs(826) <= a or b;
    layer1_outputs(827) <= '0';
    layer1_outputs(828) <= not (a and b);
    layer1_outputs(829) <= not (a and b);
    layer1_outputs(830) <= not b;
    layer1_outputs(831) <= not b or a;
    layer1_outputs(832) <= not b or a;
    layer1_outputs(833) <= a or b;
    layer1_outputs(834) <= a and b;
    layer1_outputs(835) <= not a or b;
    layer1_outputs(836) <= a;
    layer1_outputs(837) <= '0';
    layer1_outputs(838) <= b;
    layer1_outputs(839) <= not (a or b);
    layer1_outputs(840) <= a;
    layer1_outputs(841) <= not (a or b);
    layer1_outputs(842) <= b and not a;
    layer1_outputs(843) <= a xor b;
    layer1_outputs(844) <= a xor b;
    layer1_outputs(845) <= a;
    layer1_outputs(846) <= not a;
    layer1_outputs(847) <= not (a xor b);
    layer1_outputs(848) <= '1';
    layer1_outputs(849) <= '1';
    layer1_outputs(850) <= a and not b;
    layer1_outputs(851) <= '0';
    layer1_outputs(852) <= not b or a;
    layer1_outputs(853) <= '1';
    layer1_outputs(854) <= a and not b;
    layer1_outputs(855) <= not (a or b);
    layer1_outputs(856) <= b;
    layer1_outputs(857) <= not b;
    layer1_outputs(858) <= b;
    layer1_outputs(859) <= '1';
    layer1_outputs(860) <= not (a or b);
    layer1_outputs(861) <= not a or b;
    layer1_outputs(862) <= b;
    layer1_outputs(863) <= '1';
    layer1_outputs(864) <= b;
    layer1_outputs(865) <= not a or b;
    layer1_outputs(866) <= not (a and b);
    layer1_outputs(867) <= a or b;
    layer1_outputs(868) <= b and not a;
    layer1_outputs(869) <= '0';
    layer1_outputs(870) <= '1';
    layer1_outputs(871) <= not (a or b);
    layer1_outputs(872) <= b;
    layer1_outputs(873) <= not a or b;
    layer1_outputs(874) <= a;
    layer1_outputs(875) <= not a or b;
    layer1_outputs(876) <= not (a and b);
    layer1_outputs(877) <= '0';
    layer1_outputs(878) <= a;
    layer1_outputs(879) <= b and not a;
    layer1_outputs(880) <= a and not b;
    layer1_outputs(881) <= '1';
    layer1_outputs(882) <= a and not b;
    layer1_outputs(883) <= not a;
    layer1_outputs(884) <= a and not b;
    layer1_outputs(885) <= not b or a;
    layer1_outputs(886) <= not a;
    layer1_outputs(887) <= '1';
    layer1_outputs(888) <= not (a xor b);
    layer1_outputs(889) <= a and not b;
    layer1_outputs(890) <= '0';
    layer1_outputs(891) <= not (a or b);
    layer1_outputs(892) <= '1';
    layer1_outputs(893) <= not (a and b);
    layer1_outputs(894) <= b;
    layer1_outputs(895) <= not a or b;
    layer1_outputs(896) <= a;
    layer1_outputs(897) <= b;
    layer1_outputs(898) <= not b;
    layer1_outputs(899) <= not b;
    layer1_outputs(900) <= not (a or b);
    layer1_outputs(901) <= '0';
    layer1_outputs(902) <= not (a xor b);
    layer1_outputs(903) <= not (a or b);
    layer1_outputs(904) <= not a;
    layer1_outputs(905) <= not a;
    layer1_outputs(906) <= not a;
    layer1_outputs(907) <= b and not a;
    layer1_outputs(908) <= a;
    layer1_outputs(909) <= '1';
    layer1_outputs(910) <= not b;
    layer1_outputs(911) <= not a or b;
    layer1_outputs(912) <= not a;
    layer1_outputs(913) <= not a;
    layer1_outputs(914) <= not a or b;
    layer1_outputs(915) <= not a;
    layer1_outputs(916) <= a or b;
    layer1_outputs(917) <= b and not a;
    layer1_outputs(918) <= not (a or b);
    layer1_outputs(919) <= a or b;
    layer1_outputs(920) <= a and b;
    layer1_outputs(921) <= not (a or b);
    layer1_outputs(922) <= not (a and b);
    layer1_outputs(923) <= '1';
    layer1_outputs(924) <= a and b;
    layer1_outputs(925) <= not b or a;
    layer1_outputs(926) <= b;
    layer1_outputs(927) <= not (a xor b);
    layer1_outputs(928) <= a or b;
    layer1_outputs(929) <= '0';
    layer1_outputs(930) <= a or b;
    layer1_outputs(931) <= b and not a;
    layer1_outputs(932) <= b and not a;
    layer1_outputs(933) <= a or b;
    layer1_outputs(934) <= a and not b;
    layer1_outputs(935) <= '0';
    layer1_outputs(936) <= b and not a;
    layer1_outputs(937) <= not (a and b);
    layer1_outputs(938) <= not b or a;
    layer1_outputs(939) <= not b;
    layer1_outputs(940) <= not (a and b);
    layer1_outputs(941) <= a or b;
    layer1_outputs(942) <= a and not b;
    layer1_outputs(943) <= '0';
    layer1_outputs(944) <= '0';
    layer1_outputs(945) <= not (a xor b);
    layer1_outputs(946) <= not (a and b);
    layer1_outputs(947) <= b and not a;
    layer1_outputs(948) <= '1';
    layer1_outputs(949) <= a and b;
    layer1_outputs(950) <= a and b;
    layer1_outputs(951) <= '1';
    layer1_outputs(952) <= not a;
    layer1_outputs(953) <= not a or b;
    layer1_outputs(954) <= not b or a;
    layer1_outputs(955) <= not b;
    layer1_outputs(956) <= not (a and b);
    layer1_outputs(957) <= b and not a;
    layer1_outputs(958) <= not (a and b);
    layer1_outputs(959) <= b and not a;
    layer1_outputs(960) <= b;
    layer1_outputs(961) <= a and not b;
    layer1_outputs(962) <= a and not b;
    layer1_outputs(963) <= not a;
    layer1_outputs(964) <= b;
    layer1_outputs(965) <= b and not a;
    layer1_outputs(966) <= not (a or b);
    layer1_outputs(967) <= a and b;
    layer1_outputs(968) <= not a or b;
    layer1_outputs(969) <= a;
    layer1_outputs(970) <= b;
    layer1_outputs(971) <= '1';
    layer1_outputs(972) <= not b;
    layer1_outputs(973) <= '0';
    layer1_outputs(974) <= '0';
    layer1_outputs(975) <= not b;
    layer1_outputs(976) <= a or b;
    layer1_outputs(977) <= not a or b;
    layer1_outputs(978) <= not a;
    layer1_outputs(979) <= not (a or b);
    layer1_outputs(980) <= not (a or b);
    layer1_outputs(981) <= b;
    layer1_outputs(982) <= '1';
    layer1_outputs(983) <= not a or b;
    layer1_outputs(984) <= not (a or b);
    layer1_outputs(985) <= a and b;
    layer1_outputs(986) <= not b;
    layer1_outputs(987) <= not (a and b);
    layer1_outputs(988) <= not a;
    layer1_outputs(989) <= b and not a;
    layer1_outputs(990) <= a and b;
    layer1_outputs(991) <= '1';
    layer1_outputs(992) <= a and not b;
    layer1_outputs(993) <= not (a or b);
    layer1_outputs(994) <= not (a and b);
    layer1_outputs(995) <= '1';
    layer1_outputs(996) <= a and b;
    layer1_outputs(997) <= a xor b;
    layer1_outputs(998) <= not (a and b);
    layer1_outputs(999) <= '0';
    layer1_outputs(1000) <= '0';
    layer1_outputs(1001) <= a and b;
    layer1_outputs(1002) <= a and b;
    layer1_outputs(1003) <= not (a xor b);
    layer1_outputs(1004) <= b and not a;
    layer1_outputs(1005) <= not (a or b);
    layer1_outputs(1006) <= a or b;
    layer1_outputs(1007) <= a and not b;
    layer1_outputs(1008) <= not b or a;
    layer1_outputs(1009) <= b and not a;
    layer1_outputs(1010) <= a or b;
    layer1_outputs(1011) <= not a;
    layer1_outputs(1012) <= not b or a;
    layer1_outputs(1013) <= '1';
    layer1_outputs(1014) <= '0';
    layer1_outputs(1015) <= not (a or b);
    layer1_outputs(1016) <= a and not b;
    layer1_outputs(1017) <= not (a or b);
    layer1_outputs(1018) <= not (a or b);
    layer1_outputs(1019) <= a or b;
    layer1_outputs(1020) <= not b;
    layer1_outputs(1021) <= not a or b;
    layer1_outputs(1022) <= not (a and b);
    layer1_outputs(1023) <= '0';
    layer1_outputs(1024) <= '1';
    layer1_outputs(1025) <= a and b;
    layer1_outputs(1026) <= '0';
    layer1_outputs(1027) <= not a or b;
    layer1_outputs(1028) <= not a;
    layer1_outputs(1029) <= a or b;
    layer1_outputs(1030) <= not (a and b);
    layer1_outputs(1031) <= b and not a;
    layer1_outputs(1032) <= b;
    layer1_outputs(1033) <= not (a or b);
    layer1_outputs(1034) <= not b or a;
    layer1_outputs(1035) <= not (a and b);
    layer1_outputs(1036) <= a or b;
    layer1_outputs(1037) <= '1';
    layer1_outputs(1038) <= a and not b;
    layer1_outputs(1039) <= '1';
    layer1_outputs(1040) <= a;
    layer1_outputs(1041) <= a;
    layer1_outputs(1042) <= '0';
    layer1_outputs(1043) <= '0';
    layer1_outputs(1044) <= a and b;
    layer1_outputs(1045) <= a;
    layer1_outputs(1046) <= a and not b;
    layer1_outputs(1047) <= a and not b;
    layer1_outputs(1048) <= b and not a;
    layer1_outputs(1049) <= '0';
    layer1_outputs(1050) <= not (a and b);
    layer1_outputs(1051) <= b;
    layer1_outputs(1052) <= a or b;
    layer1_outputs(1053) <= not a or b;
    layer1_outputs(1054) <= '1';
    layer1_outputs(1055) <= a and not b;
    layer1_outputs(1056) <= not a or b;
    layer1_outputs(1057) <= not (a and b);
    layer1_outputs(1058) <= a xor b;
    layer1_outputs(1059) <= a and b;
    layer1_outputs(1060) <= a and not b;
    layer1_outputs(1061) <= not a;
    layer1_outputs(1062) <= b and not a;
    layer1_outputs(1063) <= not (a and b);
    layer1_outputs(1064) <= a and not b;
    layer1_outputs(1065) <= not b or a;
    layer1_outputs(1066) <= a xor b;
    layer1_outputs(1067) <= not b;
    layer1_outputs(1068) <= not (a or b);
    layer1_outputs(1069) <= a or b;
    layer1_outputs(1070) <= not (a and b);
    layer1_outputs(1071) <= b;
    layer1_outputs(1072) <= not (a and b);
    layer1_outputs(1073) <= '1';
    layer1_outputs(1074) <= '0';
    layer1_outputs(1075) <= not (a and b);
    layer1_outputs(1076) <= '1';
    layer1_outputs(1077) <= not (a xor b);
    layer1_outputs(1078) <= not (a or b);
    layer1_outputs(1079) <= not a or b;
    layer1_outputs(1080) <= '0';
    layer1_outputs(1081) <= a;
    layer1_outputs(1082) <= not a;
    layer1_outputs(1083) <= not a;
    layer1_outputs(1084) <= not (a and b);
    layer1_outputs(1085) <= '0';
    layer1_outputs(1086) <= a;
    layer1_outputs(1087) <= a or b;
    layer1_outputs(1088) <= '1';
    layer1_outputs(1089) <= a xor b;
    layer1_outputs(1090) <= b;
    layer1_outputs(1091) <= a and b;
    layer1_outputs(1092) <= a or b;
    layer1_outputs(1093) <= a and not b;
    layer1_outputs(1094) <= not a or b;
    layer1_outputs(1095) <= not a;
    layer1_outputs(1096) <= not a or b;
    layer1_outputs(1097) <= not b;
    layer1_outputs(1098) <= not (a xor b);
    layer1_outputs(1099) <= '1';
    layer1_outputs(1100) <= not (a and b);
    layer1_outputs(1101) <= not b;
    layer1_outputs(1102) <= not a or b;
    layer1_outputs(1103) <= '0';
    layer1_outputs(1104) <= '0';
    layer1_outputs(1105) <= '1';
    layer1_outputs(1106) <= not a;
    layer1_outputs(1107) <= not (a and b);
    layer1_outputs(1108) <= a or b;
    layer1_outputs(1109) <= '0';
    layer1_outputs(1110) <= not a;
    layer1_outputs(1111) <= not (a and b);
    layer1_outputs(1112) <= not a or b;
    layer1_outputs(1113) <= not (a or b);
    layer1_outputs(1114) <= not (a and b);
    layer1_outputs(1115) <= not a or b;
    layer1_outputs(1116) <= a or b;
    layer1_outputs(1117) <= a and b;
    layer1_outputs(1118) <= not b;
    layer1_outputs(1119) <= a xor b;
    layer1_outputs(1120) <= a and not b;
    layer1_outputs(1121) <= b;
    layer1_outputs(1122) <= not a or b;
    layer1_outputs(1123) <= not b;
    layer1_outputs(1124) <= a xor b;
    layer1_outputs(1125) <= a and not b;
    layer1_outputs(1126) <= '0';
    layer1_outputs(1127) <= a;
    layer1_outputs(1128) <= a;
    layer1_outputs(1129) <= not b;
    layer1_outputs(1130) <= '1';
    layer1_outputs(1131) <= not (a or b);
    layer1_outputs(1132) <= not b;
    layer1_outputs(1133) <= not a or b;
    layer1_outputs(1134) <= not a;
    layer1_outputs(1135) <= not a or b;
    layer1_outputs(1136) <= '1';
    layer1_outputs(1137) <= '1';
    layer1_outputs(1138) <= a xor b;
    layer1_outputs(1139) <= '0';
    layer1_outputs(1140) <= b and not a;
    layer1_outputs(1141) <= b and not a;
    layer1_outputs(1142) <= b;
    layer1_outputs(1143) <= '0';
    layer1_outputs(1144) <= '0';
    layer1_outputs(1145) <= a;
    layer1_outputs(1146) <= not b;
    layer1_outputs(1147) <= not (a and b);
    layer1_outputs(1148) <= '0';
    layer1_outputs(1149) <= not a or b;
    layer1_outputs(1150) <= b;
    layer1_outputs(1151) <= not b;
    layer1_outputs(1152) <= not (a and b);
    layer1_outputs(1153) <= a and b;
    layer1_outputs(1154) <= not b or a;
    layer1_outputs(1155) <= '1';
    layer1_outputs(1156) <= '0';
    layer1_outputs(1157) <= not (a or b);
    layer1_outputs(1158) <= a;
    layer1_outputs(1159) <= '0';
    layer1_outputs(1160) <= a and b;
    layer1_outputs(1161) <= '1';
    layer1_outputs(1162) <= a xor b;
    layer1_outputs(1163) <= a and b;
    layer1_outputs(1164) <= a and b;
    layer1_outputs(1165) <= not (a xor b);
    layer1_outputs(1166) <= a xor b;
    layer1_outputs(1167) <= not a or b;
    layer1_outputs(1168) <= '0';
    layer1_outputs(1169) <= '0';
    layer1_outputs(1170) <= a or b;
    layer1_outputs(1171) <= '1';
    layer1_outputs(1172) <= a;
    layer1_outputs(1173) <= not a;
    layer1_outputs(1174) <= '0';
    layer1_outputs(1175) <= not (a or b);
    layer1_outputs(1176) <= '1';
    layer1_outputs(1177) <= not (a or b);
    layer1_outputs(1178) <= b;
    layer1_outputs(1179) <= '0';
    layer1_outputs(1180) <= a or b;
    layer1_outputs(1181) <= not b or a;
    layer1_outputs(1182) <= not a;
    layer1_outputs(1183) <= not b or a;
    layer1_outputs(1184) <= not b;
    layer1_outputs(1185) <= b;
    layer1_outputs(1186) <= a xor b;
    layer1_outputs(1187) <= '1';
    layer1_outputs(1188) <= a xor b;
    layer1_outputs(1189) <= '1';
    layer1_outputs(1190) <= a or b;
    layer1_outputs(1191) <= not b;
    layer1_outputs(1192) <= b and not a;
    layer1_outputs(1193) <= b and not a;
    layer1_outputs(1194) <= not (a and b);
    layer1_outputs(1195) <= a and b;
    layer1_outputs(1196) <= not (a and b);
    layer1_outputs(1197) <= '0';
    layer1_outputs(1198) <= a xor b;
    layer1_outputs(1199) <= a or b;
    layer1_outputs(1200) <= not (a and b);
    layer1_outputs(1201) <= not (a or b);
    layer1_outputs(1202) <= not a;
    layer1_outputs(1203) <= a and b;
    layer1_outputs(1204) <= not b;
    layer1_outputs(1205) <= a and b;
    layer1_outputs(1206) <= b and not a;
    layer1_outputs(1207) <= a;
    layer1_outputs(1208) <= a xor b;
    layer1_outputs(1209) <= a and not b;
    layer1_outputs(1210) <= a;
    layer1_outputs(1211) <= '0';
    layer1_outputs(1212) <= '1';
    layer1_outputs(1213) <= '0';
    layer1_outputs(1214) <= not a or b;
    layer1_outputs(1215) <= '0';
    layer1_outputs(1216) <= a and b;
    layer1_outputs(1217) <= a and b;
    layer1_outputs(1218) <= not (a and b);
    layer1_outputs(1219) <= '0';
    layer1_outputs(1220) <= not (a xor b);
    layer1_outputs(1221) <= '0';
    layer1_outputs(1222) <= b and not a;
    layer1_outputs(1223) <= a;
    layer1_outputs(1224) <= b and not a;
    layer1_outputs(1225) <= a and not b;
    layer1_outputs(1226) <= not a;
    layer1_outputs(1227) <= not (a and b);
    layer1_outputs(1228) <= not a or b;
    layer1_outputs(1229) <= not (a and b);
    layer1_outputs(1230) <= '0';
    layer1_outputs(1231) <= '1';
    layer1_outputs(1232) <= not b or a;
    layer1_outputs(1233) <= not b;
    layer1_outputs(1234) <= not a or b;
    layer1_outputs(1235) <= '0';
    layer1_outputs(1236) <= not (a or b);
    layer1_outputs(1237) <= not (a or b);
    layer1_outputs(1238) <= b and not a;
    layer1_outputs(1239) <= '1';
    layer1_outputs(1240) <= '1';
    layer1_outputs(1241) <= a and not b;
    layer1_outputs(1242) <= not b;
    layer1_outputs(1243) <= a and not b;
    layer1_outputs(1244) <= not b or a;
    layer1_outputs(1245) <= '1';
    layer1_outputs(1246) <= a and not b;
    layer1_outputs(1247) <= '0';
    layer1_outputs(1248) <= not b or a;
    layer1_outputs(1249) <= not (a xor b);
    layer1_outputs(1250) <= not a or b;
    layer1_outputs(1251) <= a and b;
    layer1_outputs(1252) <= not (a or b);
    layer1_outputs(1253) <= a xor b;
    layer1_outputs(1254) <= not (a and b);
    layer1_outputs(1255) <= '1';
    layer1_outputs(1256) <= b and not a;
    layer1_outputs(1257) <= not a or b;
    layer1_outputs(1258) <= not a or b;
    layer1_outputs(1259) <= b and not a;
    layer1_outputs(1260) <= not a or b;
    layer1_outputs(1261) <= '1';
    layer1_outputs(1262) <= not b;
    layer1_outputs(1263) <= '0';
    layer1_outputs(1264) <= not (a or b);
    layer1_outputs(1265) <= not (a or b);
    layer1_outputs(1266) <= a;
    layer1_outputs(1267) <= not (a xor b);
    layer1_outputs(1268) <= '1';
    layer1_outputs(1269) <= not b or a;
    layer1_outputs(1270) <= a and not b;
    layer1_outputs(1271) <= a;
    layer1_outputs(1272) <= not (a or b);
    layer1_outputs(1273) <= not a;
    layer1_outputs(1274) <= not a;
    layer1_outputs(1275) <= b and not a;
    layer1_outputs(1276) <= not (a and b);
    layer1_outputs(1277) <= a and b;
    layer1_outputs(1278) <= a and b;
    layer1_outputs(1279) <= not (a and b);
    layer1_outputs(1280) <= not b;
    layer1_outputs(1281) <= '1';
    layer1_outputs(1282) <= a and not b;
    layer1_outputs(1283) <= not a;
    layer1_outputs(1284) <= a or b;
    layer1_outputs(1285) <= not b or a;
    layer1_outputs(1286) <= a or b;
    layer1_outputs(1287) <= not b;
    layer1_outputs(1288) <= not b;
    layer1_outputs(1289) <= not (a or b);
    layer1_outputs(1290) <= a;
    layer1_outputs(1291) <= '1';
    layer1_outputs(1292) <= '1';
    layer1_outputs(1293) <= not (a or b);
    layer1_outputs(1294) <= '0';
    layer1_outputs(1295) <= not b;
    layer1_outputs(1296) <= not (a and b);
    layer1_outputs(1297) <= a and not b;
    layer1_outputs(1298) <= not a;
    layer1_outputs(1299) <= not a or b;
    layer1_outputs(1300) <= b and not a;
    layer1_outputs(1301) <= a or b;
    layer1_outputs(1302) <= not (a xor b);
    layer1_outputs(1303) <= '1';
    layer1_outputs(1304) <= b;
    layer1_outputs(1305) <= not (a or b);
    layer1_outputs(1306) <= '1';
    layer1_outputs(1307) <= b and not a;
    layer1_outputs(1308) <= not a or b;
    layer1_outputs(1309) <= not b or a;
    layer1_outputs(1310) <= not (a and b);
    layer1_outputs(1311) <= a and b;
    layer1_outputs(1312) <= not a or b;
    layer1_outputs(1313) <= a xor b;
    layer1_outputs(1314) <= a or b;
    layer1_outputs(1315) <= '1';
    layer1_outputs(1316) <= '0';
    layer1_outputs(1317) <= '0';
    layer1_outputs(1318) <= not (a and b);
    layer1_outputs(1319) <= not b;
    layer1_outputs(1320) <= b;
    layer1_outputs(1321) <= a;
    layer1_outputs(1322) <= not b;
    layer1_outputs(1323) <= b;
    layer1_outputs(1324) <= not a or b;
    layer1_outputs(1325) <= a or b;
    layer1_outputs(1326) <= a or b;
    layer1_outputs(1327) <= a or b;
    layer1_outputs(1328) <= a and not b;
    layer1_outputs(1329) <= '1';
    layer1_outputs(1330) <= a;
    layer1_outputs(1331) <= a;
    layer1_outputs(1332) <= not a;
    layer1_outputs(1333) <= not (a and b);
    layer1_outputs(1334) <= b;
    layer1_outputs(1335) <= a;
    layer1_outputs(1336) <= a and b;
    layer1_outputs(1337) <= '1';
    layer1_outputs(1338) <= not b or a;
    layer1_outputs(1339) <= not a or b;
    layer1_outputs(1340) <= a xor b;
    layer1_outputs(1341) <= not (a or b);
    layer1_outputs(1342) <= not b;
    layer1_outputs(1343) <= a;
    layer1_outputs(1344) <= '1';
    layer1_outputs(1345) <= b and not a;
    layer1_outputs(1346) <= not a or b;
    layer1_outputs(1347) <= '1';
    layer1_outputs(1348) <= '0';
    layer1_outputs(1349) <= b;
    layer1_outputs(1350) <= not b or a;
    layer1_outputs(1351) <= b and not a;
    layer1_outputs(1352) <= '0';
    layer1_outputs(1353) <= a and b;
    layer1_outputs(1354) <= not (a or b);
    layer1_outputs(1355) <= a and not b;
    layer1_outputs(1356) <= a or b;
    layer1_outputs(1357) <= not (a and b);
    layer1_outputs(1358) <= a xor b;
    layer1_outputs(1359) <= not (a or b);
    layer1_outputs(1360) <= not a;
    layer1_outputs(1361) <= a xor b;
    layer1_outputs(1362) <= a;
    layer1_outputs(1363) <= a;
    layer1_outputs(1364) <= b and not a;
    layer1_outputs(1365) <= '1';
    layer1_outputs(1366) <= b and not a;
    layer1_outputs(1367) <= a;
    layer1_outputs(1368) <= a and b;
    layer1_outputs(1369) <= a and b;
    layer1_outputs(1370) <= not (a xor b);
    layer1_outputs(1371) <= '0';
    layer1_outputs(1372) <= a and not b;
    layer1_outputs(1373) <= not b or a;
    layer1_outputs(1374) <= '1';
    layer1_outputs(1375) <= b and not a;
    layer1_outputs(1376) <= not a;
    layer1_outputs(1377) <= b and not a;
    layer1_outputs(1378) <= not (a xor b);
    layer1_outputs(1379) <= not (a and b);
    layer1_outputs(1380) <= not (a and b);
    layer1_outputs(1381) <= b and not a;
    layer1_outputs(1382) <= a and b;
    layer1_outputs(1383) <= not b;
    layer1_outputs(1384) <= '1';
    layer1_outputs(1385) <= '1';
    layer1_outputs(1386) <= not b;
    layer1_outputs(1387) <= '0';
    layer1_outputs(1388) <= a and b;
    layer1_outputs(1389) <= not b;
    layer1_outputs(1390) <= '1';
    layer1_outputs(1391) <= '0';
    layer1_outputs(1392) <= not b or a;
    layer1_outputs(1393) <= a and b;
    layer1_outputs(1394) <= b and not a;
    layer1_outputs(1395) <= b;
    layer1_outputs(1396) <= a or b;
    layer1_outputs(1397) <= not (a xor b);
    layer1_outputs(1398) <= a xor b;
    layer1_outputs(1399) <= a and not b;
    layer1_outputs(1400) <= a or b;
    layer1_outputs(1401) <= not (a and b);
    layer1_outputs(1402) <= '0';
    layer1_outputs(1403) <= '1';
    layer1_outputs(1404) <= '1';
    layer1_outputs(1405) <= '0';
    layer1_outputs(1406) <= a;
    layer1_outputs(1407) <= b and not a;
    layer1_outputs(1408) <= not (a and b);
    layer1_outputs(1409) <= '0';
    layer1_outputs(1410) <= a and not b;
    layer1_outputs(1411) <= not a;
    layer1_outputs(1412) <= a and not b;
    layer1_outputs(1413) <= not a;
    layer1_outputs(1414) <= a or b;
    layer1_outputs(1415) <= a or b;
    layer1_outputs(1416) <= not b or a;
    layer1_outputs(1417) <= '1';
    layer1_outputs(1418) <= not (a or b);
    layer1_outputs(1419) <= b and not a;
    layer1_outputs(1420) <= b and not a;
    layer1_outputs(1421) <= a or b;
    layer1_outputs(1422) <= '0';
    layer1_outputs(1423) <= a;
    layer1_outputs(1424) <= a;
    layer1_outputs(1425) <= not a or b;
    layer1_outputs(1426) <= not a or b;
    layer1_outputs(1427) <= a;
    layer1_outputs(1428) <= b;
    layer1_outputs(1429) <= a xor b;
    layer1_outputs(1430) <= not b;
    layer1_outputs(1431) <= not (a xor b);
    layer1_outputs(1432) <= a xor b;
    layer1_outputs(1433) <= '0';
    layer1_outputs(1434) <= b and not a;
    layer1_outputs(1435) <= not (a xor b);
    layer1_outputs(1436) <= a and b;
    layer1_outputs(1437) <= not (a or b);
    layer1_outputs(1438) <= not b;
    layer1_outputs(1439) <= not a or b;
    layer1_outputs(1440) <= a or b;
    layer1_outputs(1441) <= a and b;
    layer1_outputs(1442) <= not (a or b);
    layer1_outputs(1443) <= not (a and b);
    layer1_outputs(1444) <= a;
    layer1_outputs(1445) <= not b;
    layer1_outputs(1446) <= a and not b;
    layer1_outputs(1447) <= not (a and b);
    layer1_outputs(1448) <= not a or b;
    layer1_outputs(1449) <= not b or a;
    layer1_outputs(1450) <= b;
    layer1_outputs(1451) <= '1';
    layer1_outputs(1452) <= a and b;
    layer1_outputs(1453) <= a or b;
    layer1_outputs(1454) <= '1';
    layer1_outputs(1455) <= not a;
    layer1_outputs(1456) <= not b;
    layer1_outputs(1457) <= not a;
    layer1_outputs(1458) <= b;
    layer1_outputs(1459) <= a and not b;
    layer1_outputs(1460) <= a or b;
    layer1_outputs(1461) <= not (a or b);
    layer1_outputs(1462) <= '1';
    layer1_outputs(1463) <= not a;
    layer1_outputs(1464) <= '1';
    layer1_outputs(1465) <= a and b;
    layer1_outputs(1466) <= not (a or b);
    layer1_outputs(1467) <= not b;
    layer1_outputs(1468) <= '0';
    layer1_outputs(1469) <= not (a and b);
    layer1_outputs(1470) <= '1';
    layer1_outputs(1471) <= '1';
    layer1_outputs(1472) <= a and b;
    layer1_outputs(1473) <= not a or b;
    layer1_outputs(1474) <= a xor b;
    layer1_outputs(1475) <= not a or b;
    layer1_outputs(1476) <= a and b;
    layer1_outputs(1477) <= not (a and b);
    layer1_outputs(1478) <= not b;
    layer1_outputs(1479) <= not (a and b);
    layer1_outputs(1480) <= not a or b;
    layer1_outputs(1481) <= not a or b;
    layer1_outputs(1482) <= '0';
    layer1_outputs(1483) <= b;
    layer1_outputs(1484) <= not (a and b);
    layer1_outputs(1485) <= not (a and b);
    layer1_outputs(1486) <= not (a and b);
    layer1_outputs(1487) <= a and not b;
    layer1_outputs(1488) <= not a or b;
    layer1_outputs(1489) <= a and not b;
    layer1_outputs(1490) <= b;
    layer1_outputs(1491) <= b and not a;
    layer1_outputs(1492) <= '1';
    layer1_outputs(1493) <= a and b;
    layer1_outputs(1494) <= b and not a;
    layer1_outputs(1495) <= '0';
    layer1_outputs(1496) <= a;
    layer1_outputs(1497) <= not b;
    layer1_outputs(1498) <= '0';
    layer1_outputs(1499) <= b;
    layer1_outputs(1500) <= a xor b;
    layer1_outputs(1501) <= a or b;
    layer1_outputs(1502) <= a and b;
    layer1_outputs(1503) <= '1';
    layer1_outputs(1504) <= not b or a;
    layer1_outputs(1505) <= not b;
    layer1_outputs(1506) <= not (a or b);
    layer1_outputs(1507) <= '0';
    layer1_outputs(1508) <= a or b;
    layer1_outputs(1509) <= not (a and b);
    layer1_outputs(1510) <= a and not b;
    layer1_outputs(1511) <= b and not a;
    layer1_outputs(1512) <= b;
    layer1_outputs(1513) <= not (a and b);
    layer1_outputs(1514) <= a and not b;
    layer1_outputs(1515) <= b and not a;
    layer1_outputs(1516) <= not b;
    layer1_outputs(1517) <= a and b;
    layer1_outputs(1518) <= not (a and b);
    layer1_outputs(1519) <= a and not b;
    layer1_outputs(1520) <= '0';
    layer1_outputs(1521) <= not a or b;
    layer1_outputs(1522) <= not b;
    layer1_outputs(1523) <= not (a and b);
    layer1_outputs(1524) <= '0';
    layer1_outputs(1525) <= not b;
    layer1_outputs(1526) <= a or b;
    layer1_outputs(1527) <= '1';
    layer1_outputs(1528) <= not (a or b);
    layer1_outputs(1529) <= not b or a;
    layer1_outputs(1530) <= not (a or b);
    layer1_outputs(1531) <= b and not a;
    layer1_outputs(1532) <= '0';
    layer1_outputs(1533) <= not b or a;
    layer1_outputs(1534) <= not (a and b);
    layer1_outputs(1535) <= b and not a;
    layer1_outputs(1536) <= not b;
    layer1_outputs(1537) <= a;
    layer1_outputs(1538) <= not a or b;
    layer1_outputs(1539) <= not (a and b);
    layer1_outputs(1540) <= not a;
    layer1_outputs(1541) <= not (a xor b);
    layer1_outputs(1542) <= not (a and b);
    layer1_outputs(1543) <= a or b;
    layer1_outputs(1544) <= a and b;
    layer1_outputs(1545) <= not a;
    layer1_outputs(1546) <= not (a xor b);
    layer1_outputs(1547) <= b;
    layer1_outputs(1548) <= b and not a;
    layer1_outputs(1549) <= not b;
    layer1_outputs(1550) <= '0';
    layer1_outputs(1551) <= not a or b;
    layer1_outputs(1552) <= not b;
    layer1_outputs(1553) <= a and b;
    layer1_outputs(1554) <= not (a and b);
    layer1_outputs(1555) <= not (a or b);
    layer1_outputs(1556) <= a and not b;
    layer1_outputs(1557) <= not a or b;
    layer1_outputs(1558) <= '0';
    layer1_outputs(1559) <= not (a and b);
    layer1_outputs(1560) <= not (a or b);
    layer1_outputs(1561) <= b and not a;
    layer1_outputs(1562) <= a and not b;
    layer1_outputs(1563) <= a and not b;
    layer1_outputs(1564) <= b;
    layer1_outputs(1565) <= a;
    layer1_outputs(1566) <= not b or a;
    layer1_outputs(1567) <= a and not b;
    layer1_outputs(1568) <= '1';
    layer1_outputs(1569) <= b;
    layer1_outputs(1570) <= not (a xor b);
    layer1_outputs(1571) <= not b or a;
    layer1_outputs(1572) <= not b;
    layer1_outputs(1573) <= a and not b;
    layer1_outputs(1574) <= b and not a;
    layer1_outputs(1575) <= not b;
    layer1_outputs(1576) <= '0';
    layer1_outputs(1577) <= not b or a;
    layer1_outputs(1578) <= '0';
    layer1_outputs(1579) <= '1';
    layer1_outputs(1580) <= not a or b;
    layer1_outputs(1581) <= a and not b;
    layer1_outputs(1582) <= a or b;
    layer1_outputs(1583) <= b;
    layer1_outputs(1584) <= not b or a;
    layer1_outputs(1585) <= not b or a;
    layer1_outputs(1586) <= b and not a;
    layer1_outputs(1587) <= not (a or b);
    layer1_outputs(1588) <= not (a and b);
    layer1_outputs(1589) <= a or b;
    layer1_outputs(1590) <= '0';
    layer1_outputs(1591) <= '1';
    layer1_outputs(1592) <= '0';
    layer1_outputs(1593) <= not a or b;
    layer1_outputs(1594) <= not (a xor b);
    layer1_outputs(1595) <= '0';
    layer1_outputs(1596) <= not a or b;
    layer1_outputs(1597) <= '1';
    layer1_outputs(1598) <= a and not b;
    layer1_outputs(1599) <= not a;
    layer1_outputs(1600) <= not a or b;
    layer1_outputs(1601) <= not b;
    layer1_outputs(1602) <= '1';
    layer1_outputs(1603) <= not (a and b);
    layer1_outputs(1604) <= not b;
    layer1_outputs(1605) <= not b or a;
    layer1_outputs(1606) <= a and b;
    layer1_outputs(1607) <= '1';
    layer1_outputs(1608) <= b;
    layer1_outputs(1609) <= b;
    layer1_outputs(1610) <= a;
    layer1_outputs(1611) <= not b;
    layer1_outputs(1612) <= not (a and b);
    layer1_outputs(1613) <= '0';
    layer1_outputs(1614) <= not (a and b);
    layer1_outputs(1615) <= '1';
    layer1_outputs(1616) <= not a or b;
    layer1_outputs(1617) <= a;
    layer1_outputs(1618) <= a;
    layer1_outputs(1619) <= b and not a;
    layer1_outputs(1620) <= a;
    layer1_outputs(1621) <= a xor b;
    layer1_outputs(1622) <= not (a or b);
    layer1_outputs(1623) <= '1';
    layer1_outputs(1624) <= a;
    layer1_outputs(1625) <= '1';
    layer1_outputs(1626) <= not a or b;
    layer1_outputs(1627) <= a and not b;
    layer1_outputs(1628) <= a and not b;
    layer1_outputs(1629) <= '1';
    layer1_outputs(1630) <= a and not b;
    layer1_outputs(1631) <= not b or a;
    layer1_outputs(1632) <= not (a and b);
    layer1_outputs(1633) <= b and not a;
    layer1_outputs(1634) <= b;
    layer1_outputs(1635) <= b and not a;
    layer1_outputs(1636) <= a and not b;
    layer1_outputs(1637) <= b and not a;
    layer1_outputs(1638) <= a xor b;
    layer1_outputs(1639) <= '0';
    layer1_outputs(1640) <= '0';
    layer1_outputs(1641) <= '1';
    layer1_outputs(1642) <= '1';
    layer1_outputs(1643) <= a or b;
    layer1_outputs(1644) <= not b or a;
    layer1_outputs(1645) <= not a;
    layer1_outputs(1646) <= not b or a;
    layer1_outputs(1647) <= not (a or b);
    layer1_outputs(1648) <= '0';
    layer1_outputs(1649) <= not a or b;
    layer1_outputs(1650) <= not a or b;
    layer1_outputs(1651) <= '0';
    layer1_outputs(1652) <= not b;
    layer1_outputs(1653) <= a or b;
    layer1_outputs(1654) <= not b;
    layer1_outputs(1655) <= a xor b;
    layer1_outputs(1656) <= b;
    layer1_outputs(1657) <= '0';
    layer1_outputs(1658) <= a;
    layer1_outputs(1659) <= not a;
    layer1_outputs(1660) <= not b or a;
    layer1_outputs(1661) <= not a;
    layer1_outputs(1662) <= a and not b;
    layer1_outputs(1663) <= not b;
    layer1_outputs(1664) <= a or b;
    layer1_outputs(1665) <= a and b;
    layer1_outputs(1666) <= b and not a;
    layer1_outputs(1667) <= '1';
    layer1_outputs(1668) <= not a;
    layer1_outputs(1669) <= b;
    layer1_outputs(1670) <= b and not a;
    layer1_outputs(1671) <= not (a and b);
    layer1_outputs(1672) <= b;
    layer1_outputs(1673) <= b;
    layer1_outputs(1674) <= a and b;
    layer1_outputs(1675) <= not a or b;
    layer1_outputs(1676) <= '1';
    layer1_outputs(1677) <= b;
    layer1_outputs(1678) <= '1';
    layer1_outputs(1679) <= not a;
    layer1_outputs(1680) <= b and not a;
    layer1_outputs(1681) <= b;
    layer1_outputs(1682) <= a and not b;
    layer1_outputs(1683) <= b;
    layer1_outputs(1684) <= '1';
    layer1_outputs(1685) <= a and b;
    layer1_outputs(1686) <= a and b;
    layer1_outputs(1687) <= not b;
    layer1_outputs(1688) <= not a or b;
    layer1_outputs(1689) <= a;
    layer1_outputs(1690) <= '0';
    layer1_outputs(1691) <= not b or a;
    layer1_outputs(1692) <= b and not a;
    layer1_outputs(1693) <= a and not b;
    layer1_outputs(1694) <= not a or b;
    layer1_outputs(1695) <= a and b;
    layer1_outputs(1696) <= not (a and b);
    layer1_outputs(1697) <= a and b;
    layer1_outputs(1698) <= a and not b;
    layer1_outputs(1699) <= a xor b;
    layer1_outputs(1700) <= a and not b;
    layer1_outputs(1701) <= '0';
    layer1_outputs(1702) <= '0';
    layer1_outputs(1703) <= a or b;
    layer1_outputs(1704) <= not b or a;
    layer1_outputs(1705) <= not b;
    layer1_outputs(1706) <= b;
    layer1_outputs(1707) <= a or b;
    layer1_outputs(1708) <= a xor b;
    layer1_outputs(1709) <= not a;
    layer1_outputs(1710) <= b and not a;
    layer1_outputs(1711) <= not (a or b);
    layer1_outputs(1712) <= a;
    layer1_outputs(1713) <= not (a or b);
    layer1_outputs(1714) <= b and not a;
    layer1_outputs(1715) <= not a;
    layer1_outputs(1716) <= not (a or b);
    layer1_outputs(1717) <= not (a and b);
    layer1_outputs(1718) <= not (a or b);
    layer1_outputs(1719) <= a and b;
    layer1_outputs(1720) <= not b;
    layer1_outputs(1721) <= a;
    layer1_outputs(1722) <= a and not b;
    layer1_outputs(1723) <= not b or a;
    layer1_outputs(1724) <= '1';
    layer1_outputs(1725) <= a and b;
    layer1_outputs(1726) <= not b or a;
    layer1_outputs(1727) <= a;
    layer1_outputs(1728) <= a or b;
    layer1_outputs(1729) <= not (a and b);
    layer1_outputs(1730) <= a and not b;
    layer1_outputs(1731) <= '1';
    layer1_outputs(1732) <= '0';
    layer1_outputs(1733) <= not (a xor b);
    layer1_outputs(1734) <= '1';
    layer1_outputs(1735) <= not b or a;
    layer1_outputs(1736) <= a or b;
    layer1_outputs(1737) <= a and not b;
    layer1_outputs(1738) <= '1';
    layer1_outputs(1739) <= a and b;
    layer1_outputs(1740) <= not (a or b);
    layer1_outputs(1741) <= not (a or b);
    layer1_outputs(1742) <= a or b;
    layer1_outputs(1743) <= b;
    layer1_outputs(1744) <= a;
    layer1_outputs(1745) <= not a or b;
    layer1_outputs(1746) <= '1';
    layer1_outputs(1747) <= '1';
    layer1_outputs(1748) <= '0';
    layer1_outputs(1749) <= not (a and b);
    layer1_outputs(1750) <= b;
    layer1_outputs(1751) <= not (a or b);
    layer1_outputs(1752) <= not a;
    layer1_outputs(1753) <= '1';
    layer1_outputs(1754) <= a and not b;
    layer1_outputs(1755) <= a and b;
    layer1_outputs(1756) <= a or b;
    layer1_outputs(1757) <= '1';
    layer1_outputs(1758) <= not b;
    layer1_outputs(1759) <= '1';
    layer1_outputs(1760) <= a and b;
    layer1_outputs(1761) <= not a;
    layer1_outputs(1762) <= '0';
    layer1_outputs(1763) <= '0';
    layer1_outputs(1764) <= a and b;
    layer1_outputs(1765) <= not (a or b);
    layer1_outputs(1766) <= a;
    layer1_outputs(1767) <= '0';
    layer1_outputs(1768) <= a;
    layer1_outputs(1769) <= not b or a;
    layer1_outputs(1770) <= a xor b;
    layer1_outputs(1771) <= not (a and b);
    layer1_outputs(1772) <= not b;
    layer1_outputs(1773) <= a and not b;
    layer1_outputs(1774) <= a or b;
    layer1_outputs(1775) <= '1';
    layer1_outputs(1776) <= not a;
    layer1_outputs(1777) <= b;
    layer1_outputs(1778) <= '0';
    layer1_outputs(1779) <= b and not a;
    layer1_outputs(1780) <= not b or a;
    layer1_outputs(1781) <= not b or a;
    layer1_outputs(1782) <= a;
    layer1_outputs(1783) <= '0';
    layer1_outputs(1784) <= not a;
    layer1_outputs(1785) <= not a;
    layer1_outputs(1786) <= not a;
    layer1_outputs(1787) <= '1';
    layer1_outputs(1788) <= b and not a;
    layer1_outputs(1789) <= not (a or b);
    layer1_outputs(1790) <= not (a and b);
    layer1_outputs(1791) <= a or b;
    layer1_outputs(1792) <= a;
    layer1_outputs(1793) <= a;
    layer1_outputs(1794) <= not a or b;
    layer1_outputs(1795) <= not b or a;
    layer1_outputs(1796) <= not a or b;
    layer1_outputs(1797) <= not a;
    layer1_outputs(1798) <= a or b;
    layer1_outputs(1799) <= not b;
    layer1_outputs(1800) <= '0';
    layer1_outputs(1801) <= not b;
    layer1_outputs(1802) <= a and not b;
    layer1_outputs(1803) <= '0';
    layer1_outputs(1804) <= a;
    layer1_outputs(1805) <= not b or a;
    layer1_outputs(1806) <= not (a and b);
    layer1_outputs(1807) <= a xor b;
    layer1_outputs(1808) <= not b;
    layer1_outputs(1809) <= a xor b;
    layer1_outputs(1810) <= not (a and b);
    layer1_outputs(1811) <= not a;
    layer1_outputs(1812) <= not b or a;
    layer1_outputs(1813) <= b and not a;
    layer1_outputs(1814) <= a and b;
    layer1_outputs(1815) <= not (a or b);
    layer1_outputs(1816) <= b;
    layer1_outputs(1817) <= a and not b;
    layer1_outputs(1818) <= '0';
    layer1_outputs(1819) <= not b or a;
    layer1_outputs(1820) <= a and not b;
    layer1_outputs(1821) <= '1';
    layer1_outputs(1822) <= a and not b;
    layer1_outputs(1823) <= not a or b;
    layer1_outputs(1824) <= '0';
    layer1_outputs(1825) <= not b;
    layer1_outputs(1826) <= a and b;
    layer1_outputs(1827) <= a;
    layer1_outputs(1828) <= not (a or b);
    layer1_outputs(1829) <= not b or a;
    layer1_outputs(1830) <= not (a and b);
    layer1_outputs(1831) <= a;
    layer1_outputs(1832) <= a or b;
    layer1_outputs(1833) <= not a;
    layer1_outputs(1834) <= not b;
    layer1_outputs(1835) <= '1';
    layer1_outputs(1836) <= not b;
    layer1_outputs(1837) <= '0';
    layer1_outputs(1838) <= not a;
    layer1_outputs(1839) <= not a or b;
    layer1_outputs(1840) <= '0';
    layer1_outputs(1841) <= not b or a;
    layer1_outputs(1842) <= not b;
    layer1_outputs(1843) <= a;
    layer1_outputs(1844) <= not (a or b);
    layer1_outputs(1845) <= not a;
    layer1_outputs(1846) <= b;
    layer1_outputs(1847) <= not a or b;
    layer1_outputs(1848) <= not a or b;
    layer1_outputs(1849) <= a or b;
    layer1_outputs(1850) <= not a or b;
    layer1_outputs(1851) <= '1';
    layer1_outputs(1852) <= '1';
    layer1_outputs(1853) <= a or b;
    layer1_outputs(1854) <= not b or a;
    layer1_outputs(1855) <= not a;
    layer1_outputs(1856) <= a and b;
    layer1_outputs(1857) <= not b;
    layer1_outputs(1858) <= a and b;
    layer1_outputs(1859) <= '1';
    layer1_outputs(1860) <= b;
    layer1_outputs(1861) <= not a or b;
    layer1_outputs(1862) <= a and not b;
    layer1_outputs(1863) <= not (a or b);
    layer1_outputs(1864) <= a and not b;
    layer1_outputs(1865) <= not a;
    layer1_outputs(1866) <= not (a or b);
    layer1_outputs(1867) <= not a;
    layer1_outputs(1868) <= not a or b;
    layer1_outputs(1869) <= a and not b;
    layer1_outputs(1870) <= b and not a;
    layer1_outputs(1871) <= not (a or b);
    layer1_outputs(1872) <= a and not b;
    layer1_outputs(1873) <= b and not a;
    layer1_outputs(1874) <= '1';
    layer1_outputs(1875) <= not b or a;
    layer1_outputs(1876) <= not a or b;
    layer1_outputs(1877) <= not (a or b);
    layer1_outputs(1878) <= '0';
    layer1_outputs(1879) <= b and not a;
    layer1_outputs(1880) <= a and b;
    layer1_outputs(1881) <= not (a or b);
    layer1_outputs(1882) <= a or b;
    layer1_outputs(1883) <= a and not b;
    layer1_outputs(1884) <= not (a or b);
    layer1_outputs(1885) <= not b;
    layer1_outputs(1886) <= not a;
    layer1_outputs(1887) <= not b or a;
    layer1_outputs(1888) <= b;
    layer1_outputs(1889) <= '0';
    layer1_outputs(1890) <= a and b;
    layer1_outputs(1891) <= not b;
    layer1_outputs(1892) <= '0';
    layer1_outputs(1893) <= not b or a;
    layer1_outputs(1894) <= not b;
    layer1_outputs(1895) <= a and not b;
    layer1_outputs(1896) <= not b or a;
    layer1_outputs(1897) <= a;
    layer1_outputs(1898) <= not a;
    layer1_outputs(1899) <= not a;
    layer1_outputs(1900) <= a or b;
    layer1_outputs(1901) <= '0';
    layer1_outputs(1902) <= not b or a;
    layer1_outputs(1903) <= '0';
    layer1_outputs(1904) <= b and not a;
    layer1_outputs(1905) <= b and not a;
    layer1_outputs(1906) <= a;
    layer1_outputs(1907) <= a and not b;
    layer1_outputs(1908) <= a and b;
    layer1_outputs(1909) <= not a or b;
    layer1_outputs(1910) <= a and not b;
    layer1_outputs(1911) <= '1';
    layer1_outputs(1912) <= '1';
    layer1_outputs(1913) <= not b;
    layer1_outputs(1914) <= not a;
    layer1_outputs(1915) <= a and b;
    layer1_outputs(1916) <= '1';
    layer1_outputs(1917) <= not b or a;
    layer1_outputs(1918) <= not (a or b);
    layer1_outputs(1919) <= not (a and b);
    layer1_outputs(1920) <= not (a and b);
    layer1_outputs(1921) <= not (a and b);
    layer1_outputs(1922) <= not a;
    layer1_outputs(1923) <= not b;
    layer1_outputs(1924) <= not b;
    layer1_outputs(1925) <= '0';
    layer1_outputs(1926) <= not (a or b);
    layer1_outputs(1927) <= a;
    layer1_outputs(1928) <= a and not b;
    layer1_outputs(1929) <= not (a or b);
    layer1_outputs(1930) <= not (a or b);
    layer1_outputs(1931) <= b;
    layer1_outputs(1932) <= '1';
    layer1_outputs(1933) <= not a or b;
    layer1_outputs(1934) <= not a;
    layer1_outputs(1935) <= '0';
    layer1_outputs(1936) <= '1';
    layer1_outputs(1937) <= '0';
    layer1_outputs(1938) <= not a or b;
    layer1_outputs(1939) <= '0';
    layer1_outputs(1940) <= not b;
    layer1_outputs(1941) <= not b or a;
    layer1_outputs(1942) <= not b or a;
    layer1_outputs(1943) <= a and not b;
    layer1_outputs(1944) <= a and b;
    layer1_outputs(1945) <= a or b;
    layer1_outputs(1946) <= a;
    layer1_outputs(1947) <= not b or a;
    layer1_outputs(1948) <= '1';
    layer1_outputs(1949) <= a and not b;
    layer1_outputs(1950) <= a;
    layer1_outputs(1951) <= not a or b;
    layer1_outputs(1952) <= not b or a;
    layer1_outputs(1953) <= b;
    layer1_outputs(1954) <= b;
    layer1_outputs(1955) <= not (a and b);
    layer1_outputs(1956) <= a or b;
    layer1_outputs(1957) <= '1';
    layer1_outputs(1958) <= not b;
    layer1_outputs(1959) <= '0';
    layer1_outputs(1960) <= not a;
    layer1_outputs(1961) <= '1';
    layer1_outputs(1962) <= b and not a;
    layer1_outputs(1963) <= a or b;
    layer1_outputs(1964) <= '0';
    layer1_outputs(1965) <= not (a and b);
    layer1_outputs(1966) <= a and b;
    layer1_outputs(1967) <= a and not b;
    layer1_outputs(1968) <= not (a xor b);
    layer1_outputs(1969) <= not b;
    layer1_outputs(1970) <= '1';
    layer1_outputs(1971) <= a xor b;
    layer1_outputs(1972) <= not a or b;
    layer1_outputs(1973) <= '1';
    layer1_outputs(1974) <= b and not a;
    layer1_outputs(1975) <= a xor b;
    layer1_outputs(1976) <= '0';
    layer1_outputs(1977) <= a;
    layer1_outputs(1978) <= '1';
    layer1_outputs(1979) <= a or b;
    layer1_outputs(1980) <= not b;
    layer1_outputs(1981) <= a or b;
    layer1_outputs(1982) <= a and not b;
    layer1_outputs(1983) <= b and not a;
    layer1_outputs(1984) <= not b or a;
    layer1_outputs(1985) <= a and b;
    layer1_outputs(1986) <= not (a or b);
    layer1_outputs(1987) <= '1';
    layer1_outputs(1988) <= a or b;
    layer1_outputs(1989) <= b;
    layer1_outputs(1990) <= '0';
    layer1_outputs(1991) <= a;
    layer1_outputs(1992) <= not a or b;
    layer1_outputs(1993) <= a and b;
    layer1_outputs(1994) <= a;
    layer1_outputs(1995) <= not b or a;
    layer1_outputs(1996) <= not b or a;
    layer1_outputs(1997) <= not (a or b);
    layer1_outputs(1998) <= b and not a;
    layer1_outputs(1999) <= a xor b;
    layer1_outputs(2000) <= a xor b;
    layer1_outputs(2001) <= a and b;
    layer1_outputs(2002) <= b and not a;
    layer1_outputs(2003) <= not (a and b);
    layer1_outputs(2004) <= '1';
    layer1_outputs(2005) <= a;
    layer1_outputs(2006) <= '0';
    layer1_outputs(2007) <= not (a and b);
    layer1_outputs(2008) <= not b or a;
    layer1_outputs(2009) <= not (a and b);
    layer1_outputs(2010) <= not b or a;
    layer1_outputs(2011) <= '1';
    layer1_outputs(2012) <= not b or a;
    layer1_outputs(2013) <= b;
    layer1_outputs(2014) <= a or b;
    layer1_outputs(2015) <= a and not b;
    layer1_outputs(2016) <= not a or b;
    layer1_outputs(2017) <= a or b;
    layer1_outputs(2018) <= '1';
    layer1_outputs(2019) <= not (a and b);
    layer1_outputs(2020) <= not b or a;
    layer1_outputs(2021) <= b and not a;
    layer1_outputs(2022) <= a xor b;
    layer1_outputs(2023) <= a;
    layer1_outputs(2024) <= '1';
    layer1_outputs(2025) <= not a;
    layer1_outputs(2026) <= a and b;
    layer1_outputs(2027) <= not a or b;
    layer1_outputs(2028) <= not (a and b);
    layer1_outputs(2029) <= b;
    layer1_outputs(2030) <= a and b;
    layer1_outputs(2031) <= a xor b;
    layer1_outputs(2032) <= not b;
    layer1_outputs(2033) <= a or b;
    layer1_outputs(2034) <= a xor b;
    layer1_outputs(2035) <= '0';
    layer1_outputs(2036) <= not (a and b);
    layer1_outputs(2037) <= not (a and b);
    layer1_outputs(2038) <= '1';
    layer1_outputs(2039) <= not (a and b);
    layer1_outputs(2040) <= a xor b;
    layer1_outputs(2041) <= '0';
    layer1_outputs(2042) <= a and not b;
    layer1_outputs(2043) <= '0';
    layer1_outputs(2044) <= a and not b;
    layer1_outputs(2045) <= not b or a;
    layer1_outputs(2046) <= '1';
    layer1_outputs(2047) <= not (a xor b);
    layer1_outputs(2048) <= not (a and b);
    layer1_outputs(2049) <= not (a and b);
    layer1_outputs(2050) <= not b;
    layer1_outputs(2051) <= '1';
    layer1_outputs(2052) <= a and b;
    layer1_outputs(2053) <= '0';
    layer1_outputs(2054) <= a or b;
    layer1_outputs(2055) <= b;
    layer1_outputs(2056) <= not (a xor b);
    layer1_outputs(2057) <= '1';
    layer1_outputs(2058) <= b;
    layer1_outputs(2059) <= a and not b;
    layer1_outputs(2060) <= b;
    layer1_outputs(2061) <= not a or b;
    layer1_outputs(2062) <= a and b;
    layer1_outputs(2063) <= a and not b;
    layer1_outputs(2064) <= '1';
    layer1_outputs(2065) <= '0';
    layer1_outputs(2066) <= a and not b;
    layer1_outputs(2067) <= not b or a;
    layer1_outputs(2068) <= a and not b;
    layer1_outputs(2069) <= b and not a;
    layer1_outputs(2070) <= a and b;
    layer1_outputs(2071) <= a and not b;
    layer1_outputs(2072) <= not (a and b);
    layer1_outputs(2073) <= not (a and b);
    layer1_outputs(2074) <= not (a or b);
    layer1_outputs(2075) <= a;
    layer1_outputs(2076) <= '1';
    layer1_outputs(2077) <= not (a or b);
    layer1_outputs(2078) <= b and not a;
    layer1_outputs(2079) <= not b or a;
    layer1_outputs(2080) <= not a;
    layer1_outputs(2081) <= a or b;
    layer1_outputs(2082) <= '1';
    layer1_outputs(2083) <= '1';
    layer1_outputs(2084) <= '0';
    layer1_outputs(2085) <= '0';
    layer1_outputs(2086) <= not b or a;
    layer1_outputs(2087) <= a and b;
    layer1_outputs(2088) <= not (a or b);
    layer1_outputs(2089) <= not b or a;
    layer1_outputs(2090) <= not a or b;
    layer1_outputs(2091) <= not a;
    layer1_outputs(2092) <= '1';
    layer1_outputs(2093) <= a and b;
    layer1_outputs(2094) <= a and b;
    layer1_outputs(2095) <= b and not a;
    layer1_outputs(2096) <= a or b;
    layer1_outputs(2097) <= not (a and b);
    layer1_outputs(2098) <= a and b;
    layer1_outputs(2099) <= not b or a;
    layer1_outputs(2100) <= not b or a;
    layer1_outputs(2101) <= not b;
    layer1_outputs(2102) <= not (a or b);
    layer1_outputs(2103) <= not a or b;
    layer1_outputs(2104) <= '0';
    layer1_outputs(2105) <= '0';
    layer1_outputs(2106) <= b;
    layer1_outputs(2107) <= not (a xor b);
    layer1_outputs(2108) <= a or b;
    layer1_outputs(2109) <= not (a and b);
    layer1_outputs(2110) <= not b or a;
    layer1_outputs(2111) <= b and not a;
    layer1_outputs(2112) <= '0';
    layer1_outputs(2113) <= not b or a;
    layer1_outputs(2114) <= '0';
    layer1_outputs(2115) <= '0';
    layer1_outputs(2116) <= b and not a;
    layer1_outputs(2117) <= a and not b;
    layer1_outputs(2118) <= not (a or b);
    layer1_outputs(2119) <= not a;
    layer1_outputs(2120) <= a;
    layer1_outputs(2121) <= b and not a;
    layer1_outputs(2122) <= b;
    layer1_outputs(2123) <= '1';
    layer1_outputs(2124) <= not (a and b);
    layer1_outputs(2125) <= not (a or b);
    layer1_outputs(2126) <= not a or b;
    layer1_outputs(2127) <= not (a or b);
    layer1_outputs(2128) <= a;
    layer1_outputs(2129) <= '0';
    layer1_outputs(2130) <= not (a and b);
    layer1_outputs(2131) <= b;
    layer1_outputs(2132) <= not (a xor b);
    layer1_outputs(2133) <= a and b;
    layer1_outputs(2134) <= b;
    layer1_outputs(2135) <= '0';
    layer1_outputs(2136) <= a and not b;
    layer1_outputs(2137) <= not b or a;
    layer1_outputs(2138) <= a and not b;
    layer1_outputs(2139) <= not b or a;
    layer1_outputs(2140) <= '1';
    layer1_outputs(2141) <= not b or a;
    layer1_outputs(2142) <= not a or b;
    layer1_outputs(2143) <= '0';
    layer1_outputs(2144) <= not b;
    layer1_outputs(2145) <= not b;
    layer1_outputs(2146) <= a and not b;
    layer1_outputs(2147) <= not b or a;
    layer1_outputs(2148) <= not a or b;
    layer1_outputs(2149) <= not (a or b);
    layer1_outputs(2150) <= not a or b;
    layer1_outputs(2151) <= not (a xor b);
    layer1_outputs(2152) <= not (a xor b);
    layer1_outputs(2153) <= not (a or b);
    layer1_outputs(2154) <= not a;
    layer1_outputs(2155) <= a;
    layer1_outputs(2156) <= not (a and b);
    layer1_outputs(2157) <= a or b;
    layer1_outputs(2158) <= not a;
    layer1_outputs(2159) <= a;
    layer1_outputs(2160) <= not a;
    layer1_outputs(2161) <= not (a and b);
    layer1_outputs(2162) <= not a or b;
    layer1_outputs(2163) <= '0';
    layer1_outputs(2164) <= b;
    layer1_outputs(2165) <= b;
    layer1_outputs(2166) <= '1';
    layer1_outputs(2167) <= not (a and b);
    layer1_outputs(2168) <= not (a and b);
    layer1_outputs(2169) <= a and b;
    layer1_outputs(2170) <= '1';
    layer1_outputs(2171) <= not (a xor b);
    layer1_outputs(2172) <= '0';
    layer1_outputs(2173) <= b and not a;
    layer1_outputs(2174) <= b;
    layer1_outputs(2175) <= a or b;
    layer1_outputs(2176) <= a;
    layer1_outputs(2177) <= b;
    layer1_outputs(2178) <= a and b;
    layer1_outputs(2179) <= not (a xor b);
    layer1_outputs(2180) <= a or b;
    layer1_outputs(2181) <= not b;
    layer1_outputs(2182) <= a and b;
    layer1_outputs(2183) <= b and not a;
    layer1_outputs(2184) <= not b;
    layer1_outputs(2185) <= not a;
    layer1_outputs(2186) <= b;
    layer1_outputs(2187) <= not b;
    layer1_outputs(2188) <= not (a and b);
    layer1_outputs(2189) <= not a;
    layer1_outputs(2190) <= b and not a;
    layer1_outputs(2191) <= not a or b;
    layer1_outputs(2192) <= not b or a;
    layer1_outputs(2193) <= not b or a;
    layer1_outputs(2194) <= a and b;
    layer1_outputs(2195) <= b;
    layer1_outputs(2196) <= b and not a;
    layer1_outputs(2197) <= b;
    layer1_outputs(2198) <= not a;
    layer1_outputs(2199) <= not (a xor b);
    layer1_outputs(2200) <= not (a or b);
    layer1_outputs(2201) <= '0';
    layer1_outputs(2202) <= '1';
    layer1_outputs(2203) <= b and not a;
    layer1_outputs(2204) <= b and not a;
    layer1_outputs(2205) <= '1';
    layer1_outputs(2206) <= '0';
    layer1_outputs(2207) <= a and b;
    layer1_outputs(2208) <= a;
    layer1_outputs(2209) <= a;
    layer1_outputs(2210) <= not (a and b);
    layer1_outputs(2211) <= not b or a;
    layer1_outputs(2212) <= not b;
    layer1_outputs(2213) <= a;
    layer1_outputs(2214) <= b;
    layer1_outputs(2215) <= not a or b;
    layer1_outputs(2216) <= not (a or b);
    layer1_outputs(2217) <= '1';
    layer1_outputs(2218) <= '0';
    layer1_outputs(2219) <= '0';
    layer1_outputs(2220) <= a and b;
    layer1_outputs(2221) <= '1';
    layer1_outputs(2222) <= '0';
    layer1_outputs(2223) <= not (a and b);
    layer1_outputs(2224) <= not b;
    layer1_outputs(2225) <= '1';
    layer1_outputs(2226) <= b and not a;
    layer1_outputs(2227) <= '0';
    layer1_outputs(2228) <= '0';
    layer1_outputs(2229) <= not (a or b);
    layer1_outputs(2230) <= '0';
    layer1_outputs(2231) <= not (a and b);
    layer1_outputs(2232) <= not (a and b);
    layer1_outputs(2233) <= b and not a;
    layer1_outputs(2234) <= b and not a;
    layer1_outputs(2235) <= not b;
    layer1_outputs(2236) <= a or b;
    layer1_outputs(2237) <= not b or a;
    layer1_outputs(2238) <= '0';
    layer1_outputs(2239) <= not b or a;
    layer1_outputs(2240) <= not (a and b);
    layer1_outputs(2241) <= not (a and b);
    layer1_outputs(2242) <= '1';
    layer1_outputs(2243) <= a and b;
    layer1_outputs(2244) <= not (a or b);
    layer1_outputs(2245) <= not (a and b);
    layer1_outputs(2246) <= b;
    layer1_outputs(2247) <= '1';
    layer1_outputs(2248) <= a;
    layer1_outputs(2249) <= a;
    layer1_outputs(2250) <= not b;
    layer1_outputs(2251) <= '1';
    layer1_outputs(2252) <= a and not b;
    layer1_outputs(2253) <= a and b;
    layer1_outputs(2254) <= not (a xor b);
    layer1_outputs(2255) <= '1';
    layer1_outputs(2256) <= a and not b;
    layer1_outputs(2257) <= '1';
    layer1_outputs(2258) <= not b or a;
    layer1_outputs(2259) <= b and not a;
    layer1_outputs(2260) <= not (a and b);
    layer1_outputs(2261) <= a xor b;
    layer1_outputs(2262) <= not (a and b);
    layer1_outputs(2263) <= '0';
    layer1_outputs(2264) <= not b;
    layer1_outputs(2265) <= a or b;
    layer1_outputs(2266) <= a and b;
    layer1_outputs(2267) <= not a;
    layer1_outputs(2268) <= not (a xor b);
    layer1_outputs(2269) <= '1';
    layer1_outputs(2270) <= '1';
    layer1_outputs(2271) <= not a or b;
    layer1_outputs(2272) <= b;
    layer1_outputs(2273) <= not (a or b);
    layer1_outputs(2274) <= not b or a;
    layer1_outputs(2275) <= b and not a;
    layer1_outputs(2276) <= not b or a;
    layer1_outputs(2277) <= '0';
    layer1_outputs(2278) <= b and not a;
    layer1_outputs(2279) <= a or b;
    layer1_outputs(2280) <= not a;
    layer1_outputs(2281) <= b and not a;
    layer1_outputs(2282) <= not a;
    layer1_outputs(2283) <= a xor b;
    layer1_outputs(2284) <= not (a or b);
    layer1_outputs(2285) <= '0';
    layer1_outputs(2286) <= b;
    layer1_outputs(2287) <= b;
    layer1_outputs(2288) <= not b;
    layer1_outputs(2289) <= b;
    layer1_outputs(2290) <= a;
    layer1_outputs(2291) <= '1';
    layer1_outputs(2292) <= not b or a;
    layer1_outputs(2293) <= not a or b;
    layer1_outputs(2294) <= not (a and b);
    layer1_outputs(2295) <= a;
    layer1_outputs(2296) <= not b or a;
    layer1_outputs(2297) <= a and b;
    layer1_outputs(2298) <= not (a and b);
    layer1_outputs(2299) <= a and b;
    layer1_outputs(2300) <= a or b;
    layer1_outputs(2301) <= not (a and b);
    layer1_outputs(2302) <= b and not a;
    layer1_outputs(2303) <= '1';
    layer1_outputs(2304) <= b;
    layer1_outputs(2305) <= a;
    layer1_outputs(2306) <= b and not a;
    layer1_outputs(2307) <= a and not b;
    layer1_outputs(2308) <= b and not a;
    layer1_outputs(2309) <= b and not a;
    layer1_outputs(2310) <= not (a and b);
    layer1_outputs(2311) <= not b;
    layer1_outputs(2312) <= a;
    layer1_outputs(2313) <= a and b;
    layer1_outputs(2314) <= not a;
    layer1_outputs(2315) <= not b;
    layer1_outputs(2316) <= not (a or b);
    layer1_outputs(2317) <= not a or b;
    layer1_outputs(2318) <= not a or b;
    layer1_outputs(2319) <= not b or a;
    layer1_outputs(2320) <= not (a and b);
    layer1_outputs(2321) <= a and b;
    layer1_outputs(2322) <= not b;
    layer1_outputs(2323) <= b and not a;
    layer1_outputs(2324) <= not a or b;
    layer1_outputs(2325) <= not (a and b);
    layer1_outputs(2326) <= not (a or b);
    layer1_outputs(2327) <= b;
    layer1_outputs(2328) <= a and not b;
    layer1_outputs(2329) <= a and b;
    layer1_outputs(2330) <= not (a xor b);
    layer1_outputs(2331) <= not b or a;
    layer1_outputs(2332) <= b;
    layer1_outputs(2333) <= b and not a;
    layer1_outputs(2334) <= b and not a;
    layer1_outputs(2335) <= not (a or b);
    layer1_outputs(2336) <= not a or b;
    layer1_outputs(2337) <= not a;
    layer1_outputs(2338) <= not (a or b);
    layer1_outputs(2339) <= not b or a;
    layer1_outputs(2340) <= a or b;
    layer1_outputs(2341) <= '0';
    layer1_outputs(2342) <= '1';
    layer1_outputs(2343) <= '0';
    layer1_outputs(2344) <= b;
    layer1_outputs(2345) <= a;
    layer1_outputs(2346) <= a xor b;
    layer1_outputs(2347) <= a or b;
    layer1_outputs(2348) <= a and not b;
    layer1_outputs(2349) <= a and b;
    layer1_outputs(2350) <= not b;
    layer1_outputs(2351) <= not b or a;
    layer1_outputs(2352) <= '0';
    layer1_outputs(2353) <= a and b;
    layer1_outputs(2354) <= b;
    layer1_outputs(2355) <= '0';
    layer1_outputs(2356) <= not (a and b);
    layer1_outputs(2357) <= '1';
    layer1_outputs(2358) <= not a;
    layer1_outputs(2359) <= '1';
    layer1_outputs(2360) <= '0';
    layer1_outputs(2361) <= not a;
    layer1_outputs(2362) <= not (a or b);
    layer1_outputs(2363) <= '1';
    layer1_outputs(2364) <= a and b;
    layer1_outputs(2365) <= '1';
    layer1_outputs(2366) <= b and not a;
    layer1_outputs(2367) <= b;
    layer1_outputs(2368) <= b and not a;
    layer1_outputs(2369) <= '0';
    layer1_outputs(2370) <= not a;
    layer1_outputs(2371) <= '1';
    layer1_outputs(2372) <= a or b;
    layer1_outputs(2373) <= '0';
    layer1_outputs(2374) <= not (a or b);
    layer1_outputs(2375) <= '0';
    layer1_outputs(2376) <= not b;
    layer1_outputs(2377) <= not a;
    layer1_outputs(2378) <= '0';
    layer1_outputs(2379) <= not b or a;
    layer1_outputs(2380) <= '1';
    layer1_outputs(2381) <= '1';
    layer1_outputs(2382) <= not a or b;
    layer1_outputs(2383) <= a and b;
    layer1_outputs(2384) <= a or b;
    layer1_outputs(2385) <= a;
    layer1_outputs(2386) <= a or b;
    layer1_outputs(2387) <= '1';
    layer1_outputs(2388) <= a;
    layer1_outputs(2389) <= not b or a;
    layer1_outputs(2390) <= not a;
    layer1_outputs(2391) <= not b or a;
    layer1_outputs(2392) <= not b;
    layer1_outputs(2393) <= not (a or b);
    layer1_outputs(2394) <= b and not a;
    layer1_outputs(2395) <= b and not a;
    layer1_outputs(2396) <= not (a or b);
    layer1_outputs(2397) <= a or b;
    layer1_outputs(2398) <= not a or b;
    layer1_outputs(2399) <= not a;
    layer1_outputs(2400) <= a and not b;
    layer1_outputs(2401) <= a and b;
    layer1_outputs(2402) <= not (a xor b);
    layer1_outputs(2403) <= not b or a;
    layer1_outputs(2404) <= '1';
    layer1_outputs(2405) <= not b or a;
    layer1_outputs(2406) <= b and not a;
    layer1_outputs(2407) <= '1';
    layer1_outputs(2408) <= a xor b;
    layer1_outputs(2409) <= a and not b;
    layer1_outputs(2410) <= a and b;
    layer1_outputs(2411) <= '1';
    layer1_outputs(2412) <= b;
    layer1_outputs(2413) <= a and not b;
    layer1_outputs(2414) <= not (a and b);
    layer1_outputs(2415) <= not a;
    layer1_outputs(2416) <= '0';
    layer1_outputs(2417) <= '1';
    layer1_outputs(2418) <= a and b;
    layer1_outputs(2419) <= b and not a;
    layer1_outputs(2420) <= b and not a;
    layer1_outputs(2421) <= a;
    layer1_outputs(2422) <= '0';
    layer1_outputs(2423) <= not (a xor b);
    layer1_outputs(2424) <= '1';
    layer1_outputs(2425) <= not (a or b);
    layer1_outputs(2426) <= not (a or b);
    layer1_outputs(2427) <= '0';
    layer1_outputs(2428) <= not b or a;
    layer1_outputs(2429) <= not (a and b);
    layer1_outputs(2430) <= not a;
    layer1_outputs(2431) <= not b;
    layer1_outputs(2432) <= a;
    layer1_outputs(2433) <= a or b;
    layer1_outputs(2434) <= a;
    layer1_outputs(2435) <= not (a or b);
    layer1_outputs(2436) <= b;
    layer1_outputs(2437) <= not a;
    layer1_outputs(2438) <= a and b;
    layer1_outputs(2439) <= '1';
    layer1_outputs(2440) <= not a;
    layer1_outputs(2441) <= '1';
    layer1_outputs(2442) <= not b or a;
    layer1_outputs(2443) <= '0';
    layer1_outputs(2444) <= a and b;
    layer1_outputs(2445) <= not a;
    layer1_outputs(2446) <= '1';
    layer1_outputs(2447) <= not b;
    layer1_outputs(2448) <= not (a and b);
    layer1_outputs(2449) <= not (a or b);
    layer1_outputs(2450) <= a or b;
    layer1_outputs(2451) <= a and not b;
    layer1_outputs(2452) <= '0';
    layer1_outputs(2453) <= a;
    layer1_outputs(2454) <= not (a or b);
    layer1_outputs(2455) <= '1';
    layer1_outputs(2456) <= not a;
    layer1_outputs(2457) <= a or b;
    layer1_outputs(2458) <= b and not a;
    layer1_outputs(2459) <= a or b;
    layer1_outputs(2460) <= not b;
    layer1_outputs(2461) <= not a or b;
    layer1_outputs(2462) <= not (a or b);
    layer1_outputs(2463) <= not a or b;
    layer1_outputs(2464) <= '0';
    layer1_outputs(2465) <= not b or a;
    layer1_outputs(2466) <= a or b;
    layer1_outputs(2467) <= not b or a;
    layer1_outputs(2468) <= not a;
    layer1_outputs(2469) <= '1';
    layer1_outputs(2470) <= a and not b;
    layer1_outputs(2471) <= a;
    layer1_outputs(2472) <= a or b;
    layer1_outputs(2473) <= b and not a;
    layer1_outputs(2474) <= a;
    layer1_outputs(2475) <= not (a and b);
    layer1_outputs(2476) <= not (a or b);
    layer1_outputs(2477) <= not b;
    layer1_outputs(2478) <= '1';
    layer1_outputs(2479) <= '0';
    layer1_outputs(2480) <= not a or b;
    layer1_outputs(2481) <= b and not a;
    layer1_outputs(2482) <= not b or a;
    layer1_outputs(2483) <= not (a and b);
    layer1_outputs(2484) <= not a;
    layer1_outputs(2485) <= not b;
    layer1_outputs(2486) <= not a or b;
    layer1_outputs(2487) <= not b or a;
    layer1_outputs(2488) <= '0';
    layer1_outputs(2489) <= not a;
    layer1_outputs(2490) <= not (a and b);
    layer1_outputs(2491) <= not b;
    layer1_outputs(2492) <= not (a and b);
    layer1_outputs(2493) <= b and not a;
    layer1_outputs(2494) <= b;
    layer1_outputs(2495) <= '0';
    layer1_outputs(2496) <= '0';
    layer1_outputs(2497) <= not a or b;
    layer1_outputs(2498) <= b;
    layer1_outputs(2499) <= a or b;
    layer1_outputs(2500) <= not (a and b);
    layer1_outputs(2501) <= not a or b;
    layer1_outputs(2502) <= a or b;
    layer1_outputs(2503) <= '0';
    layer1_outputs(2504) <= b;
    layer1_outputs(2505) <= not b or a;
    layer1_outputs(2506) <= not b;
    layer1_outputs(2507) <= b and not a;
    layer1_outputs(2508) <= not b or a;
    layer1_outputs(2509) <= '0';
    layer1_outputs(2510) <= not (a and b);
    layer1_outputs(2511) <= not (a and b);
    layer1_outputs(2512) <= not b or a;
    layer1_outputs(2513) <= a and b;
    layer1_outputs(2514) <= a xor b;
    layer1_outputs(2515) <= not a or b;
    layer1_outputs(2516) <= '1';
    layer1_outputs(2517) <= a and b;
    layer1_outputs(2518) <= not a;
    layer1_outputs(2519) <= '1';
    layer1_outputs(2520) <= a and b;
    layer1_outputs(2521) <= a and not b;
    layer1_outputs(2522) <= not (a xor b);
    layer1_outputs(2523) <= a;
    layer1_outputs(2524) <= '1';
    layer1_outputs(2525) <= not b or a;
    layer1_outputs(2526) <= not a;
    layer1_outputs(2527) <= a;
    layer1_outputs(2528) <= '0';
    layer1_outputs(2529) <= a and not b;
    layer1_outputs(2530) <= not b or a;
    layer1_outputs(2531) <= not a or b;
    layer1_outputs(2532) <= not (a or b);
    layer1_outputs(2533) <= not (a and b);
    layer1_outputs(2534) <= a or b;
    layer1_outputs(2535) <= not b or a;
    layer1_outputs(2536) <= a and b;
    layer1_outputs(2537) <= a or b;
    layer1_outputs(2538) <= '1';
    layer1_outputs(2539) <= a and not b;
    layer1_outputs(2540) <= a or b;
    layer1_outputs(2541) <= '0';
    layer1_outputs(2542) <= a or b;
    layer1_outputs(2543) <= a and not b;
    layer1_outputs(2544) <= not (a or b);
    layer1_outputs(2545) <= b and not a;
    layer1_outputs(2546) <= '0';
    layer1_outputs(2547) <= b and not a;
    layer1_outputs(2548) <= a xor b;
    layer1_outputs(2549) <= a and b;
    layer1_outputs(2550) <= b;
    layer1_outputs(2551) <= not a or b;
    layer1_outputs(2552) <= '0';
    layer1_outputs(2553) <= not a;
    layer1_outputs(2554) <= a or b;
    layer1_outputs(2555) <= '0';
    layer1_outputs(2556) <= b;
    layer1_outputs(2557) <= a or b;
    layer1_outputs(2558) <= not a;
    layer1_outputs(2559) <= b;
    layer1_outputs(2560) <= b;
    layer1_outputs(2561) <= not a;
    layer1_outputs(2562) <= '0';
    layer1_outputs(2563) <= not b or a;
    layer1_outputs(2564) <= '0';
    layer1_outputs(2565) <= b and not a;
    layer1_outputs(2566) <= not (a or b);
    layer1_outputs(2567) <= '1';
    layer1_outputs(2568) <= b;
    layer1_outputs(2569) <= b and not a;
    layer1_outputs(2570) <= a and not b;
    layer1_outputs(2571) <= a xor b;
    layer1_outputs(2572) <= a and b;
    layer1_outputs(2573) <= b and not a;
    layer1_outputs(2574) <= a;
    layer1_outputs(2575) <= not (a or b);
    layer1_outputs(2576) <= a and b;
    layer1_outputs(2577) <= a and b;
    layer1_outputs(2578) <= not (a xor b);
    layer1_outputs(2579) <= a and b;
    layer1_outputs(2580) <= not a or b;
    layer1_outputs(2581) <= b;
    layer1_outputs(2582) <= '1';
    layer1_outputs(2583) <= '1';
    layer1_outputs(2584) <= a xor b;
    layer1_outputs(2585) <= not b;
    layer1_outputs(2586) <= not b or a;
    layer1_outputs(2587) <= not b;
    layer1_outputs(2588) <= '1';
    layer1_outputs(2589) <= '0';
    layer1_outputs(2590) <= b;
    layer1_outputs(2591) <= '0';
    layer1_outputs(2592) <= not (a and b);
    layer1_outputs(2593) <= not (a and b);
    layer1_outputs(2594) <= a xor b;
    layer1_outputs(2595) <= '1';
    layer1_outputs(2596) <= '0';
    layer1_outputs(2597) <= a or b;
    layer1_outputs(2598) <= not b;
    layer1_outputs(2599) <= a;
    layer1_outputs(2600) <= not a or b;
    layer1_outputs(2601) <= a xor b;
    layer1_outputs(2602) <= a and b;
    layer1_outputs(2603) <= not b or a;
    layer1_outputs(2604) <= '0';
    layer1_outputs(2605) <= b and not a;
    layer1_outputs(2606) <= a;
    layer1_outputs(2607) <= not b;
    layer1_outputs(2608) <= not (a and b);
    layer1_outputs(2609) <= not b or a;
    layer1_outputs(2610) <= b and not a;
    layer1_outputs(2611) <= not a;
    layer1_outputs(2612) <= '1';
    layer1_outputs(2613) <= not b or a;
    layer1_outputs(2614) <= b and not a;
    layer1_outputs(2615) <= b and not a;
    layer1_outputs(2616) <= not a or b;
    layer1_outputs(2617) <= not (a xor b);
    layer1_outputs(2618) <= not (a or b);
    layer1_outputs(2619) <= not b;
    layer1_outputs(2620) <= b and not a;
    layer1_outputs(2621) <= '0';
    layer1_outputs(2622) <= not b;
    layer1_outputs(2623) <= not b;
    layer1_outputs(2624) <= a and not b;
    layer1_outputs(2625) <= a;
    layer1_outputs(2626) <= a and b;
    layer1_outputs(2627) <= not b or a;
    layer1_outputs(2628) <= '0';
    layer1_outputs(2629) <= b and not a;
    layer1_outputs(2630) <= not (a or b);
    layer1_outputs(2631) <= '1';
    layer1_outputs(2632) <= a and b;
    layer1_outputs(2633) <= a or b;
    layer1_outputs(2634) <= not a or b;
    layer1_outputs(2635) <= not (a or b);
    layer1_outputs(2636) <= not (a or b);
    layer1_outputs(2637) <= not b;
    layer1_outputs(2638) <= a and b;
    layer1_outputs(2639) <= '0';
    layer1_outputs(2640) <= not b or a;
    layer1_outputs(2641) <= a and not b;
    layer1_outputs(2642) <= not a;
    layer1_outputs(2643) <= not a or b;
    layer1_outputs(2644) <= not b or a;
    layer1_outputs(2645) <= a or b;
    layer1_outputs(2646) <= a and b;
    layer1_outputs(2647) <= not (a xor b);
    layer1_outputs(2648) <= b;
    layer1_outputs(2649) <= not a;
    layer1_outputs(2650) <= a and b;
    layer1_outputs(2651) <= not b;
    layer1_outputs(2652) <= b and not a;
    layer1_outputs(2653) <= b;
    layer1_outputs(2654) <= not a;
    layer1_outputs(2655) <= not a or b;
    layer1_outputs(2656) <= not (a and b);
    layer1_outputs(2657) <= not (a and b);
    layer1_outputs(2658) <= a and b;
    layer1_outputs(2659) <= not b;
    layer1_outputs(2660) <= not b;
    layer1_outputs(2661) <= a or b;
    layer1_outputs(2662) <= '0';
    layer1_outputs(2663) <= a or b;
    layer1_outputs(2664) <= not (a and b);
    layer1_outputs(2665) <= a and not b;
    layer1_outputs(2666) <= '1';
    layer1_outputs(2667) <= b and not a;
    layer1_outputs(2668) <= '1';
    layer1_outputs(2669) <= '1';
    layer1_outputs(2670) <= not b or a;
    layer1_outputs(2671) <= not b or a;
    layer1_outputs(2672) <= not a;
    layer1_outputs(2673) <= not b;
    layer1_outputs(2674) <= not (a xor b);
    layer1_outputs(2675) <= a and b;
    layer1_outputs(2676) <= a;
    layer1_outputs(2677) <= not b;
    layer1_outputs(2678) <= not b or a;
    layer1_outputs(2679) <= a and not b;
    layer1_outputs(2680) <= not b or a;
    layer1_outputs(2681) <= not b or a;
    layer1_outputs(2682) <= not (a and b);
    layer1_outputs(2683) <= a and not b;
    layer1_outputs(2684) <= '0';
    layer1_outputs(2685) <= b;
    layer1_outputs(2686) <= not a or b;
    layer1_outputs(2687) <= not b or a;
    layer1_outputs(2688) <= a;
    layer1_outputs(2689) <= '0';
    layer1_outputs(2690) <= '1';
    layer1_outputs(2691) <= '0';
    layer1_outputs(2692) <= not (a and b);
    layer1_outputs(2693) <= '1';
    layer1_outputs(2694) <= not (a and b);
    layer1_outputs(2695) <= b;
    layer1_outputs(2696) <= '0';
    layer1_outputs(2697) <= b and not a;
    layer1_outputs(2698) <= '0';
    layer1_outputs(2699) <= not a or b;
    layer1_outputs(2700) <= not b or a;
    layer1_outputs(2701) <= b and not a;
    layer1_outputs(2702) <= a;
    layer1_outputs(2703) <= a or b;
    layer1_outputs(2704) <= b and not a;
    layer1_outputs(2705) <= not b;
    layer1_outputs(2706) <= a or b;
    layer1_outputs(2707) <= b;
    layer1_outputs(2708) <= '1';
    layer1_outputs(2709) <= a;
    layer1_outputs(2710) <= a and b;
    layer1_outputs(2711) <= b and not a;
    layer1_outputs(2712) <= not a or b;
    layer1_outputs(2713) <= '1';
    layer1_outputs(2714) <= not b or a;
    layer1_outputs(2715) <= a or b;
    layer1_outputs(2716) <= '0';
    layer1_outputs(2717) <= a and not b;
    layer1_outputs(2718) <= '0';
    layer1_outputs(2719) <= '1';
    layer1_outputs(2720) <= not b;
    layer1_outputs(2721) <= a;
    layer1_outputs(2722) <= b and not a;
    layer1_outputs(2723) <= '1';
    layer1_outputs(2724) <= not b or a;
    layer1_outputs(2725) <= b;
    layer1_outputs(2726) <= not a;
    layer1_outputs(2727) <= a or b;
    layer1_outputs(2728) <= a and not b;
    layer1_outputs(2729) <= not b or a;
    layer1_outputs(2730) <= a and b;
    layer1_outputs(2731) <= not b or a;
    layer1_outputs(2732) <= not a or b;
    layer1_outputs(2733) <= '0';
    layer1_outputs(2734) <= b;
    layer1_outputs(2735) <= not (a and b);
    layer1_outputs(2736) <= not a;
    layer1_outputs(2737) <= not (a and b);
    layer1_outputs(2738) <= a and b;
    layer1_outputs(2739) <= a and b;
    layer1_outputs(2740) <= a xor b;
    layer1_outputs(2741) <= not (a xor b);
    layer1_outputs(2742) <= b;
    layer1_outputs(2743) <= '1';
    layer1_outputs(2744) <= not a or b;
    layer1_outputs(2745) <= not (a or b);
    layer1_outputs(2746) <= '0';
    layer1_outputs(2747) <= not (a or b);
    layer1_outputs(2748) <= a and b;
    layer1_outputs(2749) <= not b or a;
    layer1_outputs(2750) <= not (a or b);
    layer1_outputs(2751) <= '1';
    layer1_outputs(2752) <= b and not a;
    layer1_outputs(2753) <= not a or b;
    layer1_outputs(2754) <= not a;
    layer1_outputs(2755) <= '0';
    layer1_outputs(2756) <= not (a and b);
    layer1_outputs(2757) <= not (a or b);
    layer1_outputs(2758) <= b and not a;
    layer1_outputs(2759) <= not (a and b);
    layer1_outputs(2760) <= a and not b;
    layer1_outputs(2761) <= a and b;
    layer1_outputs(2762) <= not a or b;
    layer1_outputs(2763) <= '0';
    layer1_outputs(2764) <= '0';
    layer1_outputs(2765) <= a;
    layer1_outputs(2766) <= a and b;
    layer1_outputs(2767) <= not (a xor b);
    layer1_outputs(2768) <= a and not b;
    layer1_outputs(2769) <= not b or a;
    layer1_outputs(2770) <= '0';
    layer1_outputs(2771) <= not b;
    layer1_outputs(2772) <= '0';
    layer1_outputs(2773) <= not b or a;
    layer1_outputs(2774) <= not (a or b);
    layer1_outputs(2775) <= not (a or b);
    layer1_outputs(2776) <= '0';
    layer1_outputs(2777) <= a or b;
    layer1_outputs(2778) <= a xor b;
    layer1_outputs(2779) <= a;
    layer1_outputs(2780) <= not b or a;
    layer1_outputs(2781) <= a and b;
    layer1_outputs(2782) <= not a;
    layer1_outputs(2783) <= '0';
    layer1_outputs(2784) <= not (a and b);
    layer1_outputs(2785) <= a and not b;
    layer1_outputs(2786) <= b and not a;
    layer1_outputs(2787) <= b;
    layer1_outputs(2788) <= not a;
    layer1_outputs(2789) <= a and not b;
    layer1_outputs(2790) <= a and not b;
    layer1_outputs(2791) <= a or b;
    layer1_outputs(2792) <= not b or a;
    layer1_outputs(2793) <= not (a and b);
    layer1_outputs(2794) <= a and not b;
    layer1_outputs(2795) <= a and b;
    layer1_outputs(2796) <= not a;
    layer1_outputs(2797) <= '1';
    layer1_outputs(2798) <= not b or a;
    layer1_outputs(2799) <= a or b;
    layer1_outputs(2800) <= b;
    layer1_outputs(2801) <= a and not b;
    layer1_outputs(2802) <= not (a and b);
    layer1_outputs(2803) <= a or b;
    layer1_outputs(2804) <= b and not a;
    layer1_outputs(2805) <= not a;
    layer1_outputs(2806) <= '1';
    layer1_outputs(2807) <= not a or b;
    layer1_outputs(2808) <= not (a and b);
    layer1_outputs(2809) <= a or b;
    layer1_outputs(2810) <= not (a or b);
    layer1_outputs(2811) <= not b;
    layer1_outputs(2812) <= not b or a;
    layer1_outputs(2813) <= '0';
    layer1_outputs(2814) <= not a or b;
    layer1_outputs(2815) <= not a or b;
    layer1_outputs(2816) <= not b or a;
    layer1_outputs(2817) <= not (a and b);
    layer1_outputs(2818) <= not (a and b);
    layer1_outputs(2819) <= not (a or b);
    layer1_outputs(2820) <= a;
    layer1_outputs(2821) <= a and not b;
    layer1_outputs(2822) <= a and not b;
    layer1_outputs(2823) <= a xor b;
    layer1_outputs(2824) <= not b or a;
    layer1_outputs(2825) <= a and b;
    layer1_outputs(2826) <= a and b;
    layer1_outputs(2827) <= a and b;
    layer1_outputs(2828) <= not (a and b);
    layer1_outputs(2829) <= b;
    layer1_outputs(2830) <= '0';
    layer1_outputs(2831) <= not b or a;
    layer1_outputs(2832) <= '0';
    layer1_outputs(2833) <= b and not a;
    layer1_outputs(2834) <= '0';
    layer1_outputs(2835) <= not (a and b);
    layer1_outputs(2836) <= '1';
    layer1_outputs(2837) <= not (a and b);
    layer1_outputs(2838) <= '1';
    layer1_outputs(2839) <= not (a or b);
    layer1_outputs(2840) <= a and b;
    layer1_outputs(2841) <= '0';
    layer1_outputs(2842) <= a xor b;
    layer1_outputs(2843) <= not a or b;
    layer1_outputs(2844) <= not a or b;
    layer1_outputs(2845) <= not (a or b);
    layer1_outputs(2846) <= '1';
    layer1_outputs(2847) <= not a or b;
    layer1_outputs(2848) <= not (a or b);
    layer1_outputs(2849) <= '1';
    layer1_outputs(2850) <= '1';
    layer1_outputs(2851) <= a and not b;
    layer1_outputs(2852) <= '0';
    layer1_outputs(2853) <= '0';
    layer1_outputs(2854) <= not (a and b);
    layer1_outputs(2855) <= not a;
    layer1_outputs(2856) <= b and not a;
    layer1_outputs(2857) <= b;
    layer1_outputs(2858) <= a;
    layer1_outputs(2859) <= '0';
    layer1_outputs(2860) <= not a;
    layer1_outputs(2861) <= not a or b;
    layer1_outputs(2862) <= not (a and b);
    layer1_outputs(2863) <= not a;
    layer1_outputs(2864) <= not (a and b);
    layer1_outputs(2865) <= a and not b;
    layer1_outputs(2866) <= a and not b;
    layer1_outputs(2867) <= not a or b;
    layer1_outputs(2868) <= not b;
    layer1_outputs(2869) <= not b;
    layer1_outputs(2870) <= not a;
    layer1_outputs(2871) <= a and b;
    layer1_outputs(2872) <= b;
    layer1_outputs(2873) <= a;
    layer1_outputs(2874) <= a or b;
    layer1_outputs(2875) <= not a;
    layer1_outputs(2876) <= '1';
    layer1_outputs(2877) <= a and not b;
    layer1_outputs(2878) <= '1';
    layer1_outputs(2879) <= not (a and b);
    layer1_outputs(2880) <= b;
    layer1_outputs(2881) <= '0';
    layer1_outputs(2882) <= not a;
    layer1_outputs(2883) <= a and b;
    layer1_outputs(2884) <= '0';
    layer1_outputs(2885) <= not (a and b);
    layer1_outputs(2886) <= a;
    layer1_outputs(2887) <= not (a and b);
    layer1_outputs(2888) <= not (a xor b);
    layer1_outputs(2889) <= '1';
    layer1_outputs(2890) <= a and not b;
    layer1_outputs(2891) <= not a or b;
    layer1_outputs(2892) <= a;
    layer1_outputs(2893) <= '1';
    layer1_outputs(2894) <= not a;
    layer1_outputs(2895) <= b;
    layer1_outputs(2896) <= a xor b;
    layer1_outputs(2897) <= not b or a;
    layer1_outputs(2898) <= not (a or b);
    layer1_outputs(2899) <= a xor b;
    layer1_outputs(2900) <= b;
    layer1_outputs(2901) <= a;
    layer1_outputs(2902) <= '1';
    layer1_outputs(2903) <= a or b;
    layer1_outputs(2904) <= '0';
    layer1_outputs(2905) <= not b;
    layer1_outputs(2906) <= a xor b;
    layer1_outputs(2907) <= not a or b;
    layer1_outputs(2908) <= not (a xor b);
    layer1_outputs(2909) <= a or b;
    layer1_outputs(2910) <= '1';
    layer1_outputs(2911) <= not a or b;
    layer1_outputs(2912) <= not a or b;
    layer1_outputs(2913) <= b and not a;
    layer1_outputs(2914) <= a and not b;
    layer1_outputs(2915) <= not a or b;
    layer1_outputs(2916) <= not a or b;
    layer1_outputs(2917) <= b and not a;
    layer1_outputs(2918) <= not (a or b);
    layer1_outputs(2919) <= not b;
    layer1_outputs(2920) <= a and not b;
    layer1_outputs(2921) <= b and not a;
    layer1_outputs(2922) <= not b;
    layer1_outputs(2923) <= b;
    layer1_outputs(2924) <= not (a and b);
    layer1_outputs(2925) <= not (a or b);
    layer1_outputs(2926) <= '1';
    layer1_outputs(2927) <= a or b;
    layer1_outputs(2928) <= not a or b;
    layer1_outputs(2929) <= b and not a;
    layer1_outputs(2930) <= a and b;
    layer1_outputs(2931) <= '1';
    layer1_outputs(2932) <= a or b;
    layer1_outputs(2933) <= '0';
    layer1_outputs(2934) <= not a;
    layer1_outputs(2935) <= not (a or b);
    layer1_outputs(2936) <= not b or a;
    layer1_outputs(2937) <= not b;
    layer1_outputs(2938) <= not (a xor b);
    layer1_outputs(2939) <= not a;
    layer1_outputs(2940) <= not (a and b);
    layer1_outputs(2941) <= not b or a;
    layer1_outputs(2942) <= not (a and b);
    layer1_outputs(2943) <= not b or a;
    layer1_outputs(2944) <= '1';
    layer1_outputs(2945) <= b and not a;
    layer1_outputs(2946) <= not (a xor b);
    layer1_outputs(2947) <= '1';
    layer1_outputs(2948) <= a and b;
    layer1_outputs(2949) <= not b or a;
    layer1_outputs(2950) <= a or b;
    layer1_outputs(2951) <= a and b;
    layer1_outputs(2952) <= not a;
    layer1_outputs(2953) <= a;
    layer1_outputs(2954) <= a;
    layer1_outputs(2955) <= not (a and b);
    layer1_outputs(2956) <= a and not b;
    layer1_outputs(2957) <= not a or b;
    layer1_outputs(2958) <= '0';
    layer1_outputs(2959) <= not a or b;
    layer1_outputs(2960) <= not (a xor b);
    layer1_outputs(2961) <= not b;
    layer1_outputs(2962) <= a or b;
    layer1_outputs(2963) <= not b or a;
    layer1_outputs(2964) <= '0';
    layer1_outputs(2965) <= '1';
    layer1_outputs(2966) <= '1';
    layer1_outputs(2967) <= a or b;
    layer1_outputs(2968) <= not a or b;
    layer1_outputs(2969) <= a;
    layer1_outputs(2970) <= a or b;
    layer1_outputs(2971) <= b;
    layer1_outputs(2972) <= a and b;
    layer1_outputs(2973) <= '1';
    layer1_outputs(2974) <= a and not b;
    layer1_outputs(2975) <= b and not a;
    layer1_outputs(2976) <= not (a and b);
    layer1_outputs(2977) <= not (a xor b);
    layer1_outputs(2978) <= b and not a;
    layer1_outputs(2979) <= a and b;
    layer1_outputs(2980) <= a and b;
    layer1_outputs(2981) <= a and b;
    layer1_outputs(2982) <= b and not a;
    layer1_outputs(2983) <= a;
    layer1_outputs(2984) <= not (a or b);
    layer1_outputs(2985) <= b;
    layer1_outputs(2986) <= a and not b;
    layer1_outputs(2987) <= a or b;
    layer1_outputs(2988) <= not a;
    layer1_outputs(2989) <= not a or b;
    layer1_outputs(2990) <= b;
    layer1_outputs(2991) <= not (a and b);
    layer1_outputs(2992) <= a and not b;
    layer1_outputs(2993) <= not b;
    layer1_outputs(2994) <= not (a or b);
    layer1_outputs(2995) <= b;
    layer1_outputs(2996) <= a and not b;
    layer1_outputs(2997) <= a and b;
    layer1_outputs(2998) <= not (a and b);
    layer1_outputs(2999) <= not (a or b);
    layer1_outputs(3000) <= a and b;
    layer1_outputs(3001) <= not (a and b);
    layer1_outputs(3002) <= not a;
    layer1_outputs(3003) <= not a;
    layer1_outputs(3004) <= a and not b;
    layer1_outputs(3005) <= b and not a;
    layer1_outputs(3006) <= a or b;
    layer1_outputs(3007) <= b;
    layer1_outputs(3008) <= '0';
    layer1_outputs(3009) <= '0';
    layer1_outputs(3010) <= a or b;
    layer1_outputs(3011) <= not (a or b);
    layer1_outputs(3012) <= not (a xor b);
    layer1_outputs(3013) <= a and b;
    layer1_outputs(3014) <= a or b;
    layer1_outputs(3015) <= not b;
    layer1_outputs(3016) <= not b;
    layer1_outputs(3017) <= '0';
    layer1_outputs(3018) <= not (a and b);
    layer1_outputs(3019) <= not b;
    layer1_outputs(3020) <= not b;
    layer1_outputs(3021) <= a and b;
    layer1_outputs(3022) <= not b or a;
    layer1_outputs(3023) <= not a or b;
    layer1_outputs(3024) <= '1';
    layer1_outputs(3025) <= a;
    layer1_outputs(3026) <= b and not a;
    layer1_outputs(3027) <= not (a or b);
    layer1_outputs(3028) <= '1';
    layer1_outputs(3029) <= not b or a;
    layer1_outputs(3030) <= not (a or b);
    layer1_outputs(3031) <= '0';
    layer1_outputs(3032) <= a;
    layer1_outputs(3033) <= a and b;
    layer1_outputs(3034) <= '0';
    layer1_outputs(3035) <= a or b;
    layer1_outputs(3036) <= b and not a;
    layer1_outputs(3037) <= '0';
    layer1_outputs(3038) <= b;
    layer1_outputs(3039) <= a and b;
    layer1_outputs(3040) <= not b or a;
    layer1_outputs(3041) <= '0';
    layer1_outputs(3042) <= not a or b;
    layer1_outputs(3043) <= not (a and b);
    layer1_outputs(3044) <= not (a and b);
    layer1_outputs(3045) <= '1';
    layer1_outputs(3046) <= a;
    layer1_outputs(3047) <= '1';
    layer1_outputs(3048) <= a and not b;
    layer1_outputs(3049) <= b;
    layer1_outputs(3050) <= not b or a;
    layer1_outputs(3051) <= not (a or b);
    layer1_outputs(3052) <= '1';
    layer1_outputs(3053) <= not a;
    layer1_outputs(3054) <= not (a or b);
    layer1_outputs(3055) <= not b;
    layer1_outputs(3056) <= '1';
    layer1_outputs(3057) <= not b;
    layer1_outputs(3058) <= '1';
    layer1_outputs(3059) <= '1';
    layer1_outputs(3060) <= a;
    layer1_outputs(3061) <= not b or a;
    layer1_outputs(3062) <= b;
    layer1_outputs(3063) <= a;
    layer1_outputs(3064) <= not b;
    layer1_outputs(3065) <= a;
    layer1_outputs(3066) <= a;
    layer1_outputs(3067) <= b;
    layer1_outputs(3068) <= not a or b;
    layer1_outputs(3069) <= a and b;
    layer1_outputs(3070) <= not a or b;
    layer1_outputs(3071) <= a and b;
    layer1_outputs(3072) <= not (a or b);
    layer1_outputs(3073) <= a and not b;
    layer1_outputs(3074) <= a or b;
    layer1_outputs(3075) <= a or b;
    layer1_outputs(3076) <= not b;
    layer1_outputs(3077) <= b;
    layer1_outputs(3078) <= b and not a;
    layer1_outputs(3079) <= a or b;
    layer1_outputs(3080) <= not b or a;
    layer1_outputs(3081) <= not a or b;
    layer1_outputs(3082) <= not b or a;
    layer1_outputs(3083) <= not a or b;
    layer1_outputs(3084) <= not a;
    layer1_outputs(3085) <= not a;
    layer1_outputs(3086) <= not a;
    layer1_outputs(3087) <= '0';
    layer1_outputs(3088) <= a and b;
    layer1_outputs(3089) <= a and not b;
    layer1_outputs(3090) <= not b or a;
    layer1_outputs(3091) <= '1';
    layer1_outputs(3092) <= '1';
    layer1_outputs(3093) <= a;
    layer1_outputs(3094) <= a or b;
    layer1_outputs(3095) <= b;
    layer1_outputs(3096) <= not (a xor b);
    layer1_outputs(3097) <= '1';
    layer1_outputs(3098) <= not a;
    layer1_outputs(3099) <= not b;
    layer1_outputs(3100) <= not a;
    layer1_outputs(3101) <= not b or a;
    layer1_outputs(3102) <= a;
    layer1_outputs(3103) <= '0';
    layer1_outputs(3104) <= a;
    layer1_outputs(3105) <= b;
    layer1_outputs(3106) <= a and b;
    layer1_outputs(3107) <= not b;
    layer1_outputs(3108) <= '1';
    layer1_outputs(3109) <= not (a and b);
    layer1_outputs(3110) <= a;
    layer1_outputs(3111) <= a and not b;
    layer1_outputs(3112) <= not a;
    layer1_outputs(3113) <= not (a or b);
    layer1_outputs(3114) <= not a or b;
    layer1_outputs(3115) <= '0';
    layer1_outputs(3116) <= not a or b;
    layer1_outputs(3117) <= not (a and b);
    layer1_outputs(3118) <= not a;
    layer1_outputs(3119) <= b;
    layer1_outputs(3120) <= a;
    layer1_outputs(3121) <= not (a xor b);
    layer1_outputs(3122) <= not (a and b);
    layer1_outputs(3123) <= a;
    layer1_outputs(3124) <= '0';
    layer1_outputs(3125) <= '0';
    layer1_outputs(3126) <= a;
    layer1_outputs(3127) <= not b;
    layer1_outputs(3128) <= a or b;
    layer1_outputs(3129) <= not b or a;
    layer1_outputs(3130) <= '1';
    layer1_outputs(3131) <= '1';
    layer1_outputs(3132) <= b;
    layer1_outputs(3133) <= not (a xor b);
    layer1_outputs(3134) <= b and not a;
    layer1_outputs(3135) <= '0';
    layer1_outputs(3136) <= a and not b;
    layer1_outputs(3137) <= a and not b;
    layer1_outputs(3138) <= not (a or b);
    layer1_outputs(3139) <= not b or a;
    layer1_outputs(3140) <= '0';
    layer1_outputs(3141) <= b;
    layer1_outputs(3142) <= '0';
    layer1_outputs(3143) <= '0';
    layer1_outputs(3144) <= b and not a;
    layer1_outputs(3145) <= a and not b;
    layer1_outputs(3146) <= a or b;
    layer1_outputs(3147) <= not (a or b);
    layer1_outputs(3148) <= a and not b;
    layer1_outputs(3149) <= '1';
    layer1_outputs(3150) <= not a or b;
    layer1_outputs(3151) <= a and not b;
    layer1_outputs(3152) <= '1';
    layer1_outputs(3153) <= not a or b;
    layer1_outputs(3154) <= '1';
    layer1_outputs(3155) <= b;
    layer1_outputs(3156) <= a;
    layer1_outputs(3157) <= b;
    layer1_outputs(3158) <= not b;
    layer1_outputs(3159) <= not (a or b);
    layer1_outputs(3160) <= '1';
    layer1_outputs(3161) <= '0';
    layer1_outputs(3162) <= b and not a;
    layer1_outputs(3163) <= not a or b;
    layer1_outputs(3164) <= not (a and b);
    layer1_outputs(3165) <= b and not a;
    layer1_outputs(3166) <= not b or a;
    layer1_outputs(3167) <= not (a and b);
    layer1_outputs(3168) <= not (a or b);
    layer1_outputs(3169) <= not b;
    layer1_outputs(3170) <= b and not a;
    layer1_outputs(3171) <= '0';
    layer1_outputs(3172) <= not (a or b);
    layer1_outputs(3173) <= not a;
    layer1_outputs(3174) <= '1';
    layer1_outputs(3175) <= b;
    layer1_outputs(3176) <= '0';
    layer1_outputs(3177) <= a and b;
    layer1_outputs(3178) <= a;
    layer1_outputs(3179) <= '0';
    layer1_outputs(3180) <= not (a xor b);
    layer1_outputs(3181) <= b and not a;
    layer1_outputs(3182) <= b and not a;
    layer1_outputs(3183) <= b and not a;
    layer1_outputs(3184) <= '1';
    layer1_outputs(3185) <= not (a and b);
    layer1_outputs(3186) <= not (a or b);
    layer1_outputs(3187) <= not a;
    layer1_outputs(3188) <= a or b;
    layer1_outputs(3189) <= not (a or b);
    layer1_outputs(3190) <= '0';
    layer1_outputs(3191) <= '0';
    layer1_outputs(3192) <= a and b;
    layer1_outputs(3193) <= a;
    layer1_outputs(3194) <= a and not b;
    layer1_outputs(3195) <= not b or a;
    layer1_outputs(3196) <= a and not b;
    layer1_outputs(3197) <= a and not b;
    layer1_outputs(3198) <= a and not b;
    layer1_outputs(3199) <= a or b;
    layer1_outputs(3200) <= '1';
    layer1_outputs(3201) <= not b or a;
    layer1_outputs(3202) <= a and b;
    layer1_outputs(3203) <= not (a or b);
    layer1_outputs(3204) <= '1';
    layer1_outputs(3205) <= b;
    layer1_outputs(3206) <= a and b;
    layer1_outputs(3207) <= '1';
    layer1_outputs(3208) <= a and b;
    layer1_outputs(3209) <= b;
    layer1_outputs(3210) <= a and b;
    layer1_outputs(3211) <= not (a and b);
    layer1_outputs(3212) <= not a;
    layer1_outputs(3213) <= a and not b;
    layer1_outputs(3214) <= b;
    layer1_outputs(3215) <= '1';
    layer1_outputs(3216) <= '1';
    layer1_outputs(3217) <= '1';
    layer1_outputs(3218) <= a and not b;
    layer1_outputs(3219) <= a or b;
    layer1_outputs(3220) <= a or b;
    layer1_outputs(3221) <= '1';
    layer1_outputs(3222) <= b;
    layer1_outputs(3223) <= not (a and b);
    layer1_outputs(3224) <= not (a or b);
    layer1_outputs(3225) <= a or b;
    layer1_outputs(3226) <= b;
    layer1_outputs(3227) <= not a;
    layer1_outputs(3228) <= a and not b;
    layer1_outputs(3229) <= not b or a;
    layer1_outputs(3230) <= a;
    layer1_outputs(3231) <= not (a or b);
    layer1_outputs(3232) <= not b;
    layer1_outputs(3233) <= not (a or b);
    layer1_outputs(3234) <= '1';
    layer1_outputs(3235) <= b;
    layer1_outputs(3236) <= not a or b;
    layer1_outputs(3237) <= not (a and b);
    layer1_outputs(3238) <= not (a or b);
    layer1_outputs(3239) <= a;
    layer1_outputs(3240) <= a and b;
    layer1_outputs(3241) <= '0';
    layer1_outputs(3242) <= a or b;
    layer1_outputs(3243) <= a or b;
    layer1_outputs(3244) <= a and b;
    layer1_outputs(3245) <= a xor b;
    layer1_outputs(3246) <= a;
    layer1_outputs(3247) <= a;
    layer1_outputs(3248) <= a;
    layer1_outputs(3249) <= a and not b;
    layer1_outputs(3250) <= '1';
    layer1_outputs(3251) <= '0';
    layer1_outputs(3252) <= not b;
    layer1_outputs(3253) <= not b or a;
    layer1_outputs(3254) <= '1';
    layer1_outputs(3255) <= not b;
    layer1_outputs(3256) <= a;
    layer1_outputs(3257) <= a or b;
    layer1_outputs(3258) <= a and not b;
    layer1_outputs(3259) <= not b or a;
    layer1_outputs(3260) <= b and not a;
    layer1_outputs(3261) <= a;
    layer1_outputs(3262) <= a and not b;
    layer1_outputs(3263) <= b;
    layer1_outputs(3264) <= b and not a;
    layer1_outputs(3265) <= a and not b;
    layer1_outputs(3266) <= a;
    layer1_outputs(3267) <= not b or a;
    layer1_outputs(3268) <= a and b;
    layer1_outputs(3269) <= not (a and b);
    layer1_outputs(3270) <= b and not a;
    layer1_outputs(3271) <= a;
    layer1_outputs(3272) <= a xor b;
    layer1_outputs(3273) <= '0';
    layer1_outputs(3274) <= not (a or b);
    layer1_outputs(3275) <= b;
    layer1_outputs(3276) <= '0';
    layer1_outputs(3277) <= not b;
    layer1_outputs(3278) <= a and b;
    layer1_outputs(3279) <= a or b;
    layer1_outputs(3280) <= not a;
    layer1_outputs(3281) <= '1';
    layer1_outputs(3282) <= '1';
    layer1_outputs(3283) <= not (a and b);
    layer1_outputs(3284) <= not (a and b);
    layer1_outputs(3285) <= a;
    layer1_outputs(3286) <= a xor b;
    layer1_outputs(3287) <= b and not a;
    layer1_outputs(3288) <= b and not a;
    layer1_outputs(3289) <= a and not b;
    layer1_outputs(3290) <= not (a and b);
    layer1_outputs(3291) <= not a;
    layer1_outputs(3292) <= not a;
    layer1_outputs(3293) <= not a or b;
    layer1_outputs(3294) <= '1';
    layer1_outputs(3295) <= not (a and b);
    layer1_outputs(3296) <= not b or a;
    layer1_outputs(3297) <= not a;
    layer1_outputs(3298) <= not b or a;
    layer1_outputs(3299) <= not (a or b);
    layer1_outputs(3300) <= a and not b;
    layer1_outputs(3301) <= a xor b;
    layer1_outputs(3302) <= not a;
    layer1_outputs(3303) <= '0';
    layer1_outputs(3304) <= a or b;
    layer1_outputs(3305) <= a;
    layer1_outputs(3306) <= not (a xor b);
    layer1_outputs(3307) <= a;
    layer1_outputs(3308) <= not a or b;
    layer1_outputs(3309) <= '0';
    layer1_outputs(3310) <= not a;
    layer1_outputs(3311) <= '1';
    layer1_outputs(3312) <= a;
    layer1_outputs(3313) <= a;
    layer1_outputs(3314) <= a and b;
    layer1_outputs(3315) <= not (a or b);
    layer1_outputs(3316) <= not (a xor b);
    layer1_outputs(3317) <= '0';
    layer1_outputs(3318) <= not (a or b);
    layer1_outputs(3319) <= not b;
    layer1_outputs(3320) <= not (a and b);
    layer1_outputs(3321) <= a or b;
    layer1_outputs(3322) <= not b;
    layer1_outputs(3323) <= '0';
    layer1_outputs(3324) <= not a;
    layer1_outputs(3325) <= not b or a;
    layer1_outputs(3326) <= a and b;
    layer1_outputs(3327) <= b and not a;
    layer1_outputs(3328) <= a and b;
    layer1_outputs(3329) <= a and not b;
    layer1_outputs(3330) <= not b or a;
    layer1_outputs(3331) <= not a;
    layer1_outputs(3332) <= not (a and b);
    layer1_outputs(3333) <= a or b;
    layer1_outputs(3334) <= not a or b;
    layer1_outputs(3335) <= not a or b;
    layer1_outputs(3336) <= '1';
    layer1_outputs(3337) <= b;
    layer1_outputs(3338) <= not a or b;
    layer1_outputs(3339) <= a and b;
    layer1_outputs(3340) <= '0';
    layer1_outputs(3341) <= a and not b;
    layer1_outputs(3342) <= not (a or b);
    layer1_outputs(3343) <= not (a and b);
    layer1_outputs(3344) <= '1';
    layer1_outputs(3345) <= not a or b;
    layer1_outputs(3346) <= not b or a;
    layer1_outputs(3347) <= not a or b;
    layer1_outputs(3348) <= '0';
    layer1_outputs(3349) <= not (a and b);
    layer1_outputs(3350) <= '0';
    layer1_outputs(3351) <= not b;
    layer1_outputs(3352) <= b and not a;
    layer1_outputs(3353) <= '1';
    layer1_outputs(3354) <= a;
    layer1_outputs(3355) <= b and not a;
    layer1_outputs(3356) <= not b;
    layer1_outputs(3357) <= a and b;
    layer1_outputs(3358) <= not b;
    layer1_outputs(3359) <= b and not a;
    layer1_outputs(3360) <= not (a and b);
    layer1_outputs(3361) <= not a or b;
    layer1_outputs(3362) <= a and b;
    layer1_outputs(3363) <= a and b;
    layer1_outputs(3364) <= b and not a;
    layer1_outputs(3365) <= not a;
    layer1_outputs(3366) <= not (a and b);
    layer1_outputs(3367) <= a and b;
    layer1_outputs(3368) <= not b or a;
    layer1_outputs(3369) <= a or b;
    layer1_outputs(3370) <= '1';
    layer1_outputs(3371) <= '1';
    layer1_outputs(3372) <= not (a xor b);
    layer1_outputs(3373) <= not a;
    layer1_outputs(3374) <= not a;
    layer1_outputs(3375) <= '1';
    layer1_outputs(3376) <= not a or b;
    layer1_outputs(3377) <= not a or b;
    layer1_outputs(3378) <= not b;
    layer1_outputs(3379) <= not (a and b);
    layer1_outputs(3380) <= a and not b;
    layer1_outputs(3381) <= '0';
    layer1_outputs(3382) <= '1';
    layer1_outputs(3383) <= not (a or b);
    layer1_outputs(3384) <= not b or a;
    layer1_outputs(3385) <= not b or a;
    layer1_outputs(3386) <= a or b;
    layer1_outputs(3387) <= not (a xor b);
    layer1_outputs(3388) <= not b or a;
    layer1_outputs(3389) <= b;
    layer1_outputs(3390) <= '1';
    layer1_outputs(3391) <= a and not b;
    layer1_outputs(3392) <= not b or a;
    layer1_outputs(3393) <= a or b;
    layer1_outputs(3394) <= '0';
    layer1_outputs(3395) <= not (a and b);
    layer1_outputs(3396) <= not a;
    layer1_outputs(3397) <= not (a and b);
    layer1_outputs(3398) <= a and not b;
    layer1_outputs(3399) <= b and not a;
    layer1_outputs(3400) <= '0';
    layer1_outputs(3401) <= not b or a;
    layer1_outputs(3402) <= not b;
    layer1_outputs(3403) <= not b;
    layer1_outputs(3404) <= not a or b;
    layer1_outputs(3405) <= '0';
    layer1_outputs(3406) <= a and not b;
    layer1_outputs(3407) <= not (a and b);
    layer1_outputs(3408) <= not b or a;
    layer1_outputs(3409) <= not a;
    layer1_outputs(3410) <= b;
    layer1_outputs(3411) <= '0';
    layer1_outputs(3412) <= not (a or b);
    layer1_outputs(3413) <= not (a and b);
    layer1_outputs(3414) <= b and not a;
    layer1_outputs(3415) <= not b;
    layer1_outputs(3416) <= a and b;
    layer1_outputs(3417) <= not (a and b);
    layer1_outputs(3418) <= '1';
    layer1_outputs(3419) <= a and b;
    layer1_outputs(3420) <= not a or b;
    layer1_outputs(3421) <= not (a and b);
    layer1_outputs(3422) <= b and not a;
    layer1_outputs(3423) <= '0';
    layer1_outputs(3424) <= a;
    layer1_outputs(3425) <= not (a and b);
    layer1_outputs(3426) <= not (a and b);
    layer1_outputs(3427) <= not a or b;
    layer1_outputs(3428) <= a and not b;
    layer1_outputs(3429) <= not b or a;
    layer1_outputs(3430) <= a and not b;
    layer1_outputs(3431) <= a or b;
    layer1_outputs(3432) <= not b or a;
    layer1_outputs(3433) <= b and not a;
    layer1_outputs(3434) <= not a or b;
    layer1_outputs(3435) <= not b or a;
    layer1_outputs(3436) <= not (a or b);
    layer1_outputs(3437) <= a xor b;
    layer1_outputs(3438) <= a;
    layer1_outputs(3439) <= a and not b;
    layer1_outputs(3440) <= a and b;
    layer1_outputs(3441) <= not a or b;
    layer1_outputs(3442) <= not a;
    layer1_outputs(3443) <= a and not b;
    layer1_outputs(3444) <= b and not a;
    layer1_outputs(3445) <= '1';
    layer1_outputs(3446) <= b and not a;
    layer1_outputs(3447) <= not b or a;
    layer1_outputs(3448) <= a;
    layer1_outputs(3449) <= a;
    layer1_outputs(3450) <= a and b;
    layer1_outputs(3451) <= b;
    layer1_outputs(3452) <= not (a or b);
    layer1_outputs(3453) <= '1';
    layer1_outputs(3454) <= a and b;
    layer1_outputs(3455) <= '1';
    layer1_outputs(3456) <= a and b;
    layer1_outputs(3457) <= not a;
    layer1_outputs(3458) <= '1';
    layer1_outputs(3459) <= '0';
    layer1_outputs(3460) <= b;
    layer1_outputs(3461) <= not (a or b);
    layer1_outputs(3462) <= not b or a;
    layer1_outputs(3463) <= '0';
    layer1_outputs(3464) <= not (a and b);
    layer1_outputs(3465) <= not a or b;
    layer1_outputs(3466) <= '0';
    layer1_outputs(3467) <= not a or b;
    layer1_outputs(3468) <= a or b;
    layer1_outputs(3469) <= not b or a;
    layer1_outputs(3470) <= a xor b;
    layer1_outputs(3471) <= not (a or b);
    layer1_outputs(3472) <= a;
    layer1_outputs(3473) <= '1';
    layer1_outputs(3474) <= a xor b;
    layer1_outputs(3475) <= '0';
    layer1_outputs(3476) <= a and b;
    layer1_outputs(3477) <= a or b;
    layer1_outputs(3478) <= '0';
    layer1_outputs(3479) <= a and b;
    layer1_outputs(3480) <= not b or a;
    layer1_outputs(3481) <= a xor b;
    layer1_outputs(3482) <= '1';
    layer1_outputs(3483) <= a xor b;
    layer1_outputs(3484) <= '0';
    layer1_outputs(3485) <= a or b;
    layer1_outputs(3486) <= not a;
    layer1_outputs(3487) <= not a;
    layer1_outputs(3488) <= not (a or b);
    layer1_outputs(3489) <= a or b;
    layer1_outputs(3490) <= '1';
    layer1_outputs(3491) <= not (a xor b);
    layer1_outputs(3492) <= b and not a;
    layer1_outputs(3493) <= not (a or b);
    layer1_outputs(3494) <= b;
    layer1_outputs(3495) <= '1';
    layer1_outputs(3496) <= not b or a;
    layer1_outputs(3497) <= not (a xor b);
    layer1_outputs(3498) <= a or b;
    layer1_outputs(3499) <= not a or b;
    layer1_outputs(3500) <= b;
    layer1_outputs(3501) <= not (a xor b);
    layer1_outputs(3502) <= b and not a;
    layer1_outputs(3503) <= '1';
    layer1_outputs(3504) <= '1';
    layer1_outputs(3505) <= b;
    layer1_outputs(3506) <= not b;
    layer1_outputs(3507) <= not b;
    layer1_outputs(3508) <= b and not a;
    layer1_outputs(3509) <= not (a xor b);
    layer1_outputs(3510) <= '1';
    layer1_outputs(3511) <= not (a xor b);
    layer1_outputs(3512) <= b;
    layer1_outputs(3513) <= a and b;
    layer1_outputs(3514) <= not b or a;
    layer1_outputs(3515) <= not b or a;
    layer1_outputs(3516) <= '0';
    layer1_outputs(3517) <= b and not a;
    layer1_outputs(3518) <= '0';
    layer1_outputs(3519) <= a and b;
    layer1_outputs(3520) <= '1';
    layer1_outputs(3521) <= '1';
    layer1_outputs(3522) <= not b or a;
    layer1_outputs(3523) <= a xor b;
    layer1_outputs(3524) <= not b or a;
    layer1_outputs(3525) <= a and not b;
    layer1_outputs(3526) <= '0';
    layer1_outputs(3527) <= '1';
    layer1_outputs(3528) <= '1';
    layer1_outputs(3529) <= not a;
    layer1_outputs(3530) <= not a or b;
    layer1_outputs(3531) <= a and b;
    layer1_outputs(3532) <= not (a or b);
    layer1_outputs(3533) <= b;
    layer1_outputs(3534) <= b and not a;
    layer1_outputs(3535) <= not (a or b);
    layer1_outputs(3536) <= not (a xor b);
    layer1_outputs(3537) <= a and b;
    layer1_outputs(3538) <= a and b;
    layer1_outputs(3539) <= '1';
    layer1_outputs(3540) <= a and not b;
    layer1_outputs(3541) <= a and b;
    layer1_outputs(3542) <= a or b;
    layer1_outputs(3543) <= '0';
    layer1_outputs(3544) <= b and not a;
    layer1_outputs(3545) <= not b;
    layer1_outputs(3546) <= '0';
    layer1_outputs(3547) <= a or b;
    layer1_outputs(3548) <= a or b;
    layer1_outputs(3549) <= not (a and b);
    layer1_outputs(3550) <= not a;
    layer1_outputs(3551) <= not b or a;
    layer1_outputs(3552) <= '1';
    layer1_outputs(3553) <= not b;
    layer1_outputs(3554) <= '0';
    layer1_outputs(3555) <= not (a or b);
    layer1_outputs(3556) <= not a;
    layer1_outputs(3557) <= a and b;
    layer1_outputs(3558) <= '0';
    layer1_outputs(3559) <= not (a and b);
    layer1_outputs(3560) <= '1';
    layer1_outputs(3561) <= '0';
    layer1_outputs(3562) <= a or b;
    layer1_outputs(3563) <= a and not b;
    layer1_outputs(3564) <= a;
    layer1_outputs(3565) <= not b or a;
    layer1_outputs(3566) <= '1';
    layer1_outputs(3567) <= not b or a;
    layer1_outputs(3568) <= not b or a;
    layer1_outputs(3569) <= '1';
    layer1_outputs(3570) <= a;
    layer1_outputs(3571) <= a or b;
    layer1_outputs(3572) <= not (a or b);
    layer1_outputs(3573) <= b;
    layer1_outputs(3574) <= '0';
    layer1_outputs(3575) <= not (a and b);
    layer1_outputs(3576) <= '1';
    layer1_outputs(3577) <= not a;
    layer1_outputs(3578) <= b and not a;
    layer1_outputs(3579) <= a;
    layer1_outputs(3580) <= not a or b;
    layer1_outputs(3581) <= not (a or b);
    layer1_outputs(3582) <= '1';
    layer1_outputs(3583) <= not b;
    layer1_outputs(3584) <= not (a and b);
    layer1_outputs(3585) <= not (a and b);
    layer1_outputs(3586) <= a and b;
    layer1_outputs(3587) <= a;
    layer1_outputs(3588) <= a and not b;
    layer1_outputs(3589) <= not b;
    layer1_outputs(3590) <= a and not b;
    layer1_outputs(3591) <= not a;
    layer1_outputs(3592) <= a xor b;
    layer1_outputs(3593) <= not (a xor b);
    layer1_outputs(3594) <= a or b;
    layer1_outputs(3595) <= a and b;
    layer1_outputs(3596) <= '1';
    layer1_outputs(3597) <= not a or b;
    layer1_outputs(3598) <= not (a and b);
    layer1_outputs(3599) <= not b or a;
    layer1_outputs(3600) <= not b or a;
    layer1_outputs(3601) <= b and not a;
    layer1_outputs(3602) <= a and not b;
    layer1_outputs(3603) <= not (a and b);
    layer1_outputs(3604) <= not b;
    layer1_outputs(3605) <= '0';
    layer1_outputs(3606) <= b and not a;
    layer1_outputs(3607) <= not (a and b);
    layer1_outputs(3608) <= not a;
    layer1_outputs(3609) <= a and b;
    layer1_outputs(3610) <= b and not a;
    layer1_outputs(3611) <= not b or a;
    layer1_outputs(3612) <= b and not a;
    layer1_outputs(3613) <= not a or b;
    layer1_outputs(3614) <= not (a and b);
    layer1_outputs(3615) <= not b or a;
    layer1_outputs(3616) <= '1';
    layer1_outputs(3617) <= not a;
    layer1_outputs(3618) <= b;
    layer1_outputs(3619) <= a and b;
    layer1_outputs(3620) <= a and not b;
    layer1_outputs(3621) <= '0';
    layer1_outputs(3622) <= b;
    layer1_outputs(3623) <= not a;
    layer1_outputs(3624) <= '1';
    layer1_outputs(3625) <= not a;
    layer1_outputs(3626) <= a;
    layer1_outputs(3627) <= not a or b;
    layer1_outputs(3628) <= not b;
    layer1_outputs(3629) <= a and not b;
    layer1_outputs(3630) <= a;
    layer1_outputs(3631) <= a and not b;
    layer1_outputs(3632) <= b;
    layer1_outputs(3633) <= a xor b;
    layer1_outputs(3634) <= not a;
    layer1_outputs(3635) <= a and b;
    layer1_outputs(3636) <= b and not a;
    layer1_outputs(3637) <= '1';
    layer1_outputs(3638) <= '0';
    layer1_outputs(3639) <= a and b;
    layer1_outputs(3640) <= b;
    layer1_outputs(3641) <= not b;
    layer1_outputs(3642) <= not (a xor b);
    layer1_outputs(3643) <= '0';
    layer1_outputs(3644) <= '0';
    layer1_outputs(3645) <= a and b;
    layer1_outputs(3646) <= a xor b;
    layer1_outputs(3647) <= not (a and b);
    layer1_outputs(3648) <= not a;
    layer1_outputs(3649) <= a and b;
    layer1_outputs(3650) <= not (a xor b);
    layer1_outputs(3651) <= not (a or b);
    layer1_outputs(3652) <= b;
    layer1_outputs(3653) <= b and not a;
    layer1_outputs(3654) <= a or b;
    layer1_outputs(3655) <= not b or a;
    layer1_outputs(3656) <= '0';
    layer1_outputs(3657) <= '0';
    layer1_outputs(3658) <= b;
    layer1_outputs(3659) <= a;
    layer1_outputs(3660) <= not (a and b);
    layer1_outputs(3661) <= b and not a;
    layer1_outputs(3662) <= a;
    layer1_outputs(3663) <= a or b;
    layer1_outputs(3664) <= not (a and b);
    layer1_outputs(3665) <= not b or a;
    layer1_outputs(3666) <= a or b;
    layer1_outputs(3667) <= a;
    layer1_outputs(3668) <= a and b;
    layer1_outputs(3669) <= '1';
    layer1_outputs(3670) <= a or b;
    layer1_outputs(3671) <= b and not a;
    layer1_outputs(3672) <= not b or a;
    layer1_outputs(3673) <= not a or b;
    layer1_outputs(3674) <= not (a and b);
    layer1_outputs(3675) <= b;
    layer1_outputs(3676) <= '1';
    layer1_outputs(3677) <= not a or b;
    layer1_outputs(3678) <= not a;
    layer1_outputs(3679) <= not (a or b);
    layer1_outputs(3680) <= b;
    layer1_outputs(3681) <= b;
    layer1_outputs(3682) <= b;
    layer1_outputs(3683) <= not a;
    layer1_outputs(3684) <= not (a xor b);
    layer1_outputs(3685) <= not (a and b);
    layer1_outputs(3686) <= not a;
    layer1_outputs(3687) <= '0';
    layer1_outputs(3688) <= not a or b;
    layer1_outputs(3689) <= b and not a;
    layer1_outputs(3690) <= a and not b;
    layer1_outputs(3691) <= b;
    layer1_outputs(3692) <= not a;
    layer1_outputs(3693) <= b;
    layer1_outputs(3694) <= not a;
    layer1_outputs(3695) <= not b or a;
    layer1_outputs(3696) <= '1';
    layer1_outputs(3697) <= not (a or b);
    layer1_outputs(3698) <= not b or a;
    layer1_outputs(3699) <= not (a or b);
    layer1_outputs(3700) <= '1';
    layer1_outputs(3701) <= a or b;
    layer1_outputs(3702) <= not (a and b);
    layer1_outputs(3703) <= '1';
    layer1_outputs(3704) <= '0';
    layer1_outputs(3705) <= '0';
    layer1_outputs(3706) <= not b or a;
    layer1_outputs(3707) <= a and not b;
    layer1_outputs(3708) <= a and b;
    layer1_outputs(3709) <= a or b;
    layer1_outputs(3710) <= not b;
    layer1_outputs(3711) <= not (a and b);
    layer1_outputs(3712) <= a xor b;
    layer1_outputs(3713) <= a and not b;
    layer1_outputs(3714) <= not (a and b);
    layer1_outputs(3715) <= not a;
    layer1_outputs(3716) <= a and b;
    layer1_outputs(3717) <= '1';
    layer1_outputs(3718) <= not a;
    layer1_outputs(3719) <= not a or b;
    layer1_outputs(3720) <= a;
    layer1_outputs(3721) <= '1';
    layer1_outputs(3722) <= not b or a;
    layer1_outputs(3723) <= not (a and b);
    layer1_outputs(3724) <= not (a or b);
    layer1_outputs(3725) <= a;
    layer1_outputs(3726) <= a and b;
    layer1_outputs(3727) <= a and b;
    layer1_outputs(3728) <= a and b;
    layer1_outputs(3729) <= not b;
    layer1_outputs(3730) <= b and not a;
    layer1_outputs(3731) <= not (a and b);
    layer1_outputs(3732) <= b;
    layer1_outputs(3733) <= a or b;
    layer1_outputs(3734) <= '0';
    layer1_outputs(3735) <= '0';
    layer1_outputs(3736) <= not a;
    layer1_outputs(3737) <= b;
    layer1_outputs(3738) <= not (a and b);
    layer1_outputs(3739) <= a;
    layer1_outputs(3740) <= not (a and b);
    layer1_outputs(3741) <= not a or b;
    layer1_outputs(3742) <= a or b;
    layer1_outputs(3743) <= a;
    layer1_outputs(3744) <= not a;
    layer1_outputs(3745) <= not a or b;
    layer1_outputs(3746) <= '1';
    layer1_outputs(3747) <= '0';
    layer1_outputs(3748) <= not a or b;
    layer1_outputs(3749) <= not a;
    layer1_outputs(3750) <= not (a or b);
    layer1_outputs(3751) <= a and b;
    layer1_outputs(3752) <= b and not a;
    layer1_outputs(3753) <= '0';
    layer1_outputs(3754) <= not (a or b);
    layer1_outputs(3755) <= b and not a;
    layer1_outputs(3756) <= a or b;
    layer1_outputs(3757) <= a and not b;
    layer1_outputs(3758) <= a and b;
    layer1_outputs(3759) <= '1';
    layer1_outputs(3760) <= b and not a;
    layer1_outputs(3761) <= not b or a;
    layer1_outputs(3762) <= '1';
    layer1_outputs(3763) <= not b or a;
    layer1_outputs(3764) <= '0';
    layer1_outputs(3765) <= a and not b;
    layer1_outputs(3766) <= not b;
    layer1_outputs(3767) <= not (a or b);
    layer1_outputs(3768) <= '0';
    layer1_outputs(3769) <= '1';
    layer1_outputs(3770) <= a and not b;
    layer1_outputs(3771) <= not (a and b);
    layer1_outputs(3772) <= b and not a;
    layer1_outputs(3773) <= not (a and b);
    layer1_outputs(3774) <= not a or b;
    layer1_outputs(3775) <= '0';
    layer1_outputs(3776) <= b;
    layer1_outputs(3777) <= not (a or b);
    layer1_outputs(3778) <= a or b;
    layer1_outputs(3779) <= a and not b;
    layer1_outputs(3780) <= '0';
    layer1_outputs(3781) <= a;
    layer1_outputs(3782) <= not b or a;
    layer1_outputs(3783) <= a and b;
    layer1_outputs(3784) <= not (a or b);
    layer1_outputs(3785) <= not (a and b);
    layer1_outputs(3786) <= b;
    layer1_outputs(3787) <= not b or a;
    layer1_outputs(3788) <= not a or b;
    layer1_outputs(3789) <= b and not a;
    layer1_outputs(3790) <= '1';
    layer1_outputs(3791) <= not b or a;
    layer1_outputs(3792) <= b and not a;
    layer1_outputs(3793) <= not (a or b);
    layer1_outputs(3794) <= not (a or b);
    layer1_outputs(3795) <= a or b;
    layer1_outputs(3796) <= not b;
    layer1_outputs(3797) <= not (a and b);
    layer1_outputs(3798) <= not b;
    layer1_outputs(3799) <= b;
    layer1_outputs(3800) <= a or b;
    layer1_outputs(3801) <= '0';
    layer1_outputs(3802) <= not (a or b);
    layer1_outputs(3803) <= b;
    layer1_outputs(3804) <= a and not b;
    layer1_outputs(3805) <= not (a and b);
    layer1_outputs(3806) <= a or b;
    layer1_outputs(3807) <= not a or b;
    layer1_outputs(3808) <= not (a or b);
    layer1_outputs(3809) <= '0';
    layer1_outputs(3810) <= a and not b;
    layer1_outputs(3811) <= '1';
    layer1_outputs(3812) <= '1';
    layer1_outputs(3813) <= a;
    layer1_outputs(3814) <= b and not a;
    layer1_outputs(3815) <= a or b;
    layer1_outputs(3816) <= b and not a;
    layer1_outputs(3817) <= '0';
    layer1_outputs(3818) <= b and not a;
    layer1_outputs(3819) <= '1';
    layer1_outputs(3820) <= '0';
    layer1_outputs(3821) <= a or b;
    layer1_outputs(3822) <= '0';
    layer1_outputs(3823) <= a;
    layer1_outputs(3824) <= '0';
    layer1_outputs(3825) <= b;
    layer1_outputs(3826) <= a and b;
    layer1_outputs(3827) <= '1';
    layer1_outputs(3828) <= '0';
    layer1_outputs(3829) <= '0';
    layer1_outputs(3830) <= '0';
    layer1_outputs(3831) <= b;
    layer1_outputs(3832) <= a xor b;
    layer1_outputs(3833) <= b;
    layer1_outputs(3834) <= b and not a;
    layer1_outputs(3835) <= not b or a;
    layer1_outputs(3836) <= a and b;
    layer1_outputs(3837) <= not a;
    layer1_outputs(3838) <= not b;
    layer1_outputs(3839) <= b;
    layer1_outputs(3840) <= '0';
    layer1_outputs(3841) <= a and b;
    layer1_outputs(3842) <= not a or b;
    layer1_outputs(3843) <= not (a and b);
    layer1_outputs(3844) <= a or b;
    layer1_outputs(3845) <= '1';
    layer1_outputs(3846) <= b and not a;
    layer1_outputs(3847) <= not (a and b);
    layer1_outputs(3848) <= not (a and b);
    layer1_outputs(3849) <= '1';
    layer1_outputs(3850) <= not b;
    layer1_outputs(3851) <= not a;
    layer1_outputs(3852) <= not a or b;
    layer1_outputs(3853) <= '1';
    layer1_outputs(3854) <= a or b;
    layer1_outputs(3855) <= not a;
    layer1_outputs(3856) <= not (a and b);
    layer1_outputs(3857) <= not (a and b);
    layer1_outputs(3858) <= a or b;
    layer1_outputs(3859) <= a;
    layer1_outputs(3860) <= not a or b;
    layer1_outputs(3861) <= b;
    layer1_outputs(3862) <= not b or a;
    layer1_outputs(3863) <= '1';
    layer1_outputs(3864) <= a and b;
    layer1_outputs(3865) <= not a;
    layer1_outputs(3866) <= not (a or b);
    layer1_outputs(3867) <= not a or b;
    layer1_outputs(3868) <= '0';
    layer1_outputs(3869) <= '1';
    layer1_outputs(3870) <= a and b;
    layer1_outputs(3871) <= '1';
    layer1_outputs(3872) <= '1';
    layer1_outputs(3873) <= not a;
    layer1_outputs(3874) <= a and b;
    layer1_outputs(3875) <= a or b;
    layer1_outputs(3876) <= not b or a;
    layer1_outputs(3877) <= '0';
    layer1_outputs(3878) <= not a;
    layer1_outputs(3879) <= not b;
    layer1_outputs(3880) <= a and not b;
    layer1_outputs(3881) <= not (a or b);
    layer1_outputs(3882) <= not (a or b);
    layer1_outputs(3883) <= b and not a;
    layer1_outputs(3884) <= not a or b;
    layer1_outputs(3885) <= a;
    layer1_outputs(3886) <= not a;
    layer1_outputs(3887) <= not (a or b);
    layer1_outputs(3888) <= a or b;
    layer1_outputs(3889) <= not a;
    layer1_outputs(3890) <= '0';
    layer1_outputs(3891) <= a or b;
    layer1_outputs(3892) <= b and not a;
    layer1_outputs(3893) <= not (a or b);
    layer1_outputs(3894) <= a or b;
    layer1_outputs(3895) <= not (a and b);
    layer1_outputs(3896) <= not (a or b);
    layer1_outputs(3897) <= a and not b;
    layer1_outputs(3898) <= b;
    layer1_outputs(3899) <= '1';
    layer1_outputs(3900) <= a and b;
    layer1_outputs(3901) <= not (a or b);
    layer1_outputs(3902) <= a and not b;
    layer1_outputs(3903) <= '1';
    layer1_outputs(3904) <= a and not b;
    layer1_outputs(3905) <= not a;
    layer1_outputs(3906) <= not (a or b);
    layer1_outputs(3907) <= a and b;
    layer1_outputs(3908) <= not (a or b);
    layer1_outputs(3909) <= '1';
    layer1_outputs(3910) <= not b or a;
    layer1_outputs(3911) <= b;
    layer1_outputs(3912) <= not b or a;
    layer1_outputs(3913) <= not (a and b);
    layer1_outputs(3914) <= not (a and b);
    layer1_outputs(3915) <= '1';
    layer1_outputs(3916) <= b and not a;
    layer1_outputs(3917) <= b;
    layer1_outputs(3918) <= a and not b;
    layer1_outputs(3919) <= not (a or b);
    layer1_outputs(3920) <= b and not a;
    layer1_outputs(3921) <= '0';
    layer1_outputs(3922) <= '0';
    layer1_outputs(3923) <= not a;
    layer1_outputs(3924) <= not b or a;
    layer1_outputs(3925) <= a and not b;
    layer1_outputs(3926) <= not (a and b);
    layer1_outputs(3927) <= b and not a;
    layer1_outputs(3928) <= a or b;
    layer1_outputs(3929) <= not a;
    layer1_outputs(3930) <= '1';
    layer1_outputs(3931) <= b and not a;
    layer1_outputs(3932) <= a or b;
    layer1_outputs(3933) <= b;
    layer1_outputs(3934) <= not b;
    layer1_outputs(3935) <= a and not b;
    layer1_outputs(3936) <= b;
    layer1_outputs(3937) <= a xor b;
    layer1_outputs(3938) <= not a;
    layer1_outputs(3939) <= b;
    layer1_outputs(3940) <= b;
    layer1_outputs(3941) <= not a or b;
    layer1_outputs(3942) <= b;
    layer1_outputs(3943) <= a and not b;
    layer1_outputs(3944) <= '0';
    layer1_outputs(3945) <= a and b;
    layer1_outputs(3946) <= not a or b;
    layer1_outputs(3947) <= '0';
    layer1_outputs(3948) <= b;
    layer1_outputs(3949) <= b and not a;
    layer1_outputs(3950) <= a;
    layer1_outputs(3951) <= '0';
    layer1_outputs(3952) <= a;
    layer1_outputs(3953) <= not (a and b);
    layer1_outputs(3954) <= b and not a;
    layer1_outputs(3955) <= a and not b;
    layer1_outputs(3956) <= not (a or b);
    layer1_outputs(3957) <= not b;
    layer1_outputs(3958) <= a;
    layer1_outputs(3959) <= not (a and b);
    layer1_outputs(3960) <= not a or b;
    layer1_outputs(3961) <= a or b;
    layer1_outputs(3962) <= b;
    layer1_outputs(3963) <= not a;
    layer1_outputs(3964) <= '0';
    layer1_outputs(3965) <= b;
    layer1_outputs(3966) <= a and not b;
    layer1_outputs(3967) <= '0';
    layer1_outputs(3968) <= '0';
    layer1_outputs(3969) <= '1';
    layer1_outputs(3970) <= a xor b;
    layer1_outputs(3971) <= a and b;
    layer1_outputs(3972) <= not (a and b);
    layer1_outputs(3973) <= a;
    layer1_outputs(3974) <= not a or b;
    layer1_outputs(3975) <= not b or a;
    layer1_outputs(3976) <= '0';
    layer1_outputs(3977) <= b;
    layer1_outputs(3978) <= not b;
    layer1_outputs(3979) <= not b;
    layer1_outputs(3980) <= not b or a;
    layer1_outputs(3981) <= not (a and b);
    layer1_outputs(3982) <= b;
    layer1_outputs(3983) <= a or b;
    layer1_outputs(3984) <= b;
    layer1_outputs(3985) <= '0';
    layer1_outputs(3986) <= not (a or b);
    layer1_outputs(3987) <= not a;
    layer1_outputs(3988) <= not b;
    layer1_outputs(3989) <= not a or b;
    layer1_outputs(3990) <= b;
    layer1_outputs(3991) <= not b or a;
    layer1_outputs(3992) <= '1';
    layer1_outputs(3993) <= not b;
    layer1_outputs(3994) <= not b or a;
    layer1_outputs(3995) <= not b or a;
    layer1_outputs(3996) <= not a or b;
    layer1_outputs(3997) <= not (a and b);
    layer1_outputs(3998) <= a and not b;
    layer1_outputs(3999) <= b and not a;
    layer1_outputs(4000) <= '1';
    layer1_outputs(4001) <= a and b;
    layer1_outputs(4002) <= b;
    layer1_outputs(4003) <= b and not a;
    layer1_outputs(4004) <= a xor b;
    layer1_outputs(4005) <= '0';
    layer1_outputs(4006) <= a and b;
    layer1_outputs(4007) <= a and b;
    layer1_outputs(4008) <= not (a and b);
    layer1_outputs(4009) <= b and not a;
    layer1_outputs(4010) <= not b or a;
    layer1_outputs(4011) <= not b or a;
    layer1_outputs(4012) <= not b or a;
    layer1_outputs(4013) <= not (a or b);
    layer1_outputs(4014) <= a and not b;
    layer1_outputs(4015) <= b;
    layer1_outputs(4016) <= not b or a;
    layer1_outputs(4017) <= b and not a;
    layer1_outputs(4018) <= '0';
    layer1_outputs(4019) <= '1';
    layer1_outputs(4020) <= '0';
    layer1_outputs(4021) <= b and not a;
    layer1_outputs(4022) <= '1';
    layer1_outputs(4023) <= not a;
    layer1_outputs(4024) <= not b;
    layer1_outputs(4025) <= not b or a;
    layer1_outputs(4026) <= '1';
    layer1_outputs(4027) <= '1';
    layer1_outputs(4028) <= '0';
    layer1_outputs(4029) <= b and not a;
    layer1_outputs(4030) <= a;
    layer1_outputs(4031) <= a and not b;
    layer1_outputs(4032) <= a and not b;
    layer1_outputs(4033) <= b;
    layer1_outputs(4034) <= b and not a;
    layer1_outputs(4035) <= '0';
    layer1_outputs(4036) <= not (a or b);
    layer1_outputs(4037) <= b;
    layer1_outputs(4038) <= b;
    layer1_outputs(4039) <= not (a or b);
    layer1_outputs(4040) <= '0';
    layer1_outputs(4041) <= a and not b;
    layer1_outputs(4042) <= not (a and b);
    layer1_outputs(4043) <= not (a or b);
    layer1_outputs(4044) <= not a or b;
    layer1_outputs(4045) <= not (a or b);
    layer1_outputs(4046) <= not b or a;
    layer1_outputs(4047) <= b and not a;
    layer1_outputs(4048) <= '1';
    layer1_outputs(4049) <= a;
    layer1_outputs(4050) <= not (a or b);
    layer1_outputs(4051) <= '0';
    layer1_outputs(4052) <= not b;
    layer1_outputs(4053) <= not (a and b);
    layer1_outputs(4054) <= a or b;
    layer1_outputs(4055) <= '0';
    layer1_outputs(4056) <= not a;
    layer1_outputs(4057) <= not (a and b);
    layer1_outputs(4058) <= '1';
    layer1_outputs(4059) <= '1';
    layer1_outputs(4060) <= a and not b;
    layer1_outputs(4061) <= a xor b;
    layer1_outputs(4062) <= not b;
    layer1_outputs(4063) <= '1';
    layer1_outputs(4064) <= not a;
    layer1_outputs(4065) <= not a;
    layer1_outputs(4066) <= a and b;
    layer1_outputs(4067) <= not (a xor b);
    layer1_outputs(4068) <= a or b;
    layer1_outputs(4069) <= not b;
    layer1_outputs(4070) <= '1';
    layer1_outputs(4071) <= not (a and b);
    layer1_outputs(4072) <= b and not a;
    layer1_outputs(4073) <= '0';
    layer1_outputs(4074) <= a;
    layer1_outputs(4075) <= not (a and b);
    layer1_outputs(4076) <= not a or b;
    layer1_outputs(4077) <= not b or a;
    layer1_outputs(4078) <= not a or b;
    layer1_outputs(4079) <= a and b;
    layer1_outputs(4080) <= '1';
    layer1_outputs(4081) <= not a or b;
    layer1_outputs(4082) <= '1';
    layer1_outputs(4083) <= a and b;
    layer1_outputs(4084) <= a and b;
    layer1_outputs(4085) <= b and not a;
    layer1_outputs(4086) <= '1';
    layer1_outputs(4087) <= a and b;
    layer1_outputs(4088) <= not (a and b);
    layer1_outputs(4089) <= '0';
    layer1_outputs(4090) <= a or b;
    layer1_outputs(4091) <= not b or a;
    layer1_outputs(4092) <= not b or a;
    layer1_outputs(4093) <= '0';
    layer1_outputs(4094) <= a and not b;
    layer1_outputs(4095) <= '0';
    layer1_outputs(4096) <= not b;
    layer1_outputs(4097) <= not (a and b);
    layer1_outputs(4098) <= not (a and b);
    layer1_outputs(4099) <= '0';
    layer1_outputs(4100) <= not b;
    layer1_outputs(4101) <= '1';
    layer1_outputs(4102) <= a or b;
    layer1_outputs(4103) <= not (a and b);
    layer1_outputs(4104) <= not a or b;
    layer1_outputs(4105) <= a and not b;
    layer1_outputs(4106) <= b;
    layer1_outputs(4107) <= not b;
    layer1_outputs(4108) <= not (a and b);
    layer1_outputs(4109) <= not b;
    layer1_outputs(4110) <= not a;
    layer1_outputs(4111) <= a;
    layer1_outputs(4112) <= not a;
    layer1_outputs(4113) <= not (a or b);
    layer1_outputs(4114) <= not b or a;
    layer1_outputs(4115) <= a and not b;
    layer1_outputs(4116) <= b and not a;
    layer1_outputs(4117) <= not (a and b);
    layer1_outputs(4118) <= a or b;
    layer1_outputs(4119) <= not a;
    layer1_outputs(4120) <= a or b;
    layer1_outputs(4121) <= '0';
    layer1_outputs(4122) <= not a or b;
    layer1_outputs(4123) <= a;
    layer1_outputs(4124) <= not b;
    layer1_outputs(4125) <= not b;
    layer1_outputs(4126) <= not b or a;
    layer1_outputs(4127) <= a and not b;
    layer1_outputs(4128) <= not a or b;
    layer1_outputs(4129) <= not (a and b);
    layer1_outputs(4130) <= not (a xor b);
    layer1_outputs(4131) <= not b or a;
    layer1_outputs(4132) <= a and not b;
    layer1_outputs(4133) <= not a or b;
    layer1_outputs(4134) <= b and not a;
    layer1_outputs(4135) <= '1';
    layer1_outputs(4136) <= b;
    layer1_outputs(4137) <= not a;
    layer1_outputs(4138) <= not a or b;
    layer1_outputs(4139) <= a and not b;
    layer1_outputs(4140) <= '0';
    layer1_outputs(4141) <= a;
    layer1_outputs(4142) <= a or b;
    layer1_outputs(4143) <= '0';
    layer1_outputs(4144) <= not b or a;
    layer1_outputs(4145) <= not b;
    layer1_outputs(4146) <= not a or b;
    layer1_outputs(4147) <= a;
    layer1_outputs(4148) <= a or b;
    layer1_outputs(4149) <= not a;
    layer1_outputs(4150) <= not b or a;
    layer1_outputs(4151) <= a and not b;
    layer1_outputs(4152) <= a;
    layer1_outputs(4153) <= not b or a;
    layer1_outputs(4154) <= b;
    layer1_outputs(4155) <= '0';
    layer1_outputs(4156) <= not (a xor b);
    layer1_outputs(4157) <= not (a or b);
    layer1_outputs(4158) <= not b;
    layer1_outputs(4159) <= not a or b;
    layer1_outputs(4160) <= a;
    layer1_outputs(4161) <= a or b;
    layer1_outputs(4162) <= not b;
    layer1_outputs(4163) <= not b or a;
    layer1_outputs(4164) <= a xor b;
    layer1_outputs(4165) <= a;
    layer1_outputs(4166) <= not b;
    layer1_outputs(4167) <= a;
    layer1_outputs(4168) <= not b;
    layer1_outputs(4169) <= a;
    layer1_outputs(4170) <= '0';
    layer1_outputs(4171) <= a or b;
    layer1_outputs(4172) <= b;
    layer1_outputs(4173) <= a and not b;
    layer1_outputs(4174) <= a and not b;
    layer1_outputs(4175) <= b and not a;
    layer1_outputs(4176) <= not b;
    layer1_outputs(4177) <= a;
    layer1_outputs(4178) <= b;
    layer1_outputs(4179) <= a and not b;
    layer1_outputs(4180) <= not a or b;
    layer1_outputs(4181) <= not (a and b);
    layer1_outputs(4182) <= '0';
    layer1_outputs(4183) <= '0';
    layer1_outputs(4184) <= a or b;
    layer1_outputs(4185) <= '0';
    layer1_outputs(4186) <= b;
    layer1_outputs(4187) <= not (a and b);
    layer1_outputs(4188) <= not (a or b);
    layer1_outputs(4189) <= a and not b;
    layer1_outputs(4190) <= b and not a;
    layer1_outputs(4191) <= not a;
    layer1_outputs(4192) <= '1';
    layer1_outputs(4193) <= '0';
    layer1_outputs(4194) <= not a or b;
    layer1_outputs(4195) <= not b or a;
    layer1_outputs(4196) <= not (a and b);
    layer1_outputs(4197) <= a and b;
    layer1_outputs(4198) <= a or b;
    layer1_outputs(4199) <= not b or a;
    layer1_outputs(4200) <= not a or b;
    layer1_outputs(4201) <= a;
    layer1_outputs(4202) <= not a or b;
    layer1_outputs(4203) <= not b;
    layer1_outputs(4204) <= not (a or b);
    layer1_outputs(4205) <= not (a or b);
    layer1_outputs(4206) <= not b;
    layer1_outputs(4207) <= '1';
    layer1_outputs(4208) <= not b or a;
    layer1_outputs(4209) <= b and not a;
    layer1_outputs(4210) <= a and not b;
    layer1_outputs(4211) <= a and not b;
    layer1_outputs(4212) <= a and b;
    layer1_outputs(4213) <= not (a or b);
    layer1_outputs(4214) <= a xor b;
    layer1_outputs(4215) <= not a or b;
    layer1_outputs(4216) <= a or b;
    layer1_outputs(4217) <= not (a and b);
    layer1_outputs(4218) <= b and not a;
    layer1_outputs(4219) <= not (a or b);
    layer1_outputs(4220) <= '1';
    layer1_outputs(4221) <= '0';
    layer1_outputs(4222) <= a or b;
    layer1_outputs(4223) <= not a or b;
    layer1_outputs(4224) <= not (a or b);
    layer1_outputs(4225) <= b;
    layer1_outputs(4226) <= not b;
    layer1_outputs(4227) <= a and b;
    layer1_outputs(4228) <= not a;
    layer1_outputs(4229) <= not b;
    layer1_outputs(4230) <= not a or b;
    layer1_outputs(4231) <= b and not a;
    layer1_outputs(4232) <= not (a and b);
    layer1_outputs(4233) <= not (a and b);
    layer1_outputs(4234) <= not (a and b);
    layer1_outputs(4235) <= a and not b;
    layer1_outputs(4236) <= '0';
    layer1_outputs(4237) <= '1';
    layer1_outputs(4238) <= '0';
    layer1_outputs(4239) <= not b;
    layer1_outputs(4240) <= '0';
    layer1_outputs(4241) <= not a;
    layer1_outputs(4242) <= a;
    layer1_outputs(4243) <= not a or b;
    layer1_outputs(4244) <= not a or b;
    layer1_outputs(4245) <= b and not a;
    layer1_outputs(4246) <= a or b;
    layer1_outputs(4247) <= not b or a;
    layer1_outputs(4248) <= not b or a;
    layer1_outputs(4249) <= not (a xor b);
    layer1_outputs(4250) <= a;
    layer1_outputs(4251) <= a and not b;
    layer1_outputs(4252) <= not b;
    layer1_outputs(4253) <= b;
    layer1_outputs(4254) <= '0';
    layer1_outputs(4255) <= not a;
    layer1_outputs(4256) <= not a;
    layer1_outputs(4257) <= b;
    layer1_outputs(4258) <= not a or b;
    layer1_outputs(4259) <= a and b;
    layer1_outputs(4260) <= a or b;
    layer1_outputs(4261) <= not (a xor b);
    layer1_outputs(4262) <= b and not a;
    layer1_outputs(4263) <= a or b;
    layer1_outputs(4264) <= '0';
    layer1_outputs(4265) <= not b;
    layer1_outputs(4266) <= a or b;
    layer1_outputs(4267) <= a xor b;
    layer1_outputs(4268) <= a and not b;
    layer1_outputs(4269) <= '0';
    layer1_outputs(4270) <= a and b;
    layer1_outputs(4271) <= not b;
    layer1_outputs(4272) <= a;
    layer1_outputs(4273) <= a or b;
    layer1_outputs(4274) <= not b or a;
    layer1_outputs(4275) <= a or b;
    layer1_outputs(4276) <= a and not b;
    layer1_outputs(4277) <= not b or a;
    layer1_outputs(4278) <= a or b;
    layer1_outputs(4279) <= '1';
    layer1_outputs(4280) <= not b;
    layer1_outputs(4281) <= b and not a;
    layer1_outputs(4282) <= not (a or b);
    layer1_outputs(4283) <= b and not a;
    layer1_outputs(4284) <= not a;
    layer1_outputs(4285) <= not b or a;
    layer1_outputs(4286) <= not b;
    layer1_outputs(4287) <= a;
    layer1_outputs(4288) <= '1';
    layer1_outputs(4289) <= not a or b;
    layer1_outputs(4290) <= '1';
    layer1_outputs(4291) <= '1';
    layer1_outputs(4292) <= '0';
    layer1_outputs(4293) <= a or b;
    layer1_outputs(4294) <= not (a and b);
    layer1_outputs(4295) <= '0';
    layer1_outputs(4296) <= '0';
    layer1_outputs(4297) <= not (a or b);
    layer1_outputs(4298) <= a and b;
    layer1_outputs(4299) <= a and b;
    layer1_outputs(4300) <= not b or a;
    layer1_outputs(4301) <= a or b;
    layer1_outputs(4302) <= '1';
    layer1_outputs(4303) <= a and not b;
    layer1_outputs(4304) <= a and b;
    layer1_outputs(4305) <= a and b;
    layer1_outputs(4306) <= a xor b;
    layer1_outputs(4307) <= a xor b;
    layer1_outputs(4308) <= a or b;
    layer1_outputs(4309) <= not (a and b);
    layer1_outputs(4310) <= '0';
    layer1_outputs(4311) <= a;
    layer1_outputs(4312) <= a and not b;
    layer1_outputs(4313) <= not a or b;
    layer1_outputs(4314) <= not (a and b);
    layer1_outputs(4315) <= not (a and b);
    layer1_outputs(4316) <= not (a xor b);
    layer1_outputs(4317) <= '1';
    layer1_outputs(4318) <= b and not a;
    layer1_outputs(4319) <= '1';
    layer1_outputs(4320) <= '1';
    layer1_outputs(4321) <= a and not b;
    layer1_outputs(4322) <= '0';
    layer1_outputs(4323) <= '0';
    layer1_outputs(4324) <= a and b;
    layer1_outputs(4325) <= not (a or b);
    layer1_outputs(4326) <= a;
    layer1_outputs(4327) <= not a or b;
    layer1_outputs(4328) <= b;
    layer1_outputs(4329) <= not b;
    layer1_outputs(4330) <= '0';
    layer1_outputs(4331) <= a xor b;
    layer1_outputs(4332) <= a or b;
    layer1_outputs(4333) <= not b;
    layer1_outputs(4334) <= '0';
    layer1_outputs(4335) <= a and not b;
    layer1_outputs(4336) <= not b;
    layer1_outputs(4337) <= '1';
    layer1_outputs(4338) <= not a;
    layer1_outputs(4339) <= a and not b;
    layer1_outputs(4340) <= b;
    layer1_outputs(4341) <= not a;
    layer1_outputs(4342) <= a xor b;
    layer1_outputs(4343) <= not a;
    layer1_outputs(4344) <= not a;
    layer1_outputs(4345) <= not (a and b);
    layer1_outputs(4346) <= '1';
    layer1_outputs(4347) <= '1';
    layer1_outputs(4348) <= a and b;
    layer1_outputs(4349) <= '1';
    layer1_outputs(4350) <= not (a or b);
    layer1_outputs(4351) <= not a;
    layer1_outputs(4352) <= a and not b;
    layer1_outputs(4353) <= a;
    layer1_outputs(4354) <= not (a and b);
    layer1_outputs(4355) <= not (a and b);
    layer1_outputs(4356) <= not b;
    layer1_outputs(4357) <= '1';
    layer1_outputs(4358) <= not a;
    layer1_outputs(4359) <= a and b;
    layer1_outputs(4360) <= '0';
    layer1_outputs(4361) <= a xor b;
    layer1_outputs(4362) <= '1';
    layer1_outputs(4363) <= a or b;
    layer1_outputs(4364) <= not (a or b);
    layer1_outputs(4365) <= not b or a;
    layer1_outputs(4366) <= b and not a;
    layer1_outputs(4367) <= not a;
    layer1_outputs(4368) <= not (a and b);
    layer1_outputs(4369) <= not b or a;
    layer1_outputs(4370) <= not b;
    layer1_outputs(4371) <= not (a or b);
    layer1_outputs(4372) <= b;
    layer1_outputs(4373) <= not b;
    layer1_outputs(4374) <= a;
    layer1_outputs(4375) <= b;
    layer1_outputs(4376) <= a and b;
    layer1_outputs(4377) <= '0';
    layer1_outputs(4378) <= '0';
    layer1_outputs(4379) <= not a or b;
    layer1_outputs(4380) <= a;
    layer1_outputs(4381) <= not (a or b);
    layer1_outputs(4382) <= '1';
    layer1_outputs(4383) <= b;
    layer1_outputs(4384) <= not b;
    layer1_outputs(4385) <= '0';
    layer1_outputs(4386) <= b and not a;
    layer1_outputs(4387) <= not b;
    layer1_outputs(4388) <= not a or b;
    layer1_outputs(4389) <= a or b;
    layer1_outputs(4390) <= not a or b;
    layer1_outputs(4391) <= a and b;
    layer1_outputs(4392) <= not b or a;
    layer1_outputs(4393) <= not (a or b);
    layer1_outputs(4394) <= a or b;
    layer1_outputs(4395) <= not (a and b);
    layer1_outputs(4396) <= a and b;
    layer1_outputs(4397) <= a;
    layer1_outputs(4398) <= not a or b;
    layer1_outputs(4399) <= b and not a;
    layer1_outputs(4400) <= '1';
    layer1_outputs(4401) <= not (a or b);
    layer1_outputs(4402) <= a;
    layer1_outputs(4403) <= not a or b;
    layer1_outputs(4404) <= not b;
    layer1_outputs(4405) <= b and not a;
    layer1_outputs(4406) <= b and not a;
    layer1_outputs(4407) <= a and b;
    layer1_outputs(4408) <= a;
    layer1_outputs(4409) <= a or b;
    layer1_outputs(4410) <= not (a and b);
    layer1_outputs(4411) <= a xor b;
    layer1_outputs(4412) <= '0';
    layer1_outputs(4413) <= a and not b;
    layer1_outputs(4414) <= not a;
    layer1_outputs(4415) <= a and b;
    layer1_outputs(4416) <= '1';
    layer1_outputs(4417) <= b;
    layer1_outputs(4418) <= a;
    layer1_outputs(4419) <= a and b;
    layer1_outputs(4420) <= not (a or b);
    layer1_outputs(4421) <= not (a and b);
    layer1_outputs(4422) <= not (a or b);
    layer1_outputs(4423) <= a and not b;
    layer1_outputs(4424) <= a;
    layer1_outputs(4425) <= a and b;
    layer1_outputs(4426) <= b;
    layer1_outputs(4427) <= a and b;
    layer1_outputs(4428) <= '1';
    layer1_outputs(4429) <= b;
    layer1_outputs(4430) <= '0';
    layer1_outputs(4431) <= a and b;
    layer1_outputs(4432) <= b;
    layer1_outputs(4433) <= not a;
    layer1_outputs(4434) <= not b;
    layer1_outputs(4435) <= not (a and b);
    layer1_outputs(4436) <= not b or a;
    layer1_outputs(4437) <= not (a or b);
    layer1_outputs(4438) <= a or b;
    layer1_outputs(4439) <= not b or a;
    layer1_outputs(4440) <= not b;
    layer1_outputs(4441) <= not a;
    layer1_outputs(4442) <= '1';
    layer1_outputs(4443) <= a and not b;
    layer1_outputs(4444) <= '0';
    layer1_outputs(4445) <= b and not a;
    layer1_outputs(4446) <= not a or b;
    layer1_outputs(4447) <= not (a and b);
    layer1_outputs(4448) <= not (a or b);
    layer1_outputs(4449) <= a and not b;
    layer1_outputs(4450) <= not (a and b);
    layer1_outputs(4451) <= a;
    layer1_outputs(4452) <= not (a and b);
    layer1_outputs(4453) <= not (a and b);
    layer1_outputs(4454) <= not (a and b);
    layer1_outputs(4455) <= not (a xor b);
    layer1_outputs(4456) <= not (a and b);
    layer1_outputs(4457) <= a and b;
    layer1_outputs(4458) <= not a;
    layer1_outputs(4459) <= b;
    layer1_outputs(4460) <= a or b;
    layer1_outputs(4461) <= b;
    layer1_outputs(4462) <= a and not b;
    layer1_outputs(4463) <= a and not b;
    layer1_outputs(4464) <= a;
    layer1_outputs(4465) <= '0';
    layer1_outputs(4466) <= not b or a;
    layer1_outputs(4467) <= a;
    layer1_outputs(4468) <= a;
    layer1_outputs(4469) <= b;
    layer1_outputs(4470) <= not (a and b);
    layer1_outputs(4471) <= '0';
    layer1_outputs(4472) <= a and b;
    layer1_outputs(4473) <= not (a or b);
    layer1_outputs(4474) <= not (a or b);
    layer1_outputs(4475) <= b and not a;
    layer1_outputs(4476) <= not b;
    layer1_outputs(4477) <= not b;
    layer1_outputs(4478) <= b;
    layer1_outputs(4479) <= b;
    layer1_outputs(4480) <= not a or b;
    layer1_outputs(4481) <= '0';
    layer1_outputs(4482) <= a;
    layer1_outputs(4483) <= a;
    layer1_outputs(4484) <= a;
    layer1_outputs(4485) <= not (a or b);
    layer1_outputs(4486) <= a and b;
    layer1_outputs(4487) <= not (a or b);
    layer1_outputs(4488) <= a or b;
    layer1_outputs(4489) <= a xor b;
    layer1_outputs(4490) <= not b;
    layer1_outputs(4491) <= not (a or b);
    layer1_outputs(4492) <= '1';
    layer1_outputs(4493) <= not a or b;
    layer1_outputs(4494) <= a or b;
    layer1_outputs(4495) <= a;
    layer1_outputs(4496) <= a and b;
    layer1_outputs(4497) <= b;
    layer1_outputs(4498) <= not (a and b);
    layer1_outputs(4499) <= a and b;
    layer1_outputs(4500) <= not a or b;
    layer1_outputs(4501) <= a and b;
    layer1_outputs(4502) <= b and not a;
    layer1_outputs(4503) <= not a or b;
    layer1_outputs(4504) <= '1';
    layer1_outputs(4505) <= not a or b;
    layer1_outputs(4506) <= '1';
    layer1_outputs(4507) <= not b or a;
    layer1_outputs(4508) <= a;
    layer1_outputs(4509) <= not (a and b);
    layer1_outputs(4510) <= a and b;
    layer1_outputs(4511) <= not (a or b);
    layer1_outputs(4512) <= not a;
    layer1_outputs(4513) <= a and not b;
    layer1_outputs(4514) <= not b or a;
    layer1_outputs(4515) <= b and not a;
    layer1_outputs(4516) <= not (a and b);
    layer1_outputs(4517) <= not b or a;
    layer1_outputs(4518) <= '0';
    layer1_outputs(4519) <= not a or b;
    layer1_outputs(4520) <= b;
    layer1_outputs(4521) <= '1';
    layer1_outputs(4522) <= a xor b;
    layer1_outputs(4523) <= a or b;
    layer1_outputs(4524) <= b and not a;
    layer1_outputs(4525) <= b and not a;
    layer1_outputs(4526) <= not (a and b);
    layer1_outputs(4527) <= a xor b;
    layer1_outputs(4528) <= not b or a;
    layer1_outputs(4529) <= a or b;
    layer1_outputs(4530) <= b and not a;
    layer1_outputs(4531) <= a and b;
    layer1_outputs(4532) <= not (a and b);
    layer1_outputs(4533) <= '1';
    layer1_outputs(4534) <= not a;
    layer1_outputs(4535) <= a;
    layer1_outputs(4536) <= a or b;
    layer1_outputs(4537) <= '0';
    layer1_outputs(4538) <= not b or a;
    layer1_outputs(4539) <= '1';
    layer1_outputs(4540) <= not (a or b);
    layer1_outputs(4541) <= a and not b;
    layer1_outputs(4542) <= '0';
    layer1_outputs(4543) <= not b or a;
    layer1_outputs(4544) <= '0';
    layer1_outputs(4545) <= a and b;
    layer1_outputs(4546) <= not a;
    layer1_outputs(4547) <= '0';
    layer1_outputs(4548) <= a and not b;
    layer1_outputs(4549) <= not (a xor b);
    layer1_outputs(4550) <= '0';
    layer1_outputs(4551) <= not (a or b);
    layer1_outputs(4552) <= not (a xor b);
    layer1_outputs(4553) <= a or b;
    layer1_outputs(4554) <= b;
    layer1_outputs(4555) <= a or b;
    layer1_outputs(4556) <= not (a or b);
    layer1_outputs(4557) <= not (a xor b);
    layer1_outputs(4558) <= b and not a;
    layer1_outputs(4559) <= not (a and b);
    layer1_outputs(4560) <= a and not b;
    layer1_outputs(4561) <= a;
    layer1_outputs(4562) <= a or b;
    layer1_outputs(4563) <= a and b;
    layer1_outputs(4564) <= '0';
    layer1_outputs(4565) <= '0';
    layer1_outputs(4566) <= a and not b;
    layer1_outputs(4567) <= not b or a;
    layer1_outputs(4568) <= not a;
    layer1_outputs(4569) <= not b or a;
    layer1_outputs(4570) <= b;
    layer1_outputs(4571) <= a xor b;
    layer1_outputs(4572) <= '1';
    layer1_outputs(4573) <= not a or b;
    layer1_outputs(4574) <= a and b;
    layer1_outputs(4575) <= not a or b;
    layer1_outputs(4576) <= a or b;
    layer1_outputs(4577) <= not a;
    layer1_outputs(4578) <= a or b;
    layer1_outputs(4579) <= '0';
    layer1_outputs(4580) <= '0';
    layer1_outputs(4581) <= not (a and b);
    layer1_outputs(4582) <= not a or b;
    layer1_outputs(4583) <= not b or a;
    layer1_outputs(4584) <= a and b;
    layer1_outputs(4585) <= b;
    layer1_outputs(4586) <= a and not b;
    layer1_outputs(4587) <= a and not b;
    layer1_outputs(4588) <= not (a or b);
    layer1_outputs(4589) <= '1';
    layer1_outputs(4590) <= a;
    layer1_outputs(4591) <= not (a or b);
    layer1_outputs(4592) <= a;
    layer1_outputs(4593) <= '0';
    layer1_outputs(4594) <= not (a and b);
    layer1_outputs(4595) <= not (a or b);
    layer1_outputs(4596) <= b;
    layer1_outputs(4597) <= not (a xor b);
    layer1_outputs(4598) <= not a or b;
    layer1_outputs(4599) <= a;
    layer1_outputs(4600) <= a and not b;
    layer1_outputs(4601) <= not a or b;
    layer1_outputs(4602) <= a;
    layer1_outputs(4603) <= not b;
    layer1_outputs(4604) <= not b;
    layer1_outputs(4605) <= not (a or b);
    layer1_outputs(4606) <= a xor b;
    layer1_outputs(4607) <= '0';
    layer1_outputs(4608) <= not a;
    layer1_outputs(4609) <= a and not b;
    layer1_outputs(4610) <= not b or a;
    layer1_outputs(4611) <= not (a xor b);
    layer1_outputs(4612) <= a;
    layer1_outputs(4613) <= not b or a;
    layer1_outputs(4614) <= '0';
    layer1_outputs(4615) <= b;
    layer1_outputs(4616) <= not b;
    layer1_outputs(4617) <= b and not a;
    layer1_outputs(4618) <= '1';
    layer1_outputs(4619) <= a and not b;
    layer1_outputs(4620) <= a and not b;
    layer1_outputs(4621) <= not b;
    layer1_outputs(4622) <= b;
    layer1_outputs(4623) <= a and b;
    layer1_outputs(4624) <= b;
    layer1_outputs(4625) <= '1';
    layer1_outputs(4626) <= not (a or b);
    layer1_outputs(4627) <= not b or a;
    layer1_outputs(4628) <= a and b;
    layer1_outputs(4629) <= not a;
    layer1_outputs(4630) <= a xor b;
    layer1_outputs(4631) <= a and not b;
    layer1_outputs(4632) <= not b;
    layer1_outputs(4633) <= not b;
    layer1_outputs(4634) <= a and b;
    layer1_outputs(4635) <= not (a or b);
    layer1_outputs(4636) <= '1';
    layer1_outputs(4637) <= a;
    layer1_outputs(4638) <= b and not a;
    layer1_outputs(4639) <= a and not b;
    layer1_outputs(4640) <= not a;
    layer1_outputs(4641) <= not b or a;
    layer1_outputs(4642) <= b and not a;
    layer1_outputs(4643) <= '1';
    layer1_outputs(4644) <= not b;
    layer1_outputs(4645) <= a;
    layer1_outputs(4646) <= not b;
    layer1_outputs(4647) <= not a;
    layer1_outputs(4648) <= not b;
    layer1_outputs(4649) <= not a or b;
    layer1_outputs(4650) <= '0';
    layer1_outputs(4651) <= '1';
    layer1_outputs(4652) <= b and not a;
    layer1_outputs(4653) <= not a;
    layer1_outputs(4654) <= a and b;
    layer1_outputs(4655) <= a and not b;
    layer1_outputs(4656) <= not b;
    layer1_outputs(4657) <= '0';
    layer1_outputs(4658) <= '0';
    layer1_outputs(4659) <= not (a and b);
    layer1_outputs(4660) <= a and b;
    layer1_outputs(4661) <= '1';
    layer1_outputs(4662) <= '1';
    layer1_outputs(4663) <= not (a and b);
    layer1_outputs(4664) <= not b or a;
    layer1_outputs(4665) <= a and b;
    layer1_outputs(4666) <= not b;
    layer1_outputs(4667) <= not (a xor b);
    layer1_outputs(4668) <= a or b;
    layer1_outputs(4669) <= b and not a;
    layer1_outputs(4670) <= b and not a;
    layer1_outputs(4671) <= '1';
    layer1_outputs(4672) <= a and b;
    layer1_outputs(4673) <= b and not a;
    layer1_outputs(4674) <= a and not b;
    layer1_outputs(4675) <= a or b;
    layer1_outputs(4676) <= a or b;
    layer1_outputs(4677) <= '0';
    layer1_outputs(4678) <= not b;
    layer1_outputs(4679) <= a xor b;
    layer1_outputs(4680) <= not b or a;
    layer1_outputs(4681) <= not b;
    layer1_outputs(4682) <= b and not a;
    layer1_outputs(4683) <= '1';
    layer1_outputs(4684) <= not a or b;
    layer1_outputs(4685) <= a or b;
    layer1_outputs(4686) <= not b or a;
    layer1_outputs(4687) <= a or b;
    layer1_outputs(4688) <= '1';
    layer1_outputs(4689) <= '1';
    layer1_outputs(4690) <= not a or b;
    layer1_outputs(4691) <= '0';
    layer1_outputs(4692) <= a xor b;
    layer1_outputs(4693) <= a;
    layer1_outputs(4694) <= a and b;
    layer1_outputs(4695) <= '0';
    layer1_outputs(4696) <= b and not a;
    layer1_outputs(4697) <= '0';
    layer1_outputs(4698) <= '1';
    layer1_outputs(4699) <= b;
    layer1_outputs(4700) <= '0';
    layer1_outputs(4701) <= '1';
    layer1_outputs(4702) <= a and not b;
    layer1_outputs(4703) <= not b or a;
    layer1_outputs(4704) <= not b;
    layer1_outputs(4705) <= not a or b;
    layer1_outputs(4706) <= b and not a;
    layer1_outputs(4707) <= '0';
    layer1_outputs(4708) <= a or b;
    layer1_outputs(4709) <= b and not a;
    layer1_outputs(4710) <= not (a or b);
    layer1_outputs(4711) <= not b or a;
    layer1_outputs(4712) <= '0';
    layer1_outputs(4713) <= a xor b;
    layer1_outputs(4714) <= b;
    layer1_outputs(4715) <= not b;
    layer1_outputs(4716) <= a;
    layer1_outputs(4717) <= not a or b;
    layer1_outputs(4718) <= not (a or b);
    layer1_outputs(4719) <= a or b;
    layer1_outputs(4720) <= b and not a;
    layer1_outputs(4721) <= a and not b;
    layer1_outputs(4722) <= not a;
    layer1_outputs(4723) <= a and not b;
    layer1_outputs(4724) <= not (a or b);
    layer1_outputs(4725) <= a and not b;
    layer1_outputs(4726) <= a or b;
    layer1_outputs(4727) <= not (a and b);
    layer1_outputs(4728) <= not a or b;
    layer1_outputs(4729) <= '1';
    layer1_outputs(4730) <= a and b;
    layer1_outputs(4731) <= a;
    layer1_outputs(4732) <= '0';
    layer1_outputs(4733) <= not b;
    layer1_outputs(4734) <= not b;
    layer1_outputs(4735) <= not a or b;
    layer1_outputs(4736) <= not b;
    layer1_outputs(4737) <= not (a or b);
    layer1_outputs(4738) <= '0';
    layer1_outputs(4739) <= not (a and b);
    layer1_outputs(4740) <= not b or a;
    layer1_outputs(4741) <= '1';
    layer1_outputs(4742) <= not (a or b);
    layer1_outputs(4743) <= a;
    layer1_outputs(4744) <= not b or a;
    layer1_outputs(4745) <= '0';
    layer1_outputs(4746) <= not b or a;
    layer1_outputs(4747) <= '0';
    layer1_outputs(4748) <= not a;
    layer1_outputs(4749) <= not (a and b);
    layer1_outputs(4750) <= a;
    layer1_outputs(4751) <= a or b;
    layer1_outputs(4752) <= not (a xor b);
    layer1_outputs(4753) <= b and not a;
    layer1_outputs(4754) <= not (a or b);
    layer1_outputs(4755) <= not a or b;
    layer1_outputs(4756) <= not (a and b);
    layer1_outputs(4757) <= '1';
    layer1_outputs(4758) <= not a;
    layer1_outputs(4759) <= '0';
    layer1_outputs(4760) <= not (a and b);
    layer1_outputs(4761) <= a and not b;
    layer1_outputs(4762) <= not (a and b);
    layer1_outputs(4763) <= a and b;
    layer1_outputs(4764) <= a xor b;
    layer1_outputs(4765) <= '0';
    layer1_outputs(4766) <= not (a or b);
    layer1_outputs(4767) <= a and not b;
    layer1_outputs(4768) <= a or b;
    layer1_outputs(4769) <= a or b;
    layer1_outputs(4770) <= not (a xor b);
    layer1_outputs(4771) <= b and not a;
    layer1_outputs(4772) <= a and not b;
    layer1_outputs(4773) <= a xor b;
    layer1_outputs(4774) <= not (a xor b);
    layer1_outputs(4775) <= not (a and b);
    layer1_outputs(4776) <= not b or a;
    layer1_outputs(4777) <= '1';
    layer1_outputs(4778) <= a and b;
    layer1_outputs(4779) <= '0';
    layer1_outputs(4780) <= '1';
    layer1_outputs(4781) <= not a;
    layer1_outputs(4782) <= '0';
    layer1_outputs(4783) <= a and b;
    layer1_outputs(4784) <= a;
    layer1_outputs(4785) <= a;
    layer1_outputs(4786) <= '1';
    layer1_outputs(4787) <= '1';
    layer1_outputs(4788) <= '0';
    layer1_outputs(4789) <= not (a or b);
    layer1_outputs(4790) <= not (a and b);
    layer1_outputs(4791) <= a or b;
    layer1_outputs(4792) <= a and b;
    layer1_outputs(4793) <= a or b;
    layer1_outputs(4794) <= not b or a;
    layer1_outputs(4795) <= not a;
    layer1_outputs(4796) <= b and not a;
    layer1_outputs(4797) <= b and not a;
    layer1_outputs(4798) <= a and b;
    layer1_outputs(4799) <= not (a and b);
    layer1_outputs(4800) <= b;
    layer1_outputs(4801) <= '0';
    layer1_outputs(4802) <= b and not a;
    layer1_outputs(4803) <= a and b;
    layer1_outputs(4804) <= a and b;
    layer1_outputs(4805) <= not b;
    layer1_outputs(4806) <= '1';
    layer1_outputs(4807) <= a and not b;
    layer1_outputs(4808) <= not a or b;
    layer1_outputs(4809) <= not (a and b);
    layer1_outputs(4810) <= not (a xor b);
    layer1_outputs(4811) <= not (a and b);
    layer1_outputs(4812) <= b;
    layer1_outputs(4813) <= '0';
    layer1_outputs(4814) <= not (a and b);
    layer1_outputs(4815) <= not (a and b);
    layer1_outputs(4816) <= not b or a;
    layer1_outputs(4817) <= '1';
    layer1_outputs(4818) <= b;
    layer1_outputs(4819) <= b and not a;
    layer1_outputs(4820) <= not a;
    layer1_outputs(4821) <= not (a or b);
    layer1_outputs(4822) <= '0';
    layer1_outputs(4823) <= '1';
    layer1_outputs(4824) <= not a;
    layer1_outputs(4825) <= not (a or b);
    layer1_outputs(4826) <= '0';
    layer1_outputs(4827) <= '0';
    layer1_outputs(4828) <= not (a and b);
    layer1_outputs(4829) <= b and not a;
    layer1_outputs(4830) <= '0';
    layer1_outputs(4831) <= b;
    layer1_outputs(4832) <= a and not b;
    layer1_outputs(4833) <= '1';
    layer1_outputs(4834) <= '1';
    layer1_outputs(4835) <= not b;
    layer1_outputs(4836) <= '1';
    layer1_outputs(4837) <= a or b;
    layer1_outputs(4838) <= '1';
    layer1_outputs(4839) <= a and b;
    layer1_outputs(4840) <= a or b;
    layer1_outputs(4841) <= a;
    layer1_outputs(4842) <= a and b;
    layer1_outputs(4843) <= '1';
    layer1_outputs(4844) <= not (a and b);
    layer1_outputs(4845) <= a and not b;
    layer1_outputs(4846) <= b and not a;
    layer1_outputs(4847) <= a;
    layer1_outputs(4848) <= not b;
    layer1_outputs(4849) <= a and b;
    layer1_outputs(4850) <= not a or b;
    layer1_outputs(4851) <= a and not b;
    layer1_outputs(4852) <= b;
    layer1_outputs(4853) <= b and not a;
    layer1_outputs(4854) <= '1';
    layer1_outputs(4855) <= a and not b;
    layer1_outputs(4856) <= '0';
    layer1_outputs(4857) <= not (a or b);
    layer1_outputs(4858) <= a and b;
    layer1_outputs(4859) <= a or b;
    layer1_outputs(4860) <= a;
    layer1_outputs(4861) <= b;
    layer1_outputs(4862) <= b and not a;
    layer1_outputs(4863) <= a and not b;
    layer1_outputs(4864) <= '0';
    layer1_outputs(4865) <= not b or a;
    layer1_outputs(4866) <= a;
    layer1_outputs(4867) <= not a;
    layer1_outputs(4868) <= '1';
    layer1_outputs(4869) <= a;
    layer1_outputs(4870) <= a and not b;
    layer1_outputs(4871) <= not b or a;
    layer1_outputs(4872) <= a and not b;
    layer1_outputs(4873) <= not b or a;
    layer1_outputs(4874) <= a;
    layer1_outputs(4875) <= a and not b;
    layer1_outputs(4876) <= not b or a;
    layer1_outputs(4877) <= a and not b;
    layer1_outputs(4878) <= not a or b;
    layer1_outputs(4879) <= b;
    layer1_outputs(4880) <= not a or b;
    layer1_outputs(4881) <= not (a or b);
    layer1_outputs(4882) <= not (a or b);
    layer1_outputs(4883) <= not a or b;
    layer1_outputs(4884) <= not (a xor b);
    layer1_outputs(4885) <= not (a and b);
    layer1_outputs(4886) <= not (a and b);
    layer1_outputs(4887) <= a and b;
    layer1_outputs(4888) <= not b or a;
    layer1_outputs(4889) <= b and not a;
    layer1_outputs(4890) <= not (a xor b);
    layer1_outputs(4891) <= '1';
    layer1_outputs(4892) <= a and not b;
    layer1_outputs(4893) <= a;
    layer1_outputs(4894) <= not b or a;
    layer1_outputs(4895) <= a xor b;
    layer1_outputs(4896) <= a and b;
    layer1_outputs(4897) <= not (a or b);
    layer1_outputs(4898) <= '1';
    layer1_outputs(4899) <= a;
    layer1_outputs(4900) <= '0';
    layer1_outputs(4901) <= a;
    layer1_outputs(4902) <= '1';
    layer1_outputs(4903) <= not b or a;
    layer1_outputs(4904) <= a or b;
    layer1_outputs(4905) <= b and not a;
    layer1_outputs(4906) <= a;
    layer1_outputs(4907) <= a xor b;
    layer1_outputs(4908) <= '0';
    layer1_outputs(4909) <= '0';
    layer1_outputs(4910) <= not a or b;
    layer1_outputs(4911) <= '0';
    layer1_outputs(4912) <= not a;
    layer1_outputs(4913) <= not (a and b);
    layer1_outputs(4914) <= '0';
    layer1_outputs(4915) <= a and not b;
    layer1_outputs(4916) <= b and not a;
    layer1_outputs(4917) <= a and b;
    layer1_outputs(4918) <= '1';
    layer1_outputs(4919) <= '1';
    layer1_outputs(4920) <= not a;
    layer1_outputs(4921) <= not (a and b);
    layer1_outputs(4922) <= b and not a;
    layer1_outputs(4923) <= '0';
    layer1_outputs(4924) <= a and not b;
    layer1_outputs(4925) <= not b;
    layer1_outputs(4926) <= a and b;
    layer1_outputs(4927) <= b;
    layer1_outputs(4928) <= '0';
    layer1_outputs(4929) <= '1';
    layer1_outputs(4930) <= b and not a;
    layer1_outputs(4931) <= not a;
    layer1_outputs(4932) <= a and b;
    layer1_outputs(4933) <= a and not b;
    layer1_outputs(4934) <= not b or a;
    layer1_outputs(4935) <= not a or b;
    layer1_outputs(4936) <= a xor b;
    layer1_outputs(4937) <= not (a or b);
    layer1_outputs(4938) <= '1';
    layer1_outputs(4939) <= not b or a;
    layer1_outputs(4940) <= a;
    layer1_outputs(4941) <= not a or b;
    layer1_outputs(4942) <= '1';
    layer1_outputs(4943) <= not a or b;
    layer1_outputs(4944) <= not b;
    layer1_outputs(4945) <= '1';
    layer1_outputs(4946) <= not (a or b);
    layer1_outputs(4947) <= a and b;
    layer1_outputs(4948) <= '1';
    layer1_outputs(4949) <= not a;
    layer1_outputs(4950) <= a and not b;
    layer1_outputs(4951) <= b;
    layer1_outputs(4952) <= not (a xor b);
    layer1_outputs(4953) <= a and not b;
    layer1_outputs(4954) <= not a;
    layer1_outputs(4955) <= not (a and b);
    layer1_outputs(4956) <= '1';
    layer1_outputs(4957) <= '0';
    layer1_outputs(4958) <= b;
    layer1_outputs(4959) <= not a or b;
    layer1_outputs(4960) <= a and not b;
    layer1_outputs(4961) <= a and not b;
    layer1_outputs(4962) <= not a or b;
    layer1_outputs(4963) <= not a or b;
    layer1_outputs(4964) <= not a or b;
    layer1_outputs(4965) <= b and not a;
    layer1_outputs(4966) <= a;
    layer1_outputs(4967) <= b;
    layer1_outputs(4968) <= b and not a;
    layer1_outputs(4969) <= not a or b;
    layer1_outputs(4970) <= not b;
    layer1_outputs(4971) <= a;
    layer1_outputs(4972) <= not b;
    layer1_outputs(4973) <= '1';
    layer1_outputs(4974) <= b and not a;
    layer1_outputs(4975) <= '0';
    layer1_outputs(4976) <= not (a or b);
    layer1_outputs(4977) <= a and not b;
    layer1_outputs(4978) <= a and not b;
    layer1_outputs(4979) <= a and b;
    layer1_outputs(4980) <= not b or a;
    layer1_outputs(4981) <= '1';
    layer1_outputs(4982) <= a or b;
    layer1_outputs(4983) <= not (a or b);
    layer1_outputs(4984) <= a and b;
    layer1_outputs(4985) <= '0';
    layer1_outputs(4986) <= b;
    layer1_outputs(4987) <= a and not b;
    layer1_outputs(4988) <= a and not b;
    layer1_outputs(4989) <= b and not a;
    layer1_outputs(4990) <= not (a or b);
    layer1_outputs(4991) <= a;
    layer1_outputs(4992) <= a or b;
    layer1_outputs(4993) <= not a or b;
    layer1_outputs(4994) <= a and b;
    layer1_outputs(4995) <= a and not b;
    layer1_outputs(4996) <= not b;
    layer1_outputs(4997) <= b;
    layer1_outputs(4998) <= a;
    layer1_outputs(4999) <= '1';
    layer1_outputs(5000) <= not (a xor b);
    layer1_outputs(5001) <= not b or a;
    layer1_outputs(5002) <= '0';
    layer1_outputs(5003) <= b and not a;
    layer1_outputs(5004) <= a and b;
    layer1_outputs(5005) <= b and not a;
    layer1_outputs(5006) <= not (a or b);
    layer1_outputs(5007) <= '0';
    layer1_outputs(5008) <= a;
    layer1_outputs(5009) <= not b;
    layer1_outputs(5010) <= a and not b;
    layer1_outputs(5011) <= not b or a;
    layer1_outputs(5012) <= a;
    layer1_outputs(5013) <= not (a xor b);
    layer1_outputs(5014) <= a and b;
    layer1_outputs(5015) <= a and not b;
    layer1_outputs(5016) <= a and not b;
    layer1_outputs(5017) <= not b;
    layer1_outputs(5018) <= '1';
    layer1_outputs(5019) <= not a or b;
    layer1_outputs(5020) <= a or b;
    layer1_outputs(5021) <= not b or a;
    layer1_outputs(5022) <= '0';
    layer1_outputs(5023) <= '1';
    layer1_outputs(5024) <= b and not a;
    layer1_outputs(5025) <= '1';
    layer1_outputs(5026) <= a xor b;
    layer1_outputs(5027) <= b and not a;
    layer1_outputs(5028) <= '0';
    layer1_outputs(5029) <= not a or b;
    layer1_outputs(5030) <= a and b;
    layer1_outputs(5031) <= '1';
    layer1_outputs(5032) <= not a;
    layer1_outputs(5033) <= not (a and b);
    layer1_outputs(5034) <= '0';
    layer1_outputs(5035) <= not a or b;
    layer1_outputs(5036) <= a;
    layer1_outputs(5037) <= a or b;
    layer1_outputs(5038) <= b;
    layer1_outputs(5039) <= a;
    layer1_outputs(5040) <= not (a and b);
    layer1_outputs(5041) <= '1';
    layer1_outputs(5042) <= not b or a;
    layer1_outputs(5043) <= not a;
    layer1_outputs(5044) <= not (a or b);
    layer1_outputs(5045) <= not a;
    layer1_outputs(5046) <= not a;
    layer1_outputs(5047) <= not b;
    layer1_outputs(5048) <= not (a and b);
    layer1_outputs(5049) <= a;
    layer1_outputs(5050) <= b;
    layer1_outputs(5051) <= not (a and b);
    layer1_outputs(5052) <= '1';
    layer1_outputs(5053) <= '0';
    layer1_outputs(5054) <= not b;
    layer1_outputs(5055) <= not a;
    layer1_outputs(5056) <= a and not b;
    layer1_outputs(5057) <= b;
    layer1_outputs(5058) <= a and not b;
    layer1_outputs(5059) <= a and b;
    layer1_outputs(5060) <= not (a and b);
    layer1_outputs(5061) <= not (a and b);
    layer1_outputs(5062) <= not a or b;
    layer1_outputs(5063) <= b;
    layer1_outputs(5064) <= a and not b;
    layer1_outputs(5065) <= b;
    layer1_outputs(5066) <= not (a or b);
    layer1_outputs(5067) <= b;
    layer1_outputs(5068) <= not (a and b);
    layer1_outputs(5069) <= not (a or b);
    layer1_outputs(5070) <= a and b;
    layer1_outputs(5071) <= a or b;
    layer1_outputs(5072) <= b;
    layer1_outputs(5073) <= not a or b;
    layer1_outputs(5074) <= not b or a;
    layer1_outputs(5075) <= '1';
    layer1_outputs(5076) <= a;
    layer1_outputs(5077) <= b;
    layer1_outputs(5078) <= not a or b;
    layer1_outputs(5079) <= '1';
    layer1_outputs(5080) <= not a;
    layer1_outputs(5081) <= a or b;
    layer1_outputs(5082) <= not a or b;
    layer1_outputs(5083) <= '0';
    layer1_outputs(5084) <= b;
    layer1_outputs(5085) <= not a or b;
    layer1_outputs(5086) <= '1';
    layer1_outputs(5087) <= '1';
    layer1_outputs(5088) <= not (a and b);
    layer1_outputs(5089) <= a and b;
    layer1_outputs(5090) <= not (a or b);
    layer1_outputs(5091) <= b and not a;
    layer1_outputs(5092) <= not a or b;
    layer1_outputs(5093) <= '0';
    layer1_outputs(5094) <= not (a and b);
    layer1_outputs(5095) <= not b;
    layer1_outputs(5096) <= a;
    layer1_outputs(5097) <= not a;
    layer1_outputs(5098) <= a and b;
    layer1_outputs(5099) <= '0';
    layer1_outputs(5100) <= b and not a;
    layer1_outputs(5101) <= not (a xor b);
    layer1_outputs(5102) <= b;
    layer1_outputs(5103) <= not a;
    layer1_outputs(5104) <= not b or a;
    layer1_outputs(5105) <= b and not a;
    layer1_outputs(5106) <= not a;
    layer1_outputs(5107) <= not (a or b);
    layer1_outputs(5108) <= a;
    layer1_outputs(5109) <= not b or a;
    layer1_outputs(5110) <= not a or b;
    layer1_outputs(5111) <= a and not b;
    layer1_outputs(5112) <= '0';
    layer1_outputs(5113) <= not (a and b);
    layer1_outputs(5114) <= a and b;
    layer1_outputs(5115) <= a;
    layer1_outputs(5116) <= not a;
    layer1_outputs(5117) <= a and b;
    layer1_outputs(5118) <= a and b;
    layer1_outputs(5119) <= not a or b;
    layer2_outputs(0) <= a;
    layer2_outputs(1) <= a or b;
    layer2_outputs(2) <= a and not b;
    layer2_outputs(3) <= a or b;
    layer2_outputs(4) <= not b;
    layer2_outputs(5) <= a and not b;
    layer2_outputs(6) <= a and not b;
    layer2_outputs(7) <= a and not b;
    layer2_outputs(8) <= a or b;
    layer2_outputs(9) <= not (a and b);
    layer2_outputs(10) <= a;
    layer2_outputs(11) <= not (a or b);
    layer2_outputs(12) <= a and not b;
    layer2_outputs(13) <= a or b;
    layer2_outputs(14) <= not a or b;
    layer2_outputs(15) <= not (a and b);
    layer2_outputs(16) <= a and not b;
    layer2_outputs(17) <= not a or b;
    layer2_outputs(18) <= not b or a;
    layer2_outputs(19) <= '0';
    layer2_outputs(20) <= not (a and b);
    layer2_outputs(21) <= b and not a;
    layer2_outputs(22) <= not (a and b);
    layer2_outputs(23) <= not a or b;
    layer2_outputs(24) <= a or b;
    layer2_outputs(25) <= '0';
    layer2_outputs(26) <= not (a xor b);
    layer2_outputs(27) <= a and not b;
    layer2_outputs(28) <= not b or a;
    layer2_outputs(29) <= '0';
    layer2_outputs(30) <= b and not a;
    layer2_outputs(31) <= '1';
    layer2_outputs(32) <= not b or a;
    layer2_outputs(33) <= a and not b;
    layer2_outputs(34) <= not (a and b);
    layer2_outputs(35) <= a or b;
    layer2_outputs(36) <= not b or a;
    layer2_outputs(37) <= a and not b;
    layer2_outputs(38) <= '0';
    layer2_outputs(39) <= '0';
    layer2_outputs(40) <= not b or a;
    layer2_outputs(41) <= a and not b;
    layer2_outputs(42) <= not a;
    layer2_outputs(43) <= '0';
    layer2_outputs(44) <= a;
    layer2_outputs(45) <= not (a and b);
    layer2_outputs(46) <= '0';
    layer2_outputs(47) <= '0';
    layer2_outputs(48) <= a or b;
    layer2_outputs(49) <= not a or b;
    layer2_outputs(50) <= not b or a;
    layer2_outputs(51) <= '0';
    layer2_outputs(52) <= b and not a;
    layer2_outputs(53) <= a;
    layer2_outputs(54) <= a;
    layer2_outputs(55) <= not (a and b);
    layer2_outputs(56) <= a and b;
    layer2_outputs(57) <= b and not a;
    layer2_outputs(58) <= not b;
    layer2_outputs(59) <= not (a or b);
    layer2_outputs(60) <= a and b;
    layer2_outputs(61) <= '0';
    layer2_outputs(62) <= '1';
    layer2_outputs(63) <= not a;
    layer2_outputs(64) <= not a or b;
    layer2_outputs(65) <= not a or b;
    layer2_outputs(66) <= not (a and b);
    layer2_outputs(67) <= not (a or b);
    layer2_outputs(68) <= a or b;
    layer2_outputs(69) <= not b or a;
    layer2_outputs(70) <= a;
    layer2_outputs(71) <= a or b;
    layer2_outputs(72) <= not a;
    layer2_outputs(73) <= not b or a;
    layer2_outputs(74) <= '1';
    layer2_outputs(75) <= '1';
    layer2_outputs(76) <= not b;
    layer2_outputs(77) <= b;
    layer2_outputs(78) <= not a or b;
    layer2_outputs(79) <= '1';
    layer2_outputs(80) <= not (a xor b);
    layer2_outputs(81) <= not a or b;
    layer2_outputs(82) <= '0';
    layer2_outputs(83) <= '1';
    layer2_outputs(84) <= b and not a;
    layer2_outputs(85) <= a;
    layer2_outputs(86) <= not (a and b);
    layer2_outputs(87) <= not b;
    layer2_outputs(88) <= '1';
    layer2_outputs(89) <= a and not b;
    layer2_outputs(90) <= not b;
    layer2_outputs(91) <= a;
    layer2_outputs(92) <= a and b;
    layer2_outputs(93) <= not b;
    layer2_outputs(94) <= a and not b;
    layer2_outputs(95) <= b;
    layer2_outputs(96) <= '0';
    layer2_outputs(97) <= not b or a;
    layer2_outputs(98) <= not a;
    layer2_outputs(99) <= '1';
    layer2_outputs(100) <= not (a and b);
    layer2_outputs(101) <= not (a and b);
    layer2_outputs(102) <= a;
    layer2_outputs(103) <= not a;
    layer2_outputs(104) <= b;
    layer2_outputs(105) <= a and not b;
    layer2_outputs(106) <= not (a and b);
    layer2_outputs(107) <= '0';
    layer2_outputs(108) <= a and b;
    layer2_outputs(109) <= not (a or b);
    layer2_outputs(110) <= a xor b;
    layer2_outputs(111) <= not a or b;
    layer2_outputs(112) <= not a;
    layer2_outputs(113) <= b;
    layer2_outputs(114) <= a and b;
    layer2_outputs(115) <= not b or a;
    layer2_outputs(116) <= not a;
    layer2_outputs(117) <= not b;
    layer2_outputs(118) <= not (a and b);
    layer2_outputs(119) <= a;
    layer2_outputs(120) <= not b or a;
    layer2_outputs(121) <= not b;
    layer2_outputs(122) <= a xor b;
    layer2_outputs(123) <= b;
    layer2_outputs(124) <= b;
    layer2_outputs(125) <= a or b;
    layer2_outputs(126) <= not b;
    layer2_outputs(127) <= b;
    layer2_outputs(128) <= a and b;
    layer2_outputs(129) <= a;
    layer2_outputs(130) <= '0';
    layer2_outputs(131) <= not a;
    layer2_outputs(132) <= '0';
    layer2_outputs(133) <= not (a and b);
    layer2_outputs(134) <= not b or a;
    layer2_outputs(135) <= '1';
    layer2_outputs(136) <= a and not b;
    layer2_outputs(137) <= a or b;
    layer2_outputs(138) <= a or b;
    layer2_outputs(139) <= a and not b;
    layer2_outputs(140) <= not (a or b);
    layer2_outputs(141) <= '0';
    layer2_outputs(142) <= '0';
    layer2_outputs(143) <= a and b;
    layer2_outputs(144) <= not b or a;
    layer2_outputs(145) <= b and not a;
    layer2_outputs(146) <= not a or b;
    layer2_outputs(147) <= not b or a;
    layer2_outputs(148) <= '0';
    layer2_outputs(149) <= b and not a;
    layer2_outputs(150) <= '0';
    layer2_outputs(151) <= a;
    layer2_outputs(152) <= a;
    layer2_outputs(153) <= a and not b;
    layer2_outputs(154) <= b and not a;
    layer2_outputs(155) <= a xor b;
    layer2_outputs(156) <= b and not a;
    layer2_outputs(157) <= a or b;
    layer2_outputs(158) <= b;
    layer2_outputs(159) <= '1';
    layer2_outputs(160) <= a and b;
    layer2_outputs(161) <= not a or b;
    layer2_outputs(162) <= a or b;
    layer2_outputs(163) <= b and not a;
    layer2_outputs(164) <= not (a and b);
    layer2_outputs(165) <= '1';
    layer2_outputs(166) <= a and not b;
    layer2_outputs(167) <= b and not a;
    layer2_outputs(168) <= not (a or b);
    layer2_outputs(169) <= b and not a;
    layer2_outputs(170) <= b and not a;
    layer2_outputs(171) <= a and b;
    layer2_outputs(172) <= '0';
    layer2_outputs(173) <= not a or b;
    layer2_outputs(174) <= not a;
    layer2_outputs(175) <= not (a and b);
    layer2_outputs(176) <= a and b;
    layer2_outputs(177) <= b;
    layer2_outputs(178) <= '0';
    layer2_outputs(179) <= not a or b;
    layer2_outputs(180) <= not (a and b);
    layer2_outputs(181) <= a and not b;
    layer2_outputs(182) <= b and not a;
    layer2_outputs(183) <= not (a and b);
    layer2_outputs(184) <= a and b;
    layer2_outputs(185) <= not (a or b);
    layer2_outputs(186) <= a and b;
    layer2_outputs(187) <= a or b;
    layer2_outputs(188) <= not (a or b);
    layer2_outputs(189) <= not a;
    layer2_outputs(190) <= not (a or b);
    layer2_outputs(191) <= a and b;
    layer2_outputs(192) <= '0';
    layer2_outputs(193) <= a and b;
    layer2_outputs(194) <= not b;
    layer2_outputs(195) <= not (a and b);
    layer2_outputs(196) <= not a;
    layer2_outputs(197) <= b;
    layer2_outputs(198) <= a and not b;
    layer2_outputs(199) <= not (a or b);
    layer2_outputs(200) <= '0';
    layer2_outputs(201) <= not a or b;
    layer2_outputs(202) <= a and not b;
    layer2_outputs(203) <= '0';
    layer2_outputs(204) <= b and not a;
    layer2_outputs(205) <= a;
    layer2_outputs(206) <= b;
    layer2_outputs(207) <= not b;
    layer2_outputs(208) <= '0';
    layer2_outputs(209) <= a xor b;
    layer2_outputs(210) <= a xor b;
    layer2_outputs(211) <= not b or a;
    layer2_outputs(212) <= a and b;
    layer2_outputs(213) <= not a or b;
    layer2_outputs(214) <= not a;
    layer2_outputs(215) <= not (a xor b);
    layer2_outputs(216) <= a;
    layer2_outputs(217) <= not b or a;
    layer2_outputs(218) <= a;
    layer2_outputs(219) <= not a or b;
    layer2_outputs(220) <= '0';
    layer2_outputs(221) <= '0';
    layer2_outputs(222) <= b and not a;
    layer2_outputs(223) <= a or b;
    layer2_outputs(224) <= a and b;
    layer2_outputs(225) <= not b;
    layer2_outputs(226) <= a;
    layer2_outputs(227) <= not a or b;
    layer2_outputs(228) <= not a or b;
    layer2_outputs(229) <= '1';
    layer2_outputs(230) <= a or b;
    layer2_outputs(231) <= '1';
    layer2_outputs(232) <= b and not a;
    layer2_outputs(233) <= not b;
    layer2_outputs(234) <= a or b;
    layer2_outputs(235) <= not (a or b);
    layer2_outputs(236) <= not a;
    layer2_outputs(237) <= not (a or b);
    layer2_outputs(238) <= b;
    layer2_outputs(239) <= a and b;
    layer2_outputs(240) <= a and b;
    layer2_outputs(241) <= '1';
    layer2_outputs(242) <= not b or a;
    layer2_outputs(243) <= not (a and b);
    layer2_outputs(244) <= not a or b;
    layer2_outputs(245) <= not b;
    layer2_outputs(246) <= b;
    layer2_outputs(247) <= not b or a;
    layer2_outputs(248) <= not b;
    layer2_outputs(249) <= a;
    layer2_outputs(250) <= a;
    layer2_outputs(251) <= b and not a;
    layer2_outputs(252) <= not (a or b);
    layer2_outputs(253) <= a and b;
    layer2_outputs(254) <= not b;
    layer2_outputs(255) <= not (a xor b);
    layer2_outputs(256) <= a;
    layer2_outputs(257) <= not a;
    layer2_outputs(258) <= not a or b;
    layer2_outputs(259) <= not b;
    layer2_outputs(260) <= not b;
    layer2_outputs(261) <= not (a and b);
    layer2_outputs(262) <= not b;
    layer2_outputs(263) <= b;
    layer2_outputs(264) <= not a;
    layer2_outputs(265) <= not (a or b);
    layer2_outputs(266) <= a and not b;
    layer2_outputs(267) <= not b;
    layer2_outputs(268) <= a or b;
    layer2_outputs(269) <= a or b;
    layer2_outputs(270) <= b;
    layer2_outputs(271) <= '0';
    layer2_outputs(272) <= b and not a;
    layer2_outputs(273) <= b;
    layer2_outputs(274) <= a;
    layer2_outputs(275) <= not a or b;
    layer2_outputs(276) <= not b or a;
    layer2_outputs(277) <= not b or a;
    layer2_outputs(278) <= b;
    layer2_outputs(279) <= not b;
    layer2_outputs(280) <= not b;
    layer2_outputs(281) <= b;
    layer2_outputs(282) <= not (a or b);
    layer2_outputs(283) <= a and not b;
    layer2_outputs(284) <= a and b;
    layer2_outputs(285) <= '1';
    layer2_outputs(286) <= not b or a;
    layer2_outputs(287) <= not (a xor b);
    layer2_outputs(288) <= not (a and b);
    layer2_outputs(289) <= not (a or b);
    layer2_outputs(290) <= not (a or b);
    layer2_outputs(291) <= a and not b;
    layer2_outputs(292) <= '0';
    layer2_outputs(293) <= not b;
    layer2_outputs(294) <= not (a or b);
    layer2_outputs(295) <= '0';
    layer2_outputs(296) <= not (a xor b);
    layer2_outputs(297) <= not b;
    layer2_outputs(298) <= not a or b;
    layer2_outputs(299) <= b;
    layer2_outputs(300) <= b and not a;
    layer2_outputs(301) <= not (a and b);
    layer2_outputs(302) <= '0';
    layer2_outputs(303) <= b;
    layer2_outputs(304) <= not (a or b);
    layer2_outputs(305) <= not b or a;
    layer2_outputs(306) <= a;
    layer2_outputs(307) <= not (a or b);
    layer2_outputs(308) <= b;
    layer2_outputs(309) <= not b;
    layer2_outputs(310) <= not (a and b);
    layer2_outputs(311) <= a and b;
    layer2_outputs(312) <= a xor b;
    layer2_outputs(313) <= not b or a;
    layer2_outputs(314) <= not (a and b);
    layer2_outputs(315) <= not b;
    layer2_outputs(316) <= not (a or b);
    layer2_outputs(317) <= not b;
    layer2_outputs(318) <= not b;
    layer2_outputs(319) <= a;
    layer2_outputs(320) <= a;
    layer2_outputs(321) <= a xor b;
    layer2_outputs(322) <= not a or b;
    layer2_outputs(323) <= not b or a;
    layer2_outputs(324) <= a;
    layer2_outputs(325) <= '0';
    layer2_outputs(326) <= '1';
    layer2_outputs(327) <= not b or a;
    layer2_outputs(328) <= not a or b;
    layer2_outputs(329) <= not b;
    layer2_outputs(330) <= not (a and b);
    layer2_outputs(331) <= not a or b;
    layer2_outputs(332) <= not a;
    layer2_outputs(333) <= a and not b;
    layer2_outputs(334) <= not (a and b);
    layer2_outputs(335) <= b;
    layer2_outputs(336) <= b and not a;
    layer2_outputs(337) <= not a;
    layer2_outputs(338) <= '1';
    layer2_outputs(339) <= not b;
    layer2_outputs(340) <= not (a or b);
    layer2_outputs(341) <= not b;
    layer2_outputs(342) <= not b or a;
    layer2_outputs(343) <= not a or b;
    layer2_outputs(344) <= not b or a;
    layer2_outputs(345) <= not b;
    layer2_outputs(346) <= b;
    layer2_outputs(347) <= not (a or b);
    layer2_outputs(348) <= a or b;
    layer2_outputs(349) <= not b or a;
    layer2_outputs(350) <= not (a and b);
    layer2_outputs(351) <= not b;
    layer2_outputs(352) <= a and not b;
    layer2_outputs(353) <= b;
    layer2_outputs(354) <= b;
    layer2_outputs(355) <= a and not b;
    layer2_outputs(356) <= a;
    layer2_outputs(357) <= b;
    layer2_outputs(358) <= '0';
    layer2_outputs(359) <= a and not b;
    layer2_outputs(360) <= not a;
    layer2_outputs(361) <= not b or a;
    layer2_outputs(362) <= not b or a;
    layer2_outputs(363) <= not a or b;
    layer2_outputs(364) <= not a;
    layer2_outputs(365) <= not b;
    layer2_outputs(366) <= '0';
    layer2_outputs(367) <= '1';
    layer2_outputs(368) <= a and not b;
    layer2_outputs(369) <= not a;
    layer2_outputs(370) <= not (a or b);
    layer2_outputs(371) <= not (a and b);
    layer2_outputs(372) <= not (a and b);
    layer2_outputs(373) <= not a;
    layer2_outputs(374) <= not (a and b);
    layer2_outputs(375) <= a or b;
    layer2_outputs(376) <= '0';
    layer2_outputs(377) <= a or b;
    layer2_outputs(378) <= b;
    layer2_outputs(379) <= a and b;
    layer2_outputs(380) <= a and b;
    layer2_outputs(381) <= not (a or b);
    layer2_outputs(382) <= not (a and b);
    layer2_outputs(383) <= a and not b;
    layer2_outputs(384) <= not b;
    layer2_outputs(385) <= not b or a;
    layer2_outputs(386) <= a and b;
    layer2_outputs(387) <= not a or b;
    layer2_outputs(388) <= not (a xor b);
    layer2_outputs(389) <= not a or b;
    layer2_outputs(390) <= not b or a;
    layer2_outputs(391) <= b and not a;
    layer2_outputs(392) <= b and not a;
    layer2_outputs(393) <= '1';
    layer2_outputs(394) <= a or b;
    layer2_outputs(395) <= not (a and b);
    layer2_outputs(396) <= not (a xor b);
    layer2_outputs(397) <= a and b;
    layer2_outputs(398) <= not (a and b);
    layer2_outputs(399) <= '1';
    layer2_outputs(400) <= not (a or b);
    layer2_outputs(401) <= a xor b;
    layer2_outputs(402) <= b and not a;
    layer2_outputs(403) <= b;
    layer2_outputs(404) <= not (a or b);
    layer2_outputs(405) <= not a;
    layer2_outputs(406) <= not (a xor b);
    layer2_outputs(407) <= not a or b;
    layer2_outputs(408) <= '0';
    layer2_outputs(409) <= not a or b;
    layer2_outputs(410) <= '1';
    layer2_outputs(411) <= not b or a;
    layer2_outputs(412) <= not (a and b);
    layer2_outputs(413) <= b and not a;
    layer2_outputs(414) <= not a or b;
    layer2_outputs(415) <= a and not b;
    layer2_outputs(416) <= not a or b;
    layer2_outputs(417) <= a and not b;
    layer2_outputs(418) <= '1';
    layer2_outputs(419) <= not a or b;
    layer2_outputs(420) <= not a or b;
    layer2_outputs(421) <= b and not a;
    layer2_outputs(422) <= not (a or b);
    layer2_outputs(423) <= not b;
    layer2_outputs(424) <= not b or a;
    layer2_outputs(425) <= '1';
    layer2_outputs(426) <= a or b;
    layer2_outputs(427) <= a and not b;
    layer2_outputs(428) <= b and not a;
    layer2_outputs(429) <= a and not b;
    layer2_outputs(430) <= a;
    layer2_outputs(431) <= not b;
    layer2_outputs(432) <= b and not a;
    layer2_outputs(433) <= a and b;
    layer2_outputs(434) <= '0';
    layer2_outputs(435) <= not a;
    layer2_outputs(436) <= a and b;
    layer2_outputs(437) <= a and not b;
    layer2_outputs(438) <= not b or a;
    layer2_outputs(439) <= not a;
    layer2_outputs(440) <= not (a or b);
    layer2_outputs(441) <= b and not a;
    layer2_outputs(442) <= b and not a;
    layer2_outputs(443) <= not (a and b);
    layer2_outputs(444) <= not a;
    layer2_outputs(445) <= b;
    layer2_outputs(446) <= a and b;
    layer2_outputs(447) <= b and not a;
    layer2_outputs(448) <= not b or a;
    layer2_outputs(449) <= a;
    layer2_outputs(450) <= b and not a;
    layer2_outputs(451) <= not a or b;
    layer2_outputs(452) <= '0';
    layer2_outputs(453) <= a;
    layer2_outputs(454) <= not a or b;
    layer2_outputs(455) <= a and b;
    layer2_outputs(456) <= a;
    layer2_outputs(457) <= '0';
    layer2_outputs(458) <= b;
    layer2_outputs(459) <= a and b;
    layer2_outputs(460) <= a or b;
    layer2_outputs(461) <= '0';
    layer2_outputs(462) <= b and not a;
    layer2_outputs(463) <= a and b;
    layer2_outputs(464) <= a or b;
    layer2_outputs(465) <= not (a xor b);
    layer2_outputs(466) <= not a;
    layer2_outputs(467) <= not b or a;
    layer2_outputs(468) <= b and not a;
    layer2_outputs(469) <= not (a or b);
    layer2_outputs(470) <= '0';
    layer2_outputs(471) <= a and not b;
    layer2_outputs(472) <= not a or b;
    layer2_outputs(473) <= b and not a;
    layer2_outputs(474) <= not (a or b);
    layer2_outputs(475) <= a and b;
    layer2_outputs(476) <= a and not b;
    layer2_outputs(477) <= '0';
    layer2_outputs(478) <= '0';
    layer2_outputs(479) <= '1';
    layer2_outputs(480) <= a and not b;
    layer2_outputs(481) <= a;
    layer2_outputs(482) <= a;
    layer2_outputs(483) <= '1';
    layer2_outputs(484) <= not b or a;
    layer2_outputs(485) <= not a or b;
    layer2_outputs(486) <= a and b;
    layer2_outputs(487) <= not a;
    layer2_outputs(488) <= not a;
    layer2_outputs(489) <= not b;
    layer2_outputs(490) <= b and not a;
    layer2_outputs(491) <= a and b;
    layer2_outputs(492) <= not (a or b);
    layer2_outputs(493) <= not (a or b);
    layer2_outputs(494) <= a;
    layer2_outputs(495) <= not a;
    layer2_outputs(496) <= '0';
    layer2_outputs(497) <= b;
    layer2_outputs(498) <= '0';
    layer2_outputs(499) <= a and not b;
    layer2_outputs(500) <= not b or a;
    layer2_outputs(501) <= not b;
    layer2_outputs(502) <= a;
    layer2_outputs(503) <= b and not a;
    layer2_outputs(504) <= not a or b;
    layer2_outputs(505) <= not (a xor b);
    layer2_outputs(506) <= a;
    layer2_outputs(507) <= a and b;
    layer2_outputs(508) <= not a;
    layer2_outputs(509) <= not b or a;
    layer2_outputs(510) <= '1';
    layer2_outputs(511) <= not (a and b);
    layer2_outputs(512) <= not (a or b);
    layer2_outputs(513) <= a;
    layer2_outputs(514) <= a or b;
    layer2_outputs(515) <= '0';
    layer2_outputs(516) <= a;
    layer2_outputs(517) <= '0';
    layer2_outputs(518) <= not b;
    layer2_outputs(519) <= not (a and b);
    layer2_outputs(520) <= a and b;
    layer2_outputs(521) <= not b or a;
    layer2_outputs(522) <= b and not a;
    layer2_outputs(523) <= '1';
    layer2_outputs(524) <= '0';
    layer2_outputs(525) <= not (a and b);
    layer2_outputs(526) <= not a;
    layer2_outputs(527) <= not b;
    layer2_outputs(528) <= a and not b;
    layer2_outputs(529) <= '0';
    layer2_outputs(530) <= not (a or b);
    layer2_outputs(531) <= not (a and b);
    layer2_outputs(532) <= not b or a;
    layer2_outputs(533) <= a;
    layer2_outputs(534) <= not (a or b);
    layer2_outputs(535) <= not a or b;
    layer2_outputs(536) <= not a or b;
    layer2_outputs(537) <= not b;
    layer2_outputs(538) <= a and not b;
    layer2_outputs(539) <= not (a and b);
    layer2_outputs(540) <= not a;
    layer2_outputs(541) <= a or b;
    layer2_outputs(542) <= not b or a;
    layer2_outputs(543) <= a;
    layer2_outputs(544) <= b;
    layer2_outputs(545) <= a and not b;
    layer2_outputs(546) <= b;
    layer2_outputs(547) <= '0';
    layer2_outputs(548) <= a or b;
    layer2_outputs(549) <= '1';
    layer2_outputs(550) <= not (a or b);
    layer2_outputs(551) <= '1';
    layer2_outputs(552) <= '1';
    layer2_outputs(553) <= not (a and b);
    layer2_outputs(554) <= not (a or b);
    layer2_outputs(555) <= '1';
    layer2_outputs(556) <= not b or a;
    layer2_outputs(557) <= not a;
    layer2_outputs(558) <= not a or b;
    layer2_outputs(559) <= b;
    layer2_outputs(560) <= not a;
    layer2_outputs(561) <= a and b;
    layer2_outputs(562) <= a and b;
    layer2_outputs(563) <= b;
    layer2_outputs(564) <= '0';
    layer2_outputs(565) <= a;
    layer2_outputs(566) <= b and not a;
    layer2_outputs(567) <= not (a and b);
    layer2_outputs(568) <= '1';
    layer2_outputs(569) <= a;
    layer2_outputs(570) <= '1';
    layer2_outputs(571) <= not a;
    layer2_outputs(572) <= '1';
    layer2_outputs(573) <= a or b;
    layer2_outputs(574) <= b and not a;
    layer2_outputs(575) <= b and not a;
    layer2_outputs(576) <= a and b;
    layer2_outputs(577) <= not b or a;
    layer2_outputs(578) <= a or b;
    layer2_outputs(579) <= a or b;
    layer2_outputs(580) <= not a;
    layer2_outputs(581) <= a or b;
    layer2_outputs(582) <= b;
    layer2_outputs(583) <= not (a or b);
    layer2_outputs(584) <= not (a or b);
    layer2_outputs(585) <= b;
    layer2_outputs(586) <= not a;
    layer2_outputs(587) <= a;
    layer2_outputs(588) <= a or b;
    layer2_outputs(589) <= not a;
    layer2_outputs(590) <= not (a or b);
    layer2_outputs(591) <= b and not a;
    layer2_outputs(592) <= a or b;
    layer2_outputs(593) <= '1';
    layer2_outputs(594) <= a or b;
    layer2_outputs(595) <= not a or b;
    layer2_outputs(596) <= not b or a;
    layer2_outputs(597) <= not b;
    layer2_outputs(598) <= '0';
    layer2_outputs(599) <= b and not a;
    layer2_outputs(600) <= b;
    layer2_outputs(601) <= a;
    layer2_outputs(602) <= b and not a;
    layer2_outputs(603) <= not b;
    layer2_outputs(604) <= not a;
    layer2_outputs(605) <= not a or b;
    layer2_outputs(606) <= '1';
    layer2_outputs(607) <= a and b;
    layer2_outputs(608) <= not b;
    layer2_outputs(609) <= a xor b;
    layer2_outputs(610) <= a and not b;
    layer2_outputs(611) <= a and not b;
    layer2_outputs(612) <= not (a xor b);
    layer2_outputs(613) <= b and not a;
    layer2_outputs(614) <= not a;
    layer2_outputs(615) <= '0';
    layer2_outputs(616) <= '1';
    layer2_outputs(617) <= a;
    layer2_outputs(618) <= not (a and b);
    layer2_outputs(619) <= '0';
    layer2_outputs(620) <= not (a or b);
    layer2_outputs(621) <= not a or b;
    layer2_outputs(622) <= not b or a;
    layer2_outputs(623) <= a;
    layer2_outputs(624) <= '0';
    layer2_outputs(625) <= b;
    layer2_outputs(626) <= '0';
    layer2_outputs(627) <= '1';
    layer2_outputs(628) <= not (a or b);
    layer2_outputs(629) <= not (a and b);
    layer2_outputs(630) <= b;
    layer2_outputs(631) <= not a or b;
    layer2_outputs(632) <= b;
    layer2_outputs(633) <= not (a or b);
    layer2_outputs(634) <= not a;
    layer2_outputs(635) <= a;
    layer2_outputs(636) <= a and not b;
    layer2_outputs(637) <= '1';
    layer2_outputs(638) <= b and not a;
    layer2_outputs(639) <= '0';
    layer2_outputs(640) <= not b;
    layer2_outputs(641) <= b and not a;
    layer2_outputs(642) <= '0';
    layer2_outputs(643) <= not b or a;
    layer2_outputs(644) <= not (a and b);
    layer2_outputs(645) <= not a;
    layer2_outputs(646) <= a and not b;
    layer2_outputs(647) <= '0';
    layer2_outputs(648) <= '1';
    layer2_outputs(649) <= not (a and b);
    layer2_outputs(650) <= a and b;
    layer2_outputs(651) <= a or b;
    layer2_outputs(652) <= not (a or b);
    layer2_outputs(653) <= a;
    layer2_outputs(654) <= not b;
    layer2_outputs(655) <= not a or b;
    layer2_outputs(656) <= b and not a;
    layer2_outputs(657) <= a xor b;
    layer2_outputs(658) <= '1';
    layer2_outputs(659) <= not b;
    layer2_outputs(660) <= not (a xor b);
    layer2_outputs(661) <= a and b;
    layer2_outputs(662) <= '0';
    layer2_outputs(663) <= '1';
    layer2_outputs(664) <= a and not b;
    layer2_outputs(665) <= '0';
    layer2_outputs(666) <= '1';
    layer2_outputs(667) <= not a or b;
    layer2_outputs(668) <= a and b;
    layer2_outputs(669) <= a and b;
    layer2_outputs(670) <= not a or b;
    layer2_outputs(671) <= not (a and b);
    layer2_outputs(672) <= a and not b;
    layer2_outputs(673) <= b;
    layer2_outputs(674) <= a or b;
    layer2_outputs(675) <= not a or b;
    layer2_outputs(676) <= a and not b;
    layer2_outputs(677) <= not a;
    layer2_outputs(678) <= a and b;
    layer2_outputs(679) <= a and not b;
    layer2_outputs(680) <= not a;
    layer2_outputs(681) <= '0';
    layer2_outputs(682) <= a or b;
    layer2_outputs(683) <= '0';
    layer2_outputs(684) <= not b;
    layer2_outputs(685) <= '0';
    layer2_outputs(686) <= '1';
    layer2_outputs(687) <= '0';
    layer2_outputs(688) <= a and b;
    layer2_outputs(689) <= a and not b;
    layer2_outputs(690) <= a and b;
    layer2_outputs(691) <= not b;
    layer2_outputs(692) <= not b;
    layer2_outputs(693) <= a and not b;
    layer2_outputs(694) <= not b;
    layer2_outputs(695) <= a;
    layer2_outputs(696) <= a and b;
    layer2_outputs(697) <= not (a and b);
    layer2_outputs(698) <= a or b;
    layer2_outputs(699) <= '1';
    layer2_outputs(700) <= not a or b;
    layer2_outputs(701) <= not (a xor b);
    layer2_outputs(702) <= not (a and b);
    layer2_outputs(703) <= not (a and b);
    layer2_outputs(704) <= not (a or b);
    layer2_outputs(705) <= not (a xor b);
    layer2_outputs(706) <= b;
    layer2_outputs(707) <= not b or a;
    layer2_outputs(708) <= b;
    layer2_outputs(709) <= '0';
    layer2_outputs(710) <= '0';
    layer2_outputs(711) <= not a;
    layer2_outputs(712) <= b and not a;
    layer2_outputs(713) <= a;
    layer2_outputs(714) <= not a;
    layer2_outputs(715) <= a or b;
    layer2_outputs(716) <= a and b;
    layer2_outputs(717) <= not (a and b);
    layer2_outputs(718) <= a and b;
    layer2_outputs(719) <= a or b;
    layer2_outputs(720) <= '1';
    layer2_outputs(721) <= a or b;
    layer2_outputs(722) <= not (a or b);
    layer2_outputs(723) <= b;
    layer2_outputs(724) <= not a;
    layer2_outputs(725) <= a;
    layer2_outputs(726) <= not a or b;
    layer2_outputs(727) <= not b;
    layer2_outputs(728) <= not a or b;
    layer2_outputs(729) <= b and not a;
    layer2_outputs(730) <= not a or b;
    layer2_outputs(731) <= not (a and b);
    layer2_outputs(732) <= a or b;
    layer2_outputs(733) <= b;
    layer2_outputs(734) <= '0';
    layer2_outputs(735) <= not a;
    layer2_outputs(736) <= a and b;
    layer2_outputs(737) <= '0';
    layer2_outputs(738) <= a or b;
    layer2_outputs(739) <= not b or a;
    layer2_outputs(740) <= not b;
    layer2_outputs(741) <= not b or a;
    layer2_outputs(742) <= not a;
    layer2_outputs(743) <= not (a and b);
    layer2_outputs(744) <= not (a or b);
    layer2_outputs(745) <= '0';
    layer2_outputs(746) <= not (a and b);
    layer2_outputs(747) <= b and not a;
    layer2_outputs(748) <= '0';
    layer2_outputs(749) <= a or b;
    layer2_outputs(750) <= not b;
    layer2_outputs(751) <= '0';
    layer2_outputs(752) <= a and not b;
    layer2_outputs(753) <= not (a and b);
    layer2_outputs(754) <= not (a and b);
    layer2_outputs(755) <= not b;
    layer2_outputs(756) <= not (a and b);
    layer2_outputs(757) <= a and not b;
    layer2_outputs(758) <= '0';
    layer2_outputs(759) <= a and not b;
    layer2_outputs(760) <= a and b;
    layer2_outputs(761) <= not (a or b);
    layer2_outputs(762) <= not (a and b);
    layer2_outputs(763) <= '0';
    layer2_outputs(764) <= a;
    layer2_outputs(765) <= a and not b;
    layer2_outputs(766) <= a and not b;
    layer2_outputs(767) <= not b;
    layer2_outputs(768) <= not a or b;
    layer2_outputs(769) <= '1';
    layer2_outputs(770) <= a;
    layer2_outputs(771) <= a and b;
    layer2_outputs(772) <= not a or b;
    layer2_outputs(773) <= not (a and b);
    layer2_outputs(774) <= b and not a;
    layer2_outputs(775) <= a and not b;
    layer2_outputs(776) <= not (a or b);
    layer2_outputs(777) <= not (a or b);
    layer2_outputs(778) <= not (a or b);
    layer2_outputs(779) <= not (a and b);
    layer2_outputs(780) <= a and b;
    layer2_outputs(781) <= '0';
    layer2_outputs(782) <= '0';
    layer2_outputs(783) <= not (a and b);
    layer2_outputs(784) <= not (a and b);
    layer2_outputs(785) <= not a or b;
    layer2_outputs(786) <= '0';
    layer2_outputs(787) <= '1';
    layer2_outputs(788) <= '1';
    layer2_outputs(789) <= not a;
    layer2_outputs(790) <= not (a xor b);
    layer2_outputs(791) <= a xor b;
    layer2_outputs(792) <= '0';
    layer2_outputs(793) <= a or b;
    layer2_outputs(794) <= a;
    layer2_outputs(795) <= a or b;
    layer2_outputs(796) <= not b or a;
    layer2_outputs(797) <= '0';
    layer2_outputs(798) <= b and not a;
    layer2_outputs(799) <= not b or a;
    layer2_outputs(800) <= b and not a;
    layer2_outputs(801) <= not a or b;
    layer2_outputs(802) <= '1';
    layer2_outputs(803) <= not b or a;
    layer2_outputs(804) <= not (a or b);
    layer2_outputs(805) <= a and b;
    layer2_outputs(806) <= not a;
    layer2_outputs(807) <= '1';
    layer2_outputs(808) <= not (a and b);
    layer2_outputs(809) <= a or b;
    layer2_outputs(810) <= '0';
    layer2_outputs(811) <= a;
    layer2_outputs(812) <= a xor b;
    layer2_outputs(813) <= '0';
    layer2_outputs(814) <= '0';
    layer2_outputs(815) <= not a;
    layer2_outputs(816) <= not b;
    layer2_outputs(817) <= not (a and b);
    layer2_outputs(818) <= a or b;
    layer2_outputs(819) <= '1';
    layer2_outputs(820) <= not (a or b);
    layer2_outputs(821) <= a and b;
    layer2_outputs(822) <= not (a or b);
    layer2_outputs(823) <= b;
    layer2_outputs(824) <= b;
    layer2_outputs(825) <= not a or b;
    layer2_outputs(826) <= a and not b;
    layer2_outputs(827) <= a and not b;
    layer2_outputs(828) <= not b or a;
    layer2_outputs(829) <= a and not b;
    layer2_outputs(830) <= '0';
    layer2_outputs(831) <= b;
    layer2_outputs(832) <= a or b;
    layer2_outputs(833) <= a or b;
    layer2_outputs(834) <= b;
    layer2_outputs(835) <= not b;
    layer2_outputs(836) <= a and b;
    layer2_outputs(837) <= b and not a;
    layer2_outputs(838) <= not a or b;
    layer2_outputs(839) <= a and not b;
    layer2_outputs(840) <= b;
    layer2_outputs(841) <= not (a xor b);
    layer2_outputs(842) <= not (a or b);
    layer2_outputs(843) <= b and not a;
    layer2_outputs(844) <= not b or a;
    layer2_outputs(845) <= '0';
    layer2_outputs(846) <= not a;
    layer2_outputs(847) <= '1';
    layer2_outputs(848) <= not a;
    layer2_outputs(849) <= a or b;
    layer2_outputs(850) <= not a or b;
    layer2_outputs(851) <= a or b;
    layer2_outputs(852) <= b and not a;
    layer2_outputs(853) <= a and not b;
    layer2_outputs(854) <= '0';
    layer2_outputs(855) <= not a or b;
    layer2_outputs(856) <= not a;
    layer2_outputs(857) <= b and not a;
    layer2_outputs(858) <= a;
    layer2_outputs(859) <= '0';
    layer2_outputs(860) <= a and b;
    layer2_outputs(861) <= not a;
    layer2_outputs(862) <= '0';
    layer2_outputs(863) <= '0';
    layer2_outputs(864) <= not a;
    layer2_outputs(865) <= not a;
    layer2_outputs(866) <= a or b;
    layer2_outputs(867) <= not b;
    layer2_outputs(868) <= b and not a;
    layer2_outputs(869) <= b;
    layer2_outputs(870) <= b;
    layer2_outputs(871) <= b;
    layer2_outputs(872) <= a or b;
    layer2_outputs(873) <= '0';
    layer2_outputs(874) <= not (a or b);
    layer2_outputs(875) <= b and not a;
    layer2_outputs(876) <= not a;
    layer2_outputs(877) <= b and not a;
    layer2_outputs(878) <= not a;
    layer2_outputs(879) <= a and b;
    layer2_outputs(880) <= not a or b;
    layer2_outputs(881) <= a and b;
    layer2_outputs(882) <= a;
    layer2_outputs(883) <= not (a and b);
    layer2_outputs(884) <= not a;
    layer2_outputs(885) <= not (a or b);
    layer2_outputs(886) <= not (a and b);
    layer2_outputs(887) <= not a or b;
    layer2_outputs(888) <= '0';
    layer2_outputs(889) <= not a or b;
    layer2_outputs(890) <= a and not b;
    layer2_outputs(891) <= not (a and b);
    layer2_outputs(892) <= not (a and b);
    layer2_outputs(893) <= b and not a;
    layer2_outputs(894) <= not (a or b);
    layer2_outputs(895) <= not b or a;
    layer2_outputs(896) <= not a;
    layer2_outputs(897) <= not b or a;
    layer2_outputs(898) <= '0';
    layer2_outputs(899) <= not a;
    layer2_outputs(900) <= a;
    layer2_outputs(901) <= not a or b;
    layer2_outputs(902) <= b and not a;
    layer2_outputs(903) <= a xor b;
    layer2_outputs(904) <= a and b;
    layer2_outputs(905) <= a or b;
    layer2_outputs(906) <= a;
    layer2_outputs(907) <= not (a and b);
    layer2_outputs(908) <= '1';
    layer2_outputs(909) <= a or b;
    layer2_outputs(910) <= '1';
    layer2_outputs(911) <= not a;
    layer2_outputs(912) <= not b or a;
    layer2_outputs(913) <= not b or a;
    layer2_outputs(914) <= not a;
    layer2_outputs(915) <= a;
    layer2_outputs(916) <= '1';
    layer2_outputs(917) <= not b or a;
    layer2_outputs(918) <= a;
    layer2_outputs(919) <= '0';
    layer2_outputs(920) <= not (a and b);
    layer2_outputs(921) <= '1';
    layer2_outputs(922) <= not b;
    layer2_outputs(923) <= b;
    layer2_outputs(924) <= a;
    layer2_outputs(925) <= not (a and b);
    layer2_outputs(926) <= not (a or b);
    layer2_outputs(927) <= not a;
    layer2_outputs(928) <= not (a or b);
    layer2_outputs(929) <= not b or a;
    layer2_outputs(930) <= not b;
    layer2_outputs(931) <= not (a or b);
    layer2_outputs(932) <= a and b;
    layer2_outputs(933) <= not a or b;
    layer2_outputs(934) <= not b or a;
    layer2_outputs(935) <= a or b;
    layer2_outputs(936) <= a or b;
    layer2_outputs(937) <= a and not b;
    layer2_outputs(938) <= not (a and b);
    layer2_outputs(939) <= not a or b;
    layer2_outputs(940) <= a or b;
    layer2_outputs(941) <= not (a and b);
    layer2_outputs(942) <= not (a and b);
    layer2_outputs(943) <= not b;
    layer2_outputs(944) <= not (a and b);
    layer2_outputs(945) <= a or b;
    layer2_outputs(946) <= a and b;
    layer2_outputs(947) <= not a;
    layer2_outputs(948) <= a or b;
    layer2_outputs(949) <= a or b;
    layer2_outputs(950) <= '0';
    layer2_outputs(951) <= b and not a;
    layer2_outputs(952) <= not a;
    layer2_outputs(953) <= not b or a;
    layer2_outputs(954) <= not b or a;
    layer2_outputs(955) <= not a or b;
    layer2_outputs(956) <= not (a or b);
    layer2_outputs(957) <= not a;
    layer2_outputs(958) <= not (a or b);
    layer2_outputs(959) <= b;
    layer2_outputs(960) <= not (a xor b);
    layer2_outputs(961) <= '1';
    layer2_outputs(962) <= b;
    layer2_outputs(963) <= b;
    layer2_outputs(964) <= '0';
    layer2_outputs(965) <= a;
    layer2_outputs(966) <= a;
    layer2_outputs(967) <= not a or b;
    layer2_outputs(968) <= a and not b;
    layer2_outputs(969) <= not a or b;
    layer2_outputs(970) <= b;
    layer2_outputs(971) <= not b or a;
    layer2_outputs(972) <= not a;
    layer2_outputs(973) <= a and b;
    layer2_outputs(974) <= a;
    layer2_outputs(975) <= not a;
    layer2_outputs(976) <= not (a and b);
    layer2_outputs(977) <= '1';
    layer2_outputs(978) <= '0';
    layer2_outputs(979) <= not (a and b);
    layer2_outputs(980) <= a and b;
    layer2_outputs(981) <= not b or a;
    layer2_outputs(982) <= not a or b;
    layer2_outputs(983) <= a;
    layer2_outputs(984) <= a;
    layer2_outputs(985) <= '1';
    layer2_outputs(986) <= b;
    layer2_outputs(987) <= not b or a;
    layer2_outputs(988) <= a or b;
    layer2_outputs(989) <= '0';
    layer2_outputs(990) <= a or b;
    layer2_outputs(991) <= not a or b;
    layer2_outputs(992) <= not b;
    layer2_outputs(993) <= a and b;
    layer2_outputs(994) <= not b or a;
    layer2_outputs(995) <= '1';
    layer2_outputs(996) <= not a or b;
    layer2_outputs(997) <= '1';
    layer2_outputs(998) <= not a;
    layer2_outputs(999) <= b;
    layer2_outputs(1000) <= b;
    layer2_outputs(1001) <= a and not b;
    layer2_outputs(1002) <= not b or a;
    layer2_outputs(1003) <= b and not a;
    layer2_outputs(1004) <= b and not a;
    layer2_outputs(1005) <= not b;
    layer2_outputs(1006) <= not (a or b);
    layer2_outputs(1007) <= '0';
    layer2_outputs(1008) <= b;
    layer2_outputs(1009) <= a and not b;
    layer2_outputs(1010) <= not a or b;
    layer2_outputs(1011) <= a;
    layer2_outputs(1012) <= b;
    layer2_outputs(1013) <= '1';
    layer2_outputs(1014) <= '0';
    layer2_outputs(1015) <= b and not a;
    layer2_outputs(1016) <= b;
    layer2_outputs(1017) <= a or b;
    layer2_outputs(1018) <= not (a or b);
    layer2_outputs(1019) <= not (a or b);
    layer2_outputs(1020) <= a and not b;
    layer2_outputs(1021) <= not a;
    layer2_outputs(1022) <= '0';
    layer2_outputs(1023) <= a;
    layer2_outputs(1024) <= b;
    layer2_outputs(1025) <= not b;
    layer2_outputs(1026) <= not b;
    layer2_outputs(1027) <= not b or a;
    layer2_outputs(1028) <= a and b;
    layer2_outputs(1029) <= not b;
    layer2_outputs(1030) <= a xor b;
    layer2_outputs(1031) <= b and not a;
    layer2_outputs(1032) <= a and not b;
    layer2_outputs(1033) <= not b or a;
    layer2_outputs(1034) <= '1';
    layer2_outputs(1035) <= not b;
    layer2_outputs(1036) <= '0';
    layer2_outputs(1037) <= b;
    layer2_outputs(1038) <= not b or a;
    layer2_outputs(1039) <= not (a or b);
    layer2_outputs(1040) <= b and not a;
    layer2_outputs(1041) <= b;
    layer2_outputs(1042) <= not a or b;
    layer2_outputs(1043) <= a or b;
    layer2_outputs(1044) <= '1';
    layer2_outputs(1045) <= not (a or b);
    layer2_outputs(1046) <= a and not b;
    layer2_outputs(1047) <= not (a or b);
    layer2_outputs(1048) <= a or b;
    layer2_outputs(1049) <= not (a or b);
    layer2_outputs(1050) <= '1';
    layer2_outputs(1051) <= b and not a;
    layer2_outputs(1052) <= a or b;
    layer2_outputs(1053) <= not (a and b);
    layer2_outputs(1054) <= a;
    layer2_outputs(1055) <= '1';
    layer2_outputs(1056) <= a or b;
    layer2_outputs(1057) <= not a;
    layer2_outputs(1058) <= b;
    layer2_outputs(1059) <= not a or b;
    layer2_outputs(1060) <= '1';
    layer2_outputs(1061) <= not (a and b);
    layer2_outputs(1062) <= b;
    layer2_outputs(1063) <= a or b;
    layer2_outputs(1064) <= not (a or b);
    layer2_outputs(1065) <= not (a and b);
    layer2_outputs(1066) <= b and not a;
    layer2_outputs(1067) <= '1';
    layer2_outputs(1068) <= not (a and b);
    layer2_outputs(1069) <= not (a and b);
    layer2_outputs(1070) <= '0';
    layer2_outputs(1071) <= a;
    layer2_outputs(1072) <= not (a and b);
    layer2_outputs(1073) <= not a or b;
    layer2_outputs(1074) <= not (a and b);
    layer2_outputs(1075) <= '1';
    layer2_outputs(1076) <= a and b;
    layer2_outputs(1077) <= b and not a;
    layer2_outputs(1078) <= not b or a;
    layer2_outputs(1079) <= '0';
    layer2_outputs(1080) <= not a or b;
    layer2_outputs(1081) <= b and not a;
    layer2_outputs(1082) <= b and not a;
    layer2_outputs(1083) <= not b;
    layer2_outputs(1084) <= not a;
    layer2_outputs(1085) <= a or b;
    layer2_outputs(1086) <= b and not a;
    layer2_outputs(1087) <= a or b;
    layer2_outputs(1088) <= b and not a;
    layer2_outputs(1089) <= not (a or b);
    layer2_outputs(1090) <= not a;
    layer2_outputs(1091) <= a or b;
    layer2_outputs(1092) <= '0';
    layer2_outputs(1093) <= not a or b;
    layer2_outputs(1094) <= not b or a;
    layer2_outputs(1095) <= '0';
    layer2_outputs(1096) <= '1';
    layer2_outputs(1097) <= not (a xor b);
    layer2_outputs(1098) <= not b;
    layer2_outputs(1099) <= b;
    layer2_outputs(1100) <= not (a and b);
    layer2_outputs(1101) <= '0';
    layer2_outputs(1102) <= '0';
    layer2_outputs(1103) <= not b;
    layer2_outputs(1104) <= a or b;
    layer2_outputs(1105) <= not (a and b);
    layer2_outputs(1106) <= not (a or b);
    layer2_outputs(1107) <= a;
    layer2_outputs(1108) <= '1';
    layer2_outputs(1109) <= '1';
    layer2_outputs(1110) <= b and not a;
    layer2_outputs(1111) <= a;
    layer2_outputs(1112) <= b and not a;
    layer2_outputs(1113) <= a and not b;
    layer2_outputs(1114) <= '1';
    layer2_outputs(1115) <= a;
    layer2_outputs(1116) <= not a or b;
    layer2_outputs(1117) <= not (a or b);
    layer2_outputs(1118) <= not (a or b);
    layer2_outputs(1119) <= not (a and b);
    layer2_outputs(1120) <= not a;
    layer2_outputs(1121) <= a and b;
    layer2_outputs(1122) <= '1';
    layer2_outputs(1123) <= b;
    layer2_outputs(1124) <= a;
    layer2_outputs(1125) <= a and b;
    layer2_outputs(1126) <= '1';
    layer2_outputs(1127) <= a and b;
    layer2_outputs(1128) <= a and b;
    layer2_outputs(1129) <= a;
    layer2_outputs(1130) <= not (a and b);
    layer2_outputs(1131) <= '0';
    layer2_outputs(1132) <= not (a xor b);
    layer2_outputs(1133) <= not (a and b);
    layer2_outputs(1134) <= '0';
    layer2_outputs(1135) <= a or b;
    layer2_outputs(1136) <= not b;
    layer2_outputs(1137) <= not b;
    layer2_outputs(1138) <= a and b;
    layer2_outputs(1139) <= not b;
    layer2_outputs(1140) <= a and b;
    layer2_outputs(1141) <= b and not a;
    layer2_outputs(1142) <= not b;
    layer2_outputs(1143) <= b;
    layer2_outputs(1144) <= not b;
    layer2_outputs(1145) <= b;
    layer2_outputs(1146) <= a or b;
    layer2_outputs(1147) <= a;
    layer2_outputs(1148) <= a and b;
    layer2_outputs(1149) <= not a;
    layer2_outputs(1150) <= not a;
    layer2_outputs(1151) <= a;
    layer2_outputs(1152) <= b and not a;
    layer2_outputs(1153) <= not b;
    layer2_outputs(1154) <= '0';
    layer2_outputs(1155) <= a and not b;
    layer2_outputs(1156) <= '1';
    layer2_outputs(1157) <= a and not b;
    layer2_outputs(1158) <= not a or b;
    layer2_outputs(1159) <= not (a and b);
    layer2_outputs(1160) <= '0';
    layer2_outputs(1161) <= a;
    layer2_outputs(1162) <= not b or a;
    layer2_outputs(1163) <= b and not a;
    layer2_outputs(1164) <= not b or a;
    layer2_outputs(1165) <= '1';
    layer2_outputs(1166) <= a xor b;
    layer2_outputs(1167) <= a and not b;
    layer2_outputs(1168) <= not b or a;
    layer2_outputs(1169) <= not b or a;
    layer2_outputs(1170) <= a and b;
    layer2_outputs(1171) <= not a or b;
    layer2_outputs(1172) <= not a;
    layer2_outputs(1173) <= '1';
    layer2_outputs(1174) <= b and not a;
    layer2_outputs(1175) <= not (a or b);
    layer2_outputs(1176) <= not a or b;
    layer2_outputs(1177) <= a xor b;
    layer2_outputs(1178) <= b;
    layer2_outputs(1179) <= not a or b;
    layer2_outputs(1180) <= not a or b;
    layer2_outputs(1181) <= not (a and b);
    layer2_outputs(1182) <= b and not a;
    layer2_outputs(1183) <= '0';
    layer2_outputs(1184) <= a or b;
    layer2_outputs(1185) <= a or b;
    layer2_outputs(1186) <= a;
    layer2_outputs(1187) <= not a or b;
    layer2_outputs(1188) <= b and not a;
    layer2_outputs(1189) <= a or b;
    layer2_outputs(1190) <= a and not b;
    layer2_outputs(1191) <= '1';
    layer2_outputs(1192) <= not a;
    layer2_outputs(1193) <= not a;
    layer2_outputs(1194) <= not (a and b);
    layer2_outputs(1195) <= not b;
    layer2_outputs(1196) <= '0';
    layer2_outputs(1197) <= a and not b;
    layer2_outputs(1198) <= b;
    layer2_outputs(1199) <= not b or a;
    layer2_outputs(1200) <= a or b;
    layer2_outputs(1201) <= not a or b;
    layer2_outputs(1202) <= '0';
    layer2_outputs(1203) <= b and not a;
    layer2_outputs(1204) <= a and not b;
    layer2_outputs(1205) <= b;
    layer2_outputs(1206) <= '0';
    layer2_outputs(1207) <= '1';
    layer2_outputs(1208) <= not b or a;
    layer2_outputs(1209) <= '1';
    layer2_outputs(1210) <= not a or b;
    layer2_outputs(1211) <= b and not a;
    layer2_outputs(1212) <= b and not a;
    layer2_outputs(1213) <= not (a and b);
    layer2_outputs(1214) <= not a;
    layer2_outputs(1215) <= not (a or b);
    layer2_outputs(1216) <= '1';
    layer2_outputs(1217) <= not (a and b);
    layer2_outputs(1218) <= not (a or b);
    layer2_outputs(1219) <= not a or b;
    layer2_outputs(1220) <= b and not a;
    layer2_outputs(1221) <= b and not a;
    layer2_outputs(1222) <= '0';
    layer2_outputs(1223) <= a and not b;
    layer2_outputs(1224) <= '1';
    layer2_outputs(1225) <= not (a or b);
    layer2_outputs(1226) <= a;
    layer2_outputs(1227) <= b;
    layer2_outputs(1228) <= '1';
    layer2_outputs(1229) <= a or b;
    layer2_outputs(1230) <= not b or a;
    layer2_outputs(1231) <= not a or b;
    layer2_outputs(1232) <= not (a or b);
    layer2_outputs(1233) <= '0';
    layer2_outputs(1234) <= a and not b;
    layer2_outputs(1235) <= b and not a;
    layer2_outputs(1236) <= a or b;
    layer2_outputs(1237) <= not b;
    layer2_outputs(1238) <= a;
    layer2_outputs(1239) <= not (a or b);
    layer2_outputs(1240) <= a;
    layer2_outputs(1241) <= b;
    layer2_outputs(1242) <= b;
    layer2_outputs(1243) <= not (a and b);
    layer2_outputs(1244) <= '1';
    layer2_outputs(1245) <= not (a or b);
    layer2_outputs(1246) <= not a or b;
    layer2_outputs(1247) <= a or b;
    layer2_outputs(1248) <= b and not a;
    layer2_outputs(1249) <= '1';
    layer2_outputs(1250) <= not b or a;
    layer2_outputs(1251) <= '1';
    layer2_outputs(1252) <= not (a and b);
    layer2_outputs(1253) <= not (a and b);
    layer2_outputs(1254) <= a and b;
    layer2_outputs(1255) <= a and not b;
    layer2_outputs(1256) <= a;
    layer2_outputs(1257) <= '0';
    layer2_outputs(1258) <= a and b;
    layer2_outputs(1259) <= not (a or b);
    layer2_outputs(1260) <= b and not a;
    layer2_outputs(1261) <= not b;
    layer2_outputs(1262) <= not b or a;
    layer2_outputs(1263) <= '1';
    layer2_outputs(1264) <= a or b;
    layer2_outputs(1265) <= not b or a;
    layer2_outputs(1266) <= not b;
    layer2_outputs(1267) <= a or b;
    layer2_outputs(1268) <= not b or a;
    layer2_outputs(1269) <= not b;
    layer2_outputs(1270) <= '1';
    layer2_outputs(1271) <= b;
    layer2_outputs(1272) <= '1';
    layer2_outputs(1273) <= '1';
    layer2_outputs(1274) <= not (a or b);
    layer2_outputs(1275) <= not b;
    layer2_outputs(1276) <= a and not b;
    layer2_outputs(1277) <= not a or b;
    layer2_outputs(1278) <= '1';
    layer2_outputs(1279) <= a and not b;
    layer2_outputs(1280) <= not (a and b);
    layer2_outputs(1281) <= not a or b;
    layer2_outputs(1282) <= not (a and b);
    layer2_outputs(1283) <= not b;
    layer2_outputs(1284) <= '1';
    layer2_outputs(1285) <= not (a or b);
    layer2_outputs(1286) <= b;
    layer2_outputs(1287) <= '1';
    layer2_outputs(1288) <= not a;
    layer2_outputs(1289) <= not (a or b);
    layer2_outputs(1290) <= b;
    layer2_outputs(1291) <= '1';
    layer2_outputs(1292) <= a;
    layer2_outputs(1293) <= a and b;
    layer2_outputs(1294) <= b and not a;
    layer2_outputs(1295) <= a and b;
    layer2_outputs(1296) <= a or b;
    layer2_outputs(1297) <= b;
    layer2_outputs(1298) <= '0';
    layer2_outputs(1299) <= not a;
    layer2_outputs(1300) <= a xor b;
    layer2_outputs(1301) <= not (a and b);
    layer2_outputs(1302) <= a;
    layer2_outputs(1303) <= '0';
    layer2_outputs(1304) <= a and not b;
    layer2_outputs(1305) <= '1';
    layer2_outputs(1306) <= '0';
    layer2_outputs(1307) <= b;
    layer2_outputs(1308) <= not a;
    layer2_outputs(1309) <= b and not a;
    layer2_outputs(1310) <= not b;
    layer2_outputs(1311) <= '1';
    layer2_outputs(1312) <= a or b;
    layer2_outputs(1313) <= b;
    layer2_outputs(1314) <= b;
    layer2_outputs(1315) <= '1';
    layer2_outputs(1316) <= not b;
    layer2_outputs(1317) <= '0';
    layer2_outputs(1318) <= b and not a;
    layer2_outputs(1319) <= not a or b;
    layer2_outputs(1320) <= a and not b;
    layer2_outputs(1321) <= a;
    layer2_outputs(1322) <= a and b;
    layer2_outputs(1323) <= '1';
    layer2_outputs(1324) <= a xor b;
    layer2_outputs(1325) <= a and b;
    layer2_outputs(1326) <= a and not b;
    layer2_outputs(1327) <= '0';
    layer2_outputs(1328) <= a;
    layer2_outputs(1329) <= '0';
    layer2_outputs(1330) <= '1';
    layer2_outputs(1331) <= not a;
    layer2_outputs(1332) <= '0';
    layer2_outputs(1333) <= a;
    layer2_outputs(1334) <= a and b;
    layer2_outputs(1335) <= not a;
    layer2_outputs(1336) <= a;
    layer2_outputs(1337) <= a and b;
    layer2_outputs(1338) <= a and not b;
    layer2_outputs(1339) <= b;
    layer2_outputs(1340) <= b and not a;
    layer2_outputs(1341) <= a and not b;
    layer2_outputs(1342) <= not b or a;
    layer2_outputs(1343) <= b;
    layer2_outputs(1344) <= not (a xor b);
    layer2_outputs(1345) <= not (a or b);
    layer2_outputs(1346) <= not (a or b);
    layer2_outputs(1347) <= a xor b;
    layer2_outputs(1348) <= a and b;
    layer2_outputs(1349) <= not a or b;
    layer2_outputs(1350) <= not b or a;
    layer2_outputs(1351) <= not a;
    layer2_outputs(1352) <= not (a or b);
    layer2_outputs(1353) <= '1';
    layer2_outputs(1354) <= b and not a;
    layer2_outputs(1355) <= not (a and b);
    layer2_outputs(1356) <= not (a or b);
    layer2_outputs(1357) <= '0';
    layer2_outputs(1358) <= b and not a;
    layer2_outputs(1359) <= not (a and b);
    layer2_outputs(1360) <= a or b;
    layer2_outputs(1361) <= not (a or b);
    layer2_outputs(1362) <= not b;
    layer2_outputs(1363) <= b and not a;
    layer2_outputs(1364) <= not a or b;
    layer2_outputs(1365) <= not b;
    layer2_outputs(1366) <= not b or a;
    layer2_outputs(1367) <= not (a or b);
    layer2_outputs(1368) <= '1';
    layer2_outputs(1369) <= not (a or b);
    layer2_outputs(1370) <= a and b;
    layer2_outputs(1371) <= a or b;
    layer2_outputs(1372) <= '1';
    layer2_outputs(1373) <= a and b;
    layer2_outputs(1374) <= '1';
    layer2_outputs(1375) <= '1';
    layer2_outputs(1376) <= '1';
    layer2_outputs(1377) <= a and b;
    layer2_outputs(1378) <= not (a xor b);
    layer2_outputs(1379) <= a and not b;
    layer2_outputs(1380) <= b and not a;
    layer2_outputs(1381) <= a or b;
    layer2_outputs(1382) <= a and not b;
    layer2_outputs(1383) <= b;
    layer2_outputs(1384) <= a and not b;
    layer2_outputs(1385) <= b;
    layer2_outputs(1386) <= b;
    layer2_outputs(1387) <= a and not b;
    layer2_outputs(1388) <= a or b;
    layer2_outputs(1389) <= not (a or b);
    layer2_outputs(1390) <= not a;
    layer2_outputs(1391) <= '1';
    layer2_outputs(1392) <= '1';
    layer2_outputs(1393) <= not (a or b);
    layer2_outputs(1394) <= not (a or b);
    layer2_outputs(1395) <= '0';
    layer2_outputs(1396) <= b and not a;
    layer2_outputs(1397) <= a;
    layer2_outputs(1398) <= a and b;
    layer2_outputs(1399) <= b;
    layer2_outputs(1400) <= not a;
    layer2_outputs(1401) <= '1';
    layer2_outputs(1402) <= not (a and b);
    layer2_outputs(1403) <= a or b;
    layer2_outputs(1404) <= not b;
    layer2_outputs(1405) <= a or b;
    layer2_outputs(1406) <= '1';
    layer2_outputs(1407) <= a;
    layer2_outputs(1408) <= '1';
    layer2_outputs(1409) <= not (a and b);
    layer2_outputs(1410) <= not b or a;
    layer2_outputs(1411) <= not a or b;
    layer2_outputs(1412) <= a;
    layer2_outputs(1413) <= a xor b;
    layer2_outputs(1414) <= not (a or b);
    layer2_outputs(1415) <= not a or b;
    layer2_outputs(1416) <= not b or a;
    layer2_outputs(1417) <= a;
    layer2_outputs(1418) <= a or b;
    layer2_outputs(1419) <= a and not b;
    layer2_outputs(1420) <= '1';
    layer2_outputs(1421) <= not a;
    layer2_outputs(1422) <= not a;
    layer2_outputs(1423) <= a;
    layer2_outputs(1424) <= '0';
    layer2_outputs(1425) <= a and not b;
    layer2_outputs(1426) <= a or b;
    layer2_outputs(1427) <= a and b;
    layer2_outputs(1428) <= b and not a;
    layer2_outputs(1429) <= not b or a;
    layer2_outputs(1430) <= not (a and b);
    layer2_outputs(1431) <= not a or b;
    layer2_outputs(1432) <= '1';
    layer2_outputs(1433) <= not (a and b);
    layer2_outputs(1434) <= '0';
    layer2_outputs(1435) <= not b or a;
    layer2_outputs(1436) <= '0';
    layer2_outputs(1437) <= '1';
    layer2_outputs(1438) <= a and b;
    layer2_outputs(1439) <= a and not b;
    layer2_outputs(1440) <= not (a and b);
    layer2_outputs(1441) <= a and not b;
    layer2_outputs(1442) <= '0';
    layer2_outputs(1443) <= '0';
    layer2_outputs(1444) <= a and not b;
    layer2_outputs(1445) <= not b;
    layer2_outputs(1446) <= '0';
    layer2_outputs(1447) <= '0';
    layer2_outputs(1448) <= not b;
    layer2_outputs(1449) <= b;
    layer2_outputs(1450) <= not b or a;
    layer2_outputs(1451) <= '0';
    layer2_outputs(1452) <= a and not b;
    layer2_outputs(1453) <= '1';
    layer2_outputs(1454) <= not b or a;
    layer2_outputs(1455) <= not (a or b);
    layer2_outputs(1456) <= a and b;
    layer2_outputs(1457) <= '0';
    layer2_outputs(1458) <= not b or a;
    layer2_outputs(1459) <= not (a and b);
    layer2_outputs(1460) <= '0';
    layer2_outputs(1461) <= not (a and b);
    layer2_outputs(1462) <= not b;
    layer2_outputs(1463) <= a and b;
    layer2_outputs(1464) <= a xor b;
    layer2_outputs(1465) <= '1';
    layer2_outputs(1466) <= not a or b;
    layer2_outputs(1467) <= '1';
    layer2_outputs(1468) <= a and b;
    layer2_outputs(1469) <= not a or b;
    layer2_outputs(1470) <= b;
    layer2_outputs(1471) <= b and not a;
    layer2_outputs(1472) <= not a;
    layer2_outputs(1473) <= not (a or b);
    layer2_outputs(1474) <= a and not b;
    layer2_outputs(1475) <= a xor b;
    layer2_outputs(1476) <= b;
    layer2_outputs(1477) <= not (a and b);
    layer2_outputs(1478) <= b and not a;
    layer2_outputs(1479) <= not (a or b);
    layer2_outputs(1480) <= not (a and b);
    layer2_outputs(1481) <= a;
    layer2_outputs(1482) <= b and not a;
    layer2_outputs(1483) <= '1';
    layer2_outputs(1484) <= a and b;
    layer2_outputs(1485) <= not (a and b);
    layer2_outputs(1486) <= a and b;
    layer2_outputs(1487) <= a and b;
    layer2_outputs(1488) <= b;
    layer2_outputs(1489) <= a and b;
    layer2_outputs(1490) <= a or b;
    layer2_outputs(1491) <= not (a or b);
    layer2_outputs(1492) <= a or b;
    layer2_outputs(1493) <= a and not b;
    layer2_outputs(1494) <= '1';
    layer2_outputs(1495) <= not (a or b);
    layer2_outputs(1496) <= '0';
    layer2_outputs(1497) <= not b or a;
    layer2_outputs(1498) <= not a;
    layer2_outputs(1499) <= not (a and b);
    layer2_outputs(1500) <= a or b;
    layer2_outputs(1501) <= '0';
    layer2_outputs(1502) <= not b or a;
    layer2_outputs(1503) <= a and not b;
    layer2_outputs(1504) <= '0';
    layer2_outputs(1505) <= not (a and b);
    layer2_outputs(1506) <= not (a or b);
    layer2_outputs(1507) <= a and b;
    layer2_outputs(1508) <= not b;
    layer2_outputs(1509) <= b;
    layer2_outputs(1510) <= a and b;
    layer2_outputs(1511) <= not b;
    layer2_outputs(1512) <= a;
    layer2_outputs(1513) <= '1';
    layer2_outputs(1514) <= a and b;
    layer2_outputs(1515) <= not b or a;
    layer2_outputs(1516) <= not b or a;
    layer2_outputs(1517) <= a and b;
    layer2_outputs(1518) <= not a;
    layer2_outputs(1519) <= '1';
    layer2_outputs(1520) <= not a or b;
    layer2_outputs(1521) <= not a;
    layer2_outputs(1522) <= not a;
    layer2_outputs(1523) <= not a or b;
    layer2_outputs(1524) <= b and not a;
    layer2_outputs(1525) <= a and not b;
    layer2_outputs(1526) <= not b;
    layer2_outputs(1527) <= b;
    layer2_outputs(1528) <= b;
    layer2_outputs(1529) <= '0';
    layer2_outputs(1530) <= a;
    layer2_outputs(1531) <= not a;
    layer2_outputs(1532) <= not b;
    layer2_outputs(1533) <= not a or b;
    layer2_outputs(1534) <= not a;
    layer2_outputs(1535) <= not b or a;
    layer2_outputs(1536) <= not a or b;
    layer2_outputs(1537) <= b;
    layer2_outputs(1538) <= a xor b;
    layer2_outputs(1539) <= '0';
    layer2_outputs(1540) <= not a;
    layer2_outputs(1541) <= b and not a;
    layer2_outputs(1542) <= b;
    layer2_outputs(1543) <= not a or b;
    layer2_outputs(1544) <= not (a or b);
    layer2_outputs(1545) <= not b or a;
    layer2_outputs(1546) <= not (a or b);
    layer2_outputs(1547) <= b and not a;
    layer2_outputs(1548) <= not (a and b);
    layer2_outputs(1549) <= '0';
    layer2_outputs(1550) <= a;
    layer2_outputs(1551) <= a and not b;
    layer2_outputs(1552) <= a or b;
    layer2_outputs(1553) <= not (a and b);
    layer2_outputs(1554) <= b;
    layer2_outputs(1555) <= b;
    layer2_outputs(1556) <= not b;
    layer2_outputs(1557) <= a and b;
    layer2_outputs(1558) <= not (a and b);
    layer2_outputs(1559) <= a and b;
    layer2_outputs(1560) <= not (a or b);
    layer2_outputs(1561) <= a and b;
    layer2_outputs(1562) <= not b;
    layer2_outputs(1563) <= not b;
    layer2_outputs(1564) <= not a or b;
    layer2_outputs(1565) <= not (a or b);
    layer2_outputs(1566) <= not b or a;
    layer2_outputs(1567) <= b;
    layer2_outputs(1568) <= '1';
    layer2_outputs(1569) <= '0';
    layer2_outputs(1570) <= a and b;
    layer2_outputs(1571) <= a and not b;
    layer2_outputs(1572) <= not b or a;
    layer2_outputs(1573) <= a;
    layer2_outputs(1574) <= not b or a;
    layer2_outputs(1575) <= not (a and b);
    layer2_outputs(1576) <= not (a and b);
    layer2_outputs(1577) <= not b;
    layer2_outputs(1578) <= not b;
    layer2_outputs(1579) <= not (a xor b);
    layer2_outputs(1580) <= a xor b;
    layer2_outputs(1581) <= not a;
    layer2_outputs(1582) <= not a or b;
    layer2_outputs(1583) <= not a;
    layer2_outputs(1584) <= not a;
    layer2_outputs(1585) <= a or b;
    layer2_outputs(1586) <= not (a xor b);
    layer2_outputs(1587) <= b and not a;
    layer2_outputs(1588) <= '0';
    layer2_outputs(1589) <= a and not b;
    layer2_outputs(1590) <= b;
    layer2_outputs(1591) <= a and not b;
    layer2_outputs(1592) <= a xor b;
    layer2_outputs(1593) <= '1';
    layer2_outputs(1594) <= a and b;
    layer2_outputs(1595) <= not b or a;
    layer2_outputs(1596) <= b and not a;
    layer2_outputs(1597) <= b;
    layer2_outputs(1598) <= a and not b;
    layer2_outputs(1599) <= not a;
    layer2_outputs(1600) <= b;
    layer2_outputs(1601) <= '0';
    layer2_outputs(1602) <= a;
    layer2_outputs(1603) <= not b or a;
    layer2_outputs(1604) <= not a;
    layer2_outputs(1605) <= b;
    layer2_outputs(1606) <= a;
    layer2_outputs(1607) <= b;
    layer2_outputs(1608) <= not b;
    layer2_outputs(1609) <= not (a and b);
    layer2_outputs(1610) <= a;
    layer2_outputs(1611) <= '1';
    layer2_outputs(1612) <= not (a or b);
    layer2_outputs(1613) <= a and not b;
    layer2_outputs(1614) <= not (a or b);
    layer2_outputs(1615) <= not a;
    layer2_outputs(1616) <= b;
    layer2_outputs(1617) <= not a or b;
    layer2_outputs(1618) <= '1';
    layer2_outputs(1619) <= a or b;
    layer2_outputs(1620) <= a and b;
    layer2_outputs(1621) <= a and not b;
    layer2_outputs(1622) <= not (a or b);
    layer2_outputs(1623) <= b;
    layer2_outputs(1624) <= not b or a;
    layer2_outputs(1625) <= a or b;
    layer2_outputs(1626) <= not b;
    layer2_outputs(1627) <= a xor b;
    layer2_outputs(1628) <= a;
    layer2_outputs(1629) <= a and not b;
    layer2_outputs(1630) <= a or b;
    layer2_outputs(1631) <= '1';
    layer2_outputs(1632) <= not a;
    layer2_outputs(1633) <= not a;
    layer2_outputs(1634) <= not a or b;
    layer2_outputs(1635) <= '0';
    layer2_outputs(1636) <= '1';
    layer2_outputs(1637) <= '1';
    layer2_outputs(1638) <= not a;
    layer2_outputs(1639) <= a and b;
    layer2_outputs(1640) <= a and b;
    layer2_outputs(1641) <= '1';
    layer2_outputs(1642) <= a and not b;
    layer2_outputs(1643) <= a or b;
    layer2_outputs(1644) <= not b or a;
    layer2_outputs(1645) <= not (a or b);
    layer2_outputs(1646) <= b;
    layer2_outputs(1647) <= not (a and b);
    layer2_outputs(1648) <= a or b;
    layer2_outputs(1649) <= '0';
    layer2_outputs(1650) <= '1';
    layer2_outputs(1651) <= not (a or b);
    layer2_outputs(1652) <= not (a or b);
    layer2_outputs(1653) <= not (a and b);
    layer2_outputs(1654) <= not a;
    layer2_outputs(1655) <= not (a or b);
    layer2_outputs(1656) <= not b or a;
    layer2_outputs(1657) <= b;
    layer2_outputs(1658) <= a or b;
    layer2_outputs(1659) <= not (a or b);
    layer2_outputs(1660) <= a;
    layer2_outputs(1661) <= a and b;
    layer2_outputs(1662) <= '1';
    layer2_outputs(1663) <= a and not b;
    layer2_outputs(1664) <= not b or a;
    layer2_outputs(1665) <= a xor b;
    layer2_outputs(1666) <= b;
    layer2_outputs(1667) <= not b or a;
    layer2_outputs(1668) <= b and not a;
    layer2_outputs(1669) <= a and b;
    layer2_outputs(1670) <= a or b;
    layer2_outputs(1671) <= a or b;
    layer2_outputs(1672) <= not a;
    layer2_outputs(1673) <= not (a xor b);
    layer2_outputs(1674) <= '1';
    layer2_outputs(1675) <= b and not a;
    layer2_outputs(1676) <= not b or a;
    layer2_outputs(1677) <= not b or a;
    layer2_outputs(1678) <= a and not b;
    layer2_outputs(1679) <= not a or b;
    layer2_outputs(1680) <= b and not a;
    layer2_outputs(1681) <= not a;
    layer2_outputs(1682) <= '1';
    layer2_outputs(1683) <= a or b;
    layer2_outputs(1684) <= not b or a;
    layer2_outputs(1685) <= a and not b;
    layer2_outputs(1686) <= '0';
    layer2_outputs(1687) <= not a or b;
    layer2_outputs(1688) <= not a or b;
    layer2_outputs(1689) <= a or b;
    layer2_outputs(1690) <= b;
    layer2_outputs(1691) <= not a or b;
    layer2_outputs(1692) <= b and not a;
    layer2_outputs(1693) <= not (a and b);
    layer2_outputs(1694) <= a or b;
    layer2_outputs(1695) <= not b;
    layer2_outputs(1696) <= a and not b;
    layer2_outputs(1697) <= not (a and b);
    layer2_outputs(1698) <= not a;
    layer2_outputs(1699) <= not (a and b);
    layer2_outputs(1700) <= not (a or b);
    layer2_outputs(1701) <= b;
    layer2_outputs(1702) <= not a or b;
    layer2_outputs(1703) <= '0';
    layer2_outputs(1704) <= not b or a;
    layer2_outputs(1705) <= not a or b;
    layer2_outputs(1706) <= a or b;
    layer2_outputs(1707) <= a or b;
    layer2_outputs(1708) <= '1';
    layer2_outputs(1709) <= '0';
    layer2_outputs(1710) <= a xor b;
    layer2_outputs(1711) <= not b or a;
    layer2_outputs(1712) <= a or b;
    layer2_outputs(1713) <= not b or a;
    layer2_outputs(1714) <= not (a or b);
    layer2_outputs(1715) <= b;
    layer2_outputs(1716) <= a;
    layer2_outputs(1717) <= not b or a;
    layer2_outputs(1718) <= not (a and b);
    layer2_outputs(1719) <= b;
    layer2_outputs(1720) <= not (a or b);
    layer2_outputs(1721) <= a;
    layer2_outputs(1722) <= not b or a;
    layer2_outputs(1723) <= not (a or b);
    layer2_outputs(1724) <= a and not b;
    layer2_outputs(1725) <= a;
    layer2_outputs(1726) <= not (a and b);
    layer2_outputs(1727) <= b;
    layer2_outputs(1728) <= a or b;
    layer2_outputs(1729) <= not a;
    layer2_outputs(1730) <= a;
    layer2_outputs(1731) <= '0';
    layer2_outputs(1732) <= a and b;
    layer2_outputs(1733) <= not a;
    layer2_outputs(1734) <= not b;
    layer2_outputs(1735) <= not a or b;
    layer2_outputs(1736) <= a and not b;
    layer2_outputs(1737) <= not (a xor b);
    layer2_outputs(1738) <= a and b;
    layer2_outputs(1739) <= '0';
    layer2_outputs(1740) <= not (a xor b);
    layer2_outputs(1741) <= b;
    layer2_outputs(1742) <= b;
    layer2_outputs(1743) <= not (a or b);
    layer2_outputs(1744) <= not (a xor b);
    layer2_outputs(1745) <= not (a and b);
    layer2_outputs(1746) <= a and b;
    layer2_outputs(1747) <= b;
    layer2_outputs(1748) <= a;
    layer2_outputs(1749) <= a;
    layer2_outputs(1750) <= a and b;
    layer2_outputs(1751) <= a;
    layer2_outputs(1752) <= a;
    layer2_outputs(1753) <= b;
    layer2_outputs(1754) <= '1';
    layer2_outputs(1755) <= b;
    layer2_outputs(1756) <= '0';
    layer2_outputs(1757) <= not (a or b);
    layer2_outputs(1758) <= b and not a;
    layer2_outputs(1759) <= '0';
    layer2_outputs(1760) <= a and not b;
    layer2_outputs(1761) <= not b or a;
    layer2_outputs(1762) <= not (a or b);
    layer2_outputs(1763) <= not (a or b);
    layer2_outputs(1764) <= a and b;
    layer2_outputs(1765) <= not (a and b);
    layer2_outputs(1766) <= not (a or b);
    layer2_outputs(1767) <= b and not a;
    layer2_outputs(1768) <= '0';
    layer2_outputs(1769) <= a and b;
    layer2_outputs(1770) <= not (a or b);
    layer2_outputs(1771) <= not a or b;
    layer2_outputs(1772) <= '0';
    layer2_outputs(1773) <= not b;
    layer2_outputs(1774) <= not (a or b);
    layer2_outputs(1775) <= b;
    layer2_outputs(1776) <= not (a and b);
    layer2_outputs(1777) <= a and not b;
    layer2_outputs(1778) <= a and b;
    layer2_outputs(1779) <= b;
    layer2_outputs(1780) <= not b;
    layer2_outputs(1781) <= '1';
    layer2_outputs(1782) <= b and not a;
    layer2_outputs(1783) <= a;
    layer2_outputs(1784) <= not b;
    layer2_outputs(1785) <= not a;
    layer2_outputs(1786) <= '1';
    layer2_outputs(1787) <= '0';
    layer2_outputs(1788) <= not b;
    layer2_outputs(1789) <= not (a or b);
    layer2_outputs(1790) <= not b;
    layer2_outputs(1791) <= not b or a;
    layer2_outputs(1792) <= a xor b;
    layer2_outputs(1793) <= a and b;
    layer2_outputs(1794) <= '0';
    layer2_outputs(1795) <= b;
    layer2_outputs(1796) <= '0';
    layer2_outputs(1797) <= '0';
    layer2_outputs(1798) <= '0';
    layer2_outputs(1799) <= '0';
    layer2_outputs(1800) <= a and not b;
    layer2_outputs(1801) <= '1';
    layer2_outputs(1802) <= '0';
    layer2_outputs(1803) <= not b or a;
    layer2_outputs(1804) <= a xor b;
    layer2_outputs(1805) <= a and b;
    layer2_outputs(1806) <= not (a or b);
    layer2_outputs(1807) <= a and not b;
    layer2_outputs(1808) <= not (a or b);
    layer2_outputs(1809) <= a and b;
    layer2_outputs(1810) <= '0';
    layer2_outputs(1811) <= not a;
    layer2_outputs(1812) <= not b;
    layer2_outputs(1813) <= not b;
    layer2_outputs(1814) <= a and not b;
    layer2_outputs(1815) <= not b or a;
    layer2_outputs(1816) <= a and not b;
    layer2_outputs(1817) <= a or b;
    layer2_outputs(1818) <= a and b;
    layer2_outputs(1819) <= not b or a;
    layer2_outputs(1820) <= not (a xor b);
    layer2_outputs(1821) <= b and not a;
    layer2_outputs(1822) <= a and b;
    layer2_outputs(1823) <= '0';
    layer2_outputs(1824) <= '0';
    layer2_outputs(1825) <= b;
    layer2_outputs(1826) <= a;
    layer2_outputs(1827) <= '1';
    layer2_outputs(1828) <= '1';
    layer2_outputs(1829) <= not b or a;
    layer2_outputs(1830) <= b and not a;
    layer2_outputs(1831) <= a and not b;
    layer2_outputs(1832) <= '1';
    layer2_outputs(1833) <= '0';
    layer2_outputs(1834) <= not (a and b);
    layer2_outputs(1835) <= b;
    layer2_outputs(1836) <= not b or a;
    layer2_outputs(1837) <= '0';
    layer2_outputs(1838) <= '1';
    layer2_outputs(1839) <= a or b;
    layer2_outputs(1840) <= a and b;
    layer2_outputs(1841) <= '1';
    layer2_outputs(1842) <= not a;
    layer2_outputs(1843) <= '0';
    layer2_outputs(1844) <= not a or b;
    layer2_outputs(1845) <= a and not b;
    layer2_outputs(1846) <= '0';
    layer2_outputs(1847) <= a or b;
    layer2_outputs(1848) <= b;
    layer2_outputs(1849) <= '1';
    layer2_outputs(1850) <= a xor b;
    layer2_outputs(1851) <= '1';
    layer2_outputs(1852) <= not b;
    layer2_outputs(1853) <= b;
    layer2_outputs(1854) <= '1';
    layer2_outputs(1855) <= '0';
    layer2_outputs(1856) <= b and not a;
    layer2_outputs(1857) <= b and not a;
    layer2_outputs(1858) <= a;
    layer2_outputs(1859) <= a and b;
    layer2_outputs(1860) <= a and not b;
    layer2_outputs(1861) <= not b or a;
    layer2_outputs(1862) <= not a;
    layer2_outputs(1863) <= not a;
    layer2_outputs(1864) <= not (a or b);
    layer2_outputs(1865) <= b;
    layer2_outputs(1866) <= a and b;
    layer2_outputs(1867) <= not b;
    layer2_outputs(1868) <= not a or b;
    layer2_outputs(1869) <= a and not b;
    layer2_outputs(1870) <= a;
    layer2_outputs(1871) <= a and b;
    layer2_outputs(1872) <= a and b;
    layer2_outputs(1873) <= not (a or b);
    layer2_outputs(1874) <= b;
    layer2_outputs(1875) <= a and not b;
    layer2_outputs(1876) <= not b;
    layer2_outputs(1877) <= not (a and b);
    layer2_outputs(1878) <= a xor b;
    layer2_outputs(1879) <= b;
    layer2_outputs(1880) <= a or b;
    layer2_outputs(1881) <= '0';
    layer2_outputs(1882) <= '1';
    layer2_outputs(1883) <= a or b;
    layer2_outputs(1884) <= not b;
    layer2_outputs(1885) <= not a or b;
    layer2_outputs(1886) <= b and not a;
    layer2_outputs(1887) <= b and not a;
    layer2_outputs(1888) <= not a;
    layer2_outputs(1889) <= '1';
    layer2_outputs(1890) <= '1';
    layer2_outputs(1891) <= not a;
    layer2_outputs(1892) <= not (a or b);
    layer2_outputs(1893) <= a xor b;
    layer2_outputs(1894) <= not b;
    layer2_outputs(1895) <= not b or a;
    layer2_outputs(1896) <= a and not b;
    layer2_outputs(1897) <= b;
    layer2_outputs(1898) <= not a;
    layer2_outputs(1899) <= a and not b;
    layer2_outputs(1900) <= not a or b;
    layer2_outputs(1901) <= a and not b;
    layer2_outputs(1902) <= a or b;
    layer2_outputs(1903) <= not a;
    layer2_outputs(1904) <= not (a or b);
    layer2_outputs(1905) <= not (a or b);
    layer2_outputs(1906) <= b;
    layer2_outputs(1907) <= a and b;
    layer2_outputs(1908) <= not b;
    layer2_outputs(1909) <= '0';
    layer2_outputs(1910) <= b and not a;
    layer2_outputs(1911) <= a or b;
    layer2_outputs(1912) <= '0';
    layer2_outputs(1913) <= '0';
    layer2_outputs(1914) <= not b or a;
    layer2_outputs(1915) <= not a or b;
    layer2_outputs(1916) <= not (a and b);
    layer2_outputs(1917) <= a and not b;
    layer2_outputs(1918) <= a and b;
    layer2_outputs(1919) <= '0';
    layer2_outputs(1920) <= a and b;
    layer2_outputs(1921) <= not (a or b);
    layer2_outputs(1922) <= b and not a;
    layer2_outputs(1923) <= not b or a;
    layer2_outputs(1924) <= not a;
    layer2_outputs(1925) <= not a or b;
    layer2_outputs(1926) <= not b;
    layer2_outputs(1927) <= '0';
    layer2_outputs(1928) <= '1';
    layer2_outputs(1929) <= a and b;
    layer2_outputs(1930) <= '0';
    layer2_outputs(1931) <= '0';
    layer2_outputs(1932) <= not a or b;
    layer2_outputs(1933) <= b and not a;
    layer2_outputs(1934) <= not b or a;
    layer2_outputs(1935) <= not b;
    layer2_outputs(1936) <= a xor b;
    layer2_outputs(1937) <= a and not b;
    layer2_outputs(1938) <= a or b;
    layer2_outputs(1939) <= not (a or b);
    layer2_outputs(1940) <= b and not a;
    layer2_outputs(1941) <= b and not a;
    layer2_outputs(1942) <= not a;
    layer2_outputs(1943) <= not b;
    layer2_outputs(1944) <= not a or b;
    layer2_outputs(1945) <= not a;
    layer2_outputs(1946) <= not (a xor b);
    layer2_outputs(1947) <= '0';
    layer2_outputs(1948) <= '0';
    layer2_outputs(1949) <= not b;
    layer2_outputs(1950) <= not a;
    layer2_outputs(1951) <= not b or a;
    layer2_outputs(1952) <= '1';
    layer2_outputs(1953) <= not a or b;
    layer2_outputs(1954) <= a and not b;
    layer2_outputs(1955) <= not (a and b);
    layer2_outputs(1956) <= not b;
    layer2_outputs(1957) <= not (a and b);
    layer2_outputs(1958) <= a xor b;
    layer2_outputs(1959) <= not b or a;
    layer2_outputs(1960) <= not b;
    layer2_outputs(1961) <= not a or b;
    layer2_outputs(1962) <= a and not b;
    layer2_outputs(1963) <= '1';
    layer2_outputs(1964) <= '0';
    layer2_outputs(1965) <= '1';
    layer2_outputs(1966) <= not a;
    layer2_outputs(1967) <= a;
    layer2_outputs(1968) <= a or b;
    layer2_outputs(1969) <= a;
    layer2_outputs(1970) <= a and not b;
    layer2_outputs(1971) <= not b or a;
    layer2_outputs(1972) <= a and not b;
    layer2_outputs(1973) <= not a or b;
    layer2_outputs(1974) <= '1';
    layer2_outputs(1975) <= not a or b;
    layer2_outputs(1976) <= not b or a;
    layer2_outputs(1977) <= a and not b;
    layer2_outputs(1978) <= not a or b;
    layer2_outputs(1979) <= not a;
    layer2_outputs(1980) <= not (a and b);
    layer2_outputs(1981) <= b;
    layer2_outputs(1982) <= '0';
    layer2_outputs(1983) <= not (a or b);
    layer2_outputs(1984) <= not (a and b);
    layer2_outputs(1985) <= a;
    layer2_outputs(1986) <= '1';
    layer2_outputs(1987) <= not b;
    layer2_outputs(1988) <= '1';
    layer2_outputs(1989) <= not (a and b);
    layer2_outputs(1990) <= not a or b;
    layer2_outputs(1991) <= not b;
    layer2_outputs(1992) <= not (a or b);
    layer2_outputs(1993) <= not (a xor b);
    layer2_outputs(1994) <= not b or a;
    layer2_outputs(1995) <= a and b;
    layer2_outputs(1996) <= not (a and b);
    layer2_outputs(1997) <= '1';
    layer2_outputs(1998) <= a;
    layer2_outputs(1999) <= not b;
    layer2_outputs(2000) <= '1';
    layer2_outputs(2001) <= b;
    layer2_outputs(2002) <= a and b;
    layer2_outputs(2003) <= '0';
    layer2_outputs(2004) <= not a or b;
    layer2_outputs(2005) <= '1';
    layer2_outputs(2006) <= not a or b;
    layer2_outputs(2007) <= not b;
    layer2_outputs(2008) <= b;
    layer2_outputs(2009) <= '1';
    layer2_outputs(2010) <= '0';
    layer2_outputs(2011) <= a or b;
    layer2_outputs(2012) <= not (a and b);
    layer2_outputs(2013) <= not b;
    layer2_outputs(2014) <= a;
    layer2_outputs(2015) <= not b or a;
    layer2_outputs(2016) <= a xor b;
    layer2_outputs(2017) <= '1';
    layer2_outputs(2018) <= b;
    layer2_outputs(2019) <= a and b;
    layer2_outputs(2020) <= b;
    layer2_outputs(2021) <= b and not a;
    layer2_outputs(2022) <= a and not b;
    layer2_outputs(2023) <= a and not b;
    layer2_outputs(2024) <= b;
    layer2_outputs(2025) <= not b or a;
    layer2_outputs(2026) <= not (a xor b);
    layer2_outputs(2027) <= a and b;
    layer2_outputs(2028) <= not b;
    layer2_outputs(2029) <= not a;
    layer2_outputs(2030) <= a and b;
    layer2_outputs(2031) <= a xor b;
    layer2_outputs(2032) <= not (a or b);
    layer2_outputs(2033) <= b;
    layer2_outputs(2034) <= '1';
    layer2_outputs(2035) <= not (a and b);
    layer2_outputs(2036) <= a and not b;
    layer2_outputs(2037) <= not b or a;
    layer2_outputs(2038) <= a and not b;
    layer2_outputs(2039) <= not (a and b);
    layer2_outputs(2040) <= not b;
    layer2_outputs(2041) <= '1';
    layer2_outputs(2042) <= '0';
    layer2_outputs(2043) <= '0';
    layer2_outputs(2044) <= not a;
    layer2_outputs(2045) <= a xor b;
    layer2_outputs(2046) <= not b;
    layer2_outputs(2047) <= not (a xor b);
    layer2_outputs(2048) <= b;
    layer2_outputs(2049) <= a or b;
    layer2_outputs(2050) <= not b or a;
    layer2_outputs(2051) <= b and not a;
    layer2_outputs(2052) <= a xor b;
    layer2_outputs(2053) <= not a;
    layer2_outputs(2054) <= '1';
    layer2_outputs(2055) <= b;
    layer2_outputs(2056) <= not a or b;
    layer2_outputs(2057) <= not b;
    layer2_outputs(2058) <= a or b;
    layer2_outputs(2059) <= a or b;
    layer2_outputs(2060) <= not (a or b);
    layer2_outputs(2061) <= '1';
    layer2_outputs(2062) <= '0';
    layer2_outputs(2063) <= not (a or b);
    layer2_outputs(2064) <= not b;
    layer2_outputs(2065) <= '1';
    layer2_outputs(2066) <= '1';
    layer2_outputs(2067) <= not (a and b);
    layer2_outputs(2068) <= not b;
    layer2_outputs(2069) <= a;
    layer2_outputs(2070) <= b and not a;
    layer2_outputs(2071) <= a or b;
    layer2_outputs(2072) <= '0';
    layer2_outputs(2073) <= a and not b;
    layer2_outputs(2074) <= a or b;
    layer2_outputs(2075) <= a or b;
    layer2_outputs(2076) <= '0';
    layer2_outputs(2077) <= not (a xor b);
    layer2_outputs(2078) <= not b;
    layer2_outputs(2079) <= b and not a;
    layer2_outputs(2080) <= a or b;
    layer2_outputs(2081) <= a and b;
    layer2_outputs(2082) <= a and not b;
    layer2_outputs(2083) <= not (a and b);
    layer2_outputs(2084) <= a and b;
    layer2_outputs(2085) <= a and b;
    layer2_outputs(2086) <= not (a or b);
    layer2_outputs(2087) <= not (a xor b);
    layer2_outputs(2088) <= '1';
    layer2_outputs(2089) <= a and b;
    layer2_outputs(2090) <= not (a or b);
    layer2_outputs(2091) <= a and b;
    layer2_outputs(2092) <= '0';
    layer2_outputs(2093) <= '0';
    layer2_outputs(2094) <= '0';
    layer2_outputs(2095) <= a and not b;
    layer2_outputs(2096) <= not a or b;
    layer2_outputs(2097) <= not a or b;
    layer2_outputs(2098) <= a and not b;
    layer2_outputs(2099) <= not b;
    layer2_outputs(2100) <= not a or b;
    layer2_outputs(2101) <= not (a and b);
    layer2_outputs(2102) <= a and b;
    layer2_outputs(2103) <= not (a and b);
    layer2_outputs(2104) <= a and b;
    layer2_outputs(2105) <= a and b;
    layer2_outputs(2106) <= b and not a;
    layer2_outputs(2107) <= a xor b;
    layer2_outputs(2108) <= not (a and b);
    layer2_outputs(2109) <= not a or b;
    layer2_outputs(2110) <= a and not b;
    layer2_outputs(2111) <= a or b;
    layer2_outputs(2112) <= '0';
    layer2_outputs(2113) <= a or b;
    layer2_outputs(2114) <= b;
    layer2_outputs(2115) <= '0';
    layer2_outputs(2116) <= a and b;
    layer2_outputs(2117) <= not a or b;
    layer2_outputs(2118) <= '1';
    layer2_outputs(2119) <= a;
    layer2_outputs(2120) <= not b;
    layer2_outputs(2121) <= b;
    layer2_outputs(2122) <= not a or b;
    layer2_outputs(2123) <= a or b;
    layer2_outputs(2124) <= not a or b;
    layer2_outputs(2125) <= not (a and b);
    layer2_outputs(2126) <= a or b;
    layer2_outputs(2127) <= a and not b;
    layer2_outputs(2128) <= not a or b;
    layer2_outputs(2129) <= '1';
    layer2_outputs(2130) <= not (a and b);
    layer2_outputs(2131) <= not (a xor b);
    layer2_outputs(2132) <= not (a and b);
    layer2_outputs(2133) <= b;
    layer2_outputs(2134) <= not a;
    layer2_outputs(2135) <= a and not b;
    layer2_outputs(2136) <= b;
    layer2_outputs(2137) <= not a or b;
    layer2_outputs(2138) <= a and not b;
    layer2_outputs(2139) <= not (a and b);
    layer2_outputs(2140) <= not a or b;
    layer2_outputs(2141) <= not (a and b);
    layer2_outputs(2142) <= not b or a;
    layer2_outputs(2143) <= b and not a;
    layer2_outputs(2144) <= a or b;
    layer2_outputs(2145) <= a and b;
    layer2_outputs(2146) <= not a;
    layer2_outputs(2147) <= not a;
    layer2_outputs(2148) <= b and not a;
    layer2_outputs(2149) <= not a;
    layer2_outputs(2150) <= a;
    layer2_outputs(2151) <= a and b;
    layer2_outputs(2152) <= a and not b;
    layer2_outputs(2153) <= b;
    layer2_outputs(2154) <= '1';
    layer2_outputs(2155) <= not a or b;
    layer2_outputs(2156) <= not b;
    layer2_outputs(2157) <= '1';
    layer2_outputs(2158) <= not (a or b);
    layer2_outputs(2159) <= a and not b;
    layer2_outputs(2160) <= not a;
    layer2_outputs(2161) <= a and not b;
    layer2_outputs(2162) <= not a or b;
    layer2_outputs(2163) <= a or b;
    layer2_outputs(2164) <= a;
    layer2_outputs(2165) <= '1';
    layer2_outputs(2166) <= a;
    layer2_outputs(2167) <= not (a or b);
    layer2_outputs(2168) <= not (a and b);
    layer2_outputs(2169) <= b and not a;
    layer2_outputs(2170) <= '0';
    layer2_outputs(2171) <= a and not b;
    layer2_outputs(2172) <= a or b;
    layer2_outputs(2173) <= '1';
    layer2_outputs(2174) <= a and not b;
    layer2_outputs(2175) <= '1';
    layer2_outputs(2176) <= b and not a;
    layer2_outputs(2177) <= not b;
    layer2_outputs(2178) <= b;
    layer2_outputs(2179) <= a or b;
    layer2_outputs(2180) <= not (a xor b);
    layer2_outputs(2181) <= a and not b;
    layer2_outputs(2182) <= a;
    layer2_outputs(2183) <= not b;
    layer2_outputs(2184) <= b;
    layer2_outputs(2185) <= '1';
    layer2_outputs(2186) <= a and not b;
    layer2_outputs(2187) <= a xor b;
    layer2_outputs(2188) <= b;
    layer2_outputs(2189) <= b and not a;
    layer2_outputs(2190) <= a or b;
    layer2_outputs(2191) <= '0';
    layer2_outputs(2192) <= not (a or b);
    layer2_outputs(2193) <= not (a and b);
    layer2_outputs(2194) <= not (a or b);
    layer2_outputs(2195) <= not a;
    layer2_outputs(2196) <= not a;
    layer2_outputs(2197) <= a and not b;
    layer2_outputs(2198) <= b and not a;
    layer2_outputs(2199) <= a or b;
    layer2_outputs(2200) <= b and not a;
    layer2_outputs(2201) <= a xor b;
    layer2_outputs(2202) <= a and b;
    layer2_outputs(2203) <= b and not a;
    layer2_outputs(2204) <= not (a or b);
    layer2_outputs(2205) <= not b;
    layer2_outputs(2206) <= not b or a;
    layer2_outputs(2207) <= a and not b;
    layer2_outputs(2208) <= a;
    layer2_outputs(2209) <= b and not a;
    layer2_outputs(2210) <= a or b;
    layer2_outputs(2211) <= a and b;
    layer2_outputs(2212) <= '1';
    layer2_outputs(2213) <= a and b;
    layer2_outputs(2214) <= '1';
    layer2_outputs(2215) <= '0';
    layer2_outputs(2216) <= '1';
    layer2_outputs(2217) <= not (a or b);
    layer2_outputs(2218) <= not b or a;
    layer2_outputs(2219) <= a or b;
    layer2_outputs(2220) <= not b;
    layer2_outputs(2221) <= b and not a;
    layer2_outputs(2222) <= '0';
    layer2_outputs(2223) <= a and b;
    layer2_outputs(2224) <= '1';
    layer2_outputs(2225) <= b;
    layer2_outputs(2226) <= not b or a;
    layer2_outputs(2227) <= not (a or b);
    layer2_outputs(2228) <= not (a and b);
    layer2_outputs(2229) <= a;
    layer2_outputs(2230) <= a and not b;
    layer2_outputs(2231) <= a and b;
    layer2_outputs(2232) <= '1';
    layer2_outputs(2233) <= not (a and b);
    layer2_outputs(2234) <= a or b;
    layer2_outputs(2235) <= not (a and b);
    layer2_outputs(2236) <= not b or a;
    layer2_outputs(2237) <= '1';
    layer2_outputs(2238) <= '0';
    layer2_outputs(2239) <= not b or a;
    layer2_outputs(2240) <= a and not b;
    layer2_outputs(2241) <= not (a or b);
    layer2_outputs(2242) <= '1';
    layer2_outputs(2243) <= not a or b;
    layer2_outputs(2244) <= '1';
    layer2_outputs(2245) <= a or b;
    layer2_outputs(2246) <= not b or a;
    layer2_outputs(2247) <= not (a or b);
    layer2_outputs(2248) <= not a;
    layer2_outputs(2249) <= a and b;
    layer2_outputs(2250) <= '0';
    layer2_outputs(2251) <= '0';
    layer2_outputs(2252) <= b;
    layer2_outputs(2253) <= not b or a;
    layer2_outputs(2254) <= a and not b;
    layer2_outputs(2255) <= not a;
    layer2_outputs(2256) <= not a;
    layer2_outputs(2257) <= a;
    layer2_outputs(2258) <= not b or a;
    layer2_outputs(2259) <= not a or b;
    layer2_outputs(2260) <= not (a or b);
    layer2_outputs(2261) <= not a or b;
    layer2_outputs(2262) <= not (a xor b);
    layer2_outputs(2263) <= '0';
    layer2_outputs(2264) <= '1';
    layer2_outputs(2265) <= '1';
    layer2_outputs(2266) <= '1';
    layer2_outputs(2267) <= b and not a;
    layer2_outputs(2268) <= not b;
    layer2_outputs(2269) <= a or b;
    layer2_outputs(2270) <= a and b;
    layer2_outputs(2271) <= a xor b;
    layer2_outputs(2272) <= not a or b;
    layer2_outputs(2273) <= a;
    layer2_outputs(2274) <= a and b;
    layer2_outputs(2275) <= a and b;
    layer2_outputs(2276) <= a;
    layer2_outputs(2277) <= a or b;
    layer2_outputs(2278) <= not (a xor b);
    layer2_outputs(2279) <= b;
    layer2_outputs(2280) <= not a or b;
    layer2_outputs(2281) <= '0';
    layer2_outputs(2282) <= b;
    layer2_outputs(2283) <= b and not a;
    layer2_outputs(2284) <= not a or b;
    layer2_outputs(2285) <= a or b;
    layer2_outputs(2286) <= not b;
    layer2_outputs(2287) <= not b;
    layer2_outputs(2288) <= a and not b;
    layer2_outputs(2289) <= not a or b;
    layer2_outputs(2290) <= a and b;
    layer2_outputs(2291) <= b;
    layer2_outputs(2292) <= not (a and b);
    layer2_outputs(2293) <= b;
    layer2_outputs(2294) <= not (a or b);
    layer2_outputs(2295) <= a xor b;
    layer2_outputs(2296) <= b;
    layer2_outputs(2297) <= a and not b;
    layer2_outputs(2298) <= a or b;
    layer2_outputs(2299) <= not a or b;
    layer2_outputs(2300) <= not a;
    layer2_outputs(2301) <= a and not b;
    layer2_outputs(2302) <= not a or b;
    layer2_outputs(2303) <= '0';
    layer2_outputs(2304) <= a and not b;
    layer2_outputs(2305) <= not (a or b);
    layer2_outputs(2306) <= a and b;
    layer2_outputs(2307) <= b;
    layer2_outputs(2308) <= not b or a;
    layer2_outputs(2309) <= not (a xor b);
    layer2_outputs(2310) <= a;
    layer2_outputs(2311) <= not (a or b);
    layer2_outputs(2312) <= not (a or b);
    layer2_outputs(2313) <= b;
    layer2_outputs(2314) <= '0';
    layer2_outputs(2315) <= a or b;
    layer2_outputs(2316) <= b and not a;
    layer2_outputs(2317) <= '0';
    layer2_outputs(2318) <= b and not a;
    layer2_outputs(2319) <= not a or b;
    layer2_outputs(2320) <= a;
    layer2_outputs(2321) <= not a or b;
    layer2_outputs(2322) <= not b or a;
    layer2_outputs(2323) <= '1';
    layer2_outputs(2324) <= a or b;
    layer2_outputs(2325) <= '0';
    layer2_outputs(2326) <= not (a and b);
    layer2_outputs(2327) <= not b;
    layer2_outputs(2328) <= a or b;
    layer2_outputs(2329) <= a or b;
    layer2_outputs(2330) <= not b or a;
    layer2_outputs(2331) <= b;
    layer2_outputs(2332) <= not a;
    layer2_outputs(2333) <= not (a or b);
    layer2_outputs(2334) <= not b or a;
    layer2_outputs(2335) <= not a;
    layer2_outputs(2336) <= not b or a;
    layer2_outputs(2337) <= '0';
    layer2_outputs(2338) <= '0';
    layer2_outputs(2339) <= '0';
    layer2_outputs(2340) <= b and not a;
    layer2_outputs(2341) <= not b or a;
    layer2_outputs(2342) <= not a or b;
    layer2_outputs(2343) <= a and b;
    layer2_outputs(2344) <= a;
    layer2_outputs(2345) <= not (a or b);
    layer2_outputs(2346) <= b;
    layer2_outputs(2347) <= '1';
    layer2_outputs(2348) <= a;
    layer2_outputs(2349) <= '1';
    layer2_outputs(2350) <= '0';
    layer2_outputs(2351) <= '0';
    layer2_outputs(2352) <= not (a or b);
    layer2_outputs(2353) <= '1';
    layer2_outputs(2354) <= not (a or b);
    layer2_outputs(2355) <= a and not b;
    layer2_outputs(2356) <= not b or a;
    layer2_outputs(2357) <= '1';
    layer2_outputs(2358) <= a and not b;
    layer2_outputs(2359) <= a and not b;
    layer2_outputs(2360) <= '0';
    layer2_outputs(2361) <= not b or a;
    layer2_outputs(2362) <= a or b;
    layer2_outputs(2363) <= a;
    layer2_outputs(2364) <= '0';
    layer2_outputs(2365) <= not (a or b);
    layer2_outputs(2366) <= not b;
    layer2_outputs(2367) <= not a or b;
    layer2_outputs(2368) <= '1';
    layer2_outputs(2369) <= not (a or b);
    layer2_outputs(2370) <= not a or b;
    layer2_outputs(2371) <= not (a xor b);
    layer2_outputs(2372) <= a or b;
    layer2_outputs(2373) <= not (a or b);
    layer2_outputs(2374) <= not (a and b);
    layer2_outputs(2375) <= not b;
    layer2_outputs(2376) <= not (a and b);
    layer2_outputs(2377) <= not b;
    layer2_outputs(2378) <= not (a and b);
    layer2_outputs(2379) <= a xor b;
    layer2_outputs(2380) <= not b or a;
    layer2_outputs(2381) <= '0';
    layer2_outputs(2382) <= b and not a;
    layer2_outputs(2383) <= a and b;
    layer2_outputs(2384) <= '0';
    layer2_outputs(2385) <= a;
    layer2_outputs(2386) <= a and not b;
    layer2_outputs(2387) <= '1';
    layer2_outputs(2388) <= '1';
    layer2_outputs(2389) <= a;
    layer2_outputs(2390) <= not b;
    layer2_outputs(2391) <= '0';
    layer2_outputs(2392) <= a and b;
    layer2_outputs(2393) <= a and not b;
    layer2_outputs(2394) <= not a or b;
    layer2_outputs(2395) <= not (a or b);
    layer2_outputs(2396) <= a and b;
    layer2_outputs(2397) <= not (a or b);
    layer2_outputs(2398) <= not a;
    layer2_outputs(2399) <= a or b;
    layer2_outputs(2400) <= a;
    layer2_outputs(2401) <= a and not b;
    layer2_outputs(2402) <= a and b;
    layer2_outputs(2403) <= not a;
    layer2_outputs(2404) <= not a or b;
    layer2_outputs(2405) <= not a;
    layer2_outputs(2406) <= not b;
    layer2_outputs(2407) <= b and not a;
    layer2_outputs(2408) <= a;
    layer2_outputs(2409) <= '1';
    layer2_outputs(2410) <= not (a and b);
    layer2_outputs(2411) <= b;
    layer2_outputs(2412) <= not b or a;
    layer2_outputs(2413) <= b and not a;
    layer2_outputs(2414) <= not (a or b);
    layer2_outputs(2415) <= b and not a;
    layer2_outputs(2416) <= b and not a;
    layer2_outputs(2417) <= not (a and b);
    layer2_outputs(2418) <= not a or b;
    layer2_outputs(2419) <= '0';
    layer2_outputs(2420) <= not (a or b);
    layer2_outputs(2421) <= a;
    layer2_outputs(2422) <= a and not b;
    layer2_outputs(2423) <= b;
    layer2_outputs(2424) <= b;
    layer2_outputs(2425) <= b and not a;
    layer2_outputs(2426) <= not (a or b);
    layer2_outputs(2427) <= not a or b;
    layer2_outputs(2428) <= '1';
    layer2_outputs(2429) <= b and not a;
    layer2_outputs(2430) <= '1';
    layer2_outputs(2431) <= not a or b;
    layer2_outputs(2432) <= '1';
    layer2_outputs(2433) <= '0';
    layer2_outputs(2434) <= not b;
    layer2_outputs(2435) <= not (a and b);
    layer2_outputs(2436) <= not b or a;
    layer2_outputs(2437) <= not b;
    layer2_outputs(2438) <= b;
    layer2_outputs(2439) <= a;
    layer2_outputs(2440) <= '1';
    layer2_outputs(2441) <= b;
    layer2_outputs(2442) <= '1';
    layer2_outputs(2443) <= a and b;
    layer2_outputs(2444) <= '0';
    layer2_outputs(2445) <= not a;
    layer2_outputs(2446) <= b;
    layer2_outputs(2447) <= not b or a;
    layer2_outputs(2448) <= not a or b;
    layer2_outputs(2449) <= a or b;
    layer2_outputs(2450) <= not a;
    layer2_outputs(2451) <= '0';
    layer2_outputs(2452) <= '1';
    layer2_outputs(2453) <= a and b;
    layer2_outputs(2454) <= b;
    layer2_outputs(2455) <= b;
    layer2_outputs(2456) <= b;
    layer2_outputs(2457) <= a;
    layer2_outputs(2458) <= a and b;
    layer2_outputs(2459) <= not (a or b);
    layer2_outputs(2460) <= not b;
    layer2_outputs(2461) <= b;
    layer2_outputs(2462) <= a and not b;
    layer2_outputs(2463) <= not a;
    layer2_outputs(2464) <= b and not a;
    layer2_outputs(2465) <= a and b;
    layer2_outputs(2466) <= '1';
    layer2_outputs(2467) <= a or b;
    layer2_outputs(2468) <= not (a or b);
    layer2_outputs(2469) <= not (a and b);
    layer2_outputs(2470) <= not (a and b);
    layer2_outputs(2471) <= '0';
    layer2_outputs(2472) <= not a or b;
    layer2_outputs(2473) <= not b;
    layer2_outputs(2474) <= a and not b;
    layer2_outputs(2475) <= not b or a;
    layer2_outputs(2476) <= '0';
    layer2_outputs(2477) <= not a;
    layer2_outputs(2478) <= b and not a;
    layer2_outputs(2479) <= '1';
    layer2_outputs(2480) <= not (a and b);
    layer2_outputs(2481) <= not a or b;
    layer2_outputs(2482) <= not a or b;
    layer2_outputs(2483) <= a and b;
    layer2_outputs(2484) <= '0';
    layer2_outputs(2485) <= b and not a;
    layer2_outputs(2486) <= not b or a;
    layer2_outputs(2487) <= not (a or b);
    layer2_outputs(2488) <= '1';
    layer2_outputs(2489) <= a and b;
    layer2_outputs(2490) <= b and not a;
    layer2_outputs(2491) <= not (a and b);
    layer2_outputs(2492) <= b and not a;
    layer2_outputs(2493) <= b;
    layer2_outputs(2494) <= a;
    layer2_outputs(2495) <= not b or a;
    layer2_outputs(2496) <= not (a xor b);
    layer2_outputs(2497) <= a;
    layer2_outputs(2498) <= b;
    layer2_outputs(2499) <= a and not b;
    layer2_outputs(2500) <= a or b;
    layer2_outputs(2501) <= not (a or b);
    layer2_outputs(2502) <= a and b;
    layer2_outputs(2503) <= '1';
    layer2_outputs(2504) <= '1';
    layer2_outputs(2505) <= not b or a;
    layer2_outputs(2506) <= not (a or b);
    layer2_outputs(2507) <= '1';
    layer2_outputs(2508) <= not (a xor b);
    layer2_outputs(2509) <= a or b;
    layer2_outputs(2510) <= not (a or b);
    layer2_outputs(2511) <= b and not a;
    layer2_outputs(2512) <= not b;
    layer2_outputs(2513) <= '1';
    layer2_outputs(2514) <= not (a or b);
    layer2_outputs(2515) <= a and not b;
    layer2_outputs(2516) <= not b;
    layer2_outputs(2517) <= '1';
    layer2_outputs(2518) <= b;
    layer2_outputs(2519) <= not a or b;
    layer2_outputs(2520) <= '1';
    layer2_outputs(2521) <= not (a xor b);
    layer2_outputs(2522) <= not a or b;
    layer2_outputs(2523) <= a or b;
    layer2_outputs(2524) <= b and not a;
    layer2_outputs(2525) <= a or b;
    layer2_outputs(2526) <= a and not b;
    layer2_outputs(2527) <= '0';
    layer2_outputs(2528) <= a and b;
    layer2_outputs(2529) <= not a;
    layer2_outputs(2530) <= not a;
    layer2_outputs(2531) <= '0';
    layer2_outputs(2532) <= not b or a;
    layer2_outputs(2533) <= not b or a;
    layer2_outputs(2534) <= not (a and b);
    layer2_outputs(2535) <= not a or b;
    layer2_outputs(2536) <= not b;
    layer2_outputs(2537) <= a and not b;
    layer2_outputs(2538) <= not (a and b);
    layer2_outputs(2539) <= a or b;
    layer2_outputs(2540) <= not b or a;
    layer2_outputs(2541) <= not b;
    layer2_outputs(2542) <= not (a xor b);
    layer2_outputs(2543) <= a or b;
    layer2_outputs(2544) <= a and not b;
    layer2_outputs(2545) <= not a or b;
    layer2_outputs(2546) <= '0';
    layer2_outputs(2547) <= not a or b;
    layer2_outputs(2548) <= not b or a;
    layer2_outputs(2549) <= not b or a;
    layer2_outputs(2550) <= '1';
    layer2_outputs(2551) <= not a or b;
    layer2_outputs(2552) <= '1';
    layer2_outputs(2553) <= '1';
    layer2_outputs(2554) <= '1';
    layer2_outputs(2555) <= not b;
    layer2_outputs(2556) <= not b;
    layer2_outputs(2557) <= '1';
    layer2_outputs(2558) <= not a or b;
    layer2_outputs(2559) <= not a or b;
    layer2_outputs(2560) <= a and b;
    layer2_outputs(2561) <= '1';
    layer2_outputs(2562) <= '1';
    layer2_outputs(2563) <= a and b;
    layer2_outputs(2564) <= a and b;
    layer2_outputs(2565) <= b and not a;
    layer2_outputs(2566) <= '1';
    layer2_outputs(2567) <= not b or a;
    layer2_outputs(2568) <= not a;
    layer2_outputs(2569) <= a and not b;
    layer2_outputs(2570) <= a xor b;
    layer2_outputs(2571) <= b and not a;
    layer2_outputs(2572) <= not b or a;
    layer2_outputs(2573) <= a or b;
    layer2_outputs(2574) <= '0';
    layer2_outputs(2575) <= not a;
    layer2_outputs(2576) <= a;
    layer2_outputs(2577) <= a and b;
    layer2_outputs(2578) <= a and b;
    layer2_outputs(2579) <= a and b;
    layer2_outputs(2580) <= '1';
    layer2_outputs(2581) <= not b or a;
    layer2_outputs(2582) <= not b;
    layer2_outputs(2583) <= a and b;
    layer2_outputs(2584) <= b;
    layer2_outputs(2585) <= a and b;
    layer2_outputs(2586) <= not a or b;
    layer2_outputs(2587) <= not a or b;
    layer2_outputs(2588) <= a or b;
    layer2_outputs(2589) <= '0';
    layer2_outputs(2590) <= '0';
    layer2_outputs(2591) <= not b;
    layer2_outputs(2592) <= not (a and b);
    layer2_outputs(2593) <= '0';
    layer2_outputs(2594) <= not a;
    layer2_outputs(2595) <= not a or b;
    layer2_outputs(2596) <= b and not a;
    layer2_outputs(2597) <= a;
    layer2_outputs(2598) <= '1';
    layer2_outputs(2599) <= not (a xor b);
    layer2_outputs(2600) <= not a or b;
    layer2_outputs(2601) <= a and b;
    layer2_outputs(2602) <= not a or b;
    layer2_outputs(2603) <= a and b;
    layer2_outputs(2604) <= b;
    layer2_outputs(2605) <= b and not a;
    layer2_outputs(2606) <= not a;
    layer2_outputs(2607) <= b;
    layer2_outputs(2608) <= '1';
    layer2_outputs(2609) <= a or b;
    layer2_outputs(2610) <= a and b;
    layer2_outputs(2611) <= a;
    layer2_outputs(2612) <= a and b;
    layer2_outputs(2613) <= not (a or b);
    layer2_outputs(2614) <= a and b;
    layer2_outputs(2615) <= not (a and b);
    layer2_outputs(2616) <= a xor b;
    layer2_outputs(2617) <= '0';
    layer2_outputs(2618) <= a or b;
    layer2_outputs(2619) <= not (a or b);
    layer2_outputs(2620) <= not (a or b);
    layer2_outputs(2621) <= a and b;
    layer2_outputs(2622) <= not a or b;
    layer2_outputs(2623) <= not (a or b);
    layer2_outputs(2624) <= b and not a;
    layer2_outputs(2625) <= not b;
    layer2_outputs(2626) <= a or b;
    layer2_outputs(2627) <= '1';
    layer2_outputs(2628) <= b;
    layer2_outputs(2629) <= '1';
    layer2_outputs(2630) <= not (a and b);
    layer2_outputs(2631) <= a xor b;
    layer2_outputs(2632) <= '1';
    layer2_outputs(2633) <= b;
    layer2_outputs(2634) <= a;
    layer2_outputs(2635) <= not a or b;
    layer2_outputs(2636) <= not (a or b);
    layer2_outputs(2637) <= b and not a;
    layer2_outputs(2638) <= a and b;
    layer2_outputs(2639) <= a and not b;
    layer2_outputs(2640) <= a and not b;
    layer2_outputs(2641) <= a and not b;
    layer2_outputs(2642) <= a and b;
    layer2_outputs(2643) <= a or b;
    layer2_outputs(2644) <= a;
    layer2_outputs(2645) <= b and not a;
    layer2_outputs(2646) <= '1';
    layer2_outputs(2647) <= b and not a;
    layer2_outputs(2648) <= not b or a;
    layer2_outputs(2649) <= a;
    layer2_outputs(2650) <= not a;
    layer2_outputs(2651) <= a or b;
    layer2_outputs(2652) <= b;
    layer2_outputs(2653) <= a xor b;
    layer2_outputs(2654) <= a or b;
    layer2_outputs(2655) <= a and b;
    layer2_outputs(2656) <= not (a xor b);
    layer2_outputs(2657) <= a and not b;
    layer2_outputs(2658) <= not b;
    layer2_outputs(2659) <= not b or a;
    layer2_outputs(2660) <= a or b;
    layer2_outputs(2661) <= not b or a;
    layer2_outputs(2662) <= '1';
    layer2_outputs(2663) <= not a;
    layer2_outputs(2664) <= a and not b;
    layer2_outputs(2665) <= not a or b;
    layer2_outputs(2666) <= '0';
    layer2_outputs(2667) <= not (a and b);
    layer2_outputs(2668) <= b;
    layer2_outputs(2669) <= b;
    layer2_outputs(2670) <= not b;
    layer2_outputs(2671) <= '0';
    layer2_outputs(2672) <= not a;
    layer2_outputs(2673) <= a or b;
    layer2_outputs(2674) <= not a or b;
    layer2_outputs(2675) <= '1';
    layer2_outputs(2676) <= '1';
    layer2_outputs(2677) <= not b or a;
    layer2_outputs(2678) <= b;
    layer2_outputs(2679) <= not (a or b);
    layer2_outputs(2680) <= '1';
    layer2_outputs(2681) <= not a or b;
    layer2_outputs(2682) <= a and b;
    layer2_outputs(2683) <= a or b;
    layer2_outputs(2684) <= not a;
    layer2_outputs(2685) <= b and not a;
    layer2_outputs(2686) <= not (a and b);
    layer2_outputs(2687) <= not b;
    layer2_outputs(2688) <= a;
    layer2_outputs(2689) <= b and not a;
    layer2_outputs(2690) <= not a;
    layer2_outputs(2691) <= '0';
    layer2_outputs(2692) <= '1';
    layer2_outputs(2693) <= not (a or b);
    layer2_outputs(2694) <= not (a or b);
    layer2_outputs(2695) <= a or b;
    layer2_outputs(2696) <= a and not b;
    layer2_outputs(2697) <= a and not b;
    layer2_outputs(2698) <= not (a or b);
    layer2_outputs(2699) <= not (a or b);
    layer2_outputs(2700) <= not (a or b);
    layer2_outputs(2701) <= b and not a;
    layer2_outputs(2702) <= not (a or b);
    layer2_outputs(2703) <= not a or b;
    layer2_outputs(2704) <= not a;
    layer2_outputs(2705) <= not (a or b);
    layer2_outputs(2706) <= not b or a;
    layer2_outputs(2707) <= a and b;
    layer2_outputs(2708) <= '0';
    layer2_outputs(2709) <= a and b;
    layer2_outputs(2710) <= not (a or b);
    layer2_outputs(2711) <= '0';
    layer2_outputs(2712) <= a;
    layer2_outputs(2713) <= '1';
    layer2_outputs(2714) <= not (a xor b);
    layer2_outputs(2715) <= a and not b;
    layer2_outputs(2716) <= not (a or b);
    layer2_outputs(2717) <= a;
    layer2_outputs(2718) <= a and b;
    layer2_outputs(2719) <= not (a or b);
    layer2_outputs(2720) <= a and b;
    layer2_outputs(2721) <= not b or a;
    layer2_outputs(2722) <= a and b;
    layer2_outputs(2723) <= b and not a;
    layer2_outputs(2724) <= not b;
    layer2_outputs(2725) <= b;
    layer2_outputs(2726) <= not a or b;
    layer2_outputs(2727) <= not a or b;
    layer2_outputs(2728) <= not a;
    layer2_outputs(2729) <= not (a and b);
    layer2_outputs(2730) <= not a or b;
    layer2_outputs(2731) <= not b;
    layer2_outputs(2732) <= not a or b;
    layer2_outputs(2733) <= '0';
    layer2_outputs(2734) <= '1';
    layer2_outputs(2735) <= not b;
    layer2_outputs(2736) <= a and not b;
    layer2_outputs(2737) <= not a;
    layer2_outputs(2738) <= '0';
    layer2_outputs(2739) <= a or b;
    layer2_outputs(2740) <= not a or b;
    layer2_outputs(2741) <= a and b;
    layer2_outputs(2742) <= not b;
    layer2_outputs(2743) <= not a or b;
    layer2_outputs(2744) <= b and not a;
    layer2_outputs(2745) <= not b;
    layer2_outputs(2746) <= not (a or b);
    layer2_outputs(2747) <= '0';
    layer2_outputs(2748) <= not (a and b);
    layer2_outputs(2749) <= not a;
    layer2_outputs(2750) <= not a or b;
    layer2_outputs(2751) <= a or b;
    layer2_outputs(2752) <= not (a or b);
    layer2_outputs(2753) <= not b;
    layer2_outputs(2754) <= a or b;
    layer2_outputs(2755) <= '0';
    layer2_outputs(2756) <= '0';
    layer2_outputs(2757) <= a and not b;
    layer2_outputs(2758) <= not a;
    layer2_outputs(2759) <= '0';
    layer2_outputs(2760) <= not (a and b);
    layer2_outputs(2761) <= b;
    layer2_outputs(2762) <= not a;
    layer2_outputs(2763) <= '1';
    layer2_outputs(2764) <= a and b;
    layer2_outputs(2765) <= not b or a;
    layer2_outputs(2766) <= not b or a;
    layer2_outputs(2767) <= not b;
    layer2_outputs(2768) <= not (a or b);
    layer2_outputs(2769) <= not (a or b);
    layer2_outputs(2770) <= '0';
    layer2_outputs(2771) <= b;
    layer2_outputs(2772) <= not (a xor b);
    layer2_outputs(2773) <= '0';
    layer2_outputs(2774) <= a and b;
    layer2_outputs(2775) <= b and not a;
    layer2_outputs(2776) <= a and not b;
    layer2_outputs(2777) <= b and not a;
    layer2_outputs(2778) <= not a;
    layer2_outputs(2779) <= not a or b;
    layer2_outputs(2780) <= not a or b;
    layer2_outputs(2781) <= a and not b;
    layer2_outputs(2782) <= b;
    layer2_outputs(2783) <= not (a and b);
    layer2_outputs(2784) <= not (a and b);
    layer2_outputs(2785) <= not a or b;
    layer2_outputs(2786) <= not (a and b);
    layer2_outputs(2787) <= a;
    layer2_outputs(2788) <= b and not a;
    layer2_outputs(2789) <= a and b;
    layer2_outputs(2790) <= not a or b;
    layer2_outputs(2791) <= '1';
    layer2_outputs(2792) <= not a or b;
    layer2_outputs(2793) <= '1';
    layer2_outputs(2794) <= b and not a;
    layer2_outputs(2795) <= not a;
    layer2_outputs(2796) <= a or b;
    layer2_outputs(2797) <= a and b;
    layer2_outputs(2798) <= a;
    layer2_outputs(2799) <= a and b;
    layer2_outputs(2800) <= '0';
    layer2_outputs(2801) <= a and not b;
    layer2_outputs(2802) <= not (a and b);
    layer2_outputs(2803) <= not b;
    layer2_outputs(2804) <= a or b;
    layer2_outputs(2805) <= a and not b;
    layer2_outputs(2806) <= a;
    layer2_outputs(2807) <= '0';
    layer2_outputs(2808) <= '0';
    layer2_outputs(2809) <= not a or b;
    layer2_outputs(2810) <= a and b;
    layer2_outputs(2811) <= not a or b;
    layer2_outputs(2812) <= a and not b;
    layer2_outputs(2813) <= a and not b;
    layer2_outputs(2814) <= a;
    layer2_outputs(2815) <= b;
    layer2_outputs(2816) <= '0';
    layer2_outputs(2817) <= a and not b;
    layer2_outputs(2818) <= not b or a;
    layer2_outputs(2819) <= '1';
    layer2_outputs(2820) <= a;
    layer2_outputs(2821) <= b and not a;
    layer2_outputs(2822) <= not (a and b);
    layer2_outputs(2823) <= '1';
    layer2_outputs(2824) <= not b;
    layer2_outputs(2825) <= '1';
    layer2_outputs(2826) <= '0';
    layer2_outputs(2827) <= a or b;
    layer2_outputs(2828) <= not b;
    layer2_outputs(2829) <= not a;
    layer2_outputs(2830) <= not b or a;
    layer2_outputs(2831) <= a;
    layer2_outputs(2832) <= not (a or b);
    layer2_outputs(2833) <= not b;
    layer2_outputs(2834) <= not b or a;
    layer2_outputs(2835) <= a and not b;
    layer2_outputs(2836) <= '0';
    layer2_outputs(2837) <= not b;
    layer2_outputs(2838) <= a and not b;
    layer2_outputs(2839) <= not b;
    layer2_outputs(2840) <= a and not b;
    layer2_outputs(2841) <= '1';
    layer2_outputs(2842) <= a or b;
    layer2_outputs(2843) <= not a;
    layer2_outputs(2844) <= b and not a;
    layer2_outputs(2845) <= not b;
    layer2_outputs(2846) <= a and not b;
    layer2_outputs(2847) <= b and not a;
    layer2_outputs(2848) <= a and b;
    layer2_outputs(2849) <= b;
    layer2_outputs(2850) <= a or b;
    layer2_outputs(2851) <= not a or b;
    layer2_outputs(2852) <= not (a or b);
    layer2_outputs(2853) <= not a;
    layer2_outputs(2854) <= not b;
    layer2_outputs(2855) <= a and b;
    layer2_outputs(2856) <= b;
    layer2_outputs(2857) <= a and b;
    layer2_outputs(2858) <= '0';
    layer2_outputs(2859) <= '1';
    layer2_outputs(2860) <= b;
    layer2_outputs(2861) <= '0';
    layer2_outputs(2862) <= a or b;
    layer2_outputs(2863) <= b and not a;
    layer2_outputs(2864) <= not a or b;
    layer2_outputs(2865) <= not (a or b);
    layer2_outputs(2866) <= not b or a;
    layer2_outputs(2867) <= a;
    layer2_outputs(2868) <= a;
    layer2_outputs(2869) <= not a;
    layer2_outputs(2870) <= not a;
    layer2_outputs(2871) <= a or b;
    layer2_outputs(2872) <= '1';
    layer2_outputs(2873) <= not b or a;
    layer2_outputs(2874) <= b and not a;
    layer2_outputs(2875) <= not (a xor b);
    layer2_outputs(2876) <= not b;
    layer2_outputs(2877) <= a;
    layer2_outputs(2878) <= a and b;
    layer2_outputs(2879) <= '0';
    layer2_outputs(2880) <= not (a and b);
    layer2_outputs(2881) <= b;
    layer2_outputs(2882) <= not a;
    layer2_outputs(2883) <= not b or a;
    layer2_outputs(2884) <= not (a or b);
    layer2_outputs(2885) <= b and not a;
    layer2_outputs(2886) <= b and not a;
    layer2_outputs(2887) <= a or b;
    layer2_outputs(2888) <= '1';
    layer2_outputs(2889) <= a or b;
    layer2_outputs(2890) <= not (a and b);
    layer2_outputs(2891) <= not (a or b);
    layer2_outputs(2892) <= not a or b;
    layer2_outputs(2893) <= a or b;
    layer2_outputs(2894) <= not a;
    layer2_outputs(2895) <= not (a or b);
    layer2_outputs(2896) <= a and b;
    layer2_outputs(2897) <= '0';
    layer2_outputs(2898) <= not a;
    layer2_outputs(2899) <= a and not b;
    layer2_outputs(2900) <= not a or b;
    layer2_outputs(2901) <= not a;
    layer2_outputs(2902) <= a and not b;
    layer2_outputs(2903) <= a and b;
    layer2_outputs(2904) <= not b;
    layer2_outputs(2905) <= a or b;
    layer2_outputs(2906) <= a and not b;
    layer2_outputs(2907) <= b and not a;
    layer2_outputs(2908) <= '1';
    layer2_outputs(2909) <= '0';
    layer2_outputs(2910) <= b and not a;
    layer2_outputs(2911) <= not (a and b);
    layer2_outputs(2912) <= not a;
    layer2_outputs(2913) <= a;
    layer2_outputs(2914) <= b and not a;
    layer2_outputs(2915) <= not a or b;
    layer2_outputs(2916) <= '1';
    layer2_outputs(2917) <= not b or a;
    layer2_outputs(2918) <= not (a or b);
    layer2_outputs(2919) <= a or b;
    layer2_outputs(2920) <= a or b;
    layer2_outputs(2921) <= not b or a;
    layer2_outputs(2922) <= not b;
    layer2_outputs(2923) <= not a;
    layer2_outputs(2924) <= not a or b;
    layer2_outputs(2925) <= b and not a;
    layer2_outputs(2926) <= a and b;
    layer2_outputs(2927) <= not (a and b);
    layer2_outputs(2928) <= '0';
    layer2_outputs(2929) <= b and not a;
    layer2_outputs(2930) <= not (a or b);
    layer2_outputs(2931) <= b;
    layer2_outputs(2932) <= '0';
    layer2_outputs(2933) <= a;
    layer2_outputs(2934) <= b;
    layer2_outputs(2935) <= a;
    layer2_outputs(2936) <= a and not b;
    layer2_outputs(2937) <= not b;
    layer2_outputs(2938) <= '0';
    layer2_outputs(2939) <= '1';
    layer2_outputs(2940) <= a;
    layer2_outputs(2941) <= not a;
    layer2_outputs(2942) <= not (a or b);
    layer2_outputs(2943) <= '0';
    layer2_outputs(2944) <= a or b;
    layer2_outputs(2945) <= b;
    layer2_outputs(2946) <= b;
    layer2_outputs(2947) <= a and b;
    layer2_outputs(2948) <= not a;
    layer2_outputs(2949) <= a;
    layer2_outputs(2950) <= a and b;
    layer2_outputs(2951) <= not a or b;
    layer2_outputs(2952) <= '0';
    layer2_outputs(2953) <= a or b;
    layer2_outputs(2954) <= not (a or b);
    layer2_outputs(2955) <= '0';
    layer2_outputs(2956) <= not (a or b);
    layer2_outputs(2957) <= not (a or b);
    layer2_outputs(2958) <= a and not b;
    layer2_outputs(2959) <= not a;
    layer2_outputs(2960) <= b;
    layer2_outputs(2961) <= a xor b;
    layer2_outputs(2962) <= not a or b;
    layer2_outputs(2963) <= not b;
    layer2_outputs(2964) <= not b;
    layer2_outputs(2965) <= not b or a;
    layer2_outputs(2966) <= a and b;
    layer2_outputs(2967) <= '0';
    layer2_outputs(2968) <= a and b;
    layer2_outputs(2969) <= b;
    layer2_outputs(2970) <= not a;
    layer2_outputs(2971) <= b;
    layer2_outputs(2972) <= not b or a;
    layer2_outputs(2973) <= a or b;
    layer2_outputs(2974) <= not (a or b);
    layer2_outputs(2975) <= '0';
    layer2_outputs(2976) <= not (a or b);
    layer2_outputs(2977) <= not (a xor b);
    layer2_outputs(2978) <= b and not a;
    layer2_outputs(2979) <= '0';
    layer2_outputs(2980) <= b;
    layer2_outputs(2981) <= b;
    layer2_outputs(2982) <= a;
    layer2_outputs(2983) <= not a;
    layer2_outputs(2984) <= not b;
    layer2_outputs(2985) <= a and not b;
    layer2_outputs(2986) <= not b or a;
    layer2_outputs(2987) <= not a;
    layer2_outputs(2988) <= b and not a;
    layer2_outputs(2989) <= a or b;
    layer2_outputs(2990) <= not (a and b);
    layer2_outputs(2991) <= '1';
    layer2_outputs(2992) <= not b or a;
    layer2_outputs(2993) <= a or b;
    layer2_outputs(2994) <= a;
    layer2_outputs(2995) <= b;
    layer2_outputs(2996) <= not b;
    layer2_outputs(2997) <= '0';
    layer2_outputs(2998) <= a and not b;
    layer2_outputs(2999) <= a or b;
    layer2_outputs(3000) <= '1';
    layer2_outputs(3001) <= not b or a;
    layer2_outputs(3002) <= '1';
    layer2_outputs(3003) <= a and b;
    layer2_outputs(3004) <= not b or a;
    layer2_outputs(3005) <= '1';
    layer2_outputs(3006) <= a;
    layer2_outputs(3007) <= not (a and b);
    layer2_outputs(3008) <= not (a or b);
    layer2_outputs(3009) <= a and not b;
    layer2_outputs(3010) <= b and not a;
    layer2_outputs(3011) <= a or b;
    layer2_outputs(3012) <= not b or a;
    layer2_outputs(3013) <= b and not a;
    layer2_outputs(3014) <= b;
    layer2_outputs(3015) <= not a;
    layer2_outputs(3016) <= not (a or b);
    layer2_outputs(3017) <= not a;
    layer2_outputs(3018) <= not (a xor b);
    layer2_outputs(3019) <= not b;
    layer2_outputs(3020) <= '0';
    layer2_outputs(3021) <= '1';
    layer2_outputs(3022) <= '1';
    layer2_outputs(3023) <= b;
    layer2_outputs(3024) <= a;
    layer2_outputs(3025) <= a and b;
    layer2_outputs(3026) <= b and not a;
    layer2_outputs(3027) <= not (a xor b);
    layer2_outputs(3028) <= not a or b;
    layer2_outputs(3029) <= b and not a;
    layer2_outputs(3030) <= a and not b;
    layer2_outputs(3031) <= not b;
    layer2_outputs(3032) <= not (a and b);
    layer2_outputs(3033) <= '1';
    layer2_outputs(3034) <= a and b;
    layer2_outputs(3035) <= not (a or b);
    layer2_outputs(3036) <= a;
    layer2_outputs(3037) <= not a or b;
    layer2_outputs(3038) <= a;
    layer2_outputs(3039) <= not b or a;
    layer2_outputs(3040) <= not (a xor b);
    layer2_outputs(3041) <= not a or b;
    layer2_outputs(3042) <= not b;
    layer2_outputs(3043) <= '0';
    layer2_outputs(3044) <= b and not a;
    layer2_outputs(3045) <= a or b;
    layer2_outputs(3046) <= '0';
    layer2_outputs(3047) <= not a or b;
    layer2_outputs(3048) <= '0';
    layer2_outputs(3049) <= not b;
    layer2_outputs(3050) <= not b;
    layer2_outputs(3051) <= b;
    layer2_outputs(3052) <= '0';
    layer2_outputs(3053) <= a and b;
    layer2_outputs(3054) <= not (a and b);
    layer2_outputs(3055) <= a or b;
    layer2_outputs(3056) <= not a or b;
    layer2_outputs(3057) <= '0';
    layer2_outputs(3058) <= a or b;
    layer2_outputs(3059) <= '1';
    layer2_outputs(3060) <= a or b;
    layer2_outputs(3061) <= b and not a;
    layer2_outputs(3062) <= a and not b;
    layer2_outputs(3063) <= not b or a;
    layer2_outputs(3064) <= not (a or b);
    layer2_outputs(3065) <= '0';
    layer2_outputs(3066) <= '1';
    layer2_outputs(3067) <= a and not b;
    layer2_outputs(3068) <= not a or b;
    layer2_outputs(3069) <= a and not b;
    layer2_outputs(3070) <= '0';
    layer2_outputs(3071) <= not (a or b);
    layer2_outputs(3072) <= not a or b;
    layer2_outputs(3073) <= not b;
    layer2_outputs(3074) <= a or b;
    layer2_outputs(3075) <= '1';
    layer2_outputs(3076) <= '0';
    layer2_outputs(3077) <= b and not a;
    layer2_outputs(3078) <= '0';
    layer2_outputs(3079) <= '1';
    layer2_outputs(3080) <= a and b;
    layer2_outputs(3081) <= not (a and b);
    layer2_outputs(3082) <= a or b;
    layer2_outputs(3083) <= not a or b;
    layer2_outputs(3084) <= a or b;
    layer2_outputs(3085) <= a and b;
    layer2_outputs(3086) <= '1';
    layer2_outputs(3087) <= '0';
    layer2_outputs(3088) <= '1';
    layer2_outputs(3089) <= '0';
    layer2_outputs(3090) <= not a or b;
    layer2_outputs(3091) <= not b;
    layer2_outputs(3092) <= not (a or b);
    layer2_outputs(3093) <= '0';
    layer2_outputs(3094) <= a;
    layer2_outputs(3095) <= a;
    layer2_outputs(3096) <= not (a or b);
    layer2_outputs(3097) <= not a or b;
    layer2_outputs(3098) <= not (a or b);
    layer2_outputs(3099) <= a;
    layer2_outputs(3100) <= b and not a;
    layer2_outputs(3101) <= a;
    layer2_outputs(3102) <= '1';
    layer2_outputs(3103) <= not (a and b);
    layer2_outputs(3104) <= not a;
    layer2_outputs(3105) <= a or b;
    layer2_outputs(3106) <= a and b;
    layer2_outputs(3107) <= b;
    layer2_outputs(3108) <= '0';
    layer2_outputs(3109) <= b and not a;
    layer2_outputs(3110) <= not (a and b);
    layer2_outputs(3111) <= not a;
    layer2_outputs(3112) <= not b;
    layer2_outputs(3113) <= '0';
    layer2_outputs(3114) <= '1';
    layer2_outputs(3115) <= not (a or b);
    layer2_outputs(3116) <= a and b;
    layer2_outputs(3117) <= not a or b;
    layer2_outputs(3118) <= not b or a;
    layer2_outputs(3119) <= '0';
    layer2_outputs(3120) <= not (a and b);
    layer2_outputs(3121) <= a or b;
    layer2_outputs(3122) <= '0';
    layer2_outputs(3123) <= not b or a;
    layer2_outputs(3124) <= not (a or b);
    layer2_outputs(3125) <= a and not b;
    layer2_outputs(3126) <= '1';
    layer2_outputs(3127) <= not b or a;
    layer2_outputs(3128) <= '1';
    layer2_outputs(3129) <= b and not a;
    layer2_outputs(3130) <= not b or a;
    layer2_outputs(3131) <= a and not b;
    layer2_outputs(3132) <= not (a and b);
    layer2_outputs(3133) <= a;
    layer2_outputs(3134) <= not b;
    layer2_outputs(3135) <= a and b;
    layer2_outputs(3136) <= b and not a;
    layer2_outputs(3137) <= not (a or b);
    layer2_outputs(3138) <= b;
    layer2_outputs(3139) <= not b or a;
    layer2_outputs(3140) <= not b;
    layer2_outputs(3141) <= not a or b;
    layer2_outputs(3142) <= '0';
    layer2_outputs(3143) <= not a or b;
    layer2_outputs(3144) <= a xor b;
    layer2_outputs(3145) <= not (a and b);
    layer2_outputs(3146) <= a or b;
    layer2_outputs(3147) <= b;
    layer2_outputs(3148) <= not a;
    layer2_outputs(3149) <= a or b;
    layer2_outputs(3150) <= '0';
    layer2_outputs(3151) <= not a;
    layer2_outputs(3152) <= b;
    layer2_outputs(3153) <= not a;
    layer2_outputs(3154) <= '0';
    layer2_outputs(3155) <= '0';
    layer2_outputs(3156) <= a and b;
    layer2_outputs(3157) <= '0';
    layer2_outputs(3158) <= not a;
    layer2_outputs(3159) <= not a;
    layer2_outputs(3160) <= '1';
    layer2_outputs(3161) <= a xor b;
    layer2_outputs(3162) <= a or b;
    layer2_outputs(3163) <= not b;
    layer2_outputs(3164) <= a and b;
    layer2_outputs(3165) <= a and not b;
    layer2_outputs(3166) <= not b or a;
    layer2_outputs(3167) <= a or b;
    layer2_outputs(3168) <= b and not a;
    layer2_outputs(3169) <= b and not a;
    layer2_outputs(3170) <= a and not b;
    layer2_outputs(3171) <= a;
    layer2_outputs(3172) <= b;
    layer2_outputs(3173) <= not a or b;
    layer2_outputs(3174) <= '1';
    layer2_outputs(3175) <= not a or b;
    layer2_outputs(3176) <= a and not b;
    layer2_outputs(3177) <= not a;
    layer2_outputs(3178) <= '1';
    layer2_outputs(3179) <= b;
    layer2_outputs(3180) <= not b or a;
    layer2_outputs(3181) <= a and b;
    layer2_outputs(3182) <= not (a and b);
    layer2_outputs(3183) <= not (a xor b);
    layer2_outputs(3184) <= '1';
    layer2_outputs(3185) <= not (a or b);
    layer2_outputs(3186) <= not (a and b);
    layer2_outputs(3187) <= a or b;
    layer2_outputs(3188) <= '1';
    layer2_outputs(3189) <= a;
    layer2_outputs(3190) <= a and not b;
    layer2_outputs(3191) <= a;
    layer2_outputs(3192) <= a and b;
    layer2_outputs(3193) <= not (a or b);
    layer2_outputs(3194) <= a;
    layer2_outputs(3195) <= not b or a;
    layer2_outputs(3196) <= a and not b;
    layer2_outputs(3197) <= '1';
    layer2_outputs(3198) <= a and b;
    layer2_outputs(3199) <= '0';
    layer2_outputs(3200) <= '0';
    layer2_outputs(3201) <= not (a or b);
    layer2_outputs(3202) <= b;
    layer2_outputs(3203) <= not b or a;
    layer2_outputs(3204) <= not (a xor b);
    layer2_outputs(3205) <= '1';
    layer2_outputs(3206) <= a and not b;
    layer2_outputs(3207) <= not b;
    layer2_outputs(3208) <= not (a xor b);
    layer2_outputs(3209) <= not a or b;
    layer2_outputs(3210) <= a;
    layer2_outputs(3211) <= b;
    layer2_outputs(3212) <= '1';
    layer2_outputs(3213) <= a or b;
    layer2_outputs(3214) <= a;
    layer2_outputs(3215) <= not (a and b);
    layer2_outputs(3216) <= '0';
    layer2_outputs(3217) <= a and b;
    layer2_outputs(3218) <= a or b;
    layer2_outputs(3219) <= not a;
    layer2_outputs(3220) <= a or b;
    layer2_outputs(3221) <= a xor b;
    layer2_outputs(3222) <= b and not a;
    layer2_outputs(3223) <= a and b;
    layer2_outputs(3224) <= '1';
    layer2_outputs(3225) <= '1';
    layer2_outputs(3226) <= not b;
    layer2_outputs(3227) <= b;
    layer2_outputs(3228) <= b;
    layer2_outputs(3229) <= not b or a;
    layer2_outputs(3230) <= b and not a;
    layer2_outputs(3231) <= a and b;
    layer2_outputs(3232) <= not b or a;
    layer2_outputs(3233) <= b and not a;
    layer2_outputs(3234) <= not (a or b);
    layer2_outputs(3235) <= a and not b;
    layer2_outputs(3236) <= '1';
    layer2_outputs(3237) <= '1';
    layer2_outputs(3238) <= b;
    layer2_outputs(3239) <= a;
    layer2_outputs(3240) <= b and not a;
    layer2_outputs(3241) <= not a or b;
    layer2_outputs(3242) <= a or b;
    layer2_outputs(3243) <= '0';
    layer2_outputs(3244) <= b;
    layer2_outputs(3245) <= a and b;
    layer2_outputs(3246) <= b and not a;
    layer2_outputs(3247) <= a;
    layer2_outputs(3248) <= a or b;
    layer2_outputs(3249) <= not b;
    layer2_outputs(3250) <= not (a or b);
    layer2_outputs(3251) <= a and not b;
    layer2_outputs(3252) <= not (a or b);
    layer2_outputs(3253) <= not a;
    layer2_outputs(3254) <= a and not b;
    layer2_outputs(3255) <= not b;
    layer2_outputs(3256) <= not (a and b);
    layer2_outputs(3257) <= '0';
    layer2_outputs(3258) <= not b;
    layer2_outputs(3259) <= not a or b;
    layer2_outputs(3260) <= not b;
    layer2_outputs(3261) <= not a;
    layer2_outputs(3262) <= not b or a;
    layer2_outputs(3263) <= not a;
    layer2_outputs(3264) <= b;
    layer2_outputs(3265) <= not (a and b);
    layer2_outputs(3266) <= b;
    layer2_outputs(3267) <= not (a or b);
    layer2_outputs(3268) <= '0';
    layer2_outputs(3269) <= b;
    layer2_outputs(3270) <= not a or b;
    layer2_outputs(3271) <= a or b;
    layer2_outputs(3272) <= a or b;
    layer2_outputs(3273) <= a;
    layer2_outputs(3274) <= a or b;
    layer2_outputs(3275) <= not a or b;
    layer2_outputs(3276) <= b and not a;
    layer2_outputs(3277) <= not (a and b);
    layer2_outputs(3278) <= '1';
    layer2_outputs(3279) <= a and b;
    layer2_outputs(3280) <= a or b;
    layer2_outputs(3281) <= not a or b;
    layer2_outputs(3282) <= b and not a;
    layer2_outputs(3283) <= not a or b;
    layer2_outputs(3284) <= not a or b;
    layer2_outputs(3285) <= a or b;
    layer2_outputs(3286) <= not b;
    layer2_outputs(3287) <= not b;
    layer2_outputs(3288) <= a;
    layer2_outputs(3289) <= a or b;
    layer2_outputs(3290) <= b;
    layer2_outputs(3291) <= a and not b;
    layer2_outputs(3292) <= '1';
    layer2_outputs(3293) <= not a or b;
    layer2_outputs(3294) <= not b;
    layer2_outputs(3295) <= a or b;
    layer2_outputs(3296) <= '1';
    layer2_outputs(3297) <= not (a or b);
    layer2_outputs(3298) <= b and not a;
    layer2_outputs(3299) <= b and not a;
    layer2_outputs(3300) <= '1';
    layer2_outputs(3301) <= '0';
    layer2_outputs(3302) <= not (a or b);
    layer2_outputs(3303) <= a and not b;
    layer2_outputs(3304) <= a or b;
    layer2_outputs(3305) <= b and not a;
    layer2_outputs(3306) <= not a or b;
    layer2_outputs(3307) <= a xor b;
    layer2_outputs(3308) <= a xor b;
    layer2_outputs(3309) <= not (a and b);
    layer2_outputs(3310) <= a and not b;
    layer2_outputs(3311) <= not b;
    layer2_outputs(3312) <= a;
    layer2_outputs(3313) <= a or b;
    layer2_outputs(3314) <= not a or b;
    layer2_outputs(3315) <= not (a or b);
    layer2_outputs(3316) <= a and not b;
    layer2_outputs(3317) <= not (a xor b);
    layer2_outputs(3318) <= '0';
    layer2_outputs(3319) <= a and not b;
    layer2_outputs(3320) <= not (a and b);
    layer2_outputs(3321) <= not (a or b);
    layer2_outputs(3322) <= b and not a;
    layer2_outputs(3323) <= '0';
    layer2_outputs(3324) <= a and b;
    layer2_outputs(3325) <= a;
    layer2_outputs(3326) <= b;
    layer2_outputs(3327) <= not b or a;
    layer2_outputs(3328) <= '1';
    layer2_outputs(3329) <= '1';
    layer2_outputs(3330) <= not b;
    layer2_outputs(3331) <= a or b;
    layer2_outputs(3332) <= '0';
    layer2_outputs(3333) <= a and b;
    layer2_outputs(3334) <= '1';
    layer2_outputs(3335) <= '1';
    layer2_outputs(3336) <= a and b;
    layer2_outputs(3337) <= a and b;
    layer2_outputs(3338) <= '0';
    layer2_outputs(3339) <= a and b;
    layer2_outputs(3340) <= not (a or b);
    layer2_outputs(3341) <= a or b;
    layer2_outputs(3342) <= b;
    layer2_outputs(3343) <= a or b;
    layer2_outputs(3344) <= a and not b;
    layer2_outputs(3345) <= not b or a;
    layer2_outputs(3346) <= '0';
    layer2_outputs(3347) <= b;
    layer2_outputs(3348) <= a or b;
    layer2_outputs(3349) <= '0';
    layer2_outputs(3350) <= not b or a;
    layer2_outputs(3351) <= not a;
    layer2_outputs(3352) <= b and not a;
    layer2_outputs(3353) <= not b or a;
    layer2_outputs(3354) <= a and not b;
    layer2_outputs(3355) <= not (a xor b);
    layer2_outputs(3356) <= not b or a;
    layer2_outputs(3357) <= '1';
    layer2_outputs(3358) <= '1';
    layer2_outputs(3359) <= b;
    layer2_outputs(3360) <= not b;
    layer2_outputs(3361) <= not b or a;
    layer2_outputs(3362) <= a xor b;
    layer2_outputs(3363) <= '1';
    layer2_outputs(3364) <= not b or a;
    layer2_outputs(3365) <= not (a or b);
    layer2_outputs(3366) <= a or b;
    layer2_outputs(3367) <= a and b;
    layer2_outputs(3368) <= not a;
    layer2_outputs(3369) <= not (a or b);
    layer2_outputs(3370) <= not (a or b);
    layer2_outputs(3371) <= not (a and b);
    layer2_outputs(3372) <= '0';
    layer2_outputs(3373) <= not b or a;
    layer2_outputs(3374) <= b;
    layer2_outputs(3375) <= a or b;
    layer2_outputs(3376) <= '0';
    layer2_outputs(3377) <= b;
    layer2_outputs(3378) <= b;
    layer2_outputs(3379) <= '1';
    layer2_outputs(3380) <= b and not a;
    layer2_outputs(3381) <= '1';
    layer2_outputs(3382) <= '0';
    layer2_outputs(3383) <= b;
    layer2_outputs(3384) <= '1';
    layer2_outputs(3385) <= not (a and b);
    layer2_outputs(3386) <= a and not b;
    layer2_outputs(3387) <= a;
    layer2_outputs(3388) <= a or b;
    layer2_outputs(3389) <= a;
    layer2_outputs(3390) <= not a or b;
    layer2_outputs(3391) <= a and b;
    layer2_outputs(3392) <= '1';
    layer2_outputs(3393) <= b and not a;
    layer2_outputs(3394) <= not (a or b);
    layer2_outputs(3395) <= not a or b;
    layer2_outputs(3396) <= '0';
    layer2_outputs(3397) <= not (a or b);
    layer2_outputs(3398) <= '0';
    layer2_outputs(3399) <= a or b;
    layer2_outputs(3400) <= a or b;
    layer2_outputs(3401) <= a and not b;
    layer2_outputs(3402) <= not a;
    layer2_outputs(3403) <= '0';
    layer2_outputs(3404) <= not a or b;
    layer2_outputs(3405) <= '1';
    layer2_outputs(3406) <= b and not a;
    layer2_outputs(3407) <= a;
    layer2_outputs(3408) <= '1';
    layer2_outputs(3409) <= a and not b;
    layer2_outputs(3410) <= '0';
    layer2_outputs(3411) <= not b;
    layer2_outputs(3412) <= '1';
    layer2_outputs(3413) <= a and b;
    layer2_outputs(3414) <= not a or b;
    layer2_outputs(3415) <= a and b;
    layer2_outputs(3416) <= a or b;
    layer2_outputs(3417) <= '0';
    layer2_outputs(3418) <= a and b;
    layer2_outputs(3419) <= a or b;
    layer2_outputs(3420) <= not a or b;
    layer2_outputs(3421) <= b;
    layer2_outputs(3422) <= not b or a;
    layer2_outputs(3423) <= not b;
    layer2_outputs(3424) <= not a or b;
    layer2_outputs(3425) <= '0';
    layer2_outputs(3426) <= not a or b;
    layer2_outputs(3427) <= a and not b;
    layer2_outputs(3428) <= a or b;
    layer2_outputs(3429) <= not b or a;
    layer2_outputs(3430) <= a and b;
    layer2_outputs(3431) <= a;
    layer2_outputs(3432) <= not b or a;
    layer2_outputs(3433) <= not a;
    layer2_outputs(3434) <= '1';
    layer2_outputs(3435) <= b and not a;
    layer2_outputs(3436) <= not (a or b);
    layer2_outputs(3437) <= not (a xor b);
    layer2_outputs(3438) <= not a;
    layer2_outputs(3439) <= a or b;
    layer2_outputs(3440) <= not a;
    layer2_outputs(3441) <= not a;
    layer2_outputs(3442) <= '1';
    layer2_outputs(3443) <= '1';
    layer2_outputs(3444) <= not (a or b);
    layer2_outputs(3445) <= not a or b;
    layer2_outputs(3446) <= not (a xor b);
    layer2_outputs(3447) <= '1';
    layer2_outputs(3448) <= not (a and b);
    layer2_outputs(3449) <= a and b;
    layer2_outputs(3450) <= '0';
    layer2_outputs(3451) <= not a;
    layer2_outputs(3452) <= not (a or b);
    layer2_outputs(3453) <= not (a or b);
    layer2_outputs(3454) <= not a;
    layer2_outputs(3455) <= a and b;
    layer2_outputs(3456) <= b;
    layer2_outputs(3457) <= a and not b;
    layer2_outputs(3458) <= '1';
    layer2_outputs(3459) <= '0';
    layer2_outputs(3460) <= not a;
    layer2_outputs(3461) <= a xor b;
    layer2_outputs(3462) <= '1';
    layer2_outputs(3463) <= a or b;
    layer2_outputs(3464) <= not (a xor b);
    layer2_outputs(3465) <= not b;
    layer2_outputs(3466) <= not b;
    layer2_outputs(3467) <= not (a and b);
    layer2_outputs(3468) <= not b;
    layer2_outputs(3469) <= not b or a;
    layer2_outputs(3470) <= not (a and b);
    layer2_outputs(3471) <= not b;
    layer2_outputs(3472) <= a and b;
    layer2_outputs(3473) <= not b or a;
    layer2_outputs(3474) <= a and b;
    layer2_outputs(3475) <= not b;
    layer2_outputs(3476) <= not (a or b);
    layer2_outputs(3477) <= not a;
    layer2_outputs(3478) <= a;
    layer2_outputs(3479) <= b and not a;
    layer2_outputs(3480) <= not b;
    layer2_outputs(3481) <= not b;
    layer2_outputs(3482) <= not a or b;
    layer2_outputs(3483) <= a or b;
    layer2_outputs(3484) <= not b or a;
    layer2_outputs(3485) <= a;
    layer2_outputs(3486) <= not a;
    layer2_outputs(3487) <= '1';
    layer2_outputs(3488) <= a and b;
    layer2_outputs(3489) <= a;
    layer2_outputs(3490) <= '1';
    layer2_outputs(3491) <= not (a and b);
    layer2_outputs(3492) <= not (a and b);
    layer2_outputs(3493) <= b and not a;
    layer2_outputs(3494) <= not a;
    layer2_outputs(3495) <= a and b;
    layer2_outputs(3496) <= b and not a;
    layer2_outputs(3497) <= not b or a;
    layer2_outputs(3498) <= a xor b;
    layer2_outputs(3499) <= a or b;
    layer2_outputs(3500) <= '1';
    layer2_outputs(3501) <= a;
    layer2_outputs(3502) <= a;
    layer2_outputs(3503) <= a and b;
    layer2_outputs(3504) <= b and not a;
    layer2_outputs(3505) <= a and b;
    layer2_outputs(3506) <= b;
    layer2_outputs(3507) <= not (a and b);
    layer2_outputs(3508) <= a and not b;
    layer2_outputs(3509) <= not (a and b);
    layer2_outputs(3510) <= a;
    layer2_outputs(3511) <= not b;
    layer2_outputs(3512) <= not (a and b);
    layer2_outputs(3513) <= a xor b;
    layer2_outputs(3514) <= not b or a;
    layer2_outputs(3515) <= b and not a;
    layer2_outputs(3516) <= a or b;
    layer2_outputs(3517) <= not a;
    layer2_outputs(3518) <= a;
    layer2_outputs(3519) <= not (a or b);
    layer2_outputs(3520) <= '1';
    layer2_outputs(3521) <= not b or a;
    layer2_outputs(3522) <= '1';
    layer2_outputs(3523) <= a and b;
    layer2_outputs(3524) <= a;
    layer2_outputs(3525) <= a and b;
    layer2_outputs(3526) <= a;
    layer2_outputs(3527) <= b and not a;
    layer2_outputs(3528) <= not a or b;
    layer2_outputs(3529) <= a and not b;
    layer2_outputs(3530) <= not a or b;
    layer2_outputs(3531) <= a and not b;
    layer2_outputs(3532) <= '1';
    layer2_outputs(3533) <= a and not b;
    layer2_outputs(3534) <= not (a and b);
    layer2_outputs(3535) <= not b;
    layer2_outputs(3536) <= not a or b;
    layer2_outputs(3537) <= a or b;
    layer2_outputs(3538) <= b;
    layer2_outputs(3539) <= b;
    layer2_outputs(3540) <= not b;
    layer2_outputs(3541) <= not b;
    layer2_outputs(3542) <= not (a or b);
    layer2_outputs(3543) <= b;
    layer2_outputs(3544) <= b and not a;
    layer2_outputs(3545) <= b;
    layer2_outputs(3546) <= not b or a;
    layer2_outputs(3547) <= not (a and b);
    layer2_outputs(3548) <= not a;
    layer2_outputs(3549) <= '1';
    layer2_outputs(3550) <= not (a or b);
    layer2_outputs(3551) <= '0';
    layer2_outputs(3552) <= a or b;
    layer2_outputs(3553) <= not (a or b);
    layer2_outputs(3554) <= not a or b;
    layer2_outputs(3555) <= '0';
    layer2_outputs(3556) <= not (a and b);
    layer2_outputs(3557) <= a;
    layer2_outputs(3558) <= b;
    layer2_outputs(3559) <= a;
    layer2_outputs(3560) <= a and not b;
    layer2_outputs(3561) <= a and not b;
    layer2_outputs(3562) <= not (a or b);
    layer2_outputs(3563) <= a;
    layer2_outputs(3564) <= not (a xor b);
    layer2_outputs(3565) <= a;
    layer2_outputs(3566) <= not b or a;
    layer2_outputs(3567) <= not (a xor b);
    layer2_outputs(3568) <= a and not b;
    layer2_outputs(3569) <= a or b;
    layer2_outputs(3570) <= '0';
    layer2_outputs(3571) <= '0';
    layer2_outputs(3572) <= a and b;
    layer2_outputs(3573) <= not b or a;
    layer2_outputs(3574) <= '0';
    layer2_outputs(3575) <= '0';
    layer2_outputs(3576) <= not b;
    layer2_outputs(3577) <= a and not b;
    layer2_outputs(3578) <= a and not b;
    layer2_outputs(3579) <= a or b;
    layer2_outputs(3580) <= a or b;
    layer2_outputs(3581) <= b;
    layer2_outputs(3582) <= not a;
    layer2_outputs(3583) <= not a;
    layer2_outputs(3584) <= '1';
    layer2_outputs(3585) <= not b;
    layer2_outputs(3586) <= not a;
    layer2_outputs(3587) <= not a or b;
    layer2_outputs(3588) <= not a or b;
    layer2_outputs(3589) <= a and not b;
    layer2_outputs(3590) <= not (a or b);
    layer2_outputs(3591) <= not b or a;
    layer2_outputs(3592) <= b;
    layer2_outputs(3593) <= a and b;
    layer2_outputs(3594) <= not (a or b);
    layer2_outputs(3595) <= not b or a;
    layer2_outputs(3596) <= not b or a;
    layer2_outputs(3597) <= a and not b;
    layer2_outputs(3598) <= not b or a;
    layer2_outputs(3599) <= '1';
    layer2_outputs(3600) <= a xor b;
    layer2_outputs(3601) <= '1';
    layer2_outputs(3602) <= not b or a;
    layer2_outputs(3603) <= not b;
    layer2_outputs(3604) <= not a;
    layer2_outputs(3605) <= not (a and b);
    layer2_outputs(3606) <= '1';
    layer2_outputs(3607) <= not (a and b);
    layer2_outputs(3608) <= b and not a;
    layer2_outputs(3609) <= b;
    layer2_outputs(3610) <= a;
    layer2_outputs(3611) <= b;
    layer2_outputs(3612) <= not (a and b);
    layer2_outputs(3613) <= '0';
    layer2_outputs(3614) <= not b or a;
    layer2_outputs(3615) <= '1';
    layer2_outputs(3616) <= b and not a;
    layer2_outputs(3617) <= b;
    layer2_outputs(3618) <= not (a and b);
    layer2_outputs(3619) <= not b or a;
    layer2_outputs(3620) <= a and not b;
    layer2_outputs(3621) <= b;
    layer2_outputs(3622) <= b and not a;
    layer2_outputs(3623) <= b;
    layer2_outputs(3624) <= b and not a;
    layer2_outputs(3625) <= not (a and b);
    layer2_outputs(3626) <= not (a or b);
    layer2_outputs(3627) <= not (a xor b);
    layer2_outputs(3628) <= a and b;
    layer2_outputs(3629) <= not b or a;
    layer2_outputs(3630) <= a and not b;
    layer2_outputs(3631) <= not (a and b);
    layer2_outputs(3632) <= not (a or b);
    layer2_outputs(3633) <= b and not a;
    layer2_outputs(3634) <= not a;
    layer2_outputs(3635) <= a and not b;
    layer2_outputs(3636) <= b;
    layer2_outputs(3637) <= not (a or b);
    layer2_outputs(3638) <= not (a xor b);
    layer2_outputs(3639) <= not b or a;
    layer2_outputs(3640) <= a and not b;
    layer2_outputs(3641) <= b and not a;
    layer2_outputs(3642) <= a or b;
    layer2_outputs(3643) <= b and not a;
    layer2_outputs(3644) <= a and b;
    layer2_outputs(3645) <= '1';
    layer2_outputs(3646) <= not a or b;
    layer2_outputs(3647) <= a xor b;
    layer2_outputs(3648) <= '0';
    layer2_outputs(3649) <= a;
    layer2_outputs(3650) <= a and not b;
    layer2_outputs(3651) <= a and b;
    layer2_outputs(3652) <= a and not b;
    layer2_outputs(3653) <= '0';
    layer2_outputs(3654) <= a and b;
    layer2_outputs(3655) <= b;
    layer2_outputs(3656) <= not (a and b);
    layer2_outputs(3657) <= not (a or b);
    layer2_outputs(3658) <= not a;
    layer2_outputs(3659) <= not a or b;
    layer2_outputs(3660) <= not b;
    layer2_outputs(3661) <= a;
    layer2_outputs(3662) <= not b;
    layer2_outputs(3663) <= not b;
    layer2_outputs(3664) <= a or b;
    layer2_outputs(3665) <= '1';
    layer2_outputs(3666) <= b;
    layer2_outputs(3667) <= b and not a;
    layer2_outputs(3668) <= a xor b;
    layer2_outputs(3669) <= a or b;
    layer2_outputs(3670) <= not b or a;
    layer2_outputs(3671) <= a and b;
    layer2_outputs(3672) <= a or b;
    layer2_outputs(3673) <= not b or a;
    layer2_outputs(3674) <= '0';
    layer2_outputs(3675) <= not (a or b);
    layer2_outputs(3676) <= not a or b;
    layer2_outputs(3677) <= not (a or b);
    layer2_outputs(3678) <= a and not b;
    layer2_outputs(3679) <= a and not b;
    layer2_outputs(3680) <= '0';
    layer2_outputs(3681) <= not b;
    layer2_outputs(3682) <= not a;
    layer2_outputs(3683) <= a and b;
    layer2_outputs(3684) <= not b or a;
    layer2_outputs(3685) <= not b or a;
    layer2_outputs(3686) <= a;
    layer2_outputs(3687) <= not b or a;
    layer2_outputs(3688) <= not a or b;
    layer2_outputs(3689) <= b and not a;
    layer2_outputs(3690) <= a or b;
    layer2_outputs(3691) <= a or b;
    layer2_outputs(3692) <= a and b;
    layer2_outputs(3693) <= not a or b;
    layer2_outputs(3694) <= b;
    layer2_outputs(3695) <= '0';
    layer2_outputs(3696) <= a;
    layer2_outputs(3697) <= a and not b;
    layer2_outputs(3698) <= a and b;
    layer2_outputs(3699) <= a;
    layer2_outputs(3700) <= a and b;
    layer2_outputs(3701) <= a;
    layer2_outputs(3702) <= not b;
    layer2_outputs(3703) <= '1';
    layer2_outputs(3704) <= a and b;
    layer2_outputs(3705) <= not b or a;
    layer2_outputs(3706) <= not b;
    layer2_outputs(3707) <= not a;
    layer2_outputs(3708) <= not a;
    layer2_outputs(3709) <= not (a or b);
    layer2_outputs(3710) <= '1';
    layer2_outputs(3711) <= not a or b;
    layer2_outputs(3712) <= not b;
    layer2_outputs(3713) <= not a or b;
    layer2_outputs(3714) <= '0';
    layer2_outputs(3715) <= not (a or b);
    layer2_outputs(3716) <= not a;
    layer2_outputs(3717) <= a and not b;
    layer2_outputs(3718) <= not (a and b);
    layer2_outputs(3719) <= not (a and b);
    layer2_outputs(3720) <= not b or a;
    layer2_outputs(3721) <= a;
    layer2_outputs(3722) <= not (a or b);
    layer2_outputs(3723) <= not b;
    layer2_outputs(3724) <= b;
    layer2_outputs(3725) <= '1';
    layer2_outputs(3726) <= '0';
    layer2_outputs(3727) <= a or b;
    layer2_outputs(3728) <= not (a xor b);
    layer2_outputs(3729) <= not b;
    layer2_outputs(3730) <= a or b;
    layer2_outputs(3731) <= a and not b;
    layer2_outputs(3732) <= not (a and b);
    layer2_outputs(3733) <= a and not b;
    layer2_outputs(3734) <= '0';
    layer2_outputs(3735) <= not (a and b);
    layer2_outputs(3736) <= not (a or b);
    layer2_outputs(3737) <= not b or a;
    layer2_outputs(3738) <= not b or a;
    layer2_outputs(3739) <= not (a and b);
    layer2_outputs(3740) <= not b or a;
    layer2_outputs(3741) <= a and b;
    layer2_outputs(3742) <= a;
    layer2_outputs(3743) <= not a or b;
    layer2_outputs(3744) <= b;
    layer2_outputs(3745) <= not (a and b);
    layer2_outputs(3746) <= a and b;
    layer2_outputs(3747) <= a xor b;
    layer2_outputs(3748) <= '1';
    layer2_outputs(3749) <= a or b;
    layer2_outputs(3750) <= '1';
    layer2_outputs(3751) <= not b or a;
    layer2_outputs(3752) <= not (a or b);
    layer2_outputs(3753) <= a;
    layer2_outputs(3754) <= not b;
    layer2_outputs(3755) <= not (a or b);
    layer2_outputs(3756) <= '0';
    layer2_outputs(3757) <= a;
    layer2_outputs(3758) <= not a or b;
    layer2_outputs(3759) <= not (a and b);
    layer2_outputs(3760) <= '0';
    layer2_outputs(3761) <= a;
    layer2_outputs(3762) <= b and not a;
    layer2_outputs(3763) <= not (a or b);
    layer2_outputs(3764) <= not a or b;
    layer2_outputs(3765) <= a or b;
    layer2_outputs(3766) <= '0';
    layer2_outputs(3767) <= a and b;
    layer2_outputs(3768) <= a;
    layer2_outputs(3769) <= a and not b;
    layer2_outputs(3770) <= not b or a;
    layer2_outputs(3771) <= b and not a;
    layer2_outputs(3772) <= a;
    layer2_outputs(3773) <= '1';
    layer2_outputs(3774) <= a xor b;
    layer2_outputs(3775) <= '1';
    layer2_outputs(3776) <= a and b;
    layer2_outputs(3777) <= a;
    layer2_outputs(3778) <= '1';
    layer2_outputs(3779) <= not (a or b);
    layer2_outputs(3780) <= '1';
    layer2_outputs(3781) <= a xor b;
    layer2_outputs(3782) <= not (a and b);
    layer2_outputs(3783) <= b and not a;
    layer2_outputs(3784) <= b;
    layer2_outputs(3785) <= b and not a;
    layer2_outputs(3786) <= not (a or b);
    layer2_outputs(3787) <= a;
    layer2_outputs(3788) <= not b;
    layer2_outputs(3789) <= a and b;
    layer2_outputs(3790) <= b and not a;
    layer2_outputs(3791) <= b and not a;
    layer2_outputs(3792) <= a;
    layer2_outputs(3793) <= b;
    layer2_outputs(3794) <= '1';
    layer2_outputs(3795) <= not b or a;
    layer2_outputs(3796) <= not (a or b);
    layer2_outputs(3797) <= b and not a;
    layer2_outputs(3798) <= not b or a;
    layer2_outputs(3799) <= a xor b;
    layer2_outputs(3800) <= b and not a;
    layer2_outputs(3801) <= b;
    layer2_outputs(3802) <= not b or a;
    layer2_outputs(3803) <= '0';
    layer2_outputs(3804) <= not (a or b);
    layer2_outputs(3805) <= not (a or b);
    layer2_outputs(3806) <= a;
    layer2_outputs(3807) <= a or b;
    layer2_outputs(3808) <= b and not a;
    layer2_outputs(3809) <= not a or b;
    layer2_outputs(3810) <= not b or a;
    layer2_outputs(3811) <= a and b;
    layer2_outputs(3812) <= not (a and b);
    layer2_outputs(3813) <= not (a and b);
    layer2_outputs(3814) <= b;
    layer2_outputs(3815) <= not a or b;
    layer2_outputs(3816) <= '0';
    layer2_outputs(3817) <= not a;
    layer2_outputs(3818) <= '0';
    layer2_outputs(3819) <= not a;
    layer2_outputs(3820) <= not a or b;
    layer2_outputs(3821) <= not a or b;
    layer2_outputs(3822) <= not b;
    layer2_outputs(3823) <= a and not b;
    layer2_outputs(3824) <= b and not a;
    layer2_outputs(3825) <= not a or b;
    layer2_outputs(3826) <= a and b;
    layer2_outputs(3827) <= a and not b;
    layer2_outputs(3828) <= not a;
    layer2_outputs(3829) <= '1';
    layer2_outputs(3830) <= a and not b;
    layer2_outputs(3831) <= a;
    layer2_outputs(3832) <= b and not a;
    layer2_outputs(3833) <= b and not a;
    layer2_outputs(3834) <= not b or a;
    layer2_outputs(3835) <= a and b;
    layer2_outputs(3836) <= not (a and b);
    layer2_outputs(3837) <= a and not b;
    layer2_outputs(3838) <= '1';
    layer2_outputs(3839) <= a;
    layer2_outputs(3840) <= not a;
    layer2_outputs(3841) <= a and b;
    layer2_outputs(3842) <= not (a and b);
    layer2_outputs(3843) <= not (a xor b);
    layer2_outputs(3844) <= b;
    layer2_outputs(3845) <= not a or b;
    layer2_outputs(3846) <= b and not a;
    layer2_outputs(3847) <= not (a or b);
    layer2_outputs(3848) <= not (a or b);
    layer2_outputs(3849) <= '0';
    layer2_outputs(3850) <= '1';
    layer2_outputs(3851) <= b and not a;
    layer2_outputs(3852) <= a;
    layer2_outputs(3853) <= not (a or b);
    layer2_outputs(3854) <= b;
    layer2_outputs(3855) <= b;
    layer2_outputs(3856) <= a and not b;
    layer2_outputs(3857) <= not a;
    layer2_outputs(3858) <= not (a and b);
    layer2_outputs(3859) <= not b or a;
    layer2_outputs(3860) <= not b or a;
    layer2_outputs(3861) <= not b or a;
    layer2_outputs(3862) <= a or b;
    layer2_outputs(3863) <= not (a or b);
    layer2_outputs(3864) <= not a or b;
    layer2_outputs(3865) <= '1';
    layer2_outputs(3866) <= not a;
    layer2_outputs(3867) <= not b;
    layer2_outputs(3868) <= not a;
    layer2_outputs(3869) <= not (a and b);
    layer2_outputs(3870) <= a xor b;
    layer2_outputs(3871) <= '1';
    layer2_outputs(3872) <= '0';
    layer2_outputs(3873) <= '0';
    layer2_outputs(3874) <= not b;
    layer2_outputs(3875) <= a and not b;
    layer2_outputs(3876) <= not b;
    layer2_outputs(3877) <= '0';
    layer2_outputs(3878) <= a;
    layer2_outputs(3879) <= '0';
    layer2_outputs(3880) <= not b or a;
    layer2_outputs(3881) <= not (a or b);
    layer2_outputs(3882) <= not a;
    layer2_outputs(3883) <= a and not b;
    layer2_outputs(3884) <= a;
    layer2_outputs(3885) <= not (a xor b);
    layer2_outputs(3886) <= '1';
    layer2_outputs(3887) <= not b;
    layer2_outputs(3888) <= a or b;
    layer2_outputs(3889) <= a xor b;
    layer2_outputs(3890) <= not a;
    layer2_outputs(3891) <= a and not b;
    layer2_outputs(3892) <= a xor b;
    layer2_outputs(3893) <= '0';
    layer2_outputs(3894) <= a xor b;
    layer2_outputs(3895) <= '0';
    layer2_outputs(3896) <= b;
    layer2_outputs(3897) <= not (a and b);
    layer2_outputs(3898) <= not (a and b);
    layer2_outputs(3899) <= '1';
    layer2_outputs(3900) <= a or b;
    layer2_outputs(3901) <= a;
    layer2_outputs(3902) <= a and not b;
    layer2_outputs(3903) <= a and b;
    layer2_outputs(3904) <= a and not b;
    layer2_outputs(3905) <= a and not b;
    layer2_outputs(3906) <= a and b;
    layer2_outputs(3907) <= '0';
    layer2_outputs(3908) <= b;
    layer2_outputs(3909) <= a and not b;
    layer2_outputs(3910) <= a;
    layer2_outputs(3911) <= a or b;
    layer2_outputs(3912) <= not b or a;
    layer2_outputs(3913) <= a or b;
    layer2_outputs(3914) <= not b or a;
    layer2_outputs(3915) <= not (a and b);
    layer2_outputs(3916) <= a;
    layer2_outputs(3917) <= not a;
    layer2_outputs(3918) <= not a;
    layer2_outputs(3919) <= not b;
    layer2_outputs(3920) <= a or b;
    layer2_outputs(3921) <= not a;
    layer2_outputs(3922) <= not a or b;
    layer2_outputs(3923) <= a or b;
    layer2_outputs(3924) <= not a or b;
    layer2_outputs(3925) <= b;
    layer2_outputs(3926) <= a and b;
    layer2_outputs(3927) <= a or b;
    layer2_outputs(3928) <= '1';
    layer2_outputs(3929) <= not a or b;
    layer2_outputs(3930) <= '0';
    layer2_outputs(3931) <= a or b;
    layer2_outputs(3932) <= a and not b;
    layer2_outputs(3933) <= '0';
    layer2_outputs(3934) <= not (a and b);
    layer2_outputs(3935) <= not (a or b);
    layer2_outputs(3936) <= '1';
    layer2_outputs(3937) <= not (a or b);
    layer2_outputs(3938) <= not b;
    layer2_outputs(3939) <= a and b;
    layer2_outputs(3940) <= a and not b;
    layer2_outputs(3941) <= a;
    layer2_outputs(3942) <= not a;
    layer2_outputs(3943) <= not a;
    layer2_outputs(3944) <= a;
    layer2_outputs(3945) <= a;
    layer2_outputs(3946) <= not a;
    layer2_outputs(3947) <= b;
    layer2_outputs(3948) <= not a or b;
    layer2_outputs(3949) <= not b;
    layer2_outputs(3950) <= '1';
    layer2_outputs(3951) <= a and not b;
    layer2_outputs(3952) <= '0';
    layer2_outputs(3953) <= b;
    layer2_outputs(3954) <= a;
    layer2_outputs(3955) <= not (a and b);
    layer2_outputs(3956) <= a xor b;
    layer2_outputs(3957) <= not b;
    layer2_outputs(3958) <= not a;
    layer2_outputs(3959) <= a and not b;
    layer2_outputs(3960) <= b and not a;
    layer2_outputs(3961) <= '1';
    layer2_outputs(3962) <= b and not a;
    layer2_outputs(3963) <= '0';
    layer2_outputs(3964) <= a and b;
    layer2_outputs(3965) <= not b;
    layer2_outputs(3966) <= '1';
    layer2_outputs(3967) <= a and not b;
    layer2_outputs(3968) <= a and b;
    layer2_outputs(3969) <= a or b;
    layer2_outputs(3970) <= '1';
    layer2_outputs(3971) <= a and b;
    layer2_outputs(3972) <= b and not a;
    layer2_outputs(3973) <= not b;
    layer2_outputs(3974) <= not (a or b);
    layer2_outputs(3975) <= not (a or b);
    layer2_outputs(3976) <= not (a and b);
    layer2_outputs(3977) <= a or b;
    layer2_outputs(3978) <= not (a and b);
    layer2_outputs(3979) <= b;
    layer2_outputs(3980) <= a and b;
    layer2_outputs(3981) <= not (a and b);
    layer2_outputs(3982) <= '1';
    layer2_outputs(3983) <= not (a or b);
    layer2_outputs(3984) <= '0';
    layer2_outputs(3985) <= not a or b;
    layer2_outputs(3986) <= a and not b;
    layer2_outputs(3987) <= a and not b;
    layer2_outputs(3988) <= not (a and b);
    layer2_outputs(3989) <= not a or b;
    layer2_outputs(3990) <= a and b;
    layer2_outputs(3991) <= '1';
    layer2_outputs(3992) <= '1';
    layer2_outputs(3993) <= '1';
    layer2_outputs(3994) <= '1';
    layer2_outputs(3995) <= a or b;
    layer2_outputs(3996) <= b and not a;
    layer2_outputs(3997) <= '0';
    layer2_outputs(3998) <= a or b;
    layer2_outputs(3999) <= '0';
    layer2_outputs(4000) <= not (a or b);
    layer2_outputs(4001) <= not (a or b);
    layer2_outputs(4002) <= not a;
    layer2_outputs(4003) <= not b or a;
    layer2_outputs(4004) <= not (a and b);
    layer2_outputs(4005) <= a or b;
    layer2_outputs(4006) <= not b;
    layer2_outputs(4007) <= not (a or b);
    layer2_outputs(4008) <= b and not a;
    layer2_outputs(4009) <= not (a or b);
    layer2_outputs(4010) <= '0';
    layer2_outputs(4011) <= not a;
    layer2_outputs(4012) <= not (a or b);
    layer2_outputs(4013) <= '0';
    layer2_outputs(4014) <= '0';
    layer2_outputs(4015) <= '1';
    layer2_outputs(4016) <= a xor b;
    layer2_outputs(4017) <= a xor b;
    layer2_outputs(4018) <= not (a and b);
    layer2_outputs(4019) <= not a or b;
    layer2_outputs(4020) <= '0';
    layer2_outputs(4021) <= not a or b;
    layer2_outputs(4022) <= not b or a;
    layer2_outputs(4023) <= a or b;
    layer2_outputs(4024) <= b;
    layer2_outputs(4025) <= not a or b;
    layer2_outputs(4026) <= '1';
    layer2_outputs(4027) <= not a;
    layer2_outputs(4028) <= '1';
    layer2_outputs(4029) <= not (a or b);
    layer2_outputs(4030) <= a and not b;
    layer2_outputs(4031) <= a and not b;
    layer2_outputs(4032) <= '1';
    layer2_outputs(4033) <= not a;
    layer2_outputs(4034) <= not b or a;
    layer2_outputs(4035) <= '1';
    layer2_outputs(4036) <= not (a xor b);
    layer2_outputs(4037) <= a and b;
    layer2_outputs(4038) <= b and not a;
    layer2_outputs(4039) <= '0';
    layer2_outputs(4040) <= '0';
    layer2_outputs(4041) <= a or b;
    layer2_outputs(4042) <= not a or b;
    layer2_outputs(4043) <= not b;
    layer2_outputs(4044) <= not a or b;
    layer2_outputs(4045) <= not (a or b);
    layer2_outputs(4046) <= not b or a;
    layer2_outputs(4047) <= not a;
    layer2_outputs(4048) <= '0';
    layer2_outputs(4049) <= not b or a;
    layer2_outputs(4050) <= a or b;
    layer2_outputs(4051) <= b;
    layer2_outputs(4052) <= not b or a;
    layer2_outputs(4053) <= a;
    layer2_outputs(4054) <= a or b;
    layer2_outputs(4055) <= not (a or b);
    layer2_outputs(4056) <= not a;
    layer2_outputs(4057) <= b;
    layer2_outputs(4058) <= not b or a;
    layer2_outputs(4059) <= '0';
    layer2_outputs(4060) <= not (a and b);
    layer2_outputs(4061) <= not b;
    layer2_outputs(4062) <= a xor b;
    layer2_outputs(4063) <= not a;
    layer2_outputs(4064) <= not b;
    layer2_outputs(4065) <= b;
    layer2_outputs(4066) <= '0';
    layer2_outputs(4067) <= a or b;
    layer2_outputs(4068) <= not (a xor b);
    layer2_outputs(4069) <= not b or a;
    layer2_outputs(4070) <= not (a and b);
    layer2_outputs(4071) <= '1';
    layer2_outputs(4072) <= not (a and b);
    layer2_outputs(4073) <= a and b;
    layer2_outputs(4074) <= not a;
    layer2_outputs(4075) <= '0';
    layer2_outputs(4076) <= a or b;
    layer2_outputs(4077) <= a and b;
    layer2_outputs(4078) <= b and not a;
    layer2_outputs(4079) <= b;
    layer2_outputs(4080) <= '1';
    layer2_outputs(4081) <= not (a and b);
    layer2_outputs(4082) <= not b or a;
    layer2_outputs(4083) <= '0';
    layer2_outputs(4084) <= b and not a;
    layer2_outputs(4085) <= a or b;
    layer2_outputs(4086) <= '0';
    layer2_outputs(4087) <= not a or b;
    layer2_outputs(4088) <= not a;
    layer2_outputs(4089) <= not b;
    layer2_outputs(4090) <= not a;
    layer2_outputs(4091) <= b;
    layer2_outputs(4092) <= not a or b;
    layer2_outputs(4093) <= not (a or b);
    layer2_outputs(4094) <= b and not a;
    layer2_outputs(4095) <= a or b;
    layer2_outputs(4096) <= a or b;
    layer2_outputs(4097) <= not (a and b);
    layer2_outputs(4098) <= not a;
    layer2_outputs(4099) <= a and b;
    layer2_outputs(4100) <= '0';
    layer2_outputs(4101) <= a and not b;
    layer2_outputs(4102) <= not b;
    layer2_outputs(4103) <= not (a and b);
    layer2_outputs(4104) <= not b or a;
    layer2_outputs(4105) <= not b;
    layer2_outputs(4106) <= '1';
    layer2_outputs(4107) <= a xor b;
    layer2_outputs(4108) <= '0';
    layer2_outputs(4109) <= b and not a;
    layer2_outputs(4110) <= not b;
    layer2_outputs(4111) <= a;
    layer2_outputs(4112) <= b;
    layer2_outputs(4113) <= a and not b;
    layer2_outputs(4114) <= a and b;
    layer2_outputs(4115) <= b;
    layer2_outputs(4116) <= '1';
    layer2_outputs(4117) <= '0';
    layer2_outputs(4118) <= a or b;
    layer2_outputs(4119) <= a and not b;
    layer2_outputs(4120) <= not b;
    layer2_outputs(4121) <= not b;
    layer2_outputs(4122) <= a or b;
    layer2_outputs(4123) <= not (a or b);
    layer2_outputs(4124) <= a and b;
    layer2_outputs(4125) <= '1';
    layer2_outputs(4126) <= '1';
    layer2_outputs(4127) <= a and b;
    layer2_outputs(4128) <= a and not b;
    layer2_outputs(4129) <= '0';
    layer2_outputs(4130) <= not b or a;
    layer2_outputs(4131) <= a or b;
    layer2_outputs(4132) <= '1';
    layer2_outputs(4133) <= not (a and b);
    layer2_outputs(4134) <= '0';
    layer2_outputs(4135) <= a;
    layer2_outputs(4136) <= b;
    layer2_outputs(4137) <= '1';
    layer2_outputs(4138) <= '1';
    layer2_outputs(4139) <= '0';
    layer2_outputs(4140) <= a and not b;
    layer2_outputs(4141) <= b;
    layer2_outputs(4142) <= not a or b;
    layer2_outputs(4143) <= '1';
    layer2_outputs(4144) <= not (a xor b);
    layer2_outputs(4145) <= not (a and b);
    layer2_outputs(4146) <= b;
    layer2_outputs(4147) <= not a or b;
    layer2_outputs(4148) <= not b or a;
    layer2_outputs(4149) <= a and not b;
    layer2_outputs(4150) <= b;
    layer2_outputs(4151) <= not (a or b);
    layer2_outputs(4152) <= not (a and b);
    layer2_outputs(4153) <= not (a and b);
    layer2_outputs(4154) <= a or b;
    layer2_outputs(4155) <= b;
    layer2_outputs(4156) <= '0';
    layer2_outputs(4157) <= not a;
    layer2_outputs(4158) <= a xor b;
    layer2_outputs(4159) <= b and not a;
    layer2_outputs(4160) <= a and b;
    layer2_outputs(4161) <= a and b;
    layer2_outputs(4162) <= not a or b;
    layer2_outputs(4163) <= not b;
    layer2_outputs(4164) <= not (a and b);
    layer2_outputs(4165) <= a and not b;
    layer2_outputs(4166) <= a xor b;
    layer2_outputs(4167) <= a xor b;
    layer2_outputs(4168) <= not (a and b);
    layer2_outputs(4169) <= not b or a;
    layer2_outputs(4170) <= '1';
    layer2_outputs(4171) <= '0';
    layer2_outputs(4172) <= a;
    layer2_outputs(4173) <= not a;
    layer2_outputs(4174) <= '0';
    layer2_outputs(4175) <= b and not a;
    layer2_outputs(4176) <= b;
    layer2_outputs(4177) <= a or b;
    layer2_outputs(4178) <= a and b;
    layer2_outputs(4179) <= a and b;
    layer2_outputs(4180) <= not b or a;
    layer2_outputs(4181) <= b;
    layer2_outputs(4182) <= '1';
    layer2_outputs(4183) <= not a;
    layer2_outputs(4184) <= not a or b;
    layer2_outputs(4185) <= not a;
    layer2_outputs(4186) <= b and not a;
    layer2_outputs(4187) <= not (a or b);
    layer2_outputs(4188) <= b;
    layer2_outputs(4189) <= not b or a;
    layer2_outputs(4190) <= '0';
    layer2_outputs(4191) <= b;
    layer2_outputs(4192) <= not (a or b);
    layer2_outputs(4193) <= a and b;
    layer2_outputs(4194) <= '0';
    layer2_outputs(4195) <= a or b;
    layer2_outputs(4196) <= a or b;
    layer2_outputs(4197) <= '0';
    layer2_outputs(4198) <= not b;
    layer2_outputs(4199) <= not a;
    layer2_outputs(4200) <= a;
    layer2_outputs(4201) <= '0';
    layer2_outputs(4202) <= not b or a;
    layer2_outputs(4203) <= '1';
    layer2_outputs(4204) <= b;
    layer2_outputs(4205) <= a and not b;
    layer2_outputs(4206) <= a;
    layer2_outputs(4207) <= a and b;
    layer2_outputs(4208) <= a xor b;
    layer2_outputs(4209) <= a and not b;
    layer2_outputs(4210) <= not a or b;
    layer2_outputs(4211) <= '0';
    layer2_outputs(4212) <= a and b;
    layer2_outputs(4213) <= not (a or b);
    layer2_outputs(4214) <= a and b;
    layer2_outputs(4215) <= a;
    layer2_outputs(4216) <= b and not a;
    layer2_outputs(4217) <= a and b;
    layer2_outputs(4218) <= not (a and b);
    layer2_outputs(4219) <= a or b;
    layer2_outputs(4220) <= not (a or b);
    layer2_outputs(4221) <= not b or a;
    layer2_outputs(4222) <= a and not b;
    layer2_outputs(4223) <= a and not b;
    layer2_outputs(4224) <= a and not b;
    layer2_outputs(4225) <= not b;
    layer2_outputs(4226) <= '0';
    layer2_outputs(4227) <= '0';
    layer2_outputs(4228) <= not (a or b);
    layer2_outputs(4229) <= a or b;
    layer2_outputs(4230) <= not a or b;
    layer2_outputs(4231) <= not b or a;
    layer2_outputs(4232) <= '1';
    layer2_outputs(4233) <= b and not a;
    layer2_outputs(4234) <= '0';
    layer2_outputs(4235) <= a;
    layer2_outputs(4236) <= not (a or b);
    layer2_outputs(4237) <= not b or a;
    layer2_outputs(4238) <= a;
    layer2_outputs(4239) <= b and not a;
    layer2_outputs(4240) <= not a;
    layer2_outputs(4241) <= b and not a;
    layer2_outputs(4242) <= not a or b;
    layer2_outputs(4243) <= b and not a;
    layer2_outputs(4244) <= '0';
    layer2_outputs(4245) <= not (a xor b);
    layer2_outputs(4246) <= '1';
    layer2_outputs(4247) <= a and b;
    layer2_outputs(4248) <= not a;
    layer2_outputs(4249) <= not (a or b);
    layer2_outputs(4250) <= not a;
    layer2_outputs(4251) <= not b or a;
    layer2_outputs(4252) <= not (a or b);
    layer2_outputs(4253) <= not b or a;
    layer2_outputs(4254) <= '1';
    layer2_outputs(4255) <= not a or b;
    layer2_outputs(4256) <= not (a or b);
    layer2_outputs(4257) <= a xor b;
    layer2_outputs(4258) <= a and not b;
    layer2_outputs(4259) <= a;
    layer2_outputs(4260) <= not b or a;
    layer2_outputs(4261) <= a;
    layer2_outputs(4262) <= not (a and b);
    layer2_outputs(4263) <= a and not b;
    layer2_outputs(4264) <= '0';
    layer2_outputs(4265) <= not a or b;
    layer2_outputs(4266) <= '0';
    layer2_outputs(4267) <= not b;
    layer2_outputs(4268) <= a and not b;
    layer2_outputs(4269) <= a;
    layer2_outputs(4270) <= not b;
    layer2_outputs(4271) <= not (a xor b);
    layer2_outputs(4272) <= '0';
    layer2_outputs(4273) <= not a or b;
    layer2_outputs(4274) <= a and not b;
    layer2_outputs(4275) <= a xor b;
    layer2_outputs(4276) <= not a or b;
    layer2_outputs(4277) <= a or b;
    layer2_outputs(4278) <= '1';
    layer2_outputs(4279) <= not b;
    layer2_outputs(4280) <= b and not a;
    layer2_outputs(4281) <= not b;
    layer2_outputs(4282) <= not b or a;
    layer2_outputs(4283) <= not b or a;
    layer2_outputs(4284) <= a and b;
    layer2_outputs(4285) <= a;
    layer2_outputs(4286) <= not (a or b);
    layer2_outputs(4287) <= not b or a;
    layer2_outputs(4288) <= not (a or b);
    layer2_outputs(4289) <= '0';
    layer2_outputs(4290) <= not (a xor b);
    layer2_outputs(4291) <= a or b;
    layer2_outputs(4292) <= a xor b;
    layer2_outputs(4293) <= '1';
    layer2_outputs(4294) <= b and not a;
    layer2_outputs(4295) <= a and b;
    layer2_outputs(4296) <= '1';
    layer2_outputs(4297) <= not a or b;
    layer2_outputs(4298) <= a;
    layer2_outputs(4299) <= a and not b;
    layer2_outputs(4300) <= not a;
    layer2_outputs(4301) <= not (a and b);
    layer2_outputs(4302) <= a and not b;
    layer2_outputs(4303) <= b and not a;
    layer2_outputs(4304) <= '0';
    layer2_outputs(4305) <= not a or b;
    layer2_outputs(4306) <= not a;
    layer2_outputs(4307) <= not b or a;
    layer2_outputs(4308) <= '1';
    layer2_outputs(4309) <= not b or a;
    layer2_outputs(4310) <= not a;
    layer2_outputs(4311) <= not b or a;
    layer2_outputs(4312) <= '0';
    layer2_outputs(4313) <= not b or a;
    layer2_outputs(4314) <= not (a or b);
    layer2_outputs(4315) <= not b or a;
    layer2_outputs(4316) <= b and not a;
    layer2_outputs(4317) <= b;
    layer2_outputs(4318) <= not (a xor b);
    layer2_outputs(4319) <= not a;
    layer2_outputs(4320) <= '1';
    layer2_outputs(4321) <= not b or a;
    layer2_outputs(4322) <= not a or b;
    layer2_outputs(4323) <= not (a and b);
    layer2_outputs(4324) <= not (a and b);
    layer2_outputs(4325) <= not a or b;
    layer2_outputs(4326) <= not b;
    layer2_outputs(4327) <= b;
    layer2_outputs(4328) <= a and not b;
    layer2_outputs(4329) <= '0';
    layer2_outputs(4330) <= '0';
    layer2_outputs(4331) <= '1';
    layer2_outputs(4332) <= not (a xor b);
    layer2_outputs(4333) <= b;
    layer2_outputs(4334) <= '0';
    layer2_outputs(4335) <= '0';
    layer2_outputs(4336) <= a xor b;
    layer2_outputs(4337) <= b;
    layer2_outputs(4338) <= b and not a;
    layer2_outputs(4339) <= a xor b;
    layer2_outputs(4340) <= a;
    layer2_outputs(4341) <= not a or b;
    layer2_outputs(4342) <= not b or a;
    layer2_outputs(4343) <= not (a or b);
    layer2_outputs(4344) <= '1';
    layer2_outputs(4345) <= a and b;
    layer2_outputs(4346) <= a or b;
    layer2_outputs(4347) <= '0';
    layer2_outputs(4348) <= not a or b;
    layer2_outputs(4349) <= not b;
    layer2_outputs(4350) <= not b;
    layer2_outputs(4351) <= not a or b;
    layer2_outputs(4352) <= b;
    layer2_outputs(4353) <= not a or b;
    layer2_outputs(4354) <= not a;
    layer2_outputs(4355) <= a and not b;
    layer2_outputs(4356) <= not (a or b);
    layer2_outputs(4357) <= a and b;
    layer2_outputs(4358) <= not b or a;
    layer2_outputs(4359) <= not b or a;
    layer2_outputs(4360) <= a and not b;
    layer2_outputs(4361) <= not (a xor b);
    layer2_outputs(4362) <= b and not a;
    layer2_outputs(4363) <= b;
    layer2_outputs(4364) <= '0';
    layer2_outputs(4365) <= a or b;
    layer2_outputs(4366) <= not (a or b);
    layer2_outputs(4367) <= b;
    layer2_outputs(4368) <= a and not b;
    layer2_outputs(4369) <= not (a and b);
    layer2_outputs(4370) <= a or b;
    layer2_outputs(4371) <= b;
    layer2_outputs(4372) <= not b;
    layer2_outputs(4373) <= not a or b;
    layer2_outputs(4374) <= not b;
    layer2_outputs(4375) <= not a or b;
    layer2_outputs(4376) <= '0';
    layer2_outputs(4377) <= b;
    layer2_outputs(4378) <= a and b;
    layer2_outputs(4379) <= '0';
    layer2_outputs(4380) <= a and b;
    layer2_outputs(4381) <= not b;
    layer2_outputs(4382) <= '0';
    layer2_outputs(4383) <= not a or b;
    layer2_outputs(4384) <= a and b;
    layer2_outputs(4385) <= a and not b;
    layer2_outputs(4386) <= not (a and b);
    layer2_outputs(4387) <= '0';
    layer2_outputs(4388) <= not (a and b);
    layer2_outputs(4389) <= a and not b;
    layer2_outputs(4390) <= b and not a;
    layer2_outputs(4391) <= not a;
    layer2_outputs(4392) <= '0';
    layer2_outputs(4393) <= not (a or b);
    layer2_outputs(4394) <= b and not a;
    layer2_outputs(4395) <= not (a xor b);
    layer2_outputs(4396) <= a and not b;
    layer2_outputs(4397) <= not (a or b);
    layer2_outputs(4398) <= not b;
    layer2_outputs(4399) <= not b;
    layer2_outputs(4400) <= not b or a;
    layer2_outputs(4401) <= not b;
    layer2_outputs(4402) <= a;
    layer2_outputs(4403) <= a and b;
    layer2_outputs(4404) <= a;
    layer2_outputs(4405) <= b and not a;
    layer2_outputs(4406) <= a or b;
    layer2_outputs(4407) <= not b;
    layer2_outputs(4408) <= '1';
    layer2_outputs(4409) <= a and not b;
    layer2_outputs(4410) <= a and not b;
    layer2_outputs(4411) <= not b;
    layer2_outputs(4412) <= not (a or b);
    layer2_outputs(4413) <= not (a or b);
    layer2_outputs(4414) <= not (a and b);
    layer2_outputs(4415) <= a;
    layer2_outputs(4416) <= not (a and b);
    layer2_outputs(4417) <= not b;
    layer2_outputs(4418) <= b and not a;
    layer2_outputs(4419) <= not b or a;
    layer2_outputs(4420) <= a and b;
    layer2_outputs(4421) <= not (a or b);
    layer2_outputs(4422) <= a;
    layer2_outputs(4423) <= a and not b;
    layer2_outputs(4424) <= '0';
    layer2_outputs(4425) <= not b or a;
    layer2_outputs(4426) <= a and not b;
    layer2_outputs(4427) <= b and not a;
    layer2_outputs(4428) <= not b or a;
    layer2_outputs(4429) <= a or b;
    layer2_outputs(4430) <= '1';
    layer2_outputs(4431) <= '0';
    layer2_outputs(4432) <= not b;
    layer2_outputs(4433) <= b and not a;
    layer2_outputs(4434) <= not (a or b);
    layer2_outputs(4435) <= '0';
    layer2_outputs(4436) <= b;
    layer2_outputs(4437) <= a and b;
    layer2_outputs(4438) <= b and not a;
    layer2_outputs(4439) <= a and not b;
    layer2_outputs(4440) <= b;
    layer2_outputs(4441) <= b;
    layer2_outputs(4442) <= a and not b;
    layer2_outputs(4443) <= b;
    layer2_outputs(4444) <= not (a xor b);
    layer2_outputs(4445) <= b;
    layer2_outputs(4446) <= '1';
    layer2_outputs(4447) <= not (a and b);
    layer2_outputs(4448) <= b;
    layer2_outputs(4449) <= not b;
    layer2_outputs(4450) <= b and not a;
    layer2_outputs(4451) <= a or b;
    layer2_outputs(4452) <= a or b;
    layer2_outputs(4453) <= not b or a;
    layer2_outputs(4454) <= a and b;
    layer2_outputs(4455) <= '0';
    layer2_outputs(4456) <= '1';
    layer2_outputs(4457) <= not a or b;
    layer2_outputs(4458) <= not b or a;
    layer2_outputs(4459) <= a;
    layer2_outputs(4460) <= a and b;
    layer2_outputs(4461) <= a;
    layer2_outputs(4462) <= '1';
    layer2_outputs(4463) <= not (a or b);
    layer2_outputs(4464) <= not (a and b);
    layer2_outputs(4465) <= '1';
    layer2_outputs(4466) <= not a or b;
    layer2_outputs(4467) <= '0';
    layer2_outputs(4468) <= b;
    layer2_outputs(4469) <= a and b;
    layer2_outputs(4470) <= b and not a;
    layer2_outputs(4471) <= a and not b;
    layer2_outputs(4472) <= not (a xor b);
    layer2_outputs(4473) <= not (a or b);
    layer2_outputs(4474) <= a;
    layer2_outputs(4475) <= a and b;
    layer2_outputs(4476) <= not (a or b);
    layer2_outputs(4477) <= a;
    layer2_outputs(4478) <= '1';
    layer2_outputs(4479) <= b;
    layer2_outputs(4480) <= '0';
    layer2_outputs(4481) <= b;
    layer2_outputs(4482) <= b;
    layer2_outputs(4483) <= a and not b;
    layer2_outputs(4484) <= not (a xor b);
    layer2_outputs(4485) <= a or b;
    layer2_outputs(4486) <= not a or b;
    layer2_outputs(4487) <= a and not b;
    layer2_outputs(4488) <= b and not a;
    layer2_outputs(4489) <= not (a and b);
    layer2_outputs(4490) <= b;
    layer2_outputs(4491) <= '0';
    layer2_outputs(4492) <= '0';
    layer2_outputs(4493) <= not b;
    layer2_outputs(4494) <= a;
    layer2_outputs(4495) <= a and b;
    layer2_outputs(4496) <= a and not b;
    layer2_outputs(4497) <= not (a and b);
    layer2_outputs(4498) <= a and not b;
    layer2_outputs(4499) <= not (a or b);
    layer2_outputs(4500) <= a and b;
    layer2_outputs(4501) <= a or b;
    layer2_outputs(4502) <= a;
    layer2_outputs(4503) <= not (a or b);
    layer2_outputs(4504) <= not b or a;
    layer2_outputs(4505) <= not (a xor b);
    layer2_outputs(4506) <= not a or b;
    layer2_outputs(4507) <= not b or a;
    layer2_outputs(4508) <= a and b;
    layer2_outputs(4509) <= a and not b;
    layer2_outputs(4510) <= '0';
    layer2_outputs(4511) <= a and b;
    layer2_outputs(4512) <= a or b;
    layer2_outputs(4513) <= not a or b;
    layer2_outputs(4514) <= a;
    layer2_outputs(4515) <= not b;
    layer2_outputs(4516) <= not (a or b);
    layer2_outputs(4517) <= b and not a;
    layer2_outputs(4518) <= '1';
    layer2_outputs(4519) <= not (a xor b);
    layer2_outputs(4520) <= not a or b;
    layer2_outputs(4521) <= not (a xor b);
    layer2_outputs(4522) <= b and not a;
    layer2_outputs(4523) <= b and not a;
    layer2_outputs(4524) <= a and not b;
    layer2_outputs(4525) <= '0';
    layer2_outputs(4526) <= b;
    layer2_outputs(4527) <= not b or a;
    layer2_outputs(4528) <= a or b;
    layer2_outputs(4529) <= a and not b;
    layer2_outputs(4530) <= '0';
    layer2_outputs(4531) <= not a;
    layer2_outputs(4532) <= a and not b;
    layer2_outputs(4533) <= '1';
    layer2_outputs(4534) <= not (a or b);
    layer2_outputs(4535) <= a and not b;
    layer2_outputs(4536) <= a or b;
    layer2_outputs(4537) <= not (a and b);
    layer2_outputs(4538) <= not b;
    layer2_outputs(4539) <= not (a or b);
    layer2_outputs(4540) <= a or b;
    layer2_outputs(4541) <= not (a and b);
    layer2_outputs(4542) <= a and b;
    layer2_outputs(4543) <= not (a and b);
    layer2_outputs(4544) <= not (a and b);
    layer2_outputs(4545) <= b and not a;
    layer2_outputs(4546) <= not b;
    layer2_outputs(4547) <= a;
    layer2_outputs(4548) <= '1';
    layer2_outputs(4549) <= b;
    layer2_outputs(4550) <= b;
    layer2_outputs(4551) <= '1';
    layer2_outputs(4552) <= a or b;
    layer2_outputs(4553) <= not a or b;
    layer2_outputs(4554) <= a and b;
    layer2_outputs(4555) <= '1';
    layer2_outputs(4556) <= a;
    layer2_outputs(4557) <= not (a or b);
    layer2_outputs(4558) <= a;
    layer2_outputs(4559) <= '0';
    layer2_outputs(4560) <= b;
    layer2_outputs(4561) <= not (a or b);
    layer2_outputs(4562) <= '1';
    layer2_outputs(4563) <= a and not b;
    layer2_outputs(4564) <= a and not b;
    layer2_outputs(4565) <= not (a and b);
    layer2_outputs(4566) <= not b or a;
    layer2_outputs(4567) <= not a or b;
    layer2_outputs(4568) <= not (a and b);
    layer2_outputs(4569) <= not b;
    layer2_outputs(4570) <= not b or a;
    layer2_outputs(4571) <= '0';
    layer2_outputs(4572) <= '1';
    layer2_outputs(4573) <= not b or a;
    layer2_outputs(4574) <= not a or b;
    layer2_outputs(4575) <= a and not b;
    layer2_outputs(4576) <= not b or a;
    layer2_outputs(4577) <= not b or a;
    layer2_outputs(4578) <= '0';
    layer2_outputs(4579) <= not b or a;
    layer2_outputs(4580) <= b and not a;
    layer2_outputs(4581) <= '1';
    layer2_outputs(4582) <= not a or b;
    layer2_outputs(4583) <= a;
    layer2_outputs(4584) <= not a;
    layer2_outputs(4585) <= a or b;
    layer2_outputs(4586) <= '0';
    layer2_outputs(4587) <= a or b;
    layer2_outputs(4588) <= not b;
    layer2_outputs(4589) <= not a;
    layer2_outputs(4590) <= a;
    layer2_outputs(4591) <= not (a or b);
    layer2_outputs(4592) <= '1';
    layer2_outputs(4593) <= not a;
    layer2_outputs(4594) <= '1';
    layer2_outputs(4595) <= b;
    layer2_outputs(4596) <= not a or b;
    layer2_outputs(4597) <= a and not b;
    layer2_outputs(4598) <= not b or a;
    layer2_outputs(4599) <= '1';
    layer2_outputs(4600) <= b;
    layer2_outputs(4601) <= '1';
    layer2_outputs(4602) <= not b or a;
    layer2_outputs(4603) <= not (a and b);
    layer2_outputs(4604) <= b and not a;
    layer2_outputs(4605) <= a or b;
    layer2_outputs(4606) <= a;
    layer2_outputs(4607) <= '1';
    layer2_outputs(4608) <= a;
    layer2_outputs(4609) <= not a;
    layer2_outputs(4610) <= a and not b;
    layer2_outputs(4611) <= not a or b;
    layer2_outputs(4612) <= not a;
    layer2_outputs(4613) <= not (a and b);
    layer2_outputs(4614) <= '0';
    layer2_outputs(4615) <= a and not b;
    layer2_outputs(4616) <= a and b;
    layer2_outputs(4617) <= a and not b;
    layer2_outputs(4618) <= a and not b;
    layer2_outputs(4619) <= not (a or b);
    layer2_outputs(4620) <= '0';
    layer2_outputs(4621) <= not b;
    layer2_outputs(4622) <= not a or b;
    layer2_outputs(4623) <= not a;
    layer2_outputs(4624) <= a and b;
    layer2_outputs(4625) <= a;
    layer2_outputs(4626) <= '1';
    layer2_outputs(4627) <= not (a and b);
    layer2_outputs(4628) <= not a or b;
    layer2_outputs(4629) <= a and not b;
    layer2_outputs(4630) <= a xor b;
    layer2_outputs(4631) <= not a or b;
    layer2_outputs(4632) <= not a or b;
    layer2_outputs(4633) <= a;
    layer2_outputs(4634) <= a;
    layer2_outputs(4635) <= not b or a;
    layer2_outputs(4636) <= '0';
    layer2_outputs(4637) <= '1';
    layer2_outputs(4638) <= '0';
    layer2_outputs(4639) <= a;
    layer2_outputs(4640) <= a and b;
    layer2_outputs(4641) <= not b or a;
    layer2_outputs(4642) <= b and not a;
    layer2_outputs(4643) <= not (a and b);
    layer2_outputs(4644) <= '1';
    layer2_outputs(4645) <= not a or b;
    layer2_outputs(4646) <= b and not a;
    layer2_outputs(4647) <= b;
    layer2_outputs(4648) <= not b;
    layer2_outputs(4649) <= not b or a;
    layer2_outputs(4650) <= a and not b;
    layer2_outputs(4651) <= a;
    layer2_outputs(4652) <= '0';
    layer2_outputs(4653) <= not a;
    layer2_outputs(4654) <= a;
    layer2_outputs(4655) <= not a;
    layer2_outputs(4656) <= b;
    layer2_outputs(4657) <= '0';
    layer2_outputs(4658) <= b and not a;
    layer2_outputs(4659) <= not b or a;
    layer2_outputs(4660) <= a;
    layer2_outputs(4661) <= '0';
    layer2_outputs(4662) <= a and not b;
    layer2_outputs(4663) <= not (a or b);
    layer2_outputs(4664) <= not a;
    layer2_outputs(4665) <= a or b;
    layer2_outputs(4666) <= a and not b;
    layer2_outputs(4667) <= not (a or b);
    layer2_outputs(4668) <= not a;
    layer2_outputs(4669) <= not (a and b);
    layer2_outputs(4670) <= a and not b;
    layer2_outputs(4671) <= '0';
    layer2_outputs(4672) <= b;
    layer2_outputs(4673) <= not b or a;
    layer2_outputs(4674) <= not (a and b);
    layer2_outputs(4675) <= b;
    layer2_outputs(4676) <= a and not b;
    layer2_outputs(4677) <= b and not a;
    layer2_outputs(4678) <= a and b;
    layer2_outputs(4679) <= not a;
    layer2_outputs(4680) <= not a or b;
    layer2_outputs(4681) <= not (a xor b);
    layer2_outputs(4682) <= b;
    layer2_outputs(4683) <= not b or a;
    layer2_outputs(4684) <= b;
    layer2_outputs(4685) <= a or b;
    layer2_outputs(4686) <= b and not a;
    layer2_outputs(4687) <= a or b;
    layer2_outputs(4688) <= a and b;
    layer2_outputs(4689) <= not a or b;
    layer2_outputs(4690) <= not a or b;
    layer2_outputs(4691) <= a;
    layer2_outputs(4692) <= not b or a;
    layer2_outputs(4693) <= '1';
    layer2_outputs(4694) <= not b;
    layer2_outputs(4695) <= not (a or b);
    layer2_outputs(4696) <= '1';
    layer2_outputs(4697) <= not (a or b);
    layer2_outputs(4698) <= not (a or b);
    layer2_outputs(4699) <= a and b;
    layer2_outputs(4700) <= not b;
    layer2_outputs(4701) <= '0';
    layer2_outputs(4702) <= a and b;
    layer2_outputs(4703) <= b and not a;
    layer2_outputs(4704) <= not (a xor b);
    layer2_outputs(4705) <= not a or b;
    layer2_outputs(4706) <= '0';
    layer2_outputs(4707) <= not (a or b);
    layer2_outputs(4708) <= not (a xor b);
    layer2_outputs(4709) <= '0';
    layer2_outputs(4710) <= b and not a;
    layer2_outputs(4711) <= a or b;
    layer2_outputs(4712) <= not a;
    layer2_outputs(4713) <= '0';
    layer2_outputs(4714) <= a xor b;
    layer2_outputs(4715) <= not a;
    layer2_outputs(4716) <= not (a and b);
    layer2_outputs(4717) <= not (a or b);
    layer2_outputs(4718) <= a and not b;
    layer2_outputs(4719) <= '1';
    layer2_outputs(4720) <= not a;
    layer2_outputs(4721) <= not (a and b);
    layer2_outputs(4722) <= not (a and b);
    layer2_outputs(4723) <= a;
    layer2_outputs(4724) <= not (a and b);
    layer2_outputs(4725) <= b;
    layer2_outputs(4726) <= not a;
    layer2_outputs(4727) <= not (a or b);
    layer2_outputs(4728) <= a and b;
    layer2_outputs(4729) <= '1';
    layer2_outputs(4730) <= '0';
    layer2_outputs(4731) <= not (a and b);
    layer2_outputs(4732) <= not (a and b);
    layer2_outputs(4733) <= not b;
    layer2_outputs(4734) <= not (a or b);
    layer2_outputs(4735) <= a or b;
    layer2_outputs(4736) <= a or b;
    layer2_outputs(4737) <= '1';
    layer2_outputs(4738) <= a;
    layer2_outputs(4739) <= a or b;
    layer2_outputs(4740) <= not (a and b);
    layer2_outputs(4741) <= not a or b;
    layer2_outputs(4742) <= not a;
    layer2_outputs(4743) <= a or b;
    layer2_outputs(4744) <= not (a or b);
    layer2_outputs(4745) <= a or b;
    layer2_outputs(4746) <= not (a and b);
    layer2_outputs(4747) <= a;
    layer2_outputs(4748) <= a and not b;
    layer2_outputs(4749) <= b;
    layer2_outputs(4750) <= not a;
    layer2_outputs(4751) <= '0';
    layer2_outputs(4752) <= a and b;
    layer2_outputs(4753) <= a and b;
    layer2_outputs(4754) <= not (a and b);
    layer2_outputs(4755) <= not b or a;
    layer2_outputs(4756) <= a;
    layer2_outputs(4757) <= a and not b;
    layer2_outputs(4758) <= not a;
    layer2_outputs(4759) <= a and not b;
    layer2_outputs(4760) <= b;
    layer2_outputs(4761) <= a or b;
    layer2_outputs(4762) <= not b or a;
    layer2_outputs(4763) <= '0';
    layer2_outputs(4764) <= b;
    layer2_outputs(4765) <= not (a or b);
    layer2_outputs(4766) <= not b;
    layer2_outputs(4767) <= not b or a;
    layer2_outputs(4768) <= a and not b;
    layer2_outputs(4769) <= '1';
    layer2_outputs(4770) <= not (a and b);
    layer2_outputs(4771) <= a or b;
    layer2_outputs(4772) <= a;
    layer2_outputs(4773) <= not b or a;
    layer2_outputs(4774) <= not (a or b);
    layer2_outputs(4775) <= b;
    layer2_outputs(4776) <= not b;
    layer2_outputs(4777) <= b;
    layer2_outputs(4778) <= b and not a;
    layer2_outputs(4779) <= a and not b;
    layer2_outputs(4780) <= a and b;
    layer2_outputs(4781) <= a;
    layer2_outputs(4782) <= not (a and b);
    layer2_outputs(4783) <= not b;
    layer2_outputs(4784) <= a or b;
    layer2_outputs(4785) <= not a or b;
    layer2_outputs(4786) <= a xor b;
    layer2_outputs(4787) <= not a or b;
    layer2_outputs(4788) <= b;
    layer2_outputs(4789) <= b and not a;
    layer2_outputs(4790) <= a and b;
    layer2_outputs(4791) <= a and not b;
    layer2_outputs(4792) <= not (a or b);
    layer2_outputs(4793) <= not a;
    layer2_outputs(4794) <= not (a and b);
    layer2_outputs(4795) <= not a or b;
    layer2_outputs(4796) <= not (a or b);
    layer2_outputs(4797) <= '0';
    layer2_outputs(4798) <= not a or b;
    layer2_outputs(4799) <= '0';
    layer2_outputs(4800) <= a and b;
    layer2_outputs(4801) <= '0';
    layer2_outputs(4802) <= '0';
    layer2_outputs(4803) <= not a or b;
    layer2_outputs(4804) <= a or b;
    layer2_outputs(4805) <= '0';
    layer2_outputs(4806) <= a;
    layer2_outputs(4807) <= '0';
    layer2_outputs(4808) <= '0';
    layer2_outputs(4809) <= not b or a;
    layer2_outputs(4810) <= b and not a;
    layer2_outputs(4811) <= a or b;
    layer2_outputs(4812) <= not a;
    layer2_outputs(4813) <= '0';
    layer2_outputs(4814) <= not a;
    layer2_outputs(4815) <= '0';
    layer2_outputs(4816) <= not a;
    layer2_outputs(4817) <= '0';
    layer2_outputs(4818) <= not (a and b);
    layer2_outputs(4819) <= '1';
    layer2_outputs(4820) <= not b;
    layer2_outputs(4821) <= '1';
    layer2_outputs(4822) <= not (a and b);
    layer2_outputs(4823) <= not b or a;
    layer2_outputs(4824) <= '1';
    layer2_outputs(4825) <= a;
    layer2_outputs(4826) <= a and b;
    layer2_outputs(4827) <= a and b;
    layer2_outputs(4828) <= b;
    layer2_outputs(4829) <= '0';
    layer2_outputs(4830) <= a and not b;
    layer2_outputs(4831) <= a or b;
    layer2_outputs(4832) <= a or b;
    layer2_outputs(4833) <= not a or b;
    layer2_outputs(4834) <= a and b;
    layer2_outputs(4835) <= '1';
    layer2_outputs(4836) <= not (a or b);
    layer2_outputs(4837) <= not b or a;
    layer2_outputs(4838) <= b;
    layer2_outputs(4839) <= not a or b;
    layer2_outputs(4840) <= not a;
    layer2_outputs(4841) <= not b;
    layer2_outputs(4842) <= not a;
    layer2_outputs(4843) <= not b;
    layer2_outputs(4844) <= b;
    layer2_outputs(4845) <= a;
    layer2_outputs(4846) <= a or b;
    layer2_outputs(4847) <= not b;
    layer2_outputs(4848) <= not (a and b);
    layer2_outputs(4849) <= '1';
    layer2_outputs(4850) <= b;
    layer2_outputs(4851) <= a and not b;
    layer2_outputs(4852) <= not b or a;
    layer2_outputs(4853) <= '0';
    layer2_outputs(4854) <= a and b;
    layer2_outputs(4855) <= not b;
    layer2_outputs(4856) <= '0';
    layer2_outputs(4857) <= b and not a;
    layer2_outputs(4858) <= not b or a;
    layer2_outputs(4859) <= a;
    layer2_outputs(4860) <= a or b;
    layer2_outputs(4861) <= a and not b;
    layer2_outputs(4862) <= not (a or b);
    layer2_outputs(4863) <= not (a and b);
    layer2_outputs(4864) <= a and b;
    layer2_outputs(4865) <= b and not a;
    layer2_outputs(4866) <= b;
    layer2_outputs(4867) <= '1';
    layer2_outputs(4868) <= '1';
    layer2_outputs(4869) <= a and not b;
    layer2_outputs(4870) <= not b;
    layer2_outputs(4871) <= not a or b;
    layer2_outputs(4872) <= a or b;
    layer2_outputs(4873) <= a or b;
    layer2_outputs(4874) <= not (a and b);
    layer2_outputs(4875) <= a;
    layer2_outputs(4876) <= '0';
    layer2_outputs(4877) <= not b;
    layer2_outputs(4878) <= a and b;
    layer2_outputs(4879) <= b;
    layer2_outputs(4880) <= a and not b;
    layer2_outputs(4881) <= '0';
    layer2_outputs(4882) <= b;
    layer2_outputs(4883) <= a and b;
    layer2_outputs(4884) <= b and not a;
    layer2_outputs(4885) <= a or b;
    layer2_outputs(4886) <= a and not b;
    layer2_outputs(4887) <= not (a and b);
    layer2_outputs(4888) <= a or b;
    layer2_outputs(4889) <= '1';
    layer2_outputs(4890) <= b and not a;
    layer2_outputs(4891) <= a and b;
    layer2_outputs(4892) <= not (a and b);
    layer2_outputs(4893) <= b;
    layer2_outputs(4894) <= a and b;
    layer2_outputs(4895) <= not (a or b);
    layer2_outputs(4896) <= '0';
    layer2_outputs(4897) <= not (a or b);
    layer2_outputs(4898) <= not a or b;
    layer2_outputs(4899) <= not b;
    layer2_outputs(4900) <= not (a or b);
    layer2_outputs(4901) <= not b or a;
    layer2_outputs(4902) <= not b or a;
    layer2_outputs(4903) <= a or b;
    layer2_outputs(4904) <= b and not a;
    layer2_outputs(4905) <= not a or b;
    layer2_outputs(4906) <= not b;
    layer2_outputs(4907) <= a;
    layer2_outputs(4908) <= '0';
    layer2_outputs(4909) <= b;
    layer2_outputs(4910) <= not (a or b);
    layer2_outputs(4911) <= not b;
    layer2_outputs(4912) <= not b or a;
    layer2_outputs(4913) <= not b;
    layer2_outputs(4914) <= '0';
    layer2_outputs(4915) <= not (a or b);
    layer2_outputs(4916) <= a and b;
    layer2_outputs(4917) <= '0';
    layer2_outputs(4918) <= b and not a;
    layer2_outputs(4919) <= '1';
    layer2_outputs(4920) <= not b or a;
    layer2_outputs(4921) <= b and not a;
    layer2_outputs(4922) <= b;
    layer2_outputs(4923) <= b and not a;
    layer2_outputs(4924) <= not a or b;
    layer2_outputs(4925) <= not b or a;
    layer2_outputs(4926) <= not (a and b);
    layer2_outputs(4927) <= a;
    layer2_outputs(4928) <= not b or a;
    layer2_outputs(4929) <= a and b;
    layer2_outputs(4930) <= not b;
    layer2_outputs(4931) <= not b or a;
    layer2_outputs(4932) <= not (a and b);
    layer2_outputs(4933) <= not b or a;
    layer2_outputs(4934) <= b;
    layer2_outputs(4935) <= not b or a;
    layer2_outputs(4936) <= not a;
    layer2_outputs(4937) <= '1';
    layer2_outputs(4938) <= not (a or b);
    layer2_outputs(4939) <= a;
    layer2_outputs(4940) <= '1';
    layer2_outputs(4941) <= not a;
    layer2_outputs(4942) <= '0';
    layer2_outputs(4943) <= b and not a;
    layer2_outputs(4944) <= '1';
    layer2_outputs(4945) <= not a;
    layer2_outputs(4946) <= b;
    layer2_outputs(4947) <= not a;
    layer2_outputs(4948) <= b;
    layer2_outputs(4949) <= a and b;
    layer2_outputs(4950) <= a or b;
    layer2_outputs(4951) <= a;
    layer2_outputs(4952) <= not b or a;
    layer2_outputs(4953) <= '1';
    layer2_outputs(4954) <= not b;
    layer2_outputs(4955) <= '0';
    layer2_outputs(4956) <= a;
    layer2_outputs(4957) <= not a;
    layer2_outputs(4958) <= not b or a;
    layer2_outputs(4959) <= not b or a;
    layer2_outputs(4960) <= not (a and b);
    layer2_outputs(4961) <= not a or b;
    layer2_outputs(4962) <= not b;
    layer2_outputs(4963) <= a or b;
    layer2_outputs(4964) <= '1';
    layer2_outputs(4965) <= not (a xor b);
    layer2_outputs(4966) <= not a;
    layer2_outputs(4967) <= '0';
    layer2_outputs(4968) <= b;
    layer2_outputs(4969) <= not b or a;
    layer2_outputs(4970) <= not a or b;
    layer2_outputs(4971) <= '1';
    layer2_outputs(4972) <= a or b;
    layer2_outputs(4973) <= '0';
    layer2_outputs(4974) <= not (a or b);
    layer2_outputs(4975) <= not (a and b);
    layer2_outputs(4976) <= b;
    layer2_outputs(4977) <= a or b;
    layer2_outputs(4978) <= '1';
    layer2_outputs(4979) <= not (a xor b);
    layer2_outputs(4980) <= a xor b;
    layer2_outputs(4981) <= not a or b;
    layer2_outputs(4982) <= not (a or b);
    layer2_outputs(4983) <= a and b;
    layer2_outputs(4984) <= not a;
    layer2_outputs(4985) <= not (a or b);
    layer2_outputs(4986) <= '1';
    layer2_outputs(4987) <= a or b;
    layer2_outputs(4988) <= not (a xor b);
    layer2_outputs(4989) <= b;
    layer2_outputs(4990) <= not (a or b);
    layer2_outputs(4991) <= a and not b;
    layer2_outputs(4992) <= not (a or b);
    layer2_outputs(4993) <= a and not b;
    layer2_outputs(4994) <= not b;
    layer2_outputs(4995) <= '0';
    layer2_outputs(4996) <= a and b;
    layer2_outputs(4997) <= not b or a;
    layer2_outputs(4998) <= not (a or b);
    layer2_outputs(4999) <= not a or b;
    layer2_outputs(5000) <= not b or a;
    layer2_outputs(5001) <= '0';
    layer2_outputs(5002) <= not (a xor b);
    layer2_outputs(5003) <= '1';
    layer2_outputs(5004) <= a and not b;
    layer2_outputs(5005) <= a and not b;
    layer2_outputs(5006) <= '1';
    layer2_outputs(5007) <= a xor b;
    layer2_outputs(5008) <= not (a and b);
    layer2_outputs(5009) <= not (a xor b);
    layer2_outputs(5010) <= not (a and b);
    layer2_outputs(5011) <= b;
    layer2_outputs(5012) <= b;
    layer2_outputs(5013) <= not (a or b);
    layer2_outputs(5014) <= not (a or b);
    layer2_outputs(5015) <= not a;
    layer2_outputs(5016) <= b and not a;
    layer2_outputs(5017) <= not (a and b);
    layer2_outputs(5018) <= not a;
    layer2_outputs(5019) <= '1';
    layer2_outputs(5020) <= a and not b;
    layer2_outputs(5021) <= a xor b;
    layer2_outputs(5022) <= not a;
    layer2_outputs(5023) <= a or b;
    layer2_outputs(5024) <= '0';
    layer2_outputs(5025) <= a xor b;
    layer2_outputs(5026) <= a or b;
    layer2_outputs(5027) <= not b;
    layer2_outputs(5028) <= a and not b;
    layer2_outputs(5029) <= a xor b;
    layer2_outputs(5030) <= b and not a;
    layer2_outputs(5031) <= not (a and b);
    layer2_outputs(5032) <= not a or b;
    layer2_outputs(5033) <= '1';
    layer2_outputs(5034) <= not a;
    layer2_outputs(5035) <= '0';
    layer2_outputs(5036) <= not a or b;
    layer2_outputs(5037) <= a or b;
    layer2_outputs(5038) <= not (a and b);
    layer2_outputs(5039) <= not a;
    layer2_outputs(5040) <= not (a or b);
    layer2_outputs(5041) <= b;
    layer2_outputs(5042) <= '1';
    layer2_outputs(5043) <= b and not a;
    layer2_outputs(5044) <= '0';
    layer2_outputs(5045) <= not a or b;
    layer2_outputs(5046) <= b;
    layer2_outputs(5047) <= b and not a;
    layer2_outputs(5048) <= b and not a;
    layer2_outputs(5049) <= not b or a;
    layer2_outputs(5050) <= not (a and b);
    layer2_outputs(5051) <= b and not a;
    layer2_outputs(5052) <= a and not b;
    layer2_outputs(5053) <= a and not b;
    layer2_outputs(5054) <= not (a or b);
    layer2_outputs(5055) <= not a;
    layer2_outputs(5056) <= not b or a;
    layer2_outputs(5057) <= a or b;
    layer2_outputs(5058) <= not a;
    layer2_outputs(5059) <= a;
    layer2_outputs(5060) <= '0';
    layer2_outputs(5061) <= a and b;
    layer2_outputs(5062) <= a and not b;
    layer2_outputs(5063) <= '1';
    layer2_outputs(5064) <= not (a or b);
    layer2_outputs(5065) <= not (a xor b);
    layer2_outputs(5066) <= '0';
    layer2_outputs(5067) <= not a;
    layer2_outputs(5068) <= not (a and b);
    layer2_outputs(5069) <= not b or a;
    layer2_outputs(5070) <= '1';
    layer2_outputs(5071) <= a;
    layer2_outputs(5072) <= not a or b;
    layer2_outputs(5073) <= b and not a;
    layer2_outputs(5074) <= not b or a;
    layer2_outputs(5075) <= not b or a;
    layer2_outputs(5076) <= a or b;
    layer2_outputs(5077) <= a and b;
    layer2_outputs(5078) <= b and not a;
    layer2_outputs(5079) <= a or b;
    layer2_outputs(5080) <= not a;
    layer2_outputs(5081) <= not a;
    layer2_outputs(5082) <= not (a or b);
    layer2_outputs(5083) <= not a;
    layer2_outputs(5084) <= '0';
    layer2_outputs(5085) <= a and b;
    layer2_outputs(5086) <= not (a xor b);
    layer2_outputs(5087) <= not b or a;
    layer2_outputs(5088) <= not b or a;
    layer2_outputs(5089) <= not (a or b);
    layer2_outputs(5090) <= a;
    layer2_outputs(5091) <= not (a or b);
    layer2_outputs(5092) <= '0';
    layer2_outputs(5093) <= a and not b;
    layer2_outputs(5094) <= a and not b;
    layer2_outputs(5095) <= not b or a;
    layer2_outputs(5096) <= not (a and b);
    layer2_outputs(5097) <= not b;
    layer2_outputs(5098) <= not (a or b);
    layer2_outputs(5099) <= a or b;
    layer2_outputs(5100) <= not b;
    layer2_outputs(5101) <= a xor b;
    layer2_outputs(5102) <= not b;
    layer2_outputs(5103) <= a and b;
    layer2_outputs(5104) <= b and not a;
    layer2_outputs(5105) <= a or b;
    layer2_outputs(5106) <= '0';
    layer2_outputs(5107) <= not a;
    layer2_outputs(5108) <= '0';
    layer2_outputs(5109) <= not (a and b);
    layer2_outputs(5110) <= not (a and b);
    layer2_outputs(5111) <= not b or a;
    layer2_outputs(5112) <= a or b;
    layer2_outputs(5113) <= not (a and b);
    layer2_outputs(5114) <= a;
    layer2_outputs(5115) <= '0';
    layer2_outputs(5116) <= '0';
    layer2_outputs(5117) <= b and not a;
    layer2_outputs(5118) <= not b or a;
    layer2_outputs(5119) <= b;
    layer3_outputs(0) <= not a;
    layer3_outputs(1) <= b and not a;
    layer3_outputs(2) <= b;
    layer3_outputs(3) <= a;
    layer3_outputs(4) <= '0';
    layer3_outputs(5) <= not (a or b);
    layer3_outputs(6) <= b;
    layer3_outputs(7) <= '1';
    layer3_outputs(8) <= a and b;
    layer3_outputs(9) <= not (a or b);
    layer3_outputs(10) <= a xor b;
    layer3_outputs(11) <= a and b;
    layer3_outputs(12) <= not (a or b);
    layer3_outputs(13) <= b;
    layer3_outputs(14) <= a and not b;
    layer3_outputs(15) <= a or b;
    layer3_outputs(16) <= not a or b;
    layer3_outputs(17) <= '0';
    layer3_outputs(18) <= not a or b;
    layer3_outputs(19) <= '0';
    layer3_outputs(20) <= not a or b;
    layer3_outputs(21) <= b;
    layer3_outputs(22) <= a or b;
    layer3_outputs(23) <= '1';
    layer3_outputs(24) <= not a or b;
    layer3_outputs(25) <= a xor b;
    layer3_outputs(26) <= '0';
    layer3_outputs(27) <= not (a or b);
    layer3_outputs(28) <= a and not b;
    layer3_outputs(29) <= b and not a;
    layer3_outputs(30) <= a and b;
    layer3_outputs(31) <= a or b;
    layer3_outputs(32) <= '0';
    layer3_outputs(33) <= not (a or b);
    layer3_outputs(34) <= a;
    layer3_outputs(35) <= not a or b;
    layer3_outputs(36) <= a or b;
    layer3_outputs(37) <= b and not a;
    layer3_outputs(38) <= a or b;
    layer3_outputs(39) <= a and b;
    layer3_outputs(40) <= a;
    layer3_outputs(41) <= a or b;
    layer3_outputs(42) <= not b;
    layer3_outputs(43) <= '0';
    layer3_outputs(44) <= not b or a;
    layer3_outputs(45) <= a and not b;
    layer3_outputs(46) <= not (a xor b);
    layer3_outputs(47) <= '0';
    layer3_outputs(48) <= not b;
    layer3_outputs(49) <= not b;
    layer3_outputs(50) <= a and b;
    layer3_outputs(51) <= not a or b;
    layer3_outputs(52) <= not a or b;
    layer3_outputs(53) <= not b;
    layer3_outputs(54) <= a;
    layer3_outputs(55) <= a;
    layer3_outputs(56) <= a;
    layer3_outputs(57) <= not b or a;
    layer3_outputs(58) <= a or b;
    layer3_outputs(59) <= a xor b;
    layer3_outputs(60) <= a;
    layer3_outputs(61) <= a and not b;
    layer3_outputs(62) <= not b;
    layer3_outputs(63) <= '0';
    layer3_outputs(64) <= not (a and b);
    layer3_outputs(65) <= '0';
    layer3_outputs(66) <= not (a xor b);
    layer3_outputs(67) <= not a or b;
    layer3_outputs(68) <= not (a or b);
    layer3_outputs(69) <= not b;
    layer3_outputs(70) <= not (a or b);
    layer3_outputs(71) <= b and not a;
    layer3_outputs(72) <= not (a xor b);
    layer3_outputs(73) <= b and not a;
    layer3_outputs(74) <= not (a and b);
    layer3_outputs(75) <= a and b;
    layer3_outputs(76) <= not a;
    layer3_outputs(77) <= not a;
    layer3_outputs(78) <= not (a or b);
    layer3_outputs(79) <= a and not b;
    layer3_outputs(80) <= not (a or b);
    layer3_outputs(81) <= not a or b;
    layer3_outputs(82) <= not (a xor b);
    layer3_outputs(83) <= not (a and b);
    layer3_outputs(84) <= a or b;
    layer3_outputs(85) <= b;
    layer3_outputs(86) <= '0';
    layer3_outputs(87) <= not (a xor b);
    layer3_outputs(88) <= not (a and b);
    layer3_outputs(89) <= b;
    layer3_outputs(90) <= a and not b;
    layer3_outputs(91) <= not a;
    layer3_outputs(92) <= a;
    layer3_outputs(93) <= not (a or b);
    layer3_outputs(94) <= '1';
    layer3_outputs(95) <= not b or a;
    layer3_outputs(96) <= not a or b;
    layer3_outputs(97) <= not (a or b);
    layer3_outputs(98) <= not b;
    layer3_outputs(99) <= not a or b;
    layer3_outputs(100) <= not (a or b);
    layer3_outputs(101) <= not (a and b);
    layer3_outputs(102) <= not b or a;
    layer3_outputs(103) <= a xor b;
    layer3_outputs(104) <= a xor b;
    layer3_outputs(105) <= b and not a;
    layer3_outputs(106) <= b and not a;
    layer3_outputs(107) <= not (a and b);
    layer3_outputs(108) <= b and not a;
    layer3_outputs(109) <= '1';
    layer3_outputs(110) <= not (a or b);
    layer3_outputs(111) <= not (a or b);
    layer3_outputs(112) <= not a;
    layer3_outputs(113) <= '0';
    layer3_outputs(114) <= a and b;
    layer3_outputs(115) <= not b or a;
    layer3_outputs(116) <= not a;
    layer3_outputs(117) <= not a;
    layer3_outputs(118) <= not a or b;
    layer3_outputs(119) <= not a;
    layer3_outputs(120) <= a;
    layer3_outputs(121) <= a;
    layer3_outputs(122) <= not (a xor b);
    layer3_outputs(123) <= a and not b;
    layer3_outputs(124) <= not b;
    layer3_outputs(125) <= '1';
    layer3_outputs(126) <= b;
    layer3_outputs(127) <= a and not b;
    layer3_outputs(128) <= b and not a;
    layer3_outputs(129) <= a and not b;
    layer3_outputs(130) <= a;
    layer3_outputs(131) <= a xor b;
    layer3_outputs(132) <= a xor b;
    layer3_outputs(133) <= not b;
    layer3_outputs(134) <= not a;
    layer3_outputs(135) <= a or b;
    layer3_outputs(136) <= b and not a;
    layer3_outputs(137) <= b and not a;
    layer3_outputs(138) <= a and not b;
    layer3_outputs(139) <= not (a and b);
    layer3_outputs(140) <= a and not b;
    layer3_outputs(141) <= '0';
    layer3_outputs(142) <= b;
    layer3_outputs(143) <= not a or b;
    layer3_outputs(144) <= not b;
    layer3_outputs(145) <= not b or a;
    layer3_outputs(146) <= '0';
    layer3_outputs(147) <= a and not b;
    layer3_outputs(148) <= not a;
    layer3_outputs(149) <= not (a and b);
    layer3_outputs(150) <= a;
    layer3_outputs(151) <= a and b;
    layer3_outputs(152) <= not b or a;
    layer3_outputs(153) <= not b;
    layer3_outputs(154) <= '1';
    layer3_outputs(155) <= a and b;
    layer3_outputs(156) <= not (a and b);
    layer3_outputs(157) <= not b or a;
    layer3_outputs(158) <= '0';
    layer3_outputs(159) <= a or b;
    layer3_outputs(160) <= a;
    layer3_outputs(161) <= a and b;
    layer3_outputs(162) <= '1';
    layer3_outputs(163) <= not a or b;
    layer3_outputs(164) <= not (a or b);
    layer3_outputs(165) <= not (a and b);
    layer3_outputs(166) <= a and b;
    layer3_outputs(167) <= a and b;
    layer3_outputs(168) <= not a or b;
    layer3_outputs(169) <= not a;
    layer3_outputs(170) <= a and not b;
    layer3_outputs(171) <= a or b;
    layer3_outputs(172) <= a and b;
    layer3_outputs(173) <= a;
    layer3_outputs(174) <= not b or a;
    layer3_outputs(175) <= a and b;
    layer3_outputs(176) <= not (a and b);
    layer3_outputs(177) <= a and not b;
    layer3_outputs(178) <= b and not a;
    layer3_outputs(179) <= not a;
    layer3_outputs(180) <= a and not b;
    layer3_outputs(181) <= b;
    layer3_outputs(182) <= b and not a;
    layer3_outputs(183) <= not a;
    layer3_outputs(184) <= '0';
    layer3_outputs(185) <= a;
    layer3_outputs(186) <= '0';
    layer3_outputs(187) <= not a;
    layer3_outputs(188) <= not b;
    layer3_outputs(189) <= not a or b;
    layer3_outputs(190) <= not b;
    layer3_outputs(191) <= b and not a;
    layer3_outputs(192) <= a and b;
    layer3_outputs(193) <= b and not a;
    layer3_outputs(194) <= not (a and b);
    layer3_outputs(195) <= b;
    layer3_outputs(196) <= not (a and b);
    layer3_outputs(197) <= not (a and b);
    layer3_outputs(198) <= a;
    layer3_outputs(199) <= not b or a;
    layer3_outputs(200) <= '0';
    layer3_outputs(201) <= b;
    layer3_outputs(202) <= a or b;
    layer3_outputs(203) <= b;
    layer3_outputs(204) <= a and b;
    layer3_outputs(205) <= b and not a;
    layer3_outputs(206) <= not a;
    layer3_outputs(207) <= a and b;
    layer3_outputs(208) <= b;
    layer3_outputs(209) <= not (a xor b);
    layer3_outputs(210) <= a or b;
    layer3_outputs(211) <= not b;
    layer3_outputs(212) <= a or b;
    layer3_outputs(213) <= '1';
    layer3_outputs(214) <= '0';
    layer3_outputs(215) <= a and not b;
    layer3_outputs(216) <= not b;
    layer3_outputs(217) <= not b or a;
    layer3_outputs(218) <= b;
    layer3_outputs(219) <= b and not a;
    layer3_outputs(220) <= b;
    layer3_outputs(221) <= '0';
    layer3_outputs(222) <= b and not a;
    layer3_outputs(223) <= not b or a;
    layer3_outputs(224) <= b;
    layer3_outputs(225) <= not b;
    layer3_outputs(226) <= a;
    layer3_outputs(227) <= b and not a;
    layer3_outputs(228) <= '1';
    layer3_outputs(229) <= not (a or b);
    layer3_outputs(230) <= not a;
    layer3_outputs(231) <= a and b;
    layer3_outputs(232) <= not (a xor b);
    layer3_outputs(233) <= not (a or b);
    layer3_outputs(234) <= '1';
    layer3_outputs(235) <= not (a or b);
    layer3_outputs(236) <= '0';
    layer3_outputs(237) <= a and b;
    layer3_outputs(238) <= not a or b;
    layer3_outputs(239) <= '1';
    layer3_outputs(240) <= a and b;
    layer3_outputs(241) <= b;
    layer3_outputs(242) <= '0';
    layer3_outputs(243) <= not a;
    layer3_outputs(244) <= not (a or b);
    layer3_outputs(245) <= not b;
    layer3_outputs(246) <= a or b;
    layer3_outputs(247) <= not b or a;
    layer3_outputs(248) <= not b or a;
    layer3_outputs(249) <= '0';
    layer3_outputs(250) <= not (a or b);
    layer3_outputs(251) <= not b or a;
    layer3_outputs(252) <= not (a or b);
    layer3_outputs(253) <= '1';
    layer3_outputs(254) <= not a;
    layer3_outputs(255) <= not (a or b);
    layer3_outputs(256) <= a or b;
    layer3_outputs(257) <= not (a and b);
    layer3_outputs(258) <= a and b;
    layer3_outputs(259) <= a and not b;
    layer3_outputs(260) <= a and b;
    layer3_outputs(261) <= b;
    layer3_outputs(262) <= not a or b;
    layer3_outputs(263) <= '1';
    layer3_outputs(264) <= a;
    layer3_outputs(265) <= '1';
    layer3_outputs(266) <= not a or b;
    layer3_outputs(267) <= a;
    layer3_outputs(268) <= not (a and b);
    layer3_outputs(269) <= b;
    layer3_outputs(270) <= not (a or b);
    layer3_outputs(271) <= not b or a;
    layer3_outputs(272) <= not (a or b);
    layer3_outputs(273) <= not (a xor b);
    layer3_outputs(274) <= a and b;
    layer3_outputs(275) <= b and not a;
    layer3_outputs(276) <= '1';
    layer3_outputs(277) <= b and not a;
    layer3_outputs(278) <= a and not b;
    layer3_outputs(279) <= a and b;
    layer3_outputs(280) <= not b;
    layer3_outputs(281) <= a and b;
    layer3_outputs(282) <= not a or b;
    layer3_outputs(283) <= not (a or b);
    layer3_outputs(284) <= not b;
    layer3_outputs(285) <= a;
    layer3_outputs(286) <= a and b;
    layer3_outputs(287) <= a and b;
    layer3_outputs(288) <= not a or b;
    layer3_outputs(289) <= not a;
    layer3_outputs(290) <= not a or b;
    layer3_outputs(291) <= '0';
    layer3_outputs(292) <= '1';
    layer3_outputs(293) <= a;
    layer3_outputs(294) <= '0';
    layer3_outputs(295) <= not (a and b);
    layer3_outputs(296) <= a and not b;
    layer3_outputs(297) <= '0';
    layer3_outputs(298) <= not a;
    layer3_outputs(299) <= not b or a;
    layer3_outputs(300) <= b;
    layer3_outputs(301) <= a and b;
    layer3_outputs(302) <= not a;
    layer3_outputs(303) <= not (a or b);
    layer3_outputs(304) <= a;
    layer3_outputs(305) <= '0';
    layer3_outputs(306) <= not a;
    layer3_outputs(307) <= b;
    layer3_outputs(308) <= not b or a;
    layer3_outputs(309) <= not b;
    layer3_outputs(310) <= a and b;
    layer3_outputs(311) <= not a;
    layer3_outputs(312) <= a and not b;
    layer3_outputs(313) <= '1';
    layer3_outputs(314) <= not a;
    layer3_outputs(315) <= a and b;
    layer3_outputs(316) <= b and not a;
    layer3_outputs(317) <= not b or a;
    layer3_outputs(318) <= a or b;
    layer3_outputs(319) <= not a;
    layer3_outputs(320) <= b and not a;
    layer3_outputs(321) <= '0';
    layer3_outputs(322) <= a xor b;
    layer3_outputs(323) <= b;
    layer3_outputs(324) <= not a;
    layer3_outputs(325) <= a and b;
    layer3_outputs(326) <= '1';
    layer3_outputs(327) <= not b;
    layer3_outputs(328) <= not b;
    layer3_outputs(329) <= not b or a;
    layer3_outputs(330) <= not (a or b);
    layer3_outputs(331) <= b;
    layer3_outputs(332) <= not a or b;
    layer3_outputs(333) <= not b or a;
    layer3_outputs(334) <= a or b;
    layer3_outputs(335) <= not b or a;
    layer3_outputs(336) <= a and b;
    layer3_outputs(337) <= a and not b;
    layer3_outputs(338) <= '0';
    layer3_outputs(339) <= not b;
    layer3_outputs(340) <= b;
    layer3_outputs(341) <= b and not a;
    layer3_outputs(342) <= not b or a;
    layer3_outputs(343) <= '1';
    layer3_outputs(344) <= '0';
    layer3_outputs(345) <= b;
    layer3_outputs(346) <= a and b;
    layer3_outputs(347) <= b and not a;
    layer3_outputs(348) <= not a or b;
    layer3_outputs(349) <= b and not a;
    layer3_outputs(350) <= not (a and b);
    layer3_outputs(351) <= not (a xor b);
    layer3_outputs(352) <= '1';
    layer3_outputs(353) <= a and not b;
    layer3_outputs(354) <= b and not a;
    layer3_outputs(355) <= a or b;
    layer3_outputs(356) <= not a or b;
    layer3_outputs(357) <= a and b;
    layer3_outputs(358) <= a;
    layer3_outputs(359) <= not b;
    layer3_outputs(360) <= b;
    layer3_outputs(361) <= b;
    layer3_outputs(362) <= a and not b;
    layer3_outputs(363) <= a;
    layer3_outputs(364) <= a and not b;
    layer3_outputs(365) <= a and not b;
    layer3_outputs(366) <= a or b;
    layer3_outputs(367) <= a and b;
    layer3_outputs(368) <= b and not a;
    layer3_outputs(369) <= not a or b;
    layer3_outputs(370) <= a;
    layer3_outputs(371) <= b;
    layer3_outputs(372) <= not a;
    layer3_outputs(373) <= not (a and b);
    layer3_outputs(374) <= a or b;
    layer3_outputs(375) <= a;
    layer3_outputs(376) <= not (a or b);
    layer3_outputs(377) <= not a or b;
    layer3_outputs(378) <= a and b;
    layer3_outputs(379) <= b and not a;
    layer3_outputs(380) <= '0';
    layer3_outputs(381) <= '0';
    layer3_outputs(382) <= not a;
    layer3_outputs(383) <= a and not b;
    layer3_outputs(384) <= b;
    layer3_outputs(385) <= not b or a;
    layer3_outputs(386) <= not (a xor b);
    layer3_outputs(387) <= not (a and b);
    layer3_outputs(388) <= a;
    layer3_outputs(389) <= not b;
    layer3_outputs(390) <= b and not a;
    layer3_outputs(391) <= '0';
    layer3_outputs(392) <= not (a or b);
    layer3_outputs(393) <= not a or b;
    layer3_outputs(394) <= a or b;
    layer3_outputs(395) <= '0';
    layer3_outputs(396) <= a and b;
    layer3_outputs(397) <= '0';
    layer3_outputs(398) <= a and not b;
    layer3_outputs(399) <= not (a and b);
    layer3_outputs(400) <= a;
    layer3_outputs(401) <= not (a or b);
    layer3_outputs(402) <= '0';
    layer3_outputs(403) <= b and not a;
    layer3_outputs(404) <= not (a and b);
    layer3_outputs(405) <= '1';
    layer3_outputs(406) <= not a or b;
    layer3_outputs(407) <= not (a xor b);
    layer3_outputs(408) <= not (a or b);
    layer3_outputs(409) <= a;
    layer3_outputs(410) <= '0';
    layer3_outputs(411) <= not a;
    layer3_outputs(412) <= b and not a;
    layer3_outputs(413) <= b and not a;
    layer3_outputs(414) <= not a or b;
    layer3_outputs(415) <= b and not a;
    layer3_outputs(416) <= not (a and b);
    layer3_outputs(417) <= not a;
    layer3_outputs(418) <= not (a and b);
    layer3_outputs(419) <= not (a and b);
    layer3_outputs(420) <= b and not a;
    layer3_outputs(421) <= not b;
    layer3_outputs(422) <= not a;
    layer3_outputs(423) <= not (a and b);
    layer3_outputs(424) <= b and not a;
    layer3_outputs(425) <= not (a and b);
    layer3_outputs(426) <= '0';
    layer3_outputs(427) <= '1';
    layer3_outputs(428) <= not (a and b);
    layer3_outputs(429) <= not a;
    layer3_outputs(430) <= a or b;
    layer3_outputs(431) <= a and b;
    layer3_outputs(432) <= b and not a;
    layer3_outputs(433) <= not a;
    layer3_outputs(434) <= '0';
    layer3_outputs(435) <= not b or a;
    layer3_outputs(436) <= '0';
    layer3_outputs(437) <= a and b;
    layer3_outputs(438) <= a;
    layer3_outputs(439) <= '0';
    layer3_outputs(440) <= a and not b;
    layer3_outputs(441) <= '0';
    layer3_outputs(442) <= a and not b;
    layer3_outputs(443) <= '1';
    layer3_outputs(444) <= a and b;
    layer3_outputs(445) <= a and b;
    layer3_outputs(446) <= not (a and b);
    layer3_outputs(447) <= not b;
    layer3_outputs(448) <= not a;
    layer3_outputs(449) <= not a;
    layer3_outputs(450) <= '0';
    layer3_outputs(451) <= '0';
    layer3_outputs(452) <= '0';
    layer3_outputs(453) <= a and b;
    layer3_outputs(454) <= a and b;
    layer3_outputs(455) <= not a or b;
    layer3_outputs(456) <= b;
    layer3_outputs(457) <= not (a or b);
    layer3_outputs(458) <= b and not a;
    layer3_outputs(459) <= not a;
    layer3_outputs(460) <= not (a or b);
    layer3_outputs(461) <= a and b;
    layer3_outputs(462) <= a xor b;
    layer3_outputs(463) <= a and not b;
    layer3_outputs(464) <= not (a and b);
    layer3_outputs(465) <= not b;
    layer3_outputs(466) <= b;
    layer3_outputs(467) <= not b or a;
    layer3_outputs(468) <= b and not a;
    layer3_outputs(469) <= not (a or b);
    layer3_outputs(470) <= '1';
    layer3_outputs(471) <= not b;
    layer3_outputs(472) <= not a or b;
    layer3_outputs(473) <= not (a or b);
    layer3_outputs(474) <= not (a and b);
    layer3_outputs(475) <= not (a and b);
    layer3_outputs(476) <= not (a or b);
    layer3_outputs(477) <= a and not b;
    layer3_outputs(478) <= '0';
    layer3_outputs(479) <= '1';
    layer3_outputs(480) <= a or b;
    layer3_outputs(481) <= a and b;
    layer3_outputs(482) <= a;
    layer3_outputs(483) <= a;
    layer3_outputs(484) <= not (a xor b);
    layer3_outputs(485) <= not (a and b);
    layer3_outputs(486) <= a or b;
    layer3_outputs(487) <= not a or b;
    layer3_outputs(488) <= b and not a;
    layer3_outputs(489) <= not (a xor b);
    layer3_outputs(490) <= '1';
    layer3_outputs(491) <= b and not a;
    layer3_outputs(492) <= not b or a;
    layer3_outputs(493) <= a or b;
    layer3_outputs(494) <= not b;
    layer3_outputs(495) <= '1';
    layer3_outputs(496) <= a xor b;
    layer3_outputs(497) <= not a or b;
    layer3_outputs(498) <= a or b;
    layer3_outputs(499) <= not b;
    layer3_outputs(500) <= a and b;
    layer3_outputs(501) <= a and b;
    layer3_outputs(502) <= not b or a;
    layer3_outputs(503) <= not (a and b);
    layer3_outputs(504) <= not a;
    layer3_outputs(505) <= not a or b;
    layer3_outputs(506) <= a and not b;
    layer3_outputs(507) <= not a;
    layer3_outputs(508) <= not (a or b);
    layer3_outputs(509) <= a or b;
    layer3_outputs(510) <= a and not b;
    layer3_outputs(511) <= b and not a;
    layer3_outputs(512) <= a and b;
    layer3_outputs(513) <= '0';
    layer3_outputs(514) <= not (a xor b);
    layer3_outputs(515) <= not a;
    layer3_outputs(516) <= b;
    layer3_outputs(517) <= not b;
    layer3_outputs(518) <= not (a and b);
    layer3_outputs(519) <= not a;
    layer3_outputs(520) <= not a;
    layer3_outputs(521) <= not b;
    layer3_outputs(522) <= b;
    layer3_outputs(523) <= not a or b;
    layer3_outputs(524) <= '0';
    layer3_outputs(525) <= b;
    layer3_outputs(526) <= b and not a;
    layer3_outputs(527) <= not (a or b);
    layer3_outputs(528) <= not (a and b);
    layer3_outputs(529) <= '1';
    layer3_outputs(530) <= b and not a;
    layer3_outputs(531) <= b and not a;
    layer3_outputs(532) <= b and not a;
    layer3_outputs(533) <= a and b;
    layer3_outputs(534) <= not (a and b);
    layer3_outputs(535) <= a;
    layer3_outputs(536) <= b;
    layer3_outputs(537) <= a;
    layer3_outputs(538) <= not b;
    layer3_outputs(539) <= not a or b;
    layer3_outputs(540) <= a xor b;
    layer3_outputs(541) <= '0';
    layer3_outputs(542) <= not (a or b);
    layer3_outputs(543) <= not b;
    layer3_outputs(544) <= not b;
    layer3_outputs(545) <= not a;
    layer3_outputs(546) <= a;
    layer3_outputs(547) <= not b;
    layer3_outputs(548) <= a and b;
    layer3_outputs(549) <= not (a or b);
    layer3_outputs(550) <= b;
    layer3_outputs(551) <= b and not a;
    layer3_outputs(552) <= not (a or b);
    layer3_outputs(553) <= b;
    layer3_outputs(554) <= a xor b;
    layer3_outputs(555) <= '0';
    layer3_outputs(556) <= not (a or b);
    layer3_outputs(557) <= b;
    layer3_outputs(558) <= a or b;
    layer3_outputs(559) <= not (a and b);
    layer3_outputs(560) <= not b;
    layer3_outputs(561) <= '0';
    layer3_outputs(562) <= b and not a;
    layer3_outputs(563) <= '1';
    layer3_outputs(564) <= a and not b;
    layer3_outputs(565) <= not a;
    layer3_outputs(566) <= not a;
    layer3_outputs(567) <= a and b;
    layer3_outputs(568) <= not (a or b);
    layer3_outputs(569) <= not (a and b);
    layer3_outputs(570) <= a or b;
    layer3_outputs(571) <= not (a and b);
    layer3_outputs(572) <= a xor b;
    layer3_outputs(573) <= not a;
    layer3_outputs(574) <= b;
    layer3_outputs(575) <= '1';
    layer3_outputs(576) <= not b or a;
    layer3_outputs(577) <= b;
    layer3_outputs(578) <= a or b;
    layer3_outputs(579) <= not a;
    layer3_outputs(580) <= not a;
    layer3_outputs(581) <= '0';
    layer3_outputs(582) <= '1';
    layer3_outputs(583) <= not (a and b);
    layer3_outputs(584) <= not a or b;
    layer3_outputs(585) <= a;
    layer3_outputs(586) <= a and not b;
    layer3_outputs(587) <= not a or b;
    layer3_outputs(588) <= '0';
    layer3_outputs(589) <= '0';
    layer3_outputs(590) <= not (a xor b);
    layer3_outputs(591) <= not b;
    layer3_outputs(592) <= b and not a;
    layer3_outputs(593) <= a and b;
    layer3_outputs(594) <= b;
    layer3_outputs(595) <= a and not b;
    layer3_outputs(596) <= a and not b;
    layer3_outputs(597) <= a and not b;
    layer3_outputs(598) <= not b;
    layer3_outputs(599) <= not a;
    layer3_outputs(600) <= b and not a;
    layer3_outputs(601) <= a and not b;
    layer3_outputs(602) <= a;
    layer3_outputs(603) <= a or b;
    layer3_outputs(604) <= a and b;
    layer3_outputs(605) <= b and not a;
    layer3_outputs(606) <= '1';
    layer3_outputs(607) <= '0';
    layer3_outputs(608) <= a and b;
    layer3_outputs(609) <= not a or b;
    layer3_outputs(610) <= not b;
    layer3_outputs(611) <= a and not b;
    layer3_outputs(612) <= not a or b;
    layer3_outputs(613) <= b and not a;
    layer3_outputs(614) <= '1';
    layer3_outputs(615) <= not (a or b);
    layer3_outputs(616) <= a or b;
    layer3_outputs(617) <= not b;
    layer3_outputs(618) <= not b or a;
    layer3_outputs(619) <= not (a or b);
    layer3_outputs(620) <= not (a and b);
    layer3_outputs(621) <= a;
    layer3_outputs(622) <= not a;
    layer3_outputs(623) <= not a or b;
    layer3_outputs(624) <= not a;
    layer3_outputs(625) <= not (a and b);
    layer3_outputs(626) <= b and not a;
    layer3_outputs(627) <= not (a or b);
    layer3_outputs(628) <= not b;
    layer3_outputs(629) <= b and not a;
    layer3_outputs(630) <= not b;
    layer3_outputs(631) <= b and not a;
    layer3_outputs(632) <= b and not a;
    layer3_outputs(633) <= a or b;
    layer3_outputs(634) <= '0';
    layer3_outputs(635) <= not b;
    layer3_outputs(636) <= not a or b;
    layer3_outputs(637) <= not a or b;
    layer3_outputs(638) <= not a or b;
    layer3_outputs(639) <= b;
    layer3_outputs(640) <= not (a and b);
    layer3_outputs(641) <= a;
    layer3_outputs(642) <= not a or b;
    layer3_outputs(643) <= a xor b;
    layer3_outputs(644) <= a;
    layer3_outputs(645) <= '1';
    layer3_outputs(646) <= not a;
    layer3_outputs(647) <= not (a and b);
    layer3_outputs(648) <= '0';
    layer3_outputs(649) <= a or b;
    layer3_outputs(650) <= a and b;
    layer3_outputs(651) <= b;
    layer3_outputs(652) <= a or b;
    layer3_outputs(653) <= a;
    layer3_outputs(654) <= '0';
    layer3_outputs(655) <= not b;
    layer3_outputs(656) <= not b or a;
    layer3_outputs(657) <= not (a or b);
    layer3_outputs(658) <= a;
    layer3_outputs(659) <= not (a and b);
    layer3_outputs(660) <= not a;
    layer3_outputs(661) <= not a;
    layer3_outputs(662) <= not b;
    layer3_outputs(663) <= not (a or b);
    layer3_outputs(664) <= a;
    layer3_outputs(665) <= not (a and b);
    layer3_outputs(666) <= not a or b;
    layer3_outputs(667) <= '1';
    layer3_outputs(668) <= b;
    layer3_outputs(669) <= not a;
    layer3_outputs(670) <= not b or a;
    layer3_outputs(671) <= not (a xor b);
    layer3_outputs(672) <= a and not b;
    layer3_outputs(673) <= not (a and b);
    layer3_outputs(674) <= '0';
    layer3_outputs(675) <= a and b;
    layer3_outputs(676) <= not b or a;
    layer3_outputs(677) <= not a;
    layer3_outputs(678) <= not (a or b);
    layer3_outputs(679) <= not (a and b);
    layer3_outputs(680) <= a or b;
    layer3_outputs(681) <= not a;
    layer3_outputs(682) <= '0';
    layer3_outputs(683) <= '1';
    layer3_outputs(684) <= not b or a;
    layer3_outputs(685) <= not (a or b);
    layer3_outputs(686) <= not b;
    layer3_outputs(687) <= a;
    layer3_outputs(688) <= a xor b;
    layer3_outputs(689) <= a or b;
    layer3_outputs(690) <= not (a or b);
    layer3_outputs(691) <= a and b;
    layer3_outputs(692) <= a xor b;
    layer3_outputs(693) <= a or b;
    layer3_outputs(694) <= not a or b;
    layer3_outputs(695) <= not (a or b);
    layer3_outputs(696) <= b;
    layer3_outputs(697) <= not (a or b);
    layer3_outputs(698) <= a and not b;
    layer3_outputs(699) <= not b;
    layer3_outputs(700) <= not a or b;
    layer3_outputs(701) <= a and not b;
    layer3_outputs(702) <= '1';
    layer3_outputs(703) <= not b;
    layer3_outputs(704) <= '0';
    layer3_outputs(705) <= not a;
    layer3_outputs(706) <= '0';
    layer3_outputs(707) <= b and not a;
    layer3_outputs(708) <= '1';
    layer3_outputs(709) <= b;
    layer3_outputs(710) <= a and not b;
    layer3_outputs(711) <= a and b;
    layer3_outputs(712) <= a;
    layer3_outputs(713) <= a and not b;
    layer3_outputs(714) <= not a;
    layer3_outputs(715) <= not a or b;
    layer3_outputs(716) <= not (a or b);
    layer3_outputs(717) <= a and b;
    layer3_outputs(718) <= b;
    layer3_outputs(719) <= '1';
    layer3_outputs(720) <= '0';
    layer3_outputs(721) <= not b;
    layer3_outputs(722) <= not a or b;
    layer3_outputs(723) <= not b;
    layer3_outputs(724) <= '0';
    layer3_outputs(725) <= '0';
    layer3_outputs(726) <= a;
    layer3_outputs(727) <= a and b;
    layer3_outputs(728) <= b and not a;
    layer3_outputs(729) <= not b or a;
    layer3_outputs(730) <= not b;
    layer3_outputs(731) <= b and not a;
    layer3_outputs(732) <= not b;
    layer3_outputs(733) <= not (a or b);
    layer3_outputs(734) <= '0';
    layer3_outputs(735) <= '1';
    layer3_outputs(736) <= '1';
    layer3_outputs(737) <= a;
    layer3_outputs(738) <= not a;
    layer3_outputs(739) <= a and not b;
    layer3_outputs(740) <= not a or b;
    layer3_outputs(741) <= '1';
    layer3_outputs(742) <= not b or a;
    layer3_outputs(743) <= '0';
    layer3_outputs(744) <= not b or a;
    layer3_outputs(745) <= '1';
    layer3_outputs(746) <= '0';
    layer3_outputs(747) <= not (a and b);
    layer3_outputs(748) <= b;
    layer3_outputs(749) <= a and not b;
    layer3_outputs(750) <= not (a or b);
    layer3_outputs(751) <= not a;
    layer3_outputs(752) <= not a or b;
    layer3_outputs(753) <= a and b;
    layer3_outputs(754) <= a;
    layer3_outputs(755) <= b;
    layer3_outputs(756) <= not (a or b);
    layer3_outputs(757) <= b and not a;
    layer3_outputs(758) <= b;
    layer3_outputs(759) <= not a;
    layer3_outputs(760) <= not a or b;
    layer3_outputs(761) <= not (a and b);
    layer3_outputs(762) <= b and not a;
    layer3_outputs(763) <= a;
    layer3_outputs(764) <= a and b;
    layer3_outputs(765) <= a and b;
    layer3_outputs(766) <= not b or a;
    layer3_outputs(767) <= '0';
    layer3_outputs(768) <= '0';
    layer3_outputs(769) <= a and b;
    layer3_outputs(770) <= not (a or b);
    layer3_outputs(771) <= not (a or b);
    layer3_outputs(772) <= not b or a;
    layer3_outputs(773) <= a and not b;
    layer3_outputs(774) <= b;
    layer3_outputs(775) <= not a or b;
    layer3_outputs(776) <= a;
    layer3_outputs(777) <= a and b;
    layer3_outputs(778) <= a and b;
    layer3_outputs(779) <= not (a xor b);
    layer3_outputs(780) <= not (a xor b);
    layer3_outputs(781) <= not b;
    layer3_outputs(782) <= not a;
    layer3_outputs(783) <= a and not b;
    layer3_outputs(784) <= '1';
    layer3_outputs(785) <= not a or b;
    layer3_outputs(786) <= a and b;
    layer3_outputs(787) <= a and b;
    layer3_outputs(788) <= not (a or b);
    layer3_outputs(789) <= not a;
    layer3_outputs(790) <= not (a and b);
    layer3_outputs(791) <= a and not b;
    layer3_outputs(792) <= not b or a;
    layer3_outputs(793) <= '0';
    layer3_outputs(794) <= b;
    layer3_outputs(795) <= a and not b;
    layer3_outputs(796) <= a xor b;
    layer3_outputs(797) <= a xor b;
    layer3_outputs(798) <= a;
    layer3_outputs(799) <= a and not b;
    layer3_outputs(800) <= b and not a;
    layer3_outputs(801) <= a and b;
    layer3_outputs(802) <= not b;
    layer3_outputs(803) <= b;
    layer3_outputs(804) <= '0';
    layer3_outputs(805) <= not a or b;
    layer3_outputs(806) <= a and b;
    layer3_outputs(807) <= not b or a;
    layer3_outputs(808) <= not a or b;
    layer3_outputs(809) <= not a;
    layer3_outputs(810) <= b and not a;
    layer3_outputs(811) <= a and not b;
    layer3_outputs(812) <= not b or a;
    layer3_outputs(813) <= not b;
    layer3_outputs(814) <= not a;
    layer3_outputs(815) <= '1';
    layer3_outputs(816) <= b;
    layer3_outputs(817) <= a and not b;
    layer3_outputs(818) <= a or b;
    layer3_outputs(819) <= not b;
    layer3_outputs(820) <= b;
    layer3_outputs(821) <= not (a or b);
    layer3_outputs(822) <= '0';
    layer3_outputs(823) <= '0';
    layer3_outputs(824) <= a xor b;
    layer3_outputs(825) <= '1';
    layer3_outputs(826) <= not (a or b);
    layer3_outputs(827) <= not b;
    layer3_outputs(828) <= a or b;
    layer3_outputs(829) <= not (a and b);
    layer3_outputs(830) <= b;
    layer3_outputs(831) <= not a or b;
    layer3_outputs(832) <= b;
    layer3_outputs(833) <= b and not a;
    layer3_outputs(834) <= not b;
    layer3_outputs(835) <= a or b;
    layer3_outputs(836) <= '1';
    layer3_outputs(837) <= not b;
    layer3_outputs(838) <= '0';
    layer3_outputs(839) <= '1';
    layer3_outputs(840) <= not a;
    layer3_outputs(841) <= b;
    layer3_outputs(842) <= '0';
    layer3_outputs(843) <= a;
    layer3_outputs(844) <= not a;
    layer3_outputs(845) <= b;
    layer3_outputs(846) <= a;
    layer3_outputs(847) <= b;
    layer3_outputs(848) <= not (a or b);
    layer3_outputs(849) <= b and not a;
    layer3_outputs(850) <= not a or b;
    layer3_outputs(851) <= not (a and b);
    layer3_outputs(852) <= a and not b;
    layer3_outputs(853) <= a xor b;
    layer3_outputs(854) <= a and not b;
    layer3_outputs(855) <= not a;
    layer3_outputs(856) <= not b;
    layer3_outputs(857) <= not b;
    layer3_outputs(858) <= not (a and b);
    layer3_outputs(859) <= not a or b;
    layer3_outputs(860) <= a and not b;
    layer3_outputs(861) <= a or b;
    layer3_outputs(862) <= a and not b;
    layer3_outputs(863) <= not b or a;
    layer3_outputs(864) <= not b;
    layer3_outputs(865) <= a or b;
    layer3_outputs(866) <= not a or b;
    layer3_outputs(867) <= not b or a;
    layer3_outputs(868) <= b and not a;
    layer3_outputs(869) <= a and not b;
    layer3_outputs(870) <= a and b;
    layer3_outputs(871) <= not (a and b);
    layer3_outputs(872) <= not b or a;
    layer3_outputs(873) <= not (a or b);
    layer3_outputs(874) <= a and b;
    layer3_outputs(875) <= b and not a;
    layer3_outputs(876) <= '0';
    layer3_outputs(877) <= '1';
    layer3_outputs(878) <= '0';
    layer3_outputs(879) <= b;
    layer3_outputs(880) <= a and b;
    layer3_outputs(881) <= '0';
    layer3_outputs(882) <= a;
    layer3_outputs(883) <= '1';
    layer3_outputs(884) <= b;
    layer3_outputs(885) <= not a or b;
    layer3_outputs(886) <= a;
    layer3_outputs(887) <= b and not a;
    layer3_outputs(888) <= not a or b;
    layer3_outputs(889) <= a and b;
    layer3_outputs(890) <= not (a and b);
    layer3_outputs(891) <= not a or b;
    layer3_outputs(892) <= not (a or b);
    layer3_outputs(893) <= a and not b;
    layer3_outputs(894) <= not (a or b);
    layer3_outputs(895) <= b;
    layer3_outputs(896) <= not a;
    layer3_outputs(897) <= a and b;
    layer3_outputs(898) <= a or b;
    layer3_outputs(899) <= '1';
    layer3_outputs(900) <= a and not b;
    layer3_outputs(901) <= a and b;
    layer3_outputs(902) <= not b or a;
    layer3_outputs(903) <= a or b;
    layer3_outputs(904) <= a xor b;
    layer3_outputs(905) <= not b;
    layer3_outputs(906) <= not (a and b);
    layer3_outputs(907) <= a and b;
    layer3_outputs(908) <= not b;
    layer3_outputs(909) <= a and not b;
    layer3_outputs(910) <= a and not b;
    layer3_outputs(911) <= not b;
    layer3_outputs(912) <= a or b;
    layer3_outputs(913) <= '0';
    layer3_outputs(914) <= '1';
    layer3_outputs(915) <= b and not a;
    layer3_outputs(916) <= '0';
    layer3_outputs(917) <= b;
    layer3_outputs(918) <= a and not b;
    layer3_outputs(919) <= b;
    layer3_outputs(920) <= b;
    layer3_outputs(921) <= a and b;
    layer3_outputs(922) <= a or b;
    layer3_outputs(923) <= a;
    layer3_outputs(924) <= not (a or b);
    layer3_outputs(925) <= b;
    layer3_outputs(926) <= not b;
    layer3_outputs(927) <= a and b;
    layer3_outputs(928) <= not b or a;
    layer3_outputs(929) <= a;
    layer3_outputs(930) <= not b or a;
    layer3_outputs(931) <= not a;
    layer3_outputs(932) <= not b;
    layer3_outputs(933) <= not b;
    layer3_outputs(934) <= not (a or b);
    layer3_outputs(935) <= '1';
    layer3_outputs(936) <= not a;
    layer3_outputs(937) <= a;
    layer3_outputs(938) <= not (a and b);
    layer3_outputs(939) <= not b;
    layer3_outputs(940) <= a and b;
    layer3_outputs(941) <= a or b;
    layer3_outputs(942) <= not a;
    layer3_outputs(943) <= a;
    layer3_outputs(944) <= b;
    layer3_outputs(945) <= b and not a;
    layer3_outputs(946) <= b;
    layer3_outputs(947) <= not a or b;
    layer3_outputs(948) <= b;
    layer3_outputs(949) <= a xor b;
    layer3_outputs(950) <= a;
    layer3_outputs(951) <= a or b;
    layer3_outputs(952) <= '1';
    layer3_outputs(953) <= not a or b;
    layer3_outputs(954) <= not a or b;
    layer3_outputs(955) <= a;
    layer3_outputs(956) <= not a or b;
    layer3_outputs(957) <= not (a and b);
    layer3_outputs(958) <= not b or a;
    layer3_outputs(959) <= a and not b;
    layer3_outputs(960) <= '0';
    layer3_outputs(961) <= not b or a;
    layer3_outputs(962) <= not (a xor b);
    layer3_outputs(963) <= '1';
    layer3_outputs(964) <= a and not b;
    layer3_outputs(965) <= b and not a;
    layer3_outputs(966) <= '0';
    layer3_outputs(967) <= '0';
    layer3_outputs(968) <= a and not b;
    layer3_outputs(969) <= '0';
    layer3_outputs(970) <= not (a or b);
    layer3_outputs(971) <= not (a xor b);
    layer3_outputs(972) <= not a or b;
    layer3_outputs(973) <= a and not b;
    layer3_outputs(974) <= not b or a;
    layer3_outputs(975) <= a xor b;
    layer3_outputs(976) <= not a;
    layer3_outputs(977) <= not a;
    layer3_outputs(978) <= a and b;
    layer3_outputs(979) <= b and not a;
    layer3_outputs(980) <= b and not a;
    layer3_outputs(981) <= a or b;
    layer3_outputs(982) <= not b;
    layer3_outputs(983) <= '0';
    layer3_outputs(984) <= not b;
    layer3_outputs(985) <= '1';
    layer3_outputs(986) <= '1';
    layer3_outputs(987) <= a xor b;
    layer3_outputs(988) <= not (a and b);
    layer3_outputs(989) <= not (a and b);
    layer3_outputs(990) <= a and not b;
    layer3_outputs(991) <= '1';
    layer3_outputs(992) <= '0';
    layer3_outputs(993) <= a or b;
    layer3_outputs(994) <= not a or b;
    layer3_outputs(995) <= a and b;
    layer3_outputs(996) <= not a or b;
    layer3_outputs(997) <= b and not a;
    layer3_outputs(998) <= not b;
    layer3_outputs(999) <= a and b;
    layer3_outputs(1000) <= not b or a;
    layer3_outputs(1001) <= not a;
    layer3_outputs(1002) <= a;
    layer3_outputs(1003) <= b;
    layer3_outputs(1004) <= a and b;
    layer3_outputs(1005) <= b and not a;
    layer3_outputs(1006) <= a and b;
    layer3_outputs(1007) <= not (a or b);
    layer3_outputs(1008) <= a or b;
    layer3_outputs(1009) <= not (a and b);
    layer3_outputs(1010) <= not b or a;
    layer3_outputs(1011) <= b and not a;
    layer3_outputs(1012) <= not b or a;
    layer3_outputs(1013) <= not (a or b);
    layer3_outputs(1014) <= b;
    layer3_outputs(1015) <= b;
    layer3_outputs(1016) <= '0';
    layer3_outputs(1017) <= not (a and b);
    layer3_outputs(1018) <= not b;
    layer3_outputs(1019) <= a and b;
    layer3_outputs(1020) <= b;
    layer3_outputs(1021) <= b;
    layer3_outputs(1022) <= a and b;
    layer3_outputs(1023) <= not b or a;
    layer3_outputs(1024) <= not a;
    layer3_outputs(1025) <= a or b;
    layer3_outputs(1026) <= a xor b;
    layer3_outputs(1027) <= not b or a;
    layer3_outputs(1028) <= a and not b;
    layer3_outputs(1029) <= a and b;
    layer3_outputs(1030) <= not (a and b);
    layer3_outputs(1031) <= a and b;
    layer3_outputs(1032) <= not b or a;
    layer3_outputs(1033) <= '0';
    layer3_outputs(1034) <= b;
    layer3_outputs(1035) <= not a or b;
    layer3_outputs(1036) <= a;
    layer3_outputs(1037) <= not b or a;
    layer3_outputs(1038) <= a and not b;
    layer3_outputs(1039) <= b and not a;
    layer3_outputs(1040) <= b and not a;
    layer3_outputs(1041) <= b and not a;
    layer3_outputs(1042) <= b;
    layer3_outputs(1043) <= '1';
    layer3_outputs(1044) <= a;
    layer3_outputs(1045) <= a xor b;
    layer3_outputs(1046) <= '0';
    layer3_outputs(1047) <= a and b;
    layer3_outputs(1048) <= '0';
    layer3_outputs(1049) <= a;
    layer3_outputs(1050) <= b and not a;
    layer3_outputs(1051) <= not b or a;
    layer3_outputs(1052) <= b;
    layer3_outputs(1053) <= b and not a;
    layer3_outputs(1054) <= '0';
    layer3_outputs(1055) <= not (a and b);
    layer3_outputs(1056) <= not b;
    layer3_outputs(1057) <= a or b;
    layer3_outputs(1058) <= a;
    layer3_outputs(1059) <= b and not a;
    layer3_outputs(1060) <= a;
    layer3_outputs(1061) <= b and not a;
    layer3_outputs(1062) <= '0';
    layer3_outputs(1063) <= a or b;
    layer3_outputs(1064) <= not (a and b);
    layer3_outputs(1065) <= '1';
    layer3_outputs(1066) <= not a;
    layer3_outputs(1067) <= a and not b;
    layer3_outputs(1068) <= a and b;
    layer3_outputs(1069) <= '1';
    layer3_outputs(1070) <= a and not b;
    layer3_outputs(1071) <= a and b;
    layer3_outputs(1072) <= not b or a;
    layer3_outputs(1073) <= not (a xor b);
    layer3_outputs(1074) <= b;
    layer3_outputs(1075) <= b and not a;
    layer3_outputs(1076) <= not a or b;
    layer3_outputs(1077) <= b and not a;
    layer3_outputs(1078) <= b and not a;
    layer3_outputs(1079) <= not a or b;
    layer3_outputs(1080) <= b;
    layer3_outputs(1081) <= '1';
    layer3_outputs(1082) <= not (a or b);
    layer3_outputs(1083) <= not b or a;
    layer3_outputs(1084) <= not (a xor b);
    layer3_outputs(1085) <= '0';
    layer3_outputs(1086) <= a and not b;
    layer3_outputs(1087) <= a and b;
    layer3_outputs(1088) <= '0';
    layer3_outputs(1089) <= not (a or b);
    layer3_outputs(1090) <= not a;
    layer3_outputs(1091) <= not (a or b);
    layer3_outputs(1092) <= a or b;
    layer3_outputs(1093) <= b and not a;
    layer3_outputs(1094) <= b and not a;
    layer3_outputs(1095) <= not (a and b);
    layer3_outputs(1096) <= a and not b;
    layer3_outputs(1097) <= not a;
    layer3_outputs(1098) <= not b or a;
    layer3_outputs(1099) <= '1';
    layer3_outputs(1100) <= '1';
    layer3_outputs(1101) <= '0';
    layer3_outputs(1102) <= not a;
    layer3_outputs(1103) <= not b or a;
    layer3_outputs(1104) <= '0';
    layer3_outputs(1105) <= not (a or b);
    layer3_outputs(1106) <= '0';
    layer3_outputs(1107) <= a and b;
    layer3_outputs(1108) <= a xor b;
    layer3_outputs(1109) <= '0';
    layer3_outputs(1110) <= a;
    layer3_outputs(1111) <= '1';
    layer3_outputs(1112) <= not b or a;
    layer3_outputs(1113) <= not (a and b);
    layer3_outputs(1114) <= not (a or b);
    layer3_outputs(1115) <= not a or b;
    layer3_outputs(1116) <= '0';
    layer3_outputs(1117) <= not a;
    layer3_outputs(1118) <= not b or a;
    layer3_outputs(1119) <= not (a xor b);
    layer3_outputs(1120) <= a;
    layer3_outputs(1121) <= '1';
    layer3_outputs(1122) <= b and not a;
    layer3_outputs(1123) <= '0';
    layer3_outputs(1124) <= '1';
    layer3_outputs(1125) <= not (a and b);
    layer3_outputs(1126) <= a or b;
    layer3_outputs(1127) <= '0';
    layer3_outputs(1128) <= not a or b;
    layer3_outputs(1129) <= b and not a;
    layer3_outputs(1130) <= b and not a;
    layer3_outputs(1131) <= not a or b;
    layer3_outputs(1132) <= a and not b;
    layer3_outputs(1133) <= a and b;
    layer3_outputs(1134) <= a;
    layer3_outputs(1135) <= a;
    layer3_outputs(1136) <= not a or b;
    layer3_outputs(1137) <= b;
    layer3_outputs(1138) <= a or b;
    layer3_outputs(1139) <= b and not a;
    layer3_outputs(1140) <= '0';
    layer3_outputs(1141) <= not (a or b);
    layer3_outputs(1142) <= not (a or b);
    layer3_outputs(1143) <= '1';
    layer3_outputs(1144) <= not a;
    layer3_outputs(1145) <= a and b;
    layer3_outputs(1146) <= not (a or b);
    layer3_outputs(1147) <= a xor b;
    layer3_outputs(1148) <= a or b;
    layer3_outputs(1149) <= a and b;
    layer3_outputs(1150) <= b;
    layer3_outputs(1151) <= '1';
    layer3_outputs(1152) <= not (a or b);
    layer3_outputs(1153) <= '1';
    layer3_outputs(1154) <= b and not a;
    layer3_outputs(1155) <= a and b;
    layer3_outputs(1156) <= not (a and b);
    layer3_outputs(1157) <= a and not b;
    layer3_outputs(1158) <= not (a and b);
    layer3_outputs(1159) <= not a or b;
    layer3_outputs(1160) <= a and b;
    layer3_outputs(1161) <= a and not b;
    layer3_outputs(1162) <= not b;
    layer3_outputs(1163) <= a and b;
    layer3_outputs(1164) <= not (a and b);
    layer3_outputs(1165) <= not (a and b);
    layer3_outputs(1166) <= a and b;
    layer3_outputs(1167) <= not a;
    layer3_outputs(1168) <= not (a xor b);
    layer3_outputs(1169) <= b and not a;
    layer3_outputs(1170) <= not (a or b);
    layer3_outputs(1171) <= not (a or b);
    layer3_outputs(1172) <= '0';
    layer3_outputs(1173) <= not b or a;
    layer3_outputs(1174) <= a and b;
    layer3_outputs(1175) <= b and not a;
    layer3_outputs(1176) <= a;
    layer3_outputs(1177) <= not b;
    layer3_outputs(1178) <= not (a and b);
    layer3_outputs(1179) <= '0';
    layer3_outputs(1180) <= a;
    layer3_outputs(1181) <= a or b;
    layer3_outputs(1182) <= a and not b;
    layer3_outputs(1183) <= not b;
    layer3_outputs(1184) <= '1';
    layer3_outputs(1185) <= '0';
    layer3_outputs(1186) <= a and not b;
    layer3_outputs(1187) <= not b;
    layer3_outputs(1188) <= a xor b;
    layer3_outputs(1189) <= not a or b;
    layer3_outputs(1190) <= a;
    layer3_outputs(1191) <= a and b;
    layer3_outputs(1192) <= '0';
    layer3_outputs(1193) <= not b or a;
    layer3_outputs(1194) <= not a;
    layer3_outputs(1195) <= a;
    layer3_outputs(1196) <= '1';
    layer3_outputs(1197) <= b and not a;
    layer3_outputs(1198) <= not (a and b);
    layer3_outputs(1199) <= not a;
    layer3_outputs(1200) <= not a or b;
    layer3_outputs(1201) <= b and not a;
    layer3_outputs(1202) <= '0';
    layer3_outputs(1203) <= not (a and b);
    layer3_outputs(1204) <= not b;
    layer3_outputs(1205) <= not (a xor b);
    layer3_outputs(1206) <= a or b;
    layer3_outputs(1207) <= not (a xor b);
    layer3_outputs(1208) <= b;
    layer3_outputs(1209) <= a or b;
    layer3_outputs(1210) <= a and b;
    layer3_outputs(1211) <= not (a or b);
    layer3_outputs(1212) <= '1';
    layer3_outputs(1213) <= '1';
    layer3_outputs(1214) <= b and not a;
    layer3_outputs(1215) <= not a;
    layer3_outputs(1216) <= b;
    layer3_outputs(1217) <= not a;
    layer3_outputs(1218) <= '0';
    layer3_outputs(1219) <= not b;
    layer3_outputs(1220) <= not (a and b);
    layer3_outputs(1221) <= not b;
    layer3_outputs(1222) <= a and not b;
    layer3_outputs(1223) <= not b or a;
    layer3_outputs(1224) <= b and not a;
    layer3_outputs(1225) <= a or b;
    layer3_outputs(1226) <= not (a and b);
    layer3_outputs(1227) <= not (a and b);
    layer3_outputs(1228) <= '0';
    layer3_outputs(1229) <= b;
    layer3_outputs(1230) <= a;
    layer3_outputs(1231) <= not (a or b);
    layer3_outputs(1232) <= not b or a;
    layer3_outputs(1233) <= '0';
    layer3_outputs(1234) <= b and not a;
    layer3_outputs(1235) <= not b;
    layer3_outputs(1236) <= a and b;
    layer3_outputs(1237) <= '1';
    layer3_outputs(1238) <= a and b;
    layer3_outputs(1239) <= not (a or b);
    layer3_outputs(1240) <= not (a and b);
    layer3_outputs(1241) <= not (a and b);
    layer3_outputs(1242) <= not b or a;
    layer3_outputs(1243) <= a and b;
    layer3_outputs(1244) <= not a or b;
    layer3_outputs(1245) <= a and b;
    layer3_outputs(1246) <= b and not a;
    layer3_outputs(1247) <= not a or b;
    layer3_outputs(1248) <= not b or a;
    layer3_outputs(1249) <= a and b;
    layer3_outputs(1250) <= b and not a;
    layer3_outputs(1251) <= a;
    layer3_outputs(1252) <= not b or a;
    layer3_outputs(1253) <= not a or b;
    layer3_outputs(1254) <= not a or b;
    layer3_outputs(1255) <= '0';
    layer3_outputs(1256) <= a and not b;
    layer3_outputs(1257) <= a and not b;
    layer3_outputs(1258) <= '0';
    layer3_outputs(1259) <= not (a or b);
    layer3_outputs(1260) <= '1';
    layer3_outputs(1261) <= a or b;
    layer3_outputs(1262) <= a and b;
    layer3_outputs(1263) <= not a or b;
    layer3_outputs(1264) <= a;
    layer3_outputs(1265) <= '0';
    layer3_outputs(1266) <= '1';
    layer3_outputs(1267) <= not (a or b);
    layer3_outputs(1268) <= b;
    layer3_outputs(1269) <= not (a or b);
    layer3_outputs(1270) <= not b;
    layer3_outputs(1271) <= not a;
    layer3_outputs(1272) <= not a;
    layer3_outputs(1273) <= '0';
    layer3_outputs(1274) <= not a or b;
    layer3_outputs(1275) <= not a;
    layer3_outputs(1276) <= a;
    layer3_outputs(1277) <= b and not a;
    layer3_outputs(1278) <= '1';
    layer3_outputs(1279) <= not a;
    layer3_outputs(1280) <= a and b;
    layer3_outputs(1281) <= not b or a;
    layer3_outputs(1282) <= not b or a;
    layer3_outputs(1283) <= a;
    layer3_outputs(1284) <= a and not b;
    layer3_outputs(1285) <= a;
    layer3_outputs(1286) <= not a or b;
    layer3_outputs(1287) <= not b;
    layer3_outputs(1288) <= b;
    layer3_outputs(1289) <= not a or b;
    layer3_outputs(1290) <= not b or a;
    layer3_outputs(1291) <= '1';
    layer3_outputs(1292) <= a and not b;
    layer3_outputs(1293) <= b and not a;
    layer3_outputs(1294) <= not b;
    layer3_outputs(1295) <= b;
    layer3_outputs(1296) <= not a or b;
    layer3_outputs(1297) <= not b;
    layer3_outputs(1298) <= not b or a;
    layer3_outputs(1299) <= a and b;
    layer3_outputs(1300) <= not b or a;
    layer3_outputs(1301) <= a and not b;
    layer3_outputs(1302) <= '0';
    layer3_outputs(1303) <= not a or b;
    layer3_outputs(1304) <= not b;
    layer3_outputs(1305) <= not a or b;
    layer3_outputs(1306) <= not a or b;
    layer3_outputs(1307) <= not b or a;
    layer3_outputs(1308) <= '1';
    layer3_outputs(1309) <= '1';
    layer3_outputs(1310) <= not a or b;
    layer3_outputs(1311) <= b;
    layer3_outputs(1312) <= a and not b;
    layer3_outputs(1313) <= b and not a;
    layer3_outputs(1314) <= a xor b;
    layer3_outputs(1315) <= a and b;
    layer3_outputs(1316) <= not b or a;
    layer3_outputs(1317) <= not b;
    layer3_outputs(1318) <= not a or b;
    layer3_outputs(1319) <= not b or a;
    layer3_outputs(1320) <= not a;
    layer3_outputs(1321) <= b;
    layer3_outputs(1322) <= not a;
    layer3_outputs(1323) <= not b;
    layer3_outputs(1324) <= not a;
    layer3_outputs(1325) <= not (a or b);
    layer3_outputs(1326) <= a and b;
    layer3_outputs(1327) <= not a;
    layer3_outputs(1328) <= '0';
    layer3_outputs(1329) <= a or b;
    layer3_outputs(1330) <= a and not b;
    layer3_outputs(1331) <= not a or b;
    layer3_outputs(1332) <= a and b;
    layer3_outputs(1333) <= not (a or b);
    layer3_outputs(1334) <= '0';
    layer3_outputs(1335) <= a and not b;
    layer3_outputs(1336) <= a and not b;
    layer3_outputs(1337) <= a and not b;
    layer3_outputs(1338) <= '1';
    layer3_outputs(1339) <= not b;
    layer3_outputs(1340) <= a or b;
    layer3_outputs(1341) <= a or b;
    layer3_outputs(1342) <= a and b;
    layer3_outputs(1343) <= not a or b;
    layer3_outputs(1344) <= not b;
    layer3_outputs(1345) <= '1';
    layer3_outputs(1346) <= not b;
    layer3_outputs(1347) <= b;
    layer3_outputs(1348) <= a;
    layer3_outputs(1349) <= '0';
    layer3_outputs(1350) <= not (a or b);
    layer3_outputs(1351) <= '0';
    layer3_outputs(1352) <= '0';
    layer3_outputs(1353) <= a and b;
    layer3_outputs(1354) <= a and b;
    layer3_outputs(1355) <= not b or a;
    layer3_outputs(1356) <= a and b;
    layer3_outputs(1357) <= '1';
    layer3_outputs(1358) <= not (a and b);
    layer3_outputs(1359) <= a;
    layer3_outputs(1360) <= not (a and b);
    layer3_outputs(1361) <= '1';
    layer3_outputs(1362) <= not b or a;
    layer3_outputs(1363) <= not a or b;
    layer3_outputs(1364) <= not (a xor b);
    layer3_outputs(1365) <= not b;
    layer3_outputs(1366) <= not b or a;
    layer3_outputs(1367) <= not a;
    layer3_outputs(1368) <= not a or b;
    layer3_outputs(1369) <= a and b;
    layer3_outputs(1370) <= '1';
    layer3_outputs(1371) <= '0';
    layer3_outputs(1372) <= a xor b;
    layer3_outputs(1373) <= b and not a;
    layer3_outputs(1374) <= a and not b;
    layer3_outputs(1375) <= not b;
    layer3_outputs(1376) <= not a;
    layer3_outputs(1377) <= not (a or b);
    layer3_outputs(1378) <= '1';
    layer3_outputs(1379) <= not (a and b);
    layer3_outputs(1380) <= a and b;
    layer3_outputs(1381) <= b;
    layer3_outputs(1382) <= a;
    layer3_outputs(1383) <= a and not b;
    layer3_outputs(1384) <= a and b;
    layer3_outputs(1385) <= not a or b;
    layer3_outputs(1386) <= not (a or b);
    layer3_outputs(1387) <= a xor b;
    layer3_outputs(1388) <= a and b;
    layer3_outputs(1389) <= a;
    layer3_outputs(1390) <= not (a and b);
    layer3_outputs(1391) <= a and not b;
    layer3_outputs(1392) <= a or b;
    layer3_outputs(1393) <= b and not a;
    layer3_outputs(1394) <= a and b;
    layer3_outputs(1395) <= b;
    layer3_outputs(1396) <= not (a and b);
    layer3_outputs(1397) <= not (a and b);
    layer3_outputs(1398) <= a;
    layer3_outputs(1399) <= not (a and b);
    layer3_outputs(1400) <= b;
    layer3_outputs(1401) <= not b;
    layer3_outputs(1402) <= a and not b;
    layer3_outputs(1403) <= '0';
    layer3_outputs(1404) <= not (a and b);
    layer3_outputs(1405) <= a and b;
    layer3_outputs(1406) <= '1';
    layer3_outputs(1407) <= a or b;
    layer3_outputs(1408) <= a or b;
    layer3_outputs(1409) <= '1';
    layer3_outputs(1410) <= not a or b;
    layer3_outputs(1411) <= '1';
    layer3_outputs(1412) <= a and not b;
    layer3_outputs(1413) <= not b;
    layer3_outputs(1414) <= b and not a;
    layer3_outputs(1415) <= b;
    layer3_outputs(1416) <= '0';
    layer3_outputs(1417) <= b and not a;
    layer3_outputs(1418) <= a and not b;
    layer3_outputs(1419) <= not a or b;
    layer3_outputs(1420) <= not a or b;
    layer3_outputs(1421) <= not a;
    layer3_outputs(1422) <= not (a or b);
    layer3_outputs(1423) <= b;
    layer3_outputs(1424) <= a and b;
    layer3_outputs(1425) <= '0';
    layer3_outputs(1426) <= not (a or b);
    layer3_outputs(1427) <= a and not b;
    layer3_outputs(1428) <= '0';
    layer3_outputs(1429) <= a xor b;
    layer3_outputs(1430) <= b and not a;
    layer3_outputs(1431) <= b and not a;
    layer3_outputs(1432) <= not (a or b);
    layer3_outputs(1433) <= '1';
    layer3_outputs(1434) <= a and not b;
    layer3_outputs(1435) <= not b;
    layer3_outputs(1436) <= '0';
    layer3_outputs(1437) <= not b or a;
    layer3_outputs(1438) <= a;
    layer3_outputs(1439) <= b;
    layer3_outputs(1440) <= not b;
    layer3_outputs(1441) <= not (a or b);
    layer3_outputs(1442) <= not (a and b);
    layer3_outputs(1443) <= not a or b;
    layer3_outputs(1444) <= not b;
    layer3_outputs(1445) <= b;
    layer3_outputs(1446) <= not b;
    layer3_outputs(1447) <= b and not a;
    layer3_outputs(1448) <= b and not a;
    layer3_outputs(1449) <= not (a or b);
    layer3_outputs(1450) <= b and not a;
    layer3_outputs(1451) <= a and b;
    layer3_outputs(1452) <= '0';
    layer3_outputs(1453) <= not a;
    layer3_outputs(1454) <= b;
    layer3_outputs(1455) <= a and not b;
    layer3_outputs(1456) <= '1';
    layer3_outputs(1457) <= not (a or b);
    layer3_outputs(1458) <= '1';
    layer3_outputs(1459) <= a;
    layer3_outputs(1460) <= not (a or b);
    layer3_outputs(1461) <= a and b;
    layer3_outputs(1462) <= a or b;
    layer3_outputs(1463) <= '1';
    layer3_outputs(1464) <= '1';
    layer3_outputs(1465) <= not a;
    layer3_outputs(1466) <= '1';
    layer3_outputs(1467) <= a or b;
    layer3_outputs(1468) <= not b;
    layer3_outputs(1469) <= a or b;
    layer3_outputs(1470) <= not (a and b);
    layer3_outputs(1471) <= b;
    layer3_outputs(1472) <= a;
    layer3_outputs(1473) <= '0';
    layer3_outputs(1474) <= not a or b;
    layer3_outputs(1475) <= not (a and b);
    layer3_outputs(1476) <= not a or b;
    layer3_outputs(1477) <= b and not a;
    layer3_outputs(1478) <= '1';
    layer3_outputs(1479) <= not (a and b);
    layer3_outputs(1480) <= b and not a;
    layer3_outputs(1481) <= b;
    layer3_outputs(1482) <= a and b;
    layer3_outputs(1483) <= not (a or b);
    layer3_outputs(1484) <= not (a or b);
    layer3_outputs(1485) <= a and not b;
    layer3_outputs(1486) <= a and not b;
    layer3_outputs(1487) <= not b;
    layer3_outputs(1488) <= not b or a;
    layer3_outputs(1489) <= not a or b;
    layer3_outputs(1490) <= not (a or b);
    layer3_outputs(1491) <= not a or b;
    layer3_outputs(1492) <= b;
    layer3_outputs(1493) <= '1';
    layer3_outputs(1494) <= a or b;
    layer3_outputs(1495) <= not (a and b);
    layer3_outputs(1496) <= not (a and b);
    layer3_outputs(1497) <= not (a or b);
    layer3_outputs(1498) <= a xor b;
    layer3_outputs(1499) <= a or b;
    layer3_outputs(1500) <= b and not a;
    layer3_outputs(1501) <= not b;
    layer3_outputs(1502) <= not (a and b);
    layer3_outputs(1503) <= a or b;
    layer3_outputs(1504) <= not a;
    layer3_outputs(1505) <= not a;
    layer3_outputs(1506) <= not (a and b);
    layer3_outputs(1507) <= a;
    layer3_outputs(1508) <= a or b;
    layer3_outputs(1509) <= b;
    layer3_outputs(1510) <= a or b;
    layer3_outputs(1511) <= not a or b;
    layer3_outputs(1512) <= a or b;
    layer3_outputs(1513) <= a and b;
    layer3_outputs(1514) <= '1';
    layer3_outputs(1515) <= a or b;
    layer3_outputs(1516) <= a;
    layer3_outputs(1517) <= not (a and b);
    layer3_outputs(1518) <= not b;
    layer3_outputs(1519) <= not b or a;
    layer3_outputs(1520) <= a;
    layer3_outputs(1521) <= not a or b;
    layer3_outputs(1522) <= a xor b;
    layer3_outputs(1523) <= b;
    layer3_outputs(1524) <= '0';
    layer3_outputs(1525) <= a and not b;
    layer3_outputs(1526) <= '0';
    layer3_outputs(1527) <= not a or b;
    layer3_outputs(1528) <= not (a xor b);
    layer3_outputs(1529) <= b and not a;
    layer3_outputs(1530) <= '0';
    layer3_outputs(1531) <= not b;
    layer3_outputs(1532) <= not (a and b);
    layer3_outputs(1533) <= not (a and b);
    layer3_outputs(1534) <= a and b;
    layer3_outputs(1535) <= '0';
    layer3_outputs(1536) <= not b or a;
    layer3_outputs(1537) <= a and not b;
    layer3_outputs(1538) <= '0';
    layer3_outputs(1539) <= '1';
    layer3_outputs(1540) <= not (a and b);
    layer3_outputs(1541) <= not (a and b);
    layer3_outputs(1542) <= not a;
    layer3_outputs(1543) <= not a or b;
    layer3_outputs(1544) <= a or b;
    layer3_outputs(1545) <= not (a and b);
    layer3_outputs(1546) <= not (a and b);
    layer3_outputs(1547) <= b and not a;
    layer3_outputs(1548) <= a and not b;
    layer3_outputs(1549) <= not b;
    layer3_outputs(1550) <= a and b;
    layer3_outputs(1551) <= a xor b;
    layer3_outputs(1552) <= '0';
    layer3_outputs(1553) <= not a or b;
    layer3_outputs(1554) <= not a;
    layer3_outputs(1555) <= b and not a;
    layer3_outputs(1556) <= a and not b;
    layer3_outputs(1557) <= '1';
    layer3_outputs(1558) <= not b or a;
    layer3_outputs(1559) <= b and not a;
    layer3_outputs(1560) <= not (a and b);
    layer3_outputs(1561) <= b;
    layer3_outputs(1562) <= not b;
    layer3_outputs(1563) <= not a or b;
    layer3_outputs(1564) <= not a;
    layer3_outputs(1565) <= not a or b;
    layer3_outputs(1566) <= b and not a;
    layer3_outputs(1567) <= '0';
    layer3_outputs(1568) <= a xor b;
    layer3_outputs(1569) <= not b;
    layer3_outputs(1570) <= b;
    layer3_outputs(1571) <= not b or a;
    layer3_outputs(1572) <= not b or a;
    layer3_outputs(1573) <= not (a and b);
    layer3_outputs(1574) <= b and not a;
    layer3_outputs(1575) <= '1';
    layer3_outputs(1576) <= '1';
    layer3_outputs(1577) <= not a;
    layer3_outputs(1578) <= '0';
    layer3_outputs(1579) <= '1';
    layer3_outputs(1580) <= b;
    layer3_outputs(1581) <= a and b;
    layer3_outputs(1582) <= b and not a;
    layer3_outputs(1583) <= b and not a;
    layer3_outputs(1584) <= a;
    layer3_outputs(1585) <= not b or a;
    layer3_outputs(1586) <= b and not a;
    layer3_outputs(1587) <= not (a and b);
    layer3_outputs(1588) <= '1';
    layer3_outputs(1589) <= a and b;
    layer3_outputs(1590) <= a and not b;
    layer3_outputs(1591) <= not b or a;
    layer3_outputs(1592) <= a and b;
    layer3_outputs(1593) <= '1';
    layer3_outputs(1594) <= a or b;
    layer3_outputs(1595) <= a;
    layer3_outputs(1596) <= b and not a;
    layer3_outputs(1597) <= a;
    layer3_outputs(1598) <= not (a and b);
    layer3_outputs(1599) <= a and b;
    layer3_outputs(1600) <= a xor b;
    layer3_outputs(1601) <= '0';
    layer3_outputs(1602) <= b and not a;
    layer3_outputs(1603) <= not b or a;
    layer3_outputs(1604) <= a and not b;
    layer3_outputs(1605) <= not a or b;
    layer3_outputs(1606) <= a and b;
    layer3_outputs(1607) <= b and not a;
    layer3_outputs(1608) <= not a;
    layer3_outputs(1609) <= '1';
    layer3_outputs(1610) <= a and b;
    layer3_outputs(1611) <= b;
    layer3_outputs(1612) <= b;
    layer3_outputs(1613) <= a or b;
    layer3_outputs(1614) <= not b;
    layer3_outputs(1615) <= a or b;
    layer3_outputs(1616) <= '1';
    layer3_outputs(1617) <= a and b;
    layer3_outputs(1618) <= '0';
    layer3_outputs(1619) <= not (a and b);
    layer3_outputs(1620) <= not b;
    layer3_outputs(1621) <= a xor b;
    layer3_outputs(1622) <= not a;
    layer3_outputs(1623) <= a;
    layer3_outputs(1624) <= a;
    layer3_outputs(1625) <= a and b;
    layer3_outputs(1626) <= not (a or b);
    layer3_outputs(1627) <= not a;
    layer3_outputs(1628) <= not a or b;
    layer3_outputs(1629) <= a and b;
    layer3_outputs(1630) <= not a or b;
    layer3_outputs(1631) <= a or b;
    layer3_outputs(1632) <= a;
    layer3_outputs(1633) <= b and not a;
    layer3_outputs(1634) <= not (a and b);
    layer3_outputs(1635) <= not a or b;
    layer3_outputs(1636) <= not (a and b);
    layer3_outputs(1637) <= not a or b;
    layer3_outputs(1638) <= not (a and b);
    layer3_outputs(1639) <= a and b;
    layer3_outputs(1640) <= not b or a;
    layer3_outputs(1641) <= b;
    layer3_outputs(1642) <= not b;
    layer3_outputs(1643) <= a or b;
    layer3_outputs(1644) <= a and b;
    layer3_outputs(1645) <= not b;
    layer3_outputs(1646) <= not b;
    layer3_outputs(1647) <= not (a or b);
    layer3_outputs(1648) <= a and b;
    layer3_outputs(1649) <= b;
    layer3_outputs(1650) <= a;
    layer3_outputs(1651) <= a and not b;
    layer3_outputs(1652) <= b;
    layer3_outputs(1653) <= not a;
    layer3_outputs(1654) <= not a;
    layer3_outputs(1655) <= a and b;
    layer3_outputs(1656) <= '1';
    layer3_outputs(1657) <= not a or b;
    layer3_outputs(1658) <= a xor b;
    layer3_outputs(1659) <= not (a xor b);
    layer3_outputs(1660) <= a and not b;
    layer3_outputs(1661) <= not a;
    layer3_outputs(1662) <= not b;
    layer3_outputs(1663) <= '0';
    layer3_outputs(1664) <= not b or a;
    layer3_outputs(1665) <= not (a or b);
    layer3_outputs(1666) <= '0';
    layer3_outputs(1667) <= not (a or b);
    layer3_outputs(1668) <= '1';
    layer3_outputs(1669) <= not (a and b);
    layer3_outputs(1670) <= not b;
    layer3_outputs(1671) <= not (a or b);
    layer3_outputs(1672) <= not b or a;
    layer3_outputs(1673) <= a;
    layer3_outputs(1674) <= not (a and b);
    layer3_outputs(1675) <= b;
    layer3_outputs(1676) <= b;
    layer3_outputs(1677) <= a;
    layer3_outputs(1678) <= not a;
    layer3_outputs(1679) <= a;
    layer3_outputs(1680) <= '1';
    layer3_outputs(1681) <= not b or a;
    layer3_outputs(1682) <= not a;
    layer3_outputs(1683) <= not (a or b);
    layer3_outputs(1684) <= a and not b;
    layer3_outputs(1685) <= not a;
    layer3_outputs(1686) <= '1';
    layer3_outputs(1687) <= '1';
    layer3_outputs(1688) <= b and not a;
    layer3_outputs(1689) <= a and not b;
    layer3_outputs(1690) <= a and b;
    layer3_outputs(1691) <= not (a and b);
    layer3_outputs(1692) <= b;
    layer3_outputs(1693) <= a;
    layer3_outputs(1694) <= a;
    layer3_outputs(1695) <= not a or b;
    layer3_outputs(1696) <= b and not a;
    layer3_outputs(1697) <= a and b;
    layer3_outputs(1698) <= a and not b;
    layer3_outputs(1699) <= '1';
    layer3_outputs(1700) <= not b;
    layer3_outputs(1701) <= not a or b;
    layer3_outputs(1702) <= '1';
    layer3_outputs(1703) <= not a or b;
    layer3_outputs(1704) <= not (a and b);
    layer3_outputs(1705) <= '1';
    layer3_outputs(1706) <= a and not b;
    layer3_outputs(1707) <= a;
    layer3_outputs(1708) <= not (a and b);
    layer3_outputs(1709) <= not b or a;
    layer3_outputs(1710) <= a and b;
    layer3_outputs(1711) <= not b or a;
    layer3_outputs(1712) <= a or b;
    layer3_outputs(1713) <= not b;
    layer3_outputs(1714) <= b and not a;
    layer3_outputs(1715) <= not b or a;
    layer3_outputs(1716) <= b;
    layer3_outputs(1717) <= not (a and b);
    layer3_outputs(1718) <= a or b;
    layer3_outputs(1719) <= not (a xor b);
    layer3_outputs(1720) <= b and not a;
    layer3_outputs(1721) <= a;
    layer3_outputs(1722) <= not a;
    layer3_outputs(1723) <= b and not a;
    layer3_outputs(1724) <= not b;
    layer3_outputs(1725) <= not (a and b);
    layer3_outputs(1726) <= a;
    layer3_outputs(1727) <= not a or b;
    layer3_outputs(1728) <= not a or b;
    layer3_outputs(1729) <= '0';
    layer3_outputs(1730) <= a;
    layer3_outputs(1731) <= not b;
    layer3_outputs(1732) <= not b;
    layer3_outputs(1733) <= not a;
    layer3_outputs(1734) <= a;
    layer3_outputs(1735) <= a or b;
    layer3_outputs(1736) <= a;
    layer3_outputs(1737) <= '0';
    layer3_outputs(1738) <= a and not b;
    layer3_outputs(1739) <= not b or a;
    layer3_outputs(1740) <= a or b;
    layer3_outputs(1741) <= '0';
    layer3_outputs(1742) <= not a or b;
    layer3_outputs(1743) <= b;
    layer3_outputs(1744) <= not (a and b);
    layer3_outputs(1745) <= a;
    layer3_outputs(1746) <= not b;
    layer3_outputs(1747) <= a;
    layer3_outputs(1748) <= a or b;
    layer3_outputs(1749) <= a;
    layer3_outputs(1750) <= '0';
    layer3_outputs(1751) <= not b;
    layer3_outputs(1752) <= a and not b;
    layer3_outputs(1753) <= b;
    layer3_outputs(1754) <= b;
    layer3_outputs(1755) <= not a;
    layer3_outputs(1756) <= a;
    layer3_outputs(1757) <= not (a or b);
    layer3_outputs(1758) <= not b or a;
    layer3_outputs(1759) <= '0';
    layer3_outputs(1760) <= not (a or b);
    layer3_outputs(1761) <= b and not a;
    layer3_outputs(1762) <= b and not a;
    layer3_outputs(1763) <= b and not a;
    layer3_outputs(1764) <= not b or a;
    layer3_outputs(1765) <= a or b;
    layer3_outputs(1766) <= a and not b;
    layer3_outputs(1767) <= not b;
    layer3_outputs(1768) <= b and not a;
    layer3_outputs(1769) <= '0';
    layer3_outputs(1770) <= b;
    layer3_outputs(1771) <= a xor b;
    layer3_outputs(1772) <= a;
    layer3_outputs(1773) <= not (a xor b);
    layer3_outputs(1774) <= not b;
    layer3_outputs(1775) <= '0';
    layer3_outputs(1776) <= a and b;
    layer3_outputs(1777) <= not b;
    layer3_outputs(1778) <= a;
    layer3_outputs(1779) <= not b;
    layer3_outputs(1780) <= '1';
    layer3_outputs(1781) <= a and b;
    layer3_outputs(1782) <= '1';
    layer3_outputs(1783) <= not a or b;
    layer3_outputs(1784) <= b;
    layer3_outputs(1785) <= not (a or b);
    layer3_outputs(1786) <= not a;
    layer3_outputs(1787) <= a and not b;
    layer3_outputs(1788) <= a and b;
    layer3_outputs(1789) <= b;
    layer3_outputs(1790) <= '0';
    layer3_outputs(1791) <= '0';
    layer3_outputs(1792) <= a and b;
    layer3_outputs(1793) <= b;
    layer3_outputs(1794) <= '1';
    layer3_outputs(1795) <= not (a and b);
    layer3_outputs(1796) <= not a;
    layer3_outputs(1797) <= not a or b;
    layer3_outputs(1798) <= not (a or b);
    layer3_outputs(1799) <= not b or a;
    layer3_outputs(1800) <= '1';
    layer3_outputs(1801) <= a and not b;
    layer3_outputs(1802) <= a or b;
    layer3_outputs(1803) <= b;
    layer3_outputs(1804) <= a and b;
    layer3_outputs(1805) <= not (a and b);
    layer3_outputs(1806) <= a;
    layer3_outputs(1807) <= a or b;
    layer3_outputs(1808) <= '1';
    layer3_outputs(1809) <= a;
    layer3_outputs(1810) <= not (a xor b);
    layer3_outputs(1811) <= '0';
    layer3_outputs(1812) <= '1';
    layer3_outputs(1813) <= a;
    layer3_outputs(1814) <= b;
    layer3_outputs(1815) <= '1';
    layer3_outputs(1816) <= a;
    layer3_outputs(1817) <= a and not b;
    layer3_outputs(1818) <= a and not b;
    layer3_outputs(1819) <= not (a and b);
    layer3_outputs(1820) <= '0';
    layer3_outputs(1821) <= not (a or b);
    layer3_outputs(1822) <= b;
    layer3_outputs(1823) <= '1';
    layer3_outputs(1824) <= '0';
    layer3_outputs(1825) <= not (a or b);
    layer3_outputs(1826) <= b and not a;
    layer3_outputs(1827) <= '0';
    layer3_outputs(1828) <= b and not a;
    layer3_outputs(1829) <= not (a and b);
    layer3_outputs(1830) <= not a or b;
    layer3_outputs(1831) <= '1';
    layer3_outputs(1832) <= not a or b;
    layer3_outputs(1833) <= b;
    layer3_outputs(1834) <= not (a xor b);
    layer3_outputs(1835) <= not (a or b);
    layer3_outputs(1836) <= a or b;
    layer3_outputs(1837) <= b and not a;
    layer3_outputs(1838) <= a and b;
    layer3_outputs(1839) <= a and not b;
    layer3_outputs(1840) <= '1';
    layer3_outputs(1841) <= not (a or b);
    layer3_outputs(1842) <= not (a or b);
    layer3_outputs(1843) <= not (a and b);
    layer3_outputs(1844) <= a and b;
    layer3_outputs(1845) <= not a;
    layer3_outputs(1846) <= a and b;
    layer3_outputs(1847) <= '1';
    layer3_outputs(1848) <= not a or b;
    layer3_outputs(1849) <= not (a or b);
    layer3_outputs(1850) <= not a;
    layer3_outputs(1851) <= b and not a;
    layer3_outputs(1852) <= '1';
    layer3_outputs(1853) <= not b or a;
    layer3_outputs(1854) <= not (a and b);
    layer3_outputs(1855) <= a or b;
    layer3_outputs(1856) <= not a;
    layer3_outputs(1857) <= a and not b;
    layer3_outputs(1858) <= b and not a;
    layer3_outputs(1859) <= not b;
    layer3_outputs(1860) <= '1';
    layer3_outputs(1861) <= not a;
    layer3_outputs(1862) <= b and not a;
    layer3_outputs(1863) <= not b or a;
    layer3_outputs(1864) <= not a;
    layer3_outputs(1865) <= not b or a;
    layer3_outputs(1866) <= '0';
    layer3_outputs(1867) <= not a;
    layer3_outputs(1868) <= '0';
    layer3_outputs(1869) <= a xor b;
    layer3_outputs(1870) <= a or b;
    layer3_outputs(1871) <= not (a and b);
    layer3_outputs(1872) <= not (a and b);
    layer3_outputs(1873) <= '1';
    layer3_outputs(1874) <= a;
    layer3_outputs(1875) <= not (a or b);
    layer3_outputs(1876) <= '0';
    layer3_outputs(1877) <= not (a or b);
    layer3_outputs(1878) <= b and not a;
    layer3_outputs(1879) <= '1';
    layer3_outputs(1880) <= '0';
    layer3_outputs(1881) <= not (a or b);
    layer3_outputs(1882) <= a and b;
    layer3_outputs(1883) <= b and not a;
    layer3_outputs(1884) <= b;
    layer3_outputs(1885) <= not a or b;
    layer3_outputs(1886) <= '1';
    layer3_outputs(1887) <= not (a or b);
    layer3_outputs(1888) <= a or b;
    layer3_outputs(1889) <= not a or b;
    layer3_outputs(1890) <= not b or a;
    layer3_outputs(1891) <= '0';
    layer3_outputs(1892) <= b and not a;
    layer3_outputs(1893) <= a or b;
    layer3_outputs(1894) <= not a;
    layer3_outputs(1895) <= a or b;
    layer3_outputs(1896) <= b;
    layer3_outputs(1897) <= a and b;
    layer3_outputs(1898) <= a or b;
    layer3_outputs(1899) <= not (a or b);
    layer3_outputs(1900) <= a or b;
    layer3_outputs(1901) <= '0';
    layer3_outputs(1902) <= a and not b;
    layer3_outputs(1903) <= not (a and b);
    layer3_outputs(1904) <= not a or b;
    layer3_outputs(1905) <= '1';
    layer3_outputs(1906) <= a and b;
    layer3_outputs(1907) <= not a or b;
    layer3_outputs(1908) <= not b or a;
    layer3_outputs(1909) <= '1';
    layer3_outputs(1910) <= a and not b;
    layer3_outputs(1911) <= '1';
    layer3_outputs(1912) <= a;
    layer3_outputs(1913) <= '1';
    layer3_outputs(1914) <= not b;
    layer3_outputs(1915) <= not (a or b);
    layer3_outputs(1916) <= not (a or b);
    layer3_outputs(1917) <= a and not b;
    layer3_outputs(1918) <= '1';
    layer3_outputs(1919) <= '0';
    layer3_outputs(1920) <= a and b;
    layer3_outputs(1921) <= a and b;
    layer3_outputs(1922) <= a and not b;
    layer3_outputs(1923) <= b;
    layer3_outputs(1924) <= '0';
    layer3_outputs(1925) <= not a;
    layer3_outputs(1926) <= not a or b;
    layer3_outputs(1927) <= a;
    layer3_outputs(1928) <= not a or b;
    layer3_outputs(1929) <= a;
    layer3_outputs(1930) <= not b or a;
    layer3_outputs(1931) <= not b;
    layer3_outputs(1932) <= not a;
    layer3_outputs(1933) <= a or b;
    layer3_outputs(1934) <= '0';
    layer3_outputs(1935) <= a and b;
    layer3_outputs(1936) <= a and not b;
    layer3_outputs(1937) <= a and not b;
    layer3_outputs(1938) <= not a;
    layer3_outputs(1939) <= not b;
    layer3_outputs(1940) <= a or b;
    layer3_outputs(1941) <= b and not a;
    layer3_outputs(1942) <= '0';
    layer3_outputs(1943) <= not (a or b);
    layer3_outputs(1944) <= not b;
    layer3_outputs(1945) <= not a or b;
    layer3_outputs(1946) <= b;
    layer3_outputs(1947) <= a or b;
    layer3_outputs(1948) <= '1';
    layer3_outputs(1949) <= b and not a;
    layer3_outputs(1950) <= b;
    layer3_outputs(1951) <= '1';
    layer3_outputs(1952) <= a xor b;
    layer3_outputs(1953) <= '0';
    layer3_outputs(1954) <= '1';
    layer3_outputs(1955) <= a or b;
    layer3_outputs(1956) <= not (a and b);
    layer3_outputs(1957) <= a or b;
    layer3_outputs(1958) <= a or b;
    layer3_outputs(1959) <= '0';
    layer3_outputs(1960) <= a;
    layer3_outputs(1961) <= a and b;
    layer3_outputs(1962) <= '1';
    layer3_outputs(1963) <= not b;
    layer3_outputs(1964) <= not a or b;
    layer3_outputs(1965) <= '1';
    layer3_outputs(1966) <= a xor b;
    layer3_outputs(1967) <= a and b;
    layer3_outputs(1968) <= not (a or b);
    layer3_outputs(1969) <= not (a xor b);
    layer3_outputs(1970) <= not (a or b);
    layer3_outputs(1971) <= a and not b;
    layer3_outputs(1972) <= a;
    layer3_outputs(1973) <= a and not b;
    layer3_outputs(1974) <= '1';
    layer3_outputs(1975) <= b and not a;
    layer3_outputs(1976) <= a or b;
    layer3_outputs(1977) <= a;
    layer3_outputs(1978) <= not (a xor b);
    layer3_outputs(1979) <= not (a and b);
    layer3_outputs(1980) <= b and not a;
    layer3_outputs(1981) <= '0';
    layer3_outputs(1982) <= not (a and b);
    layer3_outputs(1983) <= not b;
    layer3_outputs(1984) <= not b or a;
    layer3_outputs(1985) <= b and not a;
    layer3_outputs(1986) <= '0';
    layer3_outputs(1987) <= not (a or b);
    layer3_outputs(1988) <= not a or b;
    layer3_outputs(1989) <= a and b;
    layer3_outputs(1990) <= not a or b;
    layer3_outputs(1991) <= not b;
    layer3_outputs(1992) <= a;
    layer3_outputs(1993) <= a;
    layer3_outputs(1994) <= a;
    layer3_outputs(1995) <= '1';
    layer3_outputs(1996) <= a or b;
    layer3_outputs(1997) <= not a;
    layer3_outputs(1998) <= a or b;
    layer3_outputs(1999) <= not b;
    layer3_outputs(2000) <= not (a and b);
    layer3_outputs(2001) <= not (a xor b);
    layer3_outputs(2002) <= '1';
    layer3_outputs(2003) <= a or b;
    layer3_outputs(2004) <= '1';
    layer3_outputs(2005) <= a and b;
    layer3_outputs(2006) <= not b or a;
    layer3_outputs(2007) <= not (a xor b);
    layer3_outputs(2008) <= not a or b;
    layer3_outputs(2009) <= not (a and b);
    layer3_outputs(2010) <= not b;
    layer3_outputs(2011) <= a and not b;
    layer3_outputs(2012) <= not (a and b);
    layer3_outputs(2013) <= a or b;
    layer3_outputs(2014) <= '1';
    layer3_outputs(2015) <= not b or a;
    layer3_outputs(2016) <= not (a xor b);
    layer3_outputs(2017) <= not a;
    layer3_outputs(2018) <= a or b;
    layer3_outputs(2019) <= '0';
    layer3_outputs(2020) <= not (a and b);
    layer3_outputs(2021) <= a;
    layer3_outputs(2022) <= not b or a;
    layer3_outputs(2023) <= '0';
    layer3_outputs(2024) <= '1';
    layer3_outputs(2025) <= not (a and b);
    layer3_outputs(2026) <= b and not a;
    layer3_outputs(2027) <= a or b;
    layer3_outputs(2028) <= '0';
    layer3_outputs(2029) <= not (a and b);
    layer3_outputs(2030) <= not b or a;
    layer3_outputs(2031) <= '1';
    layer3_outputs(2032) <= a;
    layer3_outputs(2033) <= b;
    layer3_outputs(2034) <= a or b;
    layer3_outputs(2035) <= a and not b;
    layer3_outputs(2036) <= not (a or b);
    layer3_outputs(2037) <= '1';
    layer3_outputs(2038) <= not b;
    layer3_outputs(2039) <= not a;
    layer3_outputs(2040) <= '0';
    layer3_outputs(2041) <= a and not b;
    layer3_outputs(2042) <= not a or b;
    layer3_outputs(2043) <= not a or b;
    layer3_outputs(2044) <= not b;
    layer3_outputs(2045) <= not a;
    layer3_outputs(2046) <= a and b;
    layer3_outputs(2047) <= not a or b;
    layer3_outputs(2048) <= '0';
    layer3_outputs(2049) <= not b or a;
    layer3_outputs(2050) <= not b;
    layer3_outputs(2051) <= a or b;
    layer3_outputs(2052) <= not b or a;
    layer3_outputs(2053) <= a and b;
    layer3_outputs(2054) <= a or b;
    layer3_outputs(2055) <= not b;
    layer3_outputs(2056) <= b;
    layer3_outputs(2057) <= not (a and b);
    layer3_outputs(2058) <= not (a xor b);
    layer3_outputs(2059) <= a;
    layer3_outputs(2060) <= a;
    layer3_outputs(2061) <= not b;
    layer3_outputs(2062) <= a;
    layer3_outputs(2063) <= not b or a;
    layer3_outputs(2064) <= b;
    layer3_outputs(2065) <= '1';
    layer3_outputs(2066) <= '1';
    layer3_outputs(2067) <= b;
    layer3_outputs(2068) <= a and not b;
    layer3_outputs(2069) <= not (a or b);
    layer3_outputs(2070) <= a;
    layer3_outputs(2071) <= not (a and b);
    layer3_outputs(2072) <= '0';
    layer3_outputs(2073) <= not a or b;
    layer3_outputs(2074) <= a or b;
    layer3_outputs(2075) <= b;
    layer3_outputs(2076) <= not b or a;
    layer3_outputs(2077) <= a;
    layer3_outputs(2078) <= '0';
    layer3_outputs(2079) <= not b;
    layer3_outputs(2080) <= b;
    layer3_outputs(2081) <= not b;
    layer3_outputs(2082) <= '0';
    layer3_outputs(2083) <= not (a or b);
    layer3_outputs(2084) <= not a or b;
    layer3_outputs(2085) <= '0';
    layer3_outputs(2086) <= not a;
    layer3_outputs(2087) <= b;
    layer3_outputs(2088) <= b;
    layer3_outputs(2089) <= a or b;
    layer3_outputs(2090) <= a;
    layer3_outputs(2091) <= a or b;
    layer3_outputs(2092) <= a or b;
    layer3_outputs(2093) <= not a;
    layer3_outputs(2094) <= a xor b;
    layer3_outputs(2095) <= not b;
    layer3_outputs(2096) <= not b;
    layer3_outputs(2097) <= not (a or b);
    layer3_outputs(2098) <= not b;
    layer3_outputs(2099) <= not b or a;
    layer3_outputs(2100) <= b and not a;
    layer3_outputs(2101) <= not a;
    layer3_outputs(2102) <= a;
    layer3_outputs(2103) <= '0';
    layer3_outputs(2104) <= '1';
    layer3_outputs(2105) <= '0';
    layer3_outputs(2106) <= '0';
    layer3_outputs(2107) <= not a or b;
    layer3_outputs(2108) <= not b or a;
    layer3_outputs(2109) <= b and not a;
    layer3_outputs(2110) <= not a or b;
    layer3_outputs(2111) <= '1';
    layer3_outputs(2112) <= not (a or b);
    layer3_outputs(2113) <= not a;
    layer3_outputs(2114) <= '1';
    layer3_outputs(2115) <= '0';
    layer3_outputs(2116) <= a or b;
    layer3_outputs(2117) <= '0';
    layer3_outputs(2118) <= not b or a;
    layer3_outputs(2119) <= not b;
    layer3_outputs(2120) <= a and not b;
    layer3_outputs(2121) <= not (a and b);
    layer3_outputs(2122) <= '0';
    layer3_outputs(2123) <= '1';
    layer3_outputs(2124) <= not (a and b);
    layer3_outputs(2125) <= a;
    layer3_outputs(2126) <= b and not a;
    layer3_outputs(2127) <= a;
    layer3_outputs(2128) <= a and b;
    layer3_outputs(2129) <= not (a or b);
    layer3_outputs(2130) <= a and not b;
    layer3_outputs(2131) <= not (a and b);
    layer3_outputs(2132) <= not (a and b);
    layer3_outputs(2133) <= a;
    layer3_outputs(2134) <= not b;
    layer3_outputs(2135) <= a or b;
    layer3_outputs(2136) <= not (a or b);
    layer3_outputs(2137) <= b and not a;
    layer3_outputs(2138) <= b and not a;
    layer3_outputs(2139) <= not a;
    layer3_outputs(2140) <= a or b;
    layer3_outputs(2141) <= b and not a;
    layer3_outputs(2142) <= not b or a;
    layer3_outputs(2143) <= b;
    layer3_outputs(2144) <= a;
    layer3_outputs(2145) <= '1';
    layer3_outputs(2146) <= not a;
    layer3_outputs(2147) <= a;
    layer3_outputs(2148) <= not (a or b);
    layer3_outputs(2149) <= a and not b;
    layer3_outputs(2150) <= '1';
    layer3_outputs(2151) <= not a or b;
    layer3_outputs(2152) <= not a or b;
    layer3_outputs(2153) <= '1';
    layer3_outputs(2154) <= not a or b;
    layer3_outputs(2155) <= a;
    layer3_outputs(2156) <= a and b;
    layer3_outputs(2157) <= a and not b;
    layer3_outputs(2158) <= b;
    layer3_outputs(2159) <= not (a and b);
    layer3_outputs(2160) <= not (a and b);
    layer3_outputs(2161) <= b and not a;
    layer3_outputs(2162) <= not a or b;
    layer3_outputs(2163) <= b and not a;
    layer3_outputs(2164) <= '0';
    layer3_outputs(2165) <= '1';
    layer3_outputs(2166) <= a or b;
    layer3_outputs(2167) <= not a;
    layer3_outputs(2168) <= a or b;
    layer3_outputs(2169) <= a and b;
    layer3_outputs(2170) <= not b or a;
    layer3_outputs(2171) <= a xor b;
    layer3_outputs(2172) <= b and not a;
    layer3_outputs(2173) <= b;
    layer3_outputs(2174) <= a and not b;
    layer3_outputs(2175) <= b and not a;
    layer3_outputs(2176) <= '0';
    layer3_outputs(2177) <= a and not b;
    layer3_outputs(2178) <= not (a and b);
    layer3_outputs(2179) <= a or b;
    layer3_outputs(2180) <= a or b;
    layer3_outputs(2181) <= '1';
    layer3_outputs(2182) <= not (a and b);
    layer3_outputs(2183) <= b;
    layer3_outputs(2184) <= not (a and b);
    layer3_outputs(2185) <= a and not b;
    layer3_outputs(2186) <= '1';
    layer3_outputs(2187) <= a and b;
    layer3_outputs(2188) <= b;
    layer3_outputs(2189) <= not b or a;
    layer3_outputs(2190) <= not a;
    layer3_outputs(2191) <= '0';
    layer3_outputs(2192) <= a and not b;
    layer3_outputs(2193) <= not a;
    layer3_outputs(2194) <= a;
    layer3_outputs(2195) <= a and not b;
    layer3_outputs(2196) <= not a;
    layer3_outputs(2197) <= not a;
    layer3_outputs(2198) <= b and not a;
    layer3_outputs(2199) <= not b or a;
    layer3_outputs(2200) <= not b or a;
    layer3_outputs(2201) <= a and b;
    layer3_outputs(2202) <= not (a or b);
    layer3_outputs(2203) <= not b;
    layer3_outputs(2204) <= not a;
    layer3_outputs(2205) <= not (a xor b);
    layer3_outputs(2206) <= a and not b;
    layer3_outputs(2207) <= not b or a;
    layer3_outputs(2208) <= b and not a;
    layer3_outputs(2209) <= a or b;
    layer3_outputs(2210) <= not a;
    layer3_outputs(2211) <= a;
    layer3_outputs(2212) <= not b or a;
    layer3_outputs(2213) <= b;
    layer3_outputs(2214) <= a;
    layer3_outputs(2215) <= not b or a;
    layer3_outputs(2216) <= a and b;
    layer3_outputs(2217) <= not (a and b);
    layer3_outputs(2218) <= '0';
    layer3_outputs(2219) <= not b or a;
    layer3_outputs(2220) <= a or b;
    layer3_outputs(2221) <= a and b;
    layer3_outputs(2222) <= b;
    layer3_outputs(2223) <= not (a or b);
    layer3_outputs(2224) <= a and not b;
    layer3_outputs(2225) <= a or b;
    layer3_outputs(2226) <= a;
    layer3_outputs(2227) <= b;
    layer3_outputs(2228) <= not (a or b);
    layer3_outputs(2229) <= '1';
    layer3_outputs(2230) <= not (a and b);
    layer3_outputs(2231) <= not a or b;
    layer3_outputs(2232) <= not a or b;
    layer3_outputs(2233) <= '0';
    layer3_outputs(2234) <= not a;
    layer3_outputs(2235) <= b;
    layer3_outputs(2236) <= a and not b;
    layer3_outputs(2237) <= '0';
    layer3_outputs(2238) <= not b or a;
    layer3_outputs(2239) <= not b;
    layer3_outputs(2240) <= not a or b;
    layer3_outputs(2241) <= not (a and b);
    layer3_outputs(2242) <= b and not a;
    layer3_outputs(2243) <= a;
    layer3_outputs(2244) <= not a or b;
    layer3_outputs(2245) <= a;
    layer3_outputs(2246) <= b and not a;
    layer3_outputs(2247) <= b and not a;
    layer3_outputs(2248) <= a and b;
    layer3_outputs(2249) <= b;
    layer3_outputs(2250) <= b and not a;
    layer3_outputs(2251) <= not b;
    layer3_outputs(2252) <= b;
    layer3_outputs(2253) <= a;
    layer3_outputs(2254) <= '1';
    layer3_outputs(2255) <= a xor b;
    layer3_outputs(2256) <= not b;
    layer3_outputs(2257) <= not b;
    layer3_outputs(2258) <= not a or b;
    layer3_outputs(2259) <= '0';
    layer3_outputs(2260) <= a;
    layer3_outputs(2261) <= a and b;
    layer3_outputs(2262) <= not a;
    layer3_outputs(2263) <= a or b;
    layer3_outputs(2264) <= a;
    layer3_outputs(2265) <= '0';
    layer3_outputs(2266) <= not b or a;
    layer3_outputs(2267) <= not (a and b);
    layer3_outputs(2268) <= not a;
    layer3_outputs(2269) <= a or b;
    layer3_outputs(2270) <= '1';
    layer3_outputs(2271) <= not a;
    layer3_outputs(2272) <= b;
    layer3_outputs(2273) <= not (a and b);
    layer3_outputs(2274) <= not (a or b);
    layer3_outputs(2275) <= a;
    layer3_outputs(2276) <= not (a or b);
    layer3_outputs(2277) <= a and not b;
    layer3_outputs(2278) <= '1';
    layer3_outputs(2279) <= a and b;
    layer3_outputs(2280) <= not b;
    layer3_outputs(2281) <= a or b;
    layer3_outputs(2282) <= '1';
    layer3_outputs(2283) <= not a or b;
    layer3_outputs(2284) <= a or b;
    layer3_outputs(2285) <= not a or b;
    layer3_outputs(2286) <= not (a or b);
    layer3_outputs(2287) <= not a;
    layer3_outputs(2288) <= b;
    layer3_outputs(2289) <= not a or b;
    layer3_outputs(2290) <= a xor b;
    layer3_outputs(2291) <= '1';
    layer3_outputs(2292) <= a or b;
    layer3_outputs(2293) <= not a or b;
    layer3_outputs(2294) <= b and not a;
    layer3_outputs(2295) <= a;
    layer3_outputs(2296) <= b;
    layer3_outputs(2297) <= '1';
    layer3_outputs(2298) <= not (a xor b);
    layer3_outputs(2299) <= '1';
    layer3_outputs(2300) <= a or b;
    layer3_outputs(2301) <= a and not b;
    layer3_outputs(2302) <= not a;
    layer3_outputs(2303) <= '0';
    layer3_outputs(2304) <= b;
    layer3_outputs(2305) <= '0';
    layer3_outputs(2306) <= not b;
    layer3_outputs(2307) <= not a or b;
    layer3_outputs(2308) <= not (a or b);
    layer3_outputs(2309) <= not (a or b);
    layer3_outputs(2310) <= not b or a;
    layer3_outputs(2311) <= a and not b;
    layer3_outputs(2312) <= b;
    layer3_outputs(2313) <= '1';
    layer3_outputs(2314) <= not a;
    layer3_outputs(2315) <= b;
    layer3_outputs(2316) <= '1';
    layer3_outputs(2317) <= not a;
    layer3_outputs(2318) <= b and not a;
    layer3_outputs(2319) <= a;
    layer3_outputs(2320) <= not (a xor b);
    layer3_outputs(2321) <= '0';
    layer3_outputs(2322) <= not a or b;
    layer3_outputs(2323) <= '0';
    layer3_outputs(2324) <= not (a or b);
    layer3_outputs(2325) <= a and b;
    layer3_outputs(2326) <= not a;
    layer3_outputs(2327) <= a;
    layer3_outputs(2328) <= a and not b;
    layer3_outputs(2329) <= not a or b;
    layer3_outputs(2330) <= a or b;
    layer3_outputs(2331) <= a and b;
    layer3_outputs(2332) <= not a;
    layer3_outputs(2333) <= not (a and b);
    layer3_outputs(2334) <= not (a or b);
    layer3_outputs(2335) <= not b or a;
    layer3_outputs(2336) <= '0';
    layer3_outputs(2337) <= not (a or b);
    layer3_outputs(2338) <= not (a xor b);
    layer3_outputs(2339) <= not a;
    layer3_outputs(2340) <= not (a or b);
    layer3_outputs(2341) <= not b or a;
    layer3_outputs(2342) <= not (a or b);
    layer3_outputs(2343) <= '1';
    layer3_outputs(2344) <= a and not b;
    layer3_outputs(2345) <= a and not b;
    layer3_outputs(2346) <= b;
    layer3_outputs(2347) <= '1';
    layer3_outputs(2348) <= a;
    layer3_outputs(2349) <= not b;
    layer3_outputs(2350) <= b and not a;
    layer3_outputs(2351) <= a;
    layer3_outputs(2352) <= '1';
    layer3_outputs(2353) <= b and not a;
    layer3_outputs(2354) <= not a;
    layer3_outputs(2355) <= a and not b;
    layer3_outputs(2356) <= a and b;
    layer3_outputs(2357) <= a and b;
    layer3_outputs(2358) <= not b or a;
    layer3_outputs(2359) <= a and not b;
    layer3_outputs(2360) <= '0';
    layer3_outputs(2361) <= a and not b;
    layer3_outputs(2362) <= not (a or b);
    layer3_outputs(2363) <= a and b;
    layer3_outputs(2364) <= b and not a;
    layer3_outputs(2365) <= not (a or b);
    layer3_outputs(2366) <= '0';
    layer3_outputs(2367) <= a and b;
    layer3_outputs(2368) <= '1';
    layer3_outputs(2369) <= '0';
    layer3_outputs(2370) <= not b;
    layer3_outputs(2371) <= a and not b;
    layer3_outputs(2372) <= not b or a;
    layer3_outputs(2373) <= not b or a;
    layer3_outputs(2374) <= not b or a;
    layer3_outputs(2375) <= b and not a;
    layer3_outputs(2376) <= b and not a;
    layer3_outputs(2377) <= not b or a;
    layer3_outputs(2378) <= b;
    layer3_outputs(2379) <= b;
    layer3_outputs(2380) <= a and not b;
    layer3_outputs(2381) <= not (a or b);
    layer3_outputs(2382) <= a or b;
    layer3_outputs(2383) <= not b;
    layer3_outputs(2384) <= '1';
    layer3_outputs(2385) <= not b;
    layer3_outputs(2386) <= '1';
    layer3_outputs(2387) <= a and b;
    layer3_outputs(2388) <= not a;
    layer3_outputs(2389) <= not a or b;
    layer3_outputs(2390) <= a and not b;
    layer3_outputs(2391) <= a and not b;
    layer3_outputs(2392) <= a and b;
    layer3_outputs(2393) <= a and b;
    layer3_outputs(2394) <= '1';
    layer3_outputs(2395) <= not b or a;
    layer3_outputs(2396) <= '0';
    layer3_outputs(2397) <= '0';
    layer3_outputs(2398) <= not (a or b);
    layer3_outputs(2399) <= not a;
    layer3_outputs(2400) <= not a;
    layer3_outputs(2401) <= b;
    layer3_outputs(2402) <= not (a or b);
    layer3_outputs(2403) <= '0';
    layer3_outputs(2404) <= a and b;
    layer3_outputs(2405) <= a and not b;
    layer3_outputs(2406) <= not b or a;
    layer3_outputs(2407) <= '0';
    layer3_outputs(2408) <= not b;
    layer3_outputs(2409) <= not a or b;
    layer3_outputs(2410) <= b;
    layer3_outputs(2411) <= '1';
    layer3_outputs(2412) <= not (a or b);
    layer3_outputs(2413) <= not (a and b);
    layer3_outputs(2414) <= a or b;
    layer3_outputs(2415) <= not b;
    layer3_outputs(2416) <= not (a and b);
    layer3_outputs(2417) <= not a;
    layer3_outputs(2418) <= a and not b;
    layer3_outputs(2419) <= '0';
    layer3_outputs(2420) <= not a or b;
    layer3_outputs(2421) <= not (a or b);
    layer3_outputs(2422) <= a and not b;
    layer3_outputs(2423) <= a or b;
    layer3_outputs(2424) <= b;
    layer3_outputs(2425) <= not (a and b);
    layer3_outputs(2426) <= '0';
    layer3_outputs(2427) <= not a or b;
    layer3_outputs(2428) <= '1';
    layer3_outputs(2429) <= a or b;
    layer3_outputs(2430) <= b;
    layer3_outputs(2431) <= a or b;
    layer3_outputs(2432) <= not a or b;
    layer3_outputs(2433) <= not a;
    layer3_outputs(2434) <= b;
    layer3_outputs(2435) <= b and not a;
    layer3_outputs(2436) <= not a;
    layer3_outputs(2437) <= a and b;
    layer3_outputs(2438) <= a and b;
    layer3_outputs(2439) <= '1';
    layer3_outputs(2440) <= not a;
    layer3_outputs(2441) <= b and not a;
    layer3_outputs(2442) <= not (a and b);
    layer3_outputs(2443) <= a or b;
    layer3_outputs(2444) <= not (a xor b);
    layer3_outputs(2445) <= b;
    layer3_outputs(2446) <= not (a and b);
    layer3_outputs(2447) <= b;
    layer3_outputs(2448) <= not a or b;
    layer3_outputs(2449) <= a and not b;
    layer3_outputs(2450) <= b;
    layer3_outputs(2451) <= not (a and b);
    layer3_outputs(2452) <= a and not b;
    layer3_outputs(2453) <= not (a or b);
    layer3_outputs(2454) <= a and not b;
    layer3_outputs(2455) <= not (a or b);
    layer3_outputs(2456) <= b and not a;
    layer3_outputs(2457) <= not (a or b);
    layer3_outputs(2458) <= not (a or b);
    layer3_outputs(2459) <= not a;
    layer3_outputs(2460) <= not (a or b);
    layer3_outputs(2461) <= '1';
    layer3_outputs(2462) <= b and not a;
    layer3_outputs(2463) <= not a or b;
    layer3_outputs(2464) <= not (a and b);
    layer3_outputs(2465) <= a or b;
    layer3_outputs(2466) <= not a;
    layer3_outputs(2467) <= not a or b;
    layer3_outputs(2468) <= not (a or b);
    layer3_outputs(2469) <= not a or b;
    layer3_outputs(2470) <= '1';
    layer3_outputs(2471) <= not (a xor b);
    layer3_outputs(2472) <= not b or a;
    layer3_outputs(2473) <= not (a or b);
    layer3_outputs(2474) <= not (a and b);
    layer3_outputs(2475) <= not (a or b);
    layer3_outputs(2476) <= not a;
    layer3_outputs(2477) <= not b;
    layer3_outputs(2478) <= a or b;
    layer3_outputs(2479) <= a;
    layer3_outputs(2480) <= a or b;
    layer3_outputs(2481) <= not (a and b);
    layer3_outputs(2482) <= '0';
    layer3_outputs(2483) <= a;
    layer3_outputs(2484) <= not a or b;
    layer3_outputs(2485) <= a or b;
    layer3_outputs(2486) <= a and b;
    layer3_outputs(2487) <= a and not b;
    layer3_outputs(2488) <= not (a and b);
    layer3_outputs(2489) <= not (a or b);
    layer3_outputs(2490) <= b and not a;
    layer3_outputs(2491) <= not (a or b);
    layer3_outputs(2492) <= '1';
    layer3_outputs(2493) <= b;
    layer3_outputs(2494) <= not b or a;
    layer3_outputs(2495) <= b and not a;
    layer3_outputs(2496) <= b;
    layer3_outputs(2497) <= a and b;
    layer3_outputs(2498) <= not a;
    layer3_outputs(2499) <= a;
    layer3_outputs(2500) <= '0';
    layer3_outputs(2501) <= not b;
    layer3_outputs(2502) <= not (a or b);
    layer3_outputs(2503) <= a;
    layer3_outputs(2504) <= not b;
    layer3_outputs(2505) <= '1';
    layer3_outputs(2506) <= not a;
    layer3_outputs(2507) <= not b or a;
    layer3_outputs(2508) <= not b or a;
    layer3_outputs(2509) <= b and not a;
    layer3_outputs(2510) <= not b or a;
    layer3_outputs(2511) <= '0';
    layer3_outputs(2512) <= b;
    layer3_outputs(2513) <= a and not b;
    layer3_outputs(2514) <= not b;
    layer3_outputs(2515) <= not (a or b);
    layer3_outputs(2516) <= b;
    layer3_outputs(2517) <= a or b;
    layer3_outputs(2518) <= not a or b;
    layer3_outputs(2519) <= '1';
    layer3_outputs(2520) <= b;
    layer3_outputs(2521) <= not (a and b);
    layer3_outputs(2522) <= not a;
    layer3_outputs(2523) <= not (a and b);
    layer3_outputs(2524) <= a and b;
    layer3_outputs(2525) <= '1';
    layer3_outputs(2526) <= '0';
    layer3_outputs(2527) <= a or b;
    layer3_outputs(2528) <= '0';
    layer3_outputs(2529) <= not a or b;
    layer3_outputs(2530) <= a and not b;
    layer3_outputs(2531) <= not b or a;
    layer3_outputs(2532) <= a and not b;
    layer3_outputs(2533) <= '0';
    layer3_outputs(2534) <= not b or a;
    layer3_outputs(2535) <= '0';
    layer3_outputs(2536) <= not a or b;
    layer3_outputs(2537) <= '0';
    layer3_outputs(2538) <= not b or a;
    layer3_outputs(2539) <= '1';
    layer3_outputs(2540) <= not b or a;
    layer3_outputs(2541) <= a;
    layer3_outputs(2542) <= a and not b;
    layer3_outputs(2543) <= '1';
    layer3_outputs(2544) <= b and not a;
    layer3_outputs(2545) <= not (a and b);
    layer3_outputs(2546) <= not a or b;
    layer3_outputs(2547) <= '0';
    layer3_outputs(2548) <= a or b;
    layer3_outputs(2549) <= a or b;
    layer3_outputs(2550) <= not (a or b);
    layer3_outputs(2551) <= b;
    layer3_outputs(2552) <= a;
    layer3_outputs(2553) <= a or b;
    layer3_outputs(2554) <= not (a or b);
    layer3_outputs(2555) <= b;
    layer3_outputs(2556) <= a;
    layer3_outputs(2557) <= not (a or b);
    layer3_outputs(2558) <= not (a and b);
    layer3_outputs(2559) <= '0';
    layer3_outputs(2560) <= '1';
    layer3_outputs(2561) <= not a or b;
    layer3_outputs(2562) <= b;
    layer3_outputs(2563) <= b;
    layer3_outputs(2564) <= not (a and b);
    layer3_outputs(2565) <= not a or b;
    layer3_outputs(2566) <= not (a or b);
    layer3_outputs(2567) <= a and b;
    layer3_outputs(2568) <= '0';
    layer3_outputs(2569) <= not a or b;
    layer3_outputs(2570) <= a or b;
    layer3_outputs(2571) <= not a;
    layer3_outputs(2572) <= a or b;
    layer3_outputs(2573) <= a and not b;
    layer3_outputs(2574) <= not a or b;
    layer3_outputs(2575) <= not b;
    layer3_outputs(2576) <= '1';
    layer3_outputs(2577) <= not (a or b);
    layer3_outputs(2578) <= not b or a;
    layer3_outputs(2579) <= '0';
    layer3_outputs(2580) <= a;
    layer3_outputs(2581) <= a or b;
    layer3_outputs(2582) <= a and not b;
    layer3_outputs(2583) <= '0';
    layer3_outputs(2584) <= '1';
    layer3_outputs(2585) <= a;
    layer3_outputs(2586) <= not a;
    layer3_outputs(2587) <= a and not b;
    layer3_outputs(2588) <= a xor b;
    layer3_outputs(2589) <= '1';
    layer3_outputs(2590) <= not b or a;
    layer3_outputs(2591) <= not b;
    layer3_outputs(2592) <= b and not a;
    layer3_outputs(2593) <= not (a and b);
    layer3_outputs(2594) <= a and b;
    layer3_outputs(2595) <= not a or b;
    layer3_outputs(2596) <= '0';
    layer3_outputs(2597) <= b;
    layer3_outputs(2598) <= not (a or b);
    layer3_outputs(2599) <= not b;
    layer3_outputs(2600) <= not (a or b);
    layer3_outputs(2601) <= a and not b;
    layer3_outputs(2602) <= not (a xor b);
    layer3_outputs(2603) <= not a;
    layer3_outputs(2604) <= not a or b;
    layer3_outputs(2605) <= a and b;
    layer3_outputs(2606) <= not a;
    layer3_outputs(2607) <= b;
    layer3_outputs(2608) <= not (a or b);
    layer3_outputs(2609) <= '1';
    layer3_outputs(2610) <= not a;
    layer3_outputs(2611) <= not (a and b);
    layer3_outputs(2612) <= not b or a;
    layer3_outputs(2613) <= '0';
    layer3_outputs(2614) <= not (a or b);
    layer3_outputs(2615) <= not a;
    layer3_outputs(2616) <= not (a and b);
    layer3_outputs(2617) <= '1';
    layer3_outputs(2618) <= not (a and b);
    layer3_outputs(2619) <= a;
    layer3_outputs(2620) <= '0';
    layer3_outputs(2621) <= a;
    layer3_outputs(2622) <= b and not a;
    layer3_outputs(2623) <= not b;
    layer3_outputs(2624) <= b;
    layer3_outputs(2625) <= '1';
    layer3_outputs(2626) <= '0';
    layer3_outputs(2627) <= not b;
    layer3_outputs(2628) <= not b;
    layer3_outputs(2629) <= not (a and b);
    layer3_outputs(2630) <= a and b;
    layer3_outputs(2631) <= not b or a;
    layer3_outputs(2632) <= a and b;
    layer3_outputs(2633) <= not b;
    layer3_outputs(2634) <= '0';
    layer3_outputs(2635) <= a or b;
    layer3_outputs(2636) <= not (a or b);
    layer3_outputs(2637) <= a xor b;
    layer3_outputs(2638) <= not a;
    layer3_outputs(2639) <= b and not a;
    layer3_outputs(2640) <= a and not b;
    layer3_outputs(2641) <= not b;
    layer3_outputs(2642) <= a xor b;
    layer3_outputs(2643) <= '1';
    layer3_outputs(2644) <= b and not a;
    layer3_outputs(2645) <= '0';
    layer3_outputs(2646) <= a and not b;
    layer3_outputs(2647) <= not b or a;
    layer3_outputs(2648) <= a xor b;
    layer3_outputs(2649) <= not (a xor b);
    layer3_outputs(2650) <= not (a or b);
    layer3_outputs(2651) <= a or b;
    layer3_outputs(2652) <= a;
    layer3_outputs(2653) <= a and b;
    layer3_outputs(2654) <= a;
    layer3_outputs(2655) <= a or b;
    layer3_outputs(2656) <= not (a and b);
    layer3_outputs(2657) <= a xor b;
    layer3_outputs(2658) <= a and not b;
    layer3_outputs(2659) <= b and not a;
    layer3_outputs(2660) <= not a or b;
    layer3_outputs(2661) <= a and b;
    layer3_outputs(2662) <= a and b;
    layer3_outputs(2663) <= a and b;
    layer3_outputs(2664) <= not a;
    layer3_outputs(2665) <= b;
    layer3_outputs(2666) <= a and not b;
    layer3_outputs(2667) <= not (a and b);
    layer3_outputs(2668) <= not a or b;
    layer3_outputs(2669) <= '0';
    layer3_outputs(2670) <= a;
    layer3_outputs(2671) <= not (a and b);
    layer3_outputs(2672) <= a or b;
    layer3_outputs(2673) <= a or b;
    layer3_outputs(2674) <= a or b;
    layer3_outputs(2675) <= b and not a;
    layer3_outputs(2676) <= not (a and b);
    layer3_outputs(2677) <= a or b;
    layer3_outputs(2678) <= '1';
    layer3_outputs(2679) <= not b or a;
    layer3_outputs(2680) <= a and b;
    layer3_outputs(2681) <= not a or b;
    layer3_outputs(2682) <= a;
    layer3_outputs(2683) <= a and b;
    layer3_outputs(2684) <= b and not a;
    layer3_outputs(2685) <= '1';
    layer3_outputs(2686) <= not a or b;
    layer3_outputs(2687) <= a and b;
    layer3_outputs(2688) <= b and not a;
    layer3_outputs(2689) <= a or b;
    layer3_outputs(2690) <= a;
    layer3_outputs(2691) <= b and not a;
    layer3_outputs(2692) <= not a;
    layer3_outputs(2693) <= not a;
    layer3_outputs(2694) <= a and not b;
    layer3_outputs(2695) <= a and b;
    layer3_outputs(2696) <= '0';
    layer3_outputs(2697) <= not a;
    layer3_outputs(2698) <= a and not b;
    layer3_outputs(2699) <= a and not b;
    layer3_outputs(2700) <= a;
    layer3_outputs(2701) <= a and b;
    layer3_outputs(2702) <= a and not b;
    layer3_outputs(2703) <= b and not a;
    layer3_outputs(2704) <= a;
    layer3_outputs(2705) <= '1';
    layer3_outputs(2706) <= not (a and b);
    layer3_outputs(2707) <= a and not b;
    layer3_outputs(2708) <= '1';
    layer3_outputs(2709) <= '0';
    layer3_outputs(2710) <= not b or a;
    layer3_outputs(2711) <= not a;
    layer3_outputs(2712) <= a or b;
    layer3_outputs(2713) <= '1';
    layer3_outputs(2714) <= not b or a;
    layer3_outputs(2715) <= not (a or b);
    layer3_outputs(2716) <= not a;
    layer3_outputs(2717) <= a and b;
    layer3_outputs(2718) <= not b;
    layer3_outputs(2719) <= not a;
    layer3_outputs(2720) <= a;
    layer3_outputs(2721) <= b and not a;
    layer3_outputs(2722) <= not (a and b);
    layer3_outputs(2723) <= not (a or b);
    layer3_outputs(2724) <= a or b;
    layer3_outputs(2725) <= a or b;
    layer3_outputs(2726) <= b and not a;
    layer3_outputs(2727) <= not (a and b);
    layer3_outputs(2728) <= b and not a;
    layer3_outputs(2729) <= not b or a;
    layer3_outputs(2730) <= not a;
    layer3_outputs(2731) <= '1';
    layer3_outputs(2732) <= not a;
    layer3_outputs(2733) <= b;
    layer3_outputs(2734) <= b and not a;
    layer3_outputs(2735) <= a;
    layer3_outputs(2736) <= not (a or b);
    layer3_outputs(2737) <= a xor b;
    layer3_outputs(2738) <= not a;
    layer3_outputs(2739) <= not a or b;
    layer3_outputs(2740) <= not (a and b);
    layer3_outputs(2741) <= not (a or b);
    layer3_outputs(2742) <= a or b;
    layer3_outputs(2743) <= a or b;
    layer3_outputs(2744) <= not b or a;
    layer3_outputs(2745) <= not (a and b);
    layer3_outputs(2746) <= not b;
    layer3_outputs(2747) <= a;
    layer3_outputs(2748) <= not b or a;
    layer3_outputs(2749) <= b;
    layer3_outputs(2750) <= a and b;
    layer3_outputs(2751) <= not (a and b);
    layer3_outputs(2752) <= a;
    layer3_outputs(2753) <= not a or b;
    layer3_outputs(2754) <= not (a and b);
    layer3_outputs(2755) <= b;
    layer3_outputs(2756) <= a and not b;
    layer3_outputs(2757) <= '0';
    layer3_outputs(2758) <= b;
    layer3_outputs(2759) <= a and not b;
    layer3_outputs(2760) <= not (a or b);
    layer3_outputs(2761) <= b;
    layer3_outputs(2762) <= not b or a;
    layer3_outputs(2763) <= b;
    layer3_outputs(2764) <= not a;
    layer3_outputs(2765) <= not b or a;
    layer3_outputs(2766) <= not b;
    layer3_outputs(2767) <= '1';
    layer3_outputs(2768) <= not a or b;
    layer3_outputs(2769) <= not a;
    layer3_outputs(2770) <= not a or b;
    layer3_outputs(2771) <= a;
    layer3_outputs(2772) <= b and not a;
    layer3_outputs(2773) <= '1';
    layer3_outputs(2774) <= not b;
    layer3_outputs(2775) <= a;
    layer3_outputs(2776) <= '0';
    layer3_outputs(2777) <= '0';
    layer3_outputs(2778) <= '1';
    layer3_outputs(2779) <= not a;
    layer3_outputs(2780) <= a or b;
    layer3_outputs(2781) <= not b or a;
    layer3_outputs(2782) <= b;
    layer3_outputs(2783) <= a and b;
    layer3_outputs(2784) <= not (a or b);
    layer3_outputs(2785) <= a and b;
    layer3_outputs(2786) <= not a;
    layer3_outputs(2787) <= b;
    layer3_outputs(2788) <= not a;
    layer3_outputs(2789) <= '0';
    layer3_outputs(2790) <= a;
    layer3_outputs(2791) <= not (a or b);
    layer3_outputs(2792) <= not a;
    layer3_outputs(2793) <= b and not a;
    layer3_outputs(2794) <= a and not b;
    layer3_outputs(2795) <= a;
    layer3_outputs(2796) <= a and not b;
    layer3_outputs(2797) <= not (a or b);
    layer3_outputs(2798) <= a;
    layer3_outputs(2799) <= a and not b;
    layer3_outputs(2800) <= '0';
    layer3_outputs(2801) <= a and b;
    layer3_outputs(2802) <= a and b;
    layer3_outputs(2803) <= a or b;
    layer3_outputs(2804) <= not a or b;
    layer3_outputs(2805) <= '0';
    layer3_outputs(2806) <= a and not b;
    layer3_outputs(2807) <= not a;
    layer3_outputs(2808) <= not (a or b);
    layer3_outputs(2809) <= not b or a;
    layer3_outputs(2810) <= not (a and b);
    layer3_outputs(2811) <= a or b;
    layer3_outputs(2812) <= not (a xor b);
    layer3_outputs(2813) <= b and not a;
    layer3_outputs(2814) <= not (a xor b);
    layer3_outputs(2815) <= not b;
    layer3_outputs(2816) <= not (a or b);
    layer3_outputs(2817) <= not (a and b);
    layer3_outputs(2818) <= a and b;
    layer3_outputs(2819) <= not b;
    layer3_outputs(2820) <= a xor b;
    layer3_outputs(2821) <= not a;
    layer3_outputs(2822) <= a or b;
    layer3_outputs(2823) <= a and not b;
    layer3_outputs(2824) <= a xor b;
    layer3_outputs(2825) <= a or b;
    layer3_outputs(2826) <= a and b;
    layer3_outputs(2827) <= a and not b;
    layer3_outputs(2828) <= not a or b;
    layer3_outputs(2829) <= not (a and b);
    layer3_outputs(2830) <= '0';
    layer3_outputs(2831) <= not (a and b);
    layer3_outputs(2832) <= a or b;
    layer3_outputs(2833) <= '1';
    layer3_outputs(2834) <= b and not a;
    layer3_outputs(2835) <= a and b;
    layer3_outputs(2836) <= a;
    layer3_outputs(2837) <= a and not b;
    layer3_outputs(2838) <= not a or b;
    layer3_outputs(2839) <= b and not a;
    layer3_outputs(2840) <= a and b;
    layer3_outputs(2841) <= not b or a;
    layer3_outputs(2842) <= not b;
    layer3_outputs(2843) <= '0';
    layer3_outputs(2844) <= not a;
    layer3_outputs(2845) <= a or b;
    layer3_outputs(2846) <= '1';
    layer3_outputs(2847) <= not (a and b);
    layer3_outputs(2848) <= not (a and b);
    layer3_outputs(2849) <= a;
    layer3_outputs(2850) <= not a;
    layer3_outputs(2851) <= '0';
    layer3_outputs(2852) <= a and not b;
    layer3_outputs(2853) <= not a or b;
    layer3_outputs(2854) <= a or b;
    layer3_outputs(2855) <= '0';
    layer3_outputs(2856) <= not (a xor b);
    layer3_outputs(2857) <= not a or b;
    layer3_outputs(2858) <= not (a or b);
    layer3_outputs(2859) <= '0';
    layer3_outputs(2860) <= '0';
    layer3_outputs(2861) <= not (a or b);
    layer3_outputs(2862) <= not b;
    layer3_outputs(2863) <= '1';
    layer3_outputs(2864) <= b;
    layer3_outputs(2865) <= b;
    layer3_outputs(2866) <= not a;
    layer3_outputs(2867) <= a and not b;
    layer3_outputs(2868) <= '0';
    layer3_outputs(2869) <= a xor b;
    layer3_outputs(2870) <= not (a or b);
    layer3_outputs(2871) <= '1';
    layer3_outputs(2872) <= not b or a;
    layer3_outputs(2873) <= a and not b;
    layer3_outputs(2874) <= not a;
    layer3_outputs(2875) <= b;
    layer3_outputs(2876) <= a;
    layer3_outputs(2877) <= not b or a;
    layer3_outputs(2878) <= not a;
    layer3_outputs(2879) <= '1';
    layer3_outputs(2880) <= '0';
    layer3_outputs(2881) <= b and not a;
    layer3_outputs(2882) <= a or b;
    layer3_outputs(2883) <= '1';
    layer3_outputs(2884) <= '0';
    layer3_outputs(2885) <= b;
    layer3_outputs(2886) <= not a or b;
    layer3_outputs(2887) <= a and not b;
    layer3_outputs(2888) <= not a;
    layer3_outputs(2889) <= a and b;
    layer3_outputs(2890) <= not a or b;
    layer3_outputs(2891) <= a or b;
    layer3_outputs(2892) <= b;
    layer3_outputs(2893) <= a and not b;
    layer3_outputs(2894) <= a and not b;
    layer3_outputs(2895) <= not (a or b);
    layer3_outputs(2896) <= '0';
    layer3_outputs(2897) <= not (a and b);
    layer3_outputs(2898) <= a or b;
    layer3_outputs(2899) <= b;
    layer3_outputs(2900) <= not (a or b);
    layer3_outputs(2901) <= b;
    layer3_outputs(2902) <= a and not b;
    layer3_outputs(2903) <= not a;
    layer3_outputs(2904) <= not b;
    layer3_outputs(2905) <= a and b;
    layer3_outputs(2906) <= a and b;
    layer3_outputs(2907) <= not a;
    layer3_outputs(2908) <= '0';
    layer3_outputs(2909) <= a;
    layer3_outputs(2910) <= a;
    layer3_outputs(2911) <= not a or b;
    layer3_outputs(2912) <= not a;
    layer3_outputs(2913) <= a and b;
    layer3_outputs(2914) <= a;
    layer3_outputs(2915) <= '0';
    layer3_outputs(2916) <= not b;
    layer3_outputs(2917) <= a or b;
    layer3_outputs(2918) <= a;
    layer3_outputs(2919) <= b;
    layer3_outputs(2920) <= not a or b;
    layer3_outputs(2921) <= not a;
    layer3_outputs(2922) <= b;
    layer3_outputs(2923) <= not b;
    layer3_outputs(2924) <= a or b;
    layer3_outputs(2925) <= not b or a;
    layer3_outputs(2926) <= not b;
    layer3_outputs(2927) <= a;
    layer3_outputs(2928) <= not (a and b);
    layer3_outputs(2929) <= not b or a;
    layer3_outputs(2930) <= a and not b;
    layer3_outputs(2931) <= not (a and b);
    layer3_outputs(2932) <= a xor b;
    layer3_outputs(2933) <= not (a and b);
    layer3_outputs(2934) <= b;
    layer3_outputs(2935) <= not a or b;
    layer3_outputs(2936) <= a or b;
    layer3_outputs(2937) <= b and not a;
    layer3_outputs(2938) <= b and not a;
    layer3_outputs(2939) <= b and not a;
    layer3_outputs(2940) <= not b;
    layer3_outputs(2941) <= not a;
    layer3_outputs(2942) <= not (a and b);
    layer3_outputs(2943) <= not a or b;
    layer3_outputs(2944) <= not b or a;
    layer3_outputs(2945) <= not b or a;
    layer3_outputs(2946) <= b and not a;
    layer3_outputs(2947) <= not (a or b);
    layer3_outputs(2948) <= not a;
    layer3_outputs(2949) <= not b or a;
    layer3_outputs(2950) <= a and not b;
    layer3_outputs(2951) <= a or b;
    layer3_outputs(2952) <= '0';
    layer3_outputs(2953) <= b;
    layer3_outputs(2954) <= not b or a;
    layer3_outputs(2955) <= not (a xor b);
    layer3_outputs(2956) <= b;
    layer3_outputs(2957) <= not a;
    layer3_outputs(2958) <= b and not a;
    layer3_outputs(2959) <= a and b;
    layer3_outputs(2960) <= '1';
    layer3_outputs(2961) <= b and not a;
    layer3_outputs(2962) <= not a or b;
    layer3_outputs(2963) <= not (a or b);
    layer3_outputs(2964) <= b and not a;
    layer3_outputs(2965) <= b and not a;
    layer3_outputs(2966) <= not a;
    layer3_outputs(2967) <= not (a or b);
    layer3_outputs(2968) <= not a;
    layer3_outputs(2969) <= a;
    layer3_outputs(2970) <= not a or b;
    layer3_outputs(2971) <= b and not a;
    layer3_outputs(2972) <= not (a or b);
    layer3_outputs(2973) <= not a;
    layer3_outputs(2974) <= a and not b;
    layer3_outputs(2975) <= not b;
    layer3_outputs(2976) <= not (a or b);
    layer3_outputs(2977) <= not b;
    layer3_outputs(2978) <= '0';
    layer3_outputs(2979) <= not b or a;
    layer3_outputs(2980) <= not a;
    layer3_outputs(2981) <= a;
    layer3_outputs(2982) <= a and b;
    layer3_outputs(2983) <= a or b;
    layer3_outputs(2984) <= b;
    layer3_outputs(2985) <= '1';
    layer3_outputs(2986) <= not (a and b);
    layer3_outputs(2987) <= a;
    layer3_outputs(2988) <= not a or b;
    layer3_outputs(2989) <= '1';
    layer3_outputs(2990) <= not b;
    layer3_outputs(2991) <= '1';
    layer3_outputs(2992) <= b and not a;
    layer3_outputs(2993) <= a and b;
    layer3_outputs(2994) <= not (a and b);
    layer3_outputs(2995) <= '0';
    layer3_outputs(2996) <= a and b;
    layer3_outputs(2997) <= a and b;
    layer3_outputs(2998) <= a or b;
    layer3_outputs(2999) <= a;
    layer3_outputs(3000) <= b and not a;
    layer3_outputs(3001) <= not b;
    layer3_outputs(3002) <= not b or a;
    layer3_outputs(3003) <= '0';
    layer3_outputs(3004) <= a;
    layer3_outputs(3005) <= not b;
    layer3_outputs(3006) <= b;
    layer3_outputs(3007) <= '1';
    layer3_outputs(3008) <= not b or a;
    layer3_outputs(3009) <= b and not a;
    layer3_outputs(3010) <= a or b;
    layer3_outputs(3011) <= not (a xor b);
    layer3_outputs(3012) <= '1';
    layer3_outputs(3013) <= '1';
    layer3_outputs(3014) <= not b;
    layer3_outputs(3015) <= a xor b;
    layer3_outputs(3016) <= '1';
    layer3_outputs(3017) <= not (a and b);
    layer3_outputs(3018) <= '1';
    layer3_outputs(3019) <= not (a or b);
    layer3_outputs(3020) <= not (a and b);
    layer3_outputs(3021) <= b and not a;
    layer3_outputs(3022) <= a;
    layer3_outputs(3023) <= not a or b;
    layer3_outputs(3024) <= not b or a;
    layer3_outputs(3025) <= not a;
    layer3_outputs(3026) <= not b or a;
    layer3_outputs(3027) <= b and not a;
    layer3_outputs(3028) <= a and b;
    layer3_outputs(3029) <= not (a or b);
    layer3_outputs(3030) <= '1';
    layer3_outputs(3031) <= '0';
    layer3_outputs(3032) <= a or b;
    layer3_outputs(3033) <= a or b;
    layer3_outputs(3034) <= not b or a;
    layer3_outputs(3035) <= not b or a;
    layer3_outputs(3036) <= not b or a;
    layer3_outputs(3037) <= not (a and b);
    layer3_outputs(3038) <= a and b;
    layer3_outputs(3039) <= not a or b;
    layer3_outputs(3040) <= b and not a;
    layer3_outputs(3041) <= b;
    layer3_outputs(3042) <= not a or b;
    layer3_outputs(3043) <= not a or b;
    layer3_outputs(3044) <= a and b;
    layer3_outputs(3045) <= a or b;
    layer3_outputs(3046) <= not a;
    layer3_outputs(3047) <= not a;
    layer3_outputs(3048) <= not (a or b);
    layer3_outputs(3049) <= not b;
    layer3_outputs(3050) <= '0';
    layer3_outputs(3051) <= not (a or b);
    layer3_outputs(3052) <= not (a and b);
    layer3_outputs(3053) <= not (a or b);
    layer3_outputs(3054) <= '0';
    layer3_outputs(3055) <= a;
    layer3_outputs(3056) <= not b or a;
    layer3_outputs(3057) <= not b;
    layer3_outputs(3058) <= a and b;
    layer3_outputs(3059) <= '1';
    layer3_outputs(3060) <= a or b;
    layer3_outputs(3061) <= b and not a;
    layer3_outputs(3062) <= a;
    layer3_outputs(3063) <= not a or b;
    layer3_outputs(3064) <= b and not a;
    layer3_outputs(3065) <= not (a or b);
    layer3_outputs(3066) <= not a;
    layer3_outputs(3067) <= b and not a;
    layer3_outputs(3068) <= '0';
    layer3_outputs(3069) <= '0';
    layer3_outputs(3070) <= not b;
    layer3_outputs(3071) <= not b or a;
    layer3_outputs(3072) <= '1';
    layer3_outputs(3073) <= a xor b;
    layer3_outputs(3074) <= not a;
    layer3_outputs(3075) <= not a or b;
    layer3_outputs(3076) <= a or b;
    layer3_outputs(3077) <= '0';
    layer3_outputs(3078) <= b and not a;
    layer3_outputs(3079) <= b and not a;
    layer3_outputs(3080) <= not a;
    layer3_outputs(3081) <= b;
    layer3_outputs(3082) <= not (a xor b);
    layer3_outputs(3083) <= not (a xor b);
    layer3_outputs(3084) <= not a or b;
    layer3_outputs(3085) <= a and b;
    layer3_outputs(3086) <= a or b;
    layer3_outputs(3087) <= b and not a;
    layer3_outputs(3088) <= '1';
    layer3_outputs(3089) <= a and b;
    layer3_outputs(3090) <= not (a and b);
    layer3_outputs(3091) <= not b;
    layer3_outputs(3092) <= a and not b;
    layer3_outputs(3093) <= a or b;
    layer3_outputs(3094) <= b;
    layer3_outputs(3095) <= not a;
    layer3_outputs(3096) <= not a or b;
    layer3_outputs(3097) <= '0';
    layer3_outputs(3098) <= a and b;
    layer3_outputs(3099) <= not (a and b);
    layer3_outputs(3100) <= a and b;
    layer3_outputs(3101) <= not a or b;
    layer3_outputs(3102) <= not b;
    layer3_outputs(3103) <= b;
    layer3_outputs(3104) <= b and not a;
    layer3_outputs(3105) <= not (a or b);
    layer3_outputs(3106) <= not a;
    layer3_outputs(3107) <= not b;
    layer3_outputs(3108) <= not a or b;
    layer3_outputs(3109) <= not (a or b);
    layer3_outputs(3110) <= not b;
    layer3_outputs(3111) <= not a or b;
    layer3_outputs(3112) <= not (a and b);
    layer3_outputs(3113) <= '0';
    layer3_outputs(3114) <= not (a or b);
    layer3_outputs(3115) <= not b or a;
    layer3_outputs(3116) <= b and not a;
    layer3_outputs(3117) <= '0';
    layer3_outputs(3118) <= not a;
    layer3_outputs(3119) <= not b or a;
    layer3_outputs(3120) <= a and not b;
    layer3_outputs(3121) <= a and b;
    layer3_outputs(3122) <= a and not b;
    layer3_outputs(3123) <= a or b;
    layer3_outputs(3124) <= not b or a;
    layer3_outputs(3125) <= a;
    layer3_outputs(3126) <= '0';
    layer3_outputs(3127) <= a;
    layer3_outputs(3128) <= '0';
    layer3_outputs(3129) <= not (a and b);
    layer3_outputs(3130) <= not a or b;
    layer3_outputs(3131) <= '1';
    layer3_outputs(3132) <= a;
    layer3_outputs(3133) <= b;
    layer3_outputs(3134) <= not (a xor b);
    layer3_outputs(3135) <= a;
    layer3_outputs(3136) <= a and not b;
    layer3_outputs(3137) <= '0';
    layer3_outputs(3138) <= b and not a;
    layer3_outputs(3139) <= b;
    layer3_outputs(3140) <= not b;
    layer3_outputs(3141) <= b and not a;
    layer3_outputs(3142) <= '1';
    layer3_outputs(3143) <= not b;
    layer3_outputs(3144) <= not (a and b);
    layer3_outputs(3145) <= '0';
    layer3_outputs(3146) <= not b or a;
    layer3_outputs(3147) <= not b;
    layer3_outputs(3148) <= a or b;
    layer3_outputs(3149) <= a or b;
    layer3_outputs(3150) <= not b;
    layer3_outputs(3151) <= b;
    layer3_outputs(3152) <= '1';
    layer3_outputs(3153) <= not b;
    layer3_outputs(3154) <= '0';
    layer3_outputs(3155) <= not (a and b);
    layer3_outputs(3156) <= not (a and b);
    layer3_outputs(3157) <= '1';
    layer3_outputs(3158) <= b;
    layer3_outputs(3159) <= b;
    layer3_outputs(3160) <= not (a or b);
    layer3_outputs(3161) <= b;
    layer3_outputs(3162) <= not b or a;
    layer3_outputs(3163) <= not (a and b);
    layer3_outputs(3164) <= a xor b;
    layer3_outputs(3165) <= not b or a;
    layer3_outputs(3166) <= not a;
    layer3_outputs(3167) <= a and b;
    layer3_outputs(3168) <= not a or b;
    layer3_outputs(3169) <= not (a or b);
    layer3_outputs(3170) <= a and b;
    layer3_outputs(3171) <= not (a or b);
    layer3_outputs(3172) <= not b;
    layer3_outputs(3173) <= a or b;
    layer3_outputs(3174) <= not a or b;
    layer3_outputs(3175) <= not b;
    layer3_outputs(3176) <= not b or a;
    layer3_outputs(3177) <= a or b;
    layer3_outputs(3178) <= a;
    layer3_outputs(3179) <= not a;
    layer3_outputs(3180) <= a and not b;
    layer3_outputs(3181) <= b;
    layer3_outputs(3182) <= a and b;
    layer3_outputs(3183) <= a and b;
    layer3_outputs(3184) <= a and not b;
    layer3_outputs(3185) <= a and not b;
    layer3_outputs(3186) <= '1';
    layer3_outputs(3187) <= a and b;
    layer3_outputs(3188) <= not b;
    layer3_outputs(3189) <= not a or b;
    layer3_outputs(3190) <= b and not a;
    layer3_outputs(3191) <= '1';
    layer3_outputs(3192) <= a and b;
    layer3_outputs(3193) <= b and not a;
    layer3_outputs(3194) <= a and not b;
    layer3_outputs(3195) <= not b;
    layer3_outputs(3196) <= not b or a;
    layer3_outputs(3197) <= not a or b;
    layer3_outputs(3198) <= not a;
    layer3_outputs(3199) <= b and not a;
    layer3_outputs(3200) <= not a or b;
    layer3_outputs(3201) <= '0';
    layer3_outputs(3202) <= a xor b;
    layer3_outputs(3203) <= a and not b;
    layer3_outputs(3204) <= b and not a;
    layer3_outputs(3205) <= b and not a;
    layer3_outputs(3206) <= a or b;
    layer3_outputs(3207) <= b;
    layer3_outputs(3208) <= a and not b;
    layer3_outputs(3209) <= not (a and b);
    layer3_outputs(3210) <= not (a and b);
    layer3_outputs(3211) <= '1';
    layer3_outputs(3212) <= a xor b;
    layer3_outputs(3213) <= a and not b;
    layer3_outputs(3214) <= not b;
    layer3_outputs(3215) <= not (a and b);
    layer3_outputs(3216) <= a or b;
    layer3_outputs(3217) <= a and b;
    layer3_outputs(3218) <= a;
    layer3_outputs(3219) <= not b;
    layer3_outputs(3220) <= b and not a;
    layer3_outputs(3221) <= not (a and b);
    layer3_outputs(3222) <= not a or b;
    layer3_outputs(3223) <= '1';
    layer3_outputs(3224) <= '1';
    layer3_outputs(3225) <= a;
    layer3_outputs(3226) <= '0';
    layer3_outputs(3227) <= not (a or b);
    layer3_outputs(3228) <= not a or b;
    layer3_outputs(3229) <= not (a or b);
    layer3_outputs(3230) <= b and not a;
    layer3_outputs(3231) <= a or b;
    layer3_outputs(3232) <= not (a and b);
    layer3_outputs(3233) <= not a;
    layer3_outputs(3234) <= not b or a;
    layer3_outputs(3235) <= not (a or b);
    layer3_outputs(3236) <= a and not b;
    layer3_outputs(3237) <= a xor b;
    layer3_outputs(3238) <= a and b;
    layer3_outputs(3239) <= not b or a;
    layer3_outputs(3240) <= '0';
    layer3_outputs(3241) <= a xor b;
    layer3_outputs(3242) <= b;
    layer3_outputs(3243) <= not b or a;
    layer3_outputs(3244) <= not a;
    layer3_outputs(3245) <= '0';
    layer3_outputs(3246) <= a xor b;
    layer3_outputs(3247) <= not a or b;
    layer3_outputs(3248) <= b and not a;
    layer3_outputs(3249) <= not b or a;
    layer3_outputs(3250) <= a xor b;
    layer3_outputs(3251) <= not (a and b);
    layer3_outputs(3252) <= not (a and b);
    layer3_outputs(3253) <= b and not a;
    layer3_outputs(3254) <= b and not a;
    layer3_outputs(3255) <= a and b;
    layer3_outputs(3256) <= not (a and b);
    layer3_outputs(3257) <= not (a or b);
    layer3_outputs(3258) <= not b;
    layer3_outputs(3259) <= not b;
    layer3_outputs(3260) <= not (a xor b);
    layer3_outputs(3261) <= not a or b;
    layer3_outputs(3262) <= '0';
    layer3_outputs(3263) <= not a or b;
    layer3_outputs(3264) <= '1';
    layer3_outputs(3265) <= not (a or b);
    layer3_outputs(3266) <= b and not a;
    layer3_outputs(3267) <= '1';
    layer3_outputs(3268) <= not (a or b);
    layer3_outputs(3269) <= '1';
    layer3_outputs(3270) <= a;
    layer3_outputs(3271) <= not (a and b);
    layer3_outputs(3272) <= '1';
    layer3_outputs(3273) <= not (a and b);
    layer3_outputs(3274) <= '0';
    layer3_outputs(3275) <= not b or a;
    layer3_outputs(3276) <= not b;
    layer3_outputs(3277) <= '1';
    layer3_outputs(3278) <= not a or b;
    layer3_outputs(3279) <= a or b;
    layer3_outputs(3280) <= not a;
    layer3_outputs(3281) <= not (a and b);
    layer3_outputs(3282) <= not b;
    layer3_outputs(3283) <= a and not b;
    layer3_outputs(3284) <= b and not a;
    layer3_outputs(3285) <= not (a or b);
    layer3_outputs(3286) <= '1';
    layer3_outputs(3287) <= not b or a;
    layer3_outputs(3288) <= a xor b;
    layer3_outputs(3289) <= not (a and b);
    layer3_outputs(3290) <= a and not b;
    layer3_outputs(3291) <= not b or a;
    layer3_outputs(3292) <= '1';
    layer3_outputs(3293) <= not (a and b);
    layer3_outputs(3294) <= not (a and b);
    layer3_outputs(3295) <= a and not b;
    layer3_outputs(3296) <= not b;
    layer3_outputs(3297) <= not a;
    layer3_outputs(3298) <= '1';
    layer3_outputs(3299) <= b;
    layer3_outputs(3300) <= '1';
    layer3_outputs(3301) <= not b;
    layer3_outputs(3302) <= b and not a;
    layer3_outputs(3303) <= not a or b;
    layer3_outputs(3304) <= a;
    layer3_outputs(3305) <= a and b;
    layer3_outputs(3306) <= '1';
    layer3_outputs(3307) <= not b or a;
    layer3_outputs(3308) <= a and not b;
    layer3_outputs(3309) <= not (a or b);
    layer3_outputs(3310) <= not b or a;
    layer3_outputs(3311) <= b;
    layer3_outputs(3312) <= a and b;
    layer3_outputs(3313) <= '0';
    layer3_outputs(3314) <= b;
    layer3_outputs(3315) <= '1';
    layer3_outputs(3316) <= not a;
    layer3_outputs(3317) <= a or b;
    layer3_outputs(3318) <= '0';
    layer3_outputs(3319) <= a and not b;
    layer3_outputs(3320) <= b and not a;
    layer3_outputs(3321) <= not (a or b);
    layer3_outputs(3322) <= not b;
    layer3_outputs(3323) <= not (a or b);
    layer3_outputs(3324) <= not b;
    layer3_outputs(3325) <= a and not b;
    layer3_outputs(3326) <= b;
    layer3_outputs(3327) <= not b;
    layer3_outputs(3328) <= a;
    layer3_outputs(3329) <= not b;
    layer3_outputs(3330) <= not a;
    layer3_outputs(3331) <= a and b;
    layer3_outputs(3332) <= not a;
    layer3_outputs(3333) <= '0';
    layer3_outputs(3334) <= not (a or b);
    layer3_outputs(3335) <= '0';
    layer3_outputs(3336) <= a and not b;
    layer3_outputs(3337) <= not (a or b);
    layer3_outputs(3338) <= a and b;
    layer3_outputs(3339) <= a and b;
    layer3_outputs(3340) <= a or b;
    layer3_outputs(3341) <= not (a and b);
    layer3_outputs(3342) <= not a;
    layer3_outputs(3343) <= b;
    layer3_outputs(3344) <= b;
    layer3_outputs(3345) <= a and b;
    layer3_outputs(3346) <= not (a or b);
    layer3_outputs(3347) <= '0';
    layer3_outputs(3348) <= '0';
    layer3_outputs(3349) <= not b;
    layer3_outputs(3350) <= a and not b;
    layer3_outputs(3351) <= '0';
    layer3_outputs(3352) <= a and b;
    layer3_outputs(3353) <= not a or b;
    layer3_outputs(3354) <= not a;
    layer3_outputs(3355) <= a and not b;
    layer3_outputs(3356) <= not b or a;
    layer3_outputs(3357) <= not b or a;
    layer3_outputs(3358) <= b and not a;
    layer3_outputs(3359) <= '0';
    layer3_outputs(3360) <= not a;
    layer3_outputs(3361) <= not (a or b);
    layer3_outputs(3362) <= not b;
    layer3_outputs(3363) <= a;
    layer3_outputs(3364) <= '0';
    layer3_outputs(3365) <= a or b;
    layer3_outputs(3366) <= a;
    layer3_outputs(3367) <= a xor b;
    layer3_outputs(3368) <= a;
    layer3_outputs(3369) <= a and b;
    layer3_outputs(3370) <= '0';
    layer3_outputs(3371) <= a;
    layer3_outputs(3372) <= a and b;
    layer3_outputs(3373) <= not (a or b);
    layer3_outputs(3374) <= not b;
    layer3_outputs(3375) <= a or b;
    layer3_outputs(3376) <= b;
    layer3_outputs(3377) <= a or b;
    layer3_outputs(3378) <= not a or b;
    layer3_outputs(3379) <= '1';
    layer3_outputs(3380) <= a and b;
    layer3_outputs(3381) <= a and not b;
    layer3_outputs(3382) <= not a;
    layer3_outputs(3383) <= '1';
    layer3_outputs(3384) <= not (a or b);
    layer3_outputs(3385) <= a;
    layer3_outputs(3386) <= a and b;
    layer3_outputs(3387) <= a or b;
    layer3_outputs(3388) <= '1';
    layer3_outputs(3389) <= a and b;
    layer3_outputs(3390) <= '0';
    layer3_outputs(3391) <= b;
    layer3_outputs(3392) <= '0';
    layer3_outputs(3393) <= b;
    layer3_outputs(3394) <= not (a or b);
    layer3_outputs(3395) <= not (a or b);
    layer3_outputs(3396) <= not a or b;
    layer3_outputs(3397) <= a and b;
    layer3_outputs(3398) <= not a or b;
    layer3_outputs(3399) <= not b or a;
    layer3_outputs(3400) <= not a or b;
    layer3_outputs(3401) <= a;
    layer3_outputs(3402) <= not a or b;
    layer3_outputs(3403) <= a or b;
    layer3_outputs(3404) <= a;
    layer3_outputs(3405) <= not b;
    layer3_outputs(3406) <= a or b;
    layer3_outputs(3407) <= a or b;
    layer3_outputs(3408) <= not b or a;
    layer3_outputs(3409) <= b and not a;
    layer3_outputs(3410) <= not b;
    layer3_outputs(3411) <= not (a or b);
    layer3_outputs(3412) <= not a;
    layer3_outputs(3413) <= a and not b;
    layer3_outputs(3414) <= not b;
    layer3_outputs(3415) <= not (a and b);
    layer3_outputs(3416) <= a;
    layer3_outputs(3417) <= not b or a;
    layer3_outputs(3418) <= not b or a;
    layer3_outputs(3419) <= not a or b;
    layer3_outputs(3420) <= not b or a;
    layer3_outputs(3421) <= '0';
    layer3_outputs(3422) <= not a or b;
    layer3_outputs(3423) <= not (a or b);
    layer3_outputs(3424) <= '1';
    layer3_outputs(3425) <= not b;
    layer3_outputs(3426) <= not (a or b);
    layer3_outputs(3427) <= b;
    layer3_outputs(3428) <= b and not a;
    layer3_outputs(3429) <= b and not a;
    layer3_outputs(3430) <= a xor b;
    layer3_outputs(3431) <= a;
    layer3_outputs(3432) <= a;
    layer3_outputs(3433) <= a and not b;
    layer3_outputs(3434) <= '0';
    layer3_outputs(3435) <= not b or a;
    layer3_outputs(3436) <= not (a or b);
    layer3_outputs(3437) <= b and not a;
    layer3_outputs(3438) <= '1';
    layer3_outputs(3439) <= not b or a;
    layer3_outputs(3440) <= a and b;
    layer3_outputs(3441) <= a and b;
    layer3_outputs(3442) <= '1';
    layer3_outputs(3443) <= not a or b;
    layer3_outputs(3444) <= not b or a;
    layer3_outputs(3445) <= not (a or b);
    layer3_outputs(3446) <= a and b;
    layer3_outputs(3447) <= not a;
    layer3_outputs(3448) <= a and b;
    layer3_outputs(3449) <= b;
    layer3_outputs(3450) <= a or b;
    layer3_outputs(3451) <= a and b;
    layer3_outputs(3452) <= a;
    layer3_outputs(3453) <= not a;
    layer3_outputs(3454) <= not b or a;
    layer3_outputs(3455) <= not (a and b);
    layer3_outputs(3456) <= not a or b;
    layer3_outputs(3457) <= '0';
    layer3_outputs(3458) <= not (a and b);
    layer3_outputs(3459) <= b;
    layer3_outputs(3460) <= not a or b;
    layer3_outputs(3461) <= not (a and b);
    layer3_outputs(3462) <= b and not a;
    layer3_outputs(3463) <= not a;
    layer3_outputs(3464) <= b and not a;
    layer3_outputs(3465) <= a and not b;
    layer3_outputs(3466) <= not a or b;
    layer3_outputs(3467) <= a;
    layer3_outputs(3468) <= not (a or b);
    layer3_outputs(3469) <= not b or a;
    layer3_outputs(3470) <= a and not b;
    layer3_outputs(3471) <= '0';
    layer3_outputs(3472) <= not b or a;
    layer3_outputs(3473) <= '1';
    layer3_outputs(3474) <= a or b;
    layer3_outputs(3475) <= a or b;
    layer3_outputs(3476) <= a;
    layer3_outputs(3477) <= not b or a;
    layer3_outputs(3478) <= a and b;
    layer3_outputs(3479) <= not a or b;
    layer3_outputs(3480) <= b and not a;
    layer3_outputs(3481) <= not a or b;
    layer3_outputs(3482) <= b;
    layer3_outputs(3483) <= not b or a;
    layer3_outputs(3484) <= not b or a;
    layer3_outputs(3485) <= b;
    layer3_outputs(3486) <= a or b;
    layer3_outputs(3487) <= a;
    layer3_outputs(3488) <= a and b;
    layer3_outputs(3489) <= not b;
    layer3_outputs(3490) <= b;
    layer3_outputs(3491) <= not a;
    layer3_outputs(3492) <= b;
    layer3_outputs(3493) <= b and not a;
    layer3_outputs(3494) <= b and not a;
    layer3_outputs(3495) <= a and b;
    layer3_outputs(3496) <= a and not b;
    layer3_outputs(3497) <= not a or b;
    layer3_outputs(3498) <= not b;
    layer3_outputs(3499) <= not (a or b);
    layer3_outputs(3500) <= not b or a;
    layer3_outputs(3501) <= not (a or b);
    layer3_outputs(3502) <= a or b;
    layer3_outputs(3503) <= not (a or b);
    layer3_outputs(3504) <= not a or b;
    layer3_outputs(3505) <= not b;
    layer3_outputs(3506) <= not b or a;
    layer3_outputs(3507) <= b;
    layer3_outputs(3508) <= not (a and b);
    layer3_outputs(3509) <= a;
    layer3_outputs(3510) <= '1';
    layer3_outputs(3511) <= a xor b;
    layer3_outputs(3512) <= a and not b;
    layer3_outputs(3513) <= not (a or b);
    layer3_outputs(3514) <= a;
    layer3_outputs(3515) <= not b or a;
    layer3_outputs(3516) <= a and b;
    layer3_outputs(3517) <= not b;
    layer3_outputs(3518) <= not b;
    layer3_outputs(3519) <= a and b;
    layer3_outputs(3520) <= '0';
    layer3_outputs(3521) <= b and not a;
    layer3_outputs(3522) <= '1';
    layer3_outputs(3523) <= '1';
    layer3_outputs(3524) <= not (a or b);
    layer3_outputs(3525) <= a;
    layer3_outputs(3526) <= not (a or b);
    layer3_outputs(3527) <= not a or b;
    layer3_outputs(3528) <= not (a and b);
    layer3_outputs(3529) <= a or b;
    layer3_outputs(3530) <= b and not a;
    layer3_outputs(3531) <= '0';
    layer3_outputs(3532) <= not (a or b);
    layer3_outputs(3533) <= a or b;
    layer3_outputs(3534) <= not (a or b);
    layer3_outputs(3535) <= not a;
    layer3_outputs(3536) <= a and not b;
    layer3_outputs(3537) <= not b;
    layer3_outputs(3538) <= not (a and b);
    layer3_outputs(3539) <= '0';
    layer3_outputs(3540) <= '1';
    layer3_outputs(3541) <= not (a or b);
    layer3_outputs(3542) <= a or b;
    layer3_outputs(3543) <= b and not a;
    layer3_outputs(3544) <= b and not a;
    layer3_outputs(3545) <= '1';
    layer3_outputs(3546) <= '0';
    layer3_outputs(3547) <= b;
    layer3_outputs(3548) <= a and not b;
    layer3_outputs(3549) <= a xor b;
    layer3_outputs(3550) <= a or b;
    layer3_outputs(3551) <= '1';
    layer3_outputs(3552) <= a;
    layer3_outputs(3553) <= b;
    layer3_outputs(3554) <= a and b;
    layer3_outputs(3555) <= not (a and b);
    layer3_outputs(3556) <= not b;
    layer3_outputs(3557) <= not a;
    layer3_outputs(3558) <= a or b;
    layer3_outputs(3559) <= b and not a;
    layer3_outputs(3560) <= a or b;
    layer3_outputs(3561) <= a or b;
    layer3_outputs(3562) <= not (a or b);
    layer3_outputs(3563) <= '0';
    layer3_outputs(3564) <= not a or b;
    layer3_outputs(3565) <= a;
    layer3_outputs(3566) <= a and b;
    layer3_outputs(3567) <= '0';
    layer3_outputs(3568) <= a or b;
    layer3_outputs(3569) <= a or b;
    layer3_outputs(3570) <= a and not b;
    layer3_outputs(3571) <= b;
    layer3_outputs(3572) <= b and not a;
    layer3_outputs(3573) <= not (a or b);
    layer3_outputs(3574) <= a;
    layer3_outputs(3575) <= '1';
    layer3_outputs(3576) <= a or b;
    layer3_outputs(3577) <= '0';
    layer3_outputs(3578) <= b;
    layer3_outputs(3579) <= not a or b;
    layer3_outputs(3580) <= b and not a;
    layer3_outputs(3581) <= not (a or b);
    layer3_outputs(3582) <= not a;
    layer3_outputs(3583) <= b;
    layer3_outputs(3584) <= a and b;
    layer3_outputs(3585) <= a and not b;
    layer3_outputs(3586) <= a or b;
    layer3_outputs(3587) <= not a;
    layer3_outputs(3588) <= not (a and b);
    layer3_outputs(3589) <= '0';
    layer3_outputs(3590) <= '1';
    layer3_outputs(3591) <= not b or a;
    layer3_outputs(3592) <= '1';
    layer3_outputs(3593) <= b and not a;
    layer3_outputs(3594) <= not (a and b);
    layer3_outputs(3595) <= not a;
    layer3_outputs(3596) <= b and not a;
    layer3_outputs(3597) <= a and not b;
    layer3_outputs(3598) <= not b or a;
    layer3_outputs(3599) <= b and not a;
    layer3_outputs(3600) <= not b;
    layer3_outputs(3601) <= not a or b;
    layer3_outputs(3602) <= '1';
    layer3_outputs(3603) <= '0';
    layer3_outputs(3604) <= not a or b;
    layer3_outputs(3605) <= a and not b;
    layer3_outputs(3606) <= not (a or b);
    layer3_outputs(3607) <= b;
    layer3_outputs(3608) <= not (a or b);
    layer3_outputs(3609) <= '1';
    layer3_outputs(3610) <= a or b;
    layer3_outputs(3611) <= not (a and b);
    layer3_outputs(3612) <= not (a and b);
    layer3_outputs(3613) <= '1';
    layer3_outputs(3614) <= a and not b;
    layer3_outputs(3615) <= a and b;
    layer3_outputs(3616) <= b and not a;
    layer3_outputs(3617) <= '0';
    layer3_outputs(3618) <= not (a or b);
    layer3_outputs(3619) <= b;
    layer3_outputs(3620) <= a;
    layer3_outputs(3621) <= '0';
    layer3_outputs(3622) <= a or b;
    layer3_outputs(3623) <= not a or b;
    layer3_outputs(3624) <= a;
    layer3_outputs(3625) <= '0';
    layer3_outputs(3626) <= a and b;
    layer3_outputs(3627) <= not (a or b);
    layer3_outputs(3628) <= '0';
    layer3_outputs(3629) <= a and b;
    layer3_outputs(3630) <= not (a xor b);
    layer3_outputs(3631) <= a xor b;
    layer3_outputs(3632) <= b;
    layer3_outputs(3633) <= a or b;
    layer3_outputs(3634) <= not b or a;
    layer3_outputs(3635) <= a and b;
    layer3_outputs(3636) <= not b;
    layer3_outputs(3637) <= '1';
    layer3_outputs(3638) <= a or b;
    layer3_outputs(3639) <= not (a xor b);
    layer3_outputs(3640) <= a;
    layer3_outputs(3641) <= a and not b;
    layer3_outputs(3642) <= not (a or b);
    layer3_outputs(3643) <= b;
    layer3_outputs(3644) <= not (a and b);
    layer3_outputs(3645) <= '1';
    layer3_outputs(3646) <= a;
    layer3_outputs(3647) <= '1';
    layer3_outputs(3648) <= a;
    layer3_outputs(3649) <= not (a and b);
    layer3_outputs(3650) <= '0';
    layer3_outputs(3651) <= '0';
    layer3_outputs(3652) <= a;
    layer3_outputs(3653) <= a or b;
    layer3_outputs(3654) <= not b or a;
    layer3_outputs(3655) <= b;
    layer3_outputs(3656) <= '0';
    layer3_outputs(3657) <= '0';
    layer3_outputs(3658) <= b;
    layer3_outputs(3659) <= '1';
    layer3_outputs(3660) <= a and b;
    layer3_outputs(3661) <= b and not a;
    layer3_outputs(3662) <= a and b;
    layer3_outputs(3663) <= not (a or b);
    layer3_outputs(3664) <= a xor b;
    layer3_outputs(3665) <= not (a xor b);
    layer3_outputs(3666) <= not b or a;
    layer3_outputs(3667) <= a or b;
    layer3_outputs(3668) <= a;
    layer3_outputs(3669) <= not a;
    layer3_outputs(3670) <= a or b;
    layer3_outputs(3671) <= a and not b;
    layer3_outputs(3672) <= not a;
    layer3_outputs(3673) <= not b;
    layer3_outputs(3674) <= not (a and b);
    layer3_outputs(3675) <= a and b;
    layer3_outputs(3676) <= not a;
    layer3_outputs(3677) <= not a or b;
    layer3_outputs(3678) <= not b or a;
    layer3_outputs(3679) <= a and not b;
    layer3_outputs(3680) <= not b;
    layer3_outputs(3681) <= not a or b;
    layer3_outputs(3682) <= '1';
    layer3_outputs(3683) <= not (a or b);
    layer3_outputs(3684) <= not a or b;
    layer3_outputs(3685) <= '0';
    layer3_outputs(3686) <= not a;
    layer3_outputs(3687) <= '0';
    layer3_outputs(3688) <= not b;
    layer3_outputs(3689) <= a;
    layer3_outputs(3690) <= b;
    layer3_outputs(3691) <= '1';
    layer3_outputs(3692) <= b;
    layer3_outputs(3693) <= '1';
    layer3_outputs(3694) <= a and b;
    layer3_outputs(3695) <= a or b;
    layer3_outputs(3696) <= not b;
    layer3_outputs(3697) <= not b;
    layer3_outputs(3698) <= a and not b;
    layer3_outputs(3699) <= '1';
    layer3_outputs(3700) <= a;
    layer3_outputs(3701) <= '0';
    layer3_outputs(3702) <= b;
    layer3_outputs(3703) <= '1';
    layer3_outputs(3704) <= '0';
    layer3_outputs(3705) <= b;
    layer3_outputs(3706) <= b and not a;
    layer3_outputs(3707) <= not a or b;
    layer3_outputs(3708) <= a;
    layer3_outputs(3709) <= a or b;
    layer3_outputs(3710) <= not a or b;
    layer3_outputs(3711) <= '0';
    layer3_outputs(3712) <= b and not a;
    layer3_outputs(3713) <= not b;
    layer3_outputs(3714) <= a xor b;
    layer3_outputs(3715) <= b and not a;
    layer3_outputs(3716) <= not (a and b);
    layer3_outputs(3717) <= not a or b;
    layer3_outputs(3718) <= a xor b;
    layer3_outputs(3719) <= b;
    layer3_outputs(3720) <= not a;
    layer3_outputs(3721) <= not b or a;
    layer3_outputs(3722) <= not (a or b);
    layer3_outputs(3723) <= a and not b;
    layer3_outputs(3724) <= '0';
    layer3_outputs(3725) <= '1';
    layer3_outputs(3726) <= b and not a;
    layer3_outputs(3727) <= not b or a;
    layer3_outputs(3728) <= not b or a;
    layer3_outputs(3729) <= not a;
    layer3_outputs(3730) <= a;
    layer3_outputs(3731) <= '0';
    layer3_outputs(3732) <= '0';
    layer3_outputs(3733) <= not (a xor b);
    layer3_outputs(3734) <= '0';
    layer3_outputs(3735) <= b and not a;
    layer3_outputs(3736) <= a;
    layer3_outputs(3737) <= a and not b;
    layer3_outputs(3738) <= not (a or b);
    layer3_outputs(3739) <= not b or a;
    layer3_outputs(3740) <= b and not a;
    layer3_outputs(3741) <= b;
    layer3_outputs(3742) <= not (a and b);
    layer3_outputs(3743) <= a and not b;
    layer3_outputs(3744) <= not b or a;
    layer3_outputs(3745) <= a or b;
    layer3_outputs(3746) <= not (a or b);
    layer3_outputs(3747) <= not (a or b);
    layer3_outputs(3748) <= b and not a;
    layer3_outputs(3749) <= a or b;
    layer3_outputs(3750) <= a and b;
    layer3_outputs(3751) <= '1';
    layer3_outputs(3752) <= b;
    layer3_outputs(3753) <= not (a or b);
    layer3_outputs(3754) <= not b;
    layer3_outputs(3755) <= a or b;
    layer3_outputs(3756) <= not a;
    layer3_outputs(3757) <= not b or a;
    layer3_outputs(3758) <= not a;
    layer3_outputs(3759) <= a xor b;
    layer3_outputs(3760) <= not (a xor b);
    layer3_outputs(3761) <= not a or b;
    layer3_outputs(3762) <= '1';
    layer3_outputs(3763) <= a;
    layer3_outputs(3764) <= not (a or b);
    layer3_outputs(3765) <= a and not b;
    layer3_outputs(3766) <= a and b;
    layer3_outputs(3767) <= '1';
    layer3_outputs(3768) <= b and not a;
    layer3_outputs(3769) <= b;
    layer3_outputs(3770) <= not (a and b);
    layer3_outputs(3771) <= not (a and b);
    layer3_outputs(3772) <= not b;
    layer3_outputs(3773) <= '0';
    layer3_outputs(3774) <= '0';
    layer3_outputs(3775) <= not (a xor b);
    layer3_outputs(3776) <= not a or b;
    layer3_outputs(3777) <= not b or a;
    layer3_outputs(3778) <= not (a and b);
    layer3_outputs(3779) <= not (a and b);
    layer3_outputs(3780) <= not (a or b);
    layer3_outputs(3781) <= not b or a;
    layer3_outputs(3782) <= b;
    layer3_outputs(3783) <= not a;
    layer3_outputs(3784) <= a and not b;
    layer3_outputs(3785) <= not (a and b);
    layer3_outputs(3786) <= a xor b;
    layer3_outputs(3787) <= a and b;
    layer3_outputs(3788) <= b;
    layer3_outputs(3789) <= '1';
    layer3_outputs(3790) <= '1';
    layer3_outputs(3791) <= b;
    layer3_outputs(3792) <= not b or a;
    layer3_outputs(3793) <= not (a and b);
    layer3_outputs(3794) <= a;
    layer3_outputs(3795) <= b;
    layer3_outputs(3796) <= not a or b;
    layer3_outputs(3797) <= not (a and b);
    layer3_outputs(3798) <= a and not b;
    layer3_outputs(3799) <= b;
    layer3_outputs(3800) <= not (a or b);
    layer3_outputs(3801) <= not (a or b);
    layer3_outputs(3802) <= not b;
    layer3_outputs(3803) <= '0';
    layer3_outputs(3804) <= not (a and b);
    layer3_outputs(3805) <= a;
    layer3_outputs(3806) <= not b;
    layer3_outputs(3807) <= '1';
    layer3_outputs(3808) <= a and not b;
    layer3_outputs(3809) <= '0';
    layer3_outputs(3810) <= not b;
    layer3_outputs(3811) <= not (a xor b);
    layer3_outputs(3812) <= a xor b;
    layer3_outputs(3813) <= a and not b;
    layer3_outputs(3814) <= not b;
    layer3_outputs(3815) <= a;
    layer3_outputs(3816) <= b and not a;
    layer3_outputs(3817) <= a or b;
    layer3_outputs(3818) <= '0';
    layer3_outputs(3819) <= not b;
    layer3_outputs(3820) <= '0';
    layer3_outputs(3821) <= a or b;
    layer3_outputs(3822) <= b and not a;
    layer3_outputs(3823) <= b and not a;
    layer3_outputs(3824) <= not (a or b);
    layer3_outputs(3825) <= a;
    layer3_outputs(3826) <= not b or a;
    layer3_outputs(3827) <= not (a or b);
    layer3_outputs(3828) <= a or b;
    layer3_outputs(3829) <= not (a and b);
    layer3_outputs(3830) <= a xor b;
    layer3_outputs(3831) <= a xor b;
    layer3_outputs(3832) <= a xor b;
    layer3_outputs(3833) <= not b or a;
    layer3_outputs(3834) <= a;
    layer3_outputs(3835) <= a and not b;
    layer3_outputs(3836) <= '1';
    layer3_outputs(3837) <= not (a and b);
    layer3_outputs(3838) <= '0';
    layer3_outputs(3839) <= a and not b;
    layer3_outputs(3840) <= a and b;
    layer3_outputs(3841) <= not b or a;
    layer3_outputs(3842) <= '1';
    layer3_outputs(3843) <= not b;
    layer3_outputs(3844) <= not b;
    layer3_outputs(3845) <= '0';
    layer3_outputs(3846) <= '0';
    layer3_outputs(3847) <= '1';
    layer3_outputs(3848) <= not a or b;
    layer3_outputs(3849) <= a or b;
    layer3_outputs(3850) <= a xor b;
    layer3_outputs(3851) <= a and b;
    layer3_outputs(3852) <= a and b;
    layer3_outputs(3853) <= not a;
    layer3_outputs(3854) <= not b or a;
    layer3_outputs(3855) <= '0';
    layer3_outputs(3856) <= '1';
    layer3_outputs(3857) <= not (a or b);
    layer3_outputs(3858) <= not (a and b);
    layer3_outputs(3859) <= b;
    layer3_outputs(3860) <= not (a and b);
    layer3_outputs(3861) <= not a or b;
    layer3_outputs(3862) <= not (a or b);
    layer3_outputs(3863) <= not a;
    layer3_outputs(3864) <= b;
    layer3_outputs(3865) <= b;
    layer3_outputs(3866) <= not (a or b);
    layer3_outputs(3867) <= a and not b;
    layer3_outputs(3868) <= not a;
    layer3_outputs(3869) <= not b;
    layer3_outputs(3870) <= not b or a;
    layer3_outputs(3871) <= a and not b;
    layer3_outputs(3872) <= a and not b;
    layer3_outputs(3873) <= '1';
    layer3_outputs(3874) <= '1';
    layer3_outputs(3875) <= a or b;
    layer3_outputs(3876) <= not (a and b);
    layer3_outputs(3877) <= '1';
    layer3_outputs(3878) <= not (a xor b);
    layer3_outputs(3879) <= b and not a;
    layer3_outputs(3880) <= a;
    layer3_outputs(3881) <= a or b;
    layer3_outputs(3882) <= a and b;
    layer3_outputs(3883) <= '1';
    layer3_outputs(3884) <= not a or b;
    layer3_outputs(3885) <= not a;
    layer3_outputs(3886) <= a xor b;
    layer3_outputs(3887) <= b and not a;
    layer3_outputs(3888) <= a and b;
    layer3_outputs(3889) <= '0';
    layer3_outputs(3890) <= a or b;
    layer3_outputs(3891) <= not a;
    layer3_outputs(3892) <= a or b;
    layer3_outputs(3893) <= a;
    layer3_outputs(3894) <= not b;
    layer3_outputs(3895) <= a and b;
    layer3_outputs(3896) <= not b;
    layer3_outputs(3897) <= '1';
    layer3_outputs(3898) <= not (a or b);
    layer3_outputs(3899) <= not b;
    layer3_outputs(3900) <= '1';
    layer3_outputs(3901) <= not (a and b);
    layer3_outputs(3902) <= not a;
    layer3_outputs(3903) <= not a;
    layer3_outputs(3904) <= not b;
    layer3_outputs(3905) <= not b;
    layer3_outputs(3906) <= not a or b;
    layer3_outputs(3907) <= not b;
    layer3_outputs(3908) <= not (a or b);
    layer3_outputs(3909) <= b;
    layer3_outputs(3910) <= not b;
    layer3_outputs(3911) <= a or b;
    layer3_outputs(3912) <= b;
    layer3_outputs(3913) <= a or b;
    layer3_outputs(3914) <= '1';
    layer3_outputs(3915) <= not b or a;
    layer3_outputs(3916) <= '1';
    layer3_outputs(3917) <= b and not a;
    layer3_outputs(3918) <= '0';
    layer3_outputs(3919) <= a and not b;
    layer3_outputs(3920) <= not (a or b);
    layer3_outputs(3921) <= a xor b;
    layer3_outputs(3922) <= b;
    layer3_outputs(3923) <= not a;
    layer3_outputs(3924) <= not (a or b);
    layer3_outputs(3925) <= b;
    layer3_outputs(3926) <= a and b;
    layer3_outputs(3927) <= '0';
    layer3_outputs(3928) <= '1';
    layer3_outputs(3929) <= '1';
    layer3_outputs(3930) <= '1';
    layer3_outputs(3931) <= a and b;
    layer3_outputs(3932) <= not (a xor b);
    layer3_outputs(3933) <= '1';
    layer3_outputs(3934) <= '0';
    layer3_outputs(3935) <= b;
    layer3_outputs(3936) <= a;
    layer3_outputs(3937) <= not (a or b);
    layer3_outputs(3938) <= not (a and b);
    layer3_outputs(3939) <= not a or b;
    layer3_outputs(3940) <= '1';
    layer3_outputs(3941) <= not (a or b);
    layer3_outputs(3942) <= not (a or b);
    layer3_outputs(3943) <= not b;
    layer3_outputs(3944) <= a and b;
    layer3_outputs(3945) <= b and not a;
    layer3_outputs(3946) <= not b or a;
    layer3_outputs(3947) <= not b or a;
    layer3_outputs(3948) <= a and b;
    layer3_outputs(3949) <= '0';
    layer3_outputs(3950) <= a and b;
    layer3_outputs(3951) <= a and not b;
    layer3_outputs(3952) <= '0';
    layer3_outputs(3953) <= not a or b;
    layer3_outputs(3954) <= b and not a;
    layer3_outputs(3955) <= a or b;
    layer3_outputs(3956) <= a;
    layer3_outputs(3957) <= a and b;
    layer3_outputs(3958) <= a or b;
    layer3_outputs(3959) <= not a;
    layer3_outputs(3960) <= b;
    layer3_outputs(3961) <= not a;
    layer3_outputs(3962) <= not b or a;
    layer3_outputs(3963) <= a or b;
    layer3_outputs(3964) <= not b or a;
    layer3_outputs(3965) <= not a;
    layer3_outputs(3966) <= a and b;
    layer3_outputs(3967) <= b and not a;
    layer3_outputs(3968) <= not (a and b);
    layer3_outputs(3969) <= a;
    layer3_outputs(3970) <= b and not a;
    layer3_outputs(3971) <= a;
    layer3_outputs(3972) <= a and not b;
    layer3_outputs(3973) <= not a;
    layer3_outputs(3974) <= '1';
    layer3_outputs(3975) <= a;
    layer3_outputs(3976) <= a;
    layer3_outputs(3977) <= not (a or b);
    layer3_outputs(3978) <= '1';
    layer3_outputs(3979) <= a and b;
    layer3_outputs(3980) <= a xor b;
    layer3_outputs(3981) <= '0';
    layer3_outputs(3982) <= a;
    layer3_outputs(3983) <= not a or b;
    layer3_outputs(3984) <= '0';
    layer3_outputs(3985) <= not (a and b);
    layer3_outputs(3986) <= '1';
    layer3_outputs(3987) <= '0';
    layer3_outputs(3988) <= '0';
    layer3_outputs(3989) <= '0';
    layer3_outputs(3990) <= '1';
    layer3_outputs(3991) <= not a or b;
    layer3_outputs(3992) <= '1';
    layer3_outputs(3993) <= not (a or b);
    layer3_outputs(3994) <= not (a and b);
    layer3_outputs(3995) <= a and b;
    layer3_outputs(3996) <= a xor b;
    layer3_outputs(3997) <= a and not b;
    layer3_outputs(3998) <= not b or a;
    layer3_outputs(3999) <= not (a or b);
    layer3_outputs(4000) <= a and b;
    layer3_outputs(4001) <= not a;
    layer3_outputs(4002) <= a and b;
    layer3_outputs(4003) <= a xor b;
    layer3_outputs(4004) <= a and not b;
    layer3_outputs(4005) <= not a or b;
    layer3_outputs(4006) <= a or b;
    layer3_outputs(4007) <= '1';
    layer3_outputs(4008) <= b;
    layer3_outputs(4009) <= not (a or b);
    layer3_outputs(4010) <= not b or a;
    layer3_outputs(4011) <= '1';
    layer3_outputs(4012) <= '1';
    layer3_outputs(4013) <= not (a or b);
    layer3_outputs(4014) <= b;
    layer3_outputs(4015) <= not b or a;
    layer3_outputs(4016) <= not a;
    layer3_outputs(4017) <= b;
    layer3_outputs(4018) <= a or b;
    layer3_outputs(4019) <= '1';
    layer3_outputs(4020) <= b and not a;
    layer3_outputs(4021) <= not (a or b);
    layer3_outputs(4022) <= a or b;
    layer3_outputs(4023) <= b and not a;
    layer3_outputs(4024) <= '0';
    layer3_outputs(4025) <= a xor b;
    layer3_outputs(4026) <= not a or b;
    layer3_outputs(4027) <= not b;
    layer3_outputs(4028) <= a or b;
    layer3_outputs(4029) <= '0';
    layer3_outputs(4030) <= b;
    layer3_outputs(4031) <= '0';
    layer3_outputs(4032) <= not (a or b);
    layer3_outputs(4033) <= not a or b;
    layer3_outputs(4034) <= b;
    layer3_outputs(4035) <= b;
    layer3_outputs(4036) <= b and not a;
    layer3_outputs(4037) <= '0';
    layer3_outputs(4038) <= '0';
    layer3_outputs(4039) <= '1';
    layer3_outputs(4040) <= a and not b;
    layer3_outputs(4041) <= a;
    layer3_outputs(4042) <= a;
    layer3_outputs(4043) <= a xor b;
    layer3_outputs(4044) <= not (a and b);
    layer3_outputs(4045) <= a and b;
    layer3_outputs(4046) <= '1';
    layer3_outputs(4047) <= '1';
    layer3_outputs(4048) <= not a or b;
    layer3_outputs(4049) <= a and b;
    layer3_outputs(4050) <= not a or b;
    layer3_outputs(4051) <= a xor b;
    layer3_outputs(4052) <= a or b;
    layer3_outputs(4053) <= a or b;
    layer3_outputs(4054) <= not a or b;
    layer3_outputs(4055) <= a and not b;
    layer3_outputs(4056) <= not (a xor b);
    layer3_outputs(4057) <= b;
    layer3_outputs(4058) <= not a or b;
    layer3_outputs(4059) <= not b;
    layer3_outputs(4060) <= not (a or b);
    layer3_outputs(4061) <= not (a or b);
    layer3_outputs(4062) <= a or b;
    layer3_outputs(4063) <= a and not b;
    layer3_outputs(4064) <= b;
    layer3_outputs(4065) <= '1';
    layer3_outputs(4066) <= not a or b;
    layer3_outputs(4067) <= not b or a;
    layer3_outputs(4068) <= a or b;
    layer3_outputs(4069) <= not (a and b);
    layer3_outputs(4070) <= not (a or b);
    layer3_outputs(4071) <= b and not a;
    layer3_outputs(4072) <= b;
    layer3_outputs(4073) <= not b or a;
    layer3_outputs(4074) <= not a;
    layer3_outputs(4075) <= not b;
    layer3_outputs(4076) <= '0';
    layer3_outputs(4077) <= '1';
    layer3_outputs(4078) <= not (a or b);
    layer3_outputs(4079) <= b and not a;
    layer3_outputs(4080) <= a and not b;
    layer3_outputs(4081) <= not a or b;
    layer3_outputs(4082) <= not (a or b);
    layer3_outputs(4083) <= a and b;
    layer3_outputs(4084) <= a or b;
    layer3_outputs(4085) <= not b or a;
    layer3_outputs(4086) <= '1';
    layer3_outputs(4087) <= not (a or b);
    layer3_outputs(4088) <= b and not a;
    layer3_outputs(4089) <= not b;
    layer3_outputs(4090) <= '1';
    layer3_outputs(4091) <= a and not b;
    layer3_outputs(4092) <= a and b;
    layer3_outputs(4093) <= '0';
    layer3_outputs(4094) <= not (a or b);
    layer3_outputs(4095) <= not (a and b);
    layer3_outputs(4096) <= not a or b;
    layer3_outputs(4097) <= '1';
    layer3_outputs(4098) <= not b or a;
    layer3_outputs(4099) <= not b;
    layer3_outputs(4100) <= not (a and b);
    layer3_outputs(4101) <= not a or b;
    layer3_outputs(4102) <= not a or b;
    layer3_outputs(4103) <= b and not a;
    layer3_outputs(4104) <= not b;
    layer3_outputs(4105) <= not (a or b);
    layer3_outputs(4106) <= a or b;
    layer3_outputs(4107) <= not (a and b);
    layer3_outputs(4108) <= a or b;
    layer3_outputs(4109) <= not (a and b);
    layer3_outputs(4110) <= not (a and b);
    layer3_outputs(4111) <= not (a and b);
    layer3_outputs(4112) <= not b;
    layer3_outputs(4113) <= b;
    layer3_outputs(4114) <= a or b;
    layer3_outputs(4115) <= a or b;
    layer3_outputs(4116) <= not (a and b);
    layer3_outputs(4117) <= '1';
    layer3_outputs(4118) <= not (a or b);
    layer3_outputs(4119) <= not b or a;
    layer3_outputs(4120) <= '0';
    layer3_outputs(4121) <= b and not a;
    layer3_outputs(4122) <= not a or b;
    layer3_outputs(4123) <= not a;
    layer3_outputs(4124) <= '1';
    layer3_outputs(4125) <= not (a or b);
    layer3_outputs(4126) <= b;
    layer3_outputs(4127) <= '1';
    layer3_outputs(4128) <= not a;
    layer3_outputs(4129) <= b;
    layer3_outputs(4130) <= a and b;
    layer3_outputs(4131) <= a and b;
    layer3_outputs(4132) <= not a or b;
    layer3_outputs(4133) <= not (a or b);
    layer3_outputs(4134) <= not b or a;
    layer3_outputs(4135) <= not a or b;
    layer3_outputs(4136) <= '0';
    layer3_outputs(4137) <= a and b;
    layer3_outputs(4138) <= not a or b;
    layer3_outputs(4139) <= not b;
    layer3_outputs(4140) <= '1';
    layer3_outputs(4141) <= not b;
    layer3_outputs(4142) <= a;
    layer3_outputs(4143) <= not (a or b);
    layer3_outputs(4144) <= b and not a;
    layer3_outputs(4145) <= a or b;
    layer3_outputs(4146) <= not b or a;
    layer3_outputs(4147) <= b and not a;
    layer3_outputs(4148) <= not a or b;
    layer3_outputs(4149) <= not a or b;
    layer3_outputs(4150) <= '0';
    layer3_outputs(4151) <= not b or a;
    layer3_outputs(4152) <= a and b;
    layer3_outputs(4153) <= a;
    layer3_outputs(4154) <= not (a and b);
    layer3_outputs(4155) <= not a or b;
    layer3_outputs(4156) <= b;
    layer3_outputs(4157) <= '1';
    layer3_outputs(4158) <= not a;
    layer3_outputs(4159) <= not (a or b);
    layer3_outputs(4160) <= a and b;
    layer3_outputs(4161) <= '1';
    layer3_outputs(4162) <= not a or b;
    layer3_outputs(4163) <= '0';
    layer3_outputs(4164) <= not b;
    layer3_outputs(4165) <= not b;
    layer3_outputs(4166) <= b;
    layer3_outputs(4167) <= a or b;
    layer3_outputs(4168) <= '1';
    layer3_outputs(4169) <= b and not a;
    layer3_outputs(4170) <= '1';
    layer3_outputs(4171) <= a xor b;
    layer3_outputs(4172) <= not (a and b);
    layer3_outputs(4173) <= a and not b;
    layer3_outputs(4174) <= a or b;
    layer3_outputs(4175) <= a and not b;
    layer3_outputs(4176) <= a and not b;
    layer3_outputs(4177) <= '1';
    layer3_outputs(4178) <= not a or b;
    layer3_outputs(4179) <= '1';
    layer3_outputs(4180) <= b;
    layer3_outputs(4181) <= '1';
    layer3_outputs(4182) <= not (a and b);
    layer3_outputs(4183) <= a;
    layer3_outputs(4184) <= '1';
    layer3_outputs(4185) <= a or b;
    layer3_outputs(4186) <= '0';
    layer3_outputs(4187) <= not a or b;
    layer3_outputs(4188) <= a;
    layer3_outputs(4189) <= not b or a;
    layer3_outputs(4190) <= a and b;
    layer3_outputs(4191) <= a or b;
    layer3_outputs(4192) <= not b or a;
    layer3_outputs(4193) <= a and b;
    layer3_outputs(4194) <= b;
    layer3_outputs(4195) <= a xor b;
    layer3_outputs(4196) <= a and not b;
    layer3_outputs(4197) <= not b;
    layer3_outputs(4198) <= a and b;
    layer3_outputs(4199) <= not a or b;
    layer3_outputs(4200) <= b;
    layer3_outputs(4201) <= a and b;
    layer3_outputs(4202) <= not (a xor b);
    layer3_outputs(4203) <= not a or b;
    layer3_outputs(4204) <= not (a and b);
    layer3_outputs(4205) <= not a;
    layer3_outputs(4206) <= a xor b;
    layer3_outputs(4207) <= a or b;
    layer3_outputs(4208) <= a;
    layer3_outputs(4209) <= a or b;
    layer3_outputs(4210) <= '0';
    layer3_outputs(4211) <= a and not b;
    layer3_outputs(4212) <= not b;
    layer3_outputs(4213) <= a;
    layer3_outputs(4214) <= not a or b;
    layer3_outputs(4215) <= not a;
    layer3_outputs(4216) <= not b or a;
    layer3_outputs(4217) <= not b;
    layer3_outputs(4218) <= a or b;
    layer3_outputs(4219) <= b;
    layer3_outputs(4220) <= not b or a;
    layer3_outputs(4221) <= not (a and b);
    layer3_outputs(4222) <= '0';
    layer3_outputs(4223) <= not (a and b);
    layer3_outputs(4224) <= not b;
    layer3_outputs(4225) <= not b;
    layer3_outputs(4226) <= not (a and b);
    layer3_outputs(4227) <= a and b;
    layer3_outputs(4228) <= a and not b;
    layer3_outputs(4229) <= '0';
    layer3_outputs(4230) <= not b;
    layer3_outputs(4231) <= '1';
    layer3_outputs(4232) <= '1';
    layer3_outputs(4233) <= a or b;
    layer3_outputs(4234) <= a;
    layer3_outputs(4235) <= a xor b;
    layer3_outputs(4236) <= a or b;
    layer3_outputs(4237) <= not b;
    layer3_outputs(4238) <= not a or b;
    layer3_outputs(4239) <= a or b;
    layer3_outputs(4240) <= not b;
    layer3_outputs(4241) <= not (a and b);
    layer3_outputs(4242) <= '0';
    layer3_outputs(4243) <= a or b;
    layer3_outputs(4244) <= b;
    layer3_outputs(4245) <= a;
    layer3_outputs(4246) <= not b;
    layer3_outputs(4247) <= not a;
    layer3_outputs(4248) <= a or b;
    layer3_outputs(4249) <= b;
    layer3_outputs(4250) <= a and b;
    layer3_outputs(4251) <= a and b;
    layer3_outputs(4252) <= a or b;
    layer3_outputs(4253) <= b;
    layer3_outputs(4254) <= a xor b;
    layer3_outputs(4255) <= not b or a;
    layer3_outputs(4256) <= '0';
    layer3_outputs(4257) <= a and not b;
    layer3_outputs(4258) <= not (a and b);
    layer3_outputs(4259) <= not (a xor b);
    layer3_outputs(4260) <= not a;
    layer3_outputs(4261) <= not (a and b);
    layer3_outputs(4262) <= a and not b;
    layer3_outputs(4263) <= '1';
    layer3_outputs(4264) <= not b or a;
    layer3_outputs(4265) <= not (a and b);
    layer3_outputs(4266) <= not (a and b);
    layer3_outputs(4267) <= '0';
    layer3_outputs(4268) <= a and not b;
    layer3_outputs(4269) <= not (a or b);
    layer3_outputs(4270) <= a;
    layer3_outputs(4271) <= a and b;
    layer3_outputs(4272) <= a or b;
    layer3_outputs(4273) <= a xor b;
    layer3_outputs(4274) <= not (a or b);
    layer3_outputs(4275) <= a or b;
    layer3_outputs(4276) <= a and not b;
    layer3_outputs(4277) <= not b;
    layer3_outputs(4278) <= not (a xor b);
    layer3_outputs(4279) <= a and b;
    layer3_outputs(4280) <= not b;
    layer3_outputs(4281) <= not (a or b);
    layer3_outputs(4282) <= not a;
    layer3_outputs(4283) <= not (a or b);
    layer3_outputs(4284) <= b;
    layer3_outputs(4285) <= b;
    layer3_outputs(4286) <= not b or a;
    layer3_outputs(4287) <= a and not b;
    layer3_outputs(4288) <= a and not b;
    layer3_outputs(4289) <= not a or b;
    layer3_outputs(4290) <= not a or b;
    layer3_outputs(4291) <= b;
    layer3_outputs(4292) <= '0';
    layer3_outputs(4293) <= a or b;
    layer3_outputs(4294) <= b;
    layer3_outputs(4295) <= not (a xor b);
    layer3_outputs(4296) <= not (a or b);
    layer3_outputs(4297) <= '0';
    layer3_outputs(4298) <= not (a or b);
    layer3_outputs(4299) <= '1';
    layer3_outputs(4300) <= not b;
    layer3_outputs(4301) <= not (a or b);
    layer3_outputs(4302) <= b and not a;
    layer3_outputs(4303) <= not a or b;
    layer3_outputs(4304) <= b;
    layer3_outputs(4305) <= '0';
    layer3_outputs(4306) <= a and not b;
    layer3_outputs(4307) <= not (a xor b);
    layer3_outputs(4308) <= '0';
    layer3_outputs(4309) <= b;
    layer3_outputs(4310) <= a and b;
    layer3_outputs(4311) <= a;
    layer3_outputs(4312) <= b;
    layer3_outputs(4313) <= not b or a;
    layer3_outputs(4314) <= b and not a;
    layer3_outputs(4315) <= not a;
    layer3_outputs(4316) <= not (a and b);
    layer3_outputs(4317) <= a and not b;
    layer3_outputs(4318) <= a and not b;
    layer3_outputs(4319) <= a;
    layer3_outputs(4320) <= not a or b;
    layer3_outputs(4321) <= a and b;
    layer3_outputs(4322) <= not a or b;
    layer3_outputs(4323) <= not b or a;
    layer3_outputs(4324) <= a;
    layer3_outputs(4325) <= a and b;
    layer3_outputs(4326) <= b and not a;
    layer3_outputs(4327) <= not b;
    layer3_outputs(4328) <= a and b;
    layer3_outputs(4329) <= '1';
    layer3_outputs(4330) <= '0';
    layer3_outputs(4331) <= a;
    layer3_outputs(4332) <= b and not a;
    layer3_outputs(4333) <= a;
    layer3_outputs(4334) <= not b;
    layer3_outputs(4335) <= not b;
    layer3_outputs(4336) <= not (a or b);
    layer3_outputs(4337) <= a and not b;
    layer3_outputs(4338) <= not (a and b);
    layer3_outputs(4339) <= a and b;
    layer3_outputs(4340) <= not a or b;
    layer3_outputs(4341) <= b and not a;
    layer3_outputs(4342) <= b;
    layer3_outputs(4343) <= a;
    layer3_outputs(4344) <= not (a or b);
    layer3_outputs(4345) <= '0';
    layer3_outputs(4346) <= b and not a;
    layer3_outputs(4347) <= '0';
    layer3_outputs(4348) <= b and not a;
    layer3_outputs(4349) <= a and not b;
    layer3_outputs(4350) <= b;
    layer3_outputs(4351) <= b;
    layer3_outputs(4352) <= a;
    layer3_outputs(4353) <= not a;
    layer3_outputs(4354) <= not b or a;
    layer3_outputs(4355) <= a and not b;
    layer3_outputs(4356) <= not b;
    layer3_outputs(4357) <= a;
    layer3_outputs(4358) <= not a or b;
    layer3_outputs(4359) <= not a or b;
    layer3_outputs(4360) <= b and not a;
    layer3_outputs(4361) <= a xor b;
    layer3_outputs(4362) <= not (a and b);
    layer3_outputs(4363) <= not b;
    layer3_outputs(4364) <= not a;
    layer3_outputs(4365) <= a and not b;
    layer3_outputs(4366) <= b and not a;
    layer3_outputs(4367) <= a;
    layer3_outputs(4368) <= not b or a;
    layer3_outputs(4369) <= not a;
    layer3_outputs(4370) <= a xor b;
    layer3_outputs(4371) <= not b or a;
    layer3_outputs(4372) <= b and not a;
    layer3_outputs(4373) <= not b or a;
    layer3_outputs(4374) <= '1';
    layer3_outputs(4375) <= not b;
    layer3_outputs(4376) <= not a or b;
    layer3_outputs(4377) <= '1';
    layer3_outputs(4378) <= not a;
    layer3_outputs(4379) <= b and not a;
    layer3_outputs(4380) <= not (a or b);
    layer3_outputs(4381) <= not a;
    layer3_outputs(4382) <= '1';
    layer3_outputs(4383) <= not b or a;
    layer3_outputs(4384) <= a and b;
    layer3_outputs(4385) <= b and not a;
    layer3_outputs(4386) <= '0';
    layer3_outputs(4387) <= a and b;
    layer3_outputs(4388) <= not (a or b);
    layer3_outputs(4389) <= '1';
    layer3_outputs(4390) <= a and not b;
    layer3_outputs(4391) <= a and b;
    layer3_outputs(4392) <= not a or b;
    layer3_outputs(4393) <= not b;
    layer3_outputs(4394) <= b;
    layer3_outputs(4395) <= not (a or b);
    layer3_outputs(4396) <= a and b;
    layer3_outputs(4397) <= not a or b;
    layer3_outputs(4398) <= not a or b;
    layer3_outputs(4399) <= a or b;
    layer3_outputs(4400) <= not (a or b);
    layer3_outputs(4401) <= not (a and b);
    layer3_outputs(4402) <= '0';
    layer3_outputs(4403) <= not a or b;
    layer3_outputs(4404) <= not a;
    layer3_outputs(4405) <= not a or b;
    layer3_outputs(4406) <= not (a or b);
    layer3_outputs(4407) <= not (a and b);
    layer3_outputs(4408) <= not (a and b);
    layer3_outputs(4409) <= '1';
    layer3_outputs(4410) <= '0';
    layer3_outputs(4411) <= '1';
    layer3_outputs(4412) <= not (a and b);
    layer3_outputs(4413) <= a;
    layer3_outputs(4414) <= '0';
    layer3_outputs(4415) <= not a or b;
    layer3_outputs(4416) <= not b or a;
    layer3_outputs(4417) <= not b;
    layer3_outputs(4418) <= not a;
    layer3_outputs(4419) <= a and not b;
    layer3_outputs(4420) <= '1';
    layer3_outputs(4421) <= not (a xor b);
    layer3_outputs(4422) <= not a;
    layer3_outputs(4423) <= b and not a;
    layer3_outputs(4424) <= a;
    layer3_outputs(4425) <= b and not a;
    layer3_outputs(4426) <= not (a and b);
    layer3_outputs(4427) <= not b;
    layer3_outputs(4428) <= not (a and b);
    layer3_outputs(4429) <= not b or a;
    layer3_outputs(4430) <= a and not b;
    layer3_outputs(4431) <= not (a and b);
    layer3_outputs(4432) <= a;
    layer3_outputs(4433) <= a;
    layer3_outputs(4434) <= not a or b;
    layer3_outputs(4435) <= not b or a;
    layer3_outputs(4436) <= not a;
    layer3_outputs(4437) <= b;
    layer3_outputs(4438) <= a xor b;
    layer3_outputs(4439) <= a and b;
    layer3_outputs(4440) <= not b;
    layer3_outputs(4441) <= b;
    layer3_outputs(4442) <= '0';
    layer3_outputs(4443) <= b and not a;
    layer3_outputs(4444) <= b and not a;
    layer3_outputs(4445) <= a and not b;
    layer3_outputs(4446) <= '1';
    layer3_outputs(4447) <= not b or a;
    layer3_outputs(4448) <= a;
    layer3_outputs(4449) <= not a;
    layer3_outputs(4450) <= not b or a;
    layer3_outputs(4451) <= not a or b;
    layer3_outputs(4452) <= b and not a;
    layer3_outputs(4453) <= not a or b;
    layer3_outputs(4454) <= not (a and b);
    layer3_outputs(4455) <= not a;
    layer3_outputs(4456) <= b and not a;
    layer3_outputs(4457) <= b;
    layer3_outputs(4458) <= b;
    layer3_outputs(4459) <= b;
    layer3_outputs(4460) <= a;
    layer3_outputs(4461) <= not a;
    layer3_outputs(4462) <= a or b;
    layer3_outputs(4463) <= not (a xor b);
    layer3_outputs(4464) <= '1';
    layer3_outputs(4465) <= a;
    layer3_outputs(4466) <= not a;
    layer3_outputs(4467) <= not b or a;
    layer3_outputs(4468) <= b;
    layer3_outputs(4469) <= not b or a;
    layer3_outputs(4470) <= b;
    layer3_outputs(4471) <= '1';
    layer3_outputs(4472) <= b and not a;
    layer3_outputs(4473) <= not b;
    layer3_outputs(4474) <= a and b;
    layer3_outputs(4475) <= '1';
    layer3_outputs(4476) <= not b or a;
    layer3_outputs(4477) <= a or b;
    layer3_outputs(4478) <= a and not b;
    layer3_outputs(4479) <= not a;
    layer3_outputs(4480) <= not b;
    layer3_outputs(4481) <= not b or a;
    layer3_outputs(4482) <= not b;
    layer3_outputs(4483) <= a or b;
    layer3_outputs(4484) <= b and not a;
    layer3_outputs(4485) <= b;
    layer3_outputs(4486) <= not a or b;
    layer3_outputs(4487) <= not (a or b);
    layer3_outputs(4488) <= not (a or b);
    layer3_outputs(4489) <= b and not a;
    layer3_outputs(4490) <= not b;
    layer3_outputs(4491) <= a and not b;
    layer3_outputs(4492) <= a and not b;
    layer3_outputs(4493) <= not (a or b);
    layer3_outputs(4494) <= '0';
    layer3_outputs(4495) <= a and not b;
    layer3_outputs(4496) <= b;
    layer3_outputs(4497) <= not (a and b);
    layer3_outputs(4498) <= '0';
    layer3_outputs(4499) <= '1';
    layer3_outputs(4500) <= '0';
    layer3_outputs(4501) <= not (a or b);
    layer3_outputs(4502) <= not (a or b);
    layer3_outputs(4503) <= not a;
    layer3_outputs(4504) <= a or b;
    layer3_outputs(4505) <= not b;
    layer3_outputs(4506) <= '1';
    layer3_outputs(4507) <= '0';
    layer3_outputs(4508) <= not a;
    layer3_outputs(4509) <= not (a and b);
    layer3_outputs(4510) <= not a or b;
    layer3_outputs(4511) <= '1';
    layer3_outputs(4512) <= not a;
    layer3_outputs(4513) <= a and not b;
    layer3_outputs(4514) <= a and not b;
    layer3_outputs(4515) <= a and b;
    layer3_outputs(4516) <= not b or a;
    layer3_outputs(4517) <= a and not b;
    layer3_outputs(4518) <= not (a and b);
    layer3_outputs(4519) <= '0';
    layer3_outputs(4520) <= a;
    layer3_outputs(4521) <= a and not b;
    layer3_outputs(4522) <= b and not a;
    layer3_outputs(4523) <= not b;
    layer3_outputs(4524) <= not a;
    layer3_outputs(4525) <= a and b;
    layer3_outputs(4526) <= not b;
    layer3_outputs(4527) <= '1';
    layer3_outputs(4528) <= not b;
    layer3_outputs(4529) <= a and b;
    layer3_outputs(4530) <= a;
    layer3_outputs(4531) <= b and not a;
    layer3_outputs(4532) <= b and not a;
    layer3_outputs(4533) <= b and not a;
    layer3_outputs(4534) <= b;
    layer3_outputs(4535) <= not (a or b);
    layer3_outputs(4536) <= not (a or b);
    layer3_outputs(4537) <= a xor b;
    layer3_outputs(4538) <= not (a and b);
    layer3_outputs(4539) <= a or b;
    layer3_outputs(4540) <= b;
    layer3_outputs(4541) <= b and not a;
    layer3_outputs(4542) <= not (a xor b);
    layer3_outputs(4543) <= a;
    layer3_outputs(4544) <= not (a and b);
    layer3_outputs(4545) <= not a;
    layer3_outputs(4546) <= b;
    layer3_outputs(4547) <= '1';
    layer3_outputs(4548) <= a;
    layer3_outputs(4549) <= not a;
    layer3_outputs(4550) <= a or b;
    layer3_outputs(4551) <= not a or b;
    layer3_outputs(4552) <= not b;
    layer3_outputs(4553) <= a and not b;
    layer3_outputs(4554) <= a and b;
    layer3_outputs(4555) <= not (a and b);
    layer3_outputs(4556) <= '0';
    layer3_outputs(4557) <= a xor b;
    layer3_outputs(4558) <= '1';
    layer3_outputs(4559) <= a xor b;
    layer3_outputs(4560) <= a and b;
    layer3_outputs(4561) <= not a or b;
    layer3_outputs(4562) <= not a;
    layer3_outputs(4563) <= a;
    layer3_outputs(4564) <= not b;
    layer3_outputs(4565) <= a;
    layer3_outputs(4566) <= not (a or b);
    layer3_outputs(4567) <= b and not a;
    layer3_outputs(4568) <= a or b;
    layer3_outputs(4569) <= a xor b;
    layer3_outputs(4570) <= not b;
    layer3_outputs(4571) <= not (a or b);
    layer3_outputs(4572) <= not b;
    layer3_outputs(4573) <= not b or a;
    layer3_outputs(4574) <= not (a and b);
    layer3_outputs(4575) <= not (a or b);
    layer3_outputs(4576) <= not a or b;
    layer3_outputs(4577) <= b;
    layer3_outputs(4578) <= not a;
    layer3_outputs(4579) <= a and not b;
    layer3_outputs(4580) <= not (a xor b);
    layer3_outputs(4581) <= a and not b;
    layer3_outputs(4582) <= a or b;
    layer3_outputs(4583) <= a or b;
    layer3_outputs(4584) <= a or b;
    layer3_outputs(4585) <= a and not b;
    layer3_outputs(4586) <= not b or a;
    layer3_outputs(4587) <= not (a and b);
    layer3_outputs(4588) <= b;
    layer3_outputs(4589) <= not b;
    layer3_outputs(4590) <= not b;
    layer3_outputs(4591) <= '0';
    layer3_outputs(4592) <= a or b;
    layer3_outputs(4593) <= not a or b;
    layer3_outputs(4594) <= not b or a;
    layer3_outputs(4595) <= '0';
    layer3_outputs(4596) <= a;
    layer3_outputs(4597) <= not (a xor b);
    layer3_outputs(4598) <= not (a or b);
    layer3_outputs(4599) <= not (a and b);
    layer3_outputs(4600) <= not b;
    layer3_outputs(4601) <= a;
    layer3_outputs(4602) <= a or b;
    layer3_outputs(4603) <= a and b;
    layer3_outputs(4604) <= not b or a;
    layer3_outputs(4605) <= '0';
    layer3_outputs(4606) <= not b or a;
    layer3_outputs(4607) <= a xor b;
    layer3_outputs(4608) <= a and not b;
    layer3_outputs(4609) <= '1';
    layer3_outputs(4610) <= a or b;
    layer3_outputs(4611) <= not (a xor b);
    layer3_outputs(4612) <= not (a and b);
    layer3_outputs(4613) <= b;
    layer3_outputs(4614) <= a;
    layer3_outputs(4615) <= a or b;
    layer3_outputs(4616) <= a and b;
    layer3_outputs(4617) <= not a;
    layer3_outputs(4618) <= a;
    layer3_outputs(4619) <= b and not a;
    layer3_outputs(4620) <= '1';
    layer3_outputs(4621) <= not a or b;
    layer3_outputs(4622) <= '0';
    layer3_outputs(4623) <= not b or a;
    layer3_outputs(4624) <= not b or a;
    layer3_outputs(4625) <= not (a or b);
    layer3_outputs(4626) <= not (a or b);
    layer3_outputs(4627) <= a and not b;
    layer3_outputs(4628) <= not (a and b);
    layer3_outputs(4629) <= a and not b;
    layer3_outputs(4630) <= b and not a;
    layer3_outputs(4631) <= not a;
    layer3_outputs(4632) <= a or b;
    layer3_outputs(4633) <= not (a xor b);
    layer3_outputs(4634) <= '1';
    layer3_outputs(4635) <= not (a or b);
    layer3_outputs(4636) <= b and not a;
    layer3_outputs(4637) <= b and not a;
    layer3_outputs(4638) <= a or b;
    layer3_outputs(4639) <= not (a or b);
    layer3_outputs(4640) <= a xor b;
    layer3_outputs(4641) <= a xor b;
    layer3_outputs(4642) <= not a;
    layer3_outputs(4643) <= a or b;
    layer3_outputs(4644) <= not b;
    layer3_outputs(4645) <= not b or a;
    layer3_outputs(4646) <= not (a and b);
    layer3_outputs(4647) <= a and b;
    layer3_outputs(4648) <= a and not b;
    layer3_outputs(4649) <= a or b;
    layer3_outputs(4650) <= not a;
    layer3_outputs(4651) <= not (a and b);
    layer3_outputs(4652) <= not (a or b);
    layer3_outputs(4653) <= a and not b;
    layer3_outputs(4654) <= b and not a;
    layer3_outputs(4655) <= not (a or b);
    layer3_outputs(4656) <= not b or a;
    layer3_outputs(4657) <= not a or b;
    layer3_outputs(4658) <= a or b;
    layer3_outputs(4659) <= a;
    layer3_outputs(4660) <= not a;
    layer3_outputs(4661) <= '1';
    layer3_outputs(4662) <= not (a or b);
    layer3_outputs(4663) <= a and b;
    layer3_outputs(4664) <= not (a or b);
    layer3_outputs(4665) <= a or b;
    layer3_outputs(4666) <= b;
    layer3_outputs(4667) <= not a or b;
    layer3_outputs(4668) <= a and b;
    layer3_outputs(4669) <= not a or b;
    layer3_outputs(4670) <= a and b;
    layer3_outputs(4671) <= b;
    layer3_outputs(4672) <= a and not b;
    layer3_outputs(4673) <= not b or a;
    layer3_outputs(4674) <= not b or a;
    layer3_outputs(4675) <= not a;
    layer3_outputs(4676) <= not b or a;
    layer3_outputs(4677) <= not a or b;
    layer3_outputs(4678) <= b and not a;
    layer3_outputs(4679) <= '0';
    layer3_outputs(4680) <= not b;
    layer3_outputs(4681) <= b and not a;
    layer3_outputs(4682) <= not (a and b);
    layer3_outputs(4683) <= b and not a;
    layer3_outputs(4684) <= not b;
    layer3_outputs(4685) <= not (a and b);
    layer3_outputs(4686) <= b and not a;
    layer3_outputs(4687) <= b and not a;
    layer3_outputs(4688) <= a or b;
    layer3_outputs(4689) <= not a or b;
    layer3_outputs(4690) <= a;
    layer3_outputs(4691) <= a and not b;
    layer3_outputs(4692) <= not b;
    layer3_outputs(4693) <= '1';
    layer3_outputs(4694) <= not (a or b);
    layer3_outputs(4695) <= not (a xor b);
    layer3_outputs(4696) <= not (a xor b);
    layer3_outputs(4697) <= not b;
    layer3_outputs(4698) <= b and not a;
    layer3_outputs(4699) <= b and not a;
    layer3_outputs(4700) <= not a or b;
    layer3_outputs(4701) <= not b or a;
    layer3_outputs(4702) <= not (a xor b);
    layer3_outputs(4703) <= not a;
    layer3_outputs(4704) <= not a or b;
    layer3_outputs(4705) <= not (a or b);
    layer3_outputs(4706) <= '1';
    layer3_outputs(4707) <= not a;
    layer3_outputs(4708) <= not (a and b);
    layer3_outputs(4709) <= b and not a;
    layer3_outputs(4710) <= b and not a;
    layer3_outputs(4711) <= not (a and b);
    layer3_outputs(4712) <= not b;
    layer3_outputs(4713) <= not b or a;
    layer3_outputs(4714) <= b and not a;
    layer3_outputs(4715) <= not a;
    layer3_outputs(4716) <= '1';
    layer3_outputs(4717) <= a and not b;
    layer3_outputs(4718) <= '0';
    layer3_outputs(4719) <= '0';
    layer3_outputs(4720) <= a or b;
    layer3_outputs(4721) <= a xor b;
    layer3_outputs(4722) <= not (a or b);
    layer3_outputs(4723) <= '0';
    layer3_outputs(4724) <= not b;
    layer3_outputs(4725) <= a;
    layer3_outputs(4726) <= a and b;
    layer3_outputs(4727) <= not (a and b);
    layer3_outputs(4728) <= a and b;
    layer3_outputs(4729) <= not (a xor b);
    layer3_outputs(4730) <= b;
    layer3_outputs(4731) <= not (a and b);
    layer3_outputs(4732) <= b;
    layer3_outputs(4733) <= not b or a;
    layer3_outputs(4734) <= not a;
    layer3_outputs(4735) <= not b;
    layer3_outputs(4736) <= not (a or b);
    layer3_outputs(4737) <= a and not b;
    layer3_outputs(4738) <= not b or a;
    layer3_outputs(4739) <= not (a and b);
    layer3_outputs(4740) <= a;
    layer3_outputs(4741) <= a;
    layer3_outputs(4742) <= not (a and b);
    layer3_outputs(4743) <= not b;
    layer3_outputs(4744) <= not a;
    layer3_outputs(4745) <= '1';
    layer3_outputs(4746) <= not (a and b);
    layer3_outputs(4747) <= a and b;
    layer3_outputs(4748) <= not a;
    layer3_outputs(4749) <= not (a and b);
    layer3_outputs(4750) <= not a;
    layer3_outputs(4751) <= a and b;
    layer3_outputs(4752) <= '1';
    layer3_outputs(4753) <= b and not a;
    layer3_outputs(4754) <= a or b;
    layer3_outputs(4755) <= a;
    layer3_outputs(4756) <= a and b;
    layer3_outputs(4757) <= b;
    layer3_outputs(4758) <= a xor b;
    layer3_outputs(4759) <= '0';
    layer3_outputs(4760) <= not a or b;
    layer3_outputs(4761) <= a;
    layer3_outputs(4762) <= not a;
    layer3_outputs(4763) <= not (a or b);
    layer3_outputs(4764) <= not b;
    layer3_outputs(4765) <= '0';
    layer3_outputs(4766) <= not (a or b);
    layer3_outputs(4767) <= b;
    layer3_outputs(4768) <= not b;
    layer3_outputs(4769) <= not (a xor b);
    layer3_outputs(4770) <= not a or b;
    layer3_outputs(4771) <= not b or a;
    layer3_outputs(4772) <= b and not a;
    layer3_outputs(4773) <= a and b;
    layer3_outputs(4774) <= '1';
    layer3_outputs(4775) <= not a;
    layer3_outputs(4776) <= '1';
    layer3_outputs(4777) <= not a;
    layer3_outputs(4778) <= b and not a;
    layer3_outputs(4779) <= '0';
    layer3_outputs(4780) <= not b or a;
    layer3_outputs(4781) <= a or b;
    layer3_outputs(4782) <= not a or b;
    layer3_outputs(4783) <= not (a and b);
    layer3_outputs(4784) <= '0';
    layer3_outputs(4785) <= not (a or b);
    layer3_outputs(4786) <= not a or b;
    layer3_outputs(4787) <= not (a or b);
    layer3_outputs(4788) <= '1';
    layer3_outputs(4789) <= not (a and b);
    layer3_outputs(4790) <= '0';
    layer3_outputs(4791) <= '1';
    layer3_outputs(4792) <= a and b;
    layer3_outputs(4793) <= a and b;
    layer3_outputs(4794) <= not a;
    layer3_outputs(4795) <= b;
    layer3_outputs(4796) <= not b or a;
    layer3_outputs(4797) <= a xor b;
    layer3_outputs(4798) <= not b;
    layer3_outputs(4799) <= not (a and b);
    layer3_outputs(4800) <= a or b;
    layer3_outputs(4801) <= not b;
    layer3_outputs(4802) <= not (a and b);
    layer3_outputs(4803) <= not b or a;
    layer3_outputs(4804) <= '0';
    layer3_outputs(4805) <= a and b;
    layer3_outputs(4806) <= b and not a;
    layer3_outputs(4807) <= '1';
    layer3_outputs(4808) <= b and not a;
    layer3_outputs(4809) <= a and not b;
    layer3_outputs(4810) <= '1';
    layer3_outputs(4811) <= b;
    layer3_outputs(4812) <= not (a and b);
    layer3_outputs(4813) <= not a or b;
    layer3_outputs(4814) <= '1';
    layer3_outputs(4815) <= not a or b;
    layer3_outputs(4816) <= a and b;
    layer3_outputs(4817) <= a;
    layer3_outputs(4818) <= not (a or b);
    layer3_outputs(4819) <= not a or b;
    layer3_outputs(4820) <= not (a and b);
    layer3_outputs(4821) <= not b;
    layer3_outputs(4822) <= b and not a;
    layer3_outputs(4823) <= '1';
    layer3_outputs(4824) <= a;
    layer3_outputs(4825) <= a xor b;
    layer3_outputs(4826) <= '1';
    layer3_outputs(4827) <= not a or b;
    layer3_outputs(4828) <= a and not b;
    layer3_outputs(4829) <= a or b;
    layer3_outputs(4830) <= '1';
    layer3_outputs(4831) <= b;
    layer3_outputs(4832) <= '1';
    layer3_outputs(4833) <= a and b;
    layer3_outputs(4834) <= '1';
    layer3_outputs(4835) <= '1';
    layer3_outputs(4836) <= a and b;
    layer3_outputs(4837) <= '1';
    layer3_outputs(4838) <= not a or b;
    layer3_outputs(4839) <= b and not a;
    layer3_outputs(4840) <= not a;
    layer3_outputs(4841) <= not (a and b);
    layer3_outputs(4842) <= not b or a;
    layer3_outputs(4843) <= b and not a;
    layer3_outputs(4844) <= not a or b;
    layer3_outputs(4845) <= a and b;
    layer3_outputs(4846) <= b;
    layer3_outputs(4847) <= not a;
    layer3_outputs(4848) <= a and not b;
    layer3_outputs(4849) <= a;
    layer3_outputs(4850) <= not b or a;
    layer3_outputs(4851) <= not (a xor b);
    layer3_outputs(4852) <= '0';
    layer3_outputs(4853) <= b;
    layer3_outputs(4854) <= a;
    layer3_outputs(4855) <= not (a or b);
    layer3_outputs(4856) <= not b;
    layer3_outputs(4857) <= b;
    layer3_outputs(4858) <= not b;
    layer3_outputs(4859) <= b;
    layer3_outputs(4860) <= not a;
    layer3_outputs(4861) <= not b or a;
    layer3_outputs(4862) <= not b;
    layer3_outputs(4863) <= '0';
    layer3_outputs(4864) <= not (a or b);
    layer3_outputs(4865) <= a or b;
    layer3_outputs(4866) <= a and not b;
    layer3_outputs(4867) <= '0';
    layer3_outputs(4868) <= not a or b;
    layer3_outputs(4869) <= a;
    layer3_outputs(4870) <= b;
    layer3_outputs(4871) <= a;
    layer3_outputs(4872) <= not (a or b);
    layer3_outputs(4873) <= not (a and b);
    layer3_outputs(4874) <= b and not a;
    layer3_outputs(4875) <= a xor b;
    layer3_outputs(4876) <= not (a and b);
    layer3_outputs(4877) <= '1';
    layer3_outputs(4878) <= not (a or b);
    layer3_outputs(4879) <= not a;
    layer3_outputs(4880) <= '1';
    layer3_outputs(4881) <= not b;
    layer3_outputs(4882) <= '0';
    layer3_outputs(4883) <= a and b;
    layer3_outputs(4884) <= '1';
    layer3_outputs(4885) <= a and not b;
    layer3_outputs(4886) <= not a or b;
    layer3_outputs(4887) <= not a;
    layer3_outputs(4888) <= not (a xor b);
    layer3_outputs(4889) <= not a or b;
    layer3_outputs(4890) <= not a;
    layer3_outputs(4891) <= a xor b;
    layer3_outputs(4892) <= not b or a;
    layer3_outputs(4893) <= '0';
    layer3_outputs(4894) <= '0';
    layer3_outputs(4895) <= a and b;
    layer3_outputs(4896) <= not (a or b);
    layer3_outputs(4897) <= '1';
    layer3_outputs(4898) <= a and not b;
    layer3_outputs(4899) <= a and not b;
    layer3_outputs(4900) <= a or b;
    layer3_outputs(4901) <= not a or b;
    layer3_outputs(4902) <= not (a or b);
    layer3_outputs(4903) <= a and b;
    layer3_outputs(4904) <= not a;
    layer3_outputs(4905) <= not a or b;
    layer3_outputs(4906) <= not a or b;
    layer3_outputs(4907) <= not a;
    layer3_outputs(4908) <= b;
    layer3_outputs(4909) <= a or b;
    layer3_outputs(4910) <= not (a or b);
    layer3_outputs(4911) <= '0';
    layer3_outputs(4912) <= a or b;
    layer3_outputs(4913) <= not (a or b);
    layer3_outputs(4914) <= a;
    layer3_outputs(4915) <= a or b;
    layer3_outputs(4916) <= not (a and b);
    layer3_outputs(4917) <= a;
    layer3_outputs(4918) <= not a or b;
    layer3_outputs(4919) <= not (a and b);
    layer3_outputs(4920) <= b;
    layer3_outputs(4921) <= a xor b;
    layer3_outputs(4922) <= not a;
    layer3_outputs(4923) <= a;
    layer3_outputs(4924) <= not b;
    layer3_outputs(4925) <= a xor b;
    layer3_outputs(4926) <= a and b;
    layer3_outputs(4927) <= a or b;
    layer3_outputs(4928) <= not (a and b);
    layer3_outputs(4929) <= '1';
    layer3_outputs(4930) <= not (a or b);
    layer3_outputs(4931) <= a;
    layer3_outputs(4932) <= a and b;
    layer3_outputs(4933) <= not (a and b);
    layer3_outputs(4934) <= not a;
    layer3_outputs(4935) <= '0';
    layer3_outputs(4936) <= '1';
    layer3_outputs(4937) <= '1';
    layer3_outputs(4938) <= '0';
    layer3_outputs(4939) <= not b or a;
    layer3_outputs(4940) <= a;
    layer3_outputs(4941) <= a or b;
    layer3_outputs(4942) <= not b;
    layer3_outputs(4943) <= b;
    layer3_outputs(4944) <= '1';
    layer3_outputs(4945) <= b;
    layer3_outputs(4946) <= b;
    layer3_outputs(4947) <= not (a and b);
    layer3_outputs(4948) <= a;
    layer3_outputs(4949) <= b;
    layer3_outputs(4950) <= a and not b;
    layer3_outputs(4951) <= '1';
    layer3_outputs(4952) <= '1';
    layer3_outputs(4953) <= not b;
    layer3_outputs(4954) <= '1';
    layer3_outputs(4955) <= not (a and b);
    layer3_outputs(4956) <= '1';
    layer3_outputs(4957) <= not (a xor b);
    layer3_outputs(4958) <= not b or a;
    layer3_outputs(4959) <= not a or b;
    layer3_outputs(4960) <= '1';
    layer3_outputs(4961) <= a and b;
    layer3_outputs(4962) <= a and not b;
    layer3_outputs(4963) <= not (a and b);
    layer3_outputs(4964) <= b;
    layer3_outputs(4965) <= not b or a;
    layer3_outputs(4966) <= a;
    layer3_outputs(4967) <= not b or a;
    layer3_outputs(4968) <= b and not a;
    layer3_outputs(4969) <= a and not b;
    layer3_outputs(4970) <= b;
    layer3_outputs(4971) <= a and not b;
    layer3_outputs(4972) <= a and not b;
    layer3_outputs(4973) <= not b;
    layer3_outputs(4974) <= a;
    layer3_outputs(4975) <= not (a or b);
    layer3_outputs(4976) <= b;
    layer3_outputs(4977) <= b and not a;
    layer3_outputs(4978) <= a and b;
    layer3_outputs(4979) <= not a;
    layer3_outputs(4980) <= b and not a;
    layer3_outputs(4981) <= not (a or b);
    layer3_outputs(4982) <= '1';
    layer3_outputs(4983) <= not b or a;
    layer3_outputs(4984) <= not b or a;
    layer3_outputs(4985) <= b;
    layer3_outputs(4986) <= not b;
    layer3_outputs(4987) <= not a;
    layer3_outputs(4988) <= a and b;
    layer3_outputs(4989) <= not a;
    layer3_outputs(4990) <= '0';
    layer3_outputs(4991) <= not b;
    layer3_outputs(4992) <= '1';
    layer3_outputs(4993) <= a;
    layer3_outputs(4994) <= a xor b;
    layer3_outputs(4995) <= a xor b;
    layer3_outputs(4996) <= a;
    layer3_outputs(4997) <= not a or b;
    layer3_outputs(4998) <= not b or a;
    layer3_outputs(4999) <= a and not b;
    layer3_outputs(5000) <= a;
    layer3_outputs(5001) <= a and b;
    layer3_outputs(5002) <= not (a or b);
    layer3_outputs(5003) <= a or b;
    layer3_outputs(5004) <= not (a xor b);
    layer3_outputs(5005) <= '1';
    layer3_outputs(5006) <= a and not b;
    layer3_outputs(5007) <= a or b;
    layer3_outputs(5008) <= not (a or b);
    layer3_outputs(5009) <= b;
    layer3_outputs(5010) <= a and b;
    layer3_outputs(5011) <= not (a and b);
    layer3_outputs(5012) <= a and b;
    layer3_outputs(5013) <= not a or b;
    layer3_outputs(5014) <= not b or a;
    layer3_outputs(5015) <= not b;
    layer3_outputs(5016) <= b;
    layer3_outputs(5017) <= '0';
    layer3_outputs(5018) <= '0';
    layer3_outputs(5019) <= not b;
    layer3_outputs(5020) <= not a;
    layer3_outputs(5021) <= '1';
    layer3_outputs(5022) <= not a or b;
    layer3_outputs(5023) <= '1';
    layer3_outputs(5024) <= not (a and b);
    layer3_outputs(5025) <= not b;
    layer3_outputs(5026) <= not a;
    layer3_outputs(5027) <= a and not b;
    layer3_outputs(5028) <= a and not b;
    layer3_outputs(5029) <= not b or a;
    layer3_outputs(5030) <= not (a and b);
    layer3_outputs(5031) <= '1';
    layer3_outputs(5032) <= b and not a;
    layer3_outputs(5033) <= not a or b;
    layer3_outputs(5034) <= not (a and b);
    layer3_outputs(5035) <= a and not b;
    layer3_outputs(5036) <= not b or a;
    layer3_outputs(5037) <= not b or a;
    layer3_outputs(5038) <= a and b;
    layer3_outputs(5039) <= '1';
    layer3_outputs(5040) <= a;
    layer3_outputs(5041) <= not b;
    layer3_outputs(5042) <= a;
    layer3_outputs(5043) <= b;
    layer3_outputs(5044) <= not a or b;
    layer3_outputs(5045) <= not b;
    layer3_outputs(5046) <= not (a or b);
    layer3_outputs(5047) <= '0';
    layer3_outputs(5048) <= '1';
    layer3_outputs(5049) <= not b or a;
    layer3_outputs(5050) <= not a;
    layer3_outputs(5051) <= b and not a;
    layer3_outputs(5052) <= '0';
    layer3_outputs(5053) <= '1';
    layer3_outputs(5054) <= not (a or b);
    layer3_outputs(5055) <= '1';
    layer3_outputs(5056) <= not a or b;
    layer3_outputs(5057) <= '1';
    layer3_outputs(5058) <= a and not b;
    layer3_outputs(5059) <= '1';
    layer3_outputs(5060) <= '0';
    layer3_outputs(5061) <= b;
    layer3_outputs(5062) <= a and not b;
    layer3_outputs(5063) <= '0';
    layer3_outputs(5064) <= not a;
    layer3_outputs(5065) <= not (a or b);
    layer3_outputs(5066) <= not b;
    layer3_outputs(5067) <= not a or b;
    layer3_outputs(5068) <= b;
    layer3_outputs(5069) <= a and not b;
    layer3_outputs(5070) <= not b;
    layer3_outputs(5071) <= not (a and b);
    layer3_outputs(5072) <= not b or a;
    layer3_outputs(5073) <= '1';
    layer3_outputs(5074) <= not b or a;
    layer3_outputs(5075) <= not b or a;
    layer3_outputs(5076) <= not (a xor b);
    layer3_outputs(5077) <= a and b;
    layer3_outputs(5078) <= a;
    layer3_outputs(5079) <= not b or a;
    layer3_outputs(5080) <= a and not b;
    layer3_outputs(5081) <= not (a xor b);
    layer3_outputs(5082) <= a;
    layer3_outputs(5083) <= '1';
    layer3_outputs(5084) <= not (a and b);
    layer3_outputs(5085) <= not b or a;
    layer3_outputs(5086) <= a xor b;
    layer3_outputs(5087) <= a;
    layer3_outputs(5088) <= a xor b;
    layer3_outputs(5089) <= a and not b;
    layer3_outputs(5090) <= a and not b;
    layer3_outputs(5091) <= b and not a;
    layer3_outputs(5092) <= not (a xor b);
    layer3_outputs(5093) <= b and not a;
    layer3_outputs(5094) <= not b;
    layer3_outputs(5095) <= a;
    layer3_outputs(5096) <= '0';
    layer3_outputs(5097) <= b;
    layer3_outputs(5098) <= a;
    layer3_outputs(5099) <= b and not a;
    layer3_outputs(5100) <= b and not a;
    layer3_outputs(5101) <= '1';
    layer3_outputs(5102) <= '1';
    layer3_outputs(5103) <= not a;
    layer3_outputs(5104) <= b;
    layer3_outputs(5105) <= '1';
    layer3_outputs(5106) <= a or b;
    layer3_outputs(5107) <= '0';
    layer3_outputs(5108) <= '1';
    layer3_outputs(5109) <= a and not b;
    layer3_outputs(5110) <= not (a or b);
    layer3_outputs(5111) <= b and not a;
    layer3_outputs(5112) <= a;
    layer3_outputs(5113) <= '0';
    layer3_outputs(5114) <= not b;
    layer3_outputs(5115) <= not (a or b);
    layer3_outputs(5116) <= a and b;
    layer3_outputs(5117) <= b and not a;
    layer3_outputs(5118) <= a and not b;
    layer3_outputs(5119) <= not a;
    layer4_outputs(0) <= '1';
    layer4_outputs(1) <= not (a or b);
    layer4_outputs(2) <= a or b;
    layer4_outputs(3) <= '1';
    layer4_outputs(4) <= a or b;
    layer4_outputs(5) <= not a;
    layer4_outputs(6) <= not a;
    layer4_outputs(7) <= '1';
    layer4_outputs(8) <= '0';
    layer4_outputs(9) <= b;
    layer4_outputs(10) <= a;
    layer4_outputs(11) <= '0';
    layer4_outputs(12) <= not b;
    layer4_outputs(13) <= a or b;
    layer4_outputs(14) <= a;
    layer4_outputs(15) <= a and not b;
    layer4_outputs(16) <= not b or a;
    layer4_outputs(17) <= a and b;
    layer4_outputs(18) <= not a or b;
    layer4_outputs(19) <= not a or b;
    layer4_outputs(20) <= not (a xor b);
    layer4_outputs(21) <= not (a or b);
    layer4_outputs(22) <= b;
    layer4_outputs(23) <= not (a and b);
    layer4_outputs(24) <= '1';
    layer4_outputs(25) <= not a;
    layer4_outputs(26) <= '0';
    layer4_outputs(27) <= '1';
    layer4_outputs(28) <= a;
    layer4_outputs(29) <= not a or b;
    layer4_outputs(30) <= not (a or b);
    layer4_outputs(31) <= a xor b;
    layer4_outputs(32) <= not b;
    layer4_outputs(33) <= a xor b;
    layer4_outputs(34) <= b;
    layer4_outputs(35) <= not (a and b);
    layer4_outputs(36) <= a and b;
    layer4_outputs(37) <= b and not a;
    layer4_outputs(38) <= not b;
    layer4_outputs(39) <= a and b;
    layer4_outputs(40) <= '0';
    layer4_outputs(41) <= a and b;
    layer4_outputs(42) <= b and not a;
    layer4_outputs(43) <= b;
    layer4_outputs(44) <= '1';
    layer4_outputs(45) <= a and b;
    layer4_outputs(46) <= a;
    layer4_outputs(47) <= a;
    layer4_outputs(48) <= not a;
    layer4_outputs(49) <= '1';
    layer4_outputs(50) <= a;
    layer4_outputs(51) <= not a or b;
    layer4_outputs(52) <= b and not a;
    layer4_outputs(53) <= not (a or b);
    layer4_outputs(54) <= not a or b;
    layer4_outputs(55) <= a xor b;
    layer4_outputs(56) <= not b or a;
    layer4_outputs(57) <= b and not a;
    layer4_outputs(58) <= '0';
    layer4_outputs(59) <= not b;
    layer4_outputs(60) <= '0';
    layer4_outputs(61) <= b;
    layer4_outputs(62) <= not (a or b);
    layer4_outputs(63) <= not a;
    layer4_outputs(64) <= '1';
    layer4_outputs(65) <= a;
    layer4_outputs(66) <= not a or b;
    layer4_outputs(67) <= not b or a;
    layer4_outputs(68) <= b and not a;
    layer4_outputs(69) <= a and not b;
    layer4_outputs(70) <= not (a or b);
    layer4_outputs(71) <= '1';
    layer4_outputs(72) <= a;
    layer4_outputs(73) <= b;
    layer4_outputs(74) <= not b or a;
    layer4_outputs(75) <= not a;
    layer4_outputs(76) <= a or b;
    layer4_outputs(77) <= '1';
    layer4_outputs(78) <= not b;
    layer4_outputs(79) <= a and not b;
    layer4_outputs(80) <= '1';
    layer4_outputs(81) <= a and not b;
    layer4_outputs(82) <= a and not b;
    layer4_outputs(83) <= a and not b;
    layer4_outputs(84) <= not (a and b);
    layer4_outputs(85) <= '1';
    layer4_outputs(86) <= a or b;
    layer4_outputs(87) <= a;
    layer4_outputs(88) <= a or b;
    layer4_outputs(89) <= not (a xor b);
    layer4_outputs(90) <= not b;
    layer4_outputs(91) <= '1';
    layer4_outputs(92) <= a and b;
    layer4_outputs(93) <= not (a and b);
    layer4_outputs(94) <= '1';
    layer4_outputs(95) <= not (a or b);
    layer4_outputs(96) <= not b;
    layer4_outputs(97) <= not b or a;
    layer4_outputs(98) <= a;
    layer4_outputs(99) <= a;
    layer4_outputs(100) <= a and not b;
    layer4_outputs(101) <= a and b;
    layer4_outputs(102) <= not (a or b);
    layer4_outputs(103) <= not b;
    layer4_outputs(104) <= not (a and b);
    layer4_outputs(105) <= a;
    layer4_outputs(106) <= '1';
    layer4_outputs(107) <= '1';
    layer4_outputs(108) <= not (a or b);
    layer4_outputs(109) <= not (a and b);
    layer4_outputs(110) <= not (a or b);
    layer4_outputs(111) <= '1';
    layer4_outputs(112) <= not (a or b);
    layer4_outputs(113) <= b;
    layer4_outputs(114) <= not b or a;
    layer4_outputs(115) <= a;
    layer4_outputs(116) <= a;
    layer4_outputs(117) <= a and not b;
    layer4_outputs(118) <= '0';
    layer4_outputs(119) <= a and b;
    layer4_outputs(120) <= not a;
    layer4_outputs(121) <= a and not b;
    layer4_outputs(122) <= a;
    layer4_outputs(123) <= not b;
    layer4_outputs(124) <= not (a and b);
    layer4_outputs(125) <= a and not b;
    layer4_outputs(126) <= b;
    layer4_outputs(127) <= not b;
    layer4_outputs(128) <= a and not b;
    layer4_outputs(129) <= a or b;
    layer4_outputs(130) <= a;
    layer4_outputs(131) <= not (a or b);
    layer4_outputs(132) <= a;
    layer4_outputs(133) <= '1';
    layer4_outputs(134) <= not (a and b);
    layer4_outputs(135) <= a;
    layer4_outputs(136) <= b and not a;
    layer4_outputs(137) <= not a or b;
    layer4_outputs(138) <= '1';
    layer4_outputs(139) <= not b;
    layer4_outputs(140) <= a and not b;
    layer4_outputs(141) <= '0';
    layer4_outputs(142) <= b and not a;
    layer4_outputs(143) <= '1';
    layer4_outputs(144) <= not a or b;
    layer4_outputs(145) <= not b;
    layer4_outputs(146) <= '1';
    layer4_outputs(147) <= '0';
    layer4_outputs(148) <= a or b;
    layer4_outputs(149) <= a and b;
    layer4_outputs(150) <= b and not a;
    layer4_outputs(151) <= not a;
    layer4_outputs(152) <= not (a or b);
    layer4_outputs(153) <= '1';
    layer4_outputs(154) <= b and not a;
    layer4_outputs(155) <= a xor b;
    layer4_outputs(156) <= not a;
    layer4_outputs(157) <= a and not b;
    layer4_outputs(158) <= a;
    layer4_outputs(159) <= not a;
    layer4_outputs(160) <= not (a and b);
    layer4_outputs(161) <= not b;
    layer4_outputs(162) <= not b;
    layer4_outputs(163) <= not a or b;
    layer4_outputs(164) <= b;
    layer4_outputs(165) <= b;
    layer4_outputs(166) <= b and not a;
    layer4_outputs(167) <= a xor b;
    layer4_outputs(168) <= not a or b;
    layer4_outputs(169) <= b;
    layer4_outputs(170) <= b;
    layer4_outputs(171) <= '1';
    layer4_outputs(172) <= '0';
    layer4_outputs(173) <= b and not a;
    layer4_outputs(174) <= b;
    layer4_outputs(175) <= not a or b;
    layer4_outputs(176) <= not (a or b);
    layer4_outputs(177) <= '0';
    layer4_outputs(178) <= a;
    layer4_outputs(179) <= not a or b;
    layer4_outputs(180) <= not (a or b);
    layer4_outputs(181) <= a and b;
    layer4_outputs(182) <= not b;
    layer4_outputs(183) <= a and b;
    layer4_outputs(184) <= not b or a;
    layer4_outputs(185) <= '0';
    layer4_outputs(186) <= a and b;
    layer4_outputs(187) <= '1';
    layer4_outputs(188) <= a;
    layer4_outputs(189) <= not b;
    layer4_outputs(190) <= b and not a;
    layer4_outputs(191) <= b and not a;
    layer4_outputs(192) <= not a or b;
    layer4_outputs(193) <= a and b;
    layer4_outputs(194) <= not b or a;
    layer4_outputs(195) <= not a or b;
    layer4_outputs(196) <= a and not b;
    layer4_outputs(197) <= '0';
    layer4_outputs(198) <= b;
    layer4_outputs(199) <= not a;
    layer4_outputs(200) <= a and not b;
    layer4_outputs(201) <= b and not a;
    layer4_outputs(202) <= a or b;
    layer4_outputs(203) <= '0';
    layer4_outputs(204) <= a or b;
    layer4_outputs(205) <= not b;
    layer4_outputs(206) <= not (a and b);
    layer4_outputs(207) <= not b;
    layer4_outputs(208) <= a and not b;
    layer4_outputs(209) <= '1';
    layer4_outputs(210) <= not a or b;
    layer4_outputs(211) <= b;
    layer4_outputs(212) <= not b;
    layer4_outputs(213) <= not b or a;
    layer4_outputs(214) <= not a or b;
    layer4_outputs(215) <= not b;
    layer4_outputs(216) <= '0';
    layer4_outputs(217) <= b;
    layer4_outputs(218) <= a and not b;
    layer4_outputs(219) <= not (a and b);
    layer4_outputs(220) <= '1';
    layer4_outputs(221) <= not b or a;
    layer4_outputs(222) <= a or b;
    layer4_outputs(223) <= a and not b;
    layer4_outputs(224) <= not (a and b);
    layer4_outputs(225) <= not b or a;
    layer4_outputs(226) <= a and b;
    layer4_outputs(227) <= not b;
    layer4_outputs(228) <= not (a and b);
    layer4_outputs(229) <= '1';
    layer4_outputs(230) <= not a or b;
    layer4_outputs(231) <= a or b;
    layer4_outputs(232) <= not (a and b);
    layer4_outputs(233) <= b;
    layer4_outputs(234) <= a;
    layer4_outputs(235) <= not a;
    layer4_outputs(236) <= not (a and b);
    layer4_outputs(237) <= b and not a;
    layer4_outputs(238) <= b;
    layer4_outputs(239) <= not b;
    layer4_outputs(240) <= not b;
    layer4_outputs(241) <= not b;
    layer4_outputs(242) <= not (a or b);
    layer4_outputs(243) <= a and not b;
    layer4_outputs(244) <= a or b;
    layer4_outputs(245) <= a or b;
    layer4_outputs(246) <= not (a or b);
    layer4_outputs(247) <= a;
    layer4_outputs(248) <= not (a or b);
    layer4_outputs(249) <= a and b;
    layer4_outputs(250) <= a;
    layer4_outputs(251) <= not (a or b);
    layer4_outputs(252) <= b;
    layer4_outputs(253) <= b;
    layer4_outputs(254) <= not (a and b);
    layer4_outputs(255) <= a and not b;
    layer4_outputs(256) <= not (a xor b);
    layer4_outputs(257) <= not b;
    layer4_outputs(258) <= b and not a;
    layer4_outputs(259) <= not a or b;
    layer4_outputs(260) <= not a;
    layer4_outputs(261) <= b and not a;
    layer4_outputs(262) <= a;
    layer4_outputs(263) <= not a or b;
    layer4_outputs(264) <= a and b;
    layer4_outputs(265) <= '0';
    layer4_outputs(266) <= not a or b;
    layer4_outputs(267) <= '0';
    layer4_outputs(268) <= b;
    layer4_outputs(269) <= b;
    layer4_outputs(270) <= not b or a;
    layer4_outputs(271) <= not a;
    layer4_outputs(272) <= not (a and b);
    layer4_outputs(273) <= not a or b;
    layer4_outputs(274) <= b and not a;
    layer4_outputs(275) <= b and not a;
    layer4_outputs(276) <= not a or b;
    layer4_outputs(277) <= not a;
    layer4_outputs(278) <= a xor b;
    layer4_outputs(279) <= not a;
    layer4_outputs(280) <= a;
    layer4_outputs(281) <= b;
    layer4_outputs(282) <= not b;
    layer4_outputs(283) <= a and b;
    layer4_outputs(284) <= not b or a;
    layer4_outputs(285) <= not a;
    layer4_outputs(286) <= not (a or b);
    layer4_outputs(287) <= b and not a;
    layer4_outputs(288) <= a or b;
    layer4_outputs(289) <= b;
    layer4_outputs(290) <= a or b;
    layer4_outputs(291) <= not a or b;
    layer4_outputs(292) <= not a or b;
    layer4_outputs(293) <= '0';
    layer4_outputs(294) <= not a;
    layer4_outputs(295) <= b and not a;
    layer4_outputs(296) <= a and not b;
    layer4_outputs(297) <= '0';
    layer4_outputs(298) <= not (a and b);
    layer4_outputs(299) <= a or b;
    layer4_outputs(300) <= not a or b;
    layer4_outputs(301) <= b;
    layer4_outputs(302) <= not (a and b);
    layer4_outputs(303) <= a xor b;
    layer4_outputs(304) <= not a;
    layer4_outputs(305) <= not b;
    layer4_outputs(306) <= not (a and b);
    layer4_outputs(307) <= not (a xor b);
    layer4_outputs(308) <= not a;
    layer4_outputs(309) <= not (a and b);
    layer4_outputs(310) <= a xor b;
    layer4_outputs(311) <= '1';
    layer4_outputs(312) <= not a;
    layer4_outputs(313) <= a;
    layer4_outputs(314) <= not (a xor b);
    layer4_outputs(315) <= not b;
    layer4_outputs(316) <= '0';
    layer4_outputs(317) <= a and b;
    layer4_outputs(318) <= '0';
    layer4_outputs(319) <= not b or a;
    layer4_outputs(320) <= b and not a;
    layer4_outputs(321) <= a and not b;
    layer4_outputs(322) <= a and not b;
    layer4_outputs(323) <= a;
    layer4_outputs(324) <= '1';
    layer4_outputs(325) <= a xor b;
    layer4_outputs(326) <= not b;
    layer4_outputs(327) <= not a or b;
    layer4_outputs(328) <= not (a and b);
    layer4_outputs(329) <= not (a and b);
    layer4_outputs(330) <= not (a or b);
    layer4_outputs(331) <= a xor b;
    layer4_outputs(332) <= b and not a;
    layer4_outputs(333) <= not a;
    layer4_outputs(334) <= '0';
    layer4_outputs(335) <= b;
    layer4_outputs(336) <= '0';
    layer4_outputs(337) <= a and b;
    layer4_outputs(338) <= a and not b;
    layer4_outputs(339) <= not a;
    layer4_outputs(340) <= not (a and b);
    layer4_outputs(341) <= a and not b;
    layer4_outputs(342) <= not (a and b);
    layer4_outputs(343) <= '1';
    layer4_outputs(344) <= a;
    layer4_outputs(345) <= not (a or b);
    layer4_outputs(346) <= a or b;
    layer4_outputs(347) <= not b;
    layer4_outputs(348) <= not (a or b);
    layer4_outputs(349) <= b and not a;
    layer4_outputs(350) <= b;
    layer4_outputs(351) <= not a;
    layer4_outputs(352) <= not b or a;
    layer4_outputs(353) <= b;
    layer4_outputs(354) <= a and not b;
    layer4_outputs(355) <= a and not b;
    layer4_outputs(356) <= b;
    layer4_outputs(357) <= a and b;
    layer4_outputs(358) <= a and not b;
    layer4_outputs(359) <= not a or b;
    layer4_outputs(360) <= b and not a;
    layer4_outputs(361) <= not a;
    layer4_outputs(362) <= a and not b;
    layer4_outputs(363) <= not (a and b);
    layer4_outputs(364) <= not a;
    layer4_outputs(365) <= not a;
    layer4_outputs(366) <= a and not b;
    layer4_outputs(367) <= not (a xor b);
    layer4_outputs(368) <= a and b;
    layer4_outputs(369) <= a or b;
    layer4_outputs(370) <= not b;
    layer4_outputs(371) <= a;
    layer4_outputs(372) <= not (a xor b);
    layer4_outputs(373) <= '0';
    layer4_outputs(374) <= a or b;
    layer4_outputs(375) <= a and not b;
    layer4_outputs(376) <= not b or a;
    layer4_outputs(377) <= a and b;
    layer4_outputs(378) <= not a;
    layer4_outputs(379) <= not b;
    layer4_outputs(380) <= not b;
    layer4_outputs(381) <= a and b;
    layer4_outputs(382) <= not a;
    layer4_outputs(383) <= a or b;
    layer4_outputs(384) <= not b;
    layer4_outputs(385) <= '1';
    layer4_outputs(386) <= a and not b;
    layer4_outputs(387) <= a or b;
    layer4_outputs(388) <= b and not a;
    layer4_outputs(389) <= not b;
    layer4_outputs(390) <= not b;
    layer4_outputs(391) <= a and b;
    layer4_outputs(392) <= b and not a;
    layer4_outputs(393) <= '0';
    layer4_outputs(394) <= a or b;
    layer4_outputs(395) <= b and not a;
    layer4_outputs(396) <= a and not b;
    layer4_outputs(397) <= a;
    layer4_outputs(398) <= a and not b;
    layer4_outputs(399) <= a;
    layer4_outputs(400) <= a and b;
    layer4_outputs(401) <= not b;
    layer4_outputs(402) <= a or b;
    layer4_outputs(403) <= a and b;
    layer4_outputs(404) <= b and not a;
    layer4_outputs(405) <= a and b;
    layer4_outputs(406) <= not (a xor b);
    layer4_outputs(407) <= not a;
    layer4_outputs(408) <= a xor b;
    layer4_outputs(409) <= a and not b;
    layer4_outputs(410) <= '0';
    layer4_outputs(411) <= b;
    layer4_outputs(412) <= '1';
    layer4_outputs(413) <= b and not a;
    layer4_outputs(414) <= a and b;
    layer4_outputs(415) <= b and not a;
    layer4_outputs(416) <= '1';
    layer4_outputs(417) <= a or b;
    layer4_outputs(418) <= a;
    layer4_outputs(419) <= a or b;
    layer4_outputs(420) <= a or b;
    layer4_outputs(421) <= not (a or b);
    layer4_outputs(422) <= not (a or b);
    layer4_outputs(423) <= not b;
    layer4_outputs(424) <= not (a and b);
    layer4_outputs(425) <= not b or a;
    layer4_outputs(426) <= b;
    layer4_outputs(427) <= b and not a;
    layer4_outputs(428) <= a;
    layer4_outputs(429) <= a and b;
    layer4_outputs(430) <= b and not a;
    layer4_outputs(431) <= '0';
    layer4_outputs(432) <= not a;
    layer4_outputs(433) <= a and not b;
    layer4_outputs(434) <= b;
    layer4_outputs(435) <= '1';
    layer4_outputs(436) <= a or b;
    layer4_outputs(437) <= a or b;
    layer4_outputs(438) <= b and not a;
    layer4_outputs(439) <= not b or a;
    layer4_outputs(440) <= a;
    layer4_outputs(441) <= not a or b;
    layer4_outputs(442) <= not b or a;
    layer4_outputs(443) <= a;
    layer4_outputs(444) <= '1';
    layer4_outputs(445) <= not (a or b);
    layer4_outputs(446) <= a or b;
    layer4_outputs(447) <= not a;
    layer4_outputs(448) <= not b;
    layer4_outputs(449) <= b;
    layer4_outputs(450) <= a and not b;
    layer4_outputs(451) <= a;
    layer4_outputs(452) <= not b;
    layer4_outputs(453) <= '1';
    layer4_outputs(454) <= b and not a;
    layer4_outputs(455) <= a and b;
    layer4_outputs(456) <= not a or b;
    layer4_outputs(457) <= not a or b;
    layer4_outputs(458) <= a or b;
    layer4_outputs(459) <= '0';
    layer4_outputs(460) <= a and b;
    layer4_outputs(461) <= a and b;
    layer4_outputs(462) <= not (a or b);
    layer4_outputs(463) <= not a or b;
    layer4_outputs(464) <= not b;
    layer4_outputs(465) <= not a or b;
    layer4_outputs(466) <= '0';
    layer4_outputs(467) <= not b or a;
    layer4_outputs(468) <= not b or a;
    layer4_outputs(469) <= not b;
    layer4_outputs(470) <= not b;
    layer4_outputs(471) <= not (a or b);
    layer4_outputs(472) <= a xor b;
    layer4_outputs(473) <= a and not b;
    layer4_outputs(474) <= not a;
    layer4_outputs(475) <= not a;
    layer4_outputs(476) <= not a or b;
    layer4_outputs(477) <= a and b;
    layer4_outputs(478) <= a xor b;
    layer4_outputs(479) <= b and not a;
    layer4_outputs(480) <= not b or a;
    layer4_outputs(481) <= not a;
    layer4_outputs(482) <= b;
    layer4_outputs(483) <= a and b;
    layer4_outputs(484) <= not (a or b);
    layer4_outputs(485) <= not (a or b);
    layer4_outputs(486) <= not b or a;
    layer4_outputs(487) <= b and not a;
    layer4_outputs(488) <= not b;
    layer4_outputs(489) <= a and not b;
    layer4_outputs(490) <= '0';
    layer4_outputs(491) <= not a;
    layer4_outputs(492) <= b and not a;
    layer4_outputs(493) <= a and b;
    layer4_outputs(494) <= not a or b;
    layer4_outputs(495) <= a or b;
    layer4_outputs(496) <= '1';
    layer4_outputs(497) <= b;
    layer4_outputs(498) <= '1';
    layer4_outputs(499) <= '0';
    layer4_outputs(500) <= not (a and b);
    layer4_outputs(501) <= not b;
    layer4_outputs(502) <= b;
    layer4_outputs(503) <= a xor b;
    layer4_outputs(504) <= not (a xor b);
    layer4_outputs(505) <= a or b;
    layer4_outputs(506) <= '0';
    layer4_outputs(507) <= a and not b;
    layer4_outputs(508) <= '0';
    layer4_outputs(509) <= '1';
    layer4_outputs(510) <= not a;
    layer4_outputs(511) <= not b or a;
    layer4_outputs(512) <= a;
    layer4_outputs(513) <= not (a and b);
    layer4_outputs(514) <= a and not b;
    layer4_outputs(515) <= a and b;
    layer4_outputs(516) <= '0';
    layer4_outputs(517) <= '1';
    layer4_outputs(518) <= not b or a;
    layer4_outputs(519) <= b and not a;
    layer4_outputs(520) <= not a or b;
    layer4_outputs(521) <= b and not a;
    layer4_outputs(522) <= a;
    layer4_outputs(523) <= '1';
    layer4_outputs(524) <= not a;
    layer4_outputs(525) <= not (a and b);
    layer4_outputs(526) <= not a or b;
    layer4_outputs(527) <= not (a and b);
    layer4_outputs(528) <= not b;
    layer4_outputs(529) <= not b or a;
    layer4_outputs(530) <= '1';
    layer4_outputs(531) <= not (a xor b);
    layer4_outputs(532) <= not a or b;
    layer4_outputs(533) <= a xor b;
    layer4_outputs(534) <= b;
    layer4_outputs(535) <= not b;
    layer4_outputs(536) <= not (a and b);
    layer4_outputs(537) <= not b;
    layer4_outputs(538) <= a;
    layer4_outputs(539) <= a and not b;
    layer4_outputs(540) <= not b or a;
    layer4_outputs(541) <= not a;
    layer4_outputs(542) <= not a or b;
    layer4_outputs(543) <= b;
    layer4_outputs(544) <= not a;
    layer4_outputs(545) <= b and not a;
    layer4_outputs(546) <= a and not b;
    layer4_outputs(547) <= b and not a;
    layer4_outputs(548) <= not b;
    layer4_outputs(549) <= not b;
    layer4_outputs(550) <= a or b;
    layer4_outputs(551) <= a and b;
    layer4_outputs(552) <= not (a or b);
    layer4_outputs(553) <= a and b;
    layer4_outputs(554) <= a;
    layer4_outputs(555) <= not (a or b);
    layer4_outputs(556) <= a;
    layer4_outputs(557) <= not a;
    layer4_outputs(558) <= a or b;
    layer4_outputs(559) <= a;
    layer4_outputs(560) <= a and b;
    layer4_outputs(561) <= not a or b;
    layer4_outputs(562) <= b;
    layer4_outputs(563) <= not (a and b);
    layer4_outputs(564) <= not a;
    layer4_outputs(565) <= '0';
    layer4_outputs(566) <= not (a or b);
    layer4_outputs(567) <= b;
    layer4_outputs(568) <= a or b;
    layer4_outputs(569) <= not b;
    layer4_outputs(570) <= not b or a;
    layer4_outputs(571) <= not a;
    layer4_outputs(572) <= not a;
    layer4_outputs(573) <= '0';
    layer4_outputs(574) <= not a or b;
    layer4_outputs(575) <= a xor b;
    layer4_outputs(576) <= not b or a;
    layer4_outputs(577) <= not (a and b);
    layer4_outputs(578) <= b and not a;
    layer4_outputs(579) <= not (a or b);
    layer4_outputs(580) <= not a or b;
    layer4_outputs(581) <= a and not b;
    layer4_outputs(582) <= '1';
    layer4_outputs(583) <= a or b;
    layer4_outputs(584) <= not b;
    layer4_outputs(585) <= not a or b;
    layer4_outputs(586) <= '1';
    layer4_outputs(587) <= a and not b;
    layer4_outputs(588) <= not a or b;
    layer4_outputs(589) <= '0';
    layer4_outputs(590) <= not (a and b);
    layer4_outputs(591) <= a;
    layer4_outputs(592) <= not b;
    layer4_outputs(593) <= a;
    layer4_outputs(594) <= a and not b;
    layer4_outputs(595) <= not a or b;
    layer4_outputs(596) <= '0';
    layer4_outputs(597) <= a;
    layer4_outputs(598) <= not b or a;
    layer4_outputs(599) <= a and not b;
    layer4_outputs(600) <= b and not a;
    layer4_outputs(601) <= not b or a;
    layer4_outputs(602) <= not a;
    layer4_outputs(603) <= b and not a;
    layer4_outputs(604) <= b and not a;
    layer4_outputs(605) <= b and not a;
    layer4_outputs(606) <= not a or b;
    layer4_outputs(607) <= b;
    layer4_outputs(608) <= not (a xor b);
    layer4_outputs(609) <= '1';
    layer4_outputs(610) <= not a;
    layer4_outputs(611) <= not b or a;
    layer4_outputs(612) <= a;
    layer4_outputs(613) <= a and not b;
    layer4_outputs(614) <= a;
    layer4_outputs(615) <= not a or b;
    layer4_outputs(616) <= not b or a;
    layer4_outputs(617) <= a;
    layer4_outputs(618) <= '0';
    layer4_outputs(619) <= not (a and b);
    layer4_outputs(620) <= not a or b;
    layer4_outputs(621) <= a or b;
    layer4_outputs(622) <= not (a or b);
    layer4_outputs(623) <= a xor b;
    layer4_outputs(624) <= a;
    layer4_outputs(625) <= not b or a;
    layer4_outputs(626) <= b;
    layer4_outputs(627) <= b;
    layer4_outputs(628) <= not a;
    layer4_outputs(629) <= b;
    layer4_outputs(630) <= not (a or b);
    layer4_outputs(631) <= not (a or b);
    layer4_outputs(632) <= '1';
    layer4_outputs(633) <= a and b;
    layer4_outputs(634) <= a xor b;
    layer4_outputs(635) <= b and not a;
    layer4_outputs(636) <= '1';
    layer4_outputs(637) <= a and b;
    layer4_outputs(638) <= not (a or b);
    layer4_outputs(639) <= not a;
    layer4_outputs(640) <= not (a or b);
    layer4_outputs(641) <= not a;
    layer4_outputs(642) <= '0';
    layer4_outputs(643) <= a;
    layer4_outputs(644) <= not (a or b);
    layer4_outputs(645) <= not (a and b);
    layer4_outputs(646) <= not (a or b);
    layer4_outputs(647) <= a or b;
    layer4_outputs(648) <= not (a or b);
    layer4_outputs(649) <= a;
    layer4_outputs(650) <= a or b;
    layer4_outputs(651) <= not a or b;
    layer4_outputs(652) <= a or b;
    layer4_outputs(653) <= not b;
    layer4_outputs(654) <= a;
    layer4_outputs(655) <= a and not b;
    layer4_outputs(656) <= a and b;
    layer4_outputs(657) <= a or b;
    layer4_outputs(658) <= '1';
    layer4_outputs(659) <= not a or b;
    layer4_outputs(660) <= b;
    layer4_outputs(661) <= not a or b;
    layer4_outputs(662) <= not b;
    layer4_outputs(663) <= not a or b;
    layer4_outputs(664) <= '0';
    layer4_outputs(665) <= b and not a;
    layer4_outputs(666) <= a;
    layer4_outputs(667) <= b;
    layer4_outputs(668) <= a and b;
    layer4_outputs(669) <= not b or a;
    layer4_outputs(670) <= a;
    layer4_outputs(671) <= b;
    layer4_outputs(672) <= not a or b;
    layer4_outputs(673) <= '1';
    layer4_outputs(674) <= a;
    layer4_outputs(675) <= not (a xor b);
    layer4_outputs(676) <= not b or a;
    layer4_outputs(677) <= a and not b;
    layer4_outputs(678) <= not b;
    layer4_outputs(679) <= not b or a;
    layer4_outputs(680) <= a and b;
    layer4_outputs(681) <= not b;
    layer4_outputs(682) <= not b;
    layer4_outputs(683) <= a and not b;
    layer4_outputs(684) <= not b or a;
    layer4_outputs(685) <= a;
    layer4_outputs(686) <= not a;
    layer4_outputs(687) <= a xor b;
    layer4_outputs(688) <= not a;
    layer4_outputs(689) <= not (a or b);
    layer4_outputs(690) <= a;
    layer4_outputs(691) <= not b or a;
    layer4_outputs(692) <= not (a or b);
    layer4_outputs(693) <= a and not b;
    layer4_outputs(694) <= a xor b;
    layer4_outputs(695) <= b and not a;
    layer4_outputs(696) <= b and not a;
    layer4_outputs(697) <= '1';
    layer4_outputs(698) <= not b;
    layer4_outputs(699) <= b;
    layer4_outputs(700) <= a;
    layer4_outputs(701) <= a and not b;
    layer4_outputs(702) <= a xor b;
    layer4_outputs(703) <= not b or a;
    layer4_outputs(704) <= b;
    layer4_outputs(705) <= not b or a;
    layer4_outputs(706) <= a or b;
    layer4_outputs(707) <= '0';
    layer4_outputs(708) <= not (a and b);
    layer4_outputs(709) <= a or b;
    layer4_outputs(710) <= '1';
    layer4_outputs(711) <= a or b;
    layer4_outputs(712) <= not b;
    layer4_outputs(713) <= not (a and b);
    layer4_outputs(714) <= not b or a;
    layer4_outputs(715) <= a xor b;
    layer4_outputs(716) <= a and b;
    layer4_outputs(717) <= '1';
    layer4_outputs(718) <= a;
    layer4_outputs(719) <= not (a xor b);
    layer4_outputs(720) <= not b;
    layer4_outputs(721) <= not (a or b);
    layer4_outputs(722) <= b and not a;
    layer4_outputs(723) <= '0';
    layer4_outputs(724) <= a or b;
    layer4_outputs(725) <= a and b;
    layer4_outputs(726) <= a and not b;
    layer4_outputs(727) <= not a;
    layer4_outputs(728) <= a xor b;
    layer4_outputs(729) <= not a;
    layer4_outputs(730) <= not b or a;
    layer4_outputs(731) <= not a or b;
    layer4_outputs(732) <= not (a xor b);
    layer4_outputs(733) <= not a;
    layer4_outputs(734) <= not b or a;
    layer4_outputs(735) <= not b;
    layer4_outputs(736) <= not (a or b);
    layer4_outputs(737) <= a;
    layer4_outputs(738) <= a and not b;
    layer4_outputs(739) <= b;
    layer4_outputs(740) <= not b;
    layer4_outputs(741) <= not (a and b);
    layer4_outputs(742) <= b;
    layer4_outputs(743) <= not (a or b);
    layer4_outputs(744) <= not a or b;
    layer4_outputs(745) <= a and not b;
    layer4_outputs(746) <= a and not b;
    layer4_outputs(747) <= b;
    layer4_outputs(748) <= '0';
    layer4_outputs(749) <= a;
    layer4_outputs(750) <= b;
    layer4_outputs(751) <= '0';
    layer4_outputs(752) <= not a;
    layer4_outputs(753) <= not b;
    layer4_outputs(754) <= not (a and b);
    layer4_outputs(755) <= b and not a;
    layer4_outputs(756) <= not (a and b);
    layer4_outputs(757) <= a and not b;
    layer4_outputs(758) <= a;
    layer4_outputs(759) <= not (a or b);
    layer4_outputs(760) <= a and b;
    layer4_outputs(761) <= not b;
    layer4_outputs(762) <= a;
    layer4_outputs(763) <= a or b;
    layer4_outputs(764) <= b and not a;
    layer4_outputs(765) <= a and not b;
    layer4_outputs(766) <= not b or a;
    layer4_outputs(767) <= b;
    layer4_outputs(768) <= not (a and b);
    layer4_outputs(769) <= not (a or b);
    layer4_outputs(770) <= a and b;
    layer4_outputs(771) <= '0';
    layer4_outputs(772) <= '1';
    layer4_outputs(773) <= a and b;
    layer4_outputs(774) <= not (a or b);
    layer4_outputs(775) <= '0';
    layer4_outputs(776) <= b;
    layer4_outputs(777) <= b;
    layer4_outputs(778) <= '0';
    layer4_outputs(779) <= a and b;
    layer4_outputs(780) <= not b;
    layer4_outputs(781) <= not b;
    layer4_outputs(782) <= not a;
    layer4_outputs(783) <= not (a or b);
    layer4_outputs(784) <= not (a or b);
    layer4_outputs(785) <= not a or b;
    layer4_outputs(786) <= not (a or b);
    layer4_outputs(787) <= not a or b;
    layer4_outputs(788) <= not b;
    layer4_outputs(789) <= '1';
    layer4_outputs(790) <= a and b;
    layer4_outputs(791) <= b;
    layer4_outputs(792) <= a and not b;
    layer4_outputs(793) <= '0';
    layer4_outputs(794) <= a;
    layer4_outputs(795) <= a and not b;
    layer4_outputs(796) <= b and not a;
    layer4_outputs(797) <= '1';
    layer4_outputs(798) <= '1';
    layer4_outputs(799) <= not b;
    layer4_outputs(800) <= b and not a;
    layer4_outputs(801) <= a or b;
    layer4_outputs(802) <= not (a or b);
    layer4_outputs(803) <= a or b;
    layer4_outputs(804) <= not b or a;
    layer4_outputs(805) <= b;
    layer4_outputs(806) <= not a or b;
    layer4_outputs(807) <= '0';
    layer4_outputs(808) <= not b;
    layer4_outputs(809) <= '1';
    layer4_outputs(810) <= a xor b;
    layer4_outputs(811) <= a and not b;
    layer4_outputs(812) <= not (a xor b);
    layer4_outputs(813) <= not a or b;
    layer4_outputs(814) <= '1';
    layer4_outputs(815) <= a or b;
    layer4_outputs(816) <= not b or a;
    layer4_outputs(817) <= a and not b;
    layer4_outputs(818) <= '0';
    layer4_outputs(819) <= not a or b;
    layer4_outputs(820) <= not b;
    layer4_outputs(821) <= a and not b;
    layer4_outputs(822) <= a and b;
    layer4_outputs(823) <= '0';
    layer4_outputs(824) <= not b;
    layer4_outputs(825) <= not b;
    layer4_outputs(826) <= a;
    layer4_outputs(827) <= '0';
    layer4_outputs(828) <= not (a xor b);
    layer4_outputs(829) <= b;
    layer4_outputs(830) <= a and not b;
    layer4_outputs(831) <= not (a or b);
    layer4_outputs(832) <= b;
    layer4_outputs(833) <= not a;
    layer4_outputs(834) <= not b or a;
    layer4_outputs(835) <= a or b;
    layer4_outputs(836) <= a xor b;
    layer4_outputs(837) <= not b;
    layer4_outputs(838) <= b;
    layer4_outputs(839) <= a and not b;
    layer4_outputs(840) <= a and b;
    layer4_outputs(841) <= a xor b;
    layer4_outputs(842) <= not b;
    layer4_outputs(843) <= not b;
    layer4_outputs(844) <= not (a and b);
    layer4_outputs(845) <= not b;
    layer4_outputs(846) <= b;
    layer4_outputs(847) <= a;
    layer4_outputs(848) <= a;
    layer4_outputs(849) <= a and not b;
    layer4_outputs(850) <= a;
    layer4_outputs(851) <= not a;
    layer4_outputs(852) <= not a or b;
    layer4_outputs(853) <= not b or a;
    layer4_outputs(854) <= '0';
    layer4_outputs(855) <= not b or a;
    layer4_outputs(856) <= '0';
    layer4_outputs(857) <= '0';
    layer4_outputs(858) <= not (a or b);
    layer4_outputs(859) <= a and b;
    layer4_outputs(860) <= '1';
    layer4_outputs(861) <= not b;
    layer4_outputs(862) <= not a;
    layer4_outputs(863) <= a and not b;
    layer4_outputs(864) <= a and b;
    layer4_outputs(865) <= not a or b;
    layer4_outputs(866) <= not b;
    layer4_outputs(867) <= b;
    layer4_outputs(868) <= '0';
    layer4_outputs(869) <= b;
    layer4_outputs(870) <= a and b;
    layer4_outputs(871) <= not a or b;
    layer4_outputs(872) <= a or b;
    layer4_outputs(873) <= b;
    layer4_outputs(874) <= not a;
    layer4_outputs(875) <= a and not b;
    layer4_outputs(876) <= a or b;
    layer4_outputs(877) <= a;
    layer4_outputs(878) <= b;
    layer4_outputs(879) <= not a;
    layer4_outputs(880) <= '1';
    layer4_outputs(881) <= a and not b;
    layer4_outputs(882) <= not b;
    layer4_outputs(883) <= a;
    layer4_outputs(884) <= not (a and b);
    layer4_outputs(885) <= not (a xor b);
    layer4_outputs(886) <= a and b;
    layer4_outputs(887) <= a or b;
    layer4_outputs(888) <= '1';
    layer4_outputs(889) <= a;
    layer4_outputs(890) <= not a or b;
    layer4_outputs(891) <= b and not a;
    layer4_outputs(892) <= not (a or b);
    layer4_outputs(893) <= not a;
    layer4_outputs(894) <= b and not a;
    layer4_outputs(895) <= a;
    layer4_outputs(896) <= not (a and b);
    layer4_outputs(897) <= a or b;
    layer4_outputs(898) <= b and not a;
    layer4_outputs(899) <= not a;
    layer4_outputs(900) <= a;
    layer4_outputs(901) <= a or b;
    layer4_outputs(902) <= a;
    layer4_outputs(903) <= a or b;
    layer4_outputs(904) <= not b or a;
    layer4_outputs(905) <= not a;
    layer4_outputs(906) <= b;
    layer4_outputs(907) <= a or b;
    layer4_outputs(908) <= a and b;
    layer4_outputs(909) <= a or b;
    layer4_outputs(910) <= a and b;
    layer4_outputs(911) <= a and not b;
    layer4_outputs(912) <= a;
    layer4_outputs(913) <= not a;
    layer4_outputs(914) <= '0';
    layer4_outputs(915) <= '1';
    layer4_outputs(916) <= a;
    layer4_outputs(917) <= b;
    layer4_outputs(918) <= b;
    layer4_outputs(919) <= '1';
    layer4_outputs(920) <= a or b;
    layer4_outputs(921) <= a;
    layer4_outputs(922) <= a or b;
    layer4_outputs(923) <= b;
    layer4_outputs(924) <= not (a xor b);
    layer4_outputs(925) <= a and not b;
    layer4_outputs(926) <= not a;
    layer4_outputs(927) <= a;
    layer4_outputs(928) <= '0';
    layer4_outputs(929) <= '0';
    layer4_outputs(930) <= not (a or b);
    layer4_outputs(931) <= a;
    layer4_outputs(932) <= a and b;
    layer4_outputs(933) <= a and not b;
    layer4_outputs(934) <= not (a or b);
    layer4_outputs(935) <= a;
    layer4_outputs(936) <= a or b;
    layer4_outputs(937) <= b;
    layer4_outputs(938) <= a;
    layer4_outputs(939) <= not b or a;
    layer4_outputs(940) <= a;
    layer4_outputs(941) <= '1';
    layer4_outputs(942) <= a and not b;
    layer4_outputs(943) <= not (a or b);
    layer4_outputs(944) <= not a;
    layer4_outputs(945) <= a and not b;
    layer4_outputs(946) <= b and not a;
    layer4_outputs(947) <= a or b;
    layer4_outputs(948) <= a;
    layer4_outputs(949) <= a and not b;
    layer4_outputs(950) <= not (a or b);
    layer4_outputs(951) <= a;
    layer4_outputs(952) <= '0';
    layer4_outputs(953) <= not b;
    layer4_outputs(954) <= a;
    layer4_outputs(955) <= b;
    layer4_outputs(956) <= not a;
    layer4_outputs(957) <= not a or b;
    layer4_outputs(958) <= not b or a;
    layer4_outputs(959) <= not (a or b);
    layer4_outputs(960) <= a or b;
    layer4_outputs(961) <= not b or a;
    layer4_outputs(962) <= not a;
    layer4_outputs(963) <= b;
    layer4_outputs(964) <= b;
    layer4_outputs(965) <= '1';
    layer4_outputs(966) <= a or b;
    layer4_outputs(967) <= a or b;
    layer4_outputs(968) <= a and b;
    layer4_outputs(969) <= not (a or b);
    layer4_outputs(970) <= not a;
    layer4_outputs(971) <= a and not b;
    layer4_outputs(972) <= not b or a;
    layer4_outputs(973) <= b and not a;
    layer4_outputs(974) <= '0';
    layer4_outputs(975) <= b and not a;
    layer4_outputs(976) <= a or b;
    layer4_outputs(977) <= '0';
    layer4_outputs(978) <= not a;
    layer4_outputs(979) <= a or b;
    layer4_outputs(980) <= a;
    layer4_outputs(981) <= not (a or b);
    layer4_outputs(982) <= not b;
    layer4_outputs(983) <= not a or b;
    layer4_outputs(984) <= a;
    layer4_outputs(985) <= a and b;
    layer4_outputs(986) <= a;
    layer4_outputs(987) <= '1';
    layer4_outputs(988) <= '1';
    layer4_outputs(989) <= not b;
    layer4_outputs(990) <= '0';
    layer4_outputs(991) <= not (a or b);
    layer4_outputs(992) <= not a or b;
    layer4_outputs(993) <= '0';
    layer4_outputs(994) <= b;
    layer4_outputs(995) <= b and not a;
    layer4_outputs(996) <= '1';
    layer4_outputs(997) <= '1';
    layer4_outputs(998) <= not a or b;
    layer4_outputs(999) <= not (a or b);
    layer4_outputs(1000) <= not a or b;
    layer4_outputs(1001) <= a or b;
    layer4_outputs(1002) <= a or b;
    layer4_outputs(1003) <= not (a and b);
    layer4_outputs(1004) <= a or b;
    layer4_outputs(1005) <= a or b;
    layer4_outputs(1006) <= a and b;
    layer4_outputs(1007) <= '0';
    layer4_outputs(1008) <= not (a xor b);
    layer4_outputs(1009) <= b and not a;
    layer4_outputs(1010) <= a;
    layer4_outputs(1011) <= a or b;
    layer4_outputs(1012) <= not (a and b);
    layer4_outputs(1013) <= a xor b;
    layer4_outputs(1014) <= not (a or b);
    layer4_outputs(1015) <= a;
    layer4_outputs(1016) <= not b or a;
    layer4_outputs(1017) <= a;
    layer4_outputs(1018) <= not b or a;
    layer4_outputs(1019) <= not b or a;
    layer4_outputs(1020) <= a and not b;
    layer4_outputs(1021) <= a and not b;
    layer4_outputs(1022) <= a or b;
    layer4_outputs(1023) <= a;
    layer4_outputs(1024) <= a or b;
    layer4_outputs(1025) <= not (a or b);
    layer4_outputs(1026) <= a and b;
    layer4_outputs(1027) <= a and b;
    layer4_outputs(1028) <= a and b;
    layer4_outputs(1029) <= a or b;
    layer4_outputs(1030) <= not a;
    layer4_outputs(1031) <= '0';
    layer4_outputs(1032) <= '0';
    layer4_outputs(1033) <= not b or a;
    layer4_outputs(1034) <= a;
    layer4_outputs(1035) <= not a or b;
    layer4_outputs(1036) <= '0';
    layer4_outputs(1037) <= b and not a;
    layer4_outputs(1038) <= a or b;
    layer4_outputs(1039) <= a;
    layer4_outputs(1040) <= a and not b;
    layer4_outputs(1041) <= not (a and b);
    layer4_outputs(1042) <= a and b;
    layer4_outputs(1043) <= not (a and b);
    layer4_outputs(1044) <= not (a or b);
    layer4_outputs(1045) <= not b or a;
    layer4_outputs(1046) <= a and not b;
    layer4_outputs(1047) <= a;
    layer4_outputs(1048) <= not a;
    layer4_outputs(1049) <= b and not a;
    layer4_outputs(1050) <= b and not a;
    layer4_outputs(1051) <= not (a and b);
    layer4_outputs(1052) <= not b;
    layer4_outputs(1053) <= '0';
    layer4_outputs(1054) <= not b;
    layer4_outputs(1055) <= a;
    layer4_outputs(1056) <= a and not b;
    layer4_outputs(1057) <= a and not b;
    layer4_outputs(1058) <= a;
    layer4_outputs(1059) <= not a or b;
    layer4_outputs(1060) <= a;
    layer4_outputs(1061) <= a and b;
    layer4_outputs(1062) <= not a or b;
    layer4_outputs(1063) <= not b;
    layer4_outputs(1064) <= not b;
    layer4_outputs(1065) <= b and not a;
    layer4_outputs(1066) <= not a;
    layer4_outputs(1067) <= b and not a;
    layer4_outputs(1068) <= a xor b;
    layer4_outputs(1069) <= a or b;
    layer4_outputs(1070) <= b and not a;
    layer4_outputs(1071) <= not (a and b);
    layer4_outputs(1072) <= b and not a;
    layer4_outputs(1073) <= a and b;
    layer4_outputs(1074) <= b;
    layer4_outputs(1075) <= a;
    layer4_outputs(1076) <= b;
    layer4_outputs(1077) <= '0';
    layer4_outputs(1078) <= not a;
    layer4_outputs(1079) <= a or b;
    layer4_outputs(1080) <= not a;
    layer4_outputs(1081) <= b;
    layer4_outputs(1082) <= b and not a;
    layer4_outputs(1083) <= not b or a;
    layer4_outputs(1084) <= not (a or b);
    layer4_outputs(1085) <= not a;
    layer4_outputs(1086) <= not (a and b);
    layer4_outputs(1087) <= b;
    layer4_outputs(1088) <= a and not b;
    layer4_outputs(1089) <= not b;
    layer4_outputs(1090) <= not b;
    layer4_outputs(1091) <= a;
    layer4_outputs(1092) <= a and not b;
    layer4_outputs(1093) <= b and not a;
    layer4_outputs(1094) <= '1';
    layer4_outputs(1095) <= not b;
    layer4_outputs(1096) <= b and not a;
    layer4_outputs(1097) <= a;
    layer4_outputs(1098) <= '1';
    layer4_outputs(1099) <= a and b;
    layer4_outputs(1100) <= not (a and b);
    layer4_outputs(1101) <= a and not b;
    layer4_outputs(1102) <= not b or a;
    layer4_outputs(1103) <= b;
    layer4_outputs(1104) <= a;
    layer4_outputs(1105) <= a and b;
    layer4_outputs(1106) <= not a or b;
    layer4_outputs(1107) <= a or b;
    layer4_outputs(1108) <= not b or a;
    layer4_outputs(1109) <= not a or b;
    layer4_outputs(1110) <= a and b;
    layer4_outputs(1111) <= not b or a;
    layer4_outputs(1112) <= b;
    layer4_outputs(1113) <= not b or a;
    layer4_outputs(1114) <= a;
    layer4_outputs(1115) <= a and not b;
    layer4_outputs(1116) <= '1';
    layer4_outputs(1117) <= b;
    layer4_outputs(1118) <= '0';
    layer4_outputs(1119) <= not a;
    layer4_outputs(1120) <= a;
    layer4_outputs(1121) <= not a or b;
    layer4_outputs(1122) <= not (a and b);
    layer4_outputs(1123) <= not a;
    layer4_outputs(1124) <= not (a or b);
    layer4_outputs(1125) <= b;
    layer4_outputs(1126) <= b and not a;
    layer4_outputs(1127) <= a and b;
    layer4_outputs(1128) <= '0';
    layer4_outputs(1129) <= '0';
    layer4_outputs(1130) <= not b or a;
    layer4_outputs(1131) <= not b or a;
    layer4_outputs(1132) <= b and not a;
    layer4_outputs(1133) <= a and not b;
    layer4_outputs(1134) <= a and not b;
    layer4_outputs(1135) <= not a;
    layer4_outputs(1136) <= not (a or b);
    layer4_outputs(1137) <= a and not b;
    layer4_outputs(1138) <= not a or b;
    layer4_outputs(1139) <= '1';
    layer4_outputs(1140) <= not (a or b);
    layer4_outputs(1141) <= a;
    layer4_outputs(1142) <= a and not b;
    layer4_outputs(1143) <= b;
    layer4_outputs(1144) <= not a;
    layer4_outputs(1145) <= not a or b;
    layer4_outputs(1146) <= not a or b;
    layer4_outputs(1147) <= a or b;
    layer4_outputs(1148) <= not (a xor b);
    layer4_outputs(1149) <= a;
    layer4_outputs(1150) <= not (a or b);
    layer4_outputs(1151) <= not (a or b);
    layer4_outputs(1152) <= a and b;
    layer4_outputs(1153) <= not a;
    layer4_outputs(1154) <= not (a or b);
    layer4_outputs(1155) <= b;
    layer4_outputs(1156) <= b and not a;
    layer4_outputs(1157) <= a;
    layer4_outputs(1158) <= a and not b;
    layer4_outputs(1159) <= not b or a;
    layer4_outputs(1160) <= b;
    layer4_outputs(1161) <= a or b;
    layer4_outputs(1162) <= a;
    layer4_outputs(1163) <= not a or b;
    layer4_outputs(1164) <= not (a or b);
    layer4_outputs(1165) <= a and b;
    layer4_outputs(1166) <= not (a or b);
    layer4_outputs(1167) <= not (a or b);
    layer4_outputs(1168) <= not b or a;
    layer4_outputs(1169) <= not (a or b);
    layer4_outputs(1170) <= not (a or b);
    layer4_outputs(1171) <= b and not a;
    layer4_outputs(1172) <= '1';
    layer4_outputs(1173) <= b;
    layer4_outputs(1174) <= b;
    layer4_outputs(1175) <= '1';
    layer4_outputs(1176) <= a and b;
    layer4_outputs(1177) <= a and not b;
    layer4_outputs(1178) <= not b;
    layer4_outputs(1179) <= not a or b;
    layer4_outputs(1180) <= not b;
    layer4_outputs(1181) <= not (a or b);
    layer4_outputs(1182) <= not a;
    layer4_outputs(1183) <= a or b;
    layer4_outputs(1184) <= '1';
    layer4_outputs(1185) <= '1';
    layer4_outputs(1186) <= a or b;
    layer4_outputs(1187) <= b and not a;
    layer4_outputs(1188) <= a and not b;
    layer4_outputs(1189) <= a xor b;
    layer4_outputs(1190) <= '0';
    layer4_outputs(1191) <= b and not a;
    layer4_outputs(1192) <= not a;
    layer4_outputs(1193) <= not b;
    layer4_outputs(1194) <= not b;
    layer4_outputs(1195) <= a and b;
    layer4_outputs(1196) <= '1';
    layer4_outputs(1197) <= a and b;
    layer4_outputs(1198) <= not (a and b);
    layer4_outputs(1199) <= a or b;
    layer4_outputs(1200) <= a and not b;
    layer4_outputs(1201) <= a or b;
    layer4_outputs(1202) <= not b;
    layer4_outputs(1203) <= '0';
    layer4_outputs(1204) <= not b or a;
    layer4_outputs(1205) <= not (a and b);
    layer4_outputs(1206) <= not (a or b);
    layer4_outputs(1207) <= not (a xor b);
    layer4_outputs(1208) <= a;
    layer4_outputs(1209) <= a and b;
    layer4_outputs(1210) <= not b;
    layer4_outputs(1211) <= b;
    layer4_outputs(1212) <= a;
    layer4_outputs(1213) <= b;
    layer4_outputs(1214) <= b;
    layer4_outputs(1215) <= a and not b;
    layer4_outputs(1216) <= b;
    layer4_outputs(1217) <= b and not a;
    layer4_outputs(1218) <= not b;
    layer4_outputs(1219) <= a and b;
    layer4_outputs(1220) <= not b or a;
    layer4_outputs(1221) <= a xor b;
    layer4_outputs(1222) <= a;
    layer4_outputs(1223) <= not a or b;
    layer4_outputs(1224) <= a xor b;
    layer4_outputs(1225) <= not a;
    layer4_outputs(1226) <= not (a and b);
    layer4_outputs(1227) <= '0';
    layer4_outputs(1228) <= a and not b;
    layer4_outputs(1229) <= not b;
    layer4_outputs(1230) <= not (a or b);
    layer4_outputs(1231) <= '0';
    layer4_outputs(1232) <= not a or b;
    layer4_outputs(1233) <= a and b;
    layer4_outputs(1234) <= not a or b;
    layer4_outputs(1235) <= not b;
    layer4_outputs(1236) <= '1';
    layer4_outputs(1237) <= not b or a;
    layer4_outputs(1238) <= not (a and b);
    layer4_outputs(1239) <= '1';
    layer4_outputs(1240) <= '1';
    layer4_outputs(1241) <= b;
    layer4_outputs(1242) <= not b;
    layer4_outputs(1243) <= b and not a;
    layer4_outputs(1244) <= a xor b;
    layer4_outputs(1245) <= '0';
    layer4_outputs(1246) <= a xor b;
    layer4_outputs(1247) <= b and not a;
    layer4_outputs(1248) <= not b;
    layer4_outputs(1249) <= not b;
    layer4_outputs(1250) <= a xor b;
    layer4_outputs(1251) <= '0';
    layer4_outputs(1252) <= '1';
    layer4_outputs(1253) <= '1';
    layer4_outputs(1254) <= a or b;
    layer4_outputs(1255) <= a xor b;
    layer4_outputs(1256) <= b and not a;
    layer4_outputs(1257) <= not a or b;
    layer4_outputs(1258) <= not a or b;
    layer4_outputs(1259) <= '0';
    layer4_outputs(1260) <= not (a or b);
    layer4_outputs(1261) <= not a;
    layer4_outputs(1262) <= b;
    layer4_outputs(1263) <= not (a or b);
    layer4_outputs(1264) <= not a;
    layer4_outputs(1265) <= a or b;
    layer4_outputs(1266) <= '0';
    layer4_outputs(1267) <= a and b;
    layer4_outputs(1268) <= not a or b;
    layer4_outputs(1269) <= '0';
    layer4_outputs(1270) <= a and not b;
    layer4_outputs(1271) <= b and not a;
    layer4_outputs(1272) <= '0';
    layer4_outputs(1273) <= not a or b;
    layer4_outputs(1274) <= not (a and b);
    layer4_outputs(1275) <= not (a or b);
    layer4_outputs(1276) <= not (a or b);
    layer4_outputs(1277) <= a and b;
    layer4_outputs(1278) <= not (a or b);
    layer4_outputs(1279) <= not (a and b);
    layer4_outputs(1280) <= not a or b;
    layer4_outputs(1281) <= b;
    layer4_outputs(1282) <= '1';
    layer4_outputs(1283) <= a and b;
    layer4_outputs(1284) <= not b;
    layer4_outputs(1285) <= b and not a;
    layer4_outputs(1286) <= a or b;
    layer4_outputs(1287) <= b;
    layer4_outputs(1288) <= not b;
    layer4_outputs(1289) <= b and not a;
    layer4_outputs(1290) <= a;
    layer4_outputs(1291) <= not b;
    layer4_outputs(1292) <= not a;
    layer4_outputs(1293) <= a xor b;
    layer4_outputs(1294) <= not a;
    layer4_outputs(1295) <= not a;
    layer4_outputs(1296) <= a and b;
    layer4_outputs(1297) <= not b;
    layer4_outputs(1298) <= not (a or b);
    layer4_outputs(1299) <= not (a and b);
    layer4_outputs(1300) <= a and not b;
    layer4_outputs(1301) <= '1';
    layer4_outputs(1302) <= '0';
    layer4_outputs(1303) <= a and not b;
    layer4_outputs(1304) <= not (a or b);
    layer4_outputs(1305) <= b;
    layer4_outputs(1306) <= not (a and b);
    layer4_outputs(1307) <= a or b;
    layer4_outputs(1308) <= not a;
    layer4_outputs(1309) <= a and not b;
    layer4_outputs(1310) <= b and not a;
    layer4_outputs(1311) <= a or b;
    layer4_outputs(1312) <= a or b;
    layer4_outputs(1313) <= b;
    layer4_outputs(1314) <= not a;
    layer4_outputs(1315) <= '0';
    layer4_outputs(1316) <= not (a or b);
    layer4_outputs(1317) <= a and not b;
    layer4_outputs(1318) <= not (a or b);
    layer4_outputs(1319) <= b;
    layer4_outputs(1320) <= b and not a;
    layer4_outputs(1321) <= not a or b;
    layer4_outputs(1322) <= '0';
    layer4_outputs(1323) <= '1';
    layer4_outputs(1324) <= not b;
    layer4_outputs(1325) <= b;
    layer4_outputs(1326) <= a or b;
    layer4_outputs(1327) <= a;
    layer4_outputs(1328) <= not (a xor b);
    layer4_outputs(1329) <= b;
    layer4_outputs(1330) <= not (a or b);
    layer4_outputs(1331) <= a and not b;
    layer4_outputs(1332) <= a;
    layer4_outputs(1333) <= b;
    layer4_outputs(1334) <= '1';
    layer4_outputs(1335) <= not b;
    layer4_outputs(1336) <= a;
    layer4_outputs(1337) <= b and not a;
    layer4_outputs(1338) <= not (a and b);
    layer4_outputs(1339) <= not a;
    layer4_outputs(1340) <= a;
    layer4_outputs(1341) <= '1';
    layer4_outputs(1342) <= not (a or b);
    layer4_outputs(1343) <= '0';
    layer4_outputs(1344) <= a and b;
    layer4_outputs(1345) <= a and not b;
    layer4_outputs(1346) <= '0';
    layer4_outputs(1347) <= b;
    layer4_outputs(1348) <= a xor b;
    layer4_outputs(1349) <= b;
    layer4_outputs(1350) <= not b or a;
    layer4_outputs(1351) <= a;
    layer4_outputs(1352) <= a;
    layer4_outputs(1353) <= not b or a;
    layer4_outputs(1354) <= not (a and b);
    layer4_outputs(1355) <= b;
    layer4_outputs(1356) <= a and not b;
    layer4_outputs(1357) <= not b or a;
    layer4_outputs(1358) <= a;
    layer4_outputs(1359) <= a;
    layer4_outputs(1360) <= a;
    layer4_outputs(1361) <= a and b;
    layer4_outputs(1362) <= a;
    layer4_outputs(1363) <= a or b;
    layer4_outputs(1364) <= not (a and b);
    layer4_outputs(1365) <= b;
    layer4_outputs(1366) <= not b or a;
    layer4_outputs(1367) <= a;
    layer4_outputs(1368) <= not b or a;
    layer4_outputs(1369) <= a;
    layer4_outputs(1370) <= a or b;
    layer4_outputs(1371) <= b and not a;
    layer4_outputs(1372) <= not a or b;
    layer4_outputs(1373) <= '0';
    layer4_outputs(1374) <= a;
    layer4_outputs(1375) <= not (a and b);
    layer4_outputs(1376) <= a and not b;
    layer4_outputs(1377) <= a;
    layer4_outputs(1378) <= b and not a;
    layer4_outputs(1379) <= not b or a;
    layer4_outputs(1380) <= '0';
    layer4_outputs(1381) <= not (a and b);
    layer4_outputs(1382) <= a and b;
    layer4_outputs(1383) <= a;
    layer4_outputs(1384) <= b and not a;
    layer4_outputs(1385) <= a;
    layer4_outputs(1386) <= a and not b;
    layer4_outputs(1387) <= a;
    layer4_outputs(1388) <= not b or a;
    layer4_outputs(1389) <= a or b;
    layer4_outputs(1390) <= not a or b;
    layer4_outputs(1391) <= a and b;
    layer4_outputs(1392) <= a;
    layer4_outputs(1393) <= not b;
    layer4_outputs(1394) <= not (a or b);
    layer4_outputs(1395) <= a;
    layer4_outputs(1396) <= b;
    layer4_outputs(1397) <= a and b;
    layer4_outputs(1398) <= not (a or b);
    layer4_outputs(1399) <= b and not a;
    layer4_outputs(1400) <= not a or b;
    layer4_outputs(1401) <= not (a and b);
    layer4_outputs(1402) <= not (a xor b);
    layer4_outputs(1403) <= not (a or b);
    layer4_outputs(1404) <= not a;
    layer4_outputs(1405) <= not a;
    layer4_outputs(1406) <= a and b;
    layer4_outputs(1407) <= b and not a;
    layer4_outputs(1408) <= not (a and b);
    layer4_outputs(1409) <= not a;
    layer4_outputs(1410) <= not b;
    layer4_outputs(1411) <= not b or a;
    layer4_outputs(1412) <= b and not a;
    layer4_outputs(1413) <= not b or a;
    layer4_outputs(1414) <= a and not b;
    layer4_outputs(1415) <= not a;
    layer4_outputs(1416) <= a or b;
    layer4_outputs(1417) <= a and b;
    layer4_outputs(1418) <= not b;
    layer4_outputs(1419) <= a and not b;
    layer4_outputs(1420) <= a;
    layer4_outputs(1421) <= a or b;
    layer4_outputs(1422) <= b and not a;
    layer4_outputs(1423) <= a xor b;
    layer4_outputs(1424) <= not (a or b);
    layer4_outputs(1425) <= '1';
    layer4_outputs(1426) <= not (a or b);
    layer4_outputs(1427) <= not (a and b);
    layer4_outputs(1428) <= b;
    layer4_outputs(1429) <= not a or b;
    layer4_outputs(1430) <= not (a and b);
    layer4_outputs(1431) <= a or b;
    layer4_outputs(1432) <= a;
    layer4_outputs(1433) <= not a;
    layer4_outputs(1434) <= not a or b;
    layer4_outputs(1435) <= not (a or b);
    layer4_outputs(1436) <= b;
    layer4_outputs(1437) <= b and not a;
    layer4_outputs(1438) <= not b or a;
    layer4_outputs(1439) <= a or b;
    layer4_outputs(1440) <= not a;
    layer4_outputs(1441) <= '1';
    layer4_outputs(1442) <= b;
    layer4_outputs(1443) <= a or b;
    layer4_outputs(1444) <= not (a and b);
    layer4_outputs(1445) <= a;
    layer4_outputs(1446) <= '1';
    layer4_outputs(1447) <= not a or b;
    layer4_outputs(1448) <= not a or b;
    layer4_outputs(1449) <= b;
    layer4_outputs(1450) <= not a;
    layer4_outputs(1451) <= '0';
    layer4_outputs(1452) <= a and b;
    layer4_outputs(1453) <= not a;
    layer4_outputs(1454) <= a xor b;
    layer4_outputs(1455) <= b;
    layer4_outputs(1456) <= not (a xor b);
    layer4_outputs(1457) <= not (a and b);
    layer4_outputs(1458) <= not a or b;
    layer4_outputs(1459) <= not a;
    layer4_outputs(1460) <= a and not b;
    layer4_outputs(1461) <= '1';
    layer4_outputs(1462) <= not b;
    layer4_outputs(1463) <= not a;
    layer4_outputs(1464) <= a and not b;
    layer4_outputs(1465) <= a;
    layer4_outputs(1466) <= a and b;
    layer4_outputs(1467) <= a xor b;
    layer4_outputs(1468) <= not a;
    layer4_outputs(1469) <= a or b;
    layer4_outputs(1470) <= '1';
    layer4_outputs(1471) <= not a or b;
    layer4_outputs(1472) <= a;
    layer4_outputs(1473) <= not (a and b);
    layer4_outputs(1474) <= b and not a;
    layer4_outputs(1475) <= not a;
    layer4_outputs(1476) <= not b;
    layer4_outputs(1477) <= '1';
    layer4_outputs(1478) <= not (a and b);
    layer4_outputs(1479) <= '1';
    layer4_outputs(1480) <= b and not a;
    layer4_outputs(1481) <= b and not a;
    layer4_outputs(1482) <= a xor b;
    layer4_outputs(1483) <= not a;
    layer4_outputs(1484) <= a or b;
    layer4_outputs(1485) <= a and not b;
    layer4_outputs(1486) <= not a or b;
    layer4_outputs(1487) <= not b or a;
    layer4_outputs(1488) <= not b or a;
    layer4_outputs(1489) <= '1';
    layer4_outputs(1490) <= a and b;
    layer4_outputs(1491) <= not a;
    layer4_outputs(1492) <= a;
    layer4_outputs(1493) <= not b;
    layer4_outputs(1494) <= a and b;
    layer4_outputs(1495) <= not (a or b);
    layer4_outputs(1496) <= not a;
    layer4_outputs(1497) <= a and b;
    layer4_outputs(1498) <= not a;
    layer4_outputs(1499) <= not (a or b);
    layer4_outputs(1500) <= not (a or b);
    layer4_outputs(1501) <= a or b;
    layer4_outputs(1502) <= a and b;
    layer4_outputs(1503) <= b and not a;
    layer4_outputs(1504) <= b and not a;
    layer4_outputs(1505) <= b;
    layer4_outputs(1506) <= not (a xor b);
    layer4_outputs(1507) <= '1';
    layer4_outputs(1508) <= '0';
    layer4_outputs(1509) <= not a;
    layer4_outputs(1510) <= a or b;
    layer4_outputs(1511) <= not (a and b);
    layer4_outputs(1512) <= a or b;
    layer4_outputs(1513) <= b and not a;
    layer4_outputs(1514) <= not (a and b);
    layer4_outputs(1515) <= a or b;
    layer4_outputs(1516) <= not b or a;
    layer4_outputs(1517) <= '0';
    layer4_outputs(1518) <= not (a and b);
    layer4_outputs(1519) <= a and not b;
    layer4_outputs(1520) <= a and not b;
    layer4_outputs(1521) <= not (a and b);
    layer4_outputs(1522) <= a or b;
    layer4_outputs(1523) <= not b or a;
    layer4_outputs(1524) <= a and not b;
    layer4_outputs(1525) <= not (a or b);
    layer4_outputs(1526) <= not (a and b);
    layer4_outputs(1527) <= not a or b;
    layer4_outputs(1528) <= b and not a;
    layer4_outputs(1529) <= a and not b;
    layer4_outputs(1530) <= '1';
    layer4_outputs(1531) <= not a or b;
    layer4_outputs(1532) <= b;
    layer4_outputs(1533) <= '1';
    layer4_outputs(1534) <= '1';
    layer4_outputs(1535) <= not (a and b);
    layer4_outputs(1536) <= a and b;
    layer4_outputs(1537) <= not (a or b);
    layer4_outputs(1538) <= b;
    layer4_outputs(1539) <= not b;
    layer4_outputs(1540) <= '1';
    layer4_outputs(1541) <= not (a xor b);
    layer4_outputs(1542) <= a and b;
    layer4_outputs(1543) <= a and b;
    layer4_outputs(1544) <= not (a and b);
    layer4_outputs(1545) <= not a or b;
    layer4_outputs(1546) <= b;
    layer4_outputs(1547) <= '0';
    layer4_outputs(1548) <= not a;
    layer4_outputs(1549) <= not b;
    layer4_outputs(1550) <= a and b;
    layer4_outputs(1551) <= a and b;
    layer4_outputs(1552) <= not (a and b);
    layer4_outputs(1553) <= not b;
    layer4_outputs(1554) <= '0';
    layer4_outputs(1555) <= not b;
    layer4_outputs(1556) <= not a;
    layer4_outputs(1557) <= not (a and b);
    layer4_outputs(1558) <= '0';
    layer4_outputs(1559) <= a and not b;
    layer4_outputs(1560) <= a;
    layer4_outputs(1561) <= not b;
    layer4_outputs(1562) <= not (a and b);
    layer4_outputs(1563) <= not (a xor b);
    layer4_outputs(1564) <= not (a or b);
    layer4_outputs(1565) <= b and not a;
    layer4_outputs(1566) <= b and not a;
    layer4_outputs(1567) <= not b or a;
    layer4_outputs(1568) <= a and b;
    layer4_outputs(1569) <= b and not a;
    layer4_outputs(1570) <= b;
    layer4_outputs(1571) <= not (a or b);
    layer4_outputs(1572) <= not a or b;
    layer4_outputs(1573) <= a or b;
    layer4_outputs(1574) <= b and not a;
    layer4_outputs(1575) <= a;
    layer4_outputs(1576) <= not b;
    layer4_outputs(1577) <= a and b;
    layer4_outputs(1578) <= a and not b;
    layer4_outputs(1579) <= a and not b;
    layer4_outputs(1580) <= not a or b;
    layer4_outputs(1581) <= not (a and b);
    layer4_outputs(1582) <= not (a xor b);
    layer4_outputs(1583) <= not (a or b);
    layer4_outputs(1584) <= not b;
    layer4_outputs(1585) <= '0';
    layer4_outputs(1586) <= '0';
    layer4_outputs(1587) <= not b;
    layer4_outputs(1588) <= b;
    layer4_outputs(1589) <= a and not b;
    layer4_outputs(1590) <= '0';
    layer4_outputs(1591) <= a or b;
    layer4_outputs(1592) <= not a or b;
    layer4_outputs(1593) <= a;
    layer4_outputs(1594) <= not (a and b);
    layer4_outputs(1595) <= a and not b;
    layer4_outputs(1596) <= not b or a;
    layer4_outputs(1597) <= a;
    layer4_outputs(1598) <= a or b;
    layer4_outputs(1599) <= not a;
    layer4_outputs(1600) <= a and not b;
    layer4_outputs(1601) <= b;
    layer4_outputs(1602) <= a and not b;
    layer4_outputs(1603) <= a;
    layer4_outputs(1604) <= a and b;
    layer4_outputs(1605) <= not a;
    layer4_outputs(1606) <= a;
    layer4_outputs(1607) <= not (a and b);
    layer4_outputs(1608) <= not (a or b);
    layer4_outputs(1609) <= a or b;
    layer4_outputs(1610) <= b;
    layer4_outputs(1611) <= a or b;
    layer4_outputs(1612) <= not b;
    layer4_outputs(1613) <= a and not b;
    layer4_outputs(1614) <= a and b;
    layer4_outputs(1615) <= not b;
    layer4_outputs(1616) <= not b or a;
    layer4_outputs(1617) <= not b;
    layer4_outputs(1618) <= not b or a;
    layer4_outputs(1619) <= not a;
    layer4_outputs(1620) <= not a;
    layer4_outputs(1621) <= a or b;
    layer4_outputs(1622) <= not a;
    layer4_outputs(1623) <= '1';
    layer4_outputs(1624) <= b and not a;
    layer4_outputs(1625) <= not b;
    layer4_outputs(1626) <= a;
    layer4_outputs(1627) <= not a or b;
    layer4_outputs(1628) <= a or b;
    layer4_outputs(1629) <= not a;
    layer4_outputs(1630) <= a and b;
    layer4_outputs(1631) <= not (a and b);
    layer4_outputs(1632) <= a and not b;
    layer4_outputs(1633) <= not (a and b);
    layer4_outputs(1634) <= not a;
    layer4_outputs(1635) <= not (a and b);
    layer4_outputs(1636) <= a or b;
    layer4_outputs(1637) <= b and not a;
    layer4_outputs(1638) <= '1';
    layer4_outputs(1639) <= not b;
    layer4_outputs(1640) <= not a;
    layer4_outputs(1641) <= a and b;
    layer4_outputs(1642) <= not b;
    layer4_outputs(1643) <= '0';
    layer4_outputs(1644) <= not b or a;
    layer4_outputs(1645) <= a and not b;
    layer4_outputs(1646) <= b;
    layer4_outputs(1647) <= a;
    layer4_outputs(1648) <= not (a xor b);
    layer4_outputs(1649) <= not a;
    layer4_outputs(1650) <= not (a and b);
    layer4_outputs(1651) <= not a;
    layer4_outputs(1652) <= a;
    layer4_outputs(1653) <= a and b;
    layer4_outputs(1654) <= not b or a;
    layer4_outputs(1655) <= not b;
    layer4_outputs(1656) <= not a or b;
    layer4_outputs(1657) <= not (a and b);
    layer4_outputs(1658) <= a xor b;
    layer4_outputs(1659) <= not b or a;
    layer4_outputs(1660) <= not (a and b);
    layer4_outputs(1661) <= '0';
    layer4_outputs(1662) <= not b;
    layer4_outputs(1663) <= a and not b;
    layer4_outputs(1664) <= not b;
    layer4_outputs(1665) <= not (a or b);
    layer4_outputs(1666) <= a or b;
    layer4_outputs(1667) <= not (a or b);
    layer4_outputs(1668) <= not b;
    layer4_outputs(1669) <= '0';
    layer4_outputs(1670) <= a and b;
    layer4_outputs(1671) <= not (a and b);
    layer4_outputs(1672) <= not (a or b);
    layer4_outputs(1673) <= not b;
    layer4_outputs(1674) <= a;
    layer4_outputs(1675) <= a and not b;
    layer4_outputs(1676) <= not a;
    layer4_outputs(1677) <= not b or a;
    layer4_outputs(1678) <= b and not a;
    layer4_outputs(1679) <= '1';
    layer4_outputs(1680) <= not b or a;
    layer4_outputs(1681) <= a and not b;
    layer4_outputs(1682) <= not (a or b);
    layer4_outputs(1683) <= b and not a;
    layer4_outputs(1684) <= not b or a;
    layer4_outputs(1685) <= '1';
    layer4_outputs(1686) <= not (a and b);
    layer4_outputs(1687) <= a xor b;
    layer4_outputs(1688) <= a;
    layer4_outputs(1689) <= not (a or b);
    layer4_outputs(1690) <= '1';
    layer4_outputs(1691) <= a and b;
    layer4_outputs(1692) <= not b;
    layer4_outputs(1693) <= not (a xor b);
    layer4_outputs(1694) <= not (a or b);
    layer4_outputs(1695) <= not a or b;
    layer4_outputs(1696) <= a and not b;
    layer4_outputs(1697) <= not (a and b);
    layer4_outputs(1698) <= a and not b;
    layer4_outputs(1699) <= not b or a;
    layer4_outputs(1700) <= a and b;
    layer4_outputs(1701) <= a and not b;
    layer4_outputs(1702) <= not a;
    layer4_outputs(1703) <= not b;
    layer4_outputs(1704) <= not (a or b);
    layer4_outputs(1705) <= not a or b;
    layer4_outputs(1706) <= '0';
    layer4_outputs(1707) <= not b;
    layer4_outputs(1708) <= not a;
    layer4_outputs(1709) <= not a;
    layer4_outputs(1710) <= b and not a;
    layer4_outputs(1711) <= not (a and b);
    layer4_outputs(1712) <= not a;
    layer4_outputs(1713) <= a xor b;
    layer4_outputs(1714) <= b and not a;
    layer4_outputs(1715) <= b;
    layer4_outputs(1716) <= a and not b;
    layer4_outputs(1717) <= b and not a;
    layer4_outputs(1718) <= not (a or b);
    layer4_outputs(1719) <= a and not b;
    layer4_outputs(1720) <= not a or b;
    layer4_outputs(1721) <= '1';
    layer4_outputs(1722) <= not a or b;
    layer4_outputs(1723) <= not (a and b);
    layer4_outputs(1724) <= a;
    layer4_outputs(1725) <= a and b;
    layer4_outputs(1726) <= '1';
    layer4_outputs(1727) <= '0';
    layer4_outputs(1728) <= b;
    layer4_outputs(1729) <= not (a or b);
    layer4_outputs(1730) <= not (a and b);
    layer4_outputs(1731) <= b;
    layer4_outputs(1732) <= not (a or b);
    layer4_outputs(1733) <= not (a or b);
    layer4_outputs(1734) <= not a;
    layer4_outputs(1735) <= a;
    layer4_outputs(1736) <= not (a xor b);
    layer4_outputs(1737) <= a and b;
    layer4_outputs(1738) <= b;
    layer4_outputs(1739) <= a and not b;
    layer4_outputs(1740) <= a;
    layer4_outputs(1741) <= not (a or b);
    layer4_outputs(1742) <= '1';
    layer4_outputs(1743) <= not b or a;
    layer4_outputs(1744) <= a and not b;
    layer4_outputs(1745) <= a;
    layer4_outputs(1746) <= not a;
    layer4_outputs(1747) <= a and not b;
    layer4_outputs(1748) <= a or b;
    layer4_outputs(1749) <= not a or b;
    layer4_outputs(1750) <= not a;
    layer4_outputs(1751) <= a or b;
    layer4_outputs(1752) <= '1';
    layer4_outputs(1753) <= a and b;
    layer4_outputs(1754) <= not (a and b);
    layer4_outputs(1755) <= not b;
    layer4_outputs(1756) <= a;
    layer4_outputs(1757) <= '0';
    layer4_outputs(1758) <= '1';
    layer4_outputs(1759) <= a or b;
    layer4_outputs(1760) <= b and not a;
    layer4_outputs(1761) <= not (a or b);
    layer4_outputs(1762) <= b;
    layer4_outputs(1763) <= not b or a;
    layer4_outputs(1764) <= a xor b;
    layer4_outputs(1765) <= a;
    layer4_outputs(1766) <= '0';
    layer4_outputs(1767) <= a and not b;
    layer4_outputs(1768) <= b and not a;
    layer4_outputs(1769) <= b;
    layer4_outputs(1770) <= not a;
    layer4_outputs(1771) <= not a;
    layer4_outputs(1772) <= b;
    layer4_outputs(1773) <= not a or b;
    layer4_outputs(1774) <= not b or a;
    layer4_outputs(1775) <= a;
    layer4_outputs(1776) <= not a;
    layer4_outputs(1777) <= not (a or b);
    layer4_outputs(1778) <= not b or a;
    layer4_outputs(1779) <= not a;
    layer4_outputs(1780) <= not b or a;
    layer4_outputs(1781) <= not b;
    layer4_outputs(1782) <= a and not b;
    layer4_outputs(1783) <= not b;
    layer4_outputs(1784) <= not b or a;
    layer4_outputs(1785) <= '0';
    layer4_outputs(1786) <= '0';
    layer4_outputs(1787) <= not b;
    layer4_outputs(1788) <= b;
    layer4_outputs(1789) <= b and not a;
    layer4_outputs(1790) <= not (a and b);
    layer4_outputs(1791) <= '1';
    layer4_outputs(1792) <= '1';
    layer4_outputs(1793) <= b and not a;
    layer4_outputs(1794) <= not (a or b);
    layer4_outputs(1795) <= not a or b;
    layer4_outputs(1796) <= not b;
    layer4_outputs(1797) <= a;
    layer4_outputs(1798) <= '1';
    layer4_outputs(1799) <= not b;
    layer4_outputs(1800) <= a and not b;
    layer4_outputs(1801) <= a and not b;
    layer4_outputs(1802) <= not (a and b);
    layer4_outputs(1803) <= not a or b;
    layer4_outputs(1804) <= not b;
    layer4_outputs(1805) <= not a;
    layer4_outputs(1806) <= b and not a;
    layer4_outputs(1807) <= a or b;
    layer4_outputs(1808) <= b and not a;
    layer4_outputs(1809) <= a;
    layer4_outputs(1810) <= a and b;
    layer4_outputs(1811) <= not (a or b);
    layer4_outputs(1812) <= not (a and b);
    layer4_outputs(1813) <= not (a or b);
    layer4_outputs(1814) <= a or b;
    layer4_outputs(1815) <= not a or b;
    layer4_outputs(1816) <= a and not b;
    layer4_outputs(1817) <= b;
    layer4_outputs(1818) <= b and not a;
    layer4_outputs(1819) <= a or b;
    layer4_outputs(1820) <= a and b;
    layer4_outputs(1821) <= '1';
    layer4_outputs(1822) <= a and not b;
    layer4_outputs(1823) <= '1';
    layer4_outputs(1824) <= not a;
    layer4_outputs(1825) <= b and not a;
    layer4_outputs(1826) <= '1';
    layer4_outputs(1827) <= a;
    layer4_outputs(1828) <= b and not a;
    layer4_outputs(1829) <= b and not a;
    layer4_outputs(1830) <= '1';
    layer4_outputs(1831) <= not a or b;
    layer4_outputs(1832) <= not b;
    layer4_outputs(1833) <= not a or b;
    layer4_outputs(1834) <= a xor b;
    layer4_outputs(1835) <= a and b;
    layer4_outputs(1836) <= not a or b;
    layer4_outputs(1837) <= not a;
    layer4_outputs(1838) <= b and not a;
    layer4_outputs(1839) <= a and b;
    layer4_outputs(1840) <= '1';
    layer4_outputs(1841) <= b and not a;
    layer4_outputs(1842) <= not (a and b);
    layer4_outputs(1843) <= not (a and b);
    layer4_outputs(1844) <= a or b;
    layer4_outputs(1845) <= a;
    layer4_outputs(1846) <= a or b;
    layer4_outputs(1847) <= not a;
    layer4_outputs(1848) <= a;
    layer4_outputs(1849) <= not (a and b);
    layer4_outputs(1850) <= not b or a;
    layer4_outputs(1851) <= a and b;
    layer4_outputs(1852) <= not b or a;
    layer4_outputs(1853) <= not b;
    layer4_outputs(1854) <= a or b;
    layer4_outputs(1855) <= a and not b;
    layer4_outputs(1856) <= not (a or b);
    layer4_outputs(1857) <= not a or b;
    layer4_outputs(1858) <= a or b;
    layer4_outputs(1859) <= not (a or b);
    layer4_outputs(1860) <= b;
    layer4_outputs(1861) <= not a or b;
    layer4_outputs(1862) <= not (a or b);
    layer4_outputs(1863) <= '1';
    layer4_outputs(1864) <= a;
    layer4_outputs(1865) <= not b;
    layer4_outputs(1866) <= a and b;
    layer4_outputs(1867) <= '1';
    layer4_outputs(1868) <= not (a xor b);
    layer4_outputs(1869) <= b;
    layer4_outputs(1870) <= not b or a;
    layer4_outputs(1871) <= a or b;
    layer4_outputs(1872) <= not a;
    layer4_outputs(1873) <= a and not b;
    layer4_outputs(1874) <= not b or a;
    layer4_outputs(1875) <= b and not a;
    layer4_outputs(1876) <= b and not a;
    layer4_outputs(1877) <= a xor b;
    layer4_outputs(1878) <= not a or b;
    layer4_outputs(1879) <= b and not a;
    layer4_outputs(1880) <= not (a xor b);
    layer4_outputs(1881) <= not (a and b);
    layer4_outputs(1882) <= a;
    layer4_outputs(1883) <= '1';
    layer4_outputs(1884) <= b and not a;
    layer4_outputs(1885) <= a and not b;
    layer4_outputs(1886) <= not (a and b);
    layer4_outputs(1887) <= not (a or b);
    layer4_outputs(1888) <= b;
    layer4_outputs(1889) <= not b;
    layer4_outputs(1890) <= a xor b;
    layer4_outputs(1891) <= not b;
    layer4_outputs(1892) <= a;
    layer4_outputs(1893) <= not b or a;
    layer4_outputs(1894) <= '1';
    layer4_outputs(1895) <= a and not b;
    layer4_outputs(1896) <= a;
    layer4_outputs(1897) <= not b;
    layer4_outputs(1898) <= not (a or b);
    layer4_outputs(1899) <= a;
    layer4_outputs(1900) <= a and not b;
    layer4_outputs(1901) <= '0';
    layer4_outputs(1902) <= not a or b;
    layer4_outputs(1903) <= not (a xor b);
    layer4_outputs(1904) <= not a;
    layer4_outputs(1905) <= a and b;
    layer4_outputs(1906) <= a xor b;
    layer4_outputs(1907) <= a and b;
    layer4_outputs(1908) <= a;
    layer4_outputs(1909) <= not a;
    layer4_outputs(1910) <= a;
    layer4_outputs(1911) <= a and not b;
    layer4_outputs(1912) <= a or b;
    layer4_outputs(1913) <= '0';
    layer4_outputs(1914) <= a or b;
    layer4_outputs(1915) <= a;
    layer4_outputs(1916) <= b;
    layer4_outputs(1917) <= not b or a;
    layer4_outputs(1918) <= a and b;
    layer4_outputs(1919) <= not (a or b);
    layer4_outputs(1920) <= a;
    layer4_outputs(1921) <= not b;
    layer4_outputs(1922) <= a or b;
    layer4_outputs(1923) <= not (a or b);
    layer4_outputs(1924) <= b and not a;
    layer4_outputs(1925) <= not b or a;
    layer4_outputs(1926) <= not a;
    layer4_outputs(1927) <= b;
    layer4_outputs(1928) <= not (a or b);
    layer4_outputs(1929) <= b;
    layer4_outputs(1930) <= not a or b;
    layer4_outputs(1931) <= not (a or b);
    layer4_outputs(1932) <= a or b;
    layer4_outputs(1933) <= '1';
    layer4_outputs(1934) <= '1';
    layer4_outputs(1935) <= not b or a;
    layer4_outputs(1936) <= not (a xor b);
    layer4_outputs(1937) <= b;
    layer4_outputs(1938) <= '1';
    layer4_outputs(1939) <= a or b;
    layer4_outputs(1940) <= not (a and b);
    layer4_outputs(1941) <= not (a and b);
    layer4_outputs(1942) <= b;
    layer4_outputs(1943) <= not b or a;
    layer4_outputs(1944) <= not a;
    layer4_outputs(1945) <= a and not b;
    layer4_outputs(1946) <= a and not b;
    layer4_outputs(1947) <= b;
    layer4_outputs(1948) <= not b or a;
    layer4_outputs(1949) <= a;
    layer4_outputs(1950) <= b;
    layer4_outputs(1951) <= a and not b;
    layer4_outputs(1952) <= a and not b;
    layer4_outputs(1953) <= not a or b;
    layer4_outputs(1954) <= not b or a;
    layer4_outputs(1955) <= a or b;
    layer4_outputs(1956) <= b and not a;
    layer4_outputs(1957) <= not (a and b);
    layer4_outputs(1958) <= not a or b;
    layer4_outputs(1959) <= '1';
    layer4_outputs(1960) <= not (a or b);
    layer4_outputs(1961) <= b;
    layer4_outputs(1962) <= '1';
    layer4_outputs(1963) <= a;
    layer4_outputs(1964) <= not (a or b);
    layer4_outputs(1965) <= not (a or b);
    layer4_outputs(1966) <= not (a xor b);
    layer4_outputs(1967) <= not b;
    layer4_outputs(1968) <= b;
    layer4_outputs(1969) <= not b;
    layer4_outputs(1970) <= not (a xor b);
    layer4_outputs(1971) <= not b or a;
    layer4_outputs(1972) <= not (a and b);
    layer4_outputs(1973) <= not (a or b);
    layer4_outputs(1974) <= b and not a;
    layer4_outputs(1975) <= a and b;
    layer4_outputs(1976) <= '1';
    layer4_outputs(1977) <= a and not b;
    layer4_outputs(1978) <= '0';
    layer4_outputs(1979) <= a and b;
    layer4_outputs(1980) <= not a or b;
    layer4_outputs(1981) <= '0';
    layer4_outputs(1982) <= b and not a;
    layer4_outputs(1983) <= not b;
    layer4_outputs(1984) <= '1';
    layer4_outputs(1985) <= a and not b;
    layer4_outputs(1986) <= not a or b;
    layer4_outputs(1987) <= a and not b;
    layer4_outputs(1988) <= not b or a;
    layer4_outputs(1989) <= a xor b;
    layer4_outputs(1990) <= b;
    layer4_outputs(1991) <= a and not b;
    layer4_outputs(1992) <= a and not b;
    layer4_outputs(1993) <= not b or a;
    layer4_outputs(1994) <= not (a and b);
    layer4_outputs(1995) <= not b;
    layer4_outputs(1996) <= '0';
    layer4_outputs(1997) <= not a or b;
    layer4_outputs(1998) <= a and b;
    layer4_outputs(1999) <= a and b;
    layer4_outputs(2000) <= not b;
    layer4_outputs(2001) <= a and not b;
    layer4_outputs(2002) <= b;
    layer4_outputs(2003) <= not a or b;
    layer4_outputs(2004) <= b;
    layer4_outputs(2005) <= a;
    layer4_outputs(2006) <= not (a and b);
    layer4_outputs(2007) <= a;
    layer4_outputs(2008) <= a and b;
    layer4_outputs(2009) <= not a or b;
    layer4_outputs(2010) <= b;
    layer4_outputs(2011) <= not b;
    layer4_outputs(2012) <= not b;
    layer4_outputs(2013) <= a and not b;
    layer4_outputs(2014) <= a and not b;
    layer4_outputs(2015) <= a;
    layer4_outputs(2016) <= a and not b;
    layer4_outputs(2017) <= not b or a;
    layer4_outputs(2018) <= '0';
    layer4_outputs(2019) <= a and not b;
    layer4_outputs(2020) <= not (a xor b);
    layer4_outputs(2021) <= not b;
    layer4_outputs(2022) <= a;
    layer4_outputs(2023) <= not a;
    layer4_outputs(2024) <= b;
    layer4_outputs(2025) <= '0';
    layer4_outputs(2026) <= a and not b;
    layer4_outputs(2027) <= '0';
    layer4_outputs(2028) <= b;
    layer4_outputs(2029) <= not (a and b);
    layer4_outputs(2030) <= not b;
    layer4_outputs(2031) <= not a;
    layer4_outputs(2032) <= a and b;
    layer4_outputs(2033) <= not a;
    layer4_outputs(2034) <= not (a or b);
    layer4_outputs(2035) <= not b or a;
    layer4_outputs(2036) <= b;
    layer4_outputs(2037) <= b;
    layer4_outputs(2038) <= not a or b;
    layer4_outputs(2039) <= not (a xor b);
    layer4_outputs(2040) <= a xor b;
    layer4_outputs(2041) <= b;
    layer4_outputs(2042) <= a;
    layer4_outputs(2043) <= a and b;
    layer4_outputs(2044) <= not (a or b);
    layer4_outputs(2045) <= not b or a;
    layer4_outputs(2046) <= a;
    layer4_outputs(2047) <= a and b;
    layer4_outputs(2048) <= not (a or b);
    layer4_outputs(2049) <= b;
    layer4_outputs(2050) <= not b;
    layer4_outputs(2051) <= a or b;
    layer4_outputs(2052) <= b;
    layer4_outputs(2053) <= not a or b;
    layer4_outputs(2054) <= b and not a;
    layer4_outputs(2055) <= a or b;
    layer4_outputs(2056) <= a and not b;
    layer4_outputs(2057) <= b;
    layer4_outputs(2058) <= a and not b;
    layer4_outputs(2059) <= a and b;
    layer4_outputs(2060) <= a;
    layer4_outputs(2061) <= not a or b;
    layer4_outputs(2062) <= '0';
    layer4_outputs(2063) <= not b or a;
    layer4_outputs(2064) <= b;
    layer4_outputs(2065) <= a;
    layer4_outputs(2066) <= not (a xor b);
    layer4_outputs(2067) <= a or b;
    layer4_outputs(2068) <= not b;
    layer4_outputs(2069) <= a or b;
    layer4_outputs(2070) <= not b;
    layer4_outputs(2071) <= a and b;
    layer4_outputs(2072) <= a or b;
    layer4_outputs(2073) <= a;
    layer4_outputs(2074) <= not a;
    layer4_outputs(2075) <= not (a and b);
    layer4_outputs(2076) <= a and not b;
    layer4_outputs(2077) <= a and b;
    layer4_outputs(2078) <= '0';
    layer4_outputs(2079) <= not b;
    layer4_outputs(2080) <= not (a or b);
    layer4_outputs(2081) <= not (a or b);
    layer4_outputs(2082) <= b and not a;
    layer4_outputs(2083) <= not b or a;
    layer4_outputs(2084) <= '0';
    layer4_outputs(2085) <= a and not b;
    layer4_outputs(2086) <= a or b;
    layer4_outputs(2087) <= a;
    layer4_outputs(2088) <= '0';
    layer4_outputs(2089) <= not b;
    layer4_outputs(2090) <= '0';
    layer4_outputs(2091) <= not (a or b);
    layer4_outputs(2092) <= not a or b;
    layer4_outputs(2093) <= not b;
    layer4_outputs(2094) <= '0';
    layer4_outputs(2095) <= '1';
    layer4_outputs(2096) <= a;
    layer4_outputs(2097) <= a and not b;
    layer4_outputs(2098) <= a;
    layer4_outputs(2099) <= not (a or b);
    layer4_outputs(2100) <= not (a or b);
    layer4_outputs(2101) <= a or b;
    layer4_outputs(2102) <= a and b;
    layer4_outputs(2103) <= b;
    layer4_outputs(2104) <= not b;
    layer4_outputs(2105) <= b;
    layer4_outputs(2106) <= a;
    layer4_outputs(2107) <= a and not b;
    layer4_outputs(2108) <= not b;
    layer4_outputs(2109) <= '1';
    layer4_outputs(2110) <= '1';
    layer4_outputs(2111) <= b and not a;
    layer4_outputs(2112) <= not b;
    layer4_outputs(2113) <= not (a xor b);
    layer4_outputs(2114) <= b and not a;
    layer4_outputs(2115) <= not (a or b);
    layer4_outputs(2116) <= not a or b;
    layer4_outputs(2117) <= not a;
    layer4_outputs(2118) <= not a;
    layer4_outputs(2119) <= not a or b;
    layer4_outputs(2120) <= a or b;
    layer4_outputs(2121) <= b and not a;
    layer4_outputs(2122) <= not a or b;
    layer4_outputs(2123) <= a and b;
    layer4_outputs(2124) <= b;
    layer4_outputs(2125) <= not a;
    layer4_outputs(2126) <= not (a or b);
    layer4_outputs(2127) <= '0';
    layer4_outputs(2128) <= a and b;
    layer4_outputs(2129) <= b and not a;
    layer4_outputs(2130) <= b;
    layer4_outputs(2131) <= not (a and b);
    layer4_outputs(2132) <= a and b;
    layer4_outputs(2133) <= a xor b;
    layer4_outputs(2134) <= not (a or b);
    layer4_outputs(2135) <= not (a and b);
    layer4_outputs(2136) <= not (a or b);
    layer4_outputs(2137) <= not a or b;
    layer4_outputs(2138) <= a and b;
    layer4_outputs(2139) <= a and b;
    layer4_outputs(2140) <= '0';
    layer4_outputs(2141) <= not b;
    layer4_outputs(2142) <= a;
    layer4_outputs(2143) <= a or b;
    layer4_outputs(2144) <= a and b;
    layer4_outputs(2145) <= a;
    layer4_outputs(2146) <= a;
    layer4_outputs(2147) <= a xor b;
    layer4_outputs(2148) <= not a or b;
    layer4_outputs(2149) <= not a or b;
    layer4_outputs(2150) <= b;
    layer4_outputs(2151) <= a and not b;
    layer4_outputs(2152) <= a and b;
    layer4_outputs(2153) <= a;
    layer4_outputs(2154) <= not (a and b);
    layer4_outputs(2155) <= a and not b;
    layer4_outputs(2156) <= not (a or b);
    layer4_outputs(2157) <= b;
    layer4_outputs(2158) <= b;
    layer4_outputs(2159) <= a;
    layer4_outputs(2160) <= '1';
    layer4_outputs(2161) <= b;
    layer4_outputs(2162) <= not b;
    layer4_outputs(2163) <= a and not b;
    layer4_outputs(2164) <= a and not b;
    layer4_outputs(2165) <= not b or a;
    layer4_outputs(2166) <= not a or b;
    layer4_outputs(2167) <= not a;
    layer4_outputs(2168) <= a and b;
    layer4_outputs(2169) <= not a or b;
    layer4_outputs(2170) <= a or b;
    layer4_outputs(2171) <= a and not b;
    layer4_outputs(2172) <= a and not b;
    layer4_outputs(2173) <= not (a or b);
    layer4_outputs(2174) <= a and not b;
    layer4_outputs(2175) <= a and b;
    layer4_outputs(2176) <= b and not a;
    layer4_outputs(2177) <= not (a and b);
    layer4_outputs(2178) <= a;
    layer4_outputs(2179) <= a;
    layer4_outputs(2180) <= '1';
    layer4_outputs(2181) <= a xor b;
    layer4_outputs(2182) <= not a or b;
    layer4_outputs(2183) <= not b or a;
    layer4_outputs(2184) <= a;
    layer4_outputs(2185) <= a and b;
    layer4_outputs(2186) <= not a or b;
    layer4_outputs(2187) <= '0';
    layer4_outputs(2188) <= a;
    layer4_outputs(2189) <= '0';
    layer4_outputs(2190) <= a and b;
    layer4_outputs(2191) <= not (a xor b);
    layer4_outputs(2192) <= a and not b;
    layer4_outputs(2193) <= not b;
    layer4_outputs(2194) <= not b or a;
    layer4_outputs(2195) <= not b or a;
    layer4_outputs(2196) <= a and b;
    layer4_outputs(2197) <= not a or b;
    layer4_outputs(2198) <= a and not b;
    layer4_outputs(2199) <= '1';
    layer4_outputs(2200) <= '1';
    layer4_outputs(2201) <= a;
    layer4_outputs(2202) <= not a;
    layer4_outputs(2203) <= b;
    layer4_outputs(2204) <= b;
    layer4_outputs(2205) <= b;
    layer4_outputs(2206) <= a and b;
    layer4_outputs(2207) <= a xor b;
    layer4_outputs(2208) <= a or b;
    layer4_outputs(2209) <= not (a and b);
    layer4_outputs(2210) <= b and not a;
    layer4_outputs(2211) <= not b;
    layer4_outputs(2212) <= not (a and b);
    layer4_outputs(2213) <= not b;
    layer4_outputs(2214) <= a or b;
    layer4_outputs(2215) <= b and not a;
    layer4_outputs(2216) <= not (a xor b);
    layer4_outputs(2217) <= not a or b;
    layer4_outputs(2218) <= '0';
    layer4_outputs(2219) <= not (a and b);
    layer4_outputs(2220) <= a and b;
    layer4_outputs(2221) <= '0';
    layer4_outputs(2222) <= b and not a;
    layer4_outputs(2223) <= not (a xor b);
    layer4_outputs(2224) <= not (a xor b);
    layer4_outputs(2225) <= b;
    layer4_outputs(2226) <= not a or b;
    layer4_outputs(2227) <= not b;
    layer4_outputs(2228) <= not (a or b);
    layer4_outputs(2229) <= a xor b;
    layer4_outputs(2230) <= '0';
    layer4_outputs(2231) <= '0';
    layer4_outputs(2232) <= not (a and b);
    layer4_outputs(2233) <= b;
    layer4_outputs(2234) <= b and not a;
    layer4_outputs(2235) <= b;
    layer4_outputs(2236) <= not (a and b);
    layer4_outputs(2237) <= b;
    layer4_outputs(2238) <= not b;
    layer4_outputs(2239) <= '0';
    layer4_outputs(2240) <= '1';
    layer4_outputs(2241) <= a;
    layer4_outputs(2242) <= not a;
    layer4_outputs(2243) <= a xor b;
    layer4_outputs(2244) <= not b or a;
    layer4_outputs(2245) <= not (a xor b);
    layer4_outputs(2246) <= not (a and b);
    layer4_outputs(2247) <= a;
    layer4_outputs(2248) <= '1';
    layer4_outputs(2249) <= not (a or b);
    layer4_outputs(2250) <= '1';
    layer4_outputs(2251) <= not a or b;
    layer4_outputs(2252) <= b;
    layer4_outputs(2253) <= a and not b;
    layer4_outputs(2254) <= a;
    layer4_outputs(2255) <= a and b;
    layer4_outputs(2256) <= not (a and b);
    layer4_outputs(2257) <= '1';
    layer4_outputs(2258) <= a xor b;
    layer4_outputs(2259) <= a;
    layer4_outputs(2260) <= a and not b;
    layer4_outputs(2261) <= not a or b;
    layer4_outputs(2262) <= not b;
    layer4_outputs(2263) <= a and b;
    layer4_outputs(2264) <= a xor b;
    layer4_outputs(2265) <= not (a or b);
    layer4_outputs(2266) <= a and not b;
    layer4_outputs(2267) <= a or b;
    layer4_outputs(2268) <= not (a xor b);
    layer4_outputs(2269) <= not (a or b);
    layer4_outputs(2270) <= not b;
    layer4_outputs(2271) <= '0';
    layer4_outputs(2272) <= not a;
    layer4_outputs(2273) <= not a;
    layer4_outputs(2274) <= a and not b;
    layer4_outputs(2275) <= a;
    layer4_outputs(2276) <= b and not a;
    layer4_outputs(2277) <= not a;
    layer4_outputs(2278) <= a xor b;
    layer4_outputs(2279) <= '0';
    layer4_outputs(2280) <= not a;
    layer4_outputs(2281) <= not a or b;
    layer4_outputs(2282) <= not a;
    layer4_outputs(2283) <= not b or a;
    layer4_outputs(2284) <= a or b;
    layer4_outputs(2285) <= not b;
    layer4_outputs(2286) <= a;
    layer4_outputs(2287) <= not (a or b);
    layer4_outputs(2288) <= not a;
    layer4_outputs(2289) <= b;
    layer4_outputs(2290) <= not a or b;
    layer4_outputs(2291) <= a or b;
    layer4_outputs(2292) <= a and b;
    layer4_outputs(2293) <= b;
    layer4_outputs(2294) <= a and b;
    layer4_outputs(2295) <= not b;
    layer4_outputs(2296) <= a or b;
    layer4_outputs(2297) <= '1';
    layer4_outputs(2298) <= not a;
    layer4_outputs(2299) <= not a;
    layer4_outputs(2300) <= a and not b;
    layer4_outputs(2301) <= not a;
    layer4_outputs(2302) <= not b or a;
    layer4_outputs(2303) <= '0';
    layer4_outputs(2304) <= a or b;
    layer4_outputs(2305) <= not (a and b);
    layer4_outputs(2306) <= not b or a;
    layer4_outputs(2307) <= not b or a;
    layer4_outputs(2308) <= '1';
    layer4_outputs(2309) <= not a or b;
    layer4_outputs(2310) <= not (a xor b);
    layer4_outputs(2311) <= b and not a;
    layer4_outputs(2312) <= not (a and b);
    layer4_outputs(2313) <= not (a or b);
    layer4_outputs(2314) <= not (a or b);
    layer4_outputs(2315) <= a and b;
    layer4_outputs(2316) <= not a or b;
    layer4_outputs(2317) <= not a or b;
    layer4_outputs(2318) <= b;
    layer4_outputs(2319) <= not (a or b);
    layer4_outputs(2320) <= not b;
    layer4_outputs(2321) <= b;
    layer4_outputs(2322) <= a xor b;
    layer4_outputs(2323) <= not (a or b);
    layer4_outputs(2324) <= not b;
    layer4_outputs(2325) <= '0';
    layer4_outputs(2326) <= b;
    layer4_outputs(2327) <= not b;
    layer4_outputs(2328) <= a;
    layer4_outputs(2329) <= a;
    layer4_outputs(2330) <= a or b;
    layer4_outputs(2331) <= not a or b;
    layer4_outputs(2332) <= '1';
    layer4_outputs(2333) <= a;
    layer4_outputs(2334) <= not b;
    layer4_outputs(2335) <= a or b;
    layer4_outputs(2336) <= b;
    layer4_outputs(2337) <= b and not a;
    layer4_outputs(2338) <= not b;
    layer4_outputs(2339) <= a;
    layer4_outputs(2340) <= not a;
    layer4_outputs(2341) <= a and not b;
    layer4_outputs(2342) <= b;
    layer4_outputs(2343) <= not a or b;
    layer4_outputs(2344) <= not (a xor b);
    layer4_outputs(2345) <= a and not b;
    layer4_outputs(2346) <= not (a and b);
    layer4_outputs(2347) <= not b;
    layer4_outputs(2348) <= a and b;
    layer4_outputs(2349) <= a and b;
    layer4_outputs(2350) <= not b or a;
    layer4_outputs(2351) <= a and not b;
    layer4_outputs(2352) <= a or b;
    layer4_outputs(2353) <= a xor b;
    layer4_outputs(2354) <= a;
    layer4_outputs(2355) <= a and not b;
    layer4_outputs(2356) <= not (a or b);
    layer4_outputs(2357) <= not a;
    layer4_outputs(2358) <= a;
    layer4_outputs(2359) <= not (a or b);
    layer4_outputs(2360) <= b;
    layer4_outputs(2361) <= a or b;
    layer4_outputs(2362) <= not (a or b);
    layer4_outputs(2363) <= not a or b;
    layer4_outputs(2364) <= a and not b;
    layer4_outputs(2365) <= not b;
    layer4_outputs(2366) <= a xor b;
    layer4_outputs(2367) <= not (a or b);
    layer4_outputs(2368) <= a and not b;
    layer4_outputs(2369) <= not a;
    layer4_outputs(2370) <= b;
    layer4_outputs(2371) <= not b;
    layer4_outputs(2372) <= not b;
    layer4_outputs(2373) <= a;
    layer4_outputs(2374) <= a;
    layer4_outputs(2375) <= not (a and b);
    layer4_outputs(2376) <= not (a and b);
    layer4_outputs(2377) <= not b or a;
    layer4_outputs(2378) <= a and b;
    layer4_outputs(2379) <= a and not b;
    layer4_outputs(2380) <= a;
    layer4_outputs(2381) <= not a or b;
    layer4_outputs(2382) <= b;
    layer4_outputs(2383) <= a and not b;
    layer4_outputs(2384) <= not a;
    layer4_outputs(2385) <= '0';
    layer4_outputs(2386) <= not a or b;
    layer4_outputs(2387) <= b and not a;
    layer4_outputs(2388) <= b;
    layer4_outputs(2389) <= a and b;
    layer4_outputs(2390) <= not a;
    layer4_outputs(2391) <= '0';
    layer4_outputs(2392) <= not b;
    layer4_outputs(2393) <= a xor b;
    layer4_outputs(2394) <= b and not a;
    layer4_outputs(2395) <= a;
    layer4_outputs(2396) <= not a or b;
    layer4_outputs(2397) <= not b;
    layer4_outputs(2398) <= a and b;
    layer4_outputs(2399) <= a and not b;
    layer4_outputs(2400) <= '1';
    layer4_outputs(2401) <= not a;
    layer4_outputs(2402) <= '1';
    layer4_outputs(2403) <= not b;
    layer4_outputs(2404) <= b and not a;
    layer4_outputs(2405) <= not a;
    layer4_outputs(2406) <= not (a or b);
    layer4_outputs(2407) <= '0';
    layer4_outputs(2408) <= a and b;
    layer4_outputs(2409) <= a and not b;
    layer4_outputs(2410) <= a;
    layer4_outputs(2411) <= a and not b;
    layer4_outputs(2412) <= a;
    layer4_outputs(2413) <= not a;
    layer4_outputs(2414) <= a and b;
    layer4_outputs(2415) <= b;
    layer4_outputs(2416) <= not (a and b);
    layer4_outputs(2417) <= b;
    layer4_outputs(2418) <= '1';
    layer4_outputs(2419) <= a and b;
    layer4_outputs(2420) <= not b or a;
    layer4_outputs(2421) <= not b or a;
    layer4_outputs(2422) <= not a or b;
    layer4_outputs(2423) <= b;
    layer4_outputs(2424) <= '1';
    layer4_outputs(2425) <= '0';
    layer4_outputs(2426) <= not (a and b);
    layer4_outputs(2427) <= '1';
    layer4_outputs(2428) <= not a;
    layer4_outputs(2429) <= b;
    layer4_outputs(2430) <= not b;
    layer4_outputs(2431) <= a xor b;
    layer4_outputs(2432) <= not b;
    layer4_outputs(2433) <= a or b;
    layer4_outputs(2434) <= not (a and b);
    layer4_outputs(2435) <= a xor b;
    layer4_outputs(2436) <= a;
    layer4_outputs(2437) <= not b or a;
    layer4_outputs(2438) <= not a;
    layer4_outputs(2439) <= b and not a;
    layer4_outputs(2440) <= not (a xor b);
    layer4_outputs(2441) <= '0';
    layer4_outputs(2442) <= not a or b;
    layer4_outputs(2443) <= '1';
    layer4_outputs(2444) <= a or b;
    layer4_outputs(2445) <= a xor b;
    layer4_outputs(2446) <= not (a and b);
    layer4_outputs(2447) <= a and not b;
    layer4_outputs(2448) <= not b;
    layer4_outputs(2449) <= a and b;
    layer4_outputs(2450) <= a and not b;
    layer4_outputs(2451) <= not b;
    layer4_outputs(2452) <= b;
    layer4_outputs(2453) <= not a;
    layer4_outputs(2454) <= '0';
    layer4_outputs(2455) <= not (a or b);
    layer4_outputs(2456) <= not a;
    layer4_outputs(2457) <= a or b;
    layer4_outputs(2458) <= not b or a;
    layer4_outputs(2459) <= not b or a;
    layer4_outputs(2460) <= a and not b;
    layer4_outputs(2461) <= a and not b;
    layer4_outputs(2462) <= not (a or b);
    layer4_outputs(2463) <= a xor b;
    layer4_outputs(2464) <= not (a or b);
    layer4_outputs(2465) <= '1';
    layer4_outputs(2466) <= '0';
    layer4_outputs(2467) <= b;
    layer4_outputs(2468) <= '1';
    layer4_outputs(2469) <= '0';
    layer4_outputs(2470) <= a and b;
    layer4_outputs(2471) <= b and not a;
    layer4_outputs(2472) <= not a;
    layer4_outputs(2473) <= not b or a;
    layer4_outputs(2474) <= '1';
    layer4_outputs(2475) <= a or b;
    layer4_outputs(2476) <= not (a or b);
    layer4_outputs(2477) <= b and not a;
    layer4_outputs(2478) <= a;
    layer4_outputs(2479) <= a or b;
    layer4_outputs(2480) <= b;
    layer4_outputs(2481) <= not (a or b);
    layer4_outputs(2482) <= not a;
    layer4_outputs(2483) <= not (a and b);
    layer4_outputs(2484) <= not a;
    layer4_outputs(2485) <= not a;
    layer4_outputs(2486) <= a or b;
    layer4_outputs(2487) <= not a;
    layer4_outputs(2488) <= not (a xor b);
    layer4_outputs(2489) <= b;
    layer4_outputs(2490) <= a xor b;
    layer4_outputs(2491) <= '1';
    layer4_outputs(2492) <= a;
    layer4_outputs(2493) <= a and not b;
    layer4_outputs(2494) <= a and b;
    layer4_outputs(2495) <= b and not a;
    layer4_outputs(2496) <= not a or b;
    layer4_outputs(2497) <= not b;
    layer4_outputs(2498) <= not (a or b);
    layer4_outputs(2499) <= '1';
    layer4_outputs(2500) <= not b;
    layer4_outputs(2501) <= not a or b;
    layer4_outputs(2502) <= '0';
    layer4_outputs(2503) <= '1';
    layer4_outputs(2504) <= '1';
    layer4_outputs(2505) <= not (a and b);
    layer4_outputs(2506) <= not (a and b);
    layer4_outputs(2507) <= a and b;
    layer4_outputs(2508) <= a and b;
    layer4_outputs(2509) <= a or b;
    layer4_outputs(2510) <= b and not a;
    layer4_outputs(2511) <= '1';
    layer4_outputs(2512) <= a and not b;
    layer4_outputs(2513) <= not (a and b);
    layer4_outputs(2514) <= a;
    layer4_outputs(2515) <= a and b;
    layer4_outputs(2516) <= a and not b;
    layer4_outputs(2517) <= '1';
    layer4_outputs(2518) <= '0';
    layer4_outputs(2519) <= not a;
    layer4_outputs(2520) <= not a;
    layer4_outputs(2521) <= not b or a;
    layer4_outputs(2522) <= a or b;
    layer4_outputs(2523) <= a and not b;
    layer4_outputs(2524) <= not b or a;
    layer4_outputs(2525) <= '0';
    layer4_outputs(2526) <= b;
    layer4_outputs(2527) <= '1';
    layer4_outputs(2528) <= a;
    layer4_outputs(2529) <= b;
    layer4_outputs(2530) <= a and not b;
    layer4_outputs(2531) <= b and not a;
    layer4_outputs(2532) <= a or b;
    layer4_outputs(2533) <= b;
    layer4_outputs(2534) <= '0';
    layer4_outputs(2535) <= b and not a;
    layer4_outputs(2536) <= a and b;
    layer4_outputs(2537) <= b and not a;
    layer4_outputs(2538) <= not a;
    layer4_outputs(2539) <= not b;
    layer4_outputs(2540) <= b and not a;
    layer4_outputs(2541) <= not b;
    layer4_outputs(2542) <= b;
    layer4_outputs(2543) <= a;
    layer4_outputs(2544) <= not (a and b);
    layer4_outputs(2545) <= '1';
    layer4_outputs(2546) <= not a or b;
    layer4_outputs(2547) <= not b or a;
    layer4_outputs(2548) <= a and b;
    layer4_outputs(2549) <= a;
    layer4_outputs(2550) <= b;
    layer4_outputs(2551) <= not a or b;
    layer4_outputs(2552) <= not a;
    layer4_outputs(2553) <= b;
    layer4_outputs(2554) <= not a or b;
    layer4_outputs(2555) <= '1';
    layer4_outputs(2556) <= not a;
    layer4_outputs(2557) <= not b or a;
    layer4_outputs(2558) <= not b;
    layer4_outputs(2559) <= b and not a;
    layer4_outputs(2560) <= b;
    layer4_outputs(2561) <= b;
    layer4_outputs(2562) <= not (a and b);
    layer4_outputs(2563) <= b and not a;
    layer4_outputs(2564) <= not b or a;
    layer4_outputs(2565) <= not a;
    layer4_outputs(2566) <= b;
    layer4_outputs(2567) <= b;
    layer4_outputs(2568) <= a and not b;
    layer4_outputs(2569) <= not (a and b);
    layer4_outputs(2570) <= a or b;
    layer4_outputs(2571) <= b;
    layer4_outputs(2572) <= b;
    layer4_outputs(2573) <= b and not a;
    layer4_outputs(2574) <= b;
    layer4_outputs(2575) <= a xor b;
    layer4_outputs(2576) <= a;
    layer4_outputs(2577) <= a and not b;
    layer4_outputs(2578) <= not b;
    layer4_outputs(2579) <= '0';
    layer4_outputs(2580) <= not b;
    layer4_outputs(2581) <= a and not b;
    layer4_outputs(2582) <= not b;
    layer4_outputs(2583) <= b and not a;
    layer4_outputs(2584) <= not b;
    layer4_outputs(2585) <= '0';
    layer4_outputs(2586) <= not b or a;
    layer4_outputs(2587) <= a and not b;
    layer4_outputs(2588) <= not b;
    layer4_outputs(2589) <= not b or a;
    layer4_outputs(2590) <= not a;
    layer4_outputs(2591) <= not (a and b);
    layer4_outputs(2592) <= not a or b;
    layer4_outputs(2593) <= '0';
    layer4_outputs(2594) <= not a;
    layer4_outputs(2595) <= b;
    layer4_outputs(2596) <= b;
    layer4_outputs(2597) <= not (a xor b);
    layer4_outputs(2598) <= not (a and b);
    layer4_outputs(2599) <= a;
    layer4_outputs(2600) <= '1';
    layer4_outputs(2601) <= not (a xor b);
    layer4_outputs(2602) <= '0';
    layer4_outputs(2603) <= a xor b;
    layer4_outputs(2604) <= a and not b;
    layer4_outputs(2605) <= not b;
    layer4_outputs(2606) <= a and b;
    layer4_outputs(2607) <= not a;
    layer4_outputs(2608) <= a or b;
    layer4_outputs(2609) <= not (a xor b);
    layer4_outputs(2610) <= a xor b;
    layer4_outputs(2611) <= not b or a;
    layer4_outputs(2612) <= '0';
    layer4_outputs(2613) <= not (a and b);
    layer4_outputs(2614) <= a or b;
    layer4_outputs(2615) <= b;
    layer4_outputs(2616) <= not (a or b);
    layer4_outputs(2617) <= a or b;
    layer4_outputs(2618) <= '0';
    layer4_outputs(2619) <= '0';
    layer4_outputs(2620) <= not a or b;
    layer4_outputs(2621) <= b and not a;
    layer4_outputs(2622) <= not a;
    layer4_outputs(2623) <= not b or a;
    layer4_outputs(2624) <= not (a xor b);
    layer4_outputs(2625) <= a and not b;
    layer4_outputs(2626) <= a and b;
    layer4_outputs(2627) <= not b;
    layer4_outputs(2628) <= not (a or b);
    layer4_outputs(2629) <= b and not a;
    layer4_outputs(2630) <= not (a and b);
    layer4_outputs(2631) <= a and b;
    layer4_outputs(2632) <= a;
    layer4_outputs(2633) <= not b;
    layer4_outputs(2634) <= not a;
    layer4_outputs(2635) <= not a;
    layer4_outputs(2636) <= not (a xor b);
    layer4_outputs(2637) <= a;
    layer4_outputs(2638) <= a;
    layer4_outputs(2639) <= b and not a;
    layer4_outputs(2640) <= '1';
    layer4_outputs(2641) <= b;
    layer4_outputs(2642) <= b and not a;
    layer4_outputs(2643) <= '0';
    layer4_outputs(2644) <= not (a or b);
    layer4_outputs(2645) <= not a or b;
    layer4_outputs(2646) <= a and b;
    layer4_outputs(2647) <= '0';
    layer4_outputs(2648) <= a;
    layer4_outputs(2649) <= not (a or b);
    layer4_outputs(2650) <= not (a and b);
    layer4_outputs(2651) <= not b;
    layer4_outputs(2652) <= a and b;
    layer4_outputs(2653) <= not b or a;
    layer4_outputs(2654) <= a;
    layer4_outputs(2655) <= '0';
    layer4_outputs(2656) <= a and b;
    layer4_outputs(2657) <= b;
    layer4_outputs(2658) <= not (a and b);
    layer4_outputs(2659) <= not a or b;
    layer4_outputs(2660) <= not (a xor b);
    layer4_outputs(2661) <= a and not b;
    layer4_outputs(2662) <= b;
    layer4_outputs(2663) <= '0';
    layer4_outputs(2664) <= '0';
    layer4_outputs(2665) <= a;
    layer4_outputs(2666) <= b and not a;
    layer4_outputs(2667) <= not (a or b);
    layer4_outputs(2668) <= not (a xor b);
    layer4_outputs(2669) <= not b;
    layer4_outputs(2670) <= b and not a;
    layer4_outputs(2671) <= not a or b;
    layer4_outputs(2672) <= not a;
    layer4_outputs(2673) <= b and not a;
    layer4_outputs(2674) <= not (a or b);
    layer4_outputs(2675) <= not a;
    layer4_outputs(2676) <= a and b;
    layer4_outputs(2677) <= not (a and b);
    layer4_outputs(2678) <= not a;
    layer4_outputs(2679) <= a or b;
    layer4_outputs(2680) <= b and not a;
    layer4_outputs(2681) <= not (a xor b);
    layer4_outputs(2682) <= not a or b;
    layer4_outputs(2683) <= b;
    layer4_outputs(2684) <= '1';
    layer4_outputs(2685) <= a;
    layer4_outputs(2686) <= a and not b;
    layer4_outputs(2687) <= not (a and b);
    layer4_outputs(2688) <= not b or a;
    layer4_outputs(2689) <= a or b;
    layer4_outputs(2690) <= not b;
    layer4_outputs(2691) <= b and not a;
    layer4_outputs(2692) <= not b;
    layer4_outputs(2693) <= '1';
    layer4_outputs(2694) <= not a or b;
    layer4_outputs(2695) <= b;
    layer4_outputs(2696) <= a and b;
    layer4_outputs(2697) <= not (a or b);
    layer4_outputs(2698) <= not (a or b);
    layer4_outputs(2699) <= a;
    layer4_outputs(2700) <= a and b;
    layer4_outputs(2701) <= a;
    layer4_outputs(2702) <= a;
    layer4_outputs(2703) <= a or b;
    layer4_outputs(2704) <= '1';
    layer4_outputs(2705) <= not (a xor b);
    layer4_outputs(2706) <= not (a and b);
    layer4_outputs(2707) <= '1';
    layer4_outputs(2708) <= a or b;
    layer4_outputs(2709) <= not (a and b);
    layer4_outputs(2710) <= not b or a;
    layer4_outputs(2711) <= not b or a;
    layer4_outputs(2712) <= b;
    layer4_outputs(2713) <= not b or a;
    layer4_outputs(2714) <= a and not b;
    layer4_outputs(2715) <= not b or a;
    layer4_outputs(2716) <= not a or b;
    layer4_outputs(2717) <= a or b;
    layer4_outputs(2718) <= not a or b;
    layer4_outputs(2719) <= a or b;
    layer4_outputs(2720) <= b and not a;
    layer4_outputs(2721) <= a or b;
    layer4_outputs(2722) <= not a;
    layer4_outputs(2723) <= a and b;
    layer4_outputs(2724) <= b and not a;
    layer4_outputs(2725) <= a;
    layer4_outputs(2726) <= b and not a;
    layer4_outputs(2727) <= not (a xor b);
    layer4_outputs(2728) <= '1';
    layer4_outputs(2729) <= a and not b;
    layer4_outputs(2730) <= a;
    layer4_outputs(2731) <= b;
    layer4_outputs(2732) <= not b;
    layer4_outputs(2733) <= not (a and b);
    layer4_outputs(2734) <= not b;
    layer4_outputs(2735) <= '0';
    layer4_outputs(2736) <= a;
    layer4_outputs(2737) <= not b;
    layer4_outputs(2738) <= a;
    layer4_outputs(2739) <= not a;
    layer4_outputs(2740) <= not b;
    layer4_outputs(2741) <= not (a and b);
    layer4_outputs(2742) <= a and not b;
    layer4_outputs(2743) <= '0';
    layer4_outputs(2744) <= '0';
    layer4_outputs(2745) <= a xor b;
    layer4_outputs(2746) <= a;
    layer4_outputs(2747) <= a;
    layer4_outputs(2748) <= not a;
    layer4_outputs(2749) <= a;
    layer4_outputs(2750) <= not (a or b);
    layer4_outputs(2751) <= a xor b;
    layer4_outputs(2752) <= not b or a;
    layer4_outputs(2753) <= '0';
    layer4_outputs(2754) <= not a;
    layer4_outputs(2755) <= a;
    layer4_outputs(2756) <= b;
    layer4_outputs(2757) <= b and not a;
    layer4_outputs(2758) <= b and not a;
    layer4_outputs(2759) <= not b or a;
    layer4_outputs(2760) <= a;
    layer4_outputs(2761) <= not (a and b);
    layer4_outputs(2762) <= a and b;
    layer4_outputs(2763) <= not b or a;
    layer4_outputs(2764) <= not a;
    layer4_outputs(2765) <= '1';
    layer4_outputs(2766) <= not a or b;
    layer4_outputs(2767) <= not a;
    layer4_outputs(2768) <= not a or b;
    layer4_outputs(2769) <= a and b;
    layer4_outputs(2770) <= b;
    layer4_outputs(2771) <= a;
    layer4_outputs(2772) <= not b;
    layer4_outputs(2773) <= not a or b;
    layer4_outputs(2774) <= a;
    layer4_outputs(2775) <= a and b;
    layer4_outputs(2776) <= b;
    layer4_outputs(2777) <= not a or b;
    layer4_outputs(2778) <= b and not a;
    layer4_outputs(2779) <= b;
    layer4_outputs(2780) <= a or b;
    layer4_outputs(2781) <= a;
    layer4_outputs(2782) <= not (a xor b);
    layer4_outputs(2783) <= a;
    layer4_outputs(2784) <= not (a and b);
    layer4_outputs(2785) <= '0';
    layer4_outputs(2786) <= '0';
    layer4_outputs(2787) <= not (a xor b);
    layer4_outputs(2788) <= a and not b;
    layer4_outputs(2789) <= a and b;
    layer4_outputs(2790) <= not (a xor b);
    layer4_outputs(2791) <= a and b;
    layer4_outputs(2792) <= not a or b;
    layer4_outputs(2793) <= a;
    layer4_outputs(2794) <= '0';
    layer4_outputs(2795) <= not (a or b);
    layer4_outputs(2796) <= not (a and b);
    layer4_outputs(2797) <= a and b;
    layer4_outputs(2798) <= not b or a;
    layer4_outputs(2799) <= not a;
    layer4_outputs(2800) <= '0';
    layer4_outputs(2801) <= a and not b;
    layer4_outputs(2802) <= '0';
    layer4_outputs(2803) <= not b;
    layer4_outputs(2804) <= a xor b;
    layer4_outputs(2805) <= not b;
    layer4_outputs(2806) <= not a;
    layer4_outputs(2807) <= a and not b;
    layer4_outputs(2808) <= '0';
    layer4_outputs(2809) <= b and not a;
    layer4_outputs(2810) <= not a or b;
    layer4_outputs(2811) <= a and b;
    layer4_outputs(2812) <= '1';
    layer4_outputs(2813) <= '0';
    layer4_outputs(2814) <= not a or b;
    layer4_outputs(2815) <= not a;
    layer4_outputs(2816) <= not (a xor b);
    layer4_outputs(2817) <= not a or b;
    layer4_outputs(2818) <= a;
    layer4_outputs(2819) <= not a or b;
    layer4_outputs(2820) <= a or b;
    layer4_outputs(2821) <= a and not b;
    layer4_outputs(2822) <= '1';
    layer4_outputs(2823) <= b;
    layer4_outputs(2824) <= not a or b;
    layer4_outputs(2825) <= not a;
    layer4_outputs(2826) <= a and not b;
    layer4_outputs(2827) <= not a or b;
    layer4_outputs(2828) <= not b or a;
    layer4_outputs(2829) <= b and not a;
    layer4_outputs(2830) <= '1';
    layer4_outputs(2831) <= not b or a;
    layer4_outputs(2832) <= not b or a;
    layer4_outputs(2833) <= a and not b;
    layer4_outputs(2834) <= '0';
    layer4_outputs(2835) <= not b;
    layer4_outputs(2836) <= a and not b;
    layer4_outputs(2837) <= not b;
    layer4_outputs(2838) <= a and b;
    layer4_outputs(2839) <= not (a and b);
    layer4_outputs(2840) <= not b or a;
    layer4_outputs(2841) <= not a or b;
    layer4_outputs(2842) <= b;
    layer4_outputs(2843) <= a and b;
    layer4_outputs(2844) <= b and not a;
    layer4_outputs(2845) <= not (a or b);
    layer4_outputs(2846) <= not a;
    layer4_outputs(2847) <= '1';
    layer4_outputs(2848) <= a and not b;
    layer4_outputs(2849) <= a;
    layer4_outputs(2850) <= '1';
    layer4_outputs(2851) <= b;
    layer4_outputs(2852) <= not b;
    layer4_outputs(2853) <= b and not a;
    layer4_outputs(2854) <= b and not a;
    layer4_outputs(2855) <= '0';
    layer4_outputs(2856) <= a or b;
    layer4_outputs(2857) <= a and not b;
    layer4_outputs(2858) <= not b;
    layer4_outputs(2859) <= b and not a;
    layer4_outputs(2860) <= not a;
    layer4_outputs(2861) <= a and not b;
    layer4_outputs(2862) <= '1';
    layer4_outputs(2863) <= a and b;
    layer4_outputs(2864) <= not a;
    layer4_outputs(2865) <= not b or a;
    layer4_outputs(2866) <= not b;
    layer4_outputs(2867) <= not a;
    layer4_outputs(2868) <= not b or a;
    layer4_outputs(2869) <= a or b;
    layer4_outputs(2870) <= not a or b;
    layer4_outputs(2871) <= not a;
    layer4_outputs(2872) <= a and b;
    layer4_outputs(2873) <= not (a or b);
    layer4_outputs(2874) <= a and not b;
    layer4_outputs(2875) <= a and b;
    layer4_outputs(2876) <= a and b;
    layer4_outputs(2877) <= a or b;
    layer4_outputs(2878) <= not b or a;
    layer4_outputs(2879) <= not (a and b);
    layer4_outputs(2880) <= a or b;
    layer4_outputs(2881) <= not (a and b);
    layer4_outputs(2882) <= '0';
    layer4_outputs(2883) <= a and not b;
    layer4_outputs(2884) <= a or b;
    layer4_outputs(2885) <= not (a or b);
    layer4_outputs(2886) <= not (a and b);
    layer4_outputs(2887) <= a and b;
    layer4_outputs(2888) <= not a or b;
    layer4_outputs(2889) <= not a or b;
    layer4_outputs(2890) <= not a;
    layer4_outputs(2891) <= not a or b;
    layer4_outputs(2892) <= not b;
    layer4_outputs(2893) <= not (a and b);
    layer4_outputs(2894) <= b and not a;
    layer4_outputs(2895) <= a and b;
    layer4_outputs(2896) <= '1';
    layer4_outputs(2897) <= not a or b;
    layer4_outputs(2898) <= a and b;
    layer4_outputs(2899) <= b;
    layer4_outputs(2900) <= not (a xor b);
    layer4_outputs(2901) <= not b;
    layer4_outputs(2902) <= not a or b;
    layer4_outputs(2903) <= not b;
    layer4_outputs(2904) <= not b or a;
    layer4_outputs(2905) <= not (a and b);
    layer4_outputs(2906) <= not a;
    layer4_outputs(2907) <= a and b;
    layer4_outputs(2908) <= '0';
    layer4_outputs(2909) <= not b or a;
    layer4_outputs(2910) <= a and not b;
    layer4_outputs(2911) <= not b or a;
    layer4_outputs(2912) <= not (a and b);
    layer4_outputs(2913) <= not (a xor b);
    layer4_outputs(2914) <= a and not b;
    layer4_outputs(2915) <= a or b;
    layer4_outputs(2916) <= b and not a;
    layer4_outputs(2917) <= not a;
    layer4_outputs(2918) <= a and b;
    layer4_outputs(2919) <= b;
    layer4_outputs(2920) <= not b;
    layer4_outputs(2921) <= not a;
    layer4_outputs(2922) <= a and not b;
    layer4_outputs(2923) <= b;
    layer4_outputs(2924) <= a xor b;
    layer4_outputs(2925) <= '1';
    layer4_outputs(2926) <= a;
    layer4_outputs(2927) <= b;
    layer4_outputs(2928) <= not (a and b);
    layer4_outputs(2929) <= not (a xor b);
    layer4_outputs(2930) <= not a;
    layer4_outputs(2931) <= not b or a;
    layer4_outputs(2932) <= not b or a;
    layer4_outputs(2933) <= a and b;
    layer4_outputs(2934) <= a;
    layer4_outputs(2935) <= '1';
    layer4_outputs(2936) <= a;
    layer4_outputs(2937) <= not (a and b);
    layer4_outputs(2938) <= not b;
    layer4_outputs(2939) <= not b or a;
    layer4_outputs(2940) <= not b;
    layer4_outputs(2941) <= a and b;
    layer4_outputs(2942) <= not a;
    layer4_outputs(2943) <= a and b;
    layer4_outputs(2944) <= b;
    layer4_outputs(2945) <= not (a or b);
    layer4_outputs(2946) <= not (a or b);
    layer4_outputs(2947) <= not a;
    layer4_outputs(2948) <= a and not b;
    layer4_outputs(2949) <= not (a and b);
    layer4_outputs(2950) <= a;
    layer4_outputs(2951) <= a;
    layer4_outputs(2952) <= b;
    layer4_outputs(2953) <= b and not a;
    layer4_outputs(2954) <= not (a or b);
    layer4_outputs(2955) <= b;
    layer4_outputs(2956) <= b and not a;
    layer4_outputs(2957) <= a and b;
    layer4_outputs(2958) <= a;
    layer4_outputs(2959) <= not b;
    layer4_outputs(2960) <= not b or a;
    layer4_outputs(2961) <= not b or a;
    layer4_outputs(2962) <= b;
    layer4_outputs(2963) <= a and not b;
    layer4_outputs(2964) <= a and b;
    layer4_outputs(2965) <= not a;
    layer4_outputs(2966) <= not a;
    layer4_outputs(2967) <= a;
    layer4_outputs(2968) <= '1';
    layer4_outputs(2969) <= not a or b;
    layer4_outputs(2970) <= b and not a;
    layer4_outputs(2971) <= a or b;
    layer4_outputs(2972) <= b and not a;
    layer4_outputs(2973) <= not a;
    layer4_outputs(2974) <= not b or a;
    layer4_outputs(2975) <= '0';
    layer4_outputs(2976) <= not (a or b);
    layer4_outputs(2977) <= '0';
    layer4_outputs(2978) <= not (a and b);
    layer4_outputs(2979) <= not (a xor b);
    layer4_outputs(2980) <= not b or a;
    layer4_outputs(2981) <= a or b;
    layer4_outputs(2982) <= not a or b;
    layer4_outputs(2983) <= '0';
    layer4_outputs(2984) <= b and not a;
    layer4_outputs(2985) <= not (a and b);
    layer4_outputs(2986) <= b;
    layer4_outputs(2987) <= '1';
    layer4_outputs(2988) <= '0';
    layer4_outputs(2989) <= '1';
    layer4_outputs(2990) <= a and not b;
    layer4_outputs(2991) <= a xor b;
    layer4_outputs(2992) <= a or b;
    layer4_outputs(2993) <= b and not a;
    layer4_outputs(2994) <= not b;
    layer4_outputs(2995) <= a and not b;
    layer4_outputs(2996) <= not b;
    layer4_outputs(2997) <= a xor b;
    layer4_outputs(2998) <= not a or b;
    layer4_outputs(2999) <= a;
    layer4_outputs(3000) <= a;
    layer4_outputs(3001) <= not a or b;
    layer4_outputs(3002) <= not b;
    layer4_outputs(3003) <= not (a or b);
    layer4_outputs(3004) <= not b or a;
    layer4_outputs(3005) <= '0';
    layer4_outputs(3006) <= a;
    layer4_outputs(3007) <= a and b;
    layer4_outputs(3008) <= not (a xor b);
    layer4_outputs(3009) <= not (a xor b);
    layer4_outputs(3010) <= a xor b;
    layer4_outputs(3011) <= '0';
    layer4_outputs(3012) <= not (a or b);
    layer4_outputs(3013) <= not a or b;
    layer4_outputs(3014) <= a and b;
    layer4_outputs(3015) <= not a;
    layer4_outputs(3016) <= not (a and b);
    layer4_outputs(3017) <= not (a or b);
    layer4_outputs(3018) <= not a or b;
    layer4_outputs(3019) <= not a;
    layer4_outputs(3020) <= b and not a;
    layer4_outputs(3021) <= not (a or b);
    layer4_outputs(3022) <= a or b;
    layer4_outputs(3023) <= not b;
    layer4_outputs(3024) <= not b;
    layer4_outputs(3025) <= a;
    layer4_outputs(3026) <= b;
    layer4_outputs(3027) <= a xor b;
    layer4_outputs(3028) <= a or b;
    layer4_outputs(3029) <= b;
    layer4_outputs(3030) <= not a or b;
    layer4_outputs(3031) <= a xor b;
    layer4_outputs(3032) <= not a;
    layer4_outputs(3033) <= not a;
    layer4_outputs(3034) <= not a or b;
    layer4_outputs(3035) <= b and not a;
    layer4_outputs(3036) <= not (a xor b);
    layer4_outputs(3037) <= not (a or b);
    layer4_outputs(3038) <= a and not b;
    layer4_outputs(3039) <= a or b;
    layer4_outputs(3040) <= not (a and b);
    layer4_outputs(3041) <= not a or b;
    layer4_outputs(3042) <= not a or b;
    layer4_outputs(3043) <= not a;
    layer4_outputs(3044) <= not b;
    layer4_outputs(3045) <= a or b;
    layer4_outputs(3046) <= not (a or b);
    layer4_outputs(3047) <= a;
    layer4_outputs(3048) <= not a or b;
    layer4_outputs(3049) <= not a or b;
    layer4_outputs(3050) <= a or b;
    layer4_outputs(3051) <= '0';
    layer4_outputs(3052) <= '0';
    layer4_outputs(3053) <= '0';
    layer4_outputs(3054) <= not b;
    layer4_outputs(3055) <= not a;
    layer4_outputs(3056) <= '0';
    layer4_outputs(3057) <= a;
    layer4_outputs(3058) <= not (a and b);
    layer4_outputs(3059) <= not b or a;
    layer4_outputs(3060) <= not a or b;
    layer4_outputs(3061) <= '1';
    layer4_outputs(3062) <= a and b;
    layer4_outputs(3063) <= '0';
    layer4_outputs(3064) <= '1';
    layer4_outputs(3065) <= not b or a;
    layer4_outputs(3066) <= b;
    layer4_outputs(3067) <= a or b;
    layer4_outputs(3068) <= a;
    layer4_outputs(3069) <= b;
    layer4_outputs(3070) <= '1';
    layer4_outputs(3071) <= a and b;
    layer4_outputs(3072) <= not (a or b);
    layer4_outputs(3073) <= a or b;
    layer4_outputs(3074) <= a and b;
    layer4_outputs(3075) <= a xor b;
    layer4_outputs(3076) <= b;
    layer4_outputs(3077) <= a;
    layer4_outputs(3078) <= a xor b;
    layer4_outputs(3079) <= a xor b;
    layer4_outputs(3080) <= a or b;
    layer4_outputs(3081) <= not b;
    layer4_outputs(3082) <= not (a and b);
    layer4_outputs(3083) <= a or b;
    layer4_outputs(3084) <= not b or a;
    layer4_outputs(3085) <= a;
    layer4_outputs(3086) <= not (a and b);
    layer4_outputs(3087) <= not a or b;
    layer4_outputs(3088) <= b;
    layer4_outputs(3089) <= not (a and b);
    layer4_outputs(3090) <= b;
    layer4_outputs(3091) <= b;
    layer4_outputs(3092) <= a and b;
    layer4_outputs(3093) <= not a or b;
    layer4_outputs(3094) <= not a or b;
    layer4_outputs(3095) <= b;
    layer4_outputs(3096) <= a;
    layer4_outputs(3097) <= a;
    layer4_outputs(3098) <= not b;
    layer4_outputs(3099) <= not b;
    layer4_outputs(3100) <= not (a xor b);
    layer4_outputs(3101) <= a;
    layer4_outputs(3102) <= b;
    layer4_outputs(3103) <= a and b;
    layer4_outputs(3104) <= b;
    layer4_outputs(3105) <= '1';
    layer4_outputs(3106) <= '0';
    layer4_outputs(3107) <= '1';
    layer4_outputs(3108) <= a and not b;
    layer4_outputs(3109) <= not a or b;
    layer4_outputs(3110) <= not a;
    layer4_outputs(3111) <= not (a or b);
    layer4_outputs(3112) <= not b or a;
    layer4_outputs(3113) <= not b;
    layer4_outputs(3114) <= b and not a;
    layer4_outputs(3115) <= '1';
    layer4_outputs(3116) <= a and b;
    layer4_outputs(3117) <= a;
    layer4_outputs(3118) <= not b or a;
    layer4_outputs(3119) <= a;
    layer4_outputs(3120) <= a or b;
    layer4_outputs(3121) <= a and not b;
    layer4_outputs(3122) <= a and not b;
    layer4_outputs(3123) <= a and b;
    layer4_outputs(3124) <= a or b;
    layer4_outputs(3125) <= '1';
    layer4_outputs(3126) <= not b or a;
    layer4_outputs(3127) <= '0';
    layer4_outputs(3128) <= not a or b;
    layer4_outputs(3129) <= not b;
    layer4_outputs(3130) <= not (a and b);
    layer4_outputs(3131) <= '1';
    layer4_outputs(3132) <= a;
    layer4_outputs(3133) <= a and not b;
    layer4_outputs(3134) <= a and not b;
    layer4_outputs(3135) <= not (a xor b);
    layer4_outputs(3136) <= b;
    layer4_outputs(3137) <= '0';
    layer4_outputs(3138) <= a or b;
    layer4_outputs(3139) <= b and not a;
    layer4_outputs(3140) <= a or b;
    layer4_outputs(3141) <= not b;
    layer4_outputs(3142) <= a and b;
    layer4_outputs(3143) <= a;
    layer4_outputs(3144) <= not b;
    layer4_outputs(3145) <= not (a xor b);
    layer4_outputs(3146) <= a and not b;
    layer4_outputs(3147) <= a or b;
    layer4_outputs(3148) <= b and not a;
    layer4_outputs(3149) <= b and not a;
    layer4_outputs(3150) <= a;
    layer4_outputs(3151) <= not (a or b);
    layer4_outputs(3152) <= a and b;
    layer4_outputs(3153) <= not b;
    layer4_outputs(3154) <= b;
    layer4_outputs(3155) <= not a;
    layer4_outputs(3156) <= not a;
    layer4_outputs(3157) <= not b;
    layer4_outputs(3158) <= not a;
    layer4_outputs(3159) <= b and not a;
    layer4_outputs(3160) <= b and not a;
    layer4_outputs(3161) <= b;
    layer4_outputs(3162) <= not a;
    layer4_outputs(3163) <= b and not a;
    layer4_outputs(3164) <= not (a or b);
    layer4_outputs(3165) <= not (a or b);
    layer4_outputs(3166) <= b and not a;
    layer4_outputs(3167) <= not b;
    layer4_outputs(3168) <= not (a or b);
    layer4_outputs(3169) <= a;
    layer4_outputs(3170) <= b and not a;
    layer4_outputs(3171) <= not (a and b);
    layer4_outputs(3172) <= a and b;
    layer4_outputs(3173) <= b and not a;
    layer4_outputs(3174) <= b and not a;
    layer4_outputs(3175) <= a or b;
    layer4_outputs(3176) <= a and not b;
    layer4_outputs(3177) <= a or b;
    layer4_outputs(3178) <= b;
    layer4_outputs(3179) <= a or b;
    layer4_outputs(3180) <= not (a or b);
    layer4_outputs(3181) <= a;
    layer4_outputs(3182) <= not a;
    layer4_outputs(3183) <= b;
    layer4_outputs(3184) <= not (a or b);
    layer4_outputs(3185) <= a and not b;
    layer4_outputs(3186) <= not a or b;
    layer4_outputs(3187) <= not (a or b);
    layer4_outputs(3188) <= not b or a;
    layer4_outputs(3189) <= a or b;
    layer4_outputs(3190) <= not a or b;
    layer4_outputs(3191) <= not b;
    layer4_outputs(3192) <= '1';
    layer4_outputs(3193) <= not b;
    layer4_outputs(3194) <= b;
    layer4_outputs(3195) <= not (a or b);
    layer4_outputs(3196) <= b;
    layer4_outputs(3197) <= '0';
    layer4_outputs(3198) <= a;
    layer4_outputs(3199) <= b and not a;
    layer4_outputs(3200) <= b and not a;
    layer4_outputs(3201) <= '1';
    layer4_outputs(3202) <= not a or b;
    layer4_outputs(3203) <= not b or a;
    layer4_outputs(3204) <= a and not b;
    layer4_outputs(3205) <= a and b;
    layer4_outputs(3206) <= not (a and b);
    layer4_outputs(3207) <= '0';
    layer4_outputs(3208) <= a or b;
    layer4_outputs(3209) <= not b or a;
    layer4_outputs(3210) <= not (a and b);
    layer4_outputs(3211) <= not (a or b);
    layer4_outputs(3212) <= a or b;
    layer4_outputs(3213) <= not b;
    layer4_outputs(3214) <= b;
    layer4_outputs(3215) <= not (a or b);
    layer4_outputs(3216) <= not (a or b);
    layer4_outputs(3217) <= not (a and b);
    layer4_outputs(3218) <= a or b;
    layer4_outputs(3219) <= a and b;
    layer4_outputs(3220) <= a and b;
    layer4_outputs(3221) <= b and not a;
    layer4_outputs(3222) <= '1';
    layer4_outputs(3223) <= a and b;
    layer4_outputs(3224) <= not a;
    layer4_outputs(3225) <= a and not b;
    layer4_outputs(3226) <= a or b;
    layer4_outputs(3227) <= a or b;
    layer4_outputs(3228) <= a or b;
    layer4_outputs(3229) <= a;
    layer4_outputs(3230) <= not b;
    layer4_outputs(3231) <= '1';
    layer4_outputs(3232) <= a and b;
    layer4_outputs(3233) <= not a;
    layer4_outputs(3234) <= not b or a;
    layer4_outputs(3235) <= b and not a;
    layer4_outputs(3236) <= b and not a;
    layer4_outputs(3237) <= not a;
    layer4_outputs(3238) <= not b;
    layer4_outputs(3239) <= b and not a;
    layer4_outputs(3240) <= '0';
    layer4_outputs(3241) <= b;
    layer4_outputs(3242) <= not b;
    layer4_outputs(3243) <= not (a or b);
    layer4_outputs(3244) <= not (a and b);
    layer4_outputs(3245) <= a;
    layer4_outputs(3246) <= a and b;
    layer4_outputs(3247) <= '1';
    layer4_outputs(3248) <= a and b;
    layer4_outputs(3249) <= not b;
    layer4_outputs(3250) <= not b;
    layer4_outputs(3251) <= a or b;
    layer4_outputs(3252) <= a or b;
    layer4_outputs(3253) <= not (a or b);
    layer4_outputs(3254) <= a and not b;
    layer4_outputs(3255) <= not a;
    layer4_outputs(3256) <= b;
    layer4_outputs(3257) <= '1';
    layer4_outputs(3258) <= a and b;
    layer4_outputs(3259) <= a or b;
    layer4_outputs(3260) <= a and b;
    layer4_outputs(3261) <= not b or a;
    layer4_outputs(3262) <= a or b;
    layer4_outputs(3263) <= a xor b;
    layer4_outputs(3264) <= not a or b;
    layer4_outputs(3265) <= not a or b;
    layer4_outputs(3266) <= '1';
    layer4_outputs(3267) <= b;
    layer4_outputs(3268) <= a;
    layer4_outputs(3269) <= a and b;
    layer4_outputs(3270) <= a;
    layer4_outputs(3271) <= a and b;
    layer4_outputs(3272) <= '0';
    layer4_outputs(3273) <= not b or a;
    layer4_outputs(3274) <= '1';
    layer4_outputs(3275) <= '0';
    layer4_outputs(3276) <= a;
    layer4_outputs(3277) <= a and b;
    layer4_outputs(3278) <= b and not a;
    layer4_outputs(3279) <= not b or a;
    layer4_outputs(3280) <= b;
    layer4_outputs(3281) <= not (a and b);
    layer4_outputs(3282) <= a;
    layer4_outputs(3283) <= not a;
    layer4_outputs(3284) <= not b or a;
    layer4_outputs(3285) <= not b or a;
    layer4_outputs(3286) <= not a or b;
    layer4_outputs(3287) <= b and not a;
    layer4_outputs(3288) <= '1';
    layer4_outputs(3289) <= a and b;
    layer4_outputs(3290) <= not (a and b);
    layer4_outputs(3291) <= not (a or b);
    layer4_outputs(3292) <= not a or b;
    layer4_outputs(3293) <= a and b;
    layer4_outputs(3294) <= a;
    layer4_outputs(3295) <= not b or a;
    layer4_outputs(3296) <= a and not b;
    layer4_outputs(3297) <= b and not a;
    layer4_outputs(3298) <= a;
    layer4_outputs(3299) <= a or b;
    layer4_outputs(3300) <= not a;
    layer4_outputs(3301) <= a;
    layer4_outputs(3302) <= not b;
    layer4_outputs(3303) <= not (a and b);
    layer4_outputs(3304) <= not a;
    layer4_outputs(3305) <= b and not a;
    layer4_outputs(3306) <= not b or a;
    layer4_outputs(3307) <= not b or a;
    layer4_outputs(3308) <= a and b;
    layer4_outputs(3309) <= b;
    layer4_outputs(3310) <= b and not a;
    layer4_outputs(3311) <= '1';
    layer4_outputs(3312) <= not (a or b);
    layer4_outputs(3313) <= not (a or b);
    layer4_outputs(3314) <= not (a or b);
    layer4_outputs(3315) <= '0';
    layer4_outputs(3316) <= a or b;
    layer4_outputs(3317) <= a;
    layer4_outputs(3318) <= b and not a;
    layer4_outputs(3319) <= not (a and b);
    layer4_outputs(3320) <= a and b;
    layer4_outputs(3321) <= a and not b;
    layer4_outputs(3322) <= not (a or b);
    layer4_outputs(3323) <= '1';
    layer4_outputs(3324) <= not b or a;
    layer4_outputs(3325) <= '1';
    layer4_outputs(3326) <= not (a xor b);
    layer4_outputs(3327) <= not a;
    layer4_outputs(3328) <= a and not b;
    layer4_outputs(3329) <= a and b;
    layer4_outputs(3330) <= a and b;
    layer4_outputs(3331) <= not (a and b);
    layer4_outputs(3332) <= not a;
    layer4_outputs(3333) <= not (a or b);
    layer4_outputs(3334) <= b;
    layer4_outputs(3335) <= not (a or b);
    layer4_outputs(3336) <= a and b;
    layer4_outputs(3337) <= '0';
    layer4_outputs(3338) <= not b or a;
    layer4_outputs(3339) <= a and b;
    layer4_outputs(3340) <= '1';
    layer4_outputs(3341) <= a and not b;
    layer4_outputs(3342) <= a;
    layer4_outputs(3343) <= not b;
    layer4_outputs(3344) <= not a;
    layer4_outputs(3345) <= b and not a;
    layer4_outputs(3346) <= not a or b;
    layer4_outputs(3347) <= '0';
    layer4_outputs(3348) <= a and not b;
    layer4_outputs(3349) <= not a or b;
    layer4_outputs(3350) <= not b;
    layer4_outputs(3351) <= a and not b;
    layer4_outputs(3352) <= not b or a;
    layer4_outputs(3353) <= not (a and b);
    layer4_outputs(3354) <= a and b;
    layer4_outputs(3355) <= a and b;
    layer4_outputs(3356) <= not a;
    layer4_outputs(3357) <= not a or b;
    layer4_outputs(3358) <= '0';
    layer4_outputs(3359) <= a and b;
    layer4_outputs(3360) <= not b or a;
    layer4_outputs(3361) <= '1';
    layer4_outputs(3362) <= a xor b;
    layer4_outputs(3363) <= b;
    layer4_outputs(3364) <= b;
    layer4_outputs(3365) <= b and not a;
    layer4_outputs(3366) <= not a;
    layer4_outputs(3367) <= not a;
    layer4_outputs(3368) <= a and not b;
    layer4_outputs(3369) <= not b or a;
    layer4_outputs(3370) <= not b or a;
    layer4_outputs(3371) <= not b or a;
    layer4_outputs(3372) <= a or b;
    layer4_outputs(3373) <= a or b;
    layer4_outputs(3374) <= b and not a;
    layer4_outputs(3375) <= b;
    layer4_outputs(3376) <= b and not a;
    layer4_outputs(3377) <= a or b;
    layer4_outputs(3378) <= not b;
    layer4_outputs(3379) <= a;
    layer4_outputs(3380) <= a or b;
    layer4_outputs(3381) <= not a;
    layer4_outputs(3382) <= a and b;
    layer4_outputs(3383) <= a and not b;
    layer4_outputs(3384) <= not (a and b);
    layer4_outputs(3385) <= b;
    layer4_outputs(3386) <= a;
    layer4_outputs(3387) <= a;
    layer4_outputs(3388) <= a and not b;
    layer4_outputs(3389) <= not b or a;
    layer4_outputs(3390) <= not (a or b);
    layer4_outputs(3391) <= b and not a;
    layer4_outputs(3392) <= a or b;
    layer4_outputs(3393) <= not (a or b);
    layer4_outputs(3394) <= '0';
    layer4_outputs(3395) <= a or b;
    layer4_outputs(3396) <= a and b;
    layer4_outputs(3397) <= not a or b;
    layer4_outputs(3398) <= a and b;
    layer4_outputs(3399) <= not b or a;
    layer4_outputs(3400) <= a or b;
    layer4_outputs(3401) <= '0';
    layer4_outputs(3402) <= a or b;
    layer4_outputs(3403) <= a;
    layer4_outputs(3404) <= a;
    layer4_outputs(3405) <= not (a or b);
    layer4_outputs(3406) <= b;
    layer4_outputs(3407) <= not b;
    layer4_outputs(3408) <= '1';
    layer4_outputs(3409) <= not a;
    layer4_outputs(3410) <= not b or a;
    layer4_outputs(3411) <= not b or a;
    layer4_outputs(3412) <= not (a or b);
    layer4_outputs(3413) <= a and not b;
    layer4_outputs(3414) <= a and b;
    layer4_outputs(3415) <= a and not b;
    layer4_outputs(3416) <= a or b;
    layer4_outputs(3417) <= '0';
    layer4_outputs(3418) <= b;
    layer4_outputs(3419) <= a and not b;
    layer4_outputs(3420) <= not b;
    layer4_outputs(3421) <= a or b;
    layer4_outputs(3422) <= a;
    layer4_outputs(3423) <= a and b;
    layer4_outputs(3424) <= a or b;
    layer4_outputs(3425) <= a;
    layer4_outputs(3426) <= not b;
    layer4_outputs(3427) <= a;
    layer4_outputs(3428) <= not b;
    layer4_outputs(3429) <= a and not b;
    layer4_outputs(3430) <= not (a or b);
    layer4_outputs(3431) <= not (a or b);
    layer4_outputs(3432) <= not b or a;
    layer4_outputs(3433) <= not a or b;
    layer4_outputs(3434) <= a;
    layer4_outputs(3435) <= not b or a;
    layer4_outputs(3436) <= '1';
    layer4_outputs(3437) <= '0';
    layer4_outputs(3438) <= '0';
    layer4_outputs(3439) <= not b;
    layer4_outputs(3440) <= not (a and b);
    layer4_outputs(3441) <= a and not b;
    layer4_outputs(3442) <= b and not a;
    layer4_outputs(3443) <= a or b;
    layer4_outputs(3444) <= a;
    layer4_outputs(3445) <= '1';
    layer4_outputs(3446) <= not (a or b);
    layer4_outputs(3447) <= not a;
    layer4_outputs(3448) <= not a or b;
    layer4_outputs(3449) <= not a;
    layer4_outputs(3450) <= not a;
    layer4_outputs(3451) <= not (a xor b);
    layer4_outputs(3452) <= '0';
    layer4_outputs(3453) <= b;
    layer4_outputs(3454) <= a and not b;
    layer4_outputs(3455) <= not a;
    layer4_outputs(3456) <= b and not a;
    layer4_outputs(3457) <= '0';
    layer4_outputs(3458) <= not b;
    layer4_outputs(3459) <= not b;
    layer4_outputs(3460) <= not a;
    layer4_outputs(3461) <= b and not a;
    layer4_outputs(3462) <= a;
    layer4_outputs(3463) <= not (a or b);
    layer4_outputs(3464) <= not a or b;
    layer4_outputs(3465) <= b;
    layer4_outputs(3466) <= a;
    layer4_outputs(3467) <= a;
    layer4_outputs(3468) <= not a or b;
    layer4_outputs(3469) <= a;
    layer4_outputs(3470) <= '0';
    layer4_outputs(3471) <= a or b;
    layer4_outputs(3472) <= not (a and b);
    layer4_outputs(3473) <= a;
    layer4_outputs(3474) <= '0';
    layer4_outputs(3475) <= a and not b;
    layer4_outputs(3476) <= not a;
    layer4_outputs(3477) <= a and not b;
    layer4_outputs(3478) <= not b or a;
    layer4_outputs(3479) <= a xor b;
    layer4_outputs(3480) <= b and not a;
    layer4_outputs(3481) <= a or b;
    layer4_outputs(3482) <= not a or b;
    layer4_outputs(3483) <= not (a or b);
    layer4_outputs(3484) <= a and not b;
    layer4_outputs(3485) <= b and not a;
    layer4_outputs(3486) <= a and b;
    layer4_outputs(3487) <= a;
    layer4_outputs(3488) <= '1';
    layer4_outputs(3489) <= a or b;
    layer4_outputs(3490) <= a and b;
    layer4_outputs(3491) <= a and not b;
    layer4_outputs(3492) <= not a;
    layer4_outputs(3493) <= not (a or b);
    layer4_outputs(3494) <= a and not b;
    layer4_outputs(3495) <= a and b;
    layer4_outputs(3496) <= '1';
    layer4_outputs(3497) <= not a or b;
    layer4_outputs(3498) <= '1';
    layer4_outputs(3499) <= not b;
    layer4_outputs(3500) <= a xor b;
    layer4_outputs(3501) <= not b;
    layer4_outputs(3502) <= not (a or b);
    layer4_outputs(3503) <= '1';
    layer4_outputs(3504) <= a;
    layer4_outputs(3505) <= not b or a;
    layer4_outputs(3506) <= b and not a;
    layer4_outputs(3507) <= a;
    layer4_outputs(3508) <= not b or a;
    layer4_outputs(3509) <= b and not a;
    layer4_outputs(3510) <= not a;
    layer4_outputs(3511) <= a and not b;
    layer4_outputs(3512) <= b;
    layer4_outputs(3513) <= not b or a;
    layer4_outputs(3514) <= a;
    layer4_outputs(3515) <= b and not a;
    layer4_outputs(3516) <= a and b;
    layer4_outputs(3517) <= not a or b;
    layer4_outputs(3518) <= b and not a;
    layer4_outputs(3519) <= not b;
    layer4_outputs(3520) <= a and not b;
    layer4_outputs(3521) <= b;
    layer4_outputs(3522) <= not b;
    layer4_outputs(3523) <= not b;
    layer4_outputs(3524) <= not a;
    layer4_outputs(3525) <= a or b;
    layer4_outputs(3526) <= '0';
    layer4_outputs(3527) <= not (a or b);
    layer4_outputs(3528) <= a;
    layer4_outputs(3529) <= not a;
    layer4_outputs(3530) <= a and not b;
    layer4_outputs(3531) <= '0';
    layer4_outputs(3532) <= not a;
    layer4_outputs(3533) <= not (a or b);
    layer4_outputs(3534) <= b and not a;
    layer4_outputs(3535) <= a and not b;
    layer4_outputs(3536) <= a;
    layer4_outputs(3537) <= not (a xor b);
    layer4_outputs(3538) <= not a or b;
    layer4_outputs(3539) <= not a or b;
    layer4_outputs(3540) <= not (a xor b);
    layer4_outputs(3541) <= not (a and b);
    layer4_outputs(3542) <= b and not a;
    layer4_outputs(3543) <= a or b;
    layer4_outputs(3544) <= not (a or b);
    layer4_outputs(3545) <= not (a or b);
    layer4_outputs(3546) <= b;
    layer4_outputs(3547) <= a and b;
    layer4_outputs(3548) <= not (a and b);
    layer4_outputs(3549) <= not b or a;
    layer4_outputs(3550) <= not b or a;
    layer4_outputs(3551) <= not a or b;
    layer4_outputs(3552) <= not b;
    layer4_outputs(3553) <= b;
    layer4_outputs(3554) <= not (a xor b);
    layer4_outputs(3555) <= a and not b;
    layer4_outputs(3556) <= a or b;
    layer4_outputs(3557) <= not (a and b);
    layer4_outputs(3558) <= a;
    layer4_outputs(3559) <= '0';
    layer4_outputs(3560) <= '0';
    layer4_outputs(3561) <= b and not a;
    layer4_outputs(3562) <= not b;
    layer4_outputs(3563) <= a;
    layer4_outputs(3564) <= b;
    layer4_outputs(3565) <= not b;
    layer4_outputs(3566) <= not (a or b);
    layer4_outputs(3567) <= a xor b;
    layer4_outputs(3568) <= not a;
    layer4_outputs(3569) <= a;
    layer4_outputs(3570) <= not (a or b);
    layer4_outputs(3571) <= not a;
    layer4_outputs(3572) <= b and not a;
    layer4_outputs(3573) <= not a;
    layer4_outputs(3574) <= a;
    layer4_outputs(3575) <= a and not b;
    layer4_outputs(3576) <= not a;
    layer4_outputs(3577) <= b and not a;
    layer4_outputs(3578) <= not b;
    layer4_outputs(3579) <= not (a and b);
    layer4_outputs(3580) <= not (a xor b);
    layer4_outputs(3581) <= '0';
    layer4_outputs(3582) <= '0';
    layer4_outputs(3583) <= not b or a;
    layer4_outputs(3584) <= not b;
    layer4_outputs(3585) <= not b or a;
    layer4_outputs(3586) <= not (a and b);
    layer4_outputs(3587) <= '0';
    layer4_outputs(3588) <= not a or b;
    layer4_outputs(3589) <= not (a xor b);
    layer4_outputs(3590) <= not b;
    layer4_outputs(3591) <= not (a or b);
    layer4_outputs(3592) <= a;
    layer4_outputs(3593) <= a;
    layer4_outputs(3594) <= not b;
    layer4_outputs(3595) <= not b or a;
    layer4_outputs(3596) <= b and not a;
    layer4_outputs(3597) <= not a;
    layer4_outputs(3598) <= '1';
    layer4_outputs(3599) <= b;
    layer4_outputs(3600) <= not a or b;
    layer4_outputs(3601) <= not b or a;
    layer4_outputs(3602) <= not (a or b);
    layer4_outputs(3603) <= a xor b;
    layer4_outputs(3604) <= '1';
    layer4_outputs(3605) <= a xor b;
    layer4_outputs(3606) <= not (a and b);
    layer4_outputs(3607) <= '1';
    layer4_outputs(3608) <= not (a xor b);
    layer4_outputs(3609) <= a;
    layer4_outputs(3610) <= not a;
    layer4_outputs(3611) <= '1';
    layer4_outputs(3612) <= not a or b;
    layer4_outputs(3613) <= not a or b;
    layer4_outputs(3614) <= not (a xor b);
    layer4_outputs(3615) <= a and not b;
    layer4_outputs(3616) <= not (a xor b);
    layer4_outputs(3617) <= not (a xor b);
    layer4_outputs(3618) <= '1';
    layer4_outputs(3619) <= b;
    layer4_outputs(3620) <= a or b;
    layer4_outputs(3621) <= not a;
    layer4_outputs(3622) <= b and not a;
    layer4_outputs(3623) <= '1';
    layer4_outputs(3624) <= a and not b;
    layer4_outputs(3625) <= '0';
    layer4_outputs(3626) <= not a;
    layer4_outputs(3627) <= a and not b;
    layer4_outputs(3628) <= not (a or b);
    layer4_outputs(3629) <= not a;
    layer4_outputs(3630) <= not a or b;
    layer4_outputs(3631) <= '1';
    layer4_outputs(3632) <= b;
    layer4_outputs(3633) <= not (a or b);
    layer4_outputs(3634) <= a and not b;
    layer4_outputs(3635) <= not (a and b);
    layer4_outputs(3636) <= '1';
    layer4_outputs(3637) <= b;
    layer4_outputs(3638) <= not a;
    layer4_outputs(3639) <= a and not b;
    layer4_outputs(3640) <= a;
    layer4_outputs(3641) <= a and not b;
    layer4_outputs(3642) <= not (a or b);
    layer4_outputs(3643) <= not b or a;
    layer4_outputs(3644) <= not (a xor b);
    layer4_outputs(3645) <= not b or a;
    layer4_outputs(3646) <= not a;
    layer4_outputs(3647) <= '0';
    layer4_outputs(3648) <= a;
    layer4_outputs(3649) <= not b or a;
    layer4_outputs(3650) <= b;
    layer4_outputs(3651) <= not a;
    layer4_outputs(3652) <= b and not a;
    layer4_outputs(3653) <= not a or b;
    layer4_outputs(3654) <= not a or b;
    layer4_outputs(3655) <= not b or a;
    layer4_outputs(3656) <= a or b;
    layer4_outputs(3657) <= b and not a;
    layer4_outputs(3658) <= b;
    layer4_outputs(3659) <= not (a or b);
    layer4_outputs(3660) <= a and not b;
    layer4_outputs(3661) <= b;
    layer4_outputs(3662) <= b and not a;
    layer4_outputs(3663) <= not (a xor b);
    layer4_outputs(3664) <= a and b;
    layer4_outputs(3665) <= b and not a;
    layer4_outputs(3666) <= b;
    layer4_outputs(3667) <= not (a or b);
    layer4_outputs(3668) <= not b;
    layer4_outputs(3669) <= not b or a;
    layer4_outputs(3670) <= b and not a;
    layer4_outputs(3671) <= a and b;
    layer4_outputs(3672) <= not (a or b);
    layer4_outputs(3673) <= b;
    layer4_outputs(3674) <= a or b;
    layer4_outputs(3675) <= not b;
    layer4_outputs(3676) <= '0';
    layer4_outputs(3677) <= not b;
    layer4_outputs(3678) <= a and not b;
    layer4_outputs(3679) <= not a or b;
    layer4_outputs(3680) <= not a or b;
    layer4_outputs(3681) <= '1';
    layer4_outputs(3682) <= a or b;
    layer4_outputs(3683) <= b;
    layer4_outputs(3684) <= a or b;
    layer4_outputs(3685) <= '1';
    layer4_outputs(3686) <= not a;
    layer4_outputs(3687) <= b and not a;
    layer4_outputs(3688) <= a;
    layer4_outputs(3689) <= a or b;
    layer4_outputs(3690) <= a;
    layer4_outputs(3691) <= not a or b;
    layer4_outputs(3692) <= not a or b;
    layer4_outputs(3693) <= a;
    layer4_outputs(3694) <= not (a and b);
    layer4_outputs(3695) <= b;
    layer4_outputs(3696) <= a or b;
    layer4_outputs(3697) <= a or b;
    layer4_outputs(3698) <= not a;
    layer4_outputs(3699) <= '0';
    layer4_outputs(3700) <= '0';
    layer4_outputs(3701) <= not (a or b);
    layer4_outputs(3702) <= not a or b;
    layer4_outputs(3703) <= not b;
    layer4_outputs(3704) <= a and not b;
    layer4_outputs(3705) <= '1';
    layer4_outputs(3706) <= not (a or b);
    layer4_outputs(3707) <= a;
    layer4_outputs(3708) <= not b or a;
    layer4_outputs(3709) <= b and not a;
    layer4_outputs(3710) <= not (a and b);
    layer4_outputs(3711) <= not (a or b);
    layer4_outputs(3712) <= a;
    layer4_outputs(3713) <= a and not b;
    layer4_outputs(3714) <= '1';
    layer4_outputs(3715) <= not (a or b);
    layer4_outputs(3716) <= not b or a;
    layer4_outputs(3717) <= not b or a;
    layer4_outputs(3718) <= a;
    layer4_outputs(3719) <= not a;
    layer4_outputs(3720) <= a or b;
    layer4_outputs(3721) <= '1';
    layer4_outputs(3722) <= a;
    layer4_outputs(3723) <= not b or a;
    layer4_outputs(3724) <= b;
    layer4_outputs(3725) <= '1';
    layer4_outputs(3726) <= b;
    layer4_outputs(3727) <= not a;
    layer4_outputs(3728) <= '1';
    layer4_outputs(3729) <= b and not a;
    layer4_outputs(3730) <= '1';
    layer4_outputs(3731) <= not b or a;
    layer4_outputs(3732) <= a and not b;
    layer4_outputs(3733) <= b and not a;
    layer4_outputs(3734) <= not (a or b);
    layer4_outputs(3735) <= a and not b;
    layer4_outputs(3736) <= a;
    layer4_outputs(3737) <= a;
    layer4_outputs(3738) <= '0';
    layer4_outputs(3739) <= not a;
    layer4_outputs(3740) <= not a;
    layer4_outputs(3741) <= '1';
    layer4_outputs(3742) <= a or b;
    layer4_outputs(3743) <= not (a and b);
    layer4_outputs(3744) <= not a or b;
    layer4_outputs(3745) <= not b or a;
    layer4_outputs(3746) <= not a or b;
    layer4_outputs(3747) <= '0';
    layer4_outputs(3748) <= not (a or b);
    layer4_outputs(3749) <= a or b;
    layer4_outputs(3750) <= not b or a;
    layer4_outputs(3751) <= not b;
    layer4_outputs(3752) <= not (a or b);
    layer4_outputs(3753) <= not b or a;
    layer4_outputs(3754) <= a;
    layer4_outputs(3755) <= a;
    layer4_outputs(3756) <= b and not a;
    layer4_outputs(3757) <= a or b;
    layer4_outputs(3758) <= not a or b;
    layer4_outputs(3759) <= not b;
    layer4_outputs(3760) <= a and not b;
    layer4_outputs(3761) <= b;
    layer4_outputs(3762) <= b;
    layer4_outputs(3763) <= not a or b;
    layer4_outputs(3764) <= '1';
    layer4_outputs(3765) <= b;
    layer4_outputs(3766) <= b;
    layer4_outputs(3767) <= not b;
    layer4_outputs(3768) <= not b;
    layer4_outputs(3769) <= b and not a;
    layer4_outputs(3770) <= a xor b;
    layer4_outputs(3771) <= not b;
    layer4_outputs(3772) <= b and not a;
    layer4_outputs(3773) <= a and not b;
    layer4_outputs(3774) <= not a;
    layer4_outputs(3775) <= a;
    layer4_outputs(3776) <= not a;
    layer4_outputs(3777) <= not (a or b);
    layer4_outputs(3778) <= a and not b;
    layer4_outputs(3779) <= b;
    layer4_outputs(3780) <= b;
    layer4_outputs(3781) <= not a;
    layer4_outputs(3782) <= b;
    layer4_outputs(3783) <= not (a and b);
    layer4_outputs(3784) <= not b;
    layer4_outputs(3785) <= not (a or b);
    layer4_outputs(3786) <= b and not a;
    layer4_outputs(3787) <= not (a and b);
    layer4_outputs(3788) <= not (a and b);
    layer4_outputs(3789) <= not (a or b);
    layer4_outputs(3790) <= not b or a;
    layer4_outputs(3791) <= not (a or b);
    layer4_outputs(3792) <= not (a or b);
    layer4_outputs(3793) <= '1';
    layer4_outputs(3794) <= not (a and b);
    layer4_outputs(3795) <= '0';
    layer4_outputs(3796) <= a or b;
    layer4_outputs(3797) <= a and b;
    layer4_outputs(3798) <= a;
    layer4_outputs(3799) <= not (a or b);
    layer4_outputs(3800) <= '1';
    layer4_outputs(3801) <= a and not b;
    layer4_outputs(3802) <= b;
    layer4_outputs(3803) <= not (a or b);
    layer4_outputs(3804) <= not (a or b);
    layer4_outputs(3805) <= not a;
    layer4_outputs(3806) <= b and not a;
    layer4_outputs(3807) <= not b;
    layer4_outputs(3808) <= '1';
    layer4_outputs(3809) <= not a or b;
    layer4_outputs(3810) <= not a or b;
    layer4_outputs(3811) <= not b or a;
    layer4_outputs(3812) <= not b;
    layer4_outputs(3813) <= not b;
    layer4_outputs(3814) <= not b;
    layer4_outputs(3815) <= not b or a;
    layer4_outputs(3816) <= '0';
    layer4_outputs(3817) <= not b;
    layer4_outputs(3818) <= not b or a;
    layer4_outputs(3819) <= b and not a;
    layer4_outputs(3820) <= not (a xor b);
    layer4_outputs(3821) <= a and b;
    layer4_outputs(3822) <= b;
    layer4_outputs(3823) <= b;
    layer4_outputs(3824) <= b and not a;
    layer4_outputs(3825) <= b and not a;
    layer4_outputs(3826) <= not a;
    layer4_outputs(3827) <= not (a xor b);
    layer4_outputs(3828) <= a and b;
    layer4_outputs(3829) <= a or b;
    layer4_outputs(3830) <= not a or b;
    layer4_outputs(3831) <= '0';
    layer4_outputs(3832) <= a;
    layer4_outputs(3833) <= a or b;
    layer4_outputs(3834) <= not b;
    layer4_outputs(3835) <= not (a or b);
    layer4_outputs(3836) <= a;
    layer4_outputs(3837) <= a and not b;
    layer4_outputs(3838) <= not (a and b);
    layer4_outputs(3839) <= a xor b;
    layer4_outputs(3840) <= not b;
    layer4_outputs(3841) <= not a;
    layer4_outputs(3842) <= not (a or b);
    layer4_outputs(3843) <= not b;
    layer4_outputs(3844) <= not b or a;
    layer4_outputs(3845) <= '0';
    layer4_outputs(3846) <= b and not a;
    layer4_outputs(3847) <= not a;
    layer4_outputs(3848) <= not (a or b);
    layer4_outputs(3849) <= b;
    layer4_outputs(3850) <= a and not b;
    layer4_outputs(3851) <= not (a and b);
    layer4_outputs(3852) <= a or b;
    layer4_outputs(3853) <= not b;
    layer4_outputs(3854) <= a;
    layer4_outputs(3855) <= not (a or b);
    layer4_outputs(3856) <= '1';
    layer4_outputs(3857) <= '0';
    layer4_outputs(3858) <= not (a and b);
    layer4_outputs(3859) <= a and b;
    layer4_outputs(3860) <= not b or a;
    layer4_outputs(3861) <= not b;
    layer4_outputs(3862) <= not (a xor b);
    layer4_outputs(3863) <= not b or a;
    layer4_outputs(3864) <= a and b;
    layer4_outputs(3865) <= b;
    layer4_outputs(3866) <= a;
    layer4_outputs(3867) <= b;
    layer4_outputs(3868) <= a and b;
    layer4_outputs(3869) <= a or b;
    layer4_outputs(3870) <= b and not a;
    layer4_outputs(3871) <= not b or a;
    layer4_outputs(3872) <= not (a or b);
    layer4_outputs(3873) <= not b or a;
    layer4_outputs(3874) <= b and not a;
    layer4_outputs(3875) <= not (a or b);
    layer4_outputs(3876) <= not b or a;
    layer4_outputs(3877) <= not (a or b);
    layer4_outputs(3878) <= a or b;
    layer4_outputs(3879) <= a or b;
    layer4_outputs(3880) <= not (a xor b);
    layer4_outputs(3881) <= a;
    layer4_outputs(3882) <= a and not b;
    layer4_outputs(3883) <= a;
    layer4_outputs(3884) <= b and not a;
    layer4_outputs(3885) <= not a or b;
    layer4_outputs(3886) <= '1';
    layer4_outputs(3887) <= not a or b;
    layer4_outputs(3888) <= a;
    layer4_outputs(3889) <= not (a xor b);
    layer4_outputs(3890) <= a xor b;
    layer4_outputs(3891) <= not (a and b);
    layer4_outputs(3892) <= not b or a;
    layer4_outputs(3893) <= a;
    layer4_outputs(3894) <= not (a xor b);
    layer4_outputs(3895) <= a;
    layer4_outputs(3896) <= a and b;
    layer4_outputs(3897) <= a and b;
    layer4_outputs(3898) <= a and b;
    layer4_outputs(3899) <= a or b;
    layer4_outputs(3900) <= '0';
    layer4_outputs(3901) <= '1';
    layer4_outputs(3902) <= '0';
    layer4_outputs(3903) <= not (a and b);
    layer4_outputs(3904) <= not (a and b);
    layer4_outputs(3905) <= not b;
    layer4_outputs(3906) <= a or b;
    layer4_outputs(3907) <= a or b;
    layer4_outputs(3908) <= not (a or b);
    layer4_outputs(3909) <= b;
    layer4_outputs(3910) <= not b or a;
    layer4_outputs(3911) <= '1';
    layer4_outputs(3912) <= a or b;
    layer4_outputs(3913) <= a or b;
    layer4_outputs(3914) <= not b;
    layer4_outputs(3915) <= a and b;
    layer4_outputs(3916) <= not a or b;
    layer4_outputs(3917) <= not a;
    layer4_outputs(3918) <= not b;
    layer4_outputs(3919) <= a;
    layer4_outputs(3920) <= not a;
    layer4_outputs(3921) <= not a;
    layer4_outputs(3922) <= not (a or b);
    layer4_outputs(3923) <= a;
    layer4_outputs(3924) <= not b or a;
    layer4_outputs(3925) <= not (a or b);
    layer4_outputs(3926) <= '1';
    layer4_outputs(3927) <= not (a or b);
    layer4_outputs(3928) <= a;
    layer4_outputs(3929) <= not (a or b);
    layer4_outputs(3930) <= b;
    layer4_outputs(3931) <= '1';
    layer4_outputs(3932) <= not b or a;
    layer4_outputs(3933) <= a xor b;
    layer4_outputs(3934) <= b;
    layer4_outputs(3935) <= not b;
    layer4_outputs(3936) <= b;
    layer4_outputs(3937) <= b;
    layer4_outputs(3938) <= not a;
    layer4_outputs(3939) <= '1';
    layer4_outputs(3940) <= not a;
    layer4_outputs(3941) <= not (a and b);
    layer4_outputs(3942) <= not (a xor b);
    layer4_outputs(3943) <= not b or a;
    layer4_outputs(3944) <= not a or b;
    layer4_outputs(3945) <= not (a and b);
    layer4_outputs(3946) <= not b or a;
    layer4_outputs(3947) <= not (a and b);
    layer4_outputs(3948) <= a;
    layer4_outputs(3949) <= not b;
    layer4_outputs(3950) <= '0';
    layer4_outputs(3951) <= b;
    layer4_outputs(3952) <= a;
    layer4_outputs(3953) <= not (a or b);
    layer4_outputs(3954) <= b and not a;
    layer4_outputs(3955) <= a or b;
    layer4_outputs(3956) <= not (a and b);
    layer4_outputs(3957) <= b;
    layer4_outputs(3958) <= a and not b;
    layer4_outputs(3959) <= a or b;
    layer4_outputs(3960) <= not a or b;
    layer4_outputs(3961) <= not a;
    layer4_outputs(3962) <= a;
    layer4_outputs(3963) <= a and b;
    layer4_outputs(3964) <= '1';
    layer4_outputs(3965) <= a and not b;
    layer4_outputs(3966) <= not (a xor b);
    layer4_outputs(3967) <= not (a xor b);
    layer4_outputs(3968) <= not (a or b);
    layer4_outputs(3969) <= a or b;
    layer4_outputs(3970) <= not (a or b);
    layer4_outputs(3971) <= b and not a;
    layer4_outputs(3972) <= a and b;
    layer4_outputs(3973) <= not (a or b);
    layer4_outputs(3974) <= a;
    layer4_outputs(3975) <= not a or b;
    layer4_outputs(3976) <= not a or b;
    layer4_outputs(3977) <= a and not b;
    layer4_outputs(3978) <= a xor b;
    layer4_outputs(3979) <= a and not b;
    layer4_outputs(3980) <= b;
    layer4_outputs(3981) <= not b;
    layer4_outputs(3982) <= not (a and b);
    layer4_outputs(3983) <= not a or b;
    layer4_outputs(3984) <= not (a and b);
    layer4_outputs(3985) <= '0';
    layer4_outputs(3986) <= b and not a;
    layer4_outputs(3987) <= b;
    layer4_outputs(3988) <= a;
    layer4_outputs(3989) <= not a;
    layer4_outputs(3990) <= b;
    layer4_outputs(3991) <= not (a and b);
    layer4_outputs(3992) <= not b;
    layer4_outputs(3993) <= '0';
    layer4_outputs(3994) <= not (a and b);
    layer4_outputs(3995) <= a and not b;
    layer4_outputs(3996) <= b;
    layer4_outputs(3997) <= not (a or b);
    layer4_outputs(3998) <= not a;
    layer4_outputs(3999) <= a or b;
    layer4_outputs(4000) <= b and not a;
    layer4_outputs(4001) <= not a;
    layer4_outputs(4002) <= not a;
    layer4_outputs(4003) <= b;
    layer4_outputs(4004) <= b;
    layer4_outputs(4005) <= b and not a;
    layer4_outputs(4006) <= a;
    layer4_outputs(4007) <= not b or a;
    layer4_outputs(4008) <= a and not b;
    layer4_outputs(4009) <= not a or b;
    layer4_outputs(4010) <= '1';
    layer4_outputs(4011) <= not b;
    layer4_outputs(4012) <= a;
    layer4_outputs(4013) <= b;
    layer4_outputs(4014) <= not (a xor b);
    layer4_outputs(4015) <= not a or b;
    layer4_outputs(4016) <= not (a or b);
    layer4_outputs(4017) <= a xor b;
    layer4_outputs(4018) <= not b or a;
    layer4_outputs(4019) <= a and b;
    layer4_outputs(4020) <= not b;
    layer4_outputs(4021) <= not a or b;
    layer4_outputs(4022) <= not (a and b);
    layer4_outputs(4023) <= a;
    layer4_outputs(4024) <= not b or a;
    layer4_outputs(4025) <= a or b;
    layer4_outputs(4026) <= a or b;
    layer4_outputs(4027) <= not b or a;
    layer4_outputs(4028) <= not a;
    layer4_outputs(4029) <= not b;
    layer4_outputs(4030) <= a and not b;
    layer4_outputs(4031) <= a and not b;
    layer4_outputs(4032) <= not b or a;
    layer4_outputs(4033) <= not a or b;
    layer4_outputs(4034) <= not b;
    layer4_outputs(4035) <= not (a xor b);
    layer4_outputs(4036) <= b;
    layer4_outputs(4037) <= '1';
    layer4_outputs(4038) <= a and not b;
    layer4_outputs(4039) <= not (a xor b);
    layer4_outputs(4040) <= not (a and b);
    layer4_outputs(4041) <= a;
    layer4_outputs(4042) <= not a;
    layer4_outputs(4043) <= b;
    layer4_outputs(4044) <= a or b;
    layer4_outputs(4045) <= not b;
    layer4_outputs(4046) <= a and not b;
    layer4_outputs(4047) <= not a;
    layer4_outputs(4048) <= a and b;
    layer4_outputs(4049) <= a or b;
    layer4_outputs(4050) <= not (a or b);
    layer4_outputs(4051) <= not (a and b);
    layer4_outputs(4052) <= '0';
    layer4_outputs(4053) <= a or b;
    layer4_outputs(4054) <= '1';
    layer4_outputs(4055) <= a;
    layer4_outputs(4056) <= not b;
    layer4_outputs(4057) <= not (a or b);
    layer4_outputs(4058) <= not a;
    layer4_outputs(4059) <= '1';
    layer4_outputs(4060) <= a;
    layer4_outputs(4061) <= a and b;
    layer4_outputs(4062) <= a;
    layer4_outputs(4063) <= not (a and b);
    layer4_outputs(4064) <= a xor b;
    layer4_outputs(4065) <= '1';
    layer4_outputs(4066) <= b and not a;
    layer4_outputs(4067) <= not b or a;
    layer4_outputs(4068) <= not (a or b);
    layer4_outputs(4069) <= not (a and b);
    layer4_outputs(4070) <= not a;
    layer4_outputs(4071) <= a and not b;
    layer4_outputs(4072) <= not a or b;
    layer4_outputs(4073) <= b and not a;
    layer4_outputs(4074) <= b;
    layer4_outputs(4075) <= not (a or b);
    layer4_outputs(4076) <= a;
    layer4_outputs(4077) <= not b or a;
    layer4_outputs(4078) <= a and not b;
    layer4_outputs(4079) <= a;
    layer4_outputs(4080) <= a and b;
    layer4_outputs(4081) <= not b;
    layer4_outputs(4082) <= not (a or b);
    layer4_outputs(4083) <= b and not a;
    layer4_outputs(4084) <= '0';
    layer4_outputs(4085) <= not a;
    layer4_outputs(4086) <= a;
    layer4_outputs(4087) <= not (a or b);
    layer4_outputs(4088) <= a and b;
    layer4_outputs(4089) <= a;
    layer4_outputs(4090) <= b and not a;
    layer4_outputs(4091) <= '0';
    layer4_outputs(4092) <= not a or b;
    layer4_outputs(4093) <= b;
    layer4_outputs(4094) <= b;
    layer4_outputs(4095) <= a and not b;
    layer4_outputs(4096) <= not a;
    layer4_outputs(4097) <= not a;
    layer4_outputs(4098) <= not b or a;
    layer4_outputs(4099) <= a and b;
    layer4_outputs(4100) <= not (a or b);
    layer4_outputs(4101) <= not a or b;
    layer4_outputs(4102) <= not (a and b);
    layer4_outputs(4103) <= a and not b;
    layer4_outputs(4104) <= not (a and b);
    layer4_outputs(4105) <= a or b;
    layer4_outputs(4106) <= a and b;
    layer4_outputs(4107) <= '0';
    layer4_outputs(4108) <= not a;
    layer4_outputs(4109) <= not b or a;
    layer4_outputs(4110) <= '0';
    layer4_outputs(4111) <= not b;
    layer4_outputs(4112) <= not (a or b);
    layer4_outputs(4113) <= a;
    layer4_outputs(4114) <= a and not b;
    layer4_outputs(4115) <= b;
    layer4_outputs(4116) <= '1';
    layer4_outputs(4117) <= a and not b;
    layer4_outputs(4118) <= a and not b;
    layer4_outputs(4119) <= b and not a;
    layer4_outputs(4120) <= not (a and b);
    layer4_outputs(4121) <= not (a xor b);
    layer4_outputs(4122) <= a and b;
    layer4_outputs(4123) <= not a or b;
    layer4_outputs(4124) <= not b;
    layer4_outputs(4125) <= not a or b;
    layer4_outputs(4126) <= not a or b;
    layer4_outputs(4127) <= a;
    layer4_outputs(4128) <= not b;
    layer4_outputs(4129) <= '1';
    layer4_outputs(4130) <= not b or a;
    layer4_outputs(4131) <= a and b;
    layer4_outputs(4132) <= '1';
    layer4_outputs(4133) <= a and not b;
    layer4_outputs(4134) <= b and not a;
    layer4_outputs(4135) <= a and not b;
    layer4_outputs(4136) <= '0';
    layer4_outputs(4137) <= not a or b;
    layer4_outputs(4138) <= not b or a;
    layer4_outputs(4139) <= not (a and b);
    layer4_outputs(4140) <= a or b;
    layer4_outputs(4141) <= not (a and b);
    layer4_outputs(4142) <= not a;
    layer4_outputs(4143) <= not (a or b);
    layer4_outputs(4144) <= a xor b;
    layer4_outputs(4145) <= not a;
    layer4_outputs(4146) <= a xor b;
    layer4_outputs(4147) <= a xor b;
    layer4_outputs(4148) <= a;
    layer4_outputs(4149) <= not b or a;
    layer4_outputs(4150) <= '0';
    layer4_outputs(4151) <= b;
    layer4_outputs(4152) <= b;
    layer4_outputs(4153) <= a xor b;
    layer4_outputs(4154) <= not a or b;
    layer4_outputs(4155) <= not (a and b);
    layer4_outputs(4156) <= not b or a;
    layer4_outputs(4157) <= not (a and b);
    layer4_outputs(4158) <= a and not b;
    layer4_outputs(4159) <= not b;
    layer4_outputs(4160) <= not (a and b);
    layer4_outputs(4161) <= not (a or b);
    layer4_outputs(4162) <= not (a and b);
    layer4_outputs(4163) <= '0';
    layer4_outputs(4164) <= not (a and b);
    layer4_outputs(4165) <= not b or a;
    layer4_outputs(4166) <= a and b;
    layer4_outputs(4167) <= a;
    layer4_outputs(4168) <= not (a and b);
    layer4_outputs(4169) <= a and b;
    layer4_outputs(4170) <= not (a and b);
    layer4_outputs(4171) <= a;
    layer4_outputs(4172) <= not (a and b);
    layer4_outputs(4173) <= not (a and b);
    layer4_outputs(4174) <= not b;
    layer4_outputs(4175) <= not (a or b);
    layer4_outputs(4176) <= not b or a;
    layer4_outputs(4177) <= b;
    layer4_outputs(4178) <= not a;
    layer4_outputs(4179) <= not a;
    layer4_outputs(4180) <= '1';
    layer4_outputs(4181) <= b;
    layer4_outputs(4182) <= not a or b;
    layer4_outputs(4183) <= a or b;
    layer4_outputs(4184) <= b;
    layer4_outputs(4185) <= not (a or b);
    layer4_outputs(4186) <= not (a and b);
    layer4_outputs(4187) <= not (a or b);
    layer4_outputs(4188) <= not a;
    layer4_outputs(4189) <= not b or a;
    layer4_outputs(4190) <= b;
    layer4_outputs(4191) <= not b;
    layer4_outputs(4192) <= not a or b;
    layer4_outputs(4193) <= a and not b;
    layer4_outputs(4194) <= not (a xor b);
    layer4_outputs(4195) <= a or b;
    layer4_outputs(4196) <= b;
    layer4_outputs(4197) <= a and not b;
    layer4_outputs(4198) <= '1';
    layer4_outputs(4199) <= '0';
    layer4_outputs(4200) <= not b or a;
    layer4_outputs(4201) <= b;
    layer4_outputs(4202) <= a or b;
    layer4_outputs(4203) <= not a or b;
    layer4_outputs(4204) <= '1';
    layer4_outputs(4205) <= not (a and b);
    layer4_outputs(4206) <= b and not a;
    layer4_outputs(4207) <= not (a or b);
    layer4_outputs(4208) <= b and not a;
    layer4_outputs(4209) <= not b;
    layer4_outputs(4210) <= a and not b;
    layer4_outputs(4211) <= a or b;
    layer4_outputs(4212) <= not a;
    layer4_outputs(4213) <= a and b;
    layer4_outputs(4214) <= '1';
    layer4_outputs(4215) <= not b;
    layer4_outputs(4216) <= a and not b;
    layer4_outputs(4217) <= not (a or b);
    layer4_outputs(4218) <= not (a and b);
    layer4_outputs(4219) <= a;
    layer4_outputs(4220) <= not b or a;
    layer4_outputs(4221) <= b and not a;
    layer4_outputs(4222) <= a;
    layer4_outputs(4223) <= not a or b;
    layer4_outputs(4224) <= b and not a;
    layer4_outputs(4225) <= '1';
    layer4_outputs(4226) <= not (a and b);
    layer4_outputs(4227) <= not (a and b);
    layer4_outputs(4228) <= a;
    layer4_outputs(4229) <= not b or a;
    layer4_outputs(4230) <= not b or a;
    layer4_outputs(4231) <= a or b;
    layer4_outputs(4232) <= a;
    layer4_outputs(4233) <= a and not b;
    layer4_outputs(4234) <= b;
    layer4_outputs(4235) <= not a or b;
    layer4_outputs(4236) <= not (a or b);
    layer4_outputs(4237) <= a xor b;
    layer4_outputs(4238) <= '1';
    layer4_outputs(4239) <= a or b;
    layer4_outputs(4240) <= a and b;
    layer4_outputs(4241) <= a;
    layer4_outputs(4242) <= not b or a;
    layer4_outputs(4243) <= a;
    layer4_outputs(4244) <= not a;
    layer4_outputs(4245) <= not (a and b);
    layer4_outputs(4246) <= a and b;
    layer4_outputs(4247) <= b;
    layer4_outputs(4248) <= a and not b;
    layer4_outputs(4249) <= '0';
    layer4_outputs(4250) <= b;
    layer4_outputs(4251) <= not b or a;
    layer4_outputs(4252) <= '0';
    layer4_outputs(4253) <= '0';
    layer4_outputs(4254) <= not a or b;
    layer4_outputs(4255) <= a;
    layer4_outputs(4256) <= a or b;
    layer4_outputs(4257) <= b;
    layer4_outputs(4258) <= a and not b;
    layer4_outputs(4259) <= a and not b;
    layer4_outputs(4260) <= a xor b;
    layer4_outputs(4261) <= a and b;
    layer4_outputs(4262) <= a and not b;
    layer4_outputs(4263) <= not a or b;
    layer4_outputs(4264) <= b and not a;
    layer4_outputs(4265) <= b;
    layer4_outputs(4266) <= not a;
    layer4_outputs(4267) <= a or b;
    layer4_outputs(4268) <= a;
    layer4_outputs(4269) <= a xor b;
    layer4_outputs(4270) <= b;
    layer4_outputs(4271) <= not b or a;
    layer4_outputs(4272) <= a and b;
    layer4_outputs(4273) <= not a or b;
    layer4_outputs(4274) <= not (a xor b);
    layer4_outputs(4275) <= a and b;
    layer4_outputs(4276) <= '0';
    layer4_outputs(4277) <= '0';
    layer4_outputs(4278) <= a and b;
    layer4_outputs(4279) <= not (a or b);
    layer4_outputs(4280) <= a or b;
    layer4_outputs(4281) <= not b or a;
    layer4_outputs(4282) <= a xor b;
    layer4_outputs(4283) <= not a;
    layer4_outputs(4284) <= a and not b;
    layer4_outputs(4285) <= a and not b;
    layer4_outputs(4286) <= not a;
    layer4_outputs(4287) <= a or b;
    layer4_outputs(4288) <= not (a or b);
    layer4_outputs(4289) <= a;
    layer4_outputs(4290) <= a and b;
    layer4_outputs(4291) <= not (a and b);
    layer4_outputs(4292) <= a;
    layer4_outputs(4293) <= not a or b;
    layer4_outputs(4294) <= a and b;
    layer4_outputs(4295) <= not b;
    layer4_outputs(4296) <= not b;
    layer4_outputs(4297) <= a or b;
    layer4_outputs(4298) <= a and not b;
    layer4_outputs(4299) <= not b;
    layer4_outputs(4300) <= '0';
    layer4_outputs(4301) <= not (a xor b);
    layer4_outputs(4302) <= not a;
    layer4_outputs(4303) <= not (a and b);
    layer4_outputs(4304) <= not a;
    layer4_outputs(4305) <= not b;
    layer4_outputs(4306) <= not b;
    layer4_outputs(4307) <= a or b;
    layer4_outputs(4308) <= b and not a;
    layer4_outputs(4309) <= b and not a;
    layer4_outputs(4310) <= a or b;
    layer4_outputs(4311) <= a or b;
    layer4_outputs(4312) <= a xor b;
    layer4_outputs(4313) <= not (a or b);
    layer4_outputs(4314) <= '1';
    layer4_outputs(4315) <= a and b;
    layer4_outputs(4316) <= not (a or b);
    layer4_outputs(4317) <= not b or a;
    layer4_outputs(4318) <= not (a or b);
    layer4_outputs(4319) <= a or b;
    layer4_outputs(4320) <= a and not b;
    layer4_outputs(4321) <= not (a or b);
    layer4_outputs(4322) <= not (a and b);
    layer4_outputs(4323) <= a xor b;
    layer4_outputs(4324) <= not b;
    layer4_outputs(4325) <= b and not a;
    layer4_outputs(4326) <= a and b;
    layer4_outputs(4327) <= not b;
    layer4_outputs(4328) <= b and not a;
    layer4_outputs(4329) <= b;
    layer4_outputs(4330) <= a;
    layer4_outputs(4331) <= not (a or b);
    layer4_outputs(4332) <= not (a and b);
    layer4_outputs(4333) <= not b;
    layer4_outputs(4334) <= a and not b;
    layer4_outputs(4335) <= '0';
    layer4_outputs(4336) <= a and not b;
    layer4_outputs(4337) <= a and not b;
    layer4_outputs(4338) <= not a;
    layer4_outputs(4339) <= not (a xor b);
    layer4_outputs(4340) <= not (a or b);
    layer4_outputs(4341) <= b and not a;
    layer4_outputs(4342) <= b;
    layer4_outputs(4343) <= '1';
    layer4_outputs(4344) <= a or b;
    layer4_outputs(4345) <= a and b;
    layer4_outputs(4346) <= a or b;
    layer4_outputs(4347) <= a or b;
    layer4_outputs(4348) <= a or b;
    layer4_outputs(4349) <= b and not a;
    layer4_outputs(4350) <= '1';
    layer4_outputs(4351) <= a;
    layer4_outputs(4352) <= '0';
    layer4_outputs(4353) <= '0';
    layer4_outputs(4354) <= a;
    layer4_outputs(4355) <= a;
    layer4_outputs(4356) <= not (a or b);
    layer4_outputs(4357) <= a;
    layer4_outputs(4358) <= b;
    layer4_outputs(4359) <= a and b;
    layer4_outputs(4360) <= a and b;
    layer4_outputs(4361) <= not a or b;
    layer4_outputs(4362) <= a and b;
    layer4_outputs(4363) <= not (a and b);
    layer4_outputs(4364) <= a;
    layer4_outputs(4365) <= b and not a;
    layer4_outputs(4366) <= not a;
    layer4_outputs(4367) <= '0';
    layer4_outputs(4368) <= not (a or b);
    layer4_outputs(4369) <= a;
    layer4_outputs(4370) <= a and not b;
    layer4_outputs(4371) <= a or b;
    layer4_outputs(4372) <= not b;
    layer4_outputs(4373) <= not a or b;
    layer4_outputs(4374) <= not (a or b);
    layer4_outputs(4375) <= not b;
    layer4_outputs(4376) <= '0';
    layer4_outputs(4377) <= a xor b;
    layer4_outputs(4378) <= not a;
    layer4_outputs(4379) <= b;
    layer4_outputs(4380) <= b;
    layer4_outputs(4381) <= b and not a;
    layer4_outputs(4382) <= a or b;
    layer4_outputs(4383) <= a;
    layer4_outputs(4384) <= not a;
    layer4_outputs(4385) <= a and not b;
    layer4_outputs(4386) <= not b;
    layer4_outputs(4387) <= '0';
    layer4_outputs(4388) <= a and b;
    layer4_outputs(4389) <= a xor b;
    layer4_outputs(4390) <= not (a and b);
    layer4_outputs(4391) <= a or b;
    layer4_outputs(4392) <= not b;
    layer4_outputs(4393) <= '0';
    layer4_outputs(4394) <= not b or a;
    layer4_outputs(4395) <= a;
    layer4_outputs(4396) <= not b;
    layer4_outputs(4397) <= not (a and b);
    layer4_outputs(4398) <= b;
    layer4_outputs(4399) <= not b or a;
    layer4_outputs(4400) <= not (a or b);
    layer4_outputs(4401) <= not a;
    layer4_outputs(4402) <= not (a and b);
    layer4_outputs(4403) <= not b;
    layer4_outputs(4404) <= a;
    layer4_outputs(4405) <= a and b;
    layer4_outputs(4406) <= a and not b;
    layer4_outputs(4407) <= not b or a;
    layer4_outputs(4408) <= '1';
    layer4_outputs(4409) <= a or b;
    layer4_outputs(4410) <= a;
    layer4_outputs(4411) <= '1';
    layer4_outputs(4412) <= '1';
    layer4_outputs(4413) <= '0';
    layer4_outputs(4414) <= a;
    layer4_outputs(4415) <= not b;
    layer4_outputs(4416) <= b and not a;
    layer4_outputs(4417) <= not b;
    layer4_outputs(4418) <= not a or b;
    layer4_outputs(4419) <= b and not a;
    layer4_outputs(4420) <= '1';
    layer4_outputs(4421) <= not (a or b);
    layer4_outputs(4422) <= a or b;
    layer4_outputs(4423) <= not b or a;
    layer4_outputs(4424) <= not a or b;
    layer4_outputs(4425) <= not (a or b);
    layer4_outputs(4426) <= not a or b;
    layer4_outputs(4427) <= not b or a;
    layer4_outputs(4428) <= a;
    layer4_outputs(4429) <= not b;
    layer4_outputs(4430) <= not (a and b);
    layer4_outputs(4431) <= b;
    layer4_outputs(4432) <= '1';
    layer4_outputs(4433) <= a;
    layer4_outputs(4434) <= b and not a;
    layer4_outputs(4435) <= a and not b;
    layer4_outputs(4436) <= b and not a;
    layer4_outputs(4437) <= b;
    layer4_outputs(4438) <= not b or a;
    layer4_outputs(4439) <= not a;
    layer4_outputs(4440) <= b;
    layer4_outputs(4441) <= a or b;
    layer4_outputs(4442) <= a or b;
    layer4_outputs(4443) <= '0';
    layer4_outputs(4444) <= a;
    layer4_outputs(4445) <= not b or a;
    layer4_outputs(4446) <= not a or b;
    layer4_outputs(4447) <= a and b;
    layer4_outputs(4448) <= not b;
    layer4_outputs(4449) <= '0';
    layer4_outputs(4450) <= not b or a;
    layer4_outputs(4451) <= not (a and b);
    layer4_outputs(4452) <= b and not a;
    layer4_outputs(4453) <= '0';
    layer4_outputs(4454) <= not b;
    layer4_outputs(4455) <= a or b;
    layer4_outputs(4456) <= a and not b;
    layer4_outputs(4457) <= a;
    layer4_outputs(4458) <= not (a and b);
    layer4_outputs(4459) <= not b or a;
    layer4_outputs(4460) <= a;
    layer4_outputs(4461) <= not b or a;
    layer4_outputs(4462) <= a;
    layer4_outputs(4463) <= a;
    layer4_outputs(4464) <= not a or b;
    layer4_outputs(4465) <= a or b;
    layer4_outputs(4466) <= a;
    layer4_outputs(4467) <= b;
    layer4_outputs(4468) <= not b;
    layer4_outputs(4469) <= not (a or b);
    layer4_outputs(4470) <= not (a and b);
    layer4_outputs(4471) <= not (a and b);
    layer4_outputs(4472) <= not b;
    layer4_outputs(4473) <= not a or b;
    layer4_outputs(4474) <= not (a and b);
    layer4_outputs(4475) <= a;
    layer4_outputs(4476) <= a;
    layer4_outputs(4477) <= a or b;
    layer4_outputs(4478) <= a and not b;
    layer4_outputs(4479) <= not a or b;
    layer4_outputs(4480) <= a and b;
    layer4_outputs(4481) <= b;
    layer4_outputs(4482) <= not (a and b);
    layer4_outputs(4483) <= a;
    layer4_outputs(4484) <= a;
    layer4_outputs(4485) <= '0';
    layer4_outputs(4486) <= not a;
    layer4_outputs(4487) <= not a or b;
    layer4_outputs(4488) <= '1';
    layer4_outputs(4489) <= not b or a;
    layer4_outputs(4490) <= not b or a;
    layer4_outputs(4491) <= a;
    layer4_outputs(4492) <= a or b;
    layer4_outputs(4493) <= not (a or b);
    layer4_outputs(4494) <= not a;
    layer4_outputs(4495) <= b;
    layer4_outputs(4496) <= not a or b;
    layer4_outputs(4497) <= not (a or b);
    layer4_outputs(4498) <= not (a or b);
    layer4_outputs(4499) <= b and not a;
    layer4_outputs(4500) <= a and b;
    layer4_outputs(4501) <= not a;
    layer4_outputs(4502) <= not b or a;
    layer4_outputs(4503) <= not b;
    layer4_outputs(4504) <= not (a and b);
    layer4_outputs(4505) <= not b;
    layer4_outputs(4506) <= not b or a;
    layer4_outputs(4507) <= a;
    layer4_outputs(4508) <= not a or b;
    layer4_outputs(4509) <= a or b;
    layer4_outputs(4510) <= a or b;
    layer4_outputs(4511) <= a;
    layer4_outputs(4512) <= a and b;
    layer4_outputs(4513) <= a;
    layer4_outputs(4514) <= not a or b;
    layer4_outputs(4515) <= b;
    layer4_outputs(4516) <= b;
    layer4_outputs(4517) <= a and not b;
    layer4_outputs(4518) <= a xor b;
    layer4_outputs(4519) <= not b or a;
    layer4_outputs(4520) <= not (a and b);
    layer4_outputs(4521) <= a xor b;
    layer4_outputs(4522) <= not (a or b);
    layer4_outputs(4523) <= b;
    layer4_outputs(4524) <= b and not a;
    layer4_outputs(4525) <= a and b;
    layer4_outputs(4526) <= not b or a;
    layer4_outputs(4527) <= '0';
    layer4_outputs(4528) <= a and b;
    layer4_outputs(4529) <= a;
    layer4_outputs(4530) <= b and not a;
    layer4_outputs(4531) <= '0';
    layer4_outputs(4532) <= a or b;
    layer4_outputs(4533) <= b and not a;
    layer4_outputs(4534) <= not b;
    layer4_outputs(4535) <= '0';
    layer4_outputs(4536) <= not b;
    layer4_outputs(4537) <= b and not a;
    layer4_outputs(4538) <= not (a or b);
    layer4_outputs(4539) <= b and not a;
    layer4_outputs(4540) <= b and not a;
    layer4_outputs(4541) <= not a or b;
    layer4_outputs(4542) <= b;
    layer4_outputs(4543) <= not a;
    layer4_outputs(4544) <= not b or a;
    layer4_outputs(4545) <= not a;
    layer4_outputs(4546) <= a;
    layer4_outputs(4547) <= a and b;
    layer4_outputs(4548) <= a;
    layer4_outputs(4549) <= not b;
    layer4_outputs(4550) <= '0';
    layer4_outputs(4551) <= b;
    layer4_outputs(4552) <= b and not a;
    layer4_outputs(4553) <= not (a and b);
    layer4_outputs(4554) <= '1';
    layer4_outputs(4555) <= not a or b;
    layer4_outputs(4556) <= not b or a;
    layer4_outputs(4557) <= '0';
    layer4_outputs(4558) <= not (a and b);
    layer4_outputs(4559) <= b;
    layer4_outputs(4560) <= a and b;
    layer4_outputs(4561) <= '1';
    layer4_outputs(4562) <= b;
    layer4_outputs(4563) <= not a or b;
    layer4_outputs(4564) <= '0';
    layer4_outputs(4565) <= not (a xor b);
    layer4_outputs(4566) <= not b or a;
    layer4_outputs(4567) <= a or b;
    layer4_outputs(4568) <= not b or a;
    layer4_outputs(4569) <= not b or a;
    layer4_outputs(4570) <= not a or b;
    layer4_outputs(4571) <= a or b;
    layer4_outputs(4572) <= a;
    layer4_outputs(4573) <= not a;
    layer4_outputs(4574) <= not a;
    layer4_outputs(4575) <= '0';
    layer4_outputs(4576) <= a or b;
    layer4_outputs(4577) <= not (a and b);
    layer4_outputs(4578) <= b and not a;
    layer4_outputs(4579) <= a and not b;
    layer4_outputs(4580) <= b and not a;
    layer4_outputs(4581) <= a;
    layer4_outputs(4582) <= a xor b;
    layer4_outputs(4583) <= '1';
    layer4_outputs(4584) <= not a or b;
    layer4_outputs(4585) <= not b or a;
    layer4_outputs(4586) <= not (a and b);
    layer4_outputs(4587) <= '0';
    layer4_outputs(4588) <= b and not a;
    layer4_outputs(4589) <= not (a or b);
    layer4_outputs(4590) <= a or b;
    layer4_outputs(4591) <= b and not a;
    layer4_outputs(4592) <= not (a and b);
    layer4_outputs(4593) <= not (a and b);
    layer4_outputs(4594) <= b and not a;
    layer4_outputs(4595) <= '0';
    layer4_outputs(4596) <= not a or b;
    layer4_outputs(4597) <= not a;
    layer4_outputs(4598) <= not b;
    layer4_outputs(4599) <= b;
    layer4_outputs(4600) <= b;
    layer4_outputs(4601) <= a and b;
    layer4_outputs(4602) <= not (a and b);
    layer4_outputs(4603) <= a;
    layer4_outputs(4604) <= not b;
    layer4_outputs(4605) <= not (a and b);
    layer4_outputs(4606) <= not b;
    layer4_outputs(4607) <= not b;
    layer4_outputs(4608) <= '1';
    layer4_outputs(4609) <= not (a or b);
    layer4_outputs(4610) <= a and not b;
    layer4_outputs(4611) <= not b or a;
    layer4_outputs(4612) <= a and b;
    layer4_outputs(4613) <= not (a or b);
    layer4_outputs(4614) <= a or b;
    layer4_outputs(4615) <= not b;
    layer4_outputs(4616) <= not (a or b);
    layer4_outputs(4617) <= not (a and b);
    layer4_outputs(4618) <= a or b;
    layer4_outputs(4619) <= a;
    layer4_outputs(4620) <= a xor b;
    layer4_outputs(4621) <= a or b;
    layer4_outputs(4622) <= '0';
    layer4_outputs(4623) <= not (a and b);
    layer4_outputs(4624) <= not b;
    layer4_outputs(4625) <= not b;
    layer4_outputs(4626) <= '0';
    layer4_outputs(4627) <= not b;
    layer4_outputs(4628) <= not b;
    layer4_outputs(4629) <= not (a and b);
    layer4_outputs(4630) <= not b or a;
    layer4_outputs(4631) <= '0';
    layer4_outputs(4632) <= '0';
    layer4_outputs(4633) <= '1';
    layer4_outputs(4634) <= a;
    layer4_outputs(4635) <= a or b;
    layer4_outputs(4636) <= not (a or b);
    layer4_outputs(4637) <= not (a or b);
    layer4_outputs(4638) <= a or b;
    layer4_outputs(4639) <= not b;
    layer4_outputs(4640) <= not b or a;
    layer4_outputs(4641) <= '1';
    layer4_outputs(4642) <= a;
    layer4_outputs(4643) <= '1';
    layer4_outputs(4644) <= b and not a;
    layer4_outputs(4645) <= b;
    layer4_outputs(4646) <= not a;
    layer4_outputs(4647) <= not (a or b);
    layer4_outputs(4648) <= b;
    layer4_outputs(4649) <= b;
    layer4_outputs(4650) <= not (a or b);
    layer4_outputs(4651) <= not b;
    layer4_outputs(4652) <= not a;
    layer4_outputs(4653) <= a or b;
    layer4_outputs(4654) <= '1';
    layer4_outputs(4655) <= not b or a;
    layer4_outputs(4656) <= a and b;
    layer4_outputs(4657) <= a and not b;
    layer4_outputs(4658) <= a and not b;
    layer4_outputs(4659) <= a;
    layer4_outputs(4660) <= not b or a;
    layer4_outputs(4661) <= a and not b;
    layer4_outputs(4662) <= b and not a;
    layer4_outputs(4663) <= b and not a;
    layer4_outputs(4664) <= not a;
    layer4_outputs(4665) <= '1';
    layer4_outputs(4666) <= '0';
    layer4_outputs(4667) <= not (a xor b);
    layer4_outputs(4668) <= a and b;
    layer4_outputs(4669) <= not a or b;
    layer4_outputs(4670) <= not a or b;
    layer4_outputs(4671) <= '1';
    layer4_outputs(4672) <= not a or b;
    layer4_outputs(4673) <= not b or a;
    layer4_outputs(4674) <= not b;
    layer4_outputs(4675) <= b and not a;
    layer4_outputs(4676) <= not b or a;
    layer4_outputs(4677) <= '1';
    layer4_outputs(4678) <= a;
    layer4_outputs(4679) <= a;
    layer4_outputs(4680) <= not (a or b);
    layer4_outputs(4681) <= '0';
    layer4_outputs(4682) <= not (a and b);
    layer4_outputs(4683) <= a;
    layer4_outputs(4684) <= a and not b;
    layer4_outputs(4685) <= b and not a;
    layer4_outputs(4686) <= not a;
    layer4_outputs(4687) <= not b or a;
    layer4_outputs(4688) <= not a or b;
    layer4_outputs(4689) <= not b;
    layer4_outputs(4690) <= a xor b;
    layer4_outputs(4691) <= not a;
    layer4_outputs(4692) <= a xor b;
    layer4_outputs(4693) <= not (a and b);
    layer4_outputs(4694) <= b and not a;
    layer4_outputs(4695) <= a and b;
    layer4_outputs(4696) <= not a or b;
    layer4_outputs(4697) <= not (a and b);
    layer4_outputs(4698) <= not a or b;
    layer4_outputs(4699) <= a;
    layer4_outputs(4700) <= a xor b;
    layer4_outputs(4701) <= a or b;
    layer4_outputs(4702) <= not (a or b);
    layer4_outputs(4703) <= a;
    layer4_outputs(4704) <= a;
    layer4_outputs(4705) <= not (a xor b);
    layer4_outputs(4706) <= a xor b;
    layer4_outputs(4707) <= a;
    layer4_outputs(4708) <= b;
    layer4_outputs(4709) <= not (a or b);
    layer4_outputs(4710) <= not (a xor b);
    layer4_outputs(4711) <= '0';
    layer4_outputs(4712) <= not a;
    layer4_outputs(4713) <= a and b;
    layer4_outputs(4714) <= not b;
    layer4_outputs(4715) <= a xor b;
    layer4_outputs(4716) <= a or b;
    layer4_outputs(4717) <= '1';
    layer4_outputs(4718) <= not a or b;
    layer4_outputs(4719) <= a;
    layer4_outputs(4720) <= not a;
    layer4_outputs(4721) <= not a;
    layer4_outputs(4722) <= '1';
    layer4_outputs(4723) <= b;
    layer4_outputs(4724) <= not a;
    layer4_outputs(4725) <= not a or b;
    layer4_outputs(4726) <= '0';
    layer4_outputs(4727) <= '0';
    layer4_outputs(4728) <= '0';
    layer4_outputs(4729) <= a and not b;
    layer4_outputs(4730) <= not a;
    layer4_outputs(4731) <= '0';
    layer4_outputs(4732) <= not a;
    layer4_outputs(4733) <= not (a or b);
    layer4_outputs(4734) <= not a;
    layer4_outputs(4735) <= b;
    layer4_outputs(4736) <= not (a xor b);
    layer4_outputs(4737) <= a xor b;
    layer4_outputs(4738) <= '0';
    layer4_outputs(4739) <= not b or a;
    layer4_outputs(4740) <= a or b;
    layer4_outputs(4741) <= a and not b;
    layer4_outputs(4742) <= '0';
    layer4_outputs(4743) <= not a;
    layer4_outputs(4744) <= a or b;
    layer4_outputs(4745) <= not (a or b);
    layer4_outputs(4746) <= not (a or b);
    layer4_outputs(4747) <= not b or a;
    layer4_outputs(4748) <= not b;
    layer4_outputs(4749) <= not a;
    layer4_outputs(4750) <= '0';
    layer4_outputs(4751) <= a;
    layer4_outputs(4752) <= a or b;
    layer4_outputs(4753) <= not b;
    layer4_outputs(4754) <= not b;
    layer4_outputs(4755) <= not a;
    layer4_outputs(4756) <= a xor b;
    layer4_outputs(4757) <= not (a or b);
    layer4_outputs(4758) <= a and b;
    layer4_outputs(4759) <= not b or a;
    layer4_outputs(4760) <= not a or b;
    layer4_outputs(4761) <= not (a and b);
    layer4_outputs(4762) <= not b;
    layer4_outputs(4763) <= '1';
    layer4_outputs(4764) <= not a or b;
    layer4_outputs(4765) <= a or b;
    layer4_outputs(4766) <= a xor b;
    layer4_outputs(4767) <= not b;
    layer4_outputs(4768) <= not (a or b);
    layer4_outputs(4769) <= not b;
    layer4_outputs(4770) <= a or b;
    layer4_outputs(4771) <= not a or b;
    layer4_outputs(4772) <= not a;
    layer4_outputs(4773) <= a xor b;
    layer4_outputs(4774) <= not (a or b);
    layer4_outputs(4775) <= '0';
    layer4_outputs(4776) <= a xor b;
    layer4_outputs(4777) <= b;
    layer4_outputs(4778) <= not b or a;
    layer4_outputs(4779) <= a and b;
    layer4_outputs(4780) <= a and not b;
    layer4_outputs(4781) <= not b or a;
    layer4_outputs(4782) <= not (a xor b);
    layer4_outputs(4783) <= not a;
    layer4_outputs(4784) <= b;
    layer4_outputs(4785) <= not a;
    layer4_outputs(4786) <= not (a or b);
    layer4_outputs(4787) <= not (a or b);
    layer4_outputs(4788) <= b;
    layer4_outputs(4789) <= a or b;
    layer4_outputs(4790) <= '1';
    layer4_outputs(4791) <= not a or b;
    layer4_outputs(4792) <= not b;
    layer4_outputs(4793) <= a;
    layer4_outputs(4794) <= a;
    layer4_outputs(4795) <= not b or a;
    layer4_outputs(4796) <= '1';
    layer4_outputs(4797) <= a and b;
    layer4_outputs(4798) <= a and not b;
    layer4_outputs(4799) <= not a;
    layer4_outputs(4800) <= a or b;
    layer4_outputs(4801) <= a or b;
    layer4_outputs(4802) <= not a;
    layer4_outputs(4803) <= not (a or b);
    layer4_outputs(4804) <= not a;
    layer4_outputs(4805) <= not b or a;
    layer4_outputs(4806) <= a and b;
    layer4_outputs(4807) <= not b or a;
    layer4_outputs(4808) <= not b or a;
    layer4_outputs(4809) <= not b or a;
    layer4_outputs(4810) <= not b;
    layer4_outputs(4811) <= not a;
    layer4_outputs(4812) <= not b;
    layer4_outputs(4813) <= a;
    layer4_outputs(4814) <= a or b;
    layer4_outputs(4815) <= not b or a;
    layer4_outputs(4816) <= not b;
    layer4_outputs(4817) <= a and not b;
    layer4_outputs(4818) <= not (a or b);
    layer4_outputs(4819) <= a;
    layer4_outputs(4820) <= not a;
    layer4_outputs(4821) <= a and b;
    layer4_outputs(4822) <= b and not a;
    layer4_outputs(4823) <= not b;
    layer4_outputs(4824) <= a;
    layer4_outputs(4825) <= a;
    layer4_outputs(4826) <= not (a or b);
    layer4_outputs(4827) <= not (a and b);
    layer4_outputs(4828) <= b and not a;
    layer4_outputs(4829) <= not b;
    layer4_outputs(4830) <= not b;
    layer4_outputs(4831) <= a and b;
    layer4_outputs(4832) <= not (a or b);
    layer4_outputs(4833) <= not a or b;
    layer4_outputs(4834) <= b and not a;
    layer4_outputs(4835) <= not b;
    layer4_outputs(4836) <= not a or b;
    layer4_outputs(4837) <= not b;
    layer4_outputs(4838) <= a;
    layer4_outputs(4839) <= not a or b;
    layer4_outputs(4840) <= not a;
    layer4_outputs(4841) <= not a;
    layer4_outputs(4842) <= a or b;
    layer4_outputs(4843) <= not b;
    layer4_outputs(4844) <= '0';
    layer4_outputs(4845) <= b and not a;
    layer4_outputs(4846) <= a and b;
    layer4_outputs(4847) <= a and not b;
    layer4_outputs(4848) <= a and not b;
    layer4_outputs(4849) <= a and b;
    layer4_outputs(4850) <= '0';
    layer4_outputs(4851) <= b and not a;
    layer4_outputs(4852) <= not (a or b);
    layer4_outputs(4853) <= b and not a;
    layer4_outputs(4854) <= a or b;
    layer4_outputs(4855) <= not a;
    layer4_outputs(4856) <= not b;
    layer4_outputs(4857) <= not b or a;
    layer4_outputs(4858) <= not (a xor b);
    layer4_outputs(4859) <= not a or b;
    layer4_outputs(4860) <= not b;
    layer4_outputs(4861) <= not (a and b);
    layer4_outputs(4862) <= not a or b;
    layer4_outputs(4863) <= b;
    layer4_outputs(4864) <= not a;
    layer4_outputs(4865) <= a or b;
    layer4_outputs(4866) <= not (a xor b);
    layer4_outputs(4867) <= not b or a;
    layer4_outputs(4868) <= not b;
    layer4_outputs(4869) <= '1';
    layer4_outputs(4870) <= not a or b;
    layer4_outputs(4871) <= not b;
    layer4_outputs(4872) <= not a;
    layer4_outputs(4873) <= a;
    layer4_outputs(4874) <= a and b;
    layer4_outputs(4875) <= '0';
    layer4_outputs(4876) <= not b;
    layer4_outputs(4877) <= not b or a;
    layer4_outputs(4878) <= a or b;
    layer4_outputs(4879) <= not b;
    layer4_outputs(4880) <= not b or a;
    layer4_outputs(4881) <= not a;
    layer4_outputs(4882) <= '1';
    layer4_outputs(4883) <= b and not a;
    layer4_outputs(4884) <= not (a and b);
    layer4_outputs(4885) <= b;
    layer4_outputs(4886) <= '0';
    layer4_outputs(4887) <= not (a or b);
    layer4_outputs(4888) <= not (a or b);
    layer4_outputs(4889) <= '0';
    layer4_outputs(4890) <= a;
    layer4_outputs(4891) <= b;
    layer4_outputs(4892) <= not b;
    layer4_outputs(4893) <= b and not a;
    layer4_outputs(4894) <= a xor b;
    layer4_outputs(4895) <= not b or a;
    layer4_outputs(4896) <= not b or a;
    layer4_outputs(4897) <= not b or a;
    layer4_outputs(4898) <= not b;
    layer4_outputs(4899) <= not b;
    layer4_outputs(4900) <= '0';
    layer4_outputs(4901) <= a or b;
    layer4_outputs(4902) <= a;
    layer4_outputs(4903) <= b and not a;
    layer4_outputs(4904) <= not a;
    layer4_outputs(4905) <= not a;
    layer4_outputs(4906) <= a and b;
    layer4_outputs(4907) <= a and b;
    layer4_outputs(4908) <= b;
    layer4_outputs(4909) <= not b;
    layer4_outputs(4910) <= '1';
    layer4_outputs(4911) <= not a;
    layer4_outputs(4912) <= not b or a;
    layer4_outputs(4913) <= '0';
    layer4_outputs(4914) <= b;
    layer4_outputs(4915) <= not b;
    layer4_outputs(4916) <= b;
    layer4_outputs(4917) <= not a or b;
    layer4_outputs(4918) <= a and not b;
    layer4_outputs(4919) <= not b or a;
    layer4_outputs(4920) <= not (a or b);
    layer4_outputs(4921) <= a and b;
    layer4_outputs(4922) <= not b;
    layer4_outputs(4923) <= a and not b;
    layer4_outputs(4924) <= a and not b;
    layer4_outputs(4925) <= a;
    layer4_outputs(4926) <= not (a and b);
    layer4_outputs(4927) <= a xor b;
    layer4_outputs(4928) <= not (a or b);
    layer4_outputs(4929) <= not a or b;
    layer4_outputs(4930) <= a and not b;
    layer4_outputs(4931) <= not (a xor b);
    layer4_outputs(4932) <= '0';
    layer4_outputs(4933) <= not b or a;
    layer4_outputs(4934) <= a;
    layer4_outputs(4935) <= not a or b;
    layer4_outputs(4936) <= a and not b;
    layer4_outputs(4937) <= not (a or b);
    layer4_outputs(4938) <= not a;
    layer4_outputs(4939) <= not b;
    layer4_outputs(4940) <= a;
    layer4_outputs(4941) <= not (a or b);
    layer4_outputs(4942) <= a and b;
    layer4_outputs(4943) <= a;
    layer4_outputs(4944) <= a and b;
    layer4_outputs(4945) <= '0';
    layer4_outputs(4946) <= not b;
    layer4_outputs(4947) <= not (a and b);
    layer4_outputs(4948) <= b;
    layer4_outputs(4949) <= not a or b;
    layer4_outputs(4950) <= '0';
    layer4_outputs(4951) <= not a or b;
    layer4_outputs(4952) <= a or b;
    layer4_outputs(4953) <= a xor b;
    layer4_outputs(4954) <= not (a or b);
    layer4_outputs(4955) <= a or b;
    layer4_outputs(4956) <= not (a and b);
    layer4_outputs(4957) <= a;
    layer4_outputs(4958) <= a;
    layer4_outputs(4959) <= not b;
    layer4_outputs(4960) <= not (a and b);
    layer4_outputs(4961) <= '0';
    layer4_outputs(4962) <= not b or a;
    layer4_outputs(4963) <= a or b;
    layer4_outputs(4964) <= a;
    layer4_outputs(4965) <= not b;
    layer4_outputs(4966) <= not b or a;
    layer4_outputs(4967) <= not (a or b);
    layer4_outputs(4968) <= not a;
    layer4_outputs(4969) <= '1';
    layer4_outputs(4970) <= b;
    layer4_outputs(4971) <= a and b;
    layer4_outputs(4972) <= not (a or b);
    layer4_outputs(4973) <= a;
    layer4_outputs(4974) <= '0';
    layer4_outputs(4975) <= not b or a;
    layer4_outputs(4976) <= not a;
    layer4_outputs(4977) <= not b or a;
    layer4_outputs(4978) <= not a;
    layer4_outputs(4979) <= not (a or b);
    layer4_outputs(4980) <= a;
    layer4_outputs(4981) <= '0';
    layer4_outputs(4982) <= not a;
    layer4_outputs(4983) <= a and b;
    layer4_outputs(4984) <= a;
    layer4_outputs(4985) <= b and not a;
    layer4_outputs(4986) <= not b;
    layer4_outputs(4987) <= b and not a;
    layer4_outputs(4988) <= a and not b;
    layer4_outputs(4989) <= a and not b;
    layer4_outputs(4990) <= b;
    layer4_outputs(4991) <= a;
    layer4_outputs(4992) <= b;
    layer4_outputs(4993) <= not (a xor b);
    layer4_outputs(4994) <= not b or a;
    layer4_outputs(4995) <= a or b;
    layer4_outputs(4996) <= not a or b;
    layer4_outputs(4997) <= '1';
    layer4_outputs(4998) <= not b;
    layer4_outputs(4999) <= not b;
    layer4_outputs(5000) <= not a or b;
    layer4_outputs(5001) <= '0';
    layer4_outputs(5002) <= '0';
    layer4_outputs(5003) <= not a or b;
    layer4_outputs(5004) <= not a or b;
    layer4_outputs(5005) <= '1';
    layer4_outputs(5006) <= a and b;
    layer4_outputs(5007) <= b;
    layer4_outputs(5008) <= a and b;
    layer4_outputs(5009) <= '1';
    layer4_outputs(5010) <= not (a or b);
    layer4_outputs(5011) <= not (a and b);
    layer4_outputs(5012) <= b;
    layer4_outputs(5013) <= '0';
    layer4_outputs(5014) <= not b or a;
    layer4_outputs(5015) <= a and b;
    layer4_outputs(5016) <= a and b;
    layer4_outputs(5017) <= b and not a;
    layer4_outputs(5018) <= a;
    layer4_outputs(5019) <= not a or b;
    layer4_outputs(5020) <= a or b;
    layer4_outputs(5021) <= a;
    layer4_outputs(5022) <= not (a or b);
    layer4_outputs(5023) <= b;
    layer4_outputs(5024) <= a and b;
    layer4_outputs(5025) <= not b;
    layer4_outputs(5026) <= not b;
    layer4_outputs(5027) <= a;
    layer4_outputs(5028) <= not b;
    layer4_outputs(5029) <= not b;
    layer4_outputs(5030) <= a and b;
    layer4_outputs(5031) <= not b or a;
    layer4_outputs(5032) <= a and b;
    layer4_outputs(5033) <= not (a and b);
    layer4_outputs(5034) <= not a or b;
    layer4_outputs(5035) <= b;
    layer4_outputs(5036) <= a and not b;
    layer4_outputs(5037) <= not b;
    layer4_outputs(5038) <= not a;
    layer4_outputs(5039) <= a or b;
    layer4_outputs(5040) <= '1';
    layer4_outputs(5041) <= b and not a;
    layer4_outputs(5042) <= a;
    layer4_outputs(5043) <= '1';
    layer4_outputs(5044) <= not (a or b);
    layer4_outputs(5045) <= a and b;
    layer4_outputs(5046) <= b;
    layer4_outputs(5047) <= not (a and b);
    layer4_outputs(5048) <= b and not a;
    layer4_outputs(5049) <= a;
    layer4_outputs(5050) <= a and not b;
    layer4_outputs(5051) <= not a;
    layer4_outputs(5052) <= not (a or b);
    layer4_outputs(5053) <= a or b;
    layer4_outputs(5054) <= a or b;
    layer4_outputs(5055) <= a;
    layer4_outputs(5056) <= '1';
    layer4_outputs(5057) <= a and not b;
    layer4_outputs(5058) <= not b;
    layer4_outputs(5059) <= '1';
    layer4_outputs(5060) <= not a or b;
    layer4_outputs(5061) <= not (a and b);
    layer4_outputs(5062) <= not b;
    layer4_outputs(5063) <= a and not b;
    layer4_outputs(5064) <= not a;
    layer4_outputs(5065) <= not a;
    layer4_outputs(5066) <= b and not a;
    layer4_outputs(5067) <= not a;
    layer4_outputs(5068) <= not (a and b);
    layer4_outputs(5069) <= '1';
    layer4_outputs(5070) <= not (a or b);
    layer4_outputs(5071) <= not b or a;
    layer4_outputs(5072) <= b and not a;
    layer4_outputs(5073) <= a;
    layer4_outputs(5074) <= b;
    layer4_outputs(5075) <= not a;
    layer4_outputs(5076) <= a or b;
    layer4_outputs(5077) <= a;
    layer4_outputs(5078) <= a and not b;
    layer4_outputs(5079) <= a and b;
    layer4_outputs(5080) <= not (a or b);
    layer4_outputs(5081) <= b;
    layer4_outputs(5082) <= not a;
    layer4_outputs(5083) <= not b or a;
    layer4_outputs(5084) <= '0';
    layer4_outputs(5085) <= not a or b;
    layer4_outputs(5086) <= '0';
    layer4_outputs(5087) <= b;
    layer4_outputs(5088) <= not (a and b);
    layer4_outputs(5089) <= not (a and b);
    layer4_outputs(5090) <= '0';
    layer4_outputs(5091) <= not a;
    layer4_outputs(5092) <= not b;
    layer4_outputs(5093) <= '1';
    layer4_outputs(5094) <= a xor b;
    layer4_outputs(5095) <= not a or b;
    layer4_outputs(5096) <= not (a and b);
    layer4_outputs(5097) <= '1';
    layer4_outputs(5098) <= b and not a;
    layer4_outputs(5099) <= b and not a;
    layer4_outputs(5100) <= not b;
    layer4_outputs(5101) <= not (a and b);
    layer4_outputs(5102) <= a or b;
    layer4_outputs(5103) <= not b;
    layer4_outputs(5104) <= '1';
    layer4_outputs(5105) <= a or b;
    layer4_outputs(5106) <= b and not a;
    layer4_outputs(5107) <= not (a and b);
    layer4_outputs(5108) <= '0';
    layer4_outputs(5109) <= '0';
    layer4_outputs(5110) <= not b;
    layer4_outputs(5111) <= not a;
    layer4_outputs(5112) <= not b or a;
    layer4_outputs(5113) <= '1';
    layer4_outputs(5114) <= a;
    layer4_outputs(5115) <= not a or b;
    layer4_outputs(5116) <= not b or a;
    layer4_outputs(5117) <= a;
    layer4_outputs(5118) <= not (a xor b);
    layer4_outputs(5119) <= '0';
    layer5_outputs(0) <= not (a or b);
    layer5_outputs(1) <= not (a and b);
    layer5_outputs(2) <= a;
    layer5_outputs(3) <= not (a or b);
    layer5_outputs(4) <= not a or b;
    layer5_outputs(5) <= not a;
    layer5_outputs(6) <= b;
    layer5_outputs(7) <= not a;
    layer5_outputs(8) <= not b;
    layer5_outputs(9) <= not (a xor b);
    layer5_outputs(10) <= not a;
    layer5_outputs(11) <= not (a xor b);
    layer5_outputs(12) <= not a;
    layer5_outputs(13) <= not (a and b);
    layer5_outputs(14) <= '1';
    layer5_outputs(15) <= a;
    layer5_outputs(16) <= b;
    layer5_outputs(17) <= b and not a;
    layer5_outputs(18) <= not b or a;
    layer5_outputs(19) <= a;
    layer5_outputs(20) <= not (a or b);
    layer5_outputs(21) <= not a;
    layer5_outputs(22) <= not (a xor b);
    layer5_outputs(23) <= '1';
    layer5_outputs(24) <= b;
    layer5_outputs(25) <= not (a and b);
    layer5_outputs(26) <= not (a and b);
    layer5_outputs(27) <= a or b;
    layer5_outputs(28) <= not (a and b);
    layer5_outputs(29) <= not b;
    layer5_outputs(30) <= not a;
    layer5_outputs(31) <= not a;
    layer5_outputs(32) <= a xor b;
    layer5_outputs(33) <= a;
    layer5_outputs(34) <= b and not a;
    layer5_outputs(35) <= not (a xor b);
    layer5_outputs(36) <= not a;
    layer5_outputs(37) <= not a;
    layer5_outputs(38) <= not b;
    layer5_outputs(39) <= not b;
    layer5_outputs(40) <= '0';
    layer5_outputs(41) <= b and not a;
    layer5_outputs(42) <= a and b;
    layer5_outputs(43) <= not (a xor b);
    layer5_outputs(44) <= b;
    layer5_outputs(45) <= not a or b;
    layer5_outputs(46) <= '0';
    layer5_outputs(47) <= a and b;
    layer5_outputs(48) <= '1';
    layer5_outputs(49) <= a and not b;
    layer5_outputs(50) <= not b or a;
    layer5_outputs(51) <= not (a and b);
    layer5_outputs(52) <= not (a and b);
    layer5_outputs(53) <= a and b;
    layer5_outputs(54) <= a and not b;
    layer5_outputs(55) <= b;
    layer5_outputs(56) <= b;
    layer5_outputs(57) <= a and not b;
    layer5_outputs(58) <= a and not b;
    layer5_outputs(59) <= not (a and b);
    layer5_outputs(60) <= not (a and b);
    layer5_outputs(61) <= a;
    layer5_outputs(62) <= not a or b;
    layer5_outputs(63) <= a or b;
    layer5_outputs(64) <= '1';
    layer5_outputs(65) <= not a or b;
    layer5_outputs(66) <= not a or b;
    layer5_outputs(67) <= a and b;
    layer5_outputs(68) <= not a;
    layer5_outputs(69) <= not a;
    layer5_outputs(70) <= b;
    layer5_outputs(71) <= '0';
    layer5_outputs(72) <= a and not b;
    layer5_outputs(73) <= not (a and b);
    layer5_outputs(74) <= a and not b;
    layer5_outputs(75) <= a and b;
    layer5_outputs(76) <= not b;
    layer5_outputs(77) <= not a;
    layer5_outputs(78) <= a and b;
    layer5_outputs(79) <= '0';
    layer5_outputs(80) <= a xor b;
    layer5_outputs(81) <= b;
    layer5_outputs(82) <= not b or a;
    layer5_outputs(83) <= b;
    layer5_outputs(84) <= '0';
    layer5_outputs(85) <= a;
    layer5_outputs(86) <= a or b;
    layer5_outputs(87) <= not b or a;
    layer5_outputs(88) <= a and not b;
    layer5_outputs(89) <= not a;
    layer5_outputs(90) <= '0';
    layer5_outputs(91) <= a and not b;
    layer5_outputs(92) <= b and not a;
    layer5_outputs(93) <= not a;
    layer5_outputs(94) <= not b;
    layer5_outputs(95) <= a;
    layer5_outputs(96) <= a and b;
    layer5_outputs(97) <= not b or a;
    layer5_outputs(98) <= not a;
    layer5_outputs(99) <= '1';
    layer5_outputs(100) <= not (a and b);
    layer5_outputs(101) <= a or b;
    layer5_outputs(102) <= a and b;
    layer5_outputs(103) <= not a;
    layer5_outputs(104) <= not b or a;
    layer5_outputs(105) <= not (a and b);
    layer5_outputs(106) <= b and not a;
    layer5_outputs(107) <= a and not b;
    layer5_outputs(108) <= not b or a;
    layer5_outputs(109) <= not b;
    layer5_outputs(110) <= a and b;
    layer5_outputs(111) <= not (a and b);
    layer5_outputs(112) <= not b;
    layer5_outputs(113) <= b;
    layer5_outputs(114) <= a and b;
    layer5_outputs(115) <= b;
    layer5_outputs(116) <= b and not a;
    layer5_outputs(117) <= b;
    layer5_outputs(118) <= b and not a;
    layer5_outputs(119) <= '1';
    layer5_outputs(120) <= not a or b;
    layer5_outputs(121) <= a or b;
    layer5_outputs(122) <= '0';
    layer5_outputs(123) <= not a or b;
    layer5_outputs(124) <= '1';
    layer5_outputs(125) <= a and not b;
    layer5_outputs(126) <= b and not a;
    layer5_outputs(127) <= not a;
    layer5_outputs(128) <= a and b;
    layer5_outputs(129) <= a and not b;
    layer5_outputs(130) <= not (a xor b);
    layer5_outputs(131) <= not a;
    layer5_outputs(132) <= not b;
    layer5_outputs(133) <= not a;
    layer5_outputs(134) <= not a;
    layer5_outputs(135) <= a and not b;
    layer5_outputs(136) <= a and b;
    layer5_outputs(137) <= not (a and b);
    layer5_outputs(138) <= not b;
    layer5_outputs(139) <= a;
    layer5_outputs(140) <= not b or a;
    layer5_outputs(141) <= b;
    layer5_outputs(142) <= a or b;
    layer5_outputs(143) <= not (a xor b);
    layer5_outputs(144) <= not a;
    layer5_outputs(145) <= a and not b;
    layer5_outputs(146) <= b;
    layer5_outputs(147) <= not a;
    layer5_outputs(148) <= not b;
    layer5_outputs(149) <= not (a xor b);
    layer5_outputs(150) <= b and not a;
    layer5_outputs(151) <= not b or a;
    layer5_outputs(152) <= b;
    layer5_outputs(153) <= a xor b;
    layer5_outputs(154) <= not b;
    layer5_outputs(155) <= a;
    layer5_outputs(156) <= '0';
    layer5_outputs(157) <= a and b;
    layer5_outputs(158) <= not (a or b);
    layer5_outputs(159) <= not b;
    layer5_outputs(160) <= a and b;
    layer5_outputs(161) <= b;
    layer5_outputs(162) <= not a or b;
    layer5_outputs(163) <= b;
    layer5_outputs(164) <= not a or b;
    layer5_outputs(165) <= a and b;
    layer5_outputs(166) <= a or b;
    layer5_outputs(167) <= a or b;
    layer5_outputs(168) <= not b;
    layer5_outputs(169) <= b and not a;
    layer5_outputs(170) <= b and not a;
    layer5_outputs(171) <= b;
    layer5_outputs(172) <= a or b;
    layer5_outputs(173) <= b and not a;
    layer5_outputs(174) <= not b or a;
    layer5_outputs(175) <= not (a xor b);
    layer5_outputs(176) <= b and not a;
    layer5_outputs(177) <= a and b;
    layer5_outputs(178) <= not b;
    layer5_outputs(179) <= b;
    layer5_outputs(180) <= not a;
    layer5_outputs(181) <= not a;
    layer5_outputs(182) <= not b;
    layer5_outputs(183) <= a xor b;
    layer5_outputs(184) <= not (a or b);
    layer5_outputs(185) <= not (a or b);
    layer5_outputs(186) <= not b;
    layer5_outputs(187) <= a or b;
    layer5_outputs(188) <= '0';
    layer5_outputs(189) <= not a;
    layer5_outputs(190) <= b;
    layer5_outputs(191) <= '1';
    layer5_outputs(192) <= a;
    layer5_outputs(193) <= not (a and b);
    layer5_outputs(194) <= not (a or b);
    layer5_outputs(195) <= not (a xor b);
    layer5_outputs(196) <= not (a xor b);
    layer5_outputs(197) <= not a;
    layer5_outputs(198) <= not (a or b);
    layer5_outputs(199) <= '1';
    layer5_outputs(200) <= not a;
    layer5_outputs(201) <= not (a xor b);
    layer5_outputs(202) <= a or b;
    layer5_outputs(203) <= a or b;
    layer5_outputs(204) <= not (a and b);
    layer5_outputs(205) <= not (a xor b);
    layer5_outputs(206) <= not b or a;
    layer5_outputs(207) <= not b;
    layer5_outputs(208) <= '1';
    layer5_outputs(209) <= not a;
    layer5_outputs(210) <= a or b;
    layer5_outputs(211) <= '0';
    layer5_outputs(212) <= not (a or b);
    layer5_outputs(213) <= a xor b;
    layer5_outputs(214) <= '1';
    layer5_outputs(215) <= not (a and b);
    layer5_outputs(216) <= b and not a;
    layer5_outputs(217) <= b and not a;
    layer5_outputs(218) <= not a or b;
    layer5_outputs(219) <= a or b;
    layer5_outputs(220) <= not b;
    layer5_outputs(221) <= a xor b;
    layer5_outputs(222) <= not (a or b);
    layer5_outputs(223) <= a xor b;
    layer5_outputs(224) <= not a or b;
    layer5_outputs(225) <= a;
    layer5_outputs(226) <= b;
    layer5_outputs(227) <= not b or a;
    layer5_outputs(228) <= '0';
    layer5_outputs(229) <= a or b;
    layer5_outputs(230) <= not b or a;
    layer5_outputs(231) <= a and not b;
    layer5_outputs(232) <= b;
    layer5_outputs(233) <= not (a xor b);
    layer5_outputs(234) <= not a or b;
    layer5_outputs(235) <= a;
    layer5_outputs(236) <= b;
    layer5_outputs(237) <= b and not a;
    layer5_outputs(238) <= not b or a;
    layer5_outputs(239) <= a xor b;
    layer5_outputs(240) <= a or b;
    layer5_outputs(241) <= a and b;
    layer5_outputs(242) <= b;
    layer5_outputs(243) <= not b;
    layer5_outputs(244) <= not a or b;
    layer5_outputs(245) <= not b or a;
    layer5_outputs(246) <= not b;
    layer5_outputs(247) <= a and not b;
    layer5_outputs(248) <= not a;
    layer5_outputs(249) <= '1';
    layer5_outputs(250) <= not a;
    layer5_outputs(251) <= not (a or b);
    layer5_outputs(252) <= a or b;
    layer5_outputs(253) <= a or b;
    layer5_outputs(254) <= a and not b;
    layer5_outputs(255) <= a and not b;
    layer5_outputs(256) <= a and b;
    layer5_outputs(257) <= not b or a;
    layer5_outputs(258) <= a and b;
    layer5_outputs(259) <= a or b;
    layer5_outputs(260) <= not (a or b);
    layer5_outputs(261) <= a and not b;
    layer5_outputs(262) <= b;
    layer5_outputs(263) <= a;
    layer5_outputs(264) <= a xor b;
    layer5_outputs(265) <= not a or b;
    layer5_outputs(266) <= b;
    layer5_outputs(267) <= not b;
    layer5_outputs(268) <= not b;
    layer5_outputs(269) <= not (a and b);
    layer5_outputs(270) <= b;
    layer5_outputs(271) <= not a;
    layer5_outputs(272) <= a;
    layer5_outputs(273) <= a;
    layer5_outputs(274) <= not b or a;
    layer5_outputs(275) <= a and not b;
    layer5_outputs(276) <= '1';
    layer5_outputs(277) <= '1';
    layer5_outputs(278) <= not a;
    layer5_outputs(279) <= a and not b;
    layer5_outputs(280) <= not b;
    layer5_outputs(281) <= not a;
    layer5_outputs(282) <= not (a or b);
    layer5_outputs(283) <= a;
    layer5_outputs(284) <= not b;
    layer5_outputs(285) <= not b;
    layer5_outputs(286) <= b;
    layer5_outputs(287) <= a and b;
    layer5_outputs(288) <= not a or b;
    layer5_outputs(289) <= not b or a;
    layer5_outputs(290) <= a xor b;
    layer5_outputs(291) <= b;
    layer5_outputs(292) <= b;
    layer5_outputs(293) <= not a;
    layer5_outputs(294) <= not a or b;
    layer5_outputs(295) <= not b or a;
    layer5_outputs(296) <= b;
    layer5_outputs(297) <= not (a or b);
    layer5_outputs(298) <= not a;
    layer5_outputs(299) <= a;
    layer5_outputs(300) <= a xor b;
    layer5_outputs(301) <= not (a and b);
    layer5_outputs(302) <= not a or b;
    layer5_outputs(303) <= not a or b;
    layer5_outputs(304) <= a and b;
    layer5_outputs(305) <= not b;
    layer5_outputs(306) <= b and not a;
    layer5_outputs(307) <= b;
    layer5_outputs(308) <= not (a and b);
    layer5_outputs(309) <= b;
    layer5_outputs(310) <= b and not a;
    layer5_outputs(311) <= not (a or b);
    layer5_outputs(312) <= a or b;
    layer5_outputs(313) <= not (a and b);
    layer5_outputs(314) <= not (a xor b);
    layer5_outputs(315) <= '0';
    layer5_outputs(316) <= not a or b;
    layer5_outputs(317) <= not (a xor b);
    layer5_outputs(318) <= a or b;
    layer5_outputs(319) <= a and b;
    layer5_outputs(320) <= a and b;
    layer5_outputs(321) <= a;
    layer5_outputs(322) <= a and b;
    layer5_outputs(323) <= b;
    layer5_outputs(324) <= a xor b;
    layer5_outputs(325) <= not (a xor b);
    layer5_outputs(326) <= not (a or b);
    layer5_outputs(327) <= a;
    layer5_outputs(328) <= not a or b;
    layer5_outputs(329) <= not a;
    layer5_outputs(330) <= a and b;
    layer5_outputs(331) <= '1';
    layer5_outputs(332) <= a;
    layer5_outputs(333) <= not (a xor b);
    layer5_outputs(334) <= not a;
    layer5_outputs(335) <= not (a or b);
    layer5_outputs(336) <= a;
    layer5_outputs(337) <= not b;
    layer5_outputs(338) <= a or b;
    layer5_outputs(339) <= a and not b;
    layer5_outputs(340) <= not (a and b);
    layer5_outputs(341) <= '0';
    layer5_outputs(342) <= not b or a;
    layer5_outputs(343) <= not b or a;
    layer5_outputs(344) <= '0';
    layer5_outputs(345) <= not (a or b);
    layer5_outputs(346) <= a or b;
    layer5_outputs(347) <= a;
    layer5_outputs(348) <= a and not b;
    layer5_outputs(349) <= not a or b;
    layer5_outputs(350) <= b and not a;
    layer5_outputs(351) <= not (a or b);
    layer5_outputs(352) <= not a;
    layer5_outputs(353) <= not (a or b);
    layer5_outputs(354) <= not a;
    layer5_outputs(355) <= a and not b;
    layer5_outputs(356) <= not a or b;
    layer5_outputs(357) <= a;
    layer5_outputs(358) <= b;
    layer5_outputs(359) <= b;
    layer5_outputs(360) <= not (a xor b);
    layer5_outputs(361) <= not (a and b);
    layer5_outputs(362) <= a or b;
    layer5_outputs(363) <= not b;
    layer5_outputs(364) <= a and not b;
    layer5_outputs(365) <= not (a xor b);
    layer5_outputs(366) <= not (a or b);
    layer5_outputs(367) <= a and b;
    layer5_outputs(368) <= a or b;
    layer5_outputs(369) <= not (a and b);
    layer5_outputs(370) <= b;
    layer5_outputs(371) <= not a;
    layer5_outputs(372) <= '1';
    layer5_outputs(373) <= a and not b;
    layer5_outputs(374) <= b and not a;
    layer5_outputs(375) <= a or b;
    layer5_outputs(376) <= not b or a;
    layer5_outputs(377) <= not (a or b);
    layer5_outputs(378) <= a and b;
    layer5_outputs(379) <= a and b;
    layer5_outputs(380) <= a xor b;
    layer5_outputs(381) <= a and not b;
    layer5_outputs(382) <= a and b;
    layer5_outputs(383) <= a and b;
    layer5_outputs(384) <= not b;
    layer5_outputs(385) <= not (a or b);
    layer5_outputs(386) <= a and not b;
    layer5_outputs(387) <= not a;
    layer5_outputs(388) <= a;
    layer5_outputs(389) <= not (a or b);
    layer5_outputs(390) <= a and not b;
    layer5_outputs(391) <= a;
    layer5_outputs(392) <= not a;
    layer5_outputs(393) <= not a or b;
    layer5_outputs(394) <= a or b;
    layer5_outputs(395) <= a;
    layer5_outputs(396) <= a or b;
    layer5_outputs(397) <= b and not a;
    layer5_outputs(398) <= not a;
    layer5_outputs(399) <= a;
    layer5_outputs(400) <= not (a and b);
    layer5_outputs(401) <= not (a and b);
    layer5_outputs(402) <= a and not b;
    layer5_outputs(403) <= not (a xor b);
    layer5_outputs(404) <= a;
    layer5_outputs(405) <= a and not b;
    layer5_outputs(406) <= not (a xor b);
    layer5_outputs(407) <= b and not a;
    layer5_outputs(408) <= '1';
    layer5_outputs(409) <= not a;
    layer5_outputs(410) <= a and b;
    layer5_outputs(411) <= '0';
    layer5_outputs(412) <= a or b;
    layer5_outputs(413) <= not a;
    layer5_outputs(414) <= a;
    layer5_outputs(415) <= a or b;
    layer5_outputs(416) <= a and not b;
    layer5_outputs(417) <= a and not b;
    layer5_outputs(418) <= not a or b;
    layer5_outputs(419) <= not b;
    layer5_outputs(420) <= not (a and b);
    layer5_outputs(421) <= not b;
    layer5_outputs(422) <= not (a xor b);
    layer5_outputs(423) <= not (a and b);
    layer5_outputs(424) <= b;
    layer5_outputs(425) <= not (a and b);
    layer5_outputs(426) <= not b;
    layer5_outputs(427) <= a xor b;
    layer5_outputs(428) <= a and not b;
    layer5_outputs(429) <= '1';
    layer5_outputs(430) <= a and b;
    layer5_outputs(431) <= '1';
    layer5_outputs(432) <= a;
    layer5_outputs(433) <= b;
    layer5_outputs(434) <= not b or a;
    layer5_outputs(435) <= not (a xor b);
    layer5_outputs(436) <= a;
    layer5_outputs(437) <= not a or b;
    layer5_outputs(438) <= b and not a;
    layer5_outputs(439) <= not (a and b);
    layer5_outputs(440) <= a and not b;
    layer5_outputs(441) <= not a;
    layer5_outputs(442) <= a and not b;
    layer5_outputs(443) <= not a;
    layer5_outputs(444) <= not b;
    layer5_outputs(445) <= not a;
    layer5_outputs(446) <= b and not a;
    layer5_outputs(447) <= a and not b;
    layer5_outputs(448) <= not (a xor b);
    layer5_outputs(449) <= not a or b;
    layer5_outputs(450) <= a;
    layer5_outputs(451) <= '1';
    layer5_outputs(452) <= not a;
    layer5_outputs(453) <= not a;
    layer5_outputs(454) <= b;
    layer5_outputs(455) <= '0';
    layer5_outputs(456) <= a xor b;
    layer5_outputs(457) <= a;
    layer5_outputs(458) <= not b or a;
    layer5_outputs(459) <= not a or b;
    layer5_outputs(460) <= a and b;
    layer5_outputs(461) <= not a;
    layer5_outputs(462) <= a and b;
    layer5_outputs(463) <= not (a xor b);
    layer5_outputs(464) <= '0';
    layer5_outputs(465) <= b;
    layer5_outputs(466) <= not (a or b);
    layer5_outputs(467) <= a or b;
    layer5_outputs(468) <= a and b;
    layer5_outputs(469) <= b;
    layer5_outputs(470) <= b;
    layer5_outputs(471) <= a and b;
    layer5_outputs(472) <= '0';
    layer5_outputs(473) <= not b;
    layer5_outputs(474) <= not b;
    layer5_outputs(475) <= a;
    layer5_outputs(476) <= a and not b;
    layer5_outputs(477) <= not (a xor b);
    layer5_outputs(478) <= not b or a;
    layer5_outputs(479) <= not b;
    layer5_outputs(480) <= not (a and b);
    layer5_outputs(481) <= '0';
    layer5_outputs(482) <= a;
    layer5_outputs(483) <= a and not b;
    layer5_outputs(484) <= a xor b;
    layer5_outputs(485) <= a and b;
    layer5_outputs(486) <= a;
    layer5_outputs(487) <= not b;
    layer5_outputs(488) <= not b;
    layer5_outputs(489) <= not b or a;
    layer5_outputs(490) <= not b or a;
    layer5_outputs(491) <= b;
    layer5_outputs(492) <= a and b;
    layer5_outputs(493) <= a and not b;
    layer5_outputs(494) <= not (a and b);
    layer5_outputs(495) <= a;
    layer5_outputs(496) <= a;
    layer5_outputs(497) <= a and b;
    layer5_outputs(498) <= a;
    layer5_outputs(499) <= not b or a;
    layer5_outputs(500) <= not b;
    layer5_outputs(501) <= a;
    layer5_outputs(502) <= a and not b;
    layer5_outputs(503) <= not b or a;
    layer5_outputs(504) <= a and not b;
    layer5_outputs(505) <= a xor b;
    layer5_outputs(506) <= not b;
    layer5_outputs(507) <= a and not b;
    layer5_outputs(508) <= '0';
    layer5_outputs(509) <= a or b;
    layer5_outputs(510) <= not b;
    layer5_outputs(511) <= b and not a;
    layer5_outputs(512) <= a or b;
    layer5_outputs(513) <= not a;
    layer5_outputs(514) <= not b or a;
    layer5_outputs(515) <= a;
    layer5_outputs(516) <= not b;
    layer5_outputs(517) <= not a or b;
    layer5_outputs(518) <= not b;
    layer5_outputs(519) <= not a;
    layer5_outputs(520) <= not b;
    layer5_outputs(521) <= b;
    layer5_outputs(522) <= not b;
    layer5_outputs(523) <= a;
    layer5_outputs(524) <= b;
    layer5_outputs(525) <= not (a or b);
    layer5_outputs(526) <= '1';
    layer5_outputs(527) <= not (a and b);
    layer5_outputs(528) <= not b or a;
    layer5_outputs(529) <= not b;
    layer5_outputs(530) <= a and not b;
    layer5_outputs(531) <= a and b;
    layer5_outputs(532) <= a;
    layer5_outputs(533) <= not a;
    layer5_outputs(534) <= b;
    layer5_outputs(535) <= a and b;
    layer5_outputs(536) <= not a;
    layer5_outputs(537) <= a or b;
    layer5_outputs(538) <= not (a xor b);
    layer5_outputs(539) <= a;
    layer5_outputs(540) <= not b;
    layer5_outputs(541) <= b and not a;
    layer5_outputs(542) <= a;
    layer5_outputs(543) <= not b or a;
    layer5_outputs(544) <= '1';
    layer5_outputs(545) <= not b or a;
    layer5_outputs(546) <= not (a xor b);
    layer5_outputs(547) <= '1';
    layer5_outputs(548) <= a;
    layer5_outputs(549) <= not a or b;
    layer5_outputs(550) <= '0';
    layer5_outputs(551) <= not b;
    layer5_outputs(552) <= b;
    layer5_outputs(553) <= a xor b;
    layer5_outputs(554) <= a;
    layer5_outputs(555) <= not a or b;
    layer5_outputs(556) <= not a or b;
    layer5_outputs(557) <= b and not a;
    layer5_outputs(558) <= '1';
    layer5_outputs(559) <= b;
    layer5_outputs(560) <= not a or b;
    layer5_outputs(561) <= a and not b;
    layer5_outputs(562) <= not (a and b);
    layer5_outputs(563) <= not b;
    layer5_outputs(564) <= b;
    layer5_outputs(565) <= not a or b;
    layer5_outputs(566) <= a;
    layer5_outputs(567) <= not (a xor b);
    layer5_outputs(568) <= a or b;
    layer5_outputs(569) <= b;
    layer5_outputs(570) <= b and not a;
    layer5_outputs(571) <= not b;
    layer5_outputs(572) <= b;
    layer5_outputs(573) <= not (a and b);
    layer5_outputs(574) <= not b;
    layer5_outputs(575) <= not a;
    layer5_outputs(576) <= a and not b;
    layer5_outputs(577) <= a and not b;
    layer5_outputs(578) <= not a or b;
    layer5_outputs(579) <= a;
    layer5_outputs(580) <= not b or a;
    layer5_outputs(581) <= not a;
    layer5_outputs(582) <= a;
    layer5_outputs(583) <= not b or a;
    layer5_outputs(584) <= not b;
    layer5_outputs(585) <= not (a and b);
    layer5_outputs(586) <= not (a xor b);
    layer5_outputs(587) <= not a;
    layer5_outputs(588) <= not a;
    layer5_outputs(589) <= not b or a;
    layer5_outputs(590) <= a;
    layer5_outputs(591) <= a or b;
    layer5_outputs(592) <= not a or b;
    layer5_outputs(593) <= b;
    layer5_outputs(594) <= not a;
    layer5_outputs(595) <= a and b;
    layer5_outputs(596) <= not (a and b);
    layer5_outputs(597) <= not (a or b);
    layer5_outputs(598) <= b;
    layer5_outputs(599) <= not a;
    layer5_outputs(600) <= not (a or b);
    layer5_outputs(601) <= b and not a;
    layer5_outputs(602) <= '0';
    layer5_outputs(603) <= a and b;
    layer5_outputs(604) <= not b;
    layer5_outputs(605) <= not b;
    layer5_outputs(606) <= b and not a;
    layer5_outputs(607) <= b;
    layer5_outputs(608) <= a;
    layer5_outputs(609) <= b;
    layer5_outputs(610) <= not a;
    layer5_outputs(611) <= not (a or b);
    layer5_outputs(612) <= not a;
    layer5_outputs(613) <= a xor b;
    layer5_outputs(614) <= b;
    layer5_outputs(615) <= not (a or b);
    layer5_outputs(616) <= a;
    layer5_outputs(617) <= not b or a;
    layer5_outputs(618) <= not (a xor b);
    layer5_outputs(619) <= not a;
    layer5_outputs(620) <= a and not b;
    layer5_outputs(621) <= b and not a;
    layer5_outputs(622) <= b;
    layer5_outputs(623) <= not b or a;
    layer5_outputs(624) <= not a or b;
    layer5_outputs(625) <= b and not a;
    layer5_outputs(626) <= a;
    layer5_outputs(627) <= not b;
    layer5_outputs(628) <= not a or b;
    layer5_outputs(629) <= not a or b;
    layer5_outputs(630) <= b;
    layer5_outputs(631) <= not b or a;
    layer5_outputs(632) <= not a or b;
    layer5_outputs(633) <= not a;
    layer5_outputs(634) <= a or b;
    layer5_outputs(635) <= not b or a;
    layer5_outputs(636) <= a or b;
    layer5_outputs(637) <= not a;
    layer5_outputs(638) <= a and b;
    layer5_outputs(639) <= a or b;
    layer5_outputs(640) <= not a;
    layer5_outputs(641) <= a or b;
    layer5_outputs(642) <= not a or b;
    layer5_outputs(643) <= b and not a;
    layer5_outputs(644) <= not a;
    layer5_outputs(645) <= not a;
    layer5_outputs(646) <= a and not b;
    layer5_outputs(647) <= not b or a;
    layer5_outputs(648) <= not (a or b);
    layer5_outputs(649) <= not b or a;
    layer5_outputs(650) <= b;
    layer5_outputs(651) <= a and not b;
    layer5_outputs(652) <= a and not b;
    layer5_outputs(653) <= '1';
    layer5_outputs(654) <= not (a xor b);
    layer5_outputs(655) <= a and b;
    layer5_outputs(656) <= not a;
    layer5_outputs(657) <= a or b;
    layer5_outputs(658) <= a xor b;
    layer5_outputs(659) <= b;
    layer5_outputs(660) <= not (a and b);
    layer5_outputs(661) <= not b;
    layer5_outputs(662) <= b;
    layer5_outputs(663) <= not (a and b);
    layer5_outputs(664) <= a;
    layer5_outputs(665) <= not b or a;
    layer5_outputs(666) <= '1';
    layer5_outputs(667) <= not b;
    layer5_outputs(668) <= a and b;
    layer5_outputs(669) <= not a or b;
    layer5_outputs(670) <= not a;
    layer5_outputs(671) <= not (a or b);
    layer5_outputs(672) <= '1';
    layer5_outputs(673) <= a and not b;
    layer5_outputs(674) <= '1';
    layer5_outputs(675) <= b;
    layer5_outputs(676) <= a;
    layer5_outputs(677) <= '1';
    layer5_outputs(678) <= a and not b;
    layer5_outputs(679) <= b and not a;
    layer5_outputs(680) <= not a or b;
    layer5_outputs(681) <= a and not b;
    layer5_outputs(682) <= a or b;
    layer5_outputs(683) <= a or b;
    layer5_outputs(684) <= a xor b;
    layer5_outputs(685) <= a or b;
    layer5_outputs(686) <= not (a xor b);
    layer5_outputs(687) <= not b;
    layer5_outputs(688) <= not (a xor b);
    layer5_outputs(689) <= not a;
    layer5_outputs(690) <= '0';
    layer5_outputs(691) <= '0';
    layer5_outputs(692) <= not (a or b);
    layer5_outputs(693) <= '1';
    layer5_outputs(694) <= a or b;
    layer5_outputs(695) <= b;
    layer5_outputs(696) <= not b;
    layer5_outputs(697) <= a and not b;
    layer5_outputs(698) <= a;
    layer5_outputs(699) <= a;
    layer5_outputs(700) <= not a;
    layer5_outputs(701) <= a or b;
    layer5_outputs(702) <= a xor b;
    layer5_outputs(703) <= a and not b;
    layer5_outputs(704) <= not (a or b);
    layer5_outputs(705) <= not b;
    layer5_outputs(706) <= not a or b;
    layer5_outputs(707) <= a and not b;
    layer5_outputs(708) <= not b;
    layer5_outputs(709) <= a and b;
    layer5_outputs(710) <= not a;
    layer5_outputs(711) <= not b or a;
    layer5_outputs(712) <= b;
    layer5_outputs(713) <= not (a or b);
    layer5_outputs(714) <= b;
    layer5_outputs(715) <= a;
    layer5_outputs(716) <= b;
    layer5_outputs(717) <= not (a xor b);
    layer5_outputs(718) <= not b or a;
    layer5_outputs(719) <= not a or b;
    layer5_outputs(720) <= not b;
    layer5_outputs(721) <= '1';
    layer5_outputs(722) <= not a;
    layer5_outputs(723) <= b;
    layer5_outputs(724) <= not (a or b);
    layer5_outputs(725) <= b and not a;
    layer5_outputs(726) <= not (a or b);
    layer5_outputs(727) <= a or b;
    layer5_outputs(728) <= not b;
    layer5_outputs(729) <= not b;
    layer5_outputs(730) <= not (a and b);
    layer5_outputs(731) <= not a;
    layer5_outputs(732) <= a xor b;
    layer5_outputs(733) <= not (a and b);
    layer5_outputs(734) <= a xor b;
    layer5_outputs(735) <= not (a or b);
    layer5_outputs(736) <= not b or a;
    layer5_outputs(737) <= a and not b;
    layer5_outputs(738) <= b and not a;
    layer5_outputs(739) <= a;
    layer5_outputs(740) <= b;
    layer5_outputs(741) <= b and not a;
    layer5_outputs(742) <= a;
    layer5_outputs(743) <= not a;
    layer5_outputs(744) <= not b;
    layer5_outputs(745) <= not (a and b);
    layer5_outputs(746) <= a;
    layer5_outputs(747) <= a and b;
    layer5_outputs(748) <= not a;
    layer5_outputs(749) <= b;
    layer5_outputs(750) <= a and b;
    layer5_outputs(751) <= a and b;
    layer5_outputs(752) <= b;
    layer5_outputs(753) <= not a or b;
    layer5_outputs(754) <= a or b;
    layer5_outputs(755) <= b and not a;
    layer5_outputs(756) <= '0';
    layer5_outputs(757) <= not a;
    layer5_outputs(758) <= not a;
    layer5_outputs(759) <= b and not a;
    layer5_outputs(760) <= b;
    layer5_outputs(761) <= not a;
    layer5_outputs(762) <= '1';
    layer5_outputs(763) <= a and b;
    layer5_outputs(764) <= a and b;
    layer5_outputs(765) <= not a;
    layer5_outputs(766) <= not (a or b);
    layer5_outputs(767) <= not b;
    layer5_outputs(768) <= a or b;
    layer5_outputs(769) <= '1';
    layer5_outputs(770) <= b;
    layer5_outputs(771) <= not (a or b);
    layer5_outputs(772) <= not a;
    layer5_outputs(773) <= not b or a;
    layer5_outputs(774) <= not (a or b);
    layer5_outputs(775) <= not (a and b);
    layer5_outputs(776) <= '1';
    layer5_outputs(777) <= '1';
    layer5_outputs(778) <= not (a xor b);
    layer5_outputs(779) <= not b or a;
    layer5_outputs(780) <= not a or b;
    layer5_outputs(781) <= b and not a;
    layer5_outputs(782) <= b;
    layer5_outputs(783) <= a and b;
    layer5_outputs(784) <= b;
    layer5_outputs(785) <= b and not a;
    layer5_outputs(786) <= a;
    layer5_outputs(787) <= a and b;
    layer5_outputs(788) <= not (a and b);
    layer5_outputs(789) <= a or b;
    layer5_outputs(790) <= '0';
    layer5_outputs(791) <= not b or a;
    layer5_outputs(792) <= '1';
    layer5_outputs(793) <= a;
    layer5_outputs(794) <= not (a or b);
    layer5_outputs(795) <= '1';
    layer5_outputs(796) <= not (a or b);
    layer5_outputs(797) <= not b or a;
    layer5_outputs(798) <= a and b;
    layer5_outputs(799) <= not a or b;
    layer5_outputs(800) <= not (a and b);
    layer5_outputs(801) <= a or b;
    layer5_outputs(802) <= '1';
    layer5_outputs(803) <= a and b;
    layer5_outputs(804) <= b and not a;
    layer5_outputs(805) <= '1';
    layer5_outputs(806) <= not (a and b);
    layer5_outputs(807) <= not (a and b);
    layer5_outputs(808) <= not b;
    layer5_outputs(809) <= b and not a;
    layer5_outputs(810) <= a and b;
    layer5_outputs(811) <= not (a or b);
    layer5_outputs(812) <= not b;
    layer5_outputs(813) <= not (a or b);
    layer5_outputs(814) <= a xor b;
    layer5_outputs(815) <= not (a or b);
    layer5_outputs(816) <= b;
    layer5_outputs(817) <= b;
    layer5_outputs(818) <= not a;
    layer5_outputs(819) <= a and b;
    layer5_outputs(820) <= '0';
    layer5_outputs(821) <= a;
    layer5_outputs(822) <= not b;
    layer5_outputs(823) <= b;
    layer5_outputs(824) <= a and b;
    layer5_outputs(825) <= a;
    layer5_outputs(826) <= a or b;
    layer5_outputs(827) <= b;
    layer5_outputs(828) <= not a or b;
    layer5_outputs(829) <= a and b;
    layer5_outputs(830) <= not b;
    layer5_outputs(831) <= a;
    layer5_outputs(832) <= not a;
    layer5_outputs(833) <= '1';
    layer5_outputs(834) <= not b or a;
    layer5_outputs(835) <= a;
    layer5_outputs(836) <= '0';
    layer5_outputs(837) <= not a or b;
    layer5_outputs(838) <= a xor b;
    layer5_outputs(839) <= not a;
    layer5_outputs(840) <= a;
    layer5_outputs(841) <= b;
    layer5_outputs(842) <= not b or a;
    layer5_outputs(843) <= not b or a;
    layer5_outputs(844) <= a and b;
    layer5_outputs(845) <= a and b;
    layer5_outputs(846) <= a;
    layer5_outputs(847) <= b and not a;
    layer5_outputs(848) <= b and not a;
    layer5_outputs(849) <= not a;
    layer5_outputs(850) <= not b;
    layer5_outputs(851) <= not (a and b);
    layer5_outputs(852) <= a xor b;
    layer5_outputs(853) <= b and not a;
    layer5_outputs(854) <= not (a xor b);
    layer5_outputs(855) <= a or b;
    layer5_outputs(856) <= a;
    layer5_outputs(857) <= b;
    layer5_outputs(858) <= not b;
    layer5_outputs(859) <= a and b;
    layer5_outputs(860) <= a and not b;
    layer5_outputs(861) <= not a;
    layer5_outputs(862) <= a or b;
    layer5_outputs(863) <= b;
    layer5_outputs(864) <= not b or a;
    layer5_outputs(865) <= not a;
    layer5_outputs(866) <= not a or b;
    layer5_outputs(867) <= '1';
    layer5_outputs(868) <= a xor b;
    layer5_outputs(869) <= not b;
    layer5_outputs(870) <= b and not a;
    layer5_outputs(871) <= b and not a;
    layer5_outputs(872) <= a and b;
    layer5_outputs(873) <= not b;
    layer5_outputs(874) <= b;
    layer5_outputs(875) <= not (a and b);
    layer5_outputs(876) <= a;
    layer5_outputs(877) <= not a;
    layer5_outputs(878) <= a and b;
    layer5_outputs(879) <= a and b;
    layer5_outputs(880) <= '0';
    layer5_outputs(881) <= b;
    layer5_outputs(882) <= not a or b;
    layer5_outputs(883) <= not b or a;
    layer5_outputs(884) <= not (a or b);
    layer5_outputs(885) <= not a or b;
    layer5_outputs(886) <= '1';
    layer5_outputs(887) <= b and not a;
    layer5_outputs(888) <= a and b;
    layer5_outputs(889) <= b;
    layer5_outputs(890) <= not (a and b);
    layer5_outputs(891) <= '0';
    layer5_outputs(892) <= a;
    layer5_outputs(893) <= a and not b;
    layer5_outputs(894) <= not b or a;
    layer5_outputs(895) <= b and not a;
    layer5_outputs(896) <= not (a xor b);
    layer5_outputs(897) <= not b;
    layer5_outputs(898) <= not b;
    layer5_outputs(899) <= not b or a;
    layer5_outputs(900) <= b;
    layer5_outputs(901) <= not a or b;
    layer5_outputs(902) <= not a or b;
    layer5_outputs(903) <= a and not b;
    layer5_outputs(904) <= a xor b;
    layer5_outputs(905) <= '1';
    layer5_outputs(906) <= '0';
    layer5_outputs(907) <= b and not a;
    layer5_outputs(908) <= a and not b;
    layer5_outputs(909) <= not b or a;
    layer5_outputs(910) <= not b or a;
    layer5_outputs(911) <= not a or b;
    layer5_outputs(912) <= b;
    layer5_outputs(913) <= a xor b;
    layer5_outputs(914) <= '0';
    layer5_outputs(915) <= a and b;
    layer5_outputs(916) <= a or b;
    layer5_outputs(917) <= a;
    layer5_outputs(918) <= b and not a;
    layer5_outputs(919) <= not b or a;
    layer5_outputs(920) <= not a or b;
    layer5_outputs(921) <= not a;
    layer5_outputs(922) <= not a;
    layer5_outputs(923) <= not b or a;
    layer5_outputs(924) <= not b or a;
    layer5_outputs(925) <= not b;
    layer5_outputs(926) <= a and not b;
    layer5_outputs(927) <= not b;
    layer5_outputs(928) <= a;
    layer5_outputs(929) <= '0';
    layer5_outputs(930) <= not b or a;
    layer5_outputs(931) <= a xor b;
    layer5_outputs(932) <= a;
    layer5_outputs(933) <= a and not b;
    layer5_outputs(934) <= a;
    layer5_outputs(935) <= not a or b;
    layer5_outputs(936) <= not b;
    layer5_outputs(937) <= not b or a;
    layer5_outputs(938) <= a xor b;
    layer5_outputs(939) <= a or b;
    layer5_outputs(940) <= a and not b;
    layer5_outputs(941) <= not b;
    layer5_outputs(942) <= '1';
    layer5_outputs(943) <= not (a or b);
    layer5_outputs(944) <= not (a and b);
    layer5_outputs(945) <= b;
    layer5_outputs(946) <= a;
    layer5_outputs(947) <= not a;
    layer5_outputs(948) <= a;
    layer5_outputs(949) <= a;
    layer5_outputs(950) <= not a;
    layer5_outputs(951) <= not (a or b);
    layer5_outputs(952) <= not (a and b);
    layer5_outputs(953) <= not a;
    layer5_outputs(954) <= not a;
    layer5_outputs(955) <= a;
    layer5_outputs(956) <= b;
    layer5_outputs(957) <= a;
    layer5_outputs(958) <= a and not b;
    layer5_outputs(959) <= not (a or b);
    layer5_outputs(960) <= a or b;
    layer5_outputs(961) <= not a;
    layer5_outputs(962) <= not a or b;
    layer5_outputs(963) <= not (a and b);
    layer5_outputs(964) <= not b or a;
    layer5_outputs(965) <= not (a and b);
    layer5_outputs(966) <= not b or a;
    layer5_outputs(967) <= not a;
    layer5_outputs(968) <= a xor b;
    layer5_outputs(969) <= not a or b;
    layer5_outputs(970) <= not b;
    layer5_outputs(971) <= a and b;
    layer5_outputs(972) <= not b;
    layer5_outputs(973) <= b;
    layer5_outputs(974) <= not (a or b);
    layer5_outputs(975) <= b;
    layer5_outputs(976) <= not a;
    layer5_outputs(977) <= not a;
    layer5_outputs(978) <= a;
    layer5_outputs(979) <= not a;
    layer5_outputs(980) <= b and not a;
    layer5_outputs(981) <= not b;
    layer5_outputs(982) <= not b;
    layer5_outputs(983) <= b;
    layer5_outputs(984) <= not b or a;
    layer5_outputs(985) <= b;
    layer5_outputs(986) <= a;
    layer5_outputs(987) <= a;
    layer5_outputs(988) <= not (a and b);
    layer5_outputs(989) <= a;
    layer5_outputs(990) <= not b;
    layer5_outputs(991) <= b and not a;
    layer5_outputs(992) <= not (a xor b);
    layer5_outputs(993) <= not b;
    layer5_outputs(994) <= not (a or b);
    layer5_outputs(995) <= not (a and b);
    layer5_outputs(996) <= not b;
    layer5_outputs(997) <= b and not a;
    layer5_outputs(998) <= b and not a;
    layer5_outputs(999) <= b;
    layer5_outputs(1000) <= a and b;
    layer5_outputs(1001) <= not b or a;
    layer5_outputs(1002) <= a or b;
    layer5_outputs(1003) <= '0';
    layer5_outputs(1004) <= not (a xor b);
    layer5_outputs(1005) <= not a;
    layer5_outputs(1006) <= a and not b;
    layer5_outputs(1007) <= not (a or b);
    layer5_outputs(1008) <= not (a or b);
    layer5_outputs(1009) <= not (a and b);
    layer5_outputs(1010) <= b;
    layer5_outputs(1011) <= not (a xor b);
    layer5_outputs(1012) <= a;
    layer5_outputs(1013) <= not b or a;
    layer5_outputs(1014) <= b and not a;
    layer5_outputs(1015) <= a or b;
    layer5_outputs(1016) <= not (a and b);
    layer5_outputs(1017) <= not (a and b);
    layer5_outputs(1018) <= a and not b;
    layer5_outputs(1019) <= a and not b;
    layer5_outputs(1020) <= not b;
    layer5_outputs(1021) <= a;
    layer5_outputs(1022) <= not b or a;
    layer5_outputs(1023) <= a and b;
    layer5_outputs(1024) <= not (a xor b);
    layer5_outputs(1025) <= not b;
    layer5_outputs(1026) <= a and b;
    layer5_outputs(1027) <= not b;
    layer5_outputs(1028) <= not a or b;
    layer5_outputs(1029) <= a and b;
    layer5_outputs(1030) <= a or b;
    layer5_outputs(1031) <= '1';
    layer5_outputs(1032) <= not (a or b);
    layer5_outputs(1033) <= a and not b;
    layer5_outputs(1034) <= b and not a;
    layer5_outputs(1035) <= a and b;
    layer5_outputs(1036) <= b and not a;
    layer5_outputs(1037) <= not (a and b);
    layer5_outputs(1038) <= '1';
    layer5_outputs(1039) <= b;
    layer5_outputs(1040) <= not b or a;
    layer5_outputs(1041) <= a;
    layer5_outputs(1042) <= b;
    layer5_outputs(1043) <= a xor b;
    layer5_outputs(1044) <= a;
    layer5_outputs(1045) <= b and not a;
    layer5_outputs(1046) <= not (a or b);
    layer5_outputs(1047) <= a and not b;
    layer5_outputs(1048) <= not b;
    layer5_outputs(1049) <= not (a xor b);
    layer5_outputs(1050) <= not a or b;
    layer5_outputs(1051) <= b and not a;
    layer5_outputs(1052) <= not (a xor b);
    layer5_outputs(1053) <= not (a xor b);
    layer5_outputs(1054) <= not b;
    layer5_outputs(1055) <= not (a and b);
    layer5_outputs(1056) <= not b;
    layer5_outputs(1057) <= a;
    layer5_outputs(1058) <= b;
    layer5_outputs(1059) <= a;
    layer5_outputs(1060) <= a or b;
    layer5_outputs(1061) <= a and b;
    layer5_outputs(1062) <= a xor b;
    layer5_outputs(1063) <= a and b;
    layer5_outputs(1064) <= b;
    layer5_outputs(1065) <= a xor b;
    layer5_outputs(1066) <= not a;
    layer5_outputs(1067) <= a;
    layer5_outputs(1068) <= '1';
    layer5_outputs(1069) <= not a;
    layer5_outputs(1070) <= not a;
    layer5_outputs(1071) <= not (a and b);
    layer5_outputs(1072) <= a and b;
    layer5_outputs(1073) <= b and not a;
    layer5_outputs(1074) <= not a;
    layer5_outputs(1075) <= not a or b;
    layer5_outputs(1076) <= not a;
    layer5_outputs(1077) <= not a or b;
    layer5_outputs(1078) <= not (a xor b);
    layer5_outputs(1079) <= b and not a;
    layer5_outputs(1080) <= b;
    layer5_outputs(1081) <= a and not b;
    layer5_outputs(1082) <= a;
    layer5_outputs(1083) <= not a or b;
    layer5_outputs(1084) <= b;
    layer5_outputs(1085) <= not b or a;
    layer5_outputs(1086) <= not b;
    layer5_outputs(1087) <= a and not b;
    layer5_outputs(1088) <= not a;
    layer5_outputs(1089) <= not b or a;
    layer5_outputs(1090) <= not a;
    layer5_outputs(1091) <= not a;
    layer5_outputs(1092) <= not a or b;
    layer5_outputs(1093) <= b;
    layer5_outputs(1094) <= a xor b;
    layer5_outputs(1095) <= b and not a;
    layer5_outputs(1096) <= a or b;
    layer5_outputs(1097) <= not a;
    layer5_outputs(1098) <= not a;
    layer5_outputs(1099) <= not (a or b);
    layer5_outputs(1100) <= '0';
    layer5_outputs(1101) <= b and not a;
    layer5_outputs(1102) <= not (a and b);
    layer5_outputs(1103) <= not a;
    layer5_outputs(1104) <= a and b;
    layer5_outputs(1105) <= not a;
    layer5_outputs(1106) <= not (a xor b);
    layer5_outputs(1107) <= not b or a;
    layer5_outputs(1108) <= not (a or b);
    layer5_outputs(1109) <= not (a and b);
    layer5_outputs(1110) <= a or b;
    layer5_outputs(1111) <= not b or a;
    layer5_outputs(1112) <= a;
    layer5_outputs(1113) <= not (a xor b);
    layer5_outputs(1114) <= not (a and b);
    layer5_outputs(1115) <= a;
    layer5_outputs(1116) <= not (a xor b);
    layer5_outputs(1117) <= a and b;
    layer5_outputs(1118) <= a;
    layer5_outputs(1119) <= not b or a;
    layer5_outputs(1120) <= a;
    layer5_outputs(1121) <= a xor b;
    layer5_outputs(1122) <= a or b;
    layer5_outputs(1123) <= not (a xor b);
    layer5_outputs(1124) <= not (a or b);
    layer5_outputs(1125) <= not (a xor b);
    layer5_outputs(1126) <= not b or a;
    layer5_outputs(1127) <= a;
    layer5_outputs(1128) <= b;
    layer5_outputs(1129) <= not b or a;
    layer5_outputs(1130) <= not a or b;
    layer5_outputs(1131) <= a and not b;
    layer5_outputs(1132) <= a and b;
    layer5_outputs(1133) <= not a or b;
    layer5_outputs(1134) <= not (a or b);
    layer5_outputs(1135) <= not (a xor b);
    layer5_outputs(1136) <= not (a xor b);
    layer5_outputs(1137) <= not (a and b);
    layer5_outputs(1138) <= a and not b;
    layer5_outputs(1139) <= not (a or b);
    layer5_outputs(1140) <= a;
    layer5_outputs(1141) <= not a;
    layer5_outputs(1142) <= a and b;
    layer5_outputs(1143) <= '0';
    layer5_outputs(1144) <= a or b;
    layer5_outputs(1145) <= not a;
    layer5_outputs(1146) <= a and not b;
    layer5_outputs(1147) <= not b or a;
    layer5_outputs(1148) <= not b;
    layer5_outputs(1149) <= not (a or b);
    layer5_outputs(1150) <= a;
    layer5_outputs(1151) <= not a;
    layer5_outputs(1152) <= not (a or b);
    layer5_outputs(1153) <= a and b;
    layer5_outputs(1154) <= a;
    layer5_outputs(1155) <= not a;
    layer5_outputs(1156) <= not a or b;
    layer5_outputs(1157) <= a;
    layer5_outputs(1158) <= a;
    layer5_outputs(1159) <= not b or a;
    layer5_outputs(1160) <= a or b;
    layer5_outputs(1161) <= a or b;
    layer5_outputs(1162) <= not (a or b);
    layer5_outputs(1163) <= not b;
    layer5_outputs(1164) <= not (a or b);
    layer5_outputs(1165) <= not (a or b);
    layer5_outputs(1166) <= not (a or b);
    layer5_outputs(1167) <= a;
    layer5_outputs(1168) <= a or b;
    layer5_outputs(1169) <= '0';
    layer5_outputs(1170) <= not (a xor b);
    layer5_outputs(1171) <= a;
    layer5_outputs(1172) <= b and not a;
    layer5_outputs(1173) <= a or b;
    layer5_outputs(1174) <= not b or a;
    layer5_outputs(1175) <= not (a or b);
    layer5_outputs(1176) <= b and not a;
    layer5_outputs(1177) <= not (a or b);
    layer5_outputs(1178) <= not b or a;
    layer5_outputs(1179) <= not (a or b);
    layer5_outputs(1180) <= a and not b;
    layer5_outputs(1181) <= b;
    layer5_outputs(1182) <= not b;
    layer5_outputs(1183) <= a and not b;
    layer5_outputs(1184) <= not (a xor b);
    layer5_outputs(1185) <= a;
    layer5_outputs(1186) <= not b;
    layer5_outputs(1187) <= not (a and b);
    layer5_outputs(1188) <= not (a or b);
    layer5_outputs(1189) <= not b or a;
    layer5_outputs(1190) <= a;
    layer5_outputs(1191) <= '1';
    layer5_outputs(1192) <= not (a or b);
    layer5_outputs(1193) <= not (a or b);
    layer5_outputs(1194) <= not a or b;
    layer5_outputs(1195) <= '0';
    layer5_outputs(1196) <= not (a or b);
    layer5_outputs(1197) <= b;
    layer5_outputs(1198) <= not (a or b);
    layer5_outputs(1199) <= not a or b;
    layer5_outputs(1200) <= b and not a;
    layer5_outputs(1201) <= a or b;
    layer5_outputs(1202) <= not a;
    layer5_outputs(1203) <= not b or a;
    layer5_outputs(1204) <= not a;
    layer5_outputs(1205) <= b;
    layer5_outputs(1206) <= not (a and b);
    layer5_outputs(1207) <= not (a xor b);
    layer5_outputs(1208) <= not a or b;
    layer5_outputs(1209) <= a and not b;
    layer5_outputs(1210) <= a;
    layer5_outputs(1211) <= b and not a;
    layer5_outputs(1212) <= '1';
    layer5_outputs(1213) <= a and not b;
    layer5_outputs(1214) <= a and b;
    layer5_outputs(1215) <= not (a and b);
    layer5_outputs(1216) <= '0';
    layer5_outputs(1217) <= a;
    layer5_outputs(1218) <= not b;
    layer5_outputs(1219) <= not a;
    layer5_outputs(1220) <= not a or b;
    layer5_outputs(1221) <= not a;
    layer5_outputs(1222) <= a xor b;
    layer5_outputs(1223) <= not (a xor b);
    layer5_outputs(1224) <= b;
    layer5_outputs(1225) <= not (a xor b);
    layer5_outputs(1226) <= not b or a;
    layer5_outputs(1227) <= a and not b;
    layer5_outputs(1228) <= a and b;
    layer5_outputs(1229) <= not (a or b);
    layer5_outputs(1230) <= not (a or b);
    layer5_outputs(1231) <= not a or b;
    layer5_outputs(1232) <= not (a and b);
    layer5_outputs(1233) <= not b;
    layer5_outputs(1234) <= not (a or b);
    layer5_outputs(1235) <= not a;
    layer5_outputs(1236) <= a;
    layer5_outputs(1237) <= b;
    layer5_outputs(1238) <= a xor b;
    layer5_outputs(1239) <= b and not a;
    layer5_outputs(1240) <= a;
    layer5_outputs(1241) <= a;
    layer5_outputs(1242) <= not b;
    layer5_outputs(1243) <= a and b;
    layer5_outputs(1244) <= a;
    layer5_outputs(1245) <= not b;
    layer5_outputs(1246) <= not a;
    layer5_outputs(1247) <= a;
    layer5_outputs(1248) <= not b;
    layer5_outputs(1249) <= '0';
    layer5_outputs(1250) <= not b or a;
    layer5_outputs(1251) <= not a;
    layer5_outputs(1252) <= not (a xor b);
    layer5_outputs(1253) <= not a;
    layer5_outputs(1254) <= b and not a;
    layer5_outputs(1255) <= a xor b;
    layer5_outputs(1256) <= a;
    layer5_outputs(1257) <= b and not a;
    layer5_outputs(1258) <= '0';
    layer5_outputs(1259) <= not (a and b);
    layer5_outputs(1260) <= not a;
    layer5_outputs(1261) <= '0';
    layer5_outputs(1262) <= not a or b;
    layer5_outputs(1263) <= a or b;
    layer5_outputs(1264) <= a xor b;
    layer5_outputs(1265) <= not a;
    layer5_outputs(1266) <= not b or a;
    layer5_outputs(1267) <= not a;
    layer5_outputs(1268) <= '1';
    layer5_outputs(1269) <= b and not a;
    layer5_outputs(1270) <= not a;
    layer5_outputs(1271) <= not a or b;
    layer5_outputs(1272) <= not a or b;
    layer5_outputs(1273) <= b;
    layer5_outputs(1274) <= '1';
    layer5_outputs(1275) <= a;
    layer5_outputs(1276) <= not b;
    layer5_outputs(1277) <= not b;
    layer5_outputs(1278) <= a and not b;
    layer5_outputs(1279) <= not a;
    layer5_outputs(1280) <= a;
    layer5_outputs(1281) <= not b;
    layer5_outputs(1282) <= b;
    layer5_outputs(1283) <= not (a or b);
    layer5_outputs(1284) <= not a;
    layer5_outputs(1285) <= a;
    layer5_outputs(1286) <= a;
    layer5_outputs(1287) <= not (a and b);
    layer5_outputs(1288) <= not a or b;
    layer5_outputs(1289) <= b and not a;
    layer5_outputs(1290) <= not (a or b);
    layer5_outputs(1291) <= not a or b;
    layer5_outputs(1292) <= b and not a;
    layer5_outputs(1293) <= '0';
    layer5_outputs(1294) <= not (a or b);
    layer5_outputs(1295) <= a xor b;
    layer5_outputs(1296) <= not b;
    layer5_outputs(1297) <= a and not b;
    layer5_outputs(1298) <= b;
    layer5_outputs(1299) <= a;
    layer5_outputs(1300) <= a and not b;
    layer5_outputs(1301) <= not a or b;
    layer5_outputs(1302) <= a;
    layer5_outputs(1303) <= a;
    layer5_outputs(1304) <= a and not b;
    layer5_outputs(1305) <= a and b;
    layer5_outputs(1306) <= b;
    layer5_outputs(1307) <= a;
    layer5_outputs(1308) <= a or b;
    layer5_outputs(1309) <= '1';
    layer5_outputs(1310) <= not (a xor b);
    layer5_outputs(1311) <= b;
    layer5_outputs(1312) <= b;
    layer5_outputs(1313) <= a xor b;
    layer5_outputs(1314) <= not (a or b);
    layer5_outputs(1315) <= not a or b;
    layer5_outputs(1316) <= not a;
    layer5_outputs(1317) <= not a or b;
    layer5_outputs(1318) <= not a;
    layer5_outputs(1319) <= a or b;
    layer5_outputs(1320) <= not (a and b);
    layer5_outputs(1321) <= a;
    layer5_outputs(1322) <= not a or b;
    layer5_outputs(1323) <= not b or a;
    layer5_outputs(1324) <= not (a or b);
    layer5_outputs(1325) <= not (a or b);
    layer5_outputs(1326) <= not (a or b);
    layer5_outputs(1327) <= a or b;
    layer5_outputs(1328) <= '0';
    layer5_outputs(1329) <= not a or b;
    layer5_outputs(1330) <= not a or b;
    layer5_outputs(1331) <= not b;
    layer5_outputs(1332) <= not b;
    layer5_outputs(1333) <= b;
    layer5_outputs(1334) <= not (a or b);
    layer5_outputs(1335) <= not (a xor b);
    layer5_outputs(1336) <= b and not a;
    layer5_outputs(1337) <= not a;
    layer5_outputs(1338) <= b;
    layer5_outputs(1339) <= not a or b;
    layer5_outputs(1340) <= not b;
    layer5_outputs(1341) <= not a;
    layer5_outputs(1342) <= a;
    layer5_outputs(1343) <= a;
    layer5_outputs(1344) <= a and not b;
    layer5_outputs(1345) <= not b;
    layer5_outputs(1346) <= a and not b;
    layer5_outputs(1347) <= a;
    layer5_outputs(1348) <= b and not a;
    layer5_outputs(1349) <= a or b;
    layer5_outputs(1350) <= not a or b;
    layer5_outputs(1351) <= not (a and b);
    layer5_outputs(1352) <= not (a or b);
    layer5_outputs(1353) <= not a or b;
    layer5_outputs(1354) <= not (a xor b);
    layer5_outputs(1355) <= not (a or b);
    layer5_outputs(1356) <= not (a and b);
    layer5_outputs(1357) <= a;
    layer5_outputs(1358) <= not a or b;
    layer5_outputs(1359) <= not (a or b);
    layer5_outputs(1360) <= not a;
    layer5_outputs(1361) <= not a;
    layer5_outputs(1362) <= '1';
    layer5_outputs(1363) <= not a;
    layer5_outputs(1364) <= a and b;
    layer5_outputs(1365) <= '0';
    layer5_outputs(1366) <= not b;
    layer5_outputs(1367) <= b;
    layer5_outputs(1368) <= a or b;
    layer5_outputs(1369) <= not a;
    layer5_outputs(1370) <= not b;
    layer5_outputs(1371) <= not b;
    layer5_outputs(1372) <= not (a and b);
    layer5_outputs(1373) <= a;
    layer5_outputs(1374) <= not a or b;
    layer5_outputs(1375) <= not a or b;
    layer5_outputs(1376) <= not a or b;
    layer5_outputs(1377) <= b and not a;
    layer5_outputs(1378) <= b;
    layer5_outputs(1379) <= b;
    layer5_outputs(1380) <= not a;
    layer5_outputs(1381) <= not (a or b);
    layer5_outputs(1382) <= a and b;
    layer5_outputs(1383) <= not a;
    layer5_outputs(1384) <= not a or b;
    layer5_outputs(1385) <= a;
    layer5_outputs(1386) <= not b or a;
    layer5_outputs(1387) <= a or b;
    layer5_outputs(1388) <= not b;
    layer5_outputs(1389) <= b;
    layer5_outputs(1390) <= not b;
    layer5_outputs(1391) <= not b;
    layer5_outputs(1392) <= a;
    layer5_outputs(1393) <= a or b;
    layer5_outputs(1394) <= a;
    layer5_outputs(1395) <= not (a and b);
    layer5_outputs(1396) <= a and not b;
    layer5_outputs(1397) <= not a or b;
    layer5_outputs(1398) <= not b;
    layer5_outputs(1399) <= a and not b;
    layer5_outputs(1400) <= a;
    layer5_outputs(1401) <= not (a xor b);
    layer5_outputs(1402) <= b;
    layer5_outputs(1403) <= not a;
    layer5_outputs(1404) <= not b;
    layer5_outputs(1405) <= not a or b;
    layer5_outputs(1406) <= a and not b;
    layer5_outputs(1407) <= not a;
    layer5_outputs(1408) <= not b;
    layer5_outputs(1409) <= a or b;
    layer5_outputs(1410) <= not b or a;
    layer5_outputs(1411) <= not a;
    layer5_outputs(1412) <= a or b;
    layer5_outputs(1413) <= a and not b;
    layer5_outputs(1414) <= '1';
    layer5_outputs(1415) <= a or b;
    layer5_outputs(1416) <= b;
    layer5_outputs(1417) <= not a or b;
    layer5_outputs(1418) <= '0';
    layer5_outputs(1419) <= b and not a;
    layer5_outputs(1420) <= not a;
    layer5_outputs(1421) <= b and not a;
    layer5_outputs(1422) <= a or b;
    layer5_outputs(1423) <= b and not a;
    layer5_outputs(1424) <= not (a and b);
    layer5_outputs(1425) <= b;
    layer5_outputs(1426) <= not b;
    layer5_outputs(1427) <= not (a and b);
    layer5_outputs(1428) <= not b or a;
    layer5_outputs(1429) <= '0';
    layer5_outputs(1430) <= not (a or b);
    layer5_outputs(1431) <= not a;
    layer5_outputs(1432) <= not b or a;
    layer5_outputs(1433) <= not a or b;
    layer5_outputs(1434) <= a and not b;
    layer5_outputs(1435) <= a and not b;
    layer5_outputs(1436) <= not a or b;
    layer5_outputs(1437) <= not (a or b);
    layer5_outputs(1438) <= not (a or b);
    layer5_outputs(1439) <= a or b;
    layer5_outputs(1440) <= a or b;
    layer5_outputs(1441) <= a or b;
    layer5_outputs(1442) <= b and not a;
    layer5_outputs(1443) <= a and b;
    layer5_outputs(1444) <= a and b;
    layer5_outputs(1445) <= not b or a;
    layer5_outputs(1446) <= not a or b;
    layer5_outputs(1447) <= '0';
    layer5_outputs(1448) <= not a or b;
    layer5_outputs(1449) <= a or b;
    layer5_outputs(1450) <= b;
    layer5_outputs(1451) <= '0';
    layer5_outputs(1452) <= a and not b;
    layer5_outputs(1453) <= b;
    layer5_outputs(1454) <= a or b;
    layer5_outputs(1455) <= not (a xor b);
    layer5_outputs(1456) <= not (a and b);
    layer5_outputs(1457) <= a and not b;
    layer5_outputs(1458) <= not a;
    layer5_outputs(1459) <= b and not a;
    layer5_outputs(1460) <= b;
    layer5_outputs(1461) <= not (a and b);
    layer5_outputs(1462) <= not b;
    layer5_outputs(1463) <= not (a and b);
    layer5_outputs(1464) <= not a;
    layer5_outputs(1465) <= not (a or b);
    layer5_outputs(1466) <= not b or a;
    layer5_outputs(1467) <= a;
    layer5_outputs(1468) <= a;
    layer5_outputs(1469) <= a and not b;
    layer5_outputs(1470) <= b;
    layer5_outputs(1471) <= a and b;
    layer5_outputs(1472) <= not (a and b);
    layer5_outputs(1473) <= '0';
    layer5_outputs(1474) <= not b;
    layer5_outputs(1475) <= not a;
    layer5_outputs(1476) <= not a;
    layer5_outputs(1477) <= not a;
    layer5_outputs(1478) <= not b;
    layer5_outputs(1479) <= not b;
    layer5_outputs(1480) <= a or b;
    layer5_outputs(1481) <= not (a or b);
    layer5_outputs(1482) <= not b;
    layer5_outputs(1483) <= '0';
    layer5_outputs(1484) <= b;
    layer5_outputs(1485) <= not (a and b);
    layer5_outputs(1486) <= not b;
    layer5_outputs(1487) <= a;
    layer5_outputs(1488) <= a and b;
    layer5_outputs(1489) <= not a or b;
    layer5_outputs(1490) <= a;
    layer5_outputs(1491) <= not (a and b);
    layer5_outputs(1492) <= '0';
    layer5_outputs(1493) <= a or b;
    layer5_outputs(1494) <= a and not b;
    layer5_outputs(1495) <= not (a or b);
    layer5_outputs(1496) <= not (a and b);
    layer5_outputs(1497) <= a or b;
    layer5_outputs(1498) <= not (a or b);
    layer5_outputs(1499) <= not (a or b);
    layer5_outputs(1500) <= not a;
    layer5_outputs(1501) <= a or b;
    layer5_outputs(1502) <= not b;
    layer5_outputs(1503) <= not b or a;
    layer5_outputs(1504) <= not a or b;
    layer5_outputs(1505) <= a and b;
    layer5_outputs(1506) <= not b or a;
    layer5_outputs(1507) <= not b;
    layer5_outputs(1508) <= not b;
    layer5_outputs(1509) <= a and not b;
    layer5_outputs(1510) <= not (a and b);
    layer5_outputs(1511) <= b;
    layer5_outputs(1512) <= b;
    layer5_outputs(1513) <= not b;
    layer5_outputs(1514) <= not a;
    layer5_outputs(1515) <= a;
    layer5_outputs(1516) <= not a;
    layer5_outputs(1517) <= a;
    layer5_outputs(1518) <= not (a or b);
    layer5_outputs(1519) <= a xor b;
    layer5_outputs(1520) <= a and b;
    layer5_outputs(1521) <= b;
    layer5_outputs(1522) <= a and b;
    layer5_outputs(1523) <= not a or b;
    layer5_outputs(1524) <= not (a and b);
    layer5_outputs(1525) <= '1';
    layer5_outputs(1526) <= not a;
    layer5_outputs(1527) <= not (a or b);
    layer5_outputs(1528) <= not a or b;
    layer5_outputs(1529) <= not b;
    layer5_outputs(1530) <= a and not b;
    layer5_outputs(1531) <= not b;
    layer5_outputs(1532) <= not a;
    layer5_outputs(1533) <= not a;
    layer5_outputs(1534) <= a and not b;
    layer5_outputs(1535) <= a;
    layer5_outputs(1536) <= not b or a;
    layer5_outputs(1537) <= not (a and b);
    layer5_outputs(1538) <= not (a and b);
    layer5_outputs(1539) <= a xor b;
    layer5_outputs(1540) <= not (a or b);
    layer5_outputs(1541) <= not b;
    layer5_outputs(1542) <= not b;
    layer5_outputs(1543) <= a and not b;
    layer5_outputs(1544) <= not a or b;
    layer5_outputs(1545) <= not a or b;
    layer5_outputs(1546) <= not (a and b);
    layer5_outputs(1547) <= b;
    layer5_outputs(1548) <= a and not b;
    layer5_outputs(1549) <= b;
    layer5_outputs(1550) <= a;
    layer5_outputs(1551) <= a;
    layer5_outputs(1552) <= a;
    layer5_outputs(1553) <= not (a and b);
    layer5_outputs(1554) <= not (a and b);
    layer5_outputs(1555) <= not a;
    layer5_outputs(1556) <= b;
    layer5_outputs(1557) <= not a;
    layer5_outputs(1558) <= b and not a;
    layer5_outputs(1559) <= a or b;
    layer5_outputs(1560) <= a;
    layer5_outputs(1561) <= '1';
    layer5_outputs(1562) <= not (a and b);
    layer5_outputs(1563) <= b;
    layer5_outputs(1564) <= not a;
    layer5_outputs(1565) <= a;
    layer5_outputs(1566) <= not a;
    layer5_outputs(1567) <= not (a or b);
    layer5_outputs(1568) <= not (a xor b);
    layer5_outputs(1569) <= a;
    layer5_outputs(1570) <= a and not b;
    layer5_outputs(1571) <= a or b;
    layer5_outputs(1572) <= a and b;
    layer5_outputs(1573) <= not b;
    layer5_outputs(1574) <= a;
    layer5_outputs(1575) <= not b;
    layer5_outputs(1576) <= not a or b;
    layer5_outputs(1577) <= a;
    layer5_outputs(1578) <= b;
    layer5_outputs(1579) <= b and not a;
    layer5_outputs(1580) <= a and b;
    layer5_outputs(1581) <= a xor b;
    layer5_outputs(1582) <= '0';
    layer5_outputs(1583) <= a;
    layer5_outputs(1584) <= a and not b;
    layer5_outputs(1585) <= b;
    layer5_outputs(1586) <= a;
    layer5_outputs(1587) <= '1';
    layer5_outputs(1588) <= '1';
    layer5_outputs(1589) <= b;
    layer5_outputs(1590) <= a and b;
    layer5_outputs(1591) <= not (a and b);
    layer5_outputs(1592) <= b;
    layer5_outputs(1593) <= not a;
    layer5_outputs(1594) <= b and not a;
    layer5_outputs(1595) <= b and not a;
    layer5_outputs(1596) <= not b;
    layer5_outputs(1597) <= not (a and b);
    layer5_outputs(1598) <= not a;
    layer5_outputs(1599) <= not (a and b);
    layer5_outputs(1600) <= a or b;
    layer5_outputs(1601) <= a and b;
    layer5_outputs(1602) <= b and not a;
    layer5_outputs(1603) <= a or b;
    layer5_outputs(1604) <= a and not b;
    layer5_outputs(1605) <= b and not a;
    layer5_outputs(1606) <= a xor b;
    layer5_outputs(1607) <= b;
    layer5_outputs(1608) <= b;
    layer5_outputs(1609) <= b and not a;
    layer5_outputs(1610) <= not (a xor b);
    layer5_outputs(1611) <= not b;
    layer5_outputs(1612) <= a;
    layer5_outputs(1613) <= not (a xor b);
    layer5_outputs(1614) <= a xor b;
    layer5_outputs(1615) <= a and b;
    layer5_outputs(1616) <= b;
    layer5_outputs(1617) <= not (a or b);
    layer5_outputs(1618) <= not a;
    layer5_outputs(1619) <= a xor b;
    layer5_outputs(1620) <= not b;
    layer5_outputs(1621) <= not a or b;
    layer5_outputs(1622) <= '0';
    layer5_outputs(1623) <= not b;
    layer5_outputs(1624) <= b;
    layer5_outputs(1625) <= '0';
    layer5_outputs(1626) <= a or b;
    layer5_outputs(1627) <= a;
    layer5_outputs(1628) <= not b or a;
    layer5_outputs(1629) <= not b;
    layer5_outputs(1630) <= b;
    layer5_outputs(1631) <= not b or a;
    layer5_outputs(1632) <= not a;
    layer5_outputs(1633) <= not b or a;
    layer5_outputs(1634) <= not a or b;
    layer5_outputs(1635) <= '1';
    layer5_outputs(1636) <= not b;
    layer5_outputs(1637) <= a and not b;
    layer5_outputs(1638) <= a;
    layer5_outputs(1639) <= not (a xor b);
    layer5_outputs(1640) <= a and not b;
    layer5_outputs(1641) <= '1';
    layer5_outputs(1642) <= not b or a;
    layer5_outputs(1643) <= a and not b;
    layer5_outputs(1644) <= not a or b;
    layer5_outputs(1645) <= a;
    layer5_outputs(1646) <= not a;
    layer5_outputs(1647) <= a xor b;
    layer5_outputs(1648) <= a and not b;
    layer5_outputs(1649) <= a or b;
    layer5_outputs(1650) <= b;
    layer5_outputs(1651) <= not a or b;
    layer5_outputs(1652) <= b;
    layer5_outputs(1653) <= not a;
    layer5_outputs(1654) <= not a or b;
    layer5_outputs(1655) <= a;
    layer5_outputs(1656) <= '1';
    layer5_outputs(1657) <= a and not b;
    layer5_outputs(1658) <= not b;
    layer5_outputs(1659) <= a and b;
    layer5_outputs(1660) <= a and b;
    layer5_outputs(1661) <= b;
    layer5_outputs(1662) <= a and b;
    layer5_outputs(1663) <= '0';
    layer5_outputs(1664) <= not b or a;
    layer5_outputs(1665) <= '0';
    layer5_outputs(1666) <= a and not b;
    layer5_outputs(1667) <= b;
    layer5_outputs(1668) <= not a;
    layer5_outputs(1669) <= not b or a;
    layer5_outputs(1670) <= not (a and b);
    layer5_outputs(1671) <= b;
    layer5_outputs(1672) <= not (a and b);
    layer5_outputs(1673) <= not a;
    layer5_outputs(1674) <= not b;
    layer5_outputs(1675) <= '0';
    layer5_outputs(1676) <= b;
    layer5_outputs(1677) <= '0';
    layer5_outputs(1678) <= not b or a;
    layer5_outputs(1679) <= '0';
    layer5_outputs(1680) <= not b or a;
    layer5_outputs(1681) <= not a;
    layer5_outputs(1682) <= b and not a;
    layer5_outputs(1683) <= not a;
    layer5_outputs(1684) <= not b;
    layer5_outputs(1685) <= b and not a;
    layer5_outputs(1686) <= b;
    layer5_outputs(1687) <= not (a and b);
    layer5_outputs(1688) <= a and b;
    layer5_outputs(1689) <= b;
    layer5_outputs(1690) <= not (a or b);
    layer5_outputs(1691) <= b;
    layer5_outputs(1692) <= b;
    layer5_outputs(1693) <= not (a and b);
    layer5_outputs(1694) <= not b;
    layer5_outputs(1695) <= '1';
    layer5_outputs(1696) <= '0';
    layer5_outputs(1697) <= not a;
    layer5_outputs(1698) <= '0';
    layer5_outputs(1699) <= not a or b;
    layer5_outputs(1700) <= a;
    layer5_outputs(1701) <= a xor b;
    layer5_outputs(1702) <= not b or a;
    layer5_outputs(1703) <= '0';
    layer5_outputs(1704) <= not a;
    layer5_outputs(1705) <= a and b;
    layer5_outputs(1706) <= not b;
    layer5_outputs(1707) <= '0';
    layer5_outputs(1708) <= b and not a;
    layer5_outputs(1709) <= b;
    layer5_outputs(1710) <= '1';
    layer5_outputs(1711) <= not (a xor b);
    layer5_outputs(1712) <= a and not b;
    layer5_outputs(1713) <= not (a or b);
    layer5_outputs(1714) <= not (a xor b);
    layer5_outputs(1715) <= b and not a;
    layer5_outputs(1716) <= not b;
    layer5_outputs(1717) <= b;
    layer5_outputs(1718) <= b;
    layer5_outputs(1719) <= '0';
    layer5_outputs(1720) <= not a;
    layer5_outputs(1721) <= not (a and b);
    layer5_outputs(1722) <= b;
    layer5_outputs(1723) <= a and b;
    layer5_outputs(1724) <= b;
    layer5_outputs(1725) <= not (a and b);
    layer5_outputs(1726) <= a or b;
    layer5_outputs(1727) <= not (a or b);
    layer5_outputs(1728) <= b;
    layer5_outputs(1729) <= not b;
    layer5_outputs(1730) <= not a or b;
    layer5_outputs(1731) <= not b or a;
    layer5_outputs(1732) <= b and not a;
    layer5_outputs(1733) <= '0';
    layer5_outputs(1734) <= not b;
    layer5_outputs(1735) <= '0';
    layer5_outputs(1736) <= b and not a;
    layer5_outputs(1737) <= b and not a;
    layer5_outputs(1738) <= a xor b;
    layer5_outputs(1739) <= not (a xor b);
    layer5_outputs(1740) <= a;
    layer5_outputs(1741) <= not b;
    layer5_outputs(1742) <= '0';
    layer5_outputs(1743) <= not b or a;
    layer5_outputs(1744) <= not a or b;
    layer5_outputs(1745) <= not a;
    layer5_outputs(1746) <= not a;
    layer5_outputs(1747) <= not (a or b);
    layer5_outputs(1748) <= not b or a;
    layer5_outputs(1749) <= a;
    layer5_outputs(1750) <= not (a and b);
    layer5_outputs(1751) <= not a;
    layer5_outputs(1752) <= b and not a;
    layer5_outputs(1753) <= not b;
    layer5_outputs(1754) <= a or b;
    layer5_outputs(1755) <= a xor b;
    layer5_outputs(1756) <= a;
    layer5_outputs(1757) <= b and not a;
    layer5_outputs(1758) <= not (a or b);
    layer5_outputs(1759) <= a and not b;
    layer5_outputs(1760) <= not a or b;
    layer5_outputs(1761) <= not a;
    layer5_outputs(1762) <= not b;
    layer5_outputs(1763) <= a;
    layer5_outputs(1764) <= b;
    layer5_outputs(1765) <= a and not b;
    layer5_outputs(1766) <= a and not b;
    layer5_outputs(1767) <= b and not a;
    layer5_outputs(1768) <= a;
    layer5_outputs(1769) <= not b;
    layer5_outputs(1770) <= not a;
    layer5_outputs(1771) <= not b;
    layer5_outputs(1772) <= not a;
    layer5_outputs(1773) <= a xor b;
    layer5_outputs(1774) <= not (a xor b);
    layer5_outputs(1775) <= '0';
    layer5_outputs(1776) <= not (a and b);
    layer5_outputs(1777) <= not a;
    layer5_outputs(1778) <= not b or a;
    layer5_outputs(1779) <= not (a and b);
    layer5_outputs(1780) <= not a;
    layer5_outputs(1781) <= a;
    layer5_outputs(1782) <= b and not a;
    layer5_outputs(1783) <= not a or b;
    layer5_outputs(1784) <= b;
    layer5_outputs(1785) <= not a or b;
    layer5_outputs(1786) <= not (a or b);
    layer5_outputs(1787) <= '0';
    layer5_outputs(1788) <= '1';
    layer5_outputs(1789) <= not b;
    layer5_outputs(1790) <= not (a and b);
    layer5_outputs(1791) <= a;
    layer5_outputs(1792) <= b;
    layer5_outputs(1793) <= not b or a;
    layer5_outputs(1794) <= a and b;
    layer5_outputs(1795) <= a and not b;
    layer5_outputs(1796) <= a;
    layer5_outputs(1797) <= a and not b;
    layer5_outputs(1798) <= not b;
    layer5_outputs(1799) <= not b;
    layer5_outputs(1800) <= not a or b;
    layer5_outputs(1801) <= a;
    layer5_outputs(1802) <= not a or b;
    layer5_outputs(1803) <= a;
    layer5_outputs(1804) <= not b;
    layer5_outputs(1805) <= b;
    layer5_outputs(1806) <= '0';
    layer5_outputs(1807) <= not b or a;
    layer5_outputs(1808) <= not (a or b);
    layer5_outputs(1809) <= not a;
    layer5_outputs(1810) <= a or b;
    layer5_outputs(1811) <= a or b;
    layer5_outputs(1812) <= b;
    layer5_outputs(1813) <= not (a xor b);
    layer5_outputs(1814) <= not b;
    layer5_outputs(1815) <= not (a or b);
    layer5_outputs(1816) <= not b or a;
    layer5_outputs(1817) <= a and b;
    layer5_outputs(1818) <= a xor b;
    layer5_outputs(1819) <= b;
    layer5_outputs(1820) <= a;
    layer5_outputs(1821) <= not b or a;
    layer5_outputs(1822) <= a xor b;
    layer5_outputs(1823) <= not (a xor b);
    layer5_outputs(1824) <= b;
    layer5_outputs(1825) <= a;
    layer5_outputs(1826) <= not a;
    layer5_outputs(1827) <= b;
    layer5_outputs(1828) <= a;
    layer5_outputs(1829) <= b and not a;
    layer5_outputs(1830) <= '0';
    layer5_outputs(1831) <= b;
    layer5_outputs(1832) <= a xor b;
    layer5_outputs(1833) <= a;
    layer5_outputs(1834) <= a and b;
    layer5_outputs(1835) <= not a;
    layer5_outputs(1836) <= a and not b;
    layer5_outputs(1837) <= '0';
    layer5_outputs(1838) <= a and not b;
    layer5_outputs(1839) <= a;
    layer5_outputs(1840) <= a or b;
    layer5_outputs(1841) <= b;
    layer5_outputs(1842) <= a xor b;
    layer5_outputs(1843) <= not (a and b);
    layer5_outputs(1844) <= not b;
    layer5_outputs(1845) <= b and not a;
    layer5_outputs(1846) <= not a or b;
    layer5_outputs(1847) <= b;
    layer5_outputs(1848) <= '0';
    layer5_outputs(1849) <= not a or b;
    layer5_outputs(1850) <= a and b;
    layer5_outputs(1851) <= a and not b;
    layer5_outputs(1852) <= not (a and b);
    layer5_outputs(1853) <= not b or a;
    layer5_outputs(1854) <= a and b;
    layer5_outputs(1855) <= b;
    layer5_outputs(1856) <= a xor b;
    layer5_outputs(1857) <= a and b;
    layer5_outputs(1858) <= a;
    layer5_outputs(1859) <= a and not b;
    layer5_outputs(1860) <= not a;
    layer5_outputs(1861) <= not (a or b);
    layer5_outputs(1862) <= not b;
    layer5_outputs(1863) <= b and not a;
    layer5_outputs(1864) <= a and not b;
    layer5_outputs(1865) <= not (a and b);
    layer5_outputs(1866) <= not (a or b);
    layer5_outputs(1867) <= not (a and b);
    layer5_outputs(1868) <= a and not b;
    layer5_outputs(1869) <= not a or b;
    layer5_outputs(1870) <= b;
    layer5_outputs(1871) <= b and not a;
    layer5_outputs(1872) <= not b;
    layer5_outputs(1873) <= a and not b;
    layer5_outputs(1874) <= not (a and b);
    layer5_outputs(1875) <= b and not a;
    layer5_outputs(1876) <= '1';
    layer5_outputs(1877) <= a and b;
    layer5_outputs(1878) <= not b or a;
    layer5_outputs(1879) <= b;
    layer5_outputs(1880) <= not (a or b);
    layer5_outputs(1881) <= b;
    layer5_outputs(1882) <= a and not b;
    layer5_outputs(1883) <= not b or a;
    layer5_outputs(1884) <= not a or b;
    layer5_outputs(1885) <= not a or b;
    layer5_outputs(1886) <= b;
    layer5_outputs(1887) <= b;
    layer5_outputs(1888) <= a and not b;
    layer5_outputs(1889) <= a xor b;
    layer5_outputs(1890) <= b;
    layer5_outputs(1891) <= not b or a;
    layer5_outputs(1892) <= b;
    layer5_outputs(1893) <= not a;
    layer5_outputs(1894) <= not b or a;
    layer5_outputs(1895) <= not (a xor b);
    layer5_outputs(1896) <= not (a or b);
    layer5_outputs(1897) <= not b;
    layer5_outputs(1898) <= not a;
    layer5_outputs(1899) <= not a or b;
    layer5_outputs(1900) <= not b;
    layer5_outputs(1901) <= a or b;
    layer5_outputs(1902) <= '0';
    layer5_outputs(1903) <= not a;
    layer5_outputs(1904) <= b;
    layer5_outputs(1905) <= a and b;
    layer5_outputs(1906) <= b and not a;
    layer5_outputs(1907) <= not b or a;
    layer5_outputs(1908) <= not (a or b);
    layer5_outputs(1909) <= a and b;
    layer5_outputs(1910) <= not b or a;
    layer5_outputs(1911) <= not b;
    layer5_outputs(1912) <= a and not b;
    layer5_outputs(1913) <= b and not a;
    layer5_outputs(1914) <= b;
    layer5_outputs(1915) <= a and not b;
    layer5_outputs(1916) <= a and not b;
    layer5_outputs(1917) <= a;
    layer5_outputs(1918) <= a and b;
    layer5_outputs(1919) <= a;
    layer5_outputs(1920) <= not b;
    layer5_outputs(1921) <= not a;
    layer5_outputs(1922) <= not a or b;
    layer5_outputs(1923) <= a;
    layer5_outputs(1924) <= not a;
    layer5_outputs(1925) <= not a or b;
    layer5_outputs(1926) <= not a;
    layer5_outputs(1927) <= a and not b;
    layer5_outputs(1928) <= not b or a;
    layer5_outputs(1929) <= a and b;
    layer5_outputs(1930) <= not (a or b);
    layer5_outputs(1931) <= not a;
    layer5_outputs(1932) <= b and not a;
    layer5_outputs(1933) <= not a;
    layer5_outputs(1934) <= not (a or b);
    layer5_outputs(1935) <= a and not b;
    layer5_outputs(1936) <= not (a or b);
    layer5_outputs(1937) <= not (a and b);
    layer5_outputs(1938) <= a and b;
    layer5_outputs(1939) <= not b or a;
    layer5_outputs(1940) <= b and not a;
    layer5_outputs(1941) <= not (a and b);
    layer5_outputs(1942) <= a and not b;
    layer5_outputs(1943) <= not b;
    layer5_outputs(1944) <= not a or b;
    layer5_outputs(1945) <= '1';
    layer5_outputs(1946) <= b and not a;
    layer5_outputs(1947) <= not (a and b);
    layer5_outputs(1948) <= b;
    layer5_outputs(1949) <= not (a xor b);
    layer5_outputs(1950) <= '1';
    layer5_outputs(1951) <= a and b;
    layer5_outputs(1952) <= a and b;
    layer5_outputs(1953) <= a or b;
    layer5_outputs(1954) <= '1';
    layer5_outputs(1955) <= a and b;
    layer5_outputs(1956) <= not a;
    layer5_outputs(1957) <= b;
    layer5_outputs(1958) <= not a;
    layer5_outputs(1959) <= not (a or b);
    layer5_outputs(1960) <= a and not b;
    layer5_outputs(1961) <= not b;
    layer5_outputs(1962) <= not (a xor b);
    layer5_outputs(1963) <= b and not a;
    layer5_outputs(1964) <= b;
    layer5_outputs(1965) <= not a or b;
    layer5_outputs(1966) <= b and not a;
    layer5_outputs(1967) <= not a;
    layer5_outputs(1968) <= not a;
    layer5_outputs(1969) <= a or b;
    layer5_outputs(1970) <= not a;
    layer5_outputs(1971) <= b;
    layer5_outputs(1972) <= not b or a;
    layer5_outputs(1973) <= a or b;
    layer5_outputs(1974) <= b;
    layer5_outputs(1975) <= a;
    layer5_outputs(1976) <= a and b;
    layer5_outputs(1977) <= a or b;
    layer5_outputs(1978) <= not b;
    layer5_outputs(1979) <= '0';
    layer5_outputs(1980) <= a;
    layer5_outputs(1981) <= a xor b;
    layer5_outputs(1982) <= not b;
    layer5_outputs(1983) <= not a;
    layer5_outputs(1984) <= a and b;
    layer5_outputs(1985) <= not b or a;
    layer5_outputs(1986) <= not b or a;
    layer5_outputs(1987) <= a and b;
    layer5_outputs(1988) <= not (a and b);
    layer5_outputs(1989) <= not b or a;
    layer5_outputs(1990) <= a;
    layer5_outputs(1991) <= b;
    layer5_outputs(1992) <= '1';
    layer5_outputs(1993) <= a and b;
    layer5_outputs(1994) <= not (a or b);
    layer5_outputs(1995) <= not b or a;
    layer5_outputs(1996) <= not b;
    layer5_outputs(1997) <= not a or b;
    layer5_outputs(1998) <= '1';
    layer5_outputs(1999) <= b and not a;
    layer5_outputs(2000) <= a or b;
    layer5_outputs(2001) <= b;
    layer5_outputs(2002) <= a and b;
    layer5_outputs(2003) <= not b;
    layer5_outputs(2004) <= a xor b;
    layer5_outputs(2005) <= not b or a;
    layer5_outputs(2006) <= not (a xor b);
    layer5_outputs(2007) <= a;
    layer5_outputs(2008) <= not (a and b);
    layer5_outputs(2009) <= a and not b;
    layer5_outputs(2010) <= not a;
    layer5_outputs(2011) <= a;
    layer5_outputs(2012) <= a xor b;
    layer5_outputs(2013) <= '1';
    layer5_outputs(2014) <= a and b;
    layer5_outputs(2015) <= b and not a;
    layer5_outputs(2016) <= not a;
    layer5_outputs(2017) <= a xor b;
    layer5_outputs(2018) <= not (a and b);
    layer5_outputs(2019) <= '1';
    layer5_outputs(2020) <= b;
    layer5_outputs(2021) <= not (a and b);
    layer5_outputs(2022) <= not a or b;
    layer5_outputs(2023) <= not a;
    layer5_outputs(2024) <= b;
    layer5_outputs(2025) <= a xor b;
    layer5_outputs(2026) <= not a or b;
    layer5_outputs(2027) <= a;
    layer5_outputs(2028) <= b;
    layer5_outputs(2029) <= b and not a;
    layer5_outputs(2030) <= a;
    layer5_outputs(2031) <= b;
    layer5_outputs(2032) <= a or b;
    layer5_outputs(2033) <= a xor b;
    layer5_outputs(2034) <= a;
    layer5_outputs(2035) <= not b;
    layer5_outputs(2036) <= not (a and b);
    layer5_outputs(2037) <= a;
    layer5_outputs(2038) <= '1';
    layer5_outputs(2039) <= a and b;
    layer5_outputs(2040) <= not (a xor b);
    layer5_outputs(2041) <= not b or a;
    layer5_outputs(2042) <= a or b;
    layer5_outputs(2043) <= not (a and b);
    layer5_outputs(2044) <= not b;
    layer5_outputs(2045) <= not a or b;
    layer5_outputs(2046) <= not a or b;
    layer5_outputs(2047) <= a and not b;
    layer5_outputs(2048) <= not b;
    layer5_outputs(2049) <= not (a xor b);
    layer5_outputs(2050) <= not (a or b);
    layer5_outputs(2051) <= b;
    layer5_outputs(2052) <= not (a and b);
    layer5_outputs(2053) <= not a;
    layer5_outputs(2054) <= a xor b;
    layer5_outputs(2055) <= not a;
    layer5_outputs(2056) <= '0';
    layer5_outputs(2057) <= a xor b;
    layer5_outputs(2058) <= not a or b;
    layer5_outputs(2059) <= a and b;
    layer5_outputs(2060) <= b and not a;
    layer5_outputs(2061) <= a and not b;
    layer5_outputs(2062) <= b;
    layer5_outputs(2063) <= a;
    layer5_outputs(2064) <= not b;
    layer5_outputs(2065) <= b;
    layer5_outputs(2066) <= a and not b;
    layer5_outputs(2067) <= a and not b;
    layer5_outputs(2068) <= not a or b;
    layer5_outputs(2069) <= not b;
    layer5_outputs(2070) <= a or b;
    layer5_outputs(2071) <= b;
    layer5_outputs(2072) <= not a;
    layer5_outputs(2073) <= a;
    layer5_outputs(2074) <= not a;
    layer5_outputs(2075) <= a;
    layer5_outputs(2076) <= not a;
    layer5_outputs(2077) <= a;
    layer5_outputs(2078) <= not (a and b);
    layer5_outputs(2079) <= a;
    layer5_outputs(2080) <= b;
    layer5_outputs(2081) <= b;
    layer5_outputs(2082) <= not a or b;
    layer5_outputs(2083) <= '0';
    layer5_outputs(2084) <= a and not b;
    layer5_outputs(2085) <= a or b;
    layer5_outputs(2086) <= not b or a;
    layer5_outputs(2087) <= not b or a;
    layer5_outputs(2088) <= not (a or b);
    layer5_outputs(2089) <= not (a or b);
    layer5_outputs(2090) <= not b;
    layer5_outputs(2091) <= not b;
    layer5_outputs(2092) <= a or b;
    layer5_outputs(2093) <= not b or a;
    layer5_outputs(2094) <= a;
    layer5_outputs(2095) <= not b;
    layer5_outputs(2096) <= not b;
    layer5_outputs(2097) <= a and not b;
    layer5_outputs(2098) <= b;
    layer5_outputs(2099) <= b;
    layer5_outputs(2100) <= b and not a;
    layer5_outputs(2101) <= a;
    layer5_outputs(2102) <= '1';
    layer5_outputs(2103) <= not b;
    layer5_outputs(2104) <= '1';
    layer5_outputs(2105) <= not (a and b);
    layer5_outputs(2106) <= a and b;
    layer5_outputs(2107) <= not b;
    layer5_outputs(2108) <= a or b;
    layer5_outputs(2109) <= not a or b;
    layer5_outputs(2110) <= a or b;
    layer5_outputs(2111) <= not a;
    layer5_outputs(2112) <= not b or a;
    layer5_outputs(2113) <= not a;
    layer5_outputs(2114) <= a and b;
    layer5_outputs(2115) <= b;
    layer5_outputs(2116) <= a;
    layer5_outputs(2117) <= a;
    layer5_outputs(2118) <= a or b;
    layer5_outputs(2119) <= not b;
    layer5_outputs(2120) <= not (a or b);
    layer5_outputs(2121) <= not (a or b);
    layer5_outputs(2122) <= b and not a;
    layer5_outputs(2123) <= a;
    layer5_outputs(2124) <= not b;
    layer5_outputs(2125) <= a and b;
    layer5_outputs(2126) <= not a or b;
    layer5_outputs(2127) <= b and not a;
    layer5_outputs(2128) <= a and not b;
    layer5_outputs(2129) <= not a;
    layer5_outputs(2130) <= a or b;
    layer5_outputs(2131) <= a;
    layer5_outputs(2132) <= a or b;
    layer5_outputs(2133) <= '1';
    layer5_outputs(2134) <= b and not a;
    layer5_outputs(2135) <= not b or a;
    layer5_outputs(2136) <= not a;
    layer5_outputs(2137) <= not b;
    layer5_outputs(2138) <= a or b;
    layer5_outputs(2139) <= not b;
    layer5_outputs(2140) <= not a;
    layer5_outputs(2141) <= '1';
    layer5_outputs(2142) <= a and b;
    layer5_outputs(2143) <= not a;
    layer5_outputs(2144) <= '0';
    layer5_outputs(2145) <= a and b;
    layer5_outputs(2146) <= a or b;
    layer5_outputs(2147) <= not b;
    layer5_outputs(2148) <= b;
    layer5_outputs(2149) <= not a or b;
    layer5_outputs(2150) <= not a or b;
    layer5_outputs(2151) <= not (a xor b);
    layer5_outputs(2152) <= not a or b;
    layer5_outputs(2153) <= not a or b;
    layer5_outputs(2154) <= b and not a;
    layer5_outputs(2155) <= b and not a;
    layer5_outputs(2156) <= '1';
    layer5_outputs(2157) <= not a or b;
    layer5_outputs(2158) <= not (a or b);
    layer5_outputs(2159) <= a and not b;
    layer5_outputs(2160) <= not (a or b);
    layer5_outputs(2161) <= '1';
    layer5_outputs(2162) <= b;
    layer5_outputs(2163) <= a and not b;
    layer5_outputs(2164) <= a xor b;
    layer5_outputs(2165) <= not b or a;
    layer5_outputs(2166) <= not (a and b);
    layer5_outputs(2167) <= b and not a;
    layer5_outputs(2168) <= b;
    layer5_outputs(2169) <= not a;
    layer5_outputs(2170) <= not a or b;
    layer5_outputs(2171) <= b;
    layer5_outputs(2172) <= not a or b;
    layer5_outputs(2173) <= '0';
    layer5_outputs(2174) <= not b;
    layer5_outputs(2175) <= a and b;
    layer5_outputs(2176) <= b and not a;
    layer5_outputs(2177) <= a and b;
    layer5_outputs(2178) <= b;
    layer5_outputs(2179) <= not b;
    layer5_outputs(2180) <= not a or b;
    layer5_outputs(2181) <= not a or b;
    layer5_outputs(2182) <= a;
    layer5_outputs(2183) <= a and b;
    layer5_outputs(2184) <= a and b;
    layer5_outputs(2185) <= a;
    layer5_outputs(2186) <= not (a xor b);
    layer5_outputs(2187) <= a xor b;
    layer5_outputs(2188) <= b;
    layer5_outputs(2189) <= not a;
    layer5_outputs(2190) <= not a;
    layer5_outputs(2191) <= a or b;
    layer5_outputs(2192) <= not a;
    layer5_outputs(2193) <= b;
    layer5_outputs(2194) <= b;
    layer5_outputs(2195) <= a and b;
    layer5_outputs(2196) <= b;
    layer5_outputs(2197) <= '1';
    layer5_outputs(2198) <= a;
    layer5_outputs(2199) <= '1';
    layer5_outputs(2200) <= a and not b;
    layer5_outputs(2201) <= not (a or b);
    layer5_outputs(2202) <= b;
    layer5_outputs(2203) <= a;
    layer5_outputs(2204) <= not a;
    layer5_outputs(2205) <= not (a or b);
    layer5_outputs(2206) <= a and not b;
    layer5_outputs(2207) <= b;
    layer5_outputs(2208) <= '0';
    layer5_outputs(2209) <= not b or a;
    layer5_outputs(2210) <= not a;
    layer5_outputs(2211) <= a and not b;
    layer5_outputs(2212) <= not a;
    layer5_outputs(2213) <= not a;
    layer5_outputs(2214) <= b and not a;
    layer5_outputs(2215) <= b;
    layer5_outputs(2216) <= b and not a;
    layer5_outputs(2217) <= not b or a;
    layer5_outputs(2218) <= b and not a;
    layer5_outputs(2219) <= a;
    layer5_outputs(2220) <= not b;
    layer5_outputs(2221) <= a xor b;
    layer5_outputs(2222) <= a or b;
    layer5_outputs(2223) <= not (a and b);
    layer5_outputs(2224) <= not a;
    layer5_outputs(2225) <= not b or a;
    layer5_outputs(2226) <= a or b;
    layer5_outputs(2227) <= b;
    layer5_outputs(2228) <= a or b;
    layer5_outputs(2229) <= '1';
    layer5_outputs(2230) <= not a or b;
    layer5_outputs(2231) <= not b;
    layer5_outputs(2232) <= not a;
    layer5_outputs(2233) <= not a;
    layer5_outputs(2234) <= not (a or b);
    layer5_outputs(2235) <= a xor b;
    layer5_outputs(2236) <= a;
    layer5_outputs(2237) <= a and b;
    layer5_outputs(2238) <= b;
    layer5_outputs(2239) <= not (a or b);
    layer5_outputs(2240) <= b and not a;
    layer5_outputs(2241) <= not (a or b);
    layer5_outputs(2242) <= not a;
    layer5_outputs(2243) <= not b or a;
    layer5_outputs(2244) <= a and not b;
    layer5_outputs(2245) <= not a;
    layer5_outputs(2246) <= not (a and b);
    layer5_outputs(2247) <= '0';
    layer5_outputs(2248) <= not (a or b);
    layer5_outputs(2249) <= a and not b;
    layer5_outputs(2250) <= not a;
    layer5_outputs(2251) <= not a or b;
    layer5_outputs(2252) <= not b;
    layer5_outputs(2253) <= not a or b;
    layer5_outputs(2254) <= not b;
    layer5_outputs(2255) <= b and not a;
    layer5_outputs(2256) <= b and not a;
    layer5_outputs(2257) <= a;
    layer5_outputs(2258) <= b and not a;
    layer5_outputs(2259) <= not b;
    layer5_outputs(2260) <= a;
    layer5_outputs(2261) <= '1';
    layer5_outputs(2262) <= not b or a;
    layer5_outputs(2263) <= not b;
    layer5_outputs(2264) <= not a or b;
    layer5_outputs(2265) <= b;
    layer5_outputs(2266) <= '0';
    layer5_outputs(2267) <= not b;
    layer5_outputs(2268) <= a xor b;
    layer5_outputs(2269) <= not a;
    layer5_outputs(2270) <= not a or b;
    layer5_outputs(2271) <= not b;
    layer5_outputs(2272) <= not b;
    layer5_outputs(2273) <= not a;
    layer5_outputs(2274) <= not b or a;
    layer5_outputs(2275) <= a;
    layer5_outputs(2276) <= b;
    layer5_outputs(2277) <= b;
    layer5_outputs(2278) <= not b;
    layer5_outputs(2279) <= not b;
    layer5_outputs(2280) <= not a;
    layer5_outputs(2281) <= a and b;
    layer5_outputs(2282) <= a and b;
    layer5_outputs(2283) <= '0';
    layer5_outputs(2284) <= not (a and b);
    layer5_outputs(2285) <= b and not a;
    layer5_outputs(2286) <= not b or a;
    layer5_outputs(2287) <= '1';
    layer5_outputs(2288) <= not a;
    layer5_outputs(2289) <= not b;
    layer5_outputs(2290) <= not (a xor b);
    layer5_outputs(2291) <= a or b;
    layer5_outputs(2292) <= b and not a;
    layer5_outputs(2293) <= b;
    layer5_outputs(2294) <= a;
    layer5_outputs(2295) <= not a;
    layer5_outputs(2296) <= b and not a;
    layer5_outputs(2297) <= b and not a;
    layer5_outputs(2298) <= b;
    layer5_outputs(2299) <= not (a and b);
    layer5_outputs(2300) <= not b or a;
    layer5_outputs(2301) <= not (a or b);
    layer5_outputs(2302) <= a;
    layer5_outputs(2303) <= a;
    layer5_outputs(2304) <= not a;
    layer5_outputs(2305) <= a;
    layer5_outputs(2306) <= b and not a;
    layer5_outputs(2307) <= not (a and b);
    layer5_outputs(2308) <= not a or b;
    layer5_outputs(2309) <= a;
    layer5_outputs(2310) <= a and not b;
    layer5_outputs(2311) <= not (a or b);
    layer5_outputs(2312) <= not (a xor b);
    layer5_outputs(2313) <= b;
    layer5_outputs(2314) <= b and not a;
    layer5_outputs(2315) <= not (a or b);
    layer5_outputs(2316) <= not a;
    layer5_outputs(2317) <= b and not a;
    layer5_outputs(2318) <= a or b;
    layer5_outputs(2319) <= not a;
    layer5_outputs(2320) <= a;
    layer5_outputs(2321) <= not b or a;
    layer5_outputs(2322) <= b;
    layer5_outputs(2323) <= not a or b;
    layer5_outputs(2324) <= b;
    layer5_outputs(2325) <= not a or b;
    layer5_outputs(2326) <= not a;
    layer5_outputs(2327) <= '1';
    layer5_outputs(2328) <= a and not b;
    layer5_outputs(2329) <= a xor b;
    layer5_outputs(2330) <= not a or b;
    layer5_outputs(2331) <= not b;
    layer5_outputs(2332) <= not a;
    layer5_outputs(2333) <= '1';
    layer5_outputs(2334) <= not b;
    layer5_outputs(2335) <= not b;
    layer5_outputs(2336) <= not b;
    layer5_outputs(2337) <= not b;
    layer5_outputs(2338) <= not a;
    layer5_outputs(2339) <= not b or a;
    layer5_outputs(2340) <= a or b;
    layer5_outputs(2341) <= a;
    layer5_outputs(2342) <= not b;
    layer5_outputs(2343) <= a xor b;
    layer5_outputs(2344) <= a and not b;
    layer5_outputs(2345) <= not b;
    layer5_outputs(2346) <= a xor b;
    layer5_outputs(2347) <= not (a or b);
    layer5_outputs(2348) <= a and not b;
    layer5_outputs(2349) <= b;
    layer5_outputs(2350) <= not (a and b);
    layer5_outputs(2351) <= b;
    layer5_outputs(2352) <= not b;
    layer5_outputs(2353) <= not b;
    layer5_outputs(2354) <= a and not b;
    layer5_outputs(2355) <= not b or a;
    layer5_outputs(2356) <= a;
    layer5_outputs(2357) <= a and not b;
    layer5_outputs(2358) <= a and not b;
    layer5_outputs(2359) <= not a or b;
    layer5_outputs(2360) <= '0';
    layer5_outputs(2361) <= not b or a;
    layer5_outputs(2362) <= '1';
    layer5_outputs(2363) <= not a;
    layer5_outputs(2364) <= not (a and b);
    layer5_outputs(2365) <= '0';
    layer5_outputs(2366) <= not b or a;
    layer5_outputs(2367) <= b and not a;
    layer5_outputs(2368) <= a;
    layer5_outputs(2369) <= not b;
    layer5_outputs(2370) <= not b or a;
    layer5_outputs(2371) <= not (a or b);
    layer5_outputs(2372) <= not (a and b);
    layer5_outputs(2373) <= a or b;
    layer5_outputs(2374) <= a;
    layer5_outputs(2375) <= b and not a;
    layer5_outputs(2376) <= a;
    layer5_outputs(2377) <= not a;
    layer5_outputs(2378) <= a or b;
    layer5_outputs(2379) <= b;
    layer5_outputs(2380) <= a;
    layer5_outputs(2381) <= b and not a;
    layer5_outputs(2382) <= not a;
    layer5_outputs(2383) <= b and not a;
    layer5_outputs(2384) <= a;
    layer5_outputs(2385) <= not (a xor b);
    layer5_outputs(2386) <= not b or a;
    layer5_outputs(2387) <= not a;
    layer5_outputs(2388) <= not a or b;
    layer5_outputs(2389) <= not (a xor b);
    layer5_outputs(2390) <= a;
    layer5_outputs(2391) <= a;
    layer5_outputs(2392) <= a and not b;
    layer5_outputs(2393) <= not (a and b);
    layer5_outputs(2394) <= a and not b;
    layer5_outputs(2395) <= b;
    layer5_outputs(2396) <= not b or a;
    layer5_outputs(2397) <= a and b;
    layer5_outputs(2398) <= a and b;
    layer5_outputs(2399) <= b and not a;
    layer5_outputs(2400) <= not b;
    layer5_outputs(2401) <= not (a or b);
    layer5_outputs(2402) <= not (a xor b);
    layer5_outputs(2403) <= not b;
    layer5_outputs(2404) <= '0';
    layer5_outputs(2405) <= not b or a;
    layer5_outputs(2406) <= a;
    layer5_outputs(2407) <= not b;
    layer5_outputs(2408) <= b;
    layer5_outputs(2409) <= not b;
    layer5_outputs(2410) <= b;
    layer5_outputs(2411) <= not a;
    layer5_outputs(2412) <= not b or a;
    layer5_outputs(2413) <= not (a or b);
    layer5_outputs(2414) <= not b or a;
    layer5_outputs(2415) <= a;
    layer5_outputs(2416) <= not (a and b);
    layer5_outputs(2417) <= b and not a;
    layer5_outputs(2418) <= not b or a;
    layer5_outputs(2419) <= not a or b;
    layer5_outputs(2420) <= a and not b;
    layer5_outputs(2421) <= a and not b;
    layer5_outputs(2422) <= b;
    layer5_outputs(2423) <= not a or b;
    layer5_outputs(2424) <= not b or a;
    layer5_outputs(2425) <= '1';
    layer5_outputs(2426) <= not b;
    layer5_outputs(2427) <= b and not a;
    layer5_outputs(2428) <= a;
    layer5_outputs(2429) <= not b or a;
    layer5_outputs(2430) <= not (a xor b);
    layer5_outputs(2431) <= not (a and b);
    layer5_outputs(2432) <= a and b;
    layer5_outputs(2433) <= not b;
    layer5_outputs(2434) <= a and b;
    layer5_outputs(2435) <= a or b;
    layer5_outputs(2436) <= b and not a;
    layer5_outputs(2437) <= not a;
    layer5_outputs(2438) <= not a;
    layer5_outputs(2439) <= a and not b;
    layer5_outputs(2440) <= not b or a;
    layer5_outputs(2441) <= not a;
    layer5_outputs(2442) <= not b or a;
    layer5_outputs(2443) <= b;
    layer5_outputs(2444) <= not a;
    layer5_outputs(2445) <= not b or a;
    layer5_outputs(2446) <= b;
    layer5_outputs(2447) <= a;
    layer5_outputs(2448) <= a xor b;
    layer5_outputs(2449) <= b and not a;
    layer5_outputs(2450) <= a and not b;
    layer5_outputs(2451) <= a or b;
    layer5_outputs(2452) <= not b or a;
    layer5_outputs(2453) <= not b or a;
    layer5_outputs(2454) <= not (a and b);
    layer5_outputs(2455) <= not b;
    layer5_outputs(2456) <= not (a xor b);
    layer5_outputs(2457) <= not a;
    layer5_outputs(2458) <= b and not a;
    layer5_outputs(2459) <= not a;
    layer5_outputs(2460) <= b and not a;
    layer5_outputs(2461) <= not b;
    layer5_outputs(2462) <= b;
    layer5_outputs(2463) <= not a;
    layer5_outputs(2464) <= not a or b;
    layer5_outputs(2465) <= '0';
    layer5_outputs(2466) <= not b;
    layer5_outputs(2467) <= a;
    layer5_outputs(2468) <= a xor b;
    layer5_outputs(2469) <= a;
    layer5_outputs(2470) <= b;
    layer5_outputs(2471) <= not b;
    layer5_outputs(2472) <= a and not b;
    layer5_outputs(2473) <= a xor b;
    layer5_outputs(2474) <= not (a and b);
    layer5_outputs(2475) <= not a or b;
    layer5_outputs(2476) <= not a or b;
    layer5_outputs(2477) <= b and not a;
    layer5_outputs(2478) <= not b;
    layer5_outputs(2479) <= a or b;
    layer5_outputs(2480) <= not b;
    layer5_outputs(2481) <= a and not b;
    layer5_outputs(2482) <= a;
    layer5_outputs(2483) <= b;
    layer5_outputs(2484) <= not b or a;
    layer5_outputs(2485) <= a or b;
    layer5_outputs(2486) <= not a;
    layer5_outputs(2487) <= b and not a;
    layer5_outputs(2488) <= not a;
    layer5_outputs(2489) <= '0';
    layer5_outputs(2490) <= not (a xor b);
    layer5_outputs(2491) <= a and not b;
    layer5_outputs(2492) <= a and b;
    layer5_outputs(2493) <= not a or b;
    layer5_outputs(2494) <= b;
    layer5_outputs(2495) <= not b;
    layer5_outputs(2496) <= '0';
    layer5_outputs(2497) <= a;
    layer5_outputs(2498) <= a and not b;
    layer5_outputs(2499) <= '1';
    layer5_outputs(2500) <= a;
    layer5_outputs(2501) <= not (a and b);
    layer5_outputs(2502) <= a and not b;
    layer5_outputs(2503) <= a and b;
    layer5_outputs(2504) <= b;
    layer5_outputs(2505) <= a;
    layer5_outputs(2506) <= '1';
    layer5_outputs(2507) <= a or b;
    layer5_outputs(2508) <= not b or a;
    layer5_outputs(2509) <= a;
    layer5_outputs(2510) <= '0';
    layer5_outputs(2511) <= not a;
    layer5_outputs(2512) <= not a;
    layer5_outputs(2513) <= a xor b;
    layer5_outputs(2514) <= not b;
    layer5_outputs(2515) <= a and not b;
    layer5_outputs(2516) <= not b;
    layer5_outputs(2517) <= a and not b;
    layer5_outputs(2518) <= b;
    layer5_outputs(2519) <= '1';
    layer5_outputs(2520) <= not (a and b);
    layer5_outputs(2521) <= a;
    layer5_outputs(2522) <= not b or a;
    layer5_outputs(2523) <= b and not a;
    layer5_outputs(2524) <= not b;
    layer5_outputs(2525) <= a or b;
    layer5_outputs(2526) <= a and b;
    layer5_outputs(2527) <= not b or a;
    layer5_outputs(2528) <= not a;
    layer5_outputs(2529) <= a and b;
    layer5_outputs(2530) <= not a;
    layer5_outputs(2531) <= a xor b;
    layer5_outputs(2532) <= not a or b;
    layer5_outputs(2533) <= not b or a;
    layer5_outputs(2534) <= a;
    layer5_outputs(2535) <= a;
    layer5_outputs(2536) <= a and b;
    layer5_outputs(2537) <= not a;
    layer5_outputs(2538) <= b and not a;
    layer5_outputs(2539) <= a and not b;
    layer5_outputs(2540) <= a;
    layer5_outputs(2541) <= b;
    layer5_outputs(2542) <= b;
    layer5_outputs(2543) <= not b;
    layer5_outputs(2544) <= '1';
    layer5_outputs(2545) <= a;
    layer5_outputs(2546) <= a;
    layer5_outputs(2547) <= b;
    layer5_outputs(2548) <= not b;
    layer5_outputs(2549) <= b and not a;
    layer5_outputs(2550) <= '0';
    layer5_outputs(2551) <= not a;
    layer5_outputs(2552) <= a and not b;
    layer5_outputs(2553) <= b and not a;
    layer5_outputs(2554) <= '0';
    layer5_outputs(2555) <= a and not b;
    layer5_outputs(2556) <= not a;
    layer5_outputs(2557) <= not a;
    layer5_outputs(2558) <= a;
    layer5_outputs(2559) <= '0';
    layer5_outputs(2560) <= a and b;
    layer5_outputs(2561) <= a and b;
    layer5_outputs(2562) <= b;
    layer5_outputs(2563) <= '0';
    layer5_outputs(2564) <= b and not a;
    layer5_outputs(2565) <= not b;
    layer5_outputs(2566) <= b;
    layer5_outputs(2567) <= not (a xor b);
    layer5_outputs(2568) <= b;
    layer5_outputs(2569) <= not a;
    layer5_outputs(2570) <= not a;
    layer5_outputs(2571) <= not (a xor b);
    layer5_outputs(2572) <= a and not b;
    layer5_outputs(2573) <= not (a or b);
    layer5_outputs(2574) <= not a;
    layer5_outputs(2575) <= '1';
    layer5_outputs(2576) <= '1';
    layer5_outputs(2577) <= not b;
    layer5_outputs(2578) <= b;
    layer5_outputs(2579) <= a;
    layer5_outputs(2580) <= a;
    layer5_outputs(2581) <= a and b;
    layer5_outputs(2582) <= b and not a;
    layer5_outputs(2583) <= b;
    layer5_outputs(2584) <= b and not a;
    layer5_outputs(2585) <= not b;
    layer5_outputs(2586) <= not b;
    layer5_outputs(2587) <= not (a or b);
    layer5_outputs(2588) <= b and not a;
    layer5_outputs(2589) <= a and not b;
    layer5_outputs(2590) <= not (a xor b);
    layer5_outputs(2591) <= not a;
    layer5_outputs(2592) <= not a;
    layer5_outputs(2593) <= b and not a;
    layer5_outputs(2594) <= not a;
    layer5_outputs(2595) <= not (a or b);
    layer5_outputs(2596) <= not a;
    layer5_outputs(2597) <= not b;
    layer5_outputs(2598) <= not (a xor b);
    layer5_outputs(2599) <= b and not a;
    layer5_outputs(2600) <= b;
    layer5_outputs(2601) <= not b or a;
    layer5_outputs(2602) <= b;
    layer5_outputs(2603) <= a;
    layer5_outputs(2604) <= a or b;
    layer5_outputs(2605) <= a xor b;
    layer5_outputs(2606) <= a or b;
    layer5_outputs(2607) <= b;
    layer5_outputs(2608) <= a xor b;
    layer5_outputs(2609) <= b;
    layer5_outputs(2610) <= not a or b;
    layer5_outputs(2611) <= not (a or b);
    layer5_outputs(2612) <= a;
    layer5_outputs(2613) <= not (a xor b);
    layer5_outputs(2614) <= a;
    layer5_outputs(2615) <= not a;
    layer5_outputs(2616) <= a or b;
    layer5_outputs(2617) <= '1';
    layer5_outputs(2618) <= not (a or b);
    layer5_outputs(2619) <= '0';
    layer5_outputs(2620) <= not (a and b);
    layer5_outputs(2621) <= not a;
    layer5_outputs(2622) <= not b or a;
    layer5_outputs(2623) <= b and not a;
    layer5_outputs(2624) <= not (a xor b);
    layer5_outputs(2625) <= not (a or b);
    layer5_outputs(2626) <= b and not a;
    layer5_outputs(2627) <= not b or a;
    layer5_outputs(2628) <= a xor b;
    layer5_outputs(2629) <= not a;
    layer5_outputs(2630) <= a or b;
    layer5_outputs(2631) <= a;
    layer5_outputs(2632) <= not a;
    layer5_outputs(2633) <= not (a and b);
    layer5_outputs(2634) <= '1';
    layer5_outputs(2635) <= b and not a;
    layer5_outputs(2636) <= not (a and b);
    layer5_outputs(2637) <= not (a and b);
    layer5_outputs(2638) <= a xor b;
    layer5_outputs(2639) <= '0';
    layer5_outputs(2640) <= not b;
    layer5_outputs(2641) <= not (a or b);
    layer5_outputs(2642) <= a or b;
    layer5_outputs(2643) <= '1';
    layer5_outputs(2644) <= a;
    layer5_outputs(2645) <= not (a and b);
    layer5_outputs(2646) <= not (a and b);
    layer5_outputs(2647) <= a xor b;
    layer5_outputs(2648) <= a and not b;
    layer5_outputs(2649) <= not b;
    layer5_outputs(2650) <= not a;
    layer5_outputs(2651) <= not b;
    layer5_outputs(2652) <= not b;
    layer5_outputs(2653) <= a or b;
    layer5_outputs(2654) <= b;
    layer5_outputs(2655) <= not b or a;
    layer5_outputs(2656) <= not b;
    layer5_outputs(2657) <= a and not b;
    layer5_outputs(2658) <= a and not b;
    layer5_outputs(2659) <= '0';
    layer5_outputs(2660) <= not (a and b);
    layer5_outputs(2661) <= a or b;
    layer5_outputs(2662) <= a and b;
    layer5_outputs(2663) <= not b;
    layer5_outputs(2664) <= not a;
    layer5_outputs(2665) <= not (a or b);
    layer5_outputs(2666) <= not a or b;
    layer5_outputs(2667) <= '1';
    layer5_outputs(2668) <= '1';
    layer5_outputs(2669) <= not b or a;
    layer5_outputs(2670) <= a xor b;
    layer5_outputs(2671) <= b;
    layer5_outputs(2672) <= a and b;
    layer5_outputs(2673) <= not a;
    layer5_outputs(2674) <= not b or a;
    layer5_outputs(2675) <= a and not b;
    layer5_outputs(2676) <= not b;
    layer5_outputs(2677) <= a or b;
    layer5_outputs(2678) <= not a;
    layer5_outputs(2679) <= not a;
    layer5_outputs(2680) <= not b or a;
    layer5_outputs(2681) <= not (a or b);
    layer5_outputs(2682) <= not (a xor b);
    layer5_outputs(2683) <= b and not a;
    layer5_outputs(2684) <= not (a xor b);
    layer5_outputs(2685) <= a or b;
    layer5_outputs(2686) <= not (a or b);
    layer5_outputs(2687) <= a and not b;
    layer5_outputs(2688) <= a and b;
    layer5_outputs(2689) <= '0';
    layer5_outputs(2690) <= not a or b;
    layer5_outputs(2691) <= not (a and b);
    layer5_outputs(2692) <= a and not b;
    layer5_outputs(2693) <= not (a or b);
    layer5_outputs(2694) <= a and b;
    layer5_outputs(2695) <= not b;
    layer5_outputs(2696) <= not (a and b);
    layer5_outputs(2697) <= a;
    layer5_outputs(2698) <= b and not a;
    layer5_outputs(2699) <= not (a or b);
    layer5_outputs(2700) <= not b;
    layer5_outputs(2701) <= a and not b;
    layer5_outputs(2702) <= a and b;
    layer5_outputs(2703) <= not (a or b);
    layer5_outputs(2704) <= a;
    layer5_outputs(2705) <= not a or b;
    layer5_outputs(2706) <= not (a or b);
    layer5_outputs(2707) <= not b;
    layer5_outputs(2708) <= b;
    layer5_outputs(2709) <= a and b;
    layer5_outputs(2710) <= not (a and b);
    layer5_outputs(2711) <= not (a and b);
    layer5_outputs(2712) <= a and not b;
    layer5_outputs(2713) <= not (a and b);
    layer5_outputs(2714) <= not (a or b);
    layer5_outputs(2715) <= not a or b;
    layer5_outputs(2716) <= a;
    layer5_outputs(2717) <= not a or b;
    layer5_outputs(2718) <= a;
    layer5_outputs(2719) <= b;
    layer5_outputs(2720) <= not a or b;
    layer5_outputs(2721) <= not (a or b);
    layer5_outputs(2722) <= not (a xor b);
    layer5_outputs(2723) <= b;
    layer5_outputs(2724) <= not b;
    layer5_outputs(2725) <= b and not a;
    layer5_outputs(2726) <= a or b;
    layer5_outputs(2727) <= a and b;
    layer5_outputs(2728) <= not (a and b);
    layer5_outputs(2729) <= b;
    layer5_outputs(2730) <= not b or a;
    layer5_outputs(2731) <= a xor b;
    layer5_outputs(2732) <= a;
    layer5_outputs(2733) <= not a;
    layer5_outputs(2734) <= not (a xor b);
    layer5_outputs(2735) <= not b;
    layer5_outputs(2736) <= b and not a;
    layer5_outputs(2737) <= not b;
    layer5_outputs(2738) <= a and not b;
    layer5_outputs(2739) <= a or b;
    layer5_outputs(2740) <= not a;
    layer5_outputs(2741) <= not a;
    layer5_outputs(2742) <= b;
    layer5_outputs(2743) <= '1';
    layer5_outputs(2744) <= b and not a;
    layer5_outputs(2745) <= b;
    layer5_outputs(2746) <= a and b;
    layer5_outputs(2747) <= not (a and b);
    layer5_outputs(2748) <= a or b;
    layer5_outputs(2749) <= not (a and b);
    layer5_outputs(2750) <= a xor b;
    layer5_outputs(2751) <= '1';
    layer5_outputs(2752) <= b;
    layer5_outputs(2753) <= a;
    layer5_outputs(2754) <= a or b;
    layer5_outputs(2755) <= b and not a;
    layer5_outputs(2756) <= not a;
    layer5_outputs(2757) <= a and not b;
    layer5_outputs(2758) <= b;
    layer5_outputs(2759) <= a and b;
    layer5_outputs(2760) <= a or b;
    layer5_outputs(2761) <= b;
    layer5_outputs(2762) <= not b;
    layer5_outputs(2763) <= b;
    layer5_outputs(2764) <= '0';
    layer5_outputs(2765) <= not b or a;
    layer5_outputs(2766) <= a and b;
    layer5_outputs(2767) <= not (a and b);
    layer5_outputs(2768) <= not a or b;
    layer5_outputs(2769) <= not b;
    layer5_outputs(2770) <= not a or b;
    layer5_outputs(2771) <= not a;
    layer5_outputs(2772) <= b;
    layer5_outputs(2773) <= not a or b;
    layer5_outputs(2774) <= not (a xor b);
    layer5_outputs(2775) <= b;
    layer5_outputs(2776) <= '1';
    layer5_outputs(2777) <= not (a or b);
    layer5_outputs(2778) <= a and not b;
    layer5_outputs(2779) <= not b or a;
    layer5_outputs(2780) <= not b;
    layer5_outputs(2781) <= b and not a;
    layer5_outputs(2782) <= not b;
    layer5_outputs(2783) <= a xor b;
    layer5_outputs(2784) <= a and b;
    layer5_outputs(2785) <= a or b;
    layer5_outputs(2786) <= b and not a;
    layer5_outputs(2787) <= b;
    layer5_outputs(2788) <= '1';
    layer5_outputs(2789) <= b and not a;
    layer5_outputs(2790) <= b;
    layer5_outputs(2791) <= a and b;
    layer5_outputs(2792) <= not b;
    layer5_outputs(2793) <= b and not a;
    layer5_outputs(2794) <= '0';
    layer5_outputs(2795) <= b;
    layer5_outputs(2796) <= a or b;
    layer5_outputs(2797) <= b and not a;
    layer5_outputs(2798) <= a and not b;
    layer5_outputs(2799) <= '1';
    layer5_outputs(2800) <= not (a or b);
    layer5_outputs(2801) <= b;
    layer5_outputs(2802) <= '1';
    layer5_outputs(2803) <= not a;
    layer5_outputs(2804) <= a and b;
    layer5_outputs(2805) <= a and not b;
    layer5_outputs(2806) <= not a or b;
    layer5_outputs(2807) <= b and not a;
    layer5_outputs(2808) <= not a;
    layer5_outputs(2809) <= a and not b;
    layer5_outputs(2810) <= a and b;
    layer5_outputs(2811) <= not (a or b);
    layer5_outputs(2812) <= a and b;
    layer5_outputs(2813) <= not a;
    layer5_outputs(2814) <= a or b;
    layer5_outputs(2815) <= a;
    layer5_outputs(2816) <= not b;
    layer5_outputs(2817) <= b;
    layer5_outputs(2818) <= b;
    layer5_outputs(2819) <= not a or b;
    layer5_outputs(2820) <= b;
    layer5_outputs(2821) <= not (a and b);
    layer5_outputs(2822) <= not (a or b);
    layer5_outputs(2823) <= not b;
    layer5_outputs(2824) <= '1';
    layer5_outputs(2825) <= b;
    layer5_outputs(2826) <= not a;
    layer5_outputs(2827) <= '0';
    layer5_outputs(2828) <= b;
    layer5_outputs(2829) <= a;
    layer5_outputs(2830) <= a;
    layer5_outputs(2831) <= not a;
    layer5_outputs(2832) <= b;
    layer5_outputs(2833) <= '0';
    layer5_outputs(2834) <= not b;
    layer5_outputs(2835) <= b;
    layer5_outputs(2836) <= not (a or b);
    layer5_outputs(2837) <= a;
    layer5_outputs(2838) <= a;
    layer5_outputs(2839) <= b and not a;
    layer5_outputs(2840) <= '1';
    layer5_outputs(2841) <= a;
    layer5_outputs(2842) <= a and b;
    layer5_outputs(2843) <= b;
    layer5_outputs(2844) <= not (a and b);
    layer5_outputs(2845) <= a xor b;
    layer5_outputs(2846) <= a and b;
    layer5_outputs(2847) <= a and not b;
    layer5_outputs(2848) <= not (a xor b);
    layer5_outputs(2849) <= a and b;
    layer5_outputs(2850) <= a and not b;
    layer5_outputs(2851) <= not b;
    layer5_outputs(2852) <= not b or a;
    layer5_outputs(2853) <= not (a and b);
    layer5_outputs(2854) <= a and b;
    layer5_outputs(2855) <= a and b;
    layer5_outputs(2856) <= a;
    layer5_outputs(2857) <= not a;
    layer5_outputs(2858) <= b;
    layer5_outputs(2859) <= not a;
    layer5_outputs(2860) <= b;
    layer5_outputs(2861) <= b;
    layer5_outputs(2862) <= a;
    layer5_outputs(2863) <= not a or b;
    layer5_outputs(2864) <= a xor b;
    layer5_outputs(2865) <= '1';
    layer5_outputs(2866) <= a and b;
    layer5_outputs(2867) <= not b or a;
    layer5_outputs(2868) <= b and not a;
    layer5_outputs(2869) <= not b;
    layer5_outputs(2870) <= not b or a;
    layer5_outputs(2871) <= a;
    layer5_outputs(2872) <= '1';
    layer5_outputs(2873) <= a and not b;
    layer5_outputs(2874) <= not b;
    layer5_outputs(2875) <= a;
    layer5_outputs(2876) <= not b;
    layer5_outputs(2877) <= b and not a;
    layer5_outputs(2878) <= b and not a;
    layer5_outputs(2879) <= not a;
    layer5_outputs(2880) <= a xor b;
    layer5_outputs(2881) <= a and not b;
    layer5_outputs(2882) <= b;
    layer5_outputs(2883) <= not a or b;
    layer5_outputs(2884) <= not (a or b);
    layer5_outputs(2885) <= not a or b;
    layer5_outputs(2886) <= not (a and b);
    layer5_outputs(2887) <= a or b;
    layer5_outputs(2888) <= b;
    layer5_outputs(2889) <= b and not a;
    layer5_outputs(2890) <= not a;
    layer5_outputs(2891) <= '0';
    layer5_outputs(2892) <= not a or b;
    layer5_outputs(2893) <= not b or a;
    layer5_outputs(2894) <= not a;
    layer5_outputs(2895) <= b;
    layer5_outputs(2896) <= a or b;
    layer5_outputs(2897) <= not (a or b);
    layer5_outputs(2898) <= a xor b;
    layer5_outputs(2899) <= b;
    layer5_outputs(2900) <= not b;
    layer5_outputs(2901) <= not (a or b);
    layer5_outputs(2902) <= a and b;
    layer5_outputs(2903) <= not b or a;
    layer5_outputs(2904) <= not b;
    layer5_outputs(2905) <= not (a and b);
    layer5_outputs(2906) <= b and not a;
    layer5_outputs(2907) <= not b;
    layer5_outputs(2908) <= a and not b;
    layer5_outputs(2909) <= b;
    layer5_outputs(2910) <= not a;
    layer5_outputs(2911) <= b;
    layer5_outputs(2912) <= b;
    layer5_outputs(2913) <= b and not a;
    layer5_outputs(2914) <= a;
    layer5_outputs(2915) <= not a;
    layer5_outputs(2916) <= a and not b;
    layer5_outputs(2917) <= a and not b;
    layer5_outputs(2918) <= a or b;
    layer5_outputs(2919) <= not a or b;
    layer5_outputs(2920) <= b;
    layer5_outputs(2921) <= not (a or b);
    layer5_outputs(2922) <= not a;
    layer5_outputs(2923) <= not a or b;
    layer5_outputs(2924) <= '0';
    layer5_outputs(2925) <= not b;
    layer5_outputs(2926) <= not a or b;
    layer5_outputs(2927) <= a;
    layer5_outputs(2928) <= '1';
    layer5_outputs(2929) <= not (a and b);
    layer5_outputs(2930) <= a or b;
    layer5_outputs(2931) <= a and b;
    layer5_outputs(2932) <= b and not a;
    layer5_outputs(2933) <= a and b;
    layer5_outputs(2934) <= not (a xor b);
    layer5_outputs(2935) <= a;
    layer5_outputs(2936) <= a or b;
    layer5_outputs(2937) <= a;
    layer5_outputs(2938) <= a and not b;
    layer5_outputs(2939) <= not b;
    layer5_outputs(2940) <= not (a xor b);
    layer5_outputs(2941) <= not b;
    layer5_outputs(2942) <= not b or a;
    layer5_outputs(2943) <= '1';
    layer5_outputs(2944) <= a or b;
    layer5_outputs(2945) <= not a;
    layer5_outputs(2946) <= '0';
    layer5_outputs(2947) <= a and not b;
    layer5_outputs(2948) <= a and not b;
    layer5_outputs(2949) <= a and not b;
    layer5_outputs(2950) <= not b;
    layer5_outputs(2951) <= not b;
    layer5_outputs(2952) <= not (a and b);
    layer5_outputs(2953) <= not a or b;
    layer5_outputs(2954) <= a or b;
    layer5_outputs(2955) <= '0';
    layer5_outputs(2956) <= not (a xor b);
    layer5_outputs(2957) <= not a or b;
    layer5_outputs(2958) <= b;
    layer5_outputs(2959) <= not b or a;
    layer5_outputs(2960) <= not b or a;
    layer5_outputs(2961) <= a;
    layer5_outputs(2962) <= not (a and b);
    layer5_outputs(2963) <= a and not b;
    layer5_outputs(2964) <= b;
    layer5_outputs(2965) <= a and b;
    layer5_outputs(2966) <= not (a or b);
    layer5_outputs(2967) <= not a;
    layer5_outputs(2968) <= a or b;
    layer5_outputs(2969) <= a xor b;
    layer5_outputs(2970) <= b;
    layer5_outputs(2971) <= not (a and b);
    layer5_outputs(2972) <= not a;
    layer5_outputs(2973) <= '0';
    layer5_outputs(2974) <= a and not b;
    layer5_outputs(2975) <= not (a xor b);
    layer5_outputs(2976) <= not a;
    layer5_outputs(2977) <= a and not b;
    layer5_outputs(2978) <= not b or a;
    layer5_outputs(2979) <= a or b;
    layer5_outputs(2980) <= not (a and b);
    layer5_outputs(2981) <= not (a xor b);
    layer5_outputs(2982) <= not b or a;
    layer5_outputs(2983) <= a xor b;
    layer5_outputs(2984) <= not b or a;
    layer5_outputs(2985) <= not b or a;
    layer5_outputs(2986) <= not a;
    layer5_outputs(2987) <= not a or b;
    layer5_outputs(2988) <= b and not a;
    layer5_outputs(2989) <= a or b;
    layer5_outputs(2990) <= not (a and b);
    layer5_outputs(2991) <= not a or b;
    layer5_outputs(2992) <= '1';
    layer5_outputs(2993) <= not (a xor b);
    layer5_outputs(2994) <= a;
    layer5_outputs(2995) <= not (a and b);
    layer5_outputs(2996) <= a;
    layer5_outputs(2997) <= a;
    layer5_outputs(2998) <= not a or b;
    layer5_outputs(2999) <= not (a or b);
    layer5_outputs(3000) <= b;
    layer5_outputs(3001) <= not b or a;
    layer5_outputs(3002) <= a;
    layer5_outputs(3003) <= not b;
    layer5_outputs(3004) <= not b or a;
    layer5_outputs(3005) <= not (a or b);
    layer5_outputs(3006) <= not (a and b);
    layer5_outputs(3007) <= not (a and b);
    layer5_outputs(3008) <= a or b;
    layer5_outputs(3009) <= not a;
    layer5_outputs(3010) <= b;
    layer5_outputs(3011) <= a xor b;
    layer5_outputs(3012) <= a and not b;
    layer5_outputs(3013) <= a and not b;
    layer5_outputs(3014) <= not b or a;
    layer5_outputs(3015) <= not b;
    layer5_outputs(3016) <= not a;
    layer5_outputs(3017) <= not a or b;
    layer5_outputs(3018) <= a and not b;
    layer5_outputs(3019) <= not (a or b);
    layer5_outputs(3020) <= not b;
    layer5_outputs(3021) <= a xor b;
    layer5_outputs(3022) <= b;
    layer5_outputs(3023) <= not b;
    layer5_outputs(3024) <= not a;
    layer5_outputs(3025) <= b;
    layer5_outputs(3026) <= '0';
    layer5_outputs(3027) <= not b;
    layer5_outputs(3028) <= a and not b;
    layer5_outputs(3029) <= not b or a;
    layer5_outputs(3030) <= not b or a;
    layer5_outputs(3031) <= not a;
    layer5_outputs(3032) <= b and not a;
    layer5_outputs(3033) <= a and not b;
    layer5_outputs(3034) <= not (a or b);
    layer5_outputs(3035) <= a and not b;
    layer5_outputs(3036) <= not b;
    layer5_outputs(3037) <= b;
    layer5_outputs(3038) <= a xor b;
    layer5_outputs(3039) <= not (a and b);
    layer5_outputs(3040) <= a;
    layer5_outputs(3041) <= not (a xor b);
    layer5_outputs(3042) <= a xor b;
    layer5_outputs(3043) <= a;
    layer5_outputs(3044) <= '0';
    layer5_outputs(3045) <= not b or a;
    layer5_outputs(3046) <= not (a or b);
    layer5_outputs(3047) <= b;
    layer5_outputs(3048) <= not a;
    layer5_outputs(3049) <= b;
    layer5_outputs(3050) <= '0';
    layer5_outputs(3051) <= not b;
    layer5_outputs(3052) <= not b;
    layer5_outputs(3053) <= not b;
    layer5_outputs(3054) <= not (a or b);
    layer5_outputs(3055) <= not a or b;
    layer5_outputs(3056) <= '1';
    layer5_outputs(3057) <= '0';
    layer5_outputs(3058) <= not (a or b);
    layer5_outputs(3059) <= not a;
    layer5_outputs(3060) <= a or b;
    layer5_outputs(3061) <= not (a xor b);
    layer5_outputs(3062) <= not b;
    layer5_outputs(3063) <= a xor b;
    layer5_outputs(3064) <= '0';
    layer5_outputs(3065) <= not (a or b);
    layer5_outputs(3066) <= not a;
    layer5_outputs(3067) <= a;
    layer5_outputs(3068) <= a and not b;
    layer5_outputs(3069) <= not (a xor b);
    layer5_outputs(3070) <= not b;
    layer5_outputs(3071) <= a and not b;
    layer5_outputs(3072) <= '1';
    layer5_outputs(3073) <= a;
    layer5_outputs(3074) <= a and not b;
    layer5_outputs(3075) <= a and not b;
    layer5_outputs(3076) <= not b;
    layer5_outputs(3077) <= not a;
    layer5_outputs(3078) <= b and not a;
    layer5_outputs(3079) <= not b;
    layer5_outputs(3080) <= a or b;
    layer5_outputs(3081) <= a and not b;
    layer5_outputs(3082) <= a or b;
    layer5_outputs(3083) <= a and not b;
    layer5_outputs(3084) <= b;
    layer5_outputs(3085) <= a and not b;
    layer5_outputs(3086) <= a and b;
    layer5_outputs(3087) <= not a;
    layer5_outputs(3088) <= a xor b;
    layer5_outputs(3089) <= a or b;
    layer5_outputs(3090) <= a;
    layer5_outputs(3091) <= a;
    layer5_outputs(3092) <= a and b;
    layer5_outputs(3093) <= b;
    layer5_outputs(3094) <= not b or a;
    layer5_outputs(3095) <= not (a or b);
    layer5_outputs(3096) <= not (a or b);
    layer5_outputs(3097) <= not (a xor b);
    layer5_outputs(3098) <= not (a xor b);
    layer5_outputs(3099) <= a or b;
    layer5_outputs(3100) <= not (a or b);
    layer5_outputs(3101) <= not a;
    layer5_outputs(3102) <= not b;
    layer5_outputs(3103) <= not a or b;
    layer5_outputs(3104) <= not a or b;
    layer5_outputs(3105) <= not b;
    layer5_outputs(3106) <= not b;
    layer5_outputs(3107) <= a xor b;
    layer5_outputs(3108) <= not a or b;
    layer5_outputs(3109) <= '0';
    layer5_outputs(3110) <= not a or b;
    layer5_outputs(3111) <= not a;
    layer5_outputs(3112) <= not (a or b);
    layer5_outputs(3113) <= not b or a;
    layer5_outputs(3114) <= not a or b;
    layer5_outputs(3115) <= a xor b;
    layer5_outputs(3116) <= a and b;
    layer5_outputs(3117) <= not a;
    layer5_outputs(3118) <= not a;
    layer5_outputs(3119) <= not a;
    layer5_outputs(3120) <= a or b;
    layer5_outputs(3121) <= not a or b;
    layer5_outputs(3122) <= not (a xor b);
    layer5_outputs(3123) <= a and not b;
    layer5_outputs(3124) <= not a;
    layer5_outputs(3125) <= not (a xor b);
    layer5_outputs(3126) <= a and not b;
    layer5_outputs(3127) <= a and b;
    layer5_outputs(3128) <= a and b;
    layer5_outputs(3129) <= a and not b;
    layer5_outputs(3130) <= a and b;
    layer5_outputs(3131) <= b;
    layer5_outputs(3132) <= not (a or b);
    layer5_outputs(3133) <= a and not b;
    layer5_outputs(3134) <= not b or a;
    layer5_outputs(3135) <= a;
    layer5_outputs(3136) <= a or b;
    layer5_outputs(3137) <= not (a xor b);
    layer5_outputs(3138) <= not a;
    layer5_outputs(3139) <= not b or a;
    layer5_outputs(3140) <= '0';
    layer5_outputs(3141) <= a or b;
    layer5_outputs(3142) <= '1';
    layer5_outputs(3143) <= not a or b;
    layer5_outputs(3144) <= not a or b;
    layer5_outputs(3145) <= not a or b;
    layer5_outputs(3146) <= b;
    layer5_outputs(3147) <= not (a xor b);
    layer5_outputs(3148) <= b;
    layer5_outputs(3149) <= not a or b;
    layer5_outputs(3150) <= a;
    layer5_outputs(3151) <= not b;
    layer5_outputs(3152) <= b;
    layer5_outputs(3153) <= not a or b;
    layer5_outputs(3154) <= not a;
    layer5_outputs(3155) <= a and not b;
    layer5_outputs(3156) <= a and b;
    layer5_outputs(3157) <= not a;
    layer5_outputs(3158) <= a and b;
    layer5_outputs(3159) <= a xor b;
    layer5_outputs(3160) <= not b;
    layer5_outputs(3161) <= not (a or b);
    layer5_outputs(3162) <= not b or a;
    layer5_outputs(3163) <= '1';
    layer5_outputs(3164) <= not b;
    layer5_outputs(3165) <= a;
    layer5_outputs(3166) <= a;
    layer5_outputs(3167) <= not b or a;
    layer5_outputs(3168) <= a xor b;
    layer5_outputs(3169) <= not (a and b);
    layer5_outputs(3170) <= not a;
    layer5_outputs(3171) <= a and b;
    layer5_outputs(3172) <= not (a or b);
    layer5_outputs(3173) <= '0';
    layer5_outputs(3174) <= not b or a;
    layer5_outputs(3175) <= not (a xor b);
    layer5_outputs(3176) <= not a or b;
    layer5_outputs(3177) <= a and not b;
    layer5_outputs(3178) <= a or b;
    layer5_outputs(3179) <= not (a or b);
    layer5_outputs(3180) <= not b;
    layer5_outputs(3181) <= a xor b;
    layer5_outputs(3182) <= not b or a;
    layer5_outputs(3183) <= not a;
    layer5_outputs(3184) <= a or b;
    layer5_outputs(3185) <= not b or a;
    layer5_outputs(3186) <= b;
    layer5_outputs(3187) <= a;
    layer5_outputs(3188) <= not a;
    layer5_outputs(3189) <= a or b;
    layer5_outputs(3190) <= '1';
    layer5_outputs(3191) <= a;
    layer5_outputs(3192) <= a;
    layer5_outputs(3193) <= a and not b;
    layer5_outputs(3194) <= not a or b;
    layer5_outputs(3195) <= not b;
    layer5_outputs(3196) <= b;
    layer5_outputs(3197) <= a;
    layer5_outputs(3198) <= b;
    layer5_outputs(3199) <= b;
    layer5_outputs(3200) <= not b;
    layer5_outputs(3201) <= a and not b;
    layer5_outputs(3202) <= not a or b;
    layer5_outputs(3203) <= not a;
    layer5_outputs(3204) <= not a or b;
    layer5_outputs(3205) <= not b;
    layer5_outputs(3206) <= not a;
    layer5_outputs(3207) <= a and b;
    layer5_outputs(3208) <= a and b;
    layer5_outputs(3209) <= not (a and b);
    layer5_outputs(3210) <= b;
    layer5_outputs(3211) <= b;
    layer5_outputs(3212) <= a xor b;
    layer5_outputs(3213) <= not (a or b);
    layer5_outputs(3214) <= not (a and b);
    layer5_outputs(3215) <= not b;
    layer5_outputs(3216) <= a and b;
    layer5_outputs(3217) <= a;
    layer5_outputs(3218) <= a xor b;
    layer5_outputs(3219) <= b and not a;
    layer5_outputs(3220) <= '0';
    layer5_outputs(3221) <= not b or a;
    layer5_outputs(3222) <= a xor b;
    layer5_outputs(3223) <= b and not a;
    layer5_outputs(3224) <= not (a or b);
    layer5_outputs(3225) <= not a or b;
    layer5_outputs(3226) <= a and b;
    layer5_outputs(3227) <= not (a and b);
    layer5_outputs(3228) <= not a or b;
    layer5_outputs(3229) <= a and not b;
    layer5_outputs(3230) <= not a;
    layer5_outputs(3231) <= b;
    layer5_outputs(3232) <= not a;
    layer5_outputs(3233) <= a and b;
    layer5_outputs(3234) <= not (a or b);
    layer5_outputs(3235) <= not (a and b);
    layer5_outputs(3236) <= not b or a;
    layer5_outputs(3237) <= not (a and b);
    layer5_outputs(3238) <= not (a and b);
    layer5_outputs(3239) <= not a;
    layer5_outputs(3240) <= not (a and b);
    layer5_outputs(3241) <= not (a and b);
    layer5_outputs(3242) <= not a or b;
    layer5_outputs(3243) <= '1';
    layer5_outputs(3244) <= not a;
    layer5_outputs(3245) <= a and not b;
    layer5_outputs(3246) <= not (a or b);
    layer5_outputs(3247) <= b;
    layer5_outputs(3248) <= a and not b;
    layer5_outputs(3249) <= b;
    layer5_outputs(3250) <= a xor b;
    layer5_outputs(3251) <= '0';
    layer5_outputs(3252) <= a xor b;
    layer5_outputs(3253) <= not (a or b);
    layer5_outputs(3254) <= not b;
    layer5_outputs(3255) <= a and b;
    layer5_outputs(3256) <= not a;
    layer5_outputs(3257) <= '1';
    layer5_outputs(3258) <= not b or a;
    layer5_outputs(3259) <= '1';
    layer5_outputs(3260) <= b and not a;
    layer5_outputs(3261) <= a or b;
    layer5_outputs(3262) <= not (a and b);
    layer5_outputs(3263) <= not a or b;
    layer5_outputs(3264) <= a or b;
    layer5_outputs(3265) <= a or b;
    layer5_outputs(3266) <= b;
    layer5_outputs(3267) <= a;
    layer5_outputs(3268) <= b;
    layer5_outputs(3269) <= not a;
    layer5_outputs(3270) <= not b;
    layer5_outputs(3271) <= not (a or b);
    layer5_outputs(3272) <= not b or a;
    layer5_outputs(3273) <= not (a or b);
    layer5_outputs(3274) <= not b;
    layer5_outputs(3275) <= a xor b;
    layer5_outputs(3276) <= not (a or b);
    layer5_outputs(3277) <= b;
    layer5_outputs(3278) <= not (a or b);
    layer5_outputs(3279) <= b;
    layer5_outputs(3280) <= a and b;
    layer5_outputs(3281) <= not b or a;
    layer5_outputs(3282) <= '0';
    layer5_outputs(3283) <= not (a and b);
    layer5_outputs(3284) <= not a;
    layer5_outputs(3285) <= a;
    layer5_outputs(3286) <= not b;
    layer5_outputs(3287) <= not b or a;
    layer5_outputs(3288) <= a or b;
    layer5_outputs(3289) <= not a or b;
    layer5_outputs(3290) <= not a;
    layer5_outputs(3291) <= '0';
    layer5_outputs(3292) <= a xor b;
    layer5_outputs(3293) <= not b or a;
    layer5_outputs(3294) <= a or b;
    layer5_outputs(3295) <= not a;
    layer5_outputs(3296) <= '0';
    layer5_outputs(3297) <= b;
    layer5_outputs(3298) <= not b;
    layer5_outputs(3299) <= not a or b;
    layer5_outputs(3300) <= b;
    layer5_outputs(3301) <= not (a and b);
    layer5_outputs(3302) <= not b;
    layer5_outputs(3303) <= a and b;
    layer5_outputs(3304) <= not a or b;
    layer5_outputs(3305) <= not b;
    layer5_outputs(3306) <= not b or a;
    layer5_outputs(3307) <= a or b;
    layer5_outputs(3308) <= a and b;
    layer5_outputs(3309) <= a xor b;
    layer5_outputs(3310) <= not (a xor b);
    layer5_outputs(3311) <= a;
    layer5_outputs(3312) <= a;
    layer5_outputs(3313) <= not (a xor b);
    layer5_outputs(3314) <= a and not b;
    layer5_outputs(3315) <= a or b;
    layer5_outputs(3316) <= not a or b;
    layer5_outputs(3317) <= a and b;
    layer5_outputs(3318) <= b;
    layer5_outputs(3319) <= not (a and b);
    layer5_outputs(3320) <= a and b;
    layer5_outputs(3321) <= '0';
    layer5_outputs(3322) <= a xor b;
    layer5_outputs(3323) <= a and not b;
    layer5_outputs(3324) <= b;
    layer5_outputs(3325) <= b;
    layer5_outputs(3326) <= not b or a;
    layer5_outputs(3327) <= not b or a;
    layer5_outputs(3328) <= b and not a;
    layer5_outputs(3329) <= not b;
    layer5_outputs(3330) <= not (a or b);
    layer5_outputs(3331) <= a and b;
    layer5_outputs(3332) <= not (a or b);
    layer5_outputs(3333) <= not (a and b);
    layer5_outputs(3334) <= not (a xor b);
    layer5_outputs(3335) <= a and b;
    layer5_outputs(3336) <= not (a or b);
    layer5_outputs(3337) <= not b;
    layer5_outputs(3338) <= b;
    layer5_outputs(3339) <= not b;
    layer5_outputs(3340) <= a;
    layer5_outputs(3341) <= not b or a;
    layer5_outputs(3342) <= a and not b;
    layer5_outputs(3343) <= not b or a;
    layer5_outputs(3344) <= not b;
    layer5_outputs(3345) <= not a;
    layer5_outputs(3346) <= b;
    layer5_outputs(3347) <= '1';
    layer5_outputs(3348) <= not b;
    layer5_outputs(3349) <= '1';
    layer5_outputs(3350) <= not (a and b);
    layer5_outputs(3351) <= not (a and b);
    layer5_outputs(3352) <= not b;
    layer5_outputs(3353) <= not a or b;
    layer5_outputs(3354) <= b;
    layer5_outputs(3355) <= '1';
    layer5_outputs(3356) <= not a or b;
    layer5_outputs(3357) <= a and b;
    layer5_outputs(3358) <= not b;
    layer5_outputs(3359) <= not a;
    layer5_outputs(3360) <= not a;
    layer5_outputs(3361) <= not a;
    layer5_outputs(3362) <= b;
    layer5_outputs(3363) <= a xor b;
    layer5_outputs(3364) <= not (a or b);
    layer5_outputs(3365) <= a and b;
    layer5_outputs(3366) <= a;
    layer5_outputs(3367) <= not b;
    layer5_outputs(3368) <= not (a and b);
    layer5_outputs(3369) <= not b;
    layer5_outputs(3370) <= a;
    layer5_outputs(3371) <= '1';
    layer5_outputs(3372) <= b and not a;
    layer5_outputs(3373) <= not (a and b);
    layer5_outputs(3374) <= a;
    layer5_outputs(3375) <= a xor b;
    layer5_outputs(3376) <= b;
    layer5_outputs(3377) <= a and b;
    layer5_outputs(3378) <= b and not a;
    layer5_outputs(3379) <= a and b;
    layer5_outputs(3380) <= not (a and b);
    layer5_outputs(3381) <= a and not b;
    layer5_outputs(3382) <= not (a and b);
    layer5_outputs(3383) <= b and not a;
    layer5_outputs(3384) <= not a;
    layer5_outputs(3385) <= not a;
    layer5_outputs(3386) <= not a;
    layer5_outputs(3387) <= not (a and b);
    layer5_outputs(3388) <= a and not b;
    layer5_outputs(3389) <= b and not a;
    layer5_outputs(3390) <= not a;
    layer5_outputs(3391) <= b and not a;
    layer5_outputs(3392) <= not a;
    layer5_outputs(3393) <= a;
    layer5_outputs(3394) <= not a or b;
    layer5_outputs(3395) <= a and not b;
    layer5_outputs(3396) <= '0';
    layer5_outputs(3397) <= b and not a;
    layer5_outputs(3398) <= not b;
    layer5_outputs(3399) <= b;
    layer5_outputs(3400) <= a and not b;
    layer5_outputs(3401) <= not b;
    layer5_outputs(3402) <= a;
    layer5_outputs(3403) <= not (a or b);
    layer5_outputs(3404) <= not (a and b);
    layer5_outputs(3405) <= not (a and b);
    layer5_outputs(3406) <= not b;
    layer5_outputs(3407) <= '0';
    layer5_outputs(3408) <= a;
    layer5_outputs(3409) <= not b;
    layer5_outputs(3410) <= b;
    layer5_outputs(3411) <= a and not b;
    layer5_outputs(3412) <= not a;
    layer5_outputs(3413) <= b and not a;
    layer5_outputs(3414) <= not a or b;
    layer5_outputs(3415) <= b;
    layer5_outputs(3416) <= not b or a;
    layer5_outputs(3417) <= a xor b;
    layer5_outputs(3418) <= '0';
    layer5_outputs(3419) <= not (a or b);
    layer5_outputs(3420) <= b;
    layer5_outputs(3421) <= not (a and b);
    layer5_outputs(3422) <= not (a and b);
    layer5_outputs(3423) <= not (a and b);
    layer5_outputs(3424) <= not (a or b);
    layer5_outputs(3425) <= not a;
    layer5_outputs(3426) <= '1';
    layer5_outputs(3427) <= b;
    layer5_outputs(3428) <= b;
    layer5_outputs(3429) <= a;
    layer5_outputs(3430) <= b;
    layer5_outputs(3431) <= not a;
    layer5_outputs(3432) <= not a;
    layer5_outputs(3433) <= not a;
    layer5_outputs(3434) <= '1';
    layer5_outputs(3435) <= not b;
    layer5_outputs(3436) <= a and b;
    layer5_outputs(3437) <= not a;
    layer5_outputs(3438) <= a;
    layer5_outputs(3439) <= not b or a;
    layer5_outputs(3440) <= b and not a;
    layer5_outputs(3441) <= not b;
    layer5_outputs(3442) <= '1';
    layer5_outputs(3443) <= not (a and b);
    layer5_outputs(3444) <= a;
    layer5_outputs(3445) <= b;
    layer5_outputs(3446) <= a and not b;
    layer5_outputs(3447) <= b and not a;
    layer5_outputs(3448) <= a and b;
    layer5_outputs(3449) <= not b;
    layer5_outputs(3450) <= a and not b;
    layer5_outputs(3451) <= a;
    layer5_outputs(3452) <= not (a or b);
    layer5_outputs(3453) <= not b or a;
    layer5_outputs(3454) <= '0';
    layer5_outputs(3455) <= b;
    layer5_outputs(3456) <= not a;
    layer5_outputs(3457) <= a;
    layer5_outputs(3458) <= a or b;
    layer5_outputs(3459) <= not a;
    layer5_outputs(3460) <= not (a or b);
    layer5_outputs(3461) <= not a or b;
    layer5_outputs(3462) <= not (a and b);
    layer5_outputs(3463) <= not a;
    layer5_outputs(3464) <= not a or b;
    layer5_outputs(3465) <= b;
    layer5_outputs(3466) <= a;
    layer5_outputs(3467) <= not a;
    layer5_outputs(3468) <= a;
    layer5_outputs(3469) <= b;
    layer5_outputs(3470) <= not b;
    layer5_outputs(3471) <= a;
    layer5_outputs(3472) <= b and not a;
    layer5_outputs(3473) <= not b;
    layer5_outputs(3474) <= a or b;
    layer5_outputs(3475) <= a and not b;
    layer5_outputs(3476) <= '1';
    layer5_outputs(3477) <= not (a xor b);
    layer5_outputs(3478) <= a and b;
    layer5_outputs(3479) <= not a or b;
    layer5_outputs(3480) <= a or b;
    layer5_outputs(3481) <= not (a or b);
    layer5_outputs(3482) <= not (a and b);
    layer5_outputs(3483) <= a;
    layer5_outputs(3484) <= not b;
    layer5_outputs(3485) <= b and not a;
    layer5_outputs(3486) <= a;
    layer5_outputs(3487) <= a and not b;
    layer5_outputs(3488) <= not b;
    layer5_outputs(3489) <= not b;
    layer5_outputs(3490) <= a and not b;
    layer5_outputs(3491) <= '0';
    layer5_outputs(3492) <= not b;
    layer5_outputs(3493) <= b and not a;
    layer5_outputs(3494) <= a and b;
    layer5_outputs(3495) <= not b or a;
    layer5_outputs(3496) <= a or b;
    layer5_outputs(3497) <= not a;
    layer5_outputs(3498) <= not b;
    layer5_outputs(3499) <= '0';
    layer5_outputs(3500) <= a;
    layer5_outputs(3501) <= a;
    layer5_outputs(3502) <= not b or a;
    layer5_outputs(3503) <= '0';
    layer5_outputs(3504) <= not (a and b);
    layer5_outputs(3505) <= not b;
    layer5_outputs(3506) <= a and not b;
    layer5_outputs(3507) <= a;
    layer5_outputs(3508) <= b;
    layer5_outputs(3509) <= '1';
    layer5_outputs(3510) <= a or b;
    layer5_outputs(3511) <= not b or a;
    layer5_outputs(3512) <= not b;
    layer5_outputs(3513) <= not b or a;
    layer5_outputs(3514) <= a and b;
    layer5_outputs(3515) <= a or b;
    layer5_outputs(3516) <= b and not a;
    layer5_outputs(3517) <= a;
    layer5_outputs(3518) <= a and not b;
    layer5_outputs(3519) <= not (a and b);
    layer5_outputs(3520) <= not a or b;
    layer5_outputs(3521) <= a;
    layer5_outputs(3522) <= a and not b;
    layer5_outputs(3523) <= a or b;
    layer5_outputs(3524) <= not (a and b);
    layer5_outputs(3525) <= b;
    layer5_outputs(3526) <= a;
    layer5_outputs(3527) <= not (a or b);
    layer5_outputs(3528) <= not (a or b);
    layer5_outputs(3529) <= b;
    layer5_outputs(3530) <= not (a and b);
    layer5_outputs(3531) <= '0';
    layer5_outputs(3532) <= not (a and b);
    layer5_outputs(3533) <= a;
    layer5_outputs(3534) <= a;
    layer5_outputs(3535) <= not a or b;
    layer5_outputs(3536) <= a and not b;
    layer5_outputs(3537) <= not (a or b);
    layer5_outputs(3538) <= not b;
    layer5_outputs(3539) <= not b;
    layer5_outputs(3540) <= a and b;
    layer5_outputs(3541) <= b and not a;
    layer5_outputs(3542) <= b;
    layer5_outputs(3543) <= '0';
    layer5_outputs(3544) <= not (a or b);
    layer5_outputs(3545) <= not a;
    layer5_outputs(3546) <= b;
    layer5_outputs(3547) <= b;
    layer5_outputs(3548) <= not b;
    layer5_outputs(3549) <= not b;
    layer5_outputs(3550) <= b;
    layer5_outputs(3551) <= a or b;
    layer5_outputs(3552) <= a;
    layer5_outputs(3553) <= b;
    layer5_outputs(3554) <= a and b;
    layer5_outputs(3555) <= a xor b;
    layer5_outputs(3556) <= b;
    layer5_outputs(3557) <= not b;
    layer5_outputs(3558) <= a or b;
    layer5_outputs(3559) <= b and not a;
    layer5_outputs(3560) <= '0';
    layer5_outputs(3561) <= b;
    layer5_outputs(3562) <= not a or b;
    layer5_outputs(3563) <= a and not b;
    layer5_outputs(3564) <= '1';
    layer5_outputs(3565) <= not b or a;
    layer5_outputs(3566) <= '0';
    layer5_outputs(3567) <= not a;
    layer5_outputs(3568) <= b;
    layer5_outputs(3569) <= not (a or b);
    layer5_outputs(3570) <= a xor b;
    layer5_outputs(3571) <= '1';
    layer5_outputs(3572) <= not (a xor b);
    layer5_outputs(3573) <= not a;
    layer5_outputs(3574) <= not (a or b);
    layer5_outputs(3575) <= not (a xor b);
    layer5_outputs(3576) <= not a;
    layer5_outputs(3577) <= a and b;
    layer5_outputs(3578) <= not a;
    layer5_outputs(3579) <= a xor b;
    layer5_outputs(3580) <= b and not a;
    layer5_outputs(3581) <= not (a and b);
    layer5_outputs(3582) <= a;
    layer5_outputs(3583) <= a;
    layer5_outputs(3584) <= not b or a;
    layer5_outputs(3585) <= '1';
    layer5_outputs(3586) <= not a;
    layer5_outputs(3587) <= not (a xor b);
    layer5_outputs(3588) <= '1';
    layer5_outputs(3589) <= not (a or b);
    layer5_outputs(3590) <= b;
    layer5_outputs(3591) <= not b or a;
    layer5_outputs(3592) <= a and not b;
    layer5_outputs(3593) <= not a;
    layer5_outputs(3594) <= not (a or b);
    layer5_outputs(3595) <= not (a or b);
    layer5_outputs(3596) <= not b;
    layer5_outputs(3597) <= not b or a;
    layer5_outputs(3598) <= a and b;
    layer5_outputs(3599) <= not b;
    layer5_outputs(3600) <= b;
    layer5_outputs(3601) <= b;
    layer5_outputs(3602) <= a;
    layer5_outputs(3603) <= a;
    layer5_outputs(3604) <= a;
    layer5_outputs(3605) <= '1';
    layer5_outputs(3606) <= a and not b;
    layer5_outputs(3607) <= a or b;
    layer5_outputs(3608) <= a and not b;
    layer5_outputs(3609) <= not a;
    layer5_outputs(3610) <= not b;
    layer5_outputs(3611) <= b and not a;
    layer5_outputs(3612) <= b;
    layer5_outputs(3613) <= '0';
    layer5_outputs(3614) <= not b;
    layer5_outputs(3615) <= not (a or b);
    layer5_outputs(3616) <= not (a and b);
    layer5_outputs(3617) <= a and b;
    layer5_outputs(3618) <= b and not a;
    layer5_outputs(3619) <= not b;
    layer5_outputs(3620) <= not a;
    layer5_outputs(3621) <= not (a xor b);
    layer5_outputs(3622) <= not b;
    layer5_outputs(3623) <= b;
    layer5_outputs(3624) <= a;
    layer5_outputs(3625) <= not a;
    layer5_outputs(3626) <= not b;
    layer5_outputs(3627) <= a;
    layer5_outputs(3628) <= a or b;
    layer5_outputs(3629) <= not (a xor b);
    layer5_outputs(3630) <= not (a or b);
    layer5_outputs(3631) <= a;
    layer5_outputs(3632) <= not a;
    layer5_outputs(3633) <= not a;
    layer5_outputs(3634) <= a;
    layer5_outputs(3635) <= not a or b;
    layer5_outputs(3636) <= '0';
    layer5_outputs(3637) <= a xor b;
    layer5_outputs(3638) <= not (a or b);
    layer5_outputs(3639) <= a;
    layer5_outputs(3640) <= not (a and b);
    layer5_outputs(3641) <= not a;
    layer5_outputs(3642) <= not a or b;
    layer5_outputs(3643) <= not (a and b);
    layer5_outputs(3644) <= b and not a;
    layer5_outputs(3645) <= not b or a;
    layer5_outputs(3646) <= a and not b;
    layer5_outputs(3647) <= not b;
    layer5_outputs(3648) <= '1';
    layer5_outputs(3649) <= b and not a;
    layer5_outputs(3650) <= not (a xor b);
    layer5_outputs(3651) <= not (a and b);
    layer5_outputs(3652) <= b;
    layer5_outputs(3653) <= not a;
    layer5_outputs(3654) <= not a;
    layer5_outputs(3655) <= b;
    layer5_outputs(3656) <= a and not b;
    layer5_outputs(3657) <= not a;
    layer5_outputs(3658) <= a and b;
    layer5_outputs(3659) <= '0';
    layer5_outputs(3660) <= '0';
    layer5_outputs(3661) <= a and not b;
    layer5_outputs(3662) <= a and b;
    layer5_outputs(3663) <= a or b;
    layer5_outputs(3664) <= not a;
    layer5_outputs(3665) <= a xor b;
    layer5_outputs(3666) <= '1';
    layer5_outputs(3667) <= a;
    layer5_outputs(3668) <= not b;
    layer5_outputs(3669) <= not b or a;
    layer5_outputs(3670) <= a and not b;
    layer5_outputs(3671) <= a and b;
    layer5_outputs(3672) <= a and b;
    layer5_outputs(3673) <= not b or a;
    layer5_outputs(3674) <= a;
    layer5_outputs(3675) <= b;
    layer5_outputs(3676) <= b;
    layer5_outputs(3677) <= '0';
    layer5_outputs(3678) <= b;
    layer5_outputs(3679) <= not b or a;
    layer5_outputs(3680) <= b;
    layer5_outputs(3681) <= a and b;
    layer5_outputs(3682) <= not b or a;
    layer5_outputs(3683) <= a xor b;
    layer5_outputs(3684) <= not a or b;
    layer5_outputs(3685) <= a xor b;
    layer5_outputs(3686) <= not a;
    layer5_outputs(3687) <= a;
    layer5_outputs(3688) <= not b;
    layer5_outputs(3689) <= a;
    layer5_outputs(3690) <= b;
    layer5_outputs(3691) <= b;
    layer5_outputs(3692) <= a;
    layer5_outputs(3693) <= b;
    layer5_outputs(3694) <= b and not a;
    layer5_outputs(3695) <= a;
    layer5_outputs(3696) <= not b;
    layer5_outputs(3697) <= a and b;
    layer5_outputs(3698) <= '1';
    layer5_outputs(3699) <= not b or a;
    layer5_outputs(3700) <= b;
    layer5_outputs(3701) <= not (a and b);
    layer5_outputs(3702) <= not b;
    layer5_outputs(3703) <= not a;
    layer5_outputs(3704) <= not b or a;
    layer5_outputs(3705) <= not b or a;
    layer5_outputs(3706) <= not a;
    layer5_outputs(3707) <= not (a xor b);
    layer5_outputs(3708) <= not (a or b);
    layer5_outputs(3709) <= not b;
    layer5_outputs(3710) <= b;
    layer5_outputs(3711) <= not a;
    layer5_outputs(3712) <= a and not b;
    layer5_outputs(3713) <= b;
    layer5_outputs(3714) <= not b or a;
    layer5_outputs(3715) <= not (a xor b);
    layer5_outputs(3716) <= not (a or b);
    layer5_outputs(3717) <= b and not a;
    layer5_outputs(3718) <= not (a or b);
    layer5_outputs(3719) <= a xor b;
    layer5_outputs(3720) <= not (a or b);
    layer5_outputs(3721) <= '0';
    layer5_outputs(3722) <= b and not a;
    layer5_outputs(3723) <= '1';
    layer5_outputs(3724) <= not (a and b);
    layer5_outputs(3725) <= not (a and b);
    layer5_outputs(3726) <= a or b;
    layer5_outputs(3727) <= a;
    layer5_outputs(3728) <= a or b;
    layer5_outputs(3729) <= not a;
    layer5_outputs(3730) <= b;
    layer5_outputs(3731) <= b and not a;
    layer5_outputs(3732) <= '0';
    layer5_outputs(3733) <= b and not a;
    layer5_outputs(3734) <= a and not b;
    layer5_outputs(3735) <= a;
    layer5_outputs(3736) <= '1';
    layer5_outputs(3737) <= b and not a;
    layer5_outputs(3738) <= a and b;
    layer5_outputs(3739) <= not b or a;
    layer5_outputs(3740) <= b and not a;
    layer5_outputs(3741) <= not a or b;
    layer5_outputs(3742) <= not (a or b);
    layer5_outputs(3743) <= not (a xor b);
    layer5_outputs(3744) <= a;
    layer5_outputs(3745) <= not a;
    layer5_outputs(3746) <= not a;
    layer5_outputs(3747) <= a xor b;
    layer5_outputs(3748) <= a and not b;
    layer5_outputs(3749) <= not a;
    layer5_outputs(3750) <= not a;
    layer5_outputs(3751) <= not a;
    layer5_outputs(3752) <= a or b;
    layer5_outputs(3753) <= b and not a;
    layer5_outputs(3754) <= not (a xor b);
    layer5_outputs(3755) <= b;
    layer5_outputs(3756) <= not (a or b);
    layer5_outputs(3757) <= a;
    layer5_outputs(3758) <= '1';
    layer5_outputs(3759) <= not b or a;
    layer5_outputs(3760) <= not b;
    layer5_outputs(3761) <= not b;
    layer5_outputs(3762) <= not a or b;
    layer5_outputs(3763) <= not b or a;
    layer5_outputs(3764) <= not a or b;
    layer5_outputs(3765) <= not a;
    layer5_outputs(3766) <= a xor b;
    layer5_outputs(3767) <= not (a xor b);
    layer5_outputs(3768) <= a or b;
    layer5_outputs(3769) <= not b or a;
    layer5_outputs(3770) <= b;
    layer5_outputs(3771) <= a or b;
    layer5_outputs(3772) <= not (a or b);
    layer5_outputs(3773) <= b and not a;
    layer5_outputs(3774) <= not (a xor b);
    layer5_outputs(3775) <= a xor b;
    layer5_outputs(3776) <= not (a or b);
    layer5_outputs(3777) <= not b or a;
    layer5_outputs(3778) <= not a or b;
    layer5_outputs(3779) <= a;
    layer5_outputs(3780) <= not a;
    layer5_outputs(3781) <= not a or b;
    layer5_outputs(3782) <= '1';
    layer5_outputs(3783) <= a;
    layer5_outputs(3784) <= a or b;
    layer5_outputs(3785) <= a and b;
    layer5_outputs(3786) <= '1';
    layer5_outputs(3787) <= not b or a;
    layer5_outputs(3788) <= not (a or b);
    layer5_outputs(3789) <= a xor b;
    layer5_outputs(3790) <= not b or a;
    layer5_outputs(3791) <= b;
    layer5_outputs(3792) <= a and b;
    layer5_outputs(3793) <= '0';
    layer5_outputs(3794) <= a and not b;
    layer5_outputs(3795) <= a;
    layer5_outputs(3796) <= '1';
    layer5_outputs(3797) <= a and not b;
    layer5_outputs(3798) <= a or b;
    layer5_outputs(3799) <= a xor b;
    layer5_outputs(3800) <= not a;
    layer5_outputs(3801) <= not a;
    layer5_outputs(3802) <= not b;
    layer5_outputs(3803) <= '0';
    layer5_outputs(3804) <= not (a and b);
    layer5_outputs(3805) <= a xor b;
    layer5_outputs(3806) <= not (a xor b);
    layer5_outputs(3807) <= a;
    layer5_outputs(3808) <= not (a or b);
    layer5_outputs(3809) <= a or b;
    layer5_outputs(3810) <= not a;
    layer5_outputs(3811) <= b;
    layer5_outputs(3812) <= not a or b;
    layer5_outputs(3813) <= a and b;
    layer5_outputs(3814) <= b and not a;
    layer5_outputs(3815) <= not (a or b);
    layer5_outputs(3816) <= not b;
    layer5_outputs(3817) <= not (a or b);
    layer5_outputs(3818) <= b and not a;
    layer5_outputs(3819) <= b and not a;
    layer5_outputs(3820) <= b;
    layer5_outputs(3821) <= not (a and b);
    layer5_outputs(3822) <= not (a and b);
    layer5_outputs(3823) <= '1';
    layer5_outputs(3824) <= not b;
    layer5_outputs(3825) <= a;
    layer5_outputs(3826) <= '1';
    layer5_outputs(3827) <= not (a and b);
    layer5_outputs(3828) <= b and not a;
    layer5_outputs(3829) <= not (a xor b);
    layer5_outputs(3830) <= b and not a;
    layer5_outputs(3831) <= b;
    layer5_outputs(3832) <= a;
    layer5_outputs(3833) <= a;
    layer5_outputs(3834) <= a or b;
    layer5_outputs(3835) <= not a or b;
    layer5_outputs(3836) <= a;
    layer5_outputs(3837) <= a and b;
    layer5_outputs(3838) <= a or b;
    layer5_outputs(3839) <= not (a xor b);
    layer5_outputs(3840) <= b;
    layer5_outputs(3841) <= not b;
    layer5_outputs(3842) <= a or b;
    layer5_outputs(3843) <= not a;
    layer5_outputs(3844) <= not b;
    layer5_outputs(3845) <= a;
    layer5_outputs(3846) <= not b;
    layer5_outputs(3847) <= a;
    layer5_outputs(3848) <= not a or b;
    layer5_outputs(3849) <= '1';
    layer5_outputs(3850) <= not a or b;
    layer5_outputs(3851) <= not (a and b);
    layer5_outputs(3852) <= a or b;
    layer5_outputs(3853) <= a or b;
    layer5_outputs(3854) <= a or b;
    layer5_outputs(3855) <= not b;
    layer5_outputs(3856) <= b;
    layer5_outputs(3857) <= not (a and b);
    layer5_outputs(3858) <= a or b;
    layer5_outputs(3859) <= a xor b;
    layer5_outputs(3860) <= a;
    layer5_outputs(3861) <= not a or b;
    layer5_outputs(3862) <= not a or b;
    layer5_outputs(3863) <= not a;
    layer5_outputs(3864) <= not b or a;
    layer5_outputs(3865) <= not (a or b);
    layer5_outputs(3866) <= not (a or b);
    layer5_outputs(3867) <= not (a and b);
    layer5_outputs(3868) <= not (a or b);
    layer5_outputs(3869) <= not b or a;
    layer5_outputs(3870) <= a;
    layer5_outputs(3871) <= a;
    layer5_outputs(3872) <= not b or a;
    layer5_outputs(3873) <= b;
    layer5_outputs(3874) <= not b or a;
    layer5_outputs(3875) <= not a;
    layer5_outputs(3876) <= a;
    layer5_outputs(3877) <= b and not a;
    layer5_outputs(3878) <= b;
    layer5_outputs(3879) <= not a or b;
    layer5_outputs(3880) <= '0';
    layer5_outputs(3881) <= not (a or b);
    layer5_outputs(3882) <= b and not a;
    layer5_outputs(3883) <= not (a xor b);
    layer5_outputs(3884) <= not (a and b);
    layer5_outputs(3885) <= a;
    layer5_outputs(3886) <= not b;
    layer5_outputs(3887) <= b;
    layer5_outputs(3888) <= not b;
    layer5_outputs(3889) <= not a or b;
    layer5_outputs(3890) <= b;
    layer5_outputs(3891) <= '1';
    layer5_outputs(3892) <= not (a or b);
    layer5_outputs(3893) <= a xor b;
    layer5_outputs(3894) <= not (a or b);
    layer5_outputs(3895) <= not b;
    layer5_outputs(3896) <= not (a or b);
    layer5_outputs(3897) <= '1';
    layer5_outputs(3898) <= a and not b;
    layer5_outputs(3899) <= '0';
    layer5_outputs(3900) <= not b or a;
    layer5_outputs(3901) <= a or b;
    layer5_outputs(3902) <= a and not b;
    layer5_outputs(3903) <= a;
    layer5_outputs(3904) <= a;
    layer5_outputs(3905) <= a;
    layer5_outputs(3906) <= '1';
    layer5_outputs(3907) <= not b;
    layer5_outputs(3908) <= a;
    layer5_outputs(3909) <= a and not b;
    layer5_outputs(3910) <= not (a or b);
    layer5_outputs(3911) <= a and not b;
    layer5_outputs(3912) <= not b;
    layer5_outputs(3913) <= a and not b;
    layer5_outputs(3914) <= not a;
    layer5_outputs(3915) <= a xor b;
    layer5_outputs(3916) <= not b;
    layer5_outputs(3917) <= '1';
    layer5_outputs(3918) <= not b;
    layer5_outputs(3919) <= b;
    layer5_outputs(3920) <= a and b;
    layer5_outputs(3921) <= b;
    layer5_outputs(3922) <= not (a or b);
    layer5_outputs(3923) <= not b or a;
    layer5_outputs(3924) <= not a;
    layer5_outputs(3925) <= b;
    layer5_outputs(3926) <= not b;
    layer5_outputs(3927) <= not (a xor b);
    layer5_outputs(3928) <= a;
    layer5_outputs(3929) <= not b or a;
    layer5_outputs(3930) <= not (a or b);
    layer5_outputs(3931) <= not (a or b);
    layer5_outputs(3932) <= a;
    layer5_outputs(3933) <= not a or b;
    layer5_outputs(3934) <= not (a or b);
    layer5_outputs(3935) <= b;
    layer5_outputs(3936) <= not b;
    layer5_outputs(3937) <= not b or a;
    layer5_outputs(3938) <= '1';
    layer5_outputs(3939) <= not a or b;
    layer5_outputs(3940) <= b and not a;
    layer5_outputs(3941) <= a;
    layer5_outputs(3942) <= not a;
    layer5_outputs(3943) <= not (a xor b);
    layer5_outputs(3944) <= a or b;
    layer5_outputs(3945) <= not (a or b);
    layer5_outputs(3946) <= not (a and b);
    layer5_outputs(3947) <= not a;
    layer5_outputs(3948) <= not (a xor b);
    layer5_outputs(3949) <= not b or a;
    layer5_outputs(3950) <= a or b;
    layer5_outputs(3951) <= b;
    layer5_outputs(3952) <= not b or a;
    layer5_outputs(3953) <= a and b;
    layer5_outputs(3954) <= '1';
    layer5_outputs(3955) <= not b or a;
    layer5_outputs(3956) <= a;
    layer5_outputs(3957) <= a;
    layer5_outputs(3958) <= not a or b;
    layer5_outputs(3959) <= not a;
    layer5_outputs(3960) <= not a;
    layer5_outputs(3961) <= a and not b;
    layer5_outputs(3962) <= a and not b;
    layer5_outputs(3963) <= a and not b;
    layer5_outputs(3964) <= not b;
    layer5_outputs(3965) <= b;
    layer5_outputs(3966) <= not (a and b);
    layer5_outputs(3967) <= b and not a;
    layer5_outputs(3968) <= not (a or b);
    layer5_outputs(3969) <= b;
    layer5_outputs(3970) <= not (a or b);
    layer5_outputs(3971) <= b and not a;
    layer5_outputs(3972) <= a and not b;
    layer5_outputs(3973) <= not b or a;
    layer5_outputs(3974) <= not (a or b);
    layer5_outputs(3975) <= a and not b;
    layer5_outputs(3976) <= not b or a;
    layer5_outputs(3977) <= a or b;
    layer5_outputs(3978) <= not (a and b);
    layer5_outputs(3979) <= a;
    layer5_outputs(3980) <= not a;
    layer5_outputs(3981) <= b;
    layer5_outputs(3982) <= not b or a;
    layer5_outputs(3983) <= b;
    layer5_outputs(3984) <= not (a or b);
    layer5_outputs(3985) <= a;
    layer5_outputs(3986) <= not b or a;
    layer5_outputs(3987) <= not (a or b);
    layer5_outputs(3988) <= a;
    layer5_outputs(3989) <= not a;
    layer5_outputs(3990) <= not (a or b);
    layer5_outputs(3991) <= a;
    layer5_outputs(3992) <= not b;
    layer5_outputs(3993) <= a xor b;
    layer5_outputs(3994) <= a and b;
    layer5_outputs(3995) <= a;
    layer5_outputs(3996) <= b;
    layer5_outputs(3997) <= not b or a;
    layer5_outputs(3998) <= not b;
    layer5_outputs(3999) <= a xor b;
    layer5_outputs(4000) <= '0';
    layer5_outputs(4001) <= not a;
    layer5_outputs(4002) <= not b;
    layer5_outputs(4003) <= not b;
    layer5_outputs(4004) <= not a;
    layer5_outputs(4005) <= b and not a;
    layer5_outputs(4006) <= a or b;
    layer5_outputs(4007) <= not a;
    layer5_outputs(4008) <= not (a and b);
    layer5_outputs(4009) <= not b;
    layer5_outputs(4010) <= b;
    layer5_outputs(4011) <= not b;
    layer5_outputs(4012) <= not (a and b);
    layer5_outputs(4013) <= a and b;
    layer5_outputs(4014) <= b and not a;
    layer5_outputs(4015) <= not b;
    layer5_outputs(4016) <= a or b;
    layer5_outputs(4017) <= a xor b;
    layer5_outputs(4018) <= not (a xor b);
    layer5_outputs(4019) <= not b;
    layer5_outputs(4020) <= not a;
    layer5_outputs(4021) <= b;
    layer5_outputs(4022) <= a;
    layer5_outputs(4023) <= b;
    layer5_outputs(4024) <= '0';
    layer5_outputs(4025) <= not b or a;
    layer5_outputs(4026) <= a;
    layer5_outputs(4027) <= a or b;
    layer5_outputs(4028) <= a and b;
    layer5_outputs(4029) <= b;
    layer5_outputs(4030) <= not (a and b);
    layer5_outputs(4031) <= b and not a;
    layer5_outputs(4032) <= not (a and b);
    layer5_outputs(4033) <= a;
    layer5_outputs(4034) <= b;
    layer5_outputs(4035) <= not a or b;
    layer5_outputs(4036) <= a;
    layer5_outputs(4037) <= a or b;
    layer5_outputs(4038) <= a;
    layer5_outputs(4039) <= a and b;
    layer5_outputs(4040) <= not b;
    layer5_outputs(4041) <= not (a or b);
    layer5_outputs(4042) <= b;
    layer5_outputs(4043) <= '0';
    layer5_outputs(4044) <= not (a or b);
    layer5_outputs(4045) <= b and not a;
    layer5_outputs(4046) <= a;
    layer5_outputs(4047) <= not a;
    layer5_outputs(4048) <= not a or b;
    layer5_outputs(4049) <= b;
    layer5_outputs(4050) <= not a;
    layer5_outputs(4051) <= not b or a;
    layer5_outputs(4052) <= not a;
    layer5_outputs(4053) <= a and b;
    layer5_outputs(4054) <= a and b;
    layer5_outputs(4055) <= not (a and b);
    layer5_outputs(4056) <= not a;
    layer5_outputs(4057) <= not (a and b);
    layer5_outputs(4058) <= not a;
    layer5_outputs(4059) <= b;
    layer5_outputs(4060) <= b and not a;
    layer5_outputs(4061) <= '1';
    layer5_outputs(4062) <= not a;
    layer5_outputs(4063) <= b and not a;
    layer5_outputs(4064) <= not b or a;
    layer5_outputs(4065) <= b and not a;
    layer5_outputs(4066) <= b and not a;
    layer5_outputs(4067) <= a and not b;
    layer5_outputs(4068) <= b and not a;
    layer5_outputs(4069) <= not b;
    layer5_outputs(4070) <= a;
    layer5_outputs(4071) <= not a or b;
    layer5_outputs(4072) <= not a or b;
    layer5_outputs(4073) <= b;
    layer5_outputs(4074) <= '0';
    layer5_outputs(4075) <= not b or a;
    layer5_outputs(4076) <= b and not a;
    layer5_outputs(4077) <= a and b;
    layer5_outputs(4078) <= b and not a;
    layer5_outputs(4079) <= not a;
    layer5_outputs(4080) <= not a or b;
    layer5_outputs(4081) <= '1';
    layer5_outputs(4082) <= not a;
    layer5_outputs(4083) <= not b or a;
    layer5_outputs(4084) <= a;
    layer5_outputs(4085) <= not (a or b);
    layer5_outputs(4086) <= a;
    layer5_outputs(4087) <= a;
    layer5_outputs(4088) <= not a;
    layer5_outputs(4089) <= not a or b;
    layer5_outputs(4090) <= '0';
    layer5_outputs(4091) <= a or b;
    layer5_outputs(4092) <= not a;
    layer5_outputs(4093) <= '0';
    layer5_outputs(4094) <= not a;
    layer5_outputs(4095) <= b;
    layer5_outputs(4096) <= a and not b;
    layer5_outputs(4097) <= not a or b;
    layer5_outputs(4098) <= a and b;
    layer5_outputs(4099) <= not b or a;
    layer5_outputs(4100) <= '1';
    layer5_outputs(4101) <= not (a and b);
    layer5_outputs(4102) <= not (a xor b);
    layer5_outputs(4103) <= a;
    layer5_outputs(4104) <= not b or a;
    layer5_outputs(4105) <= b and not a;
    layer5_outputs(4106) <= '0';
    layer5_outputs(4107) <= not b or a;
    layer5_outputs(4108) <= a;
    layer5_outputs(4109) <= not b;
    layer5_outputs(4110) <= '0';
    layer5_outputs(4111) <= a and b;
    layer5_outputs(4112) <= not b or a;
    layer5_outputs(4113) <= not (a or b);
    layer5_outputs(4114) <= not a;
    layer5_outputs(4115) <= a;
    layer5_outputs(4116) <= b;
    layer5_outputs(4117) <= not b;
    layer5_outputs(4118) <= not (a or b);
    layer5_outputs(4119) <= not b;
    layer5_outputs(4120) <= a;
    layer5_outputs(4121) <= b;
    layer5_outputs(4122) <= '0';
    layer5_outputs(4123) <= a;
    layer5_outputs(4124) <= not b;
    layer5_outputs(4125) <= not b;
    layer5_outputs(4126) <= a xor b;
    layer5_outputs(4127) <= b;
    layer5_outputs(4128) <= '1';
    layer5_outputs(4129) <= a and not b;
    layer5_outputs(4130) <= not a;
    layer5_outputs(4131) <= b;
    layer5_outputs(4132) <= not a or b;
    layer5_outputs(4133) <= not b;
    layer5_outputs(4134) <= a xor b;
    layer5_outputs(4135) <= a;
    layer5_outputs(4136) <= not a;
    layer5_outputs(4137) <= a and not b;
    layer5_outputs(4138) <= a or b;
    layer5_outputs(4139) <= '1';
    layer5_outputs(4140) <= not b;
    layer5_outputs(4141) <= b;
    layer5_outputs(4142) <= a and not b;
    layer5_outputs(4143) <= not a;
    layer5_outputs(4144) <= not b;
    layer5_outputs(4145) <= b and not a;
    layer5_outputs(4146) <= not (a xor b);
    layer5_outputs(4147) <= b;
    layer5_outputs(4148) <= a xor b;
    layer5_outputs(4149) <= '0';
    layer5_outputs(4150) <= not (a xor b);
    layer5_outputs(4151) <= b;
    layer5_outputs(4152) <= a;
    layer5_outputs(4153) <= a and b;
    layer5_outputs(4154) <= b and not a;
    layer5_outputs(4155) <= '0';
    layer5_outputs(4156) <= a and b;
    layer5_outputs(4157) <= a and not b;
    layer5_outputs(4158) <= b;
    layer5_outputs(4159) <= a and not b;
    layer5_outputs(4160) <= not a;
    layer5_outputs(4161) <= b and not a;
    layer5_outputs(4162) <= b;
    layer5_outputs(4163) <= not b;
    layer5_outputs(4164) <= not (a or b);
    layer5_outputs(4165) <= not b;
    layer5_outputs(4166) <= '1';
    layer5_outputs(4167) <= b;
    layer5_outputs(4168) <= a or b;
    layer5_outputs(4169) <= a xor b;
    layer5_outputs(4170) <= not (a or b);
    layer5_outputs(4171) <= not b;
    layer5_outputs(4172) <= not (a and b);
    layer5_outputs(4173) <= not b or a;
    layer5_outputs(4174) <= b and not a;
    layer5_outputs(4175) <= not a or b;
    layer5_outputs(4176) <= not (a xor b);
    layer5_outputs(4177) <= not a;
    layer5_outputs(4178) <= not (a xor b);
    layer5_outputs(4179) <= not b;
    layer5_outputs(4180) <= a and not b;
    layer5_outputs(4181) <= not (a and b);
    layer5_outputs(4182) <= a or b;
    layer5_outputs(4183) <= a and b;
    layer5_outputs(4184) <= a;
    layer5_outputs(4185) <= not a;
    layer5_outputs(4186) <= not (a and b);
    layer5_outputs(4187) <= b;
    layer5_outputs(4188) <= not b;
    layer5_outputs(4189) <= not (a and b);
    layer5_outputs(4190) <= '0';
    layer5_outputs(4191) <= not a or b;
    layer5_outputs(4192) <= not a or b;
    layer5_outputs(4193) <= not b;
    layer5_outputs(4194) <= not a;
    layer5_outputs(4195) <= b and not a;
    layer5_outputs(4196) <= not b;
    layer5_outputs(4197) <= not b or a;
    layer5_outputs(4198) <= a;
    layer5_outputs(4199) <= not (a or b);
    layer5_outputs(4200) <= not b or a;
    layer5_outputs(4201) <= not (a and b);
    layer5_outputs(4202) <= a and not b;
    layer5_outputs(4203) <= a and b;
    layer5_outputs(4204) <= not (a and b);
    layer5_outputs(4205) <= not a;
    layer5_outputs(4206) <= b;
    layer5_outputs(4207) <= not b or a;
    layer5_outputs(4208) <= not b or a;
    layer5_outputs(4209) <= a and not b;
    layer5_outputs(4210) <= b;
    layer5_outputs(4211) <= not b or a;
    layer5_outputs(4212) <= a or b;
    layer5_outputs(4213) <= b and not a;
    layer5_outputs(4214) <= a and b;
    layer5_outputs(4215) <= not a or b;
    layer5_outputs(4216) <= not a or b;
    layer5_outputs(4217) <= a and not b;
    layer5_outputs(4218) <= not b;
    layer5_outputs(4219) <= a and b;
    layer5_outputs(4220) <= not b;
    layer5_outputs(4221) <= not (a or b);
    layer5_outputs(4222) <= not b or a;
    layer5_outputs(4223) <= not a;
    layer5_outputs(4224) <= not a;
    layer5_outputs(4225) <= '1';
    layer5_outputs(4226) <= a and b;
    layer5_outputs(4227) <= a;
    layer5_outputs(4228) <= a xor b;
    layer5_outputs(4229) <= a or b;
    layer5_outputs(4230) <= not b or a;
    layer5_outputs(4231) <= '1';
    layer5_outputs(4232) <= b;
    layer5_outputs(4233) <= a;
    layer5_outputs(4234) <= not (a and b);
    layer5_outputs(4235) <= a and b;
    layer5_outputs(4236) <= b;
    layer5_outputs(4237) <= a and not b;
    layer5_outputs(4238) <= not (a and b);
    layer5_outputs(4239) <= b and not a;
    layer5_outputs(4240) <= a or b;
    layer5_outputs(4241) <= not (a and b);
    layer5_outputs(4242) <= not (a xor b);
    layer5_outputs(4243) <= not b or a;
    layer5_outputs(4244) <= a xor b;
    layer5_outputs(4245) <= not a or b;
    layer5_outputs(4246) <= not b or a;
    layer5_outputs(4247) <= a xor b;
    layer5_outputs(4248) <= b and not a;
    layer5_outputs(4249) <= a and b;
    layer5_outputs(4250) <= not (a or b);
    layer5_outputs(4251) <= not a;
    layer5_outputs(4252) <= a and not b;
    layer5_outputs(4253) <= not a;
    layer5_outputs(4254) <= not a or b;
    layer5_outputs(4255) <= b and not a;
    layer5_outputs(4256) <= not b or a;
    layer5_outputs(4257) <= '1';
    layer5_outputs(4258) <= b and not a;
    layer5_outputs(4259) <= b and not a;
    layer5_outputs(4260) <= b;
    layer5_outputs(4261) <= b;
    layer5_outputs(4262) <= not a;
    layer5_outputs(4263) <= not (a or b);
    layer5_outputs(4264) <= not a;
    layer5_outputs(4265) <= a xor b;
    layer5_outputs(4266) <= not a;
    layer5_outputs(4267) <= not (a or b);
    layer5_outputs(4268) <= not b or a;
    layer5_outputs(4269) <= a;
    layer5_outputs(4270) <= not a or b;
    layer5_outputs(4271) <= not a or b;
    layer5_outputs(4272) <= not a;
    layer5_outputs(4273) <= a or b;
    layer5_outputs(4274) <= not a;
    layer5_outputs(4275) <= a and b;
    layer5_outputs(4276) <= a and not b;
    layer5_outputs(4277) <= a;
    layer5_outputs(4278) <= a and not b;
    layer5_outputs(4279) <= not a or b;
    layer5_outputs(4280) <= not b;
    layer5_outputs(4281) <= '1';
    layer5_outputs(4282) <= not (a or b);
    layer5_outputs(4283) <= not b;
    layer5_outputs(4284) <= not (a and b);
    layer5_outputs(4285) <= not b;
    layer5_outputs(4286) <= not (a xor b);
    layer5_outputs(4287) <= a xor b;
    layer5_outputs(4288) <= a;
    layer5_outputs(4289) <= a or b;
    layer5_outputs(4290) <= not a or b;
    layer5_outputs(4291) <= not b;
    layer5_outputs(4292) <= not b;
    layer5_outputs(4293) <= not (a or b);
    layer5_outputs(4294) <= a;
    layer5_outputs(4295) <= not (a xor b);
    layer5_outputs(4296) <= not b or a;
    layer5_outputs(4297) <= not (a and b);
    layer5_outputs(4298) <= not b;
    layer5_outputs(4299) <= not (a xor b);
    layer5_outputs(4300) <= not (a or b);
    layer5_outputs(4301) <= not (a and b);
    layer5_outputs(4302) <= not a;
    layer5_outputs(4303) <= not b;
    layer5_outputs(4304) <= not a;
    layer5_outputs(4305) <= '1';
    layer5_outputs(4306) <= a and b;
    layer5_outputs(4307) <= '0';
    layer5_outputs(4308) <= b;
    layer5_outputs(4309) <= '1';
    layer5_outputs(4310) <= a xor b;
    layer5_outputs(4311) <= '1';
    layer5_outputs(4312) <= b;
    layer5_outputs(4313) <= not a or b;
    layer5_outputs(4314) <= b;
    layer5_outputs(4315) <= a or b;
    layer5_outputs(4316) <= a and not b;
    layer5_outputs(4317) <= not a or b;
    layer5_outputs(4318) <= b;
    layer5_outputs(4319) <= b and not a;
    layer5_outputs(4320) <= a or b;
    layer5_outputs(4321) <= not a or b;
    layer5_outputs(4322) <= a and not b;
    layer5_outputs(4323) <= a or b;
    layer5_outputs(4324) <= a or b;
    layer5_outputs(4325) <= not a;
    layer5_outputs(4326) <= not a;
    layer5_outputs(4327) <= a xor b;
    layer5_outputs(4328) <= a;
    layer5_outputs(4329) <= not b or a;
    layer5_outputs(4330) <= b;
    layer5_outputs(4331) <= '0';
    layer5_outputs(4332) <= not a;
    layer5_outputs(4333) <= b;
    layer5_outputs(4334) <= not a;
    layer5_outputs(4335) <= not b;
    layer5_outputs(4336) <= not (a or b);
    layer5_outputs(4337) <= a and b;
    layer5_outputs(4338) <= not b;
    layer5_outputs(4339) <= a and not b;
    layer5_outputs(4340) <= not b;
    layer5_outputs(4341) <= not (a or b);
    layer5_outputs(4342) <= not (a and b);
    layer5_outputs(4343) <= not (a or b);
    layer5_outputs(4344) <= a;
    layer5_outputs(4345) <= '0';
    layer5_outputs(4346) <= not (a and b);
    layer5_outputs(4347) <= not b;
    layer5_outputs(4348) <= b and not a;
    layer5_outputs(4349) <= not a;
    layer5_outputs(4350) <= b;
    layer5_outputs(4351) <= a and b;
    layer5_outputs(4352) <= b and not a;
    layer5_outputs(4353) <= not (a and b);
    layer5_outputs(4354) <= not b or a;
    layer5_outputs(4355) <= a;
    layer5_outputs(4356) <= not a;
    layer5_outputs(4357) <= a;
    layer5_outputs(4358) <= a and not b;
    layer5_outputs(4359) <= a and not b;
    layer5_outputs(4360) <= not (a and b);
    layer5_outputs(4361) <= b;
    layer5_outputs(4362) <= not b or a;
    layer5_outputs(4363) <= a xor b;
    layer5_outputs(4364) <= b;
    layer5_outputs(4365) <= '0';
    layer5_outputs(4366) <= not (a or b);
    layer5_outputs(4367) <= not (a or b);
    layer5_outputs(4368) <= b and not a;
    layer5_outputs(4369) <= '0';
    layer5_outputs(4370) <= not b;
    layer5_outputs(4371) <= '0';
    layer5_outputs(4372) <= a or b;
    layer5_outputs(4373) <= b and not a;
    layer5_outputs(4374) <= b;
    layer5_outputs(4375) <= not b or a;
    layer5_outputs(4376) <= a;
    layer5_outputs(4377) <= not a or b;
    layer5_outputs(4378) <= not (a and b);
    layer5_outputs(4379) <= not b;
    layer5_outputs(4380) <= not b;
    layer5_outputs(4381) <= not (a and b);
    layer5_outputs(4382) <= a;
    layer5_outputs(4383) <= a;
    layer5_outputs(4384) <= a and not b;
    layer5_outputs(4385) <= a;
    layer5_outputs(4386) <= a and not b;
    layer5_outputs(4387) <= '1';
    layer5_outputs(4388) <= b;
    layer5_outputs(4389) <= '1';
    layer5_outputs(4390) <= not a;
    layer5_outputs(4391) <= not (a and b);
    layer5_outputs(4392) <= a and b;
    layer5_outputs(4393) <= not a;
    layer5_outputs(4394) <= a and not b;
    layer5_outputs(4395) <= not a;
    layer5_outputs(4396) <= not b;
    layer5_outputs(4397) <= b;
    layer5_outputs(4398) <= not b or a;
    layer5_outputs(4399) <= a and not b;
    layer5_outputs(4400) <= not b;
    layer5_outputs(4401) <= '1';
    layer5_outputs(4402) <= not a;
    layer5_outputs(4403) <= not a or b;
    layer5_outputs(4404) <= a;
    layer5_outputs(4405) <= not b;
    layer5_outputs(4406) <= b;
    layer5_outputs(4407) <= not b or a;
    layer5_outputs(4408) <= not a or b;
    layer5_outputs(4409) <= not b;
    layer5_outputs(4410) <= not b;
    layer5_outputs(4411) <= not (a xor b);
    layer5_outputs(4412) <= not b or a;
    layer5_outputs(4413) <= a or b;
    layer5_outputs(4414) <= not a;
    layer5_outputs(4415) <= a;
    layer5_outputs(4416) <= a and not b;
    layer5_outputs(4417) <= not a;
    layer5_outputs(4418) <= a and b;
    layer5_outputs(4419) <= not b or a;
    layer5_outputs(4420) <= '1';
    layer5_outputs(4421) <= not b or a;
    layer5_outputs(4422) <= a;
    layer5_outputs(4423) <= not a or b;
    layer5_outputs(4424) <= a or b;
    layer5_outputs(4425) <= not (a xor b);
    layer5_outputs(4426) <= '0';
    layer5_outputs(4427) <= b;
    layer5_outputs(4428) <= not a;
    layer5_outputs(4429) <= a;
    layer5_outputs(4430) <= not (a and b);
    layer5_outputs(4431) <= a;
    layer5_outputs(4432) <= b;
    layer5_outputs(4433) <= b and not a;
    layer5_outputs(4434) <= not b;
    layer5_outputs(4435) <= b and not a;
    layer5_outputs(4436) <= b and not a;
    layer5_outputs(4437) <= b;
    layer5_outputs(4438) <= b and not a;
    layer5_outputs(4439) <= a;
    layer5_outputs(4440) <= b;
    layer5_outputs(4441) <= b;
    layer5_outputs(4442) <= not a or b;
    layer5_outputs(4443) <= not a;
    layer5_outputs(4444) <= not b;
    layer5_outputs(4445) <= a xor b;
    layer5_outputs(4446) <= a;
    layer5_outputs(4447) <= b and not a;
    layer5_outputs(4448) <= '1';
    layer5_outputs(4449) <= a and b;
    layer5_outputs(4450) <= a or b;
    layer5_outputs(4451) <= a or b;
    layer5_outputs(4452) <= a xor b;
    layer5_outputs(4453) <= a xor b;
    layer5_outputs(4454) <= not (a and b);
    layer5_outputs(4455) <= not (a and b);
    layer5_outputs(4456) <= a or b;
    layer5_outputs(4457) <= b;
    layer5_outputs(4458) <= not (a xor b);
    layer5_outputs(4459) <= not a or b;
    layer5_outputs(4460) <= not a;
    layer5_outputs(4461) <= b;
    layer5_outputs(4462) <= not a;
    layer5_outputs(4463) <= not a;
    layer5_outputs(4464) <= not a;
    layer5_outputs(4465) <= not a;
    layer5_outputs(4466) <= a;
    layer5_outputs(4467) <= a xor b;
    layer5_outputs(4468) <= a;
    layer5_outputs(4469) <= a;
    layer5_outputs(4470) <= b;
    layer5_outputs(4471) <= not a or b;
    layer5_outputs(4472) <= a;
    layer5_outputs(4473) <= b;
    layer5_outputs(4474) <= not a or b;
    layer5_outputs(4475) <= not b or a;
    layer5_outputs(4476) <= not a;
    layer5_outputs(4477) <= not a or b;
    layer5_outputs(4478) <= b;
    layer5_outputs(4479) <= not b or a;
    layer5_outputs(4480) <= a and not b;
    layer5_outputs(4481) <= not (a or b);
    layer5_outputs(4482) <= not b or a;
    layer5_outputs(4483) <= not a;
    layer5_outputs(4484) <= not a;
    layer5_outputs(4485) <= not b;
    layer5_outputs(4486) <= a and not b;
    layer5_outputs(4487) <= not b or a;
    layer5_outputs(4488) <= a and b;
    layer5_outputs(4489) <= a;
    layer5_outputs(4490) <= not a;
    layer5_outputs(4491) <= not b;
    layer5_outputs(4492) <= not (a xor b);
    layer5_outputs(4493) <= a;
    layer5_outputs(4494) <= not a or b;
    layer5_outputs(4495) <= a or b;
    layer5_outputs(4496) <= not b or a;
    layer5_outputs(4497) <= a or b;
    layer5_outputs(4498) <= not b;
    layer5_outputs(4499) <= b;
    layer5_outputs(4500) <= not b;
    layer5_outputs(4501) <= a and b;
    layer5_outputs(4502) <= not a;
    layer5_outputs(4503) <= not a or b;
    layer5_outputs(4504) <= not a or b;
    layer5_outputs(4505) <= not b;
    layer5_outputs(4506) <= b;
    layer5_outputs(4507) <= b and not a;
    layer5_outputs(4508) <= a and not b;
    layer5_outputs(4509) <= a xor b;
    layer5_outputs(4510) <= b;
    layer5_outputs(4511) <= a and b;
    layer5_outputs(4512) <= not b;
    layer5_outputs(4513) <= '1';
    layer5_outputs(4514) <= not b or a;
    layer5_outputs(4515) <= a and not b;
    layer5_outputs(4516) <= not b;
    layer5_outputs(4517) <= not b;
    layer5_outputs(4518) <= '0';
    layer5_outputs(4519) <= a and b;
    layer5_outputs(4520) <= b;
    layer5_outputs(4521) <= not (a and b);
    layer5_outputs(4522) <= b;
    layer5_outputs(4523) <= a and not b;
    layer5_outputs(4524) <= b;
    layer5_outputs(4525) <= b and not a;
    layer5_outputs(4526) <= not b or a;
    layer5_outputs(4527) <= a xor b;
    layer5_outputs(4528) <= a;
    layer5_outputs(4529) <= a and b;
    layer5_outputs(4530) <= not (a or b);
    layer5_outputs(4531) <= not (a xor b);
    layer5_outputs(4532) <= not b or a;
    layer5_outputs(4533) <= b;
    layer5_outputs(4534) <= not (a and b);
    layer5_outputs(4535) <= b;
    layer5_outputs(4536) <= b and not a;
    layer5_outputs(4537) <= not (a or b);
    layer5_outputs(4538) <= not (a and b);
    layer5_outputs(4539) <= not (a and b);
    layer5_outputs(4540) <= a xor b;
    layer5_outputs(4541) <= a or b;
    layer5_outputs(4542) <= a or b;
    layer5_outputs(4543) <= not a;
    layer5_outputs(4544) <= not b or a;
    layer5_outputs(4545) <= a or b;
    layer5_outputs(4546) <= not (a xor b);
    layer5_outputs(4547) <= a and b;
    layer5_outputs(4548) <= not b;
    layer5_outputs(4549) <= not (a or b);
    layer5_outputs(4550) <= not (a xor b);
    layer5_outputs(4551) <= not a;
    layer5_outputs(4552) <= a;
    layer5_outputs(4553) <= not b;
    layer5_outputs(4554) <= not a;
    layer5_outputs(4555) <= a;
    layer5_outputs(4556) <= '0';
    layer5_outputs(4557) <= not b or a;
    layer5_outputs(4558) <= a and b;
    layer5_outputs(4559) <= a;
    layer5_outputs(4560) <= a and not b;
    layer5_outputs(4561) <= '0';
    layer5_outputs(4562) <= not a;
    layer5_outputs(4563) <= a or b;
    layer5_outputs(4564) <= a and b;
    layer5_outputs(4565) <= not (a or b);
    layer5_outputs(4566) <= not a or b;
    layer5_outputs(4567) <= not (a or b);
    layer5_outputs(4568) <= not b;
    layer5_outputs(4569) <= not (a or b);
    layer5_outputs(4570) <= a and b;
    layer5_outputs(4571) <= not a;
    layer5_outputs(4572) <= b;
    layer5_outputs(4573) <= a xor b;
    layer5_outputs(4574) <= not a;
    layer5_outputs(4575) <= a and not b;
    layer5_outputs(4576) <= a and not b;
    layer5_outputs(4577) <= a xor b;
    layer5_outputs(4578) <= a;
    layer5_outputs(4579) <= a;
    layer5_outputs(4580) <= not (a or b);
    layer5_outputs(4581) <= a xor b;
    layer5_outputs(4582) <= not (a xor b);
    layer5_outputs(4583) <= not a;
    layer5_outputs(4584) <= not a;
    layer5_outputs(4585) <= b;
    layer5_outputs(4586) <= not b;
    layer5_outputs(4587) <= b;
    layer5_outputs(4588) <= a or b;
    layer5_outputs(4589) <= not (a or b);
    layer5_outputs(4590) <= b;
    layer5_outputs(4591) <= not (a or b);
    layer5_outputs(4592) <= not b or a;
    layer5_outputs(4593) <= a;
    layer5_outputs(4594) <= a and not b;
    layer5_outputs(4595) <= a;
    layer5_outputs(4596) <= '0';
    layer5_outputs(4597) <= a;
    layer5_outputs(4598) <= '1';
    layer5_outputs(4599) <= '1';
    layer5_outputs(4600) <= a;
    layer5_outputs(4601) <= not b or a;
    layer5_outputs(4602) <= '0';
    layer5_outputs(4603) <= not a or b;
    layer5_outputs(4604) <= not a;
    layer5_outputs(4605) <= not a;
    layer5_outputs(4606) <= '0';
    layer5_outputs(4607) <= not b or a;
    layer5_outputs(4608) <= a xor b;
    layer5_outputs(4609) <= not a or b;
    layer5_outputs(4610) <= not a;
    layer5_outputs(4611) <= not b or a;
    layer5_outputs(4612) <= '0';
    layer5_outputs(4613) <= a or b;
    layer5_outputs(4614) <= a;
    layer5_outputs(4615) <= a and not b;
    layer5_outputs(4616) <= '0';
    layer5_outputs(4617) <= not a;
    layer5_outputs(4618) <= a;
    layer5_outputs(4619) <= a and not b;
    layer5_outputs(4620) <= not (a or b);
    layer5_outputs(4621) <= not b;
    layer5_outputs(4622) <= not b or a;
    layer5_outputs(4623) <= b;
    layer5_outputs(4624) <= a;
    layer5_outputs(4625) <= a and b;
    layer5_outputs(4626) <= b;
    layer5_outputs(4627) <= not a;
    layer5_outputs(4628) <= '1';
    layer5_outputs(4629) <= not (a xor b);
    layer5_outputs(4630) <= a or b;
    layer5_outputs(4631) <= a or b;
    layer5_outputs(4632) <= not a;
    layer5_outputs(4633) <= a and b;
    layer5_outputs(4634) <= not a;
    layer5_outputs(4635) <= not a;
    layer5_outputs(4636) <= b;
    layer5_outputs(4637) <= not b;
    layer5_outputs(4638) <= a or b;
    layer5_outputs(4639) <= b;
    layer5_outputs(4640) <= '1';
    layer5_outputs(4641) <= a and not b;
    layer5_outputs(4642) <= not a;
    layer5_outputs(4643) <= a;
    layer5_outputs(4644) <= not b or a;
    layer5_outputs(4645) <= '1';
    layer5_outputs(4646) <= not a or b;
    layer5_outputs(4647) <= a and not b;
    layer5_outputs(4648) <= a and b;
    layer5_outputs(4649) <= a;
    layer5_outputs(4650) <= a or b;
    layer5_outputs(4651) <= a and not b;
    layer5_outputs(4652) <= not a;
    layer5_outputs(4653) <= not a or b;
    layer5_outputs(4654) <= not a;
    layer5_outputs(4655) <= not a or b;
    layer5_outputs(4656) <= not a or b;
    layer5_outputs(4657) <= '1';
    layer5_outputs(4658) <= a and not b;
    layer5_outputs(4659) <= not b;
    layer5_outputs(4660) <= b;
    layer5_outputs(4661) <= a;
    layer5_outputs(4662) <= not b;
    layer5_outputs(4663) <= '0';
    layer5_outputs(4664) <= a;
    layer5_outputs(4665) <= not a;
    layer5_outputs(4666) <= not b;
    layer5_outputs(4667) <= '0';
    layer5_outputs(4668) <= a and not b;
    layer5_outputs(4669) <= b;
    layer5_outputs(4670) <= b;
    layer5_outputs(4671) <= b;
    layer5_outputs(4672) <= not (a or b);
    layer5_outputs(4673) <= not (a or b);
    layer5_outputs(4674) <= not a;
    layer5_outputs(4675) <= not (a or b);
    layer5_outputs(4676) <= b and not a;
    layer5_outputs(4677) <= a and not b;
    layer5_outputs(4678) <= not b or a;
    layer5_outputs(4679) <= b and not a;
    layer5_outputs(4680) <= not (a or b);
    layer5_outputs(4681) <= a and b;
    layer5_outputs(4682) <= '0';
    layer5_outputs(4683) <= not a;
    layer5_outputs(4684) <= a and b;
    layer5_outputs(4685) <= '0';
    layer5_outputs(4686) <= not b;
    layer5_outputs(4687) <= b;
    layer5_outputs(4688) <= '1';
    layer5_outputs(4689) <= a and b;
    layer5_outputs(4690) <= a xor b;
    layer5_outputs(4691) <= not a;
    layer5_outputs(4692) <= a and not b;
    layer5_outputs(4693) <= a or b;
    layer5_outputs(4694) <= not (a xor b);
    layer5_outputs(4695) <= not a or b;
    layer5_outputs(4696) <= a or b;
    layer5_outputs(4697) <= b;
    layer5_outputs(4698) <= '0';
    layer5_outputs(4699) <= b and not a;
    layer5_outputs(4700) <= not a;
    layer5_outputs(4701) <= not (a xor b);
    layer5_outputs(4702) <= b and not a;
    layer5_outputs(4703) <= not a;
    layer5_outputs(4704) <= a and not b;
    layer5_outputs(4705) <= b;
    layer5_outputs(4706) <= not (a and b);
    layer5_outputs(4707) <= a and not b;
    layer5_outputs(4708) <= not (a or b);
    layer5_outputs(4709) <= not a;
    layer5_outputs(4710) <= not b;
    layer5_outputs(4711) <= not a;
    layer5_outputs(4712) <= not a;
    layer5_outputs(4713) <= not a;
    layer5_outputs(4714) <= not (a and b);
    layer5_outputs(4715) <= a and b;
    layer5_outputs(4716) <= not b or a;
    layer5_outputs(4717) <= a and not b;
    layer5_outputs(4718) <= not a or b;
    layer5_outputs(4719) <= a;
    layer5_outputs(4720) <= not (a xor b);
    layer5_outputs(4721) <= a;
    layer5_outputs(4722) <= not a;
    layer5_outputs(4723) <= not b;
    layer5_outputs(4724) <= not (a or b);
    layer5_outputs(4725) <= not b;
    layer5_outputs(4726) <= not a;
    layer5_outputs(4727) <= not (a or b);
    layer5_outputs(4728) <= not (a and b);
    layer5_outputs(4729) <= not (a or b);
    layer5_outputs(4730) <= '1';
    layer5_outputs(4731) <= not (a xor b);
    layer5_outputs(4732) <= not (a or b);
    layer5_outputs(4733) <= '0';
    layer5_outputs(4734) <= a and b;
    layer5_outputs(4735) <= not (a or b);
    layer5_outputs(4736) <= a or b;
    layer5_outputs(4737) <= a and b;
    layer5_outputs(4738) <= not (a and b);
    layer5_outputs(4739) <= '1';
    layer5_outputs(4740) <= a xor b;
    layer5_outputs(4741) <= b and not a;
    layer5_outputs(4742) <= not (a xor b);
    layer5_outputs(4743) <= b;
    layer5_outputs(4744) <= a xor b;
    layer5_outputs(4745) <= a;
    layer5_outputs(4746) <= not b;
    layer5_outputs(4747) <= not a;
    layer5_outputs(4748) <= b;
    layer5_outputs(4749) <= not b;
    layer5_outputs(4750) <= not a or b;
    layer5_outputs(4751) <= '0';
    layer5_outputs(4752) <= not a;
    layer5_outputs(4753) <= not (a or b);
    layer5_outputs(4754) <= b;
    layer5_outputs(4755) <= not b or a;
    layer5_outputs(4756) <= '1';
    layer5_outputs(4757) <= '1';
    layer5_outputs(4758) <= a or b;
    layer5_outputs(4759) <= not (a and b);
    layer5_outputs(4760) <= not a;
    layer5_outputs(4761) <= not a or b;
    layer5_outputs(4762) <= a or b;
    layer5_outputs(4763) <= a or b;
    layer5_outputs(4764) <= not (a or b);
    layer5_outputs(4765) <= not (a or b);
    layer5_outputs(4766) <= not a;
    layer5_outputs(4767) <= not b;
    layer5_outputs(4768) <= not (a and b);
    layer5_outputs(4769) <= not a or b;
    layer5_outputs(4770) <= a and b;
    layer5_outputs(4771) <= not b or a;
    layer5_outputs(4772) <= not (a or b);
    layer5_outputs(4773) <= b and not a;
    layer5_outputs(4774) <= b;
    layer5_outputs(4775) <= a and b;
    layer5_outputs(4776) <= b and not a;
    layer5_outputs(4777) <= b;
    layer5_outputs(4778) <= '1';
    layer5_outputs(4779) <= '1';
    layer5_outputs(4780) <= a or b;
    layer5_outputs(4781) <= a and not b;
    layer5_outputs(4782) <= not (a and b);
    layer5_outputs(4783) <= not b or a;
    layer5_outputs(4784) <= not a or b;
    layer5_outputs(4785) <= b;
    layer5_outputs(4786) <= b and not a;
    layer5_outputs(4787) <= a and b;
    layer5_outputs(4788) <= '1';
    layer5_outputs(4789) <= a;
    layer5_outputs(4790) <= not (a xor b);
    layer5_outputs(4791) <= b;
    layer5_outputs(4792) <= a and b;
    layer5_outputs(4793) <= a and b;
    layer5_outputs(4794) <= not b or a;
    layer5_outputs(4795) <= a;
    layer5_outputs(4796) <= a;
    layer5_outputs(4797) <= not a;
    layer5_outputs(4798) <= not (a or b);
    layer5_outputs(4799) <= b;
    layer5_outputs(4800) <= a and b;
    layer5_outputs(4801) <= b;
    layer5_outputs(4802) <= not (a xor b);
    layer5_outputs(4803) <= b and not a;
    layer5_outputs(4804) <= a or b;
    layer5_outputs(4805) <= not a;
    layer5_outputs(4806) <= a;
    layer5_outputs(4807) <= a;
    layer5_outputs(4808) <= not b;
    layer5_outputs(4809) <= '1';
    layer5_outputs(4810) <= b;
    layer5_outputs(4811) <= a and b;
    layer5_outputs(4812) <= a or b;
    layer5_outputs(4813) <= a;
    layer5_outputs(4814) <= not (a and b);
    layer5_outputs(4815) <= a and not b;
    layer5_outputs(4816) <= not a;
    layer5_outputs(4817) <= a and not b;
    layer5_outputs(4818) <= a or b;
    layer5_outputs(4819) <= a or b;
    layer5_outputs(4820) <= '1';
    layer5_outputs(4821) <= b;
    layer5_outputs(4822) <= a or b;
    layer5_outputs(4823) <= not a or b;
    layer5_outputs(4824) <= a and b;
    layer5_outputs(4825) <= a and b;
    layer5_outputs(4826) <= a and b;
    layer5_outputs(4827) <= not (a or b);
    layer5_outputs(4828) <= b;
    layer5_outputs(4829) <= a;
    layer5_outputs(4830) <= not a;
    layer5_outputs(4831) <= not a or b;
    layer5_outputs(4832) <= a and b;
    layer5_outputs(4833) <= not (a and b);
    layer5_outputs(4834) <= not a;
    layer5_outputs(4835) <= not b or a;
    layer5_outputs(4836) <= not b or a;
    layer5_outputs(4837) <= not a or b;
    layer5_outputs(4838) <= not a;
    layer5_outputs(4839) <= not b;
    layer5_outputs(4840) <= not b;
    layer5_outputs(4841) <= a;
    layer5_outputs(4842) <= a and not b;
    layer5_outputs(4843) <= '0';
    layer5_outputs(4844) <= '1';
    layer5_outputs(4845) <= not b;
    layer5_outputs(4846) <= b;
    layer5_outputs(4847) <= not b or a;
    layer5_outputs(4848) <= not (a and b);
    layer5_outputs(4849) <= not (a or b);
    layer5_outputs(4850) <= b;
    layer5_outputs(4851) <= a;
    layer5_outputs(4852) <= not a or b;
    layer5_outputs(4853) <= b;
    layer5_outputs(4854) <= b;
    layer5_outputs(4855) <= not (a xor b);
    layer5_outputs(4856) <= '0';
    layer5_outputs(4857) <= a and b;
    layer5_outputs(4858) <= not a or b;
    layer5_outputs(4859) <= a;
    layer5_outputs(4860) <= not a;
    layer5_outputs(4861) <= b and not a;
    layer5_outputs(4862) <= '1';
    layer5_outputs(4863) <= not a;
    layer5_outputs(4864) <= not (a or b);
    layer5_outputs(4865) <= a and not b;
    layer5_outputs(4866) <= b;
    layer5_outputs(4867) <= a;
    layer5_outputs(4868) <= a and b;
    layer5_outputs(4869) <= not b or a;
    layer5_outputs(4870) <= not a;
    layer5_outputs(4871) <= a and b;
    layer5_outputs(4872) <= a and not b;
    layer5_outputs(4873) <= a and b;
    layer5_outputs(4874) <= a;
    layer5_outputs(4875) <= a or b;
    layer5_outputs(4876) <= a;
    layer5_outputs(4877) <= a or b;
    layer5_outputs(4878) <= a and not b;
    layer5_outputs(4879) <= not a or b;
    layer5_outputs(4880) <= a;
    layer5_outputs(4881) <= not a;
    layer5_outputs(4882) <= a xor b;
    layer5_outputs(4883) <= b;
    layer5_outputs(4884) <= a;
    layer5_outputs(4885) <= not a or b;
    layer5_outputs(4886) <= '0';
    layer5_outputs(4887) <= b and not a;
    layer5_outputs(4888) <= a or b;
    layer5_outputs(4889) <= b and not a;
    layer5_outputs(4890) <= b;
    layer5_outputs(4891) <= a and not b;
    layer5_outputs(4892) <= b and not a;
    layer5_outputs(4893) <= a or b;
    layer5_outputs(4894) <= not (a or b);
    layer5_outputs(4895) <= not a;
    layer5_outputs(4896) <= b;
    layer5_outputs(4897) <= not b or a;
    layer5_outputs(4898) <= not a;
    layer5_outputs(4899) <= not a;
    layer5_outputs(4900) <= not b;
    layer5_outputs(4901) <= b;
    layer5_outputs(4902) <= not b;
    layer5_outputs(4903) <= a and b;
    layer5_outputs(4904) <= not (a and b);
    layer5_outputs(4905) <= not (a or b);
    layer5_outputs(4906) <= not (a and b);
    layer5_outputs(4907) <= not (a xor b);
    layer5_outputs(4908) <= a and not b;
    layer5_outputs(4909) <= b;
    layer5_outputs(4910) <= a;
    layer5_outputs(4911) <= b and not a;
    layer5_outputs(4912) <= not a or b;
    layer5_outputs(4913) <= not b or a;
    layer5_outputs(4914) <= a xor b;
    layer5_outputs(4915) <= b;
    layer5_outputs(4916) <= b;
    layer5_outputs(4917) <= a and not b;
    layer5_outputs(4918) <= '0';
    layer5_outputs(4919) <= not a;
    layer5_outputs(4920) <= not a;
    layer5_outputs(4921) <= not a or b;
    layer5_outputs(4922) <= not a;
    layer5_outputs(4923) <= not b or a;
    layer5_outputs(4924) <= b;
    layer5_outputs(4925) <= not (a and b);
    layer5_outputs(4926) <= b;
    layer5_outputs(4927) <= not a or b;
    layer5_outputs(4928) <= a and b;
    layer5_outputs(4929) <= not (a and b);
    layer5_outputs(4930) <= not a or b;
    layer5_outputs(4931) <= a;
    layer5_outputs(4932) <= not b or a;
    layer5_outputs(4933) <= not a or b;
    layer5_outputs(4934) <= not b or a;
    layer5_outputs(4935) <= not b;
    layer5_outputs(4936) <= a and b;
    layer5_outputs(4937) <= a or b;
    layer5_outputs(4938) <= b and not a;
    layer5_outputs(4939) <= a xor b;
    layer5_outputs(4940) <= a;
    layer5_outputs(4941) <= not a;
    layer5_outputs(4942) <= not (a or b);
    layer5_outputs(4943) <= a and not b;
    layer5_outputs(4944) <= not (a xor b);
    layer5_outputs(4945) <= b;
    layer5_outputs(4946) <= a;
    layer5_outputs(4947) <= not a;
    layer5_outputs(4948) <= a or b;
    layer5_outputs(4949) <= not (a or b);
    layer5_outputs(4950) <= a;
    layer5_outputs(4951) <= not a or b;
    layer5_outputs(4952) <= b and not a;
    layer5_outputs(4953) <= a and b;
    layer5_outputs(4954) <= not b;
    layer5_outputs(4955) <= not b;
    layer5_outputs(4956) <= a or b;
    layer5_outputs(4957) <= not b;
    layer5_outputs(4958) <= a;
    layer5_outputs(4959) <= not (a or b);
    layer5_outputs(4960) <= not a;
    layer5_outputs(4961) <= a xor b;
    layer5_outputs(4962) <= not b;
    layer5_outputs(4963) <= '1';
    layer5_outputs(4964) <= not (a xor b);
    layer5_outputs(4965) <= not a;
    layer5_outputs(4966) <= not b or a;
    layer5_outputs(4967) <= a and b;
    layer5_outputs(4968) <= a and not b;
    layer5_outputs(4969) <= b and not a;
    layer5_outputs(4970) <= not b;
    layer5_outputs(4971) <= not b;
    layer5_outputs(4972) <= a and not b;
    layer5_outputs(4973) <= not (a or b);
    layer5_outputs(4974) <= not a;
    layer5_outputs(4975) <= a and b;
    layer5_outputs(4976) <= not a;
    layer5_outputs(4977) <= b;
    layer5_outputs(4978) <= not (a or b);
    layer5_outputs(4979) <= a and not b;
    layer5_outputs(4980) <= b and not a;
    layer5_outputs(4981) <= b and not a;
    layer5_outputs(4982) <= a or b;
    layer5_outputs(4983) <= a;
    layer5_outputs(4984) <= a and not b;
    layer5_outputs(4985) <= b;
    layer5_outputs(4986) <= not a or b;
    layer5_outputs(4987) <= '1';
    layer5_outputs(4988) <= b and not a;
    layer5_outputs(4989) <= not b;
    layer5_outputs(4990) <= '1';
    layer5_outputs(4991) <= b;
    layer5_outputs(4992) <= not (a and b);
    layer5_outputs(4993) <= a and not b;
    layer5_outputs(4994) <= not (a and b);
    layer5_outputs(4995) <= a;
    layer5_outputs(4996) <= a;
    layer5_outputs(4997) <= a;
    layer5_outputs(4998) <= not (a and b);
    layer5_outputs(4999) <= not a;
    layer5_outputs(5000) <= not (a or b);
    layer5_outputs(5001) <= b;
    layer5_outputs(5002) <= a and not b;
    layer5_outputs(5003) <= a and b;
    layer5_outputs(5004) <= a and b;
    layer5_outputs(5005) <= not b;
    layer5_outputs(5006) <= b;
    layer5_outputs(5007) <= a and not b;
    layer5_outputs(5008) <= b and not a;
    layer5_outputs(5009) <= a and b;
    layer5_outputs(5010) <= '0';
    layer5_outputs(5011) <= not b;
    layer5_outputs(5012) <= '1';
    layer5_outputs(5013) <= b and not a;
    layer5_outputs(5014) <= b and not a;
    layer5_outputs(5015) <= a and b;
    layer5_outputs(5016) <= not (a and b);
    layer5_outputs(5017) <= a;
    layer5_outputs(5018) <= not b;
    layer5_outputs(5019) <= a or b;
    layer5_outputs(5020) <= a and b;
    layer5_outputs(5021) <= a and not b;
    layer5_outputs(5022) <= not (a or b);
    layer5_outputs(5023) <= a;
    layer5_outputs(5024) <= a or b;
    layer5_outputs(5025) <= a and b;
    layer5_outputs(5026) <= not b or a;
    layer5_outputs(5027) <= a and not b;
    layer5_outputs(5028) <= not b;
    layer5_outputs(5029) <= not b;
    layer5_outputs(5030) <= a and not b;
    layer5_outputs(5031) <= not (a or b);
    layer5_outputs(5032) <= not a or b;
    layer5_outputs(5033) <= '1';
    layer5_outputs(5034) <= '0';
    layer5_outputs(5035) <= not b;
    layer5_outputs(5036) <= a;
    layer5_outputs(5037) <= not b;
    layer5_outputs(5038) <= not a;
    layer5_outputs(5039) <= not b or a;
    layer5_outputs(5040) <= b;
    layer5_outputs(5041) <= not a or b;
    layer5_outputs(5042) <= not a;
    layer5_outputs(5043) <= a and b;
    layer5_outputs(5044) <= not (a xor b);
    layer5_outputs(5045) <= a and b;
    layer5_outputs(5046) <= not a;
    layer5_outputs(5047) <= not a;
    layer5_outputs(5048) <= a or b;
    layer5_outputs(5049) <= not b or a;
    layer5_outputs(5050) <= not b;
    layer5_outputs(5051) <= a and not b;
    layer5_outputs(5052) <= not a;
    layer5_outputs(5053) <= a;
    layer5_outputs(5054) <= not b or a;
    layer5_outputs(5055) <= a;
    layer5_outputs(5056) <= a and not b;
    layer5_outputs(5057) <= b;
    layer5_outputs(5058) <= a;
    layer5_outputs(5059) <= not b;
    layer5_outputs(5060) <= '0';
    layer5_outputs(5061) <= a and not b;
    layer5_outputs(5062) <= b;
    layer5_outputs(5063) <= a and not b;
    layer5_outputs(5064) <= '1';
    layer5_outputs(5065) <= a xor b;
    layer5_outputs(5066) <= not b or a;
    layer5_outputs(5067) <= '1';
    layer5_outputs(5068) <= a or b;
    layer5_outputs(5069) <= a xor b;
    layer5_outputs(5070) <= not b or a;
    layer5_outputs(5071) <= a;
    layer5_outputs(5072) <= a and not b;
    layer5_outputs(5073) <= a and b;
    layer5_outputs(5074) <= '0';
    layer5_outputs(5075) <= a xor b;
    layer5_outputs(5076) <= a xor b;
    layer5_outputs(5077) <= not b;
    layer5_outputs(5078) <= a;
    layer5_outputs(5079) <= '1';
    layer5_outputs(5080) <= b;
    layer5_outputs(5081) <= not b or a;
    layer5_outputs(5082) <= not a or b;
    layer5_outputs(5083) <= '1';
    layer5_outputs(5084) <= not b or a;
    layer5_outputs(5085) <= not b;
    layer5_outputs(5086) <= not a;
    layer5_outputs(5087) <= b;
    layer5_outputs(5088) <= a;
    layer5_outputs(5089) <= a or b;
    layer5_outputs(5090) <= a and b;
    layer5_outputs(5091) <= not (a or b);
    layer5_outputs(5092) <= not a;
    layer5_outputs(5093) <= b and not a;
    layer5_outputs(5094) <= a or b;
    layer5_outputs(5095) <= b;
    layer5_outputs(5096) <= not (a or b);
    layer5_outputs(5097) <= not b;
    layer5_outputs(5098) <= not a;
    layer5_outputs(5099) <= not (a and b);
    layer5_outputs(5100) <= not a;
    layer5_outputs(5101) <= not a or b;
    layer5_outputs(5102) <= a;
    layer5_outputs(5103) <= a or b;
    layer5_outputs(5104) <= b;
    layer5_outputs(5105) <= not (a and b);
    layer5_outputs(5106) <= a;
    layer5_outputs(5107) <= not (a xor b);
    layer5_outputs(5108) <= not b;
    layer5_outputs(5109) <= not (a or b);
    layer5_outputs(5110) <= not (a and b);
    layer5_outputs(5111) <= '1';
    layer5_outputs(5112) <= not b;
    layer5_outputs(5113) <= a or b;
    layer5_outputs(5114) <= a and not b;
    layer5_outputs(5115) <= b;
    layer5_outputs(5116) <= not b or a;
    layer5_outputs(5117) <= a;
    layer5_outputs(5118) <= a;
    layer5_outputs(5119) <= a and not b;
    layer6_outputs(0) <= a and not b;
    layer6_outputs(1) <= not (a or b);
    layer6_outputs(2) <= a and b;
    layer6_outputs(3) <= b and not a;
    layer6_outputs(4) <= not a;
    layer6_outputs(5) <= not (a and b);
    layer6_outputs(6) <= not b or a;
    layer6_outputs(7) <= a and b;
    layer6_outputs(8) <= not a or b;
    layer6_outputs(9) <= not (a or b);
    layer6_outputs(10) <= b;
    layer6_outputs(11) <= not (a or b);
    layer6_outputs(12) <= not (a xor b);
    layer6_outputs(13) <= b and not a;
    layer6_outputs(14) <= a xor b;
    layer6_outputs(15) <= not a;
    layer6_outputs(16) <= not (a xor b);
    layer6_outputs(17) <= not b;
    layer6_outputs(18) <= '1';
    layer6_outputs(19) <= not (a or b);
    layer6_outputs(20) <= not b;
    layer6_outputs(21) <= not (a or b);
    layer6_outputs(22) <= b and not a;
    layer6_outputs(23) <= not (a or b);
    layer6_outputs(24) <= a and not b;
    layer6_outputs(25) <= a xor b;
    layer6_outputs(26) <= b;
    layer6_outputs(27) <= '0';
    layer6_outputs(28) <= b;
    layer6_outputs(29) <= b and not a;
    layer6_outputs(30) <= not (a and b);
    layer6_outputs(31) <= b;
    layer6_outputs(32) <= a and b;
    layer6_outputs(33) <= '0';
    layer6_outputs(34) <= a or b;
    layer6_outputs(35) <= not b or a;
    layer6_outputs(36) <= b and not a;
    layer6_outputs(37) <= not a;
    layer6_outputs(38) <= a;
    layer6_outputs(39) <= not a;
    layer6_outputs(40) <= a;
    layer6_outputs(41) <= not b;
    layer6_outputs(42) <= not a or b;
    layer6_outputs(43) <= not b;
    layer6_outputs(44) <= not b;
    layer6_outputs(45) <= not b;
    layer6_outputs(46) <= not b;
    layer6_outputs(47) <= not a;
    layer6_outputs(48) <= not b;
    layer6_outputs(49) <= not (a and b);
    layer6_outputs(50) <= a and not b;
    layer6_outputs(51) <= a xor b;
    layer6_outputs(52) <= '0';
    layer6_outputs(53) <= a and b;
    layer6_outputs(54) <= b;
    layer6_outputs(55) <= a or b;
    layer6_outputs(56) <= b;
    layer6_outputs(57) <= not (a or b);
    layer6_outputs(58) <= not b;
    layer6_outputs(59) <= a and b;
    layer6_outputs(60) <= not (a and b);
    layer6_outputs(61) <= not (a or b);
    layer6_outputs(62) <= not (a or b);
    layer6_outputs(63) <= not (a and b);
    layer6_outputs(64) <= b;
    layer6_outputs(65) <= b;
    layer6_outputs(66) <= b and not a;
    layer6_outputs(67) <= not (a or b);
    layer6_outputs(68) <= b and not a;
    layer6_outputs(69) <= b;
    layer6_outputs(70) <= b and not a;
    layer6_outputs(71) <= not b;
    layer6_outputs(72) <= a and not b;
    layer6_outputs(73) <= a or b;
    layer6_outputs(74) <= '0';
    layer6_outputs(75) <= not a;
    layer6_outputs(76) <= not b or a;
    layer6_outputs(77) <= a and b;
    layer6_outputs(78) <= b;
    layer6_outputs(79) <= not a;
    layer6_outputs(80) <= a or b;
    layer6_outputs(81) <= not a;
    layer6_outputs(82) <= not (a or b);
    layer6_outputs(83) <= not a;
    layer6_outputs(84) <= not b;
    layer6_outputs(85) <= not b;
    layer6_outputs(86) <= not b;
    layer6_outputs(87) <= not a or b;
    layer6_outputs(88) <= b;
    layer6_outputs(89) <= not b;
    layer6_outputs(90) <= a and b;
    layer6_outputs(91) <= not (a xor b);
    layer6_outputs(92) <= a or b;
    layer6_outputs(93) <= a;
    layer6_outputs(94) <= b;
    layer6_outputs(95) <= not b;
    layer6_outputs(96) <= not b or a;
    layer6_outputs(97) <= b;
    layer6_outputs(98) <= not b;
    layer6_outputs(99) <= not a;
    layer6_outputs(100) <= b;
    layer6_outputs(101) <= not (a and b);
    layer6_outputs(102) <= a or b;
    layer6_outputs(103) <= not b;
    layer6_outputs(104) <= a xor b;
    layer6_outputs(105) <= not b or a;
    layer6_outputs(106) <= a xor b;
    layer6_outputs(107) <= not (a and b);
    layer6_outputs(108) <= a;
    layer6_outputs(109) <= not b;
    layer6_outputs(110) <= a or b;
    layer6_outputs(111) <= b;
    layer6_outputs(112) <= not b or a;
    layer6_outputs(113) <= b;
    layer6_outputs(114) <= b and not a;
    layer6_outputs(115) <= a;
    layer6_outputs(116) <= not b;
    layer6_outputs(117) <= a and not b;
    layer6_outputs(118) <= not a or b;
    layer6_outputs(119) <= '0';
    layer6_outputs(120) <= a or b;
    layer6_outputs(121) <= not a;
    layer6_outputs(122) <= not a;
    layer6_outputs(123) <= a and not b;
    layer6_outputs(124) <= not (a xor b);
    layer6_outputs(125) <= a;
    layer6_outputs(126) <= not (a or b);
    layer6_outputs(127) <= not a;
    layer6_outputs(128) <= a xor b;
    layer6_outputs(129) <= a;
    layer6_outputs(130) <= not b;
    layer6_outputs(131) <= a or b;
    layer6_outputs(132) <= not a;
    layer6_outputs(133) <= a;
    layer6_outputs(134) <= a and not b;
    layer6_outputs(135) <= not a or b;
    layer6_outputs(136) <= not a or b;
    layer6_outputs(137) <= not b;
    layer6_outputs(138) <= not b;
    layer6_outputs(139) <= not a or b;
    layer6_outputs(140) <= not a;
    layer6_outputs(141) <= a and not b;
    layer6_outputs(142) <= not a;
    layer6_outputs(143) <= not b or a;
    layer6_outputs(144) <= '1';
    layer6_outputs(145) <= b and not a;
    layer6_outputs(146) <= not b;
    layer6_outputs(147) <= a and b;
    layer6_outputs(148) <= a and not b;
    layer6_outputs(149) <= a xor b;
    layer6_outputs(150) <= a;
    layer6_outputs(151) <= not a;
    layer6_outputs(152) <= not b;
    layer6_outputs(153) <= a;
    layer6_outputs(154) <= not b or a;
    layer6_outputs(155) <= not b;
    layer6_outputs(156) <= a;
    layer6_outputs(157) <= a xor b;
    layer6_outputs(158) <= a;
    layer6_outputs(159) <= a and not b;
    layer6_outputs(160) <= b;
    layer6_outputs(161) <= not a or b;
    layer6_outputs(162) <= not b;
    layer6_outputs(163) <= not (a or b);
    layer6_outputs(164) <= not a or b;
    layer6_outputs(165) <= a;
    layer6_outputs(166) <= b;
    layer6_outputs(167) <= not a;
    layer6_outputs(168) <= a;
    layer6_outputs(169) <= a and not b;
    layer6_outputs(170) <= b;
    layer6_outputs(171) <= a;
    layer6_outputs(172) <= not b or a;
    layer6_outputs(173) <= a and not b;
    layer6_outputs(174) <= not (a xor b);
    layer6_outputs(175) <= not (a or b);
    layer6_outputs(176) <= a and not b;
    layer6_outputs(177) <= b;
    layer6_outputs(178) <= a or b;
    layer6_outputs(179) <= a or b;
    layer6_outputs(180) <= b;
    layer6_outputs(181) <= not (a or b);
    layer6_outputs(182) <= not b;
    layer6_outputs(183) <= not b or a;
    layer6_outputs(184) <= not b or a;
    layer6_outputs(185) <= not (a or b);
    layer6_outputs(186) <= not a or b;
    layer6_outputs(187) <= not (a and b);
    layer6_outputs(188) <= a and b;
    layer6_outputs(189) <= a and b;
    layer6_outputs(190) <= not b;
    layer6_outputs(191) <= '1';
    layer6_outputs(192) <= not a;
    layer6_outputs(193) <= not (a and b);
    layer6_outputs(194) <= b;
    layer6_outputs(195) <= a or b;
    layer6_outputs(196) <= not a or b;
    layer6_outputs(197) <= a or b;
    layer6_outputs(198) <= a;
    layer6_outputs(199) <= not a or b;
    layer6_outputs(200) <= not a;
    layer6_outputs(201) <= a and b;
    layer6_outputs(202) <= a xor b;
    layer6_outputs(203) <= not a or b;
    layer6_outputs(204) <= a or b;
    layer6_outputs(205) <= not b or a;
    layer6_outputs(206) <= not a;
    layer6_outputs(207) <= b;
    layer6_outputs(208) <= b;
    layer6_outputs(209) <= b;
    layer6_outputs(210) <= not a or b;
    layer6_outputs(211) <= a and not b;
    layer6_outputs(212) <= not (a xor b);
    layer6_outputs(213) <= a and b;
    layer6_outputs(214) <= not b;
    layer6_outputs(215) <= not b;
    layer6_outputs(216) <= a or b;
    layer6_outputs(217) <= a;
    layer6_outputs(218) <= a or b;
    layer6_outputs(219) <= a and not b;
    layer6_outputs(220) <= not b or a;
    layer6_outputs(221) <= not (a or b);
    layer6_outputs(222) <= not (a or b);
    layer6_outputs(223) <= not a or b;
    layer6_outputs(224) <= not b;
    layer6_outputs(225) <= not (a xor b);
    layer6_outputs(226) <= a;
    layer6_outputs(227) <= a and b;
    layer6_outputs(228) <= a or b;
    layer6_outputs(229) <= a and b;
    layer6_outputs(230) <= b;
    layer6_outputs(231) <= not a;
    layer6_outputs(232) <= a and b;
    layer6_outputs(233) <= b;
    layer6_outputs(234) <= a;
    layer6_outputs(235) <= not b;
    layer6_outputs(236) <= b and not a;
    layer6_outputs(237) <= a;
    layer6_outputs(238) <= not b;
    layer6_outputs(239) <= a and b;
    layer6_outputs(240) <= not a;
    layer6_outputs(241) <= not b or a;
    layer6_outputs(242) <= b and not a;
    layer6_outputs(243) <= a and not b;
    layer6_outputs(244) <= a or b;
    layer6_outputs(245) <= a;
    layer6_outputs(246) <= not b;
    layer6_outputs(247) <= a;
    layer6_outputs(248) <= not b;
    layer6_outputs(249) <= not b;
    layer6_outputs(250) <= a and not b;
    layer6_outputs(251) <= not b;
    layer6_outputs(252) <= not b;
    layer6_outputs(253) <= not (a and b);
    layer6_outputs(254) <= b;
    layer6_outputs(255) <= not (a and b);
    layer6_outputs(256) <= not (a and b);
    layer6_outputs(257) <= b;
    layer6_outputs(258) <= a or b;
    layer6_outputs(259) <= not b;
    layer6_outputs(260) <= not b;
    layer6_outputs(261) <= not b or a;
    layer6_outputs(262) <= a and b;
    layer6_outputs(263) <= b;
    layer6_outputs(264) <= a and not b;
    layer6_outputs(265) <= a and b;
    layer6_outputs(266) <= b;
    layer6_outputs(267) <= not b;
    layer6_outputs(268) <= not b or a;
    layer6_outputs(269) <= not b;
    layer6_outputs(270) <= a;
    layer6_outputs(271) <= a;
    layer6_outputs(272) <= not b or a;
    layer6_outputs(273) <= not a;
    layer6_outputs(274) <= a xor b;
    layer6_outputs(275) <= not b;
    layer6_outputs(276) <= not (a or b);
    layer6_outputs(277) <= not (a xor b);
    layer6_outputs(278) <= not (a or b);
    layer6_outputs(279) <= not (a xor b);
    layer6_outputs(280) <= not b;
    layer6_outputs(281) <= b and not a;
    layer6_outputs(282) <= not b or a;
    layer6_outputs(283) <= a or b;
    layer6_outputs(284) <= not (a and b);
    layer6_outputs(285) <= not a or b;
    layer6_outputs(286) <= a and not b;
    layer6_outputs(287) <= a xor b;
    layer6_outputs(288) <= a and not b;
    layer6_outputs(289) <= a;
    layer6_outputs(290) <= a or b;
    layer6_outputs(291) <= b;
    layer6_outputs(292) <= not b or a;
    layer6_outputs(293) <= not b or a;
    layer6_outputs(294) <= a or b;
    layer6_outputs(295) <= b;
    layer6_outputs(296) <= '1';
    layer6_outputs(297) <= a xor b;
    layer6_outputs(298) <= '0';
    layer6_outputs(299) <= not b or a;
    layer6_outputs(300) <= b and not a;
    layer6_outputs(301) <= not a;
    layer6_outputs(302) <= '1';
    layer6_outputs(303) <= not b;
    layer6_outputs(304) <= not a;
    layer6_outputs(305) <= not (a or b);
    layer6_outputs(306) <= not a;
    layer6_outputs(307) <= not a;
    layer6_outputs(308) <= a and not b;
    layer6_outputs(309) <= a and not b;
    layer6_outputs(310) <= a and b;
    layer6_outputs(311) <= a;
    layer6_outputs(312) <= a or b;
    layer6_outputs(313) <= a and not b;
    layer6_outputs(314) <= b;
    layer6_outputs(315) <= a and b;
    layer6_outputs(316) <= not (a xor b);
    layer6_outputs(317) <= not b or a;
    layer6_outputs(318) <= not (a xor b);
    layer6_outputs(319) <= not b or a;
    layer6_outputs(320) <= b;
    layer6_outputs(321) <= a;
    layer6_outputs(322) <= a xor b;
    layer6_outputs(323) <= not (a or b);
    layer6_outputs(324) <= a;
    layer6_outputs(325) <= b;
    layer6_outputs(326) <= not b;
    layer6_outputs(327) <= b and not a;
    layer6_outputs(328) <= not b or a;
    layer6_outputs(329) <= a and not b;
    layer6_outputs(330) <= not a or b;
    layer6_outputs(331) <= a or b;
    layer6_outputs(332) <= '1';
    layer6_outputs(333) <= not b;
    layer6_outputs(334) <= b;
    layer6_outputs(335) <= a;
    layer6_outputs(336) <= not a;
    layer6_outputs(337) <= not (a or b);
    layer6_outputs(338) <= '0';
    layer6_outputs(339) <= a;
    layer6_outputs(340) <= b;
    layer6_outputs(341) <= not b or a;
    layer6_outputs(342) <= not (a xor b);
    layer6_outputs(343) <= not b;
    layer6_outputs(344) <= b;
    layer6_outputs(345) <= a or b;
    layer6_outputs(346) <= b and not a;
    layer6_outputs(347) <= a xor b;
    layer6_outputs(348) <= a or b;
    layer6_outputs(349) <= a and not b;
    layer6_outputs(350) <= a;
    layer6_outputs(351) <= not a;
    layer6_outputs(352) <= not a;
    layer6_outputs(353) <= b;
    layer6_outputs(354) <= a or b;
    layer6_outputs(355) <= not a;
    layer6_outputs(356) <= not b;
    layer6_outputs(357) <= not a or b;
    layer6_outputs(358) <= not (a xor b);
    layer6_outputs(359) <= a;
    layer6_outputs(360) <= not a or b;
    layer6_outputs(361) <= b and not a;
    layer6_outputs(362) <= '1';
    layer6_outputs(363) <= not b or a;
    layer6_outputs(364) <= not a or b;
    layer6_outputs(365) <= a or b;
    layer6_outputs(366) <= not a or b;
    layer6_outputs(367) <= a or b;
    layer6_outputs(368) <= b;
    layer6_outputs(369) <= a and b;
    layer6_outputs(370) <= b;
    layer6_outputs(371) <= not a;
    layer6_outputs(372) <= not (a xor b);
    layer6_outputs(373) <= not a or b;
    layer6_outputs(374) <= not (a and b);
    layer6_outputs(375) <= a or b;
    layer6_outputs(376) <= not (a and b);
    layer6_outputs(377) <= a and b;
    layer6_outputs(378) <= a;
    layer6_outputs(379) <= not b or a;
    layer6_outputs(380) <= b;
    layer6_outputs(381) <= not b;
    layer6_outputs(382) <= b;
    layer6_outputs(383) <= not b;
    layer6_outputs(384) <= '0';
    layer6_outputs(385) <= a;
    layer6_outputs(386) <= not (a and b);
    layer6_outputs(387) <= b;
    layer6_outputs(388) <= a;
    layer6_outputs(389) <= not a or b;
    layer6_outputs(390) <= not a;
    layer6_outputs(391) <= not (a or b);
    layer6_outputs(392) <= not (a xor b);
    layer6_outputs(393) <= a;
    layer6_outputs(394) <= a or b;
    layer6_outputs(395) <= not b;
    layer6_outputs(396) <= a or b;
    layer6_outputs(397) <= not a;
    layer6_outputs(398) <= not (a and b);
    layer6_outputs(399) <= not b;
    layer6_outputs(400) <= not a;
    layer6_outputs(401) <= b and not a;
    layer6_outputs(402) <= a or b;
    layer6_outputs(403) <= a;
    layer6_outputs(404) <= b;
    layer6_outputs(405) <= not a;
    layer6_outputs(406) <= a and b;
    layer6_outputs(407) <= not b;
    layer6_outputs(408) <= b and not a;
    layer6_outputs(409) <= a and not b;
    layer6_outputs(410) <= a;
    layer6_outputs(411) <= not a or b;
    layer6_outputs(412) <= not (a or b);
    layer6_outputs(413) <= a or b;
    layer6_outputs(414) <= not a;
    layer6_outputs(415) <= not (a and b);
    layer6_outputs(416) <= not (a or b);
    layer6_outputs(417) <= not a;
    layer6_outputs(418) <= b and not a;
    layer6_outputs(419) <= not b or a;
    layer6_outputs(420) <= not b or a;
    layer6_outputs(421) <= not a;
    layer6_outputs(422) <= a xor b;
    layer6_outputs(423) <= not a;
    layer6_outputs(424) <= '0';
    layer6_outputs(425) <= a and not b;
    layer6_outputs(426) <= a and b;
    layer6_outputs(427) <= not b;
    layer6_outputs(428) <= a;
    layer6_outputs(429) <= not b;
    layer6_outputs(430) <= not b or a;
    layer6_outputs(431) <= b and not a;
    layer6_outputs(432) <= b;
    layer6_outputs(433) <= not a;
    layer6_outputs(434) <= not (a and b);
    layer6_outputs(435) <= not (a xor b);
    layer6_outputs(436) <= not b or a;
    layer6_outputs(437) <= not (a or b);
    layer6_outputs(438) <= a xor b;
    layer6_outputs(439) <= not a;
    layer6_outputs(440) <= not a;
    layer6_outputs(441) <= not a or b;
    layer6_outputs(442) <= not (a and b);
    layer6_outputs(443) <= not (a or b);
    layer6_outputs(444) <= not b or a;
    layer6_outputs(445) <= not b;
    layer6_outputs(446) <= not (a or b);
    layer6_outputs(447) <= b;
    layer6_outputs(448) <= not b;
    layer6_outputs(449) <= a;
    layer6_outputs(450) <= not (a or b);
    layer6_outputs(451) <= not b or a;
    layer6_outputs(452) <= b;
    layer6_outputs(453) <= a and not b;
    layer6_outputs(454) <= b;
    layer6_outputs(455) <= not b;
    layer6_outputs(456) <= not a;
    layer6_outputs(457) <= not a or b;
    layer6_outputs(458) <= not b;
    layer6_outputs(459) <= b;
    layer6_outputs(460) <= not (a xor b);
    layer6_outputs(461) <= not b;
    layer6_outputs(462) <= not (a xor b);
    layer6_outputs(463) <= a;
    layer6_outputs(464) <= a xor b;
    layer6_outputs(465) <= not a or b;
    layer6_outputs(466) <= b;
    layer6_outputs(467) <= not a or b;
    layer6_outputs(468) <= a or b;
    layer6_outputs(469) <= a;
    layer6_outputs(470) <= not (a or b);
    layer6_outputs(471) <= a and b;
    layer6_outputs(472) <= a;
    layer6_outputs(473) <= not a;
    layer6_outputs(474) <= not (a xor b);
    layer6_outputs(475) <= not (a or b);
    layer6_outputs(476) <= a and b;
    layer6_outputs(477) <= not (a and b);
    layer6_outputs(478) <= not a;
    layer6_outputs(479) <= not a;
    layer6_outputs(480) <= b;
    layer6_outputs(481) <= not a;
    layer6_outputs(482) <= a and b;
    layer6_outputs(483) <= b;
    layer6_outputs(484) <= b and not a;
    layer6_outputs(485) <= not b;
    layer6_outputs(486) <= a;
    layer6_outputs(487) <= b;
    layer6_outputs(488) <= a;
    layer6_outputs(489) <= not a or b;
    layer6_outputs(490) <= not b;
    layer6_outputs(491) <= b and not a;
    layer6_outputs(492) <= '1';
    layer6_outputs(493) <= not a;
    layer6_outputs(494) <= not (a xor b);
    layer6_outputs(495) <= b and not a;
    layer6_outputs(496) <= a xor b;
    layer6_outputs(497) <= not a;
    layer6_outputs(498) <= '1';
    layer6_outputs(499) <= b;
    layer6_outputs(500) <= not (a or b);
    layer6_outputs(501) <= not a or b;
    layer6_outputs(502) <= not b;
    layer6_outputs(503) <= not a;
    layer6_outputs(504) <= not a;
    layer6_outputs(505) <= b and not a;
    layer6_outputs(506) <= a and not b;
    layer6_outputs(507) <= not b;
    layer6_outputs(508) <= b and not a;
    layer6_outputs(509) <= b;
    layer6_outputs(510) <= a;
    layer6_outputs(511) <= not (a and b);
    layer6_outputs(512) <= a xor b;
    layer6_outputs(513) <= not (a or b);
    layer6_outputs(514) <= b;
    layer6_outputs(515) <= not (a or b);
    layer6_outputs(516) <= not a;
    layer6_outputs(517) <= not b or a;
    layer6_outputs(518) <= not a;
    layer6_outputs(519) <= a;
    layer6_outputs(520) <= b;
    layer6_outputs(521) <= not b;
    layer6_outputs(522) <= not (a xor b);
    layer6_outputs(523) <= a xor b;
    layer6_outputs(524) <= not a;
    layer6_outputs(525) <= a;
    layer6_outputs(526) <= a and b;
    layer6_outputs(527) <= not (a and b);
    layer6_outputs(528) <= a or b;
    layer6_outputs(529) <= not a or b;
    layer6_outputs(530) <= not b;
    layer6_outputs(531) <= not a or b;
    layer6_outputs(532) <= not a;
    layer6_outputs(533) <= a and b;
    layer6_outputs(534) <= not (a and b);
    layer6_outputs(535) <= a or b;
    layer6_outputs(536) <= not (a xor b);
    layer6_outputs(537) <= a;
    layer6_outputs(538) <= not (a or b);
    layer6_outputs(539) <= not b or a;
    layer6_outputs(540) <= not (a and b);
    layer6_outputs(541) <= not (a and b);
    layer6_outputs(542) <= a;
    layer6_outputs(543) <= b;
    layer6_outputs(544) <= not (a and b);
    layer6_outputs(545) <= a;
    layer6_outputs(546) <= b and not a;
    layer6_outputs(547) <= not (a or b);
    layer6_outputs(548) <= b;
    layer6_outputs(549) <= a;
    layer6_outputs(550) <= not a or b;
    layer6_outputs(551) <= b;
    layer6_outputs(552) <= not b;
    layer6_outputs(553) <= a and not b;
    layer6_outputs(554) <= not b;
    layer6_outputs(555) <= not a;
    layer6_outputs(556) <= b;
    layer6_outputs(557) <= a xor b;
    layer6_outputs(558) <= a and b;
    layer6_outputs(559) <= b;
    layer6_outputs(560) <= not b or a;
    layer6_outputs(561) <= not (a or b);
    layer6_outputs(562) <= not (a and b);
    layer6_outputs(563) <= not b;
    layer6_outputs(564) <= a;
    layer6_outputs(565) <= '1';
    layer6_outputs(566) <= b;
    layer6_outputs(567) <= not a;
    layer6_outputs(568) <= b and not a;
    layer6_outputs(569) <= not b;
    layer6_outputs(570) <= b;
    layer6_outputs(571) <= a and not b;
    layer6_outputs(572) <= not b;
    layer6_outputs(573) <= a;
    layer6_outputs(574) <= a;
    layer6_outputs(575) <= b and not a;
    layer6_outputs(576) <= b;
    layer6_outputs(577) <= not (a xor b);
    layer6_outputs(578) <= a;
    layer6_outputs(579) <= a xor b;
    layer6_outputs(580) <= not b or a;
    layer6_outputs(581) <= b and not a;
    layer6_outputs(582) <= not (a and b);
    layer6_outputs(583) <= a or b;
    layer6_outputs(584) <= not a;
    layer6_outputs(585) <= a;
    layer6_outputs(586) <= a or b;
    layer6_outputs(587) <= '0';
    layer6_outputs(588) <= not b;
    layer6_outputs(589) <= not (a and b);
    layer6_outputs(590) <= not b;
    layer6_outputs(591) <= a or b;
    layer6_outputs(592) <= not (a xor b);
    layer6_outputs(593) <= a and not b;
    layer6_outputs(594) <= not a or b;
    layer6_outputs(595) <= b and not a;
    layer6_outputs(596) <= b;
    layer6_outputs(597) <= '0';
    layer6_outputs(598) <= not b;
    layer6_outputs(599) <= not a;
    layer6_outputs(600) <= not b;
    layer6_outputs(601) <= not b;
    layer6_outputs(602) <= a or b;
    layer6_outputs(603) <= a;
    layer6_outputs(604) <= not a;
    layer6_outputs(605) <= not b or a;
    layer6_outputs(606) <= a and b;
    layer6_outputs(607) <= not a;
    layer6_outputs(608) <= not a;
    layer6_outputs(609) <= a or b;
    layer6_outputs(610) <= not b or a;
    layer6_outputs(611) <= a;
    layer6_outputs(612) <= b;
    layer6_outputs(613) <= '0';
    layer6_outputs(614) <= not b;
    layer6_outputs(615) <= not b;
    layer6_outputs(616) <= a or b;
    layer6_outputs(617) <= not b;
    layer6_outputs(618) <= a or b;
    layer6_outputs(619) <= not b;
    layer6_outputs(620) <= a;
    layer6_outputs(621) <= a;
    layer6_outputs(622) <= a;
    layer6_outputs(623) <= b and not a;
    layer6_outputs(624) <= b;
    layer6_outputs(625) <= not b or a;
    layer6_outputs(626) <= a xor b;
    layer6_outputs(627) <= not (a xor b);
    layer6_outputs(628) <= a;
    layer6_outputs(629) <= not (a or b);
    layer6_outputs(630) <= a or b;
    layer6_outputs(631) <= not (a or b);
    layer6_outputs(632) <= a;
    layer6_outputs(633) <= not (a or b);
    layer6_outputs(634) <= b;
    layer6_outputs(635) <= not a or b;
    layer6_outputs(636) <= a and not b;
    layer6_outputs(637) <= not (a or b);
    layer6_outputs(638) <= not (a or b);
    layer6_outputs(639) <= a;
    layer6_outputs(640) <= a xor b;
    layer6_outputs(641) <= not (a and b);
    layer6_outputs(642) <= not b;
    layer6_outputs(643) <= a xor b;
    layer6_outputs(644) <= not (a and b);
    layer6_outputs(645) <= not (a and b);
    layer6_outputs(646) <= not b;
    layer6_outputs(647) <= not a or b;
    layer6_outputs(648) <= not (a and b);
    layer6_outputs(649) <= not b or a;
    layer6_outputs(650) <= b;
    layer6_outputs(651) <= not b;
    layer6_outputs(652) <= b;
    layer6_outputs(653) <= not a;
    layer6_outputs(654) <= not (a and b);
    layer6_outputs(655) <= not a;
    layer6_outputs(656) <= not (a or b);
    layer6_outputs(657) <= '1';
    layer6_outputs(658) <= not (a xor b);
    layer6_outputs(659) <= not a;
    layer6_outputs(660) <= not (a and b);
    layer6_outputs(661) <= b;
    layer6_outputs(662) <= a and not b;
    layer6_outputs(663) <= not a;
    layer6_outputs(664) <= a;
    layer6_outputs(665) <= not b;
    layer6_outputs(666) <= a xor b;
    layer6_outputs(667) <= not b or a;
    layer6_outputs(668) <= not b;
    layer6_outputs(669) <= not (a and b);
    layer6_outputs(670) <= not a;
    layer6_outputs(671) <= a and b;
    layer6_outputs(672) <= b;
    layer6_outputs(673) <= not b or a;
    layer6_outputs(674) <= not a;
    layer6_outputs(675) <= b and not a;
    layer6_outputs(676) <= a and not b;
    layer6_outputs(677) <= a and not b;
    layer6_outputs(678) <= not b;
    layer6_outputs(679) <= a xor b;
    layer6_outputs(680) <= not b;
    layer6_outputs(681) <= not (a and b);
    layer6_outputs(682) <= b;
    layer6_outputs(683) <= a and not b;
    layer6_outputs(684) <= b and not a;
    layer6_outputs(685) <= not a;
    layer6_outputs(686) <= a and not b;
    layer6_outputs(687) <= not a;
    layer6_outputs(688) <= '0';
    layer6_outputs(689) <= not (a and b);
    layer6_outputs(690) <= a;
    layer6_outputs(691) <= a or b;
    layer6_outputs(692) <= a and b;
    layer6_outputs(693) <= not a;
    layer6_outputs(694) <= b;
    layer6_outputs(695) <= a;
    layer6_outputs(696) <= not (a xor b);
    layer6_outputs(697) <= not b;
    layer6_outputs(698) <= a;
    layer6_outputs(699) <= a;
    layer6_outputs(700) <= a and not b;
    layer6_outputs(701) <= a or b;
    layer6_outputs(702) <= not a or b;
    layer6_outputs(703) <= b;
    layer6_outputs(704) <= not (a or b);
    layer6_outputs(705) <= not b;
    layer6_outputs(706) <= a;
    layer6_outputs(707) <= a;
    layer6_outputs(708) <= not (a or b);
    layer6_outputs(709) <= b;
    layer6_outputs(710) <= not a;
    layer6_outputs(711) <= a and not b;
    layer6_outputs(712) <= not b or a;
    layer6_outputs(713) <= a and not b;
    layer6_outputs(714) <= not (a or b);
    layer6_outputs(715) <= b;
    layer6_outputs(716) <= a and not b;
    layer6_outputs(717) <= not a;
    layer6_outputs(718) <= b;
    layer6_outputs(719) <= '0';
    layer6_outputs(720) <= b;
    layer6_outputs(721) <= not b;
    layer6_outputs(722) <= a;
    layer6_outputs(723) <= not a;
    layer6_outputs(724) <= a xor b;
    layer6_outputs(725) <= a;
    layer6_outputs(726) <= a;
    layer6_outputs(727) <= a or b;
    layer6_outputs(728) <= not (a and b);
    layer6_outputs(729) <= a or b;
    layer6_outputs(730) <= b;
    layer6_outputs(731) <= a;
    layer6_outputs(732) <= a;
    layer6_outputs(733) <= b;
    layer6_outputs(734) <= not a;
    layer6_outputs(735) <= b;
    layer6_outputs(736) <= not a or b;
    layer6_outputs(737) <= a and b;
    layer6_outputs(738) <= a xor b;
    layer6_outputs(739) <= b;
    layer6_outputs(740) <= not b;
    layer6_outputs(741) <= not (a or b);
    layer6_outputs(742) <= a;
    layer6_outputs(743) <= not b;
    layer6_outputs(744) <= b and not a;
    layer6_outputs(745) <= not a;
    layer6_outputs(746) <= a or b;
    layer6_outputs(747) <= a and b;
    layer6_outputs(748) <= not b;
    layer6_outputs(749) <= a xor b;
    layer6_outputs(750) <= not a;
    layer6_outputs(751) <= a xor b;
    layer6_outputs(752) <= not a;
    layer6_outputs(753) <= b;
    layer6_outputs(754) <= not (a xor b);
    layer6_outputs(755) <= not b;
    layer6_outputs(756) <= not b;
    layer6_outputs(757) <= not b;
    layer6_outputs(758) <= not a or b;
    layer6_outputs(759) <= a xor b;
    layer6_outputs(760) <= not b;
    layer6_outputs(761) <= not b or a;
    layer6_outputs(762) <= '1';
    layer6_outputs(763) <= a and not b;
    layer6_outputs(764) <= '1';
    layer6_outputs(765) <= a;
    layer6_outputs(766) <= b and not a;
    layer6_outputs(767) <= not b or a;
    layer6_outputs(768) <= b and not a;
    layer6_outputs(769) <= not a;
    layer6_outputs(770) <= not (a or b);
    layer6_outputs(771) <= '1';
    layer6_outputs(772) <= b;
    layer6_outputs(773) <= not b;
    layer6_outputs(774) <= '1';
    layer6_outputs(775) <= not a;
    layer6_outputs(776) <= b;
    layer6_outputs(777) <= b and not a;
    layer6_outputs(778) <= a;
    layer6_outputs(779) <= b;
    layer6_outputs(780) <= a and not b;
    layer6_outputs(781) <= not b;
    layer6_outputs(782) <= not (a or b);
    layer6_outputs(783) <= '1';
    layer6_outputs(784) <= a or b;
    layer6_outputs(785) <= b;
    layer6_outputs(786) <= not a;
    layer6_outputs(787) <= not (a or b);
    layer6_outputs(788) <= not a;
    layer6_outputs(789) <= not a or b;
    layer6_outputs(790) <= b;
    layer6_outputs(791) <= a and not b;
    layer6_outputs(792) <= b;
    layer6_outputs(793) <= not b or a;
    layer6_outputs(794) <= not (a or b);
    layer6_outputs(795) <= a;
    layer6_outputs(796) <= not a or b;
    layer6_outputs(797) <= not (a or b);
    layer6_outputs(798) <= a and not b;
    layer6_outputs(799) <= not a;
    layer6_outputs(800) <= a;
    layer6_outputs(801) <= not b or a;
    layer6_outputs(802) <= not (a xor b);
    layer6_outputs(803) <= a;
    layer6_outputs(804) <= not b;
    layer6_outputs(805) <= b;
    layer6_outputs(806) <= a;
    layer6_outputs(807) <= b;
    layer6_outputs(808) <= not (a xor b);
    layer6_outputs(809) <= a;
    layer6_outputs(810) <= b and not a;
    layer6_outputs(811) <= '0';
    layer6_outputs(812) <= a;
    layer6_outputs(813) <= a or b;
    layer6_outputs(814) <= '0';
    layer6_outputs(815) <= not (a or b);
    layer6_outputs(816) <= b;
    layer6_outputs(817) <= not a;
    layer6_outputs(818) <= not (a and b);
    layer6_outputs(819) <= not (a and b);
    layer6_outputs(820) <= a and b;
    layer6_outputs(821) <= a and b;
    layer6_outputs(822) <= not (a or b);
    layer6_outputs(823) <= not (a xor b);
    layer6_outputs(824) <= not b;
    layer6_outputs(825) <= not (a and b);
    layer6_outputs(826) <= not a or b;
    layer6_outputs(827) <= a;
    layer6_outputs(828) <= a xor b;
    layer6_outputs(829) <= a xor b;
    layer6_outputs(830) <= not (a and b);
    layer6_outputs(831) <= not (a xor b);
    layer6_outputs(832) <= a xor b;
    layer6_outputs(833) <= not b or a;
    layer6_outputs(834) <= b and not a;
    layer6_outputs(835) <= not a;
    layer6_outputs(836) <= not b or a;
    layer6_outputs(837) <= a and b;
    layer6_outputs(838) <= b;
    layer6_outputs(839) <= a;
    layer6_outputs(840) <= not b or a;
    layer6_outputs(841) <= not b;
    layer6_outputs(842) <= not a;
    layer6_outputs(843) <= not (a xor b);
    layer6_outputs(844) <= b and not a;
    layer6_outputs(845) <= not b or a;
    layer6_outputs(846) <= not a;
    layer6_outputs(847) <= b;
    layer6_outputs(848) <= a and b;
    layer6_outputs(849) <= a or b;
    layer6_outputs(850) <= b;
    layer6_outputs(851) <= b;
    layer6_outputs(852) <= not a;
    layer6_outputs(853) <= a and not b;
    layer6_outputs(854) <= a and b;
    layer6_outputs(855) <= b and not a;
    layer6_outputs(856) <= not b;
    layer6_outputs(857) <= not (a xor b);
    layer6_outputs(858) <= '0';
    layer6_outputs(859) <= a;
    layer6_outputs(860) <= b and not a;
    layer6_outputs(861) <= not (a and b);
    layer6_outputs(862) <= a;
    layer6_outputs(863) <= not b or a;
    layer6_outputs(864) <= a and not b;
    layer6_outputs(865) <= a or b;
    layer6_outputs(866) <= a;
    layer6_outputs(867) <= not a;
    layer6_outputs(868) <= a and not b;
    layer6_outputs(869) <= not a or b;
    layer6_outputs(870) <= a and b;
    layer6_outputs(871) <= not b or a;
    layer6_outputs(872) <= a and not b;
    layer6_outputs(873) <= b and not a;
    layer6_outputs(874) <= b;
    layer6_outputs(875) <= a xor b;
    layer6_outputs(876) <= not b;
    layer6_outputs(877) <= not (a or b);
    layer6_outputs(878) <= a;
    layer6_outputs(879) <= not a or b;
    layer6_outputs(880) <= a or b;
    layer6_outputs(881) <= not a;
    layer6_outputs(882) <= not (a or b);
    layer6_outputs(883) <= a xor b;
    layer6_outputs(884) <= a and not b;
    layer6_outputs(885) <= a or b;
    layer6_outputs(886) <= not b or a;
    layer6_outputs(887) <= not (a or b);
    layer6_outputs(888) <= '1';
    layer6_outputs(889) <= not (a xor b);
    layer6_outputs(890) <= not a;
    layer6_outputs(891) <= not a or b;
    layer6_outputs(892) <= not a or b;
    layer6_outputs(893) <= not a;
    layer6_outputs(894) <= not b;
    layer6_outputs(895) <= a xor b;
    layer6_outputs(896) <= not b;
    layer6_outputs(897) <= not b;
    layer6_outputs(898) <= a and b;
    layer6_outputs(899) <= a and b;
    layer6_outputs(900) <= a;
    layer6_outputs(901) <= a and b;
    layer6_outputs(902) <= not (a and b);
    layer6_outputs(903) <= a or b;
    layer6_outputs(904) <= b and not a;
    layer6_outputs(905) <= not b;
    layer6_outputs(906) <= not b or a;
    layer6_outputs(907) <= not a;
    layer6_outputs(908) <= not a;
    layer6_outputs(909) <= not a or b;
    layer6_outputs(910) <= a;
    layer6_outputs(911) <= a and not b;
    layer6_outputs(912) <= a and b;
    layer6_outputs(913) <= not a or b;
    layer6_outputs(914) <= b;
    layer6_outputs(915) <= not a or b;
    layer6_outputs(916) <= a and not b;
    layer6_outputs(917) <= not (a or b);
    layer6_outputs(918) <= not b;
    layer6_outputs(919) <= not a;
    layer6_outputs(920) <= '1';
    layer6_outputs(921) <= b;
    layer6_outputs(922) <= a or b;
    layer6_outputs(923) <= not (a and b);
    layer6_outputs(924) <= not (a or b);
    layer6_outputs(925) <= not a;
    layer6_outputs(926) <= not a;
    layer6_outputs(927) <= b;
    layer6_outputs(928) <= a xor b;
    layer6_outputs(929) <= not a;
    layer6_outputs(930) <= not b;
    layer6_outputs(931) <= not a;
    layer6_outputs(932) <= a and not b;
    layer6_outputs(933) <= not (a xor b);
    layer6_outputs(934) <= not (a and b);
    layer6_outputs(935) <= '1';
    layer6_outputs(936) <= a and b;
    layer6_outputs(937) <= not b;
    layer6_outputs(938) <= a and b;
    layer6_outputs(939) <= a and b;
    layer6_outputs(940) <= not (a and b);
    layer6_outputs(941) <= not (a and b);
    layer6_outputs(942) <= a and not b;
    layer6_outputs(943) <= not a;
    layer6_outputs(944) <= '1';
    layer6_outputs(945) <= not a;
    layer6_outputs(946) <= not (a or b);
    layer6_outputs(947) <= not b or a;
    layer6_outputs(948) <= b and not a;
    layer6_outputs(949) <= a;
    layer6_outputs(950) <= not a or b;
    layer6_outputs(951) <= a;
    layer6_outputs(952) <= a and b;
    layer6_outputs(953) <= a and not b;
    layer6_outputs(954) <= a;
    layer6_outputs(955) <= a xor b;
    layer6_outputs(956) <= a xor b;
    layer6_outputs(957) <= not b or a;
    layer6_outputs(958) <= not b;
    layer6_outputs(959) <= not a;
    layer6_outputs(960) <= '0';
    layer6_outputs(961) <= b;
    layer6_outputs(962) <= not (a and b);
    layer6_outputs(963) <= a or b;
    layer6_outputs(964) <= not a or b;
    layer6_outputs(965) <= not (a xor b);
    layer6_outputs(966) <= a and not b;
    layer6_outputs(967) <= a;
    layer6_outputs(968) <= a and not b;
    layer6_outputs(969) <= a xor b;
    layer6_outputs(970) <= not a;
    layer6_outputs(971) <= a and not b;
    layer6_outputs(972) <= not a;
    layer6_outputs(973) <= not (a or b);
    layer6_outputs(974) <= not b;
    layer6_outputs(975) <= not (a and b);
    layer6_outputs(976) <= not a;
    layer6_outputs(977) <= a and not b;
    layer6_outputs(978) <= b and not a;
    layer6_outputs(979) <= b;
    layer6_outputs(980) <= not (a or b);
    layer6_outputs(981) <= b and not a;
    layer6_outputs(982) <= not b;
    layer6_outputs(983) <= not b;
    layer6_outputs(984) <= a and not b;
    layer6_outputs(985) <= '1';
    layer6_outputs(986) <= not a or b;
    layer6_outputs(987) <= not a;
    layer6_outputs(988) <= not b;
    layer6_outputs(989) <= not a or b;
    layer6_outputs(990) <= b;
    layer6_outputs(991) <= a and not b;
    layer6_outputs(992) <= b and not a;
    layer6_outputs(993) <= a or b;
    layer6_outputs(994) <= not b;
    layer6_outputs(995) <= a or b;
    layer6_outputs(996) <= a or b;
    layer6_outputs(997) <= a and not b;
    layer6_outputs(998) <= a and b;
    layer6_outputs(999) <= not a;
    layer6_outputs(1000) <= not b;
    layer6_outputs(1001) <= a;
    layer6_outputs(1002) <= a and not b;
    layer6_outputs(1003) <= b;
    layer6_outputs(1004) <= not (a xor b);
    layer6_outputs(1005) <= a and not b;
    layer6_outputs(1006) <= not b or a;
    layer6_outputs(1007) <= not a;
    layer6_outputs(1008) <= not a;
    layer6_outputs(1009) <= a or b;
    layer6_outputs(1010) <= not a or b;
    layer6_outputs(1011) <= a or b;
    layer6_outputs(1012) <= a xor b;
    layer6_outputs(1013) <= a and not b;
    layer6_outputs(1014) <= a and not b;
    layer6_outputs(1015) <= not a;
    layer6_outputs(1016) <= not a or b;
    layer6_outputs(1017) <= a;
    layer6_outputs(1018) <= a;
    layer6_outputs(1019) <= not b;
    layer6_outputs(1020) <= not (a and b);
    layer6_outputs(1021) <= not (a and b);
    layer6_outputs(1022) <= not (a xor b);
    layer6_outputs(1023) <= not b;
    layer6_outputs(1024) <= not (a and b);
    layer6_outputs(1025) <= a xor b;
    layer6_outputs(1026) <= not (a xor b);
    layer6_outputs(1027) <= not (a and b);
    layer6_outputs(1028) <= a and not b;
    layer6_outputs(1029) <= a;
    layer6_outputs(1030) <= not b or a;
    layer6_outputs(1031) <= not a;
    layer6_outputs(1032) <= a and not b;
    layer6_outputs(1033) <= '1';
    layer6_outputs(1034) <= a xor b;
    layer6_outputs(1035) <= b and not a;
    layer6_outputs(1036) <= a;
    layer6_outputs(1037) <= a xor b;
    layer6_outputs(1038) <= not a;
    layer6_outputs(1039) <= not (a or b);
    layer6_outputs(1040) <= a xor b;
    layer6_outputs(1041) <= not a;
    layer6_outputs(1042) <= not (a and b);
    layer6_outputs(1043) <= not (a or b);
    layer6_outputs(1044) <= b and not a;
    layer6_outputs(1045) <= b and not a;
    layer6_outputs(1046) <= '1';
    layer6_outputs(1047) <= not (a and b);
    layer6_outputs(1048) <= a and not b;
    layer6_outputs(1049) <= a and not b;
    layer6_outputs(1050) <= not b;
    layer6_outputs(1051) <= '1';
    layer6_outputs(1052) <= not a or b;
    layer6_outputs(1053) <= a and not b;
    layer6_outputs(1054) <= not b;
    layer6_outputs(1055) <= not (a or b);
    layer6_outputs(1056) <= a and not b;
    layer6_outputs(1057) <= a and not b;
    layer6_outputs(1058) <= a and not b;
    layer6_outputs(1059) <= a and b;
    layer6_outputs(1060) <= '1';
    layer6_outputs(1061) <= not b or a;
    layer6_outputs(1062) <= a;
    layer6_outputs(1063) <= not b or a;
    layer6_outputs(1064) <= not b;
    layer6_outputs(1065) <= not b;
    layer6_outputs(1066) <= b and not a;
    layer6_outputs(1067) <= not (a xor b);
    layer6_outputs(1068) <= not (a or b);
    layer6_outputs(1069) <= a and b;
    layer6_outputs(1070) <= not (a or b);
    layer6_outputs(1071) <= not b;
    layer6_outputs(1072) <= not b;
    layer6_outputs(1073) <= not b or a;
    layer6_outputs(1074) <= a;
    layer6_outputs(1075) <= b;
    layer6_outputs(1076) <= b;
    layer6_outputs(1077) <= not (a xor b);
    layer6_outputs(1078) <= not a;
    layer6_outputs(1079) <= a xor b;
    layer6_outputs(1080) <= not a;
    layer6_outputs(1081) <= a or b;
    layer6_outputs(1082) <= b and not a;
    layer6_outputs(1083) <= b;
    layer6_outputs(1084) <= b;
    layer6_outputs(1085) <= not a;
    layer6_outputs(1086) <= a and not b;
    layer6_outputs(1087) <= a and b;
    layer6_outputs(1088) <= not b;
    layer6_outputs(1089) <= not b or a;
    layer6_outputs(1090) <= not a;
    layer6_outputs(1091) <= b and not a;
    layer6_outputs(1092) <= not (a xor b);
    layer6_outputs(1093) <= not a or b;
    layer6_outputs(1094) <= '0';
    layer6_outputs(1095) <= not a;
    layer6_outputs(1096) <= a;
    layer6_outputs(1097) <= a or b;
    layer6_outputs(1098) <= '0';
    layer6_outputs(1099) <= a;
    layer6_outputs(1100) <= not a;
    layer6_outputs(1101) <= b;
    layer6_outputs(1102) <= a xor b;
    layer6_outputs(1103) <= not b or a;
    layer6_outputs(1104) <= not a;
    layer6_outputs(1105) <= a;
    layer6_outputs(1106) <= not a;
    layer6_outputs(1107) <= not b;
    layer6_outputs(1108) <= not (a and b);
    layer6_outputs(1109) <= b and not a;
    layer6_outputs(1110) <= a and b;
    layer6_outputs(1111) <= a and not b;
    layer6_outputs(1112) <= a or b;
    layer6_outputs(1113) <= not a or b;
    layer6_outputs(1114) <= a;
    layer6_outputs(1115) <= a or b;
    layer6_outputs(1116) <= not b;
    layer6_outputs(1117) <= not b;
    layer6_outputs(1118) <= b and not a;
    layer6_outputs(1119) <= a and b;
    layer6_outputs(1120) <= not (a and b);
    layer6_outputs(1121) <= a and b;
    layer6_outputs(1122) <= not (a xor b);
    layer6_outputs(1123) <= a;
    layer6_outputs(1124) <= not (a and b);
    layer6_outputs(1125) <= not b;
    layer6_outputs(1126) <= not b;
    layer6_outputs(1127) <= b and not a;
    layer6_outputs(1128) <= a and b;
    layer6_outputs(1129) <= a;
    layer6_outputs(1130) <= not a;
    layer6_outputs(1131) <= a or b;
    layer6_outputs(1132) <= b and not a;
    layer6_outputs(1133) <= a and not b;
    layer6_outputs(1134) <= a;
    layer6_outputs(1135) <= b;
    layer6_outputs(1136) <= a or b;
    layer6_outputs(1137) <= not (a or b);
    layer6_outputs(1138) <= a and b;
    layer6_outputs(1139) <= b;
    layer6_outputs(1140) <= a and b;
    layer6_outputs(1141) <= not a;
    layer6_outputs(1142) <= not a or b;
    layer6_outputs(1143) <= not (a or b);
    layer6_outputs(1144) <= a or b;
    layer6_outputs(1145) <= b;
    layer6_outputs(1146) <= b;
    layer6_outputs(1147) <= b;
    layer6_outputs(1148) <= not (a xor b);
    layer6_outputs(1149) <= a xor b;
    layer6_outputs(1150) <= not a or b;
    layer6_outputs(1151) <= a;
    layer6_outputs(1152) <= a;
    layer6_outputs(1153) <= not a or b;
    layer6_outputs(1154) <= a;
    layer6_outputs(1155) <= not a;
    layer6_outputs(1156) <= not b;
    layer6_outputs(1157) <= not a;
    layer6_outputs(1158) <= not b;
    layer6_outputs(1159) <= a or b;
    layer6_outputs(1160) <= '0';
    layer6_outputs(1161) <= not (a and b);
    layer6_outputs(1162) <= b;
    layer6_outputs(1163) <= a;
    layer6_outputs(1164) <= a or b;
    layer6_outputs(1165) <= not a;
    layer6_outputs(1166) <= not a;
    layer6_outputs(1167) <= b;
    layer6_outputs(1168) <= a and not b;
    layer6_outputs(1169) <= a xor b;
    layer6_outputs(1170) <= not (a and b);
    layer6_outputs(1171) <= b;
    layer6_outputs(1172) <= not b;
    layer6_outputs(1173) <= not (a and b);
    layer6_outputs(1174) <= a and b;
    layer6_outputs(1175) <= not (a xor b);
    layer6_outputs(1176) <= not b;
    layer6_outputs(1177) <= a or b;
    layer6_outputs(1178) <= b and not a;
    layer6_outputs(1179) <= not a;
    layer6_outputs(1180) <= not a or b;
    layer6_outputs(1181) <= not a;
    layer6_outputs(1182) <= a xor b;
    layer6_outputs(1183) <= not b;
    layer6_outputs(1184) <= '0';
    layer6_outputs(1185) <= not (a and b);
    layer6_outputs(1186) <= not b;
    layer6_outputs(1187) <= a or b;
    layer6_outputs(1188) <= not a;
    layer6_outputs(1189) <= not b or a;
    layer6_outputs(1190) <= not b or a;
    layer6_outputs(1191) <= not b;
    layer6_outputs(1192) <= b;
    layer6_outputs(1193) <= a xor b;
    layer6_outputs(1194) <= a xor b;
    layer6_outputs(1195) <= not a;
    layer6_outputs(1196) <= not b;
    layer6_outputs(1197) <= a;
    layer6_outputs(1198) <= b and not a;
    layer6_outputs(1199) <= not b;
    layer6_outputs(1200) <= not b;
    layer6_outputs(1201) <= not b;
    layer6_outputs(1202) <= b and not a;
    layer6_outputs(1203) <= a xor b;
    layer6_outputs(1204) <= not (a and b);
    layer6_outputs(1205) <= not (a xor b);
    layer6_outputs(1206) <= not a;
    layer6_outputs(1207) <= '1';
    layer6_outputs(1208) <= a;
    layer6_outputs(1209) <= not (a xor b);
    layer6_outputs(1210) <= not (a or b);
    layer6_outputs(1211) <= b and not a;
    layer6_outputs(1212) <= not b;
    layer6_outputs(1213) <= not a or b;
    layer6_outputs(1214) <= a or b;
    layer6_outputs(1215) <= a;
    layer6_outputs(1216) <= b;
    layer6_outputs(1217) <= a xor b;
    layer6_outputs(1218) <= not b;
    layer6_outputs(1219) <= a xor b;
    layer6_outputs(1220) <= not a;
    layer6_outputs(1221) <= a;
    layer6_outputs(1222) <= not a;
    layer6_outputs(1223) <= a and not b;
    layer6_outputs(1224) <= not (a and b);
    layer6_outputs(1225) <= a or b;
    layer6_outputs(1226) <= not a or b;
    layer6_outputs(1227) <= not (a and b);
    layer6_outputs(1228) <= not (a or b);
    layer6_outputs(1229) <= b and not a;
    layer6_outputs(1230) <= a xor b;
    layer6_outputs(1231) <= a;
    layer6_outputs(1232) <= b;
    layer6_outputs(1233) <= a and not b;
    layer6_outputs(1234) <= not b;
    layer6_outputs(1235) <= b;
    layer6_outputs(1236) <= not a or b;
    layer6_outputs(1237) <= a;
    layer6_outputs(1238) <= not b;
    layer6_outputs(1239) <= a;
    layer6_outputs(1240) <= not (a or b);
    layer6_outputs(1241) <= a and not b;
    layer6_outputs(1242) <= a;
    layer6_outputs(1243) <= a;
    layer6_outputs(1244) <= not a;
    layer6_outputs(1245) <= not b or a;
    layer6_outputs(1246) <= not (a or b);
    layer6_outputs(1247) <= b;
    layer6_outputs(1248) <= a or b;
    layer6_outputs(1249) <= not a;
    layer6_outputs(1250) <= not a;
    layer6_outputs(1251) <= not a;
    layer6_outputs(1252) <= not a;
    layer6_outputs(1253) <= not (a xor b);
    layer6_outputs(1254) <= a and not b;
    layer6_outputs(1255) <= not (a or b);
    layer6_outputs(1256) <= a xor b;
    layer6_outputs(1257) <= not (a and b);
    layer6_outputs(1258) <= not b;
    layer6_outputs(1259) <= not (a xor b);
    layer6_outputs(1260) <= not (a xor b);
    layer6_outputs(1261) <= not b;
    layer6_outputs(1262) <= not b;
    layer6_outputs(1263) <= b and not a;
    layer6_outputs(1264) <= b;
    layer6_outputs(1265) <= not a;
    layer6_outputs(1266) <= a;
    layer6_outputs(1267) <= a or b;
    layer6_outputs(1268) <= not a or b;
    layer6_outputs(1269) <= b and not a;
    layer6_outputs(1270) <= not (a xor b);
    layer6_outputs(1271) <= a and b;
    layer6_outputs(1272) <= not a;
    layer6_outputs(1273) <= b and not a;
    layer6_outputs(1274) <= a and not b;
    layer6_outputs(1275) <= not a or b;
    layer6_outputs(1276) <= not b;
    layer6_outputs(1277) <= not (a and b);
    layer6_outputs(1278) <= not b;
    layer6_outputs(1279) <= b;
    layer6_outputs(1280) <= a;
    layer6_outputs(1281) <= not (a and b);
    layer6_outputs(1282) <= not (a xor b);
    layer6_outputs(1283) <= a xor b;
    layer6_outputs(1284) <= not b;
    layer6_outputs(1285) <= a and b;
    layer6_outputs(1286) <= not (a or b);
    layer6_outputs(1287) <= not (a xor b);
    layer6_outputs(1288) <= not (a or b);
    layer6_outputs(1289) <= not b or a;
    layer6_outputs(1290) <= a;
    layer6_outputs(1291) <= '0';
    layer6_outputs(1292) <= not (a and b);
    layer6_outputs(1293) <= not (a and b);
    layer6_outputs(1294) <= not b;
    layer6_outputs(1295) <= a xor b;
    layer6_outputs(1296) <= a;
    layer6_outputs(1297) <= not a;
    layer6_outputs(1298) <= not (a or b);
    layer6_outputs(1299) <= not a;
    layer6_outputs(1300) <= not (a and b);
    layer6_outputs(1301) <= not (a xor b);
    layer6_outputs(1302) <= not b or a;
    layer6_outputs(1303) <= a;
    layer6_outputs(1304) <= not a;
    layer6_outputs(1305) <= not b or a;
    layer6_outputs(1306) <= a xor b;
    layer6_outputs(1307) <= '1';
    layer6_outputs(1308) <= a;
    layer6_outputs(1309) <= a;
    layer6_outputs(1310) <= not a or b;
    layer6_outputs(1311) <= b and not a;
    layer6_outputs(1312) <= not a;
    layer6_outputs(1313) <= '0';
    layer6_outputs(1314) <= not b;
    layer6_outputs(1315) <= not b;
    layer6_outputs(1316) <= not b or a;
    layer6_outputs(1317) <= not (a or b);
    layer6_outputs(1318) <= not a;
    layer6_outputs(1319) <= not a;
    layer6_outputs(1320) <= b and not a;
    layer6_outputs(1321) <= not b or a;
    layer6_outputs(1322) <= a;
    layer6_outputs(1323) <= a and b;
    layer6_outputs(1324) <= not (a or b);
    layer6_outputs(1325) <= not a;
    layer6_outputs(1326) <= a and b;
    layer6_outputs(1327) <= not (a xor b);
    layer6_outputs(1328) <= not b or a;
    layer6_outputs(1329) <= not a;
    layer6_outputs(1330) <= not a;
    layer6_outputs(1331) <= not (a and b);
    layer6_outputs(1332) <= a xor b;
    layer6_outputs(1333) <= not a or b;
    layer6_outputs(1334) <= b;
    layer6_outputs(1335) <= b;
    layer6_outputs(1336) <= not b;
    layer6_outputs(1337) <= not a or b;
    layer6_outputs(1338) <= not (a and b);
    layer6_outputs(1339) <= not (a xor b);
    layer6_outputs(1340) <= not b;
    layer6_outputs(1341) <= not a;
    layer6_outputs(1342) <= b;
    layer6_outputs(1343) <= a xor b;
    layer6_outputs(1344) <= a and b;
    layer6_outputs(1345) <= a and b;
    layer6_outputs(1346) <= a and not b;
    layer6_outputs(1347) <= a;
    layer6_outputs(1348) <= a;
    layer6_outputs(1349) <= b and not a;
    layer6_outputs(1350) <= a xor b;
    layer6_outputs(1351) <= '1';
    layer6_outputs(1352) <= a and not b;
    layer6_outputs(1353) <= a and not b;
    layer6_outputs(1354) <= '0';
    layer6_outputs(1355) <= a and not b;
    layer6_outputs(1356) <= not a;
    layer6_outputs(1357) <= not (a and b);
    layer6_outputs(1358) <= a and not b;
    layer6_outputs(1359) <= b and not a;
    layer6_outputs(1360) <= not (a and b);
    layer6_outputs(1361) <= not (a or b);
    layer6_outputs(1362) <= a and not b;
    layer6_outputs(1363) <= not a;
    layer6_outputs(1364) <= not (a or b);
    layer6_outputs(1365) <= not b;
    layer6_outputs(1366) <= a;
    layer6_outputs(1367) <= not a or b;
    layer6_outputs(1368) <= not (a and b);
    layer6_outputs(1369) <= not b;
    layer6_outputs(1370) <= not a;
    layer6_outputs(1371) <= not (a and b);
    layer6_outputs(1372) <= a;
    layer6_outputs(1373) <= a xor b;
    layer6_outputs(1374) <= a and not b;
    layer6_outputs(1375) <= a;
    layer6_outputs(1376) <= not b;
    layer6_outputs(1377) <= not b or a;
    layer6_outputs(1378) <= a xor b;
    layer6_outputs(1379) <= a;
    layer6_outputs(1380) <= not b;
    layer6_outputs(1381) <= a and b;
    layer6_outputs(1382) <= b and not a;
    layer6_outputs(1383) <= not b;
    layer6_outputs(1384) <= '0';
    layer6_outputs(1385) <= a xor b;
    layer6_outputs(1386) <= not a or b;
    layer6_outputs(1387) <= '0';
    layer6_outputs(1388) <= not (a xor b);
    layer6_outputs(1389) <= not (a xor b);
    layer6_outputs(1390) <= b and not a;
    layer6_outputs(1391) <= a and not b;
    layer6_outputs(1392) <= a;
    layer6_outputs(1393) <= not b or a;
    layer6_outputs(1394) <= b;
    layer6_outputs(1395) <= a;
    layer6_outputs(1396) <= not (a or b);
    layer6_outputs(1397) <= b and not a;
    layer6_outputs(1398) <= b;
    layer6_outputs(1399) <= a and not b;
    layer6_outputs(1400) <= not b;
    layer6_outputs(1401) <= b;
    layer6_outputs(1402) <= '1';
    layer6_outputs(1403) <= not (a or b);
    layer6_outputs(1404) <= not b;
    layer6_outputs(1405) <= a and not b;
    layer6_outputs(1406) <= not b or a;
    layer6_outputs(1407) <= a and not b;
    layer6_outputs(1408) <= b;
    layer6_outputs(1409) <= a;
    layer6_outputs(1410) <= a and not b;
    layer6_outputs(1411) <= not (a or b);
    layer6_outputs(1412) <= not a;
    layer6_outputs(1413) <= '0';
    layer6_outputs(1414) <= b;
    layer6_outputs(1415) <= not a or b;
    layer6_outputs(1416) <= b;
    layer6_outputs(1417) <= b and not a;
    layer6_outputs(1418) <= a and b;
    layer6_outputs(1419) <= not a or b;
    layer6_outputs(1420) <= a and not b;
    layer6_outputs(1421) <= a;
    layer6_outputs(1422) <= not (a or b);
    layer6_outputs(1423) <= not (a and b);
    layer6_outputs(1424) <= not b;
    layer6_outputs(1425) <= a or b;
    layer6_outputs(1426) <= a xor b;
    layer6_outputs(1427) <= not a;
    layer6_outputs(1428) <= b;
    layer6_outputs(1429) <= a;
    layer6_outputs(1430) <= a and b;
    layer6_outputs(1431) <= not (a or b);
    layer6_outputs(1432) <= b and not a;
    layer6_outputs(1433) <= not b;
    layer6_outputs(1434) <= not b;
    layer6_outputs(1435) <= not (a or b);
    layer6_outputs(1436) <= a and not b;
    layer6_outputs(1437) <= b;
    layer6_outputs(1438) <= not a;
    layer6_outputs(1439) <= a;
    layer6_outputs(1440) <= a xor b;
    layer6_outputs(1441) <= not (a xor b);
    layer6_outputs(1442) <= not b;
    layer6_outputs(1443) <= a and not b;
    layer6_outputs(1444) <= a and not b;
    layer6_outputs(1445) <= a or b;
    layer6_outputs(1446) <= not a;
    layer6_outputs(1447) <= not b or a;
    layer6_outputs(1448) <= not (a or b);
    layer6_outputs(1449) <= a;
    layer6_outputs(1450) <= a and b;
    layer6_outputs(1451) <= a;
    layer6_outputs(1452) <= not (a and b);
    layer6_outputs(1453) <= not (a xor b);
    layer6_outputs(1454) <= not (a xor b);
    layer6_outputs(1455) <= not b or a;
    layer6_outputs(1456) <= not a;
    layer6_outputs(1457) <= a or b;
    layer6_outputs(1458) <= not a;
    layer6_outputs(1459) <= '1';
    layer6_outputs(1460) <= b;
    layer6_outputs(1461) <= a and b;
    layer6_outputs(1462) <= not b or a;
    layer6_outputs(1463) <= b;
    layer6_outputs(1464) <= a and b;
    layer6_outputs(1465) <= b;
    layer6_outputs(1466) <= a;
    layer6_outputs(1467) <= a and not b;
    layer6_outputs(1468) <= not a or b;
    layer6_outputs(1469) <= b;
    layer6_outputs(1470) <= b and not a;
    layer6_outputs(1471) <= b;
    layer6_outputs(1472) <= not b;
    layer6_outputs(1473) <= not b;
    layer6_outputs(1474) <= b;
    layer6_outputs(1475) <= b;
    layer6_outputs(1476) <= a and not b;
    layer6_outputs(1477) <= not a or b;
    layer6_outputs(1478) <= not b;
    layer6_outputs(1479) <= not (a or b);
    layer6_outputs(1480) <= '1';
    layer6_outputs(1481) <= a;
    layer6_outputs(1482) <= a and not b;
    layer6_outputs(1483) <= a and b;
    layer6_outputs(1484) <= not a;
    layer6_outputs(1485) <= a xor b;
    layer6_outputs(1486) <= not b;
    layer6_outputs(1487) <= not (a and b);
    layer6_outputs(1488) <= not b;
    layer6_outputs(1489) <= not b;
    layer6_outputs(1490) <= not a or b;
    layer6_outputs(1491) <= not b;
    layer6_outputs(1492) <= not (a and b);
    layer6_outputs(1493) <= not b;
    layer6_outputs(1494) <= a;
    layer6_outputs(1495) <= a;
    layer6_outputs(1496) <= a;
    layer6_outputs(1497) <= a;
    layer6_outputs(1498) <= a and b;
    layer6_outputs(1499) <= a or b;
    layer6_outputs(1500) <= not b;
    layer6_outputs(1501) <= b;
    layer6_outputs(1502) <= b;
    layer6_outputs(1503) <= a;
    layer6_outputs(1504) <= b;
    layer6_outputs(1505) <= a and b;
    layer6_outputs(1506) <= not a;
    layer6_outputs(1507) <= a xor b;
    layer6_outputs(1508) <= not b;
    layer6_outputs(1509) <= '1';
    layer6_outputs(1510) <= b and not a;
    layer6_outputs(1511) <= b;
    layer6_outputs(1512) <= not b;
    layer6_outputs(1513) <= not b;
    layer6_outputs(1514) <= a;
    layer6_outputs(1515) <= a and not b;
    layer6_outputs(1516) <= a xor b;
    layer6_outputs(1517) <= a xor b;
    layer6_outputs(1518) <= a or b;
    layer6_outputs(1519) <= a and b;
    layer6_outputs(1520) <= not a or b;
    layer6_outputs(1521) <= not a;
    layer6_outputs(1522) <= '1';
    layer6_outputs(1523) <= not (a xor b);
    layer6_outputs(1524) <= not (a xor b);
    layer6_outputs(1525) <= a and not b;
    layer6_outputs(1526) <= a;
    layer6_outputs(1527) <= b and not a;
    layer6_outputs(1528) <= a xor b;
    layer6_outputs(1529) <= not a;
    layer6_outputs(1530) <= not a;
    layer6_outputs(1531) <= not (a or b);
    layer6_outputs(1532) <= b;
    layer6_outputs(1533) <= not a;
    layer6_outputs(1534) <= b;
    layer6_outputs(1535) <= a and not b;
    layer6_outputs(1536) <= a and not b;
    layer6_outputs(1537) <= a and not b;
    layer6_outputs(1538) <= not (a xor b);
    layer6_outputs(1539) <= not a;
    layer6_outputs(1540) <= not a;
    layer6_outputs(1541) <= a xor b;
    layer6_outputs(1542) <= not a;
    layer6_outputs(1543) <= not a;
    layer6_outputs(1544) <= '1';
    layer6_outputs(1545) <= b;
    layer6_outputs(1546) <= not (a or b);
    layer6_outputs(1547) <= not b;
    layer6_outputs(1548) <= a or b;
    layer6_outputs(1549) <= a xor b;
    layer6_outputs(1550) <= not (a and b);
    layer6_outputs(1551) <= not b or a;
    layer6_outputs(1552) <= not b;
    layer6_outputs(1553) <= '1';
    layer6_outputs(1554) <= not b;
    layer6_outputs(1555) <= a and b;
    layer6_outputs(1556) <= a and not b;
    layer6_outputs(1557) <= a xor b;
    layer6_outputs(1558) <= a;
    layer6_outputs(1559) <= a xor b;
    layer6_outputs(1560) <= not a;
    layer6_outputs(1561) <= a xor b;
    layer6_outputs(1562) <= not b;
    layer6_outputs(1563) <= not b;
    layer6_outputs(1564) <= not (a xor b);
    layer6_outputs(1565) <= not b;
    layer6_outputs(1566) <= a and b;
    layer6_outputs(1567) <= b;
    layer6_outputs(1568) <= a and not b;
    layer6_outputs(1569) <= a;
    layer6_outputs(1570) <= not (a or b);
    layer6_outputs(1571) <= not (a and b);
    layer6_outputs(1572) <= '0';
    layer6_outputs(1573) <= not a;
    layer6_outputs(1574) <= b and not a;
    layer6_outputs(1575) <= not a or b;
    layer6_outputs(1576) <= a;
    layer6_outputs(1577) <= a and b;
    layer6_outputs(1578) <= not (a and b);
    layer6_outputs(1579) <= not (a xor b);
    layer6_outputs(1580) <= b;
    layer6_outputs(1581) <= '1';
    layer6_outputs(1582) <= b;
    layer6_outputs(1583) <= '0';
    layer6_outputs(1584) <= not b;
    layer6_outputs(1585) <= a xor b;
    layer6_outputs(1586) <= b;
    layer6_outputs(1587) <= not b;
    layer6_outputs(1588) <= a and b;
    layer6_outputs(1589) <= a or b;
    layer6_outputs(1590) <= a;
    layer6_outputs(1591) <= a;
    layer6_outputs(1592) <= b and not a;
    layer6_outputs(1593) <= b and not a;
    layer6_outputs(1594) <= not b;
    layer6_outputs(1595) <= not a or b;
    layer6_outputs(1596) <= a or b;
    layer6_outputs(1597) <= a xor b;
    layer6_outputs(1598) <= not (a or b);
    layer6_outputs(1599) <= a and b;
    layer6_outputs(1600) <= b;
    layer6_outputs(1601) <= '0';
    layer6_outputs(1602) <= not (a and b);
    layer6_outputs(1603) <= not a;
    layer6_outputs(1604) <= b;
    layer6_outputs(1605) <= b;
    layer6_outputs(1606) <= a;
    layer6_outputs(1607) <= not a or b;
    layer6_outputs(1608) <= a and not b;
    layer6_outputs(1609) <= b;
    layer6_outputs(1610) <= not a or b;
    layer6_outputs(1611) <= '1';
    layer6_outputs(1612) <= not b or a;
    layer6_outputs(1613) <= a or b;
    layer6_outputs(1614) <= a or b;
    layer6_outputs(1615) <= not a or b;
    layer6_outputs(1616) <= not b;
    layer6_outputs(1617) <= a or b;
    layer6_outputs(1618) <= not (a or b);
    layer6_outputs(1619) <= a xor b;
    layer6_outputs(1620) <= a;
    layer6_outputs(1621) <= not a;
    layer6_outputs(1622) <= not (a or b);
    layer6_outputs(1623) <= not a or b;
    layer6_outputs(1624) <= not (a xor b);
    layer6_outputs(1625) <= not a;
    layer6_outputs(1626) <= not (a or b);
    layer6_outputs(1627) <= a or b;
    layer6_outputs(1628) <= not a;
    layer6_outputs(1629) <= not b;
    layer6_outputs(1630) <= a;
    layer6_outputs(1631) <= a and b;
    layer6_outputs(1632) <= b and not a;
    layer6_outputs(1633) <= a;
    layer6_outputs(1634) <= not (a or b);
    layer6_outputs(1635) <= not b or a;
    layer6_outputs(1636) <= not b;
    layer6_outputs(1637) <= a and not b;
    layer6_outputs(1638) <= a and not b;
    layer6_outputs(1639) <= b;
    layer6_outputs(1640) <= not a;
    layer6_outputs(1641) <= not a;
    layer6_outputs(1642) <= not a;
    layer6_outputs(1643) <= not b or a;
    layer6_outputs(1644) <= b;
    layer6_outputs(1645) <= a xor b;
    layer6_outputs(1646) <= not b;
    layer6_outputs(1647) <= b and not a;
    layer6_outputs(1648) <= b;
    layer6_outputs(1649) <= a;
    layer6_outputs(1650) <= a or b;
    layer6_outputs(1651) <= b;
    layer6_outputs(1652) <= not b or a;
    layer6_outputs(1653) <= a;
    layer6_outputs(1654) <= not (a or b);
    layer6_outputs(1655) <= not (a xor b);
    layer6_outputs(1656) <= b;
    layer6_outputs(1657) <= a and not b;
    layer6_outputs(1658) <= not b;
    layer6_outputs(1659) <= a;
    layer6_outputs(1660) <= a;
    layer6_outputs(1661) <= b and not a;
    layer6_outputs(1662) <= a and b;
    layer6_outputs(1663) <= a;
    layer6_outputs(1664) <= not (a or b);
    layer6_outputs(1665) <= not (a or b);
    layer6_outputs(1666) <= not b or a;
    layer6_outputs(1667) <= '1';
    layer6_outputs(1668) <= not (a xor b);
    layer6_outputs(1669) <= a;
    layer6_outputs(1670) <= not a;
    layer6_outputs(1671) <= not a;
    layer6_outputs(1672) <= a and not b;
    layer6_outputs(1673) <= a;
    layer6_outputs(1674) <= not (a or b);
    layer6_outputs(1675) <= '1';
    layer6_outputs(1676) <= not b or a;
    layer6_outputs(1677) <= not (a or b);
    layer6_outputs(1678) <= not a;
    layer6_outputs(1679) <= a;
    layer6_outputs(1680) <= not b or a;
    layer6_outputs(1681) <= not a;
    layer6_outputs(1682) <= not (a and b);
    layer6_outputs(1683) <= b;
    layer6_outputs(1684) <= not a or b;
    layer6_outputs(1685) <= b;
    layer6_outputs(1686) <= not (a and b);
    layer6_outputs(1687) <= not (a or b);
    layer6_outputs(1688) <= b;
    layer6_outputs(1689) <= b;
    layer6_outputs(1690) <= a or b;
    layer6_outputs(1691) <= not a;
    layer6_outputs(1692) <= not a;
    layer6_outputs(1693) <= not a;
    layer6_outputs(1694) <= a;
    layer6_outputs(1695) <= a or b;
    layer6_outputs(1696) <= not a;
    layer6_outputs(1697) <= b;
    layer6_outputs(1698) <= not b;
    layer6_outputs(1699) <= a;
    layer6_outputs(1700) <= not a;
    layer6_outputs(1701) <= not b;
    layer6_outputs(1702) <= a;
    layer6_outputs(1703) <= not b;
    layer6_outputs(1704) <= a and not b;
    layer6_outputs(1705) <= a and b;
    layer6_outputs(1706) <= not a;
    layer6_outputs(1707) <= not (a and b);
    layer6_outputs(1708) <= b;
    layer6_outputs(1709) <= not b;
    layer6_outputs(1710) <= not (a or b);
    layer6_outputs(1711) <= a xor b;
    layer6_outputs(1712) <= not b or a;
    layer6_outputs(1713) <= not b or a;
    layer6_outputs(1714) <= not b or a;
    layer6_outputs(1715) <= not a;
    layer6_outputs(1716) <= not b or a;
    layer6_outputs(1717) <= b;
    layer6_outputs(1718) <= not b or a;
    layer6_outputs(1719) <= a or b;
    layer6_outputs(1720) <= a and b;
    layer6_outputs(1721) <= not (a or b);
    layer6_outputs(1722) <= not b or a;
    layer6_outputs(1723) <= a;
    layer6_outputs(1724) <= a and not b;
    layer6_outputs(1725) <= a or b;
    layer6_outputs(1726) <= b and not a;
    layer6_outputs(1727) <= not (a or b);
    layer6_outputs(1728) <= not b;
    layer6_outputs(1729) <= not a;
    layer6_outputs(1730) <= not (a or b);
    layer6_outputs(1731) <= b and not a;
    layer6_outputs(1732) <= not (a and b);
    layer6_outputs(1733) <= not a;
    layer6_outputs(1734) <= a and not b;
    layer6_outputs(1735) <= a xor b;
    layer6_outputs(1736) <= not (a and b);
    layer6_outputs(1737) <= a and b;
    layer6_outputs(1738) <= not b;
    layer6_outputs(1739) <= b and not a;
    layer6_outputs(1740) <= not b or a;
    layer6_outputs(1741) <= '0';
    layer6_outputs(1742) <= not b;
    layer6_outputs(1743) <= a and b;
    layer6_outputs(1744) <= not (a xor b);
    layer6_outputs(1745) <= not a or b;
    layer6_outputs(1746) <= not a;
    layer6_outputs(1747) <= not (a xor b);
    layer6_outputs(1748) <= not a;
    layer6_outputs(1749) <= not a;
    layer6_outputs(1750) <= a and not b;
    layer6_outputs(1751) <= not a;
    layer6_outputs(1752) <= a;
    layer6_outputs(1753) <= a and b;
    layer6_outputs(1754) <= not b or a;
    layer6_outputs(1755) <= not (a and b);
    layer6_outputs(1756) <= b;
    layer6_outputs(1757) <= not a;
    layer6_outputs(1758) <= not (a or b);
    layer6_outputs(1759) <= not b;
    layer6_outputs(1760) <= b;
    layer6_outputs(1761) <= b;
    layer6_outputs(1762) <= not b;
    layer6_outputs(1763) <= not (a xor b);
    layer6_outputs(1764) <= not (a or b);
    layer6_outputs(1765) <= not a or b;
    layer6_outputs(1766) <= not a or b;
    layer6_outputs(1767) <= not (a xor b);
    layer6_outputs(1768) <= a;
    layer6_outputs(1769) <= not a;
    layer6_outputs(1770) <= not a or b;
    layer6_outputs(1771) <= a;
    layer6_outputs(1772) <= not (a or b);
    layer6_outputs(1773) <= not a;
    layer6_outputs(1774) <= not a;
    layer6_outputs(1775) <= a xor b;
    layer6_outputs(1776) <= not b;
    layer6_outputs(1777) <= a and not b;
    layer6_outputs(1778) <= a or b;
    layer6_outputs(1779) <= a and not b;
    layer6_outputs(1780) <= not (a and b);
    layer6_outputs(1781) <= not (a xor b);
    layer6_outputs(1782) <= b and not a;
    layer6_outputs(1783) <= b and not a;
    layer6_outputs(1784) <= a xor b;
    layer6_outputs(1785) <= not a;
    layer6_outputs(1786) <= not b or a;
    layer6_outputs(1787) <= a and b;
    layer6_outputs(1788) <= a and b;
    layer6_outputs(1789) <= not b or a;
    layer6_outputs(1790) <= not a or b;
    layer6_outputs(1791) <= not (a xor b);
    layer6_outputs(1792) <= not b;
    layer6_outputs(1793) <= not b or a;
    layer6_outputs(1794) <= not a;
    layer6_outputs(1795) <= not (a or b);
    layer6_outputs(1796) <= a xor b;
    layer6_outputs(1797) <= a and b;
    layer6_outputs(1798) <= a and not b;
    layer6_outputs(1799) <= '0';
    layer6_outputs(1800) <= a;
    layer6_outputs(1801) <= not a;
    layer6_outputs(1802) <= not a;
    layer6_outputs(1803) <= not a;
    layer6_outputs(1804) <= a;
    layer6_outputs(1805) <= a and b;
    layer6_outputs(1806) <= '1';
    layer6_outputs(1807) <= b;
    layer6_outputs(1808) <= not a;
    layer6_outputs(1809) <= a;
    layer6_outputs(1810) <= not a;
    layer6_outputs(1811) <= a;
    layer6_outputs(1812) <= a and b;
    layer6_outputs(1813) <= a and not b;
    layer6_outputs(1814) <= not (a and b);
    layer6_outputs(1815) <= not a;
    layer6_outputs(1816) <= not a;
    layer6_outputs(1817) <= not a;
    layer6_outputs(1818) <= a xor b;
    layer6_outputs(1819) <= a and not b;
    layer6_outputs(1820) <= b and not a;
    layer6_outputs(1821) <= not (a xor b);
    layer6_outputs(1822) <= not b;
    layer6_outputs(1823) <= a xor b;
    layer6_outputs(1824) <= a;
    layer6_outputs(1825) <= a;
    layer6_outputs(1826) <= b;
    layer6_outputs(1827) <= not (a and b);
    layer6_outputs(1828) <= not a;
    layer6_outputs(1829) <= a xor b;
    layer6_outputs(1830) <= not b or a;
    layer6_outputs(1831) <= a xor b;
    layer6_outputs(1832) <= a and b;
    layer6_outputs(1833) <= a xor b;
    layer6_outputs(1834) <= not a or b;
    layer6_outputs(1835) <= a and not b;
    layer6_outputs(1836) <= a;
    layer6_outputs(1837) <= a and b;
    layer6_outputs(1838) <= a;
    layer6_outputs(1839) <= not (a and b);
    layer6_outputs(1840) <= not a;
    layer6_outputs(1841) <= a;
    layer6_outputs(1842) <= a or b;
    layer6_outputs(1843) <= a and b;
    layer6_outputs(1844) <= a or b;
    layer6_outputs(1845) <= not (a or b);
    layer6_outputs(1846) <= not b;
    layer6_outputs(1847) <= b;
    layer6_outputs(1848) <= not (a or b);
    layer6_outputs(1849) <= not b;
    layer6_outputs(1850) <= not a;
    layer6_outputs(1851) <= a;
    layer6_outputs(1852) <= not b;
    layer6_outputs(1853) <= a and not b;
    layer6_outputs(1854) <= a and b;
    layer6_outputs(1855) <= not (a xor b);
    layer6_outputs(1856) <= b;
    layer6_outputs(1857) <= not b;
    layer6_outputs(1858) <= not (a and b);
    layer6_outputs(1859) <= a or b;
    layer6_outputs(1860) <= not a;
    layer6_outputs(1861) <= not b;
    layer6_outputs(1862) <= a and not b;
    layer6_outputs(1863) <= b and not a;
    layer6_outputs(1864) <= not (a xor b);
    layer6_outputs(1865) <= a or b;
    layer6_outputs(1866) <= not (a and b);
    layer6_outputs(1867) <= a;
    layer6_outputs(1868) <= not b;
    layer6_outputs(1869) <= not a;
    layer6_outputs(1870) <= not a or b;
    layer6_outputs(1871) <= not (a xor b);
    layer6_outputs(1872) <= '0';
    layer6_outputs(1873) <= a or b;
    layer6_outputs(1874) <= b;
    layer6_outputs(1875) <= '0';
    layer6_outputs(1876) <= not b or a;
    layer6_outputs(1877) <= not b or a;
    layer6_outputs(1878) <= not b;
    layer6_outputs(1879) <= not a or b;
    layer6_outputs(1880) <= not a;
    layer6_outputs(1881) <= not b;
    layer6_outputs(1882) <= not (a or b);
    layer6_outputs(1883) <= not a;
    layer6_outputs(1884) <= a and b;
    layer6_outputs(1885) <= not a;
    layer6_outputs(1886) <= a or b;
    layer6_outputs(1887) <= not a;
    layer6_outputs(1888) <= not b;
    layer6_outputs(1889) <= not a;
    layer6_outputs(1890) <= a xor b;
    layer6_outputs(1891) <= not b;
    layer6_outputs(1892) <= a;
    layer6_outputs(1893) <= a xor b;
    layer6_outputs(1894) <= a;
    layer6_outputs(1895) <= not (a and b);
    layer6_outputs(1896) <= a xor b;
    layer6_outputs(1897) <= not (a and b);
    layer6_outputs(1898) <= not a;
    layer6_outputs(1899) <= not (a or b);
    layer6_outputs(1900) <= not (a and b);
    layer6_outputs(1901) <= a and not b;
    layer6_outputs(1902) <= a;
    layer6_outputs(1903) <= not (a xor b);
    layer6_outputs(1904) <= not (a or b);
    layer6_outputs(1905) <= not a;
    layer6_outputs(1906) <= not b;
    layer6_outputs(1907) <= b;
    layer6_outputs(1908) <= a and b;
    layer6_outputs(1909) <= b and not a;
    layer6_outputs(1910) <= not a;
    layer6_outputs(1911) <= not a;
    layer6_outputs(1912) <= a;
    layer6_outputs(1913) <= not a;
    layer6_outputs(1914) <= a;
    layer6_outputs(1915) <= a;
    layer6_outputs(1916) <= not a or b;
    layer6_outputs(1917) <= not b or a;
    layer6_outputs(1918) <= not a or b;
    layer6_outputs(1919) <= a and b;
    layer6_outputs(1920) <= not a or b;
    layer6_outputs(1921) <= not (a and b);
    layer6_outputs(1922) <= b and not a;
    layer6_outputs(1923) <= b;
    layer6_outputs(1924) <= not a;
    layer6_outputs(1925) <= a xor b;
    layer6_outputs(1926) <= a;
    layer6_outputs(1927) <= not a or b;
    layer6_outputs(1928) <= not a;
    layer6_outputs(1929) <= not (a xor b);
    layer6_outputs(1930) <= a and not b;
    layer6_outputs(1931) <= a or b;
    layer6_outputs(1932) <= not a or b;
    layer6_outputs(1933) <= not (a and b);
    layer6_outputs(1934) <= a and not b;
    layer6_outputs(1935) <= b and not a;
    layer6_outputs(1936) <= a and not b;
    layer6_outputs(1937) <= a;
    layer6_outputs(1938) <= a or b;
    layer6_outputs(1939) <= not b or a;
    layer6_outputs(1940) <= a xor b;
    layer6_outputs(1941) <= not b;
    layer6_outputs(1942) <= a xor b;
    layer6_outputs(1943) <= not (a or b);
    layer6_outputs(1944) <= not b;
    layer6_outputs(1945) <= b;
    layer6_outputs(1946) <= a;
    layer6_outputs(1947) <= b;
    layer6_outputs(1948) <= not (a and b);
    layer6_outputs(1949) <= a and b;
    layer6_outputs(1950) <= not a;
    layer6_outputs(1951) <= not a;
    layer6_outputs(1952) <= b;
    layer6_outputs(1953) <= b;
    layer6_outputs(1954) <= '1';
    layer6_outputs(1955) <= not b or a;
    layer6_outputs(1956) <= a;
    layer6_outputs(1957) <= not (a and b);
    layer6_outputs(1958) <= a and not b;
    layer6_outputs(1959) <= a xor b;
    layer6_outputs(1960) <= b;
    layer6_outputs(1961) <= not a;
    layer6_outputs(1962) <= not (a or b);
    layer6_outputs(1963) <= not a;
    layer6_outputs(1964) <= b;
    layer6_outputs(1965) <= not (a and b);
    layer6_outputs(1966) <= not (a or b);
    layer6_outputs(1967) <= not a or b;
    layer6_outputs(1968) <= not a;
    layer6_outputs(1969) <= a;
    layer6_outputs(1970) <= '0';
    layer6_outputs(1971) <= a or b;
    layer6_outputs(1972) <= not a or b;
    layer6_outputs(1973) <= not b;
    layer6_outputs(1974) <= not b or a;
    layer6_outputs(1975) <= b and not a;
    layer6_outputs(1976) <= not b;
    layer6_outputs(1977) <= not (a and b);
    layer6_outputs(1978) <= a xor b;
    layer6_outputs(1979) <= not a;
    layer6_outputs(1980) <= not (a xor b);
    layer6_outputs(1981) <= not (a and b);
    layer6_outputs(1982) <= not a;
    layer6_outputs(1983) <= a;
    layer6_outputs(1984) <= not b;
    layer6_outputs(1985) <= not a or b;
    layer6_outputs(1986) <= not a or b;
    layer6_outputs(1987) <= a;
    layer6_outputs(1988) <= '0';
    layer6_outputs(1989) <= a and b;
    layer6_outputs(1990) <= not b;
    layer6_outputs(1991) <= a;
    layer6_outputs(1992) <= b and not a;
    layer6_outputs(1993) <= not a;
    layer6_outputs(1994) <= a;
    layer6_outputs(1995) <= b;
    layer6_outputs(1996) <= b and not a;
    layer6_outputs(1997) <= a and not b;
    layer6_outputs(1998) <= a xor b;
    layer6_outputs(1999) <= b;
    layer6_outputs(2000) <= b and not a;
    layer6_outputs(2001) <= b and not a;
    layer6_outputs(2002) <= not (a and b);
    layer6_outputs(2003) <= b;
    layer6_outputs(2004) <= '1';
    layer6_outputs(2005) <= b;
    layer6_outputs(2006) <= a;
    layer6_outputs(2007) <= a xor b;
    layer6_outputs(2008) <= a and b;
    layer6_outputs(2009) <= a and not b;
    layer6_outputs(2010) <= a or b;
    layer6_outputs(2011) <= not a;
    layer6_outputs(2012) <= not b;
    layer6_outputs(2013) <= a and b;
    layer6_outputs(2014) <= a;
    layer6_outputs(2015) <= a;
    layer6_outputs(2016) <= not a;
    layer6_outputs(2017) <= a xor b;
    layer6_outputs(2018) <= a and b;
    layer6_outputs(2019) <= not b;
    layer6_outputs(2020) <= b;
    layer6_outputs(2021) <= not (a and b);
    layer6_outputs(2022) <= not b;
    layer6_outputs(2023) <= not (a or b);
    layer6_outputs(2024) <= not b;
    layer6_outputs(2025) <= a or b;
    layer6_outputs(2026) <= not a;
    layer6_outputs(2027) <= b and not a;
    layer6_outputs(2028) <= b and not a;
    layer6_outputs(2029) <= not b or a;
    layer6_outputs(2030) <= not (a and b);
    layer6_outputs(2031) <= b;
    layer6_outputs(2032) <= not (a or b);
    layer6_outputs(2033) <= a or b;
    layer6_outputs(2034) <= b and not a;
    layer6_outputs(2035) <= b;
    layer6_outputs(2036) <= not (a or b);
    layer6_outputs(2037) <= not a or b;
    layer6_outputs(2038) <= b;
    layer6_outputs(2039) <= a xor b;
    layer6_outputs(2040) <= a or b;
    layer6_outputs(2041) <= b;
    layer6_outputs(2042) <= not (a and b);
    layer6_outputs(2043) <= not a or b;
    layer6_outputs(2044) <= a xor b;
    layer6_outputs(2045) <= a;
    layer6_outputs(2046) <= a and b;
    layer6_outputs(2047) <= not (a and b);
    layer6_outputs(2048) <= not b or a;
    layer6_outputs(2049) <= not b or a;
    layer6_outputs(2050) <= b;
    layer6_outputs(2051) <= b and not a;
    layer6_outputs(2052) <= b;
    layer6_outputs(2053) <= not a;
    layer6_outputs(2054) <= b;
    layer6_outputs(2055) <= b;
    layer6_outputs(2056) <= a xor b;
    layer6_outputs(2057) <= a and not b;
    layer6_outputs(2058) <= b;
    layer6_outputs(2059) <= a and not b;
    layer6_outputs(2060) <= not a or b;
    layer6_outputs(2061) <= b;
    layer6_outputs(2062) <= a and not b;
    layer6_outputs(2063) <= b;
    layer6_outputs(2064) <= a;
    layer6_outputs(2065) <= a xor b;
    layer6_outputs(2066) <= not a;
    layer6_outputs(2067) <= a or b;
    layer6_outputs(2068) <= a;
    layer6_outputs(2069) <= a and not b;
    layer6_outputs(2070) <= not (a or b);
    layer6_outputs(2071) <= a or b;
    layer6_outputs(2072) <= not a or b;
    layer6_outputs(2073) <= b and not a;
    layer6_outputs(2074) <= a and b;
    layer6_outputs(2075) <= b;
    layer6_outputs(2076) <= not a;
    layer6_outputs(2077) <= '0';
    layer6_outputs(2078) <= a and b;
    layer6_outputs(2079) <= not (a and b);
    layer6_outputs(2080) <= '1';
    layer6_outputs(2081) <= not (a xor b);
    layer6_outputs(2082) <= not a;
    layer6_outputs(2083) <= b and not a;
    layer6_outputs(2084) <= not a or b;
    layer6_outputs(2085) <= '1';
    layer6_outputs(2086) <= a;
    layer6_outputs(2087) <= b;
    layer6_outputs(2088) <= b and not a;
    layer6_outputs(2089) <= a xor b;
    layer6_outputs(2090) <= b;
    layer6_outputs(2091) <= not (a and b);
    layer6_outputs(2092) <= not a or b;
    layer6_outputs(2093) <= b and not a;
    layer6_outputs(2094) <= not b;
    layer6_outputs(2095) <= not a;
    layer6_outputs(2096) <= not a or b;
    layer6_outputs(2097) <= not (a or b);
    layer6_outputs(2098) <= b;
    layer6_outputs(2099) <= b;
    layer6_outputs(2100) <= not (a or b);
    layer6_outputs(2101) <= not b or a;
    layer6_outputs(2102) <= '1';
    layer6_outputs(2103) <= b;
    layer6_outputs(2104) <= b;
    layer6_outputs(2105) <= b;
    layer6_outputs(2106) <= b and not a;
    layer6_outputs(2107) <= not a;
    layer6_outputs(2108) <= b;
    layer6_outputs(2109) <= not (a xor b);
    layer6_outputs(2110) <= b;
    layer6_outputs(2111) <= a and b;
    layer6_outputs(2112) <= not a;
    layer6_outputs(2113) <= a and not b;
    layer6_outputs(2114) <= not b;
    layer6_outputs(2115) <= a or b;
    layer6_outputs(2116) <= '0';
    layer6_outputs(2117) <= a;
    layer6_outputs(2118) <= b;
    layer6_outputs(2119) <= not a;
    layer6_outputs(2120) <= b;
    layer6_outputs(2121) <= a and b;
    layer6_outputs(2122) <= not b;
    layer6_outputs(2123) <= a;
    layer6_outputs(2124) <= not a;
    layer6_outputs(2125) <= not (a xor b);
    layer6_outputs(2126) <= a or b;
    layer6_outputs(2127) <= not b or a;
    layer6_outputs(2128) <= a;
    layer6_outputs(2129) <= a;
    layer6_outputs(2130) <= b and not a;
    layer6_outputs(2131) <= not b;
    layer6_outputs(2132) <= not b or a;
    layer6_outputs(2133) <= not (a xor b);
    layer6_outputs(2134) <= not b or a;
    layer6_outputs(2135) <= a xor b;
    layer6_outputs(2136) <= not a or b;
    layer6_outputs(2137) <= a or b;
    layer6_outputs(2138) <= not (a xor b);
    layer6_outputs(2139) <= a;
    layer6_outputs(2140) <= a or b;
    layer6_outputs(2141) <= a xor b;
    layer6_outputs(2142) <= b;
    layer6_outputs(2143) <= a;
    layer6_outputs(2144) <= a;
    layer6_outputs(2145) <= a and b;
    layer6_outputs(2146) <= a;
    layer6_outputs(2147) <= b;
    layer6_outputs(2148) <= not b or a;
    layer6_outputs(2149) <= b;
    layer6_outputs(2150) <= not b;
    layer6_outputs(2151) <= a or b;
    layer6_outputs(2152) <= not b or a;
    layer6_outputs(2153) <= not b or a;
    layer6_outputs(2154) <= not (a and b);
    layer6_outputs(2155) <= a;
    layer6_outputs(2156) <= not (a and b);
    layer6_outputs(2157) <= a or b;
    layer6_outputs(2158) <= not b;
    layer6_outputs(2159) <= not b or a;
    layer6_outputs(2160) <= a;
    layer6_outputs(2161) <= a or b;
    layer6_outputs(2162) <= a and not b;
    layer6_outputs(2163) <= not (a xor b);
    layer6_outputs(2164) <= not a;
    layer6_outputs(2165) <= not (a or b);
    layer6_outputs(2166) <= a and b;
    layer6_outputs(2167) <= b;
    layer6_outputs(2168) <= a xor b;
    layer6_outputs(2169) <= not a;
    layer6_outputs(2170) <= a xor b;
    layer6_outputs(2171) <= a and b;
    layer6_outputs(2172) <= not b;
    layer6_outputs(2173) <= b and not a;
    layer6_outputs(2174) <= b;
    layer6_outputs(2175) <= not a;
    layer6_outputs(2176) <= a and not b;
    layer6_outputs(2177) <= not (a and b);
    layer6_outputs(2178) <= not b;
    layer6_outputs(2179) <= a and b;
    layer6_outputs(2180) <= b;
    layer6_outputs(2181) <= a and not b;
    layer6_outputs(2182) <= b;
    layer6_outputs(2183) <= not a;
    layer6_outputs(2184) <= a;
    layer6_outputs(2185) <= not b;
    layer6_outputs(2186) <= not (a or b);
    layer6_outputs(2187) <= not a;
    layer6_outputs(2188) <= a or b;
    layer6_outputs(2189) <= not (a and b);
    layer6_outputs(2190) <= not b or a;
    layer6_outputs(2191) <= not a or b;
    layer6_outputs(2192) <= not b;
    layer6_outputs(2193) <= not (a and b);
    layer6_outputs(2194) <= not a;
    layer6_outputs(2195) <= not a;
    layer6_outputs(2196) <= not (a or b);
    layer6_outputs(2197) <= a;
    layer6_outputs(2198) <= a and not b;
    layer6_outputs(2199) <= not b;
    layer6_outputs(2200) <= a xor b;
    layer6_outputs(2201) <= not b or a;
    layer6_outputs(2202) <= b and not a;
    layer6_outputs(2203) <= a;
    layer6_outputs(2204) <= a;
    layer6_outputs(2205) <= not a;
    layer6_outputs(2206) <= not a;
    layer6_outputs(2207) <= a xor b;
    layer6_outputs(2208) <= not a or b;
    layer6_outputs(2209) <= not a;
    layer6_outputs(2210) <= a and not b;
    layer6_outputs(2211) <= a or b;
    layer6_outputs(2212) <= not b;
    layer6_outputs(2213) <= a and b;
    layer6_outputs(2214) <= not a;
    layer6_outputs(2215) <= not b;
    layer6_outputs(2216) <= not a;
    layer6_outputs(2217) <= not a;
    layer6_outputs(2218) <= '1';
    layer6_outputs(2219) <= b and not a;
    layer6_outputs(2220) <= not (a xor b);
    layer6_outputs(2221) <= not b;
    layer6_outputs(2222) <= b;
    layer6_outputs(2223) <= a xor b;
    layer6_outputs(2224) <= a;
    layer6_outputs(2225) <= a or b;
    layer6_outputs(2226) <= b;
    layer6_outputs(2227) <= not b;
    layer6_outputs(2228) <= a and not b;
    layer6_outputs(2229) <= not a;
    layer6_outputs(2230) <= not a or b;
    layer6_outputs(2231) <= a and not b;
    layer6_outputs(2232) <= not (a and b);
    layer6_outputs(2233) <= a;
    layer6_outputs(2234) <= b and not a;
    layer6_outputs(2235) <= a and b;
    layer6_outputs(2236) <= not b;
    layer6_outputs(2237) <= not a;
    layer6_outputs(2238) <= not b or a;
    layer6_outputs(2239) <= b and not a;
    layer6_outputs(2240) <= not (a and b);
    layer6_outputs(2241) <= not a;
    layer6_outputs(2242) <= b;
    layer6_outputs(2243) <= not a;
    layer6_outputs(2244) <= '1';
    layer6_outputs(2245) <= not b or a;
    layer6_outputs(2246) <= not (a and b);
    layer6_outputs(2247) <= not b;
    layer6_outputs(2248) <= not (a xor b);
    layer6_outputs(2249) <= a or b;
    layer6_outputs(2250) <= not a;
    layer6_outputs(2251) <= '1';
    layer6_outputs(2252) <= b;
    layer6_outputs(2253) <= not a or b;
    layer6_outputs(2254) <= not (a and b);
    layer6_outputs(2255) <= not b;
    layer6_outputs(2256) <= not a or b;
    layer6_outputs(2257) <= a;
    layer6_outputs(2258) <= a;
    layer6_outputs(2259) <= not (a and b);
    layer6_outputs(2260) <= a;
    layer6_outputs(2261) <= not (a xor b);
    layer6_outputs(2262) <= not (a and b);
    layer6_outputs(2263) <= not a;
    layer6_outputs(2264) <= a and b;
    layer6_outputs(2265) <= a and b;
    layer6_outputs(2266) <= b and not a;
    layer6_outputs(2267) <= a and b;
    layer6_outputs(2268) <= b and not a;
    layer6_outputs(2269) <= not a or b;
    layer6_outputs(2270) <= b;
    layer6_outputs(2271) <= not a;
    layer6_outputs(2272) <= not b;
    layer6_outputs(2273) <= '0';
    layer6_outputs(2274) <= b;
    layer6_outputs(2275) <= not b;
    layer6_outputs(2276) <= not (a xor b);
    layer6_outputs(2277) <= not (a xor b);
    layer6_outputs(2278) <= not a;
    layer6_outputs(2279) <= not a or b;
    layer6_outputs(2280) <= a or b;
    layer6_outputs(2281) <= not b;
    layer6_outputs(2282) <= not (a and b);
    layer6_outputs(2283) <= a or b;
    layer6_outputs(2284) <= not b;
    layer6_outputs(2285) <= a and b;
    layer6_outputs(2286) <= not a;
    layer6_outputs(2287) <= not (a and b);
    layer6_outputs(2288) <= b;
    layer6_outputs(2289) <= not (a and b);
    layer6_outputs(2290) <= b and not a;
    layer6_outputs(2291) <= a and not b;
    layer6_outputs(2292) <= not a;
    layer6_outputs(2293) <= not a;
    layer6_outputs(2294) <= a or b;
    layer6_outputs(2295) <= not a;
    layer6_outputs(2296) <= not b or a;
    layer6_outputs(2297) <= a and not b;
    layer6_outputs(2298) <= not b or a;
    layer6_outputs(2299) <= a and not b;
    layer6_outputs(2300) <= a xor b;
    layer6_outputs(2301) <= not a;
    layer6_outputs(2302) <= not b or a;
    layer6_outputs(2303) <= b;
    layer6_outputs(2304) <= not (a xor b);
    layer6_outputs(2305) <= not a;
    layer6_outputs(2306) <= a;
    layer6_outputs(2307) <= not (a and b);
    layer6_outputs(2308) <= not a;
    layer6_outputs(2309) <= not (a and b);
    layer6_outputs(2310) <= not a;
    layer6_outputs(2311) <= not a or b;
    layer6_outputs(2312) <= not a;
    layer6_outputs(2313) <= not a;
    layer6_outputs(2314) <= not (a and b);
    layer6_outputs(2315) <= b;
    layer6_outputs(2316) <= not a;
    layer6_outputs(2317) <= b and not a;
    layer6_outputs(2318) <= not b or a;
    layer6_outputs(2319) <= b;
    layer6_outputs(2320) <= b and not a;
    layer6_outputs(2321) <= not a;
    layer6_outputs(2322) <= a and b;
    layer6_outputs(2323) <= b;
    layer6_outputs(2324) <= not b or a;
    layer6_outputs(2325) <= not a;
    layer6_outputs(2326) <= b;
    layer6_outputs(2327) <= not a;
    layer6_outputs(2328) <= a and b;
    layer6_outputs(2329) <= '1';
    layer6_outputs(2330) <= not a or b;
    layer6_outputs(2331) <= not a or b;
    layer6_outputs(2332) <= not b;
    layer6_outputs(2333) <= not (a or b);
    layer6_outputs(2334) <= '1';
    layer6_outputs(2335) <= not b;
    layer6_outputs(2336) <= not b or a;
    layer6_outputs(2337) <= not a;
    layer6_outputs(2338) <= a and not b;
    layer6_outputs(2339) <= not (a and b);
    layer6_outputs(2340) <= a;
    layer6_outputs(2341) <= b;
    layer6_outputs(2342) <= not a or b;
    layer6_outputs(2343) <= a or b;
    layer6_outputs(2344) <= b and not a;
    layer6_outputs(2345) <= b and not a;
    layer6_outputs(2346) <= not b or a;
    layer6_outputs(2347) <= b;
    layer6_outputs(2348) <= '0';
    layer6_outputs(2349) <= b;
    layer6_outputs(2350) <= not a or b;
    layer6_outputs(2351) <= not (a or b);
    layer6_outputs(2352) <= a and not b;
    layer6_outputs(2353) <= b and not a;
    layer6_outputs(2354) <= not (a or b);
    layer6_outputs(2355) <= '0';
    layer6_outputs(2356) <= a;
    layer6_outputs(2357) <= not a;
    layer6_outputs(2358) <= not (a or b);
    layer6_outputs(2359) <= b;
    layer6_outputs(2360) <= b and not a;
    layer6_outputs(2361) <= not a;
    layer6_outputs(2362) <= not a;
    layer6_outputs(2363) <= b;
    layer6_outputs(2364) <= a xor b;
    layer6_outputs(2365) <= not b;
    layer6_outputs(2366) <= a and b;
    layer6_outputs(2367) <= not a or b;
    layer6_outputs(2368) <= a and not b;
    layer6_outputs(2369) <= a xor b;
    layer6_outputs(2370) <= not (a or b);
    layer6_outputs(2371) <= a;
    layer6_outputs(2372) <= a and b;
    layer6_outputs(2373) <= not a or b;
    layer6_outputs(2374) <= not (a xor b);
    layer6_outputs(2375) <= b;
    layer6_outputs(2376) <= not (a or b);
    layer6_outputs(2377) <= b;
    layer6_outputs(2378) <= a;
    layer6_outputs(2379) <= not a or b;
    layer6_outputs(2380) <= b;
    layer6_outputs(2381) <= a;
    layer6_outputs(2382) <= b;
    layer6_outputs(2383) <= a;
    layer6_outputs(2384) <= a and not b;
    layer6_outputs(2385) <= a;
    layer6_outputs(2386) <= not a;
    layer6_outputs(2387) <= not b;
    layer6_outputs(2388) <= b and not a;
    layer6_outputs(2389) <= not (a xor b);
    layer6_outputs(2390) <= not a;
    layer6_outputs(2391) <= not a or b;
    layer6_outputs(2392) <= not a;
    layer6_outputs(2393) <= not a;
    layer6_outputs(2394) <= not b;
    layer6_outputs(2395) <= b and not a;
    layer6_outputs(2396) <= not (a or b);
    layer6_outputs(2397) <= not a;
    layer6_outputs(2398) <= not (a and b);
    layer6_outputs(2399) <= not b or a;
    layer6_outputs(2400) <= not b;
    layer6_outputs(2401) <= not a;
    layer6_outputs(2402) <= not b or a;
    layer6_outputs(2403) <= not a;
    layer6_outputs(2404) <= not a or b;
    layer6_outputs(2405) <= not b;
    layer6_outputs(2406) <= not a or b;
    layer6_outputs(2407) <= b;
    layer6_outputs(2408) <= not a;
    layer6_outputs(2409) <= not (a xor b);
    layer6_outputs(2410) <= a and b;
    layer6_outputs(2411) <= a xor b;
    layer6_outputs(2412) <= not (a or b);
    layer6_outputs(2413) <= not a;
    layer6_outputs(2414) <= not (a and b);
    layer6_outputs(2415) <= not a;
    layer6_outputs(2416) <= a and b;
    layer6_outputs(2417) <= a;
    layer6_outputs(2418) <= a xor b;
    layer6_outputs(2419) <= not (a and b);
    layer6_outputs(2420) <= not (a and b);
    layer6_outputs(2421) <= not a;
    layer6_outputs(2422) <= a or b;
    layer6_outputs(2423) <= not b;
    layer6_outputs(2424) <= b;
    layer6_outputs(2425) <= not (a xor b);
    layer6_outputs(2426) <= not b;
    layer6_outputs(2427) <= b;
    layer6_outputs(2428) <= a and not b;
    layer6_outputs(2429) <= a or b;
    layer6_outputs(2430) <= not (a or b);
    layer6_outputs(2431) <= b;
    layer6_outputs(2432) <= b;
    layer6_outputs(2433) <= b;
    layer6_outputs(2434) <= not (a xor b);
    layer6_outputs(2435) <= a xor b;
    layer6_outputs(2436) <= b;
    layer6_outputs(2437) <= a;
    layer6_outputs(2438) <= not b;
    layer6_outputs(2439) <= a;
    layer6_outputs(2440) <= b;
    layer6_outputs(2441) <= b and not a;
    layer6_outputs(2442) <= a;
    layer6_outputs(2443) <= not a or b;
    layer6_outputs(2444) <= a and b;
    layer6_outputs(2445) <= a;
    layer6_outputs(2446) <= not (a and b);
    layer6_outputs(2447) <= a or b;
    layer6_outputs(2448) <= a;
    layer6_outputs(2449) <= not (a or b);
    layer6_outputs(2450) <= not a;
    layer6_outputs(2451) <= a;
    layer6_outputs(2452) <= a;
    layer6_outputs(2453) <= b and not a;
    layer6_outputs(2454) <= b;
    layer6_outputs(2455) <= not a or b;
    layer6_outputs(2456) <= b;
    layer6_outputs(2457) <= not a;
    layer6_outputs(2458) <= not b;
    layer6_outputs(2459) <= a and b;
    layer6_outputs(2460) <= not a;
    layer6_outputs(2461) <= not b;
    layer6_outputs(2462) <= a xor b;
    layer6_outputs(2463) <= a or b;
    layer6_outputs(2464) <= not (a xor b);
    layer6_outputs(2465) <= not b or a;
    layer6_outputs(2466) <= b;
    layer6_outputs(2467) <= a and not b;
    layer6_outputs(2468) <= a xor b;
    layer6_outputs(2469) <= not a or b;
    layer6_outputs(2470) <= not a;
    layer6_outputs(2471) <= not b or a;
    layer6_outputs(2472) <= not a;
    layer6_outputs(2473) <= a;
    layer6_outputs(2474) <= a or b;
    layer6_outputs(2475) <= b;
    layer6_outputs(2476) <= not b or a;
    layer6_outputs(2477) <= a;
    layer6_outputs(2478) <= b;
    layer6_outputs(2479) <= not b or a;
    layer6_outputs(2480) <= not a;
    layer6_outputs(2481) <= not b;
    layer6_outputs(2482) <= a xor b;
    layer6_outputs(2483) <= not (a and b);
    layer6_outputs(2484) <= a;
    layer6_outputs(2485) <= a xor b;
    layer6_outputs(2486) <= a xor b;
    layer6_outputs(2487) <= a and not b;
    layer6_outputs(2488) <= a xor b;
    layer6_outputs(2489) <= not b or a;
    layer6_outputs(2490) <= b;
    layer6_outputs(2491) <= a;
    layer6_outputs(2492) <= not (a or b);
    layer6_outputs(2493) <= a;
    layer6_outputs(2494) <= not (a and b);
    layer6_outputs(2495) <= not (a and b);
    layer6_outputs(2496) <= not b or a;
    layer6_outputs(2497) <= not (a xor b);
    layer6_outputs(2498) <= a xor b;
    layer6_outputs(2499) <= a xor b;
    layer6_outputs(2500) <= not b;
    layer6_outputs(2501) <= not (a and b);
    layer6_outputs(2502) <= a or b;
    layer6_outputs(2503) <= a;
    layer6_outputs(2504) <= b;
    layer6_outputs(2505) <= '0';
    layer6_outputs(2506) <= not (a and b);
    layer6_outputs(2507) <= not a;
    layer6_outputs(2508) <= a xor b;
    layer6_outputs(2509) <= b and not a;
    layer6_outputs(2510) <= a xor b;
    layer6_outputs(2511) <= b;
    layer6_outputs(2512) <= not a;
    layer6_outputs(2513) <= not a or b;
    layer6_outputs(2514) <= not b;
    layer6_outputs(2515) <= not (a or b);
    layer6_outputs(2516) <= not b;
    layer6_outputs(2517) <= not b;
    layer6_outputs(2518) <= not b;
    layer6_outputs(2519) <= b and not a;
    layer6_outputs(2520) <= not (a or b);
    layer6_outputs(2521) <= not (a and b);
    layer6_outputs(2522) <= a;
    layer6_outputs(2523) <= not (a or b);
    layer6_outputs(2524) <= b;
    layer6_outputs(2525) <= a and b;
    layer6_outputs(2526) <= not (a xor b);
    layer6_outputs(2527) <= a;
    layer6_outputs(2528) <= b and not a;
    layer6_outputs(2529) <= '0';
    layer6_outputs(2530) <= b and not a;
    layer6_outputs(2531) <= a or b;
    layer6_outputs(2532) <= not b;
    layer6_outputs(2533) <= '0';
    layer6_outputs(2534) <= a or b;
    layer6_outputs(2535) <= b;
    layer6_outputs(2536) <= a and not b;
    layer6_outputs(2537) <= not (a xor b);
    layer6_outputs(2538) <= a and b;
    layer6_outputs(2539) <= not a;
    layer6_outputs(2540) <= not (a or b);
    layer6_outputs(2541) <= not (a xor b);
    layer6_outputs(2542) <= a and b;
    layer6_outputs(2543) <= a;
    layer6_outputs(2544) <= a and not b;
    layer6_outputs(2545) <= not a;
    layer6_outputs(2546) <= a;
    layer6_outputs(2547) <= a;
    layer6_outputs(2548) <= a and not b;
    layer6_outputs(2549) <= not a;
    layer6_outputs(2550) <= not (a xor b);
    layer6_outputs(2551) <= not (a or b);
    layer6_outputs(2552) <= not (a and b);
    layer6_outputs(2553) <= not b;
    layer6_outputs(2554) <= b and not a;
    layer6_outputs(2555) <= not b;
    layer6_outputs(2556) <= a and not b;
    layer6_outputs(2557) <= b and not a;
    layer6_outputs(2558) <= a or b;
    layer6_outputs(2559) <= not b;
    layer6_outputs(2560) <= not (a and b);
    layer6_outputs(2561) <= not (a and b);
    layer6_outputs(2562) <= not a;
    layer6_outputs(2563) <= not a;
    layer6_outputs(2564) <= '0';
    layer6_outputs(2565) <= not a;
    layer6_outputs(2566) <= a;
    layer6_outputs(2567) <= not (a or b);
    layer6_outputs(2568) <= b and not a;
    layer6_outputs(2569) <= not b;
    layer6_outputs(2570) <= not a;
    layer6_outputs(2571) <= a and b;
    layer6_outputs(2572) <= a and not b;
    layer6_outputs(2573) <= not b;
    layer6_outputs(2574) <= b;
    layer6_outputs(2575) <= b and not a;
    layer6_outputs(2576) <= b and not a;
    layer6_outputs(2577) <= a and b;
    layer6_outputs(2578) <= not b;
    layer6_outputs(2579) <= a and b;
    layer6_outputs(2580) <= b and not a;
    layer6_outputs(2581) <= a;
    layer6_outputs(2582) <= not (a and b);
    layer6_outputs(2583) <= a and not b;
    layer6_outputs(2584) <= a or b;
    layer6_outputs(2585) <= a and not b;
    layer6_outputs(2586) <= not (a and b);
    layer6_outputs(2587) <= not a;
    layer6_outputs(2588) <= b;
    layer6_outputs(2589) <= a or b;
    layer6_outputs(2590) <= b;
    layer6_outputs(2591) <= not (a xor b);
    layer6_outputs(2592) <= a;
    layer6_outputs(2593) <= b;
    layer6_outputs(2594) <= '0';
    layer6_outputs(2595) <= a and b;
    layer6_outputs(2596) <= b;
    layer6_outputs(2597) <= b;
    layer6_outputs(2598) <= a and not b;
    layer6_outputs(2599) <= not b or a;
    layer6_outputs(2600) <= not b;
    layer6_outputs(2601) <= a;
    layer6_outputs(2602) <= a and b;
    layer6_outputs(2603) <= not b;
    layer6_outputs(2604) <= not (a and b);
    layer6_outputs(2605) <= b;
    layer6_outputs(2606) <= not a or b;
    layer6_outputs(2607) <= not b;
    layer6_outputs(2608) <= b and not a;
    layer6_outputs(2609) <= not b or a;
    layer6_outputs(2610) <= a and not b;
    layer6_outputs(2611) <= a xor b;
    layer6_outputs(2612) <= b and not a;
    layer6_outputs(2613) <= b;
    layer6_outputs(2614) <= a xor b;
    layer6_outputs(2615) <= a or b;
    layer6_outputs(2616) <= not b or a;
    layer6_outputs(2617) <= a and b;
    layer6_outputs(2618) <= a and not b;
    layer6_outputs(2619) <= a xor b;
    layer6_outputs(2620) <= b;
    layer6_outputs(2621) <= a;
    layer6_outputs(2622) <= not b;
    layer6_outputs(2623) <= not a;
    layer6_outputs(2624) <= a xor b;
    layer6_outputs(2625) <= not a;
    layer6_outputs(2626) <= not (a and b);
    layer6_outputs(2627) <= not b or a;
    layer6_outputs(2628) <= not b;
    layer6_outputs(2629) <= a;
    layer6_outputs(2630) <= not (a and b);
    layer6_outputs(2631) <= not b;
    layer6_outputs(2632) <= not a;
    layer6_outputs(2633) <= not (a or b);
    layer6_outputs(2634) <= a;
    layer6_outputs(2635) <= a;
    layer6_outputs(2636) <= a;
    layer6_outputs(2637) <= a and b;
    layer6_outputs(2638) <= not b;
    layer6_outputs(2639) <= not a;
    layer6_outputs(2640) <= a and b;
    layer6_outputs(2641) <= a or b;
    layer6_outputs(2642) <= a;
    layer6_outputs(2643) <= a;
    layer6_outputs(2644) <= a;
    layer6_outputs(2645) <= a and not b;
    layer6_outputs(2646) <= not b;
    layer6_outputs(2647) <= not b;
    layer6_outputs(2648) <= a xor b;
    layer6_outputs(2649) <= not b;
    layer6_outputs(2650) <= not (a xor b);
    layer6_outputs(2651) <= b and not a;
    layer6_outputs(2652) <= not (a and b);
    layer6_outputs(2653) <= not (a xor b);
    layer6_outputs(2654) <= b;
    layer6_outputs(2655) <= a xor b;
    layer6_outputs(2656) <= b;
    layer6_outputs(2657) <= not a;
    layer6_outputs(2658) <= a and b;
    layer6_outputs(2659) <= not a or b;
    layer6_outputs(2660) <= a and b;
    layer6_outputs(2661) <= a;
    layer6_outputs(2662) <= not (a or b);
    layer6_outputs(2663) <= a and b;
    layer6_outputs(2664) <= b and not a;
    layer6_outputs(2665) <= b and not a;
    layer6_outputs(2666) <= not a;
    layer6_outputs(2667) <= not (a xor b);
    layer6_outputs(2668) <= not (a and b);
    layer6_outputs(2669) <= not (a and b);
    layer6_outputs(2670) <= not (a and b);
    layer6_outputs(2671) <= not b;
    layer6_outputs(2672) <= not (a and b);
    layer6_outputs(2673) <= b;
    layer6_outputs(2674) <= not (a and b);
    layer6_outputs(2675) <= b and not a;
    layer6_outputs(2676) <= b;
    layer6_outputs(2677) <= a and not b;
    layer6_outputs(2678) <= a xor b;
    layer6_outputs(2679) <= not (a xor b);
    layer6_outputs(2680) <= not a or b;
    layer6_outputs(2681) <= not a or b;
    layer6_outputs(2682) <= a or b;
    layer6_outputs(2683) <= '1';
    layer6_outputs(2684) <= not b or a;
    layer6_outputs(2685) <= '0';
    layer6_outputs(2686) <= not (a xor b);
    layer6_outputs(2687) <= not (a and b);
    layer6_outputs(2688) <= '1';
    layer6_outputs(2689) <= b and not a;
    layer6_outputs(2690) <= b and not a;
    layer6_outputs(2691) <= a and b;
    layer6_outputs(2692) <= b;
    layer6_outputs(2693) <= b and not a;
    layer6_outputs(2694) <= not (a and b);
    layer6_outputs(2695) <= not (a or b);
    layer6_outputs(2696) <= not b or a;
    layer6_outputs(2697) <= not a;
    layer6_outputs(2698) <= a and not b;
    layer6_outputs(2699) <= a;
    layer6_outputs(2700) <= a and b;
    layer6_outputs(2701) <= a xor b;
    layer6_outputs(2702) <= not b or a;
    layer6_outputs(2703) <= not b;
    layer6_outputs(2704) <= a;
    layer6_outputs(2705) <= a and not b;
    layer6_outputs(2706) <= not a;
    layer6_outputs(2707) <= not b;
    layer6_outputs(2708) <= b;
    layer6_outputs(2709) <= a;
    layer6_outputs(2710) <= a and not b;
    layer6_outputs(2711) <= a;
    layer6_outputs(2712) <= b;
    layer6_outputs(2713) <= a and not b;
    layer6_outputs(2714) <= not (a or b);
    layer6_outputs(2715) <= not (a and b);
    layer6_outputs(2716) <= not b;
    layer6_outputs(2717) <= not a;
    layer6_outputs(2718) <= not (a or b);
    layer6_outputs(2719) <= a and b;
    layer6_outputs(2720) <= a xor b;
    layer6_outputs(2721) <= a xor b;
    layer6_outputs(2722) <= b;
    layer6_outputs(2723) <= not a or b;
    layer6_outputs(2724) <= not a or b;
    layer6_outputs(2725) <= not a;
    layer6_outputs(2726) <= not a;
    layer6_outputs(2727) <= '1';
    layer6_outputs(2728) <= a or b;
    layer6_outputs(2729) <= not (a or b);
    layer6_outputs(2730) <= not (a or b);
    layer6_outputs(2731) <= not (a or b);
    layer6_outputs(2732) <= not a or b;
    layer6_outputs(2733) <= not b;
    layer6_outputs(2734) <= b;
    layer6_outputs(2735) <= b;
    layer6_outputs(2736) <= not (a or b);
    layer6_outputs(2737) <= not (a or b);
    layer6_outputs(2738) <= a and not b;
    layer6_outputs(2739) <= a and b;
    layer6_outputs(2740) <= a or b;
    layer6_outputs(2741) <= not (a and b);
    layer6_outputs(2742) <= not b;
    layer6_outputs(2743) <= b;
    layer6_outputs(2744) <= not b;
    layer6_outputs(2745) <= not b or a;
    layer6_outputs(2746) <= '1';
    layer6_outputs(2747) <= b and not a;
    layer6_outputs(2748) <= not (a or b);
    layer6_outputs(2749) <= not a or b;
    layer6_outputs(2750) <= not a;
    layer6_outputs(2751) <= not b or a;
    layer6_outputs(2752) <= b;
    layer6_outputs(2753) <= not b or a;
    layer6_outputs(2754) <= a;
    layer6_outputs(2755) <= not b;
    layer6_outputs(2756) <= not a;
    layer6_outputs(2757) <= not (a or b);
    layer6_outputs(2758) <= a;
    layer6_outputs(2759) <= b;
    layer6_outputs(2760) <= b;
    layer6_outputs(2761) <= not a;
    layer6_outputs(2762) <= not (a or b);
    layer6_outputs(2763) <= not (a xor b);
    layer6_outputs(2764) <= a xor b;
    layer6_outputs(2765) <= not (a and b);
    layer6_outputs(2766) <= not (a xor b);
    layer6_outputs(2767) <= not a or b;
    layer6_outputs(2768) <= a xor b;
    layer6_outputs(2769) <= b and not a;
    layer6_outputs(2770) <= b;
    layer6_outputs(2771) <= not (a xor b);
    layer6_outputs(2772) <= not b or a;
    layer6_outputs(2773) <= not (a and b);
    layer6_outputs(2774) <= not (a or b);
    layer6_outputs(2775) <= a and not b;
    layer6_outputs(2776) <= not a;
    layer6_outputs(2777) <= not (a or b);
    layer6_outputs(2778) <= b and not a;
    layer6_outputs(2779) <= a;
    layer6_outputs(2780) <= '1';
    layer6_outputs(2781) <= b and not a;
    layer6_outputs(2782) <= '0';
    layer6_outputs(2783) <= b and not a;
    layer6_outputs(2784) <= b;
    layer6_outputs(2785) <= a;
    layer6_outputs(2786) <= '0';
    layer6_outputs(2787) <= not a or b;
    layer6_outputs(2788) <= not b;
    layer6_outputs(2789) <= not a;
    layer6_outputs(2790) <= not b;
    layer6_outputs(2791) <= b;
    layer6_outputs(2792) <= not (a and b);
    layer6_outputs(2793) <= not a or b;
    layer6_outputs(2794) <= a;
    layer6_outputs(2795) <= a xor b;
    layer6_outputs(2796) <= not (a or b);
    layer6_outputs(2797) <= a and b;
    layer6_outputs(2798) <= not a or b;
    layer6_outputs(2799) <= not a or b;
    layer6_outputs(2800) <= not b;
    layer6_outputs(2801) <= not (a or b);
    layer6_outputs(2802) <= not a;
    layer6_outputs(2803) <= '1';
    layer6_outputs(2804) <= not b;
    layer6_outputs(2805) <= a and b;
    layer6_outputs(2806) <= a;
    layer6_outputs(2807) <= not a;
    layer6_outputs(2808) <= not (a xor b);
    layer6_outputs(2809) <= not a;
    layer6_outputs(2810) <= a and not b;
    layer6_outputs(2811) <= b;
    layer6_outputs(2812) <= '0';
    layer6_outputs(2813) <= not (a xor b);
    layer6_outputs(2814) <= not b or a;
    layer6_outputs(2815) <= b and not a;
    layer6_outputs(2816) <= '1';
    layer6_outputs(2817) <= not b;
    layer6_outputs(2818) <= not (a and b);
    layer6_outputs(2819) <= '1';
    layer6_outputs(2820) <= b;
    layer6_outputs(2821) <= a;
    layer6_outputs(2822) <= not b;
    layer6_outputs(2823) <= b and not a;
    layer6_outputs(2824) <= a and b;
    layer6_outputs(2825) <= a and not b;
    layer6_outputs(2826) <= not (a and b);
    layer6_outputs(2827) <= a xor b;
    layer6_outputs(2828) <= not b;
    layer6_outputs(2829) <= not a;
    layer6_outputs(2830) <= not (a or b);
    layer6_outputs(2831) <= a or b;
    layer6_outputs(2832) <= not a;
    layer6_outputs(2833) <= not a;
    layer6_outputs(2834) <= not (a xor b);
    layer6_outputs(2835) <= not a or b;
    layer6_outputs(2836) <= a and not b;
    layer6_outputs(2837) <= b and not a;
    layer6_outputs(2838) <= not (a or b);
    layer6_outputs(2839) <= not a;
    layer6_outputs(2840) <= not a;
    layer6_outputs(2841) <= not b;
    layer6_outputs(2842) <= b and not a;
    layer6_outputs(2843) <= a;
    layer6_outputs(2844) <= not (a and b);
    layer6_outputs(2845) <= not b;
    layer6_outputs(2846) <= not (a and b);
    layer6_outputs(2847) <= not (a xor b);
    layer6_outputs(2848) <= '1';
    layer6_outputs(2849) <= not b;
    layer6_outputs(2850) <= not (a xor b);
    layer6_outputs(2851) <= b and not a;
    layer6_outputs(2852) <= '0';
    layer6_outputs(2853) <= b;
    layer6_outputs(2854) <= a and not b;
    layer6_outputs(2855) <= not b or a;
    layer6_outputs(2856) <= not a;
    layer6_outputs(2857) <= not b;
    layer6_outputs(2858) <= not b;
    layer6_outputs(2859) <= not a;
    layer6_outputs(2860) <= b and not a;
    layer6_outputs(2861) <= a xor b;
    layer6_outputs(2862) <= a;
    layer6_outputs(2863) <= not (a or b);
    layer6_outputs(2864) <= a and b;
    layer6_outputs(2865) <= not b;
    layer6_outputs(2866) <= a xor b;
    layer6_outputs(2867) <= '1';
    layer6_outputs(2868) <= a or b;
    layer6_outputs(2869) <= a;
    layer6_outputs(2870) <= not b;
    layer6_outputs(2871) <= a;
    layer6_outputs(2872) <= a;
    layer6_outputs(2873) <= not (a and b);
    layer6_outputs(2874) <= a or b;
    layer6_outputs(2875) <= not a;
    layer6_outputs(2876) <= not a or b;
    layer6_outputs(2877) <= a;
    layer6_outputs(2878) <= not b or a;
    layer6_outputs(2879) <= a or b;
    layer6_outputs(2880) <= b;
    layer6_outputs(2881) <= '1';
    layer6_outputs(2882) <= not b;
    layer6_outputs(2883) <= a and b;
    layer6_outputs(2884) <= a;
    layer6_outputs(2885) <= a;
    layer6_outputs(2886) <= not a or b;
    layer6_outputs(2887) <= a xor b;
    layer6_outputs(2888) <= a and not b;
    layer6_outputs(2889) <= not a or b;
    layer6_outputs(2890) <= not (a and b);
    layer6_outputs(2891) <= a xor b;
    layer6_outputs(2892) <= a;
    layer6_outputs(2893) <= a and b;
    layer6_outputs(2894) <= not (a and b);
    layer6_outputs(2895) <= not (a xor b);
    layer6_outputs(2896) <= not (a xor b);
    layer6_outputs(2897) <= b and not a;
    layer6_outputs(2898) <= '1';
    layer6_outputs(2899) <= not b or a;
    layer6_outputs(2900) <= b and not a;
    layer6_outputs(2901) <= b;
    layer6_outputs(2902) <= a or b;
    layer6_outputs(2903) <= b and not a;
    layer6_outputs(2904) <= not (a xor b);
    layer6_outputs(2905) <= a and not b;
    layer6_outputs(2906) <= not (a and b);
    layer6_outputs(2907) <= a xor b;
    layer6_outputs(2908) <= a;
    layer6_outputs(2909) <= not a;
    layer6_outputs(2910) <= b;
    layer6_outputs(2911) <= b and not a;
    layer6_outputs(2912) <= not a or b;
    layer6_outputs(2913) <= not a;
    layer6_outputs(2914) <= b;
    layer6_outputs(2915) <= not b or a;
    layer6_outputs(2916) <= not a;
    layer6_outputs(2917) <= a and not b;
    layer6_outputs(2918) <= not b;
    layer6_outputs(2919) <= not b;
    layer6_outputs(2920) <= a;
    layer6_outputs(2921) <= a;
    layer6_outputs(2922) <= not b;
    layer6_outputs(2923) <= '1';
    layer6_outputs(2924) <= not (a or b);
    layer6_outputs(2925) <= not (a and b);
    layer6_outputs(2926) <= b;
    layer6_outputs(2927) <= not a;
    layer6_outputs(2928) <= a;
    layer6_outputs(2929) <= a xor b;
    layer6_outputs(2930) <= not b or a;
    layer6_outputs(2931) <= not (a or b);
    layer6_outputs(2932) <= a;
    layer6_outputs(2933) <= not (a or b);
    layer6_outputs(2934) <= not b or a;
    layer6_outputs(2935) <= a and b;
    layer6_outputs(2936) <= not a;
    layer6_outputs(2937) <= not a;
    layer6_outputs(2938) <= b;
    layer6_outputs(2939) <= not a or b;
    layer6_outputs(2940) <= a and not b;
    layer6_outputs(2941) <= not b or a;
    layer6_outputs(2942) <= a;
    layer6_outputs(2943) <= not b;
    layer6_outputs(2944) <= not b or a;
    layer6_outputs(2945) <= '1';
    layer6_outputs(2946) <= b and not a;
    layer6_outputs(2947) <= not b;
    layer6_outputs(2948) <= a and not b;
    layer6_outputs(2949) <= not b;
    layer6_outputs(2950) <= not a or b;
    layer6_outputs(2951) <= not (a xor b);
    layer6_outputs(2952) <= not (a or b);
    layer6_outputs(2953) <= '1';
    layer6_outputs(2954) <= a xor b;
    layer6_outputs(2955) <= '1';
    layer6_outputs(2956) <= a and b;
    layer6_outputs(2957) <= not b or a;
    layer6_outputs(2958) <= b;
    layer6_outputs(2959) <= b;
    layer6_outputs(2960) <= a and not b;
    layer6_outputs(2961) <= not a;
    layer6_outputs(2962) <= not (a or b);
    layer6_outputs(2963) <= not b;
    layer6_outputs(2964) <= a xor b;
    layer6_outputs(2965) <= b and not a;
    layer6_outputs(2966) <= not (a and b);
    layer6_outputs(2967) <= not b;
    layer6_outputs(2968) <= a;
    layer6_outputs(2969) <= b and not a;
    layer6_outputs(2970) <= a and not b;
    layer6_outputs(2971) <= not (a or b);
    layer6_outputs(2972) <= not b;
    layer6_outputs(2973) <= b;
    layer6_outputs(2974) <= not a;
    layer6_outputs(2975) <= b and not a;
    layer6_outputs(2976) <= not b or a;
    layer6_outputs(2977) <= not (a and b);
    layer6_outputs(2978) <= not a;
    layer6_outputs(2979) <= a xor b;
    layer6_outputs(2980) <= a xor b;
    layer6_outputs(2981) <= not a;
    layer6_outputs(2982) <= not (a and b);
    layer6_outputs(2983) <= b;
    layer6_outputs(2984) <= b and not a;
    layer6_outputs(2985) <= a and not b;
    layer6_outputs(2986) <= not (a and b);
    layer6_outputs(2987) <= b and not a;
    layer6_outputs(2988) <= not (a or b);
    layer6_outputs(2989) <= not (a xor b);
    layer6_outputs(2990) <= a;
    layer6_outputs(2991) <= b and not a;
    layer6_outputs(2992) <= a;
    layer6_outputs(2993) <= a xor b;
    layer6_outputs(2994) <= b;
    layer6_outputs(2995) <= not (a or b);
    layer6_outputs(2996) <= not a;
    layer6_outputs(2997) <= a xor b;
    layer6_outputs(2998) <= b and not a;
    layer6_outputs(2999) <= not (a and b);
    layer6_outputs(3000) <= '1';
    layer6_outputs(3001) <= not b;
    layer6_outputs(3002) <= not b or a;
    layer6_outputs(3003) <= not (a xor b);
    layer6_outputs(3004) <= a xor b;
    layer6_outputs(3005) <= not b;
    layer6_outputs(3006) <= b;
    layer6_outputs(3007) <= '1';
    layer6_outputs(3008) <= b;
    layer6_outputs(3009) <= a and not b;
    layer6_outputs(3010) <= b;
    layer6_outputs(3011) <= a;
    layer6_outputs(3012) <= not b or a;
    layer6_outputs(3013) <= b;
    layer6_outputs(3014) <= a;
    layer6_outputs(3015) <= not (a xor b);
    layer6_outputs(3016) <= not b;
    layer6_outputs(3017) <= a;
    layer6_outputs(3018) <= a and b;
    layer6_outputs(3019) <= a or b;
    layer6_outputs(3020) <= not a;
    layer6_outputs(3021) <= not a;
    layer6_outputs(3022) <= not a or b;
    layer6_outputs(3023) <= b and not a;
    layer6_outputs(3024) <= not (a and b);
    layer6_outputs(3025) <= b;
    layer6_outputs(3026) <= not b;
    layer6_outputs(3027) <= not b or a;
    layer6_outputs(3028) <= not (a and b);
    layer6_outputs(3029) <= not b;
    layer6_outputs(3030) <= a or b;
    layer6_outputs(3031) <= not (a and b);
    layer6_outputs(3032) <= not (a or b);
    layer6_outputs(3033) <= not b or a;
    layer6_outputs(3034) <= not b or a;
    layer6_outputs(3035) <= a;
    layer6_outputs(3036) <= a;
    layer6_outputs(3037) <= a;
    layer6_outputs(3038) <= a or b;
    layer6_outputs(3039) <= not (a xor b);
    layer6_outputs(3040) <= not a;
    layer6_outputs(3041) <= not (a xor b);
    layer6_outputs(3042) <= b and not a;
    layer6_outputs(3043) <= not a or b;
    layer6_outputs(3044) <= not b;
    layer6_outputs(3045) <= not a;
    layer6_outputs(3046) <= not (a xor b);
    layer6_outputs(3047) <= not a;
    layer6_outputs(3048) <= not (a and b);
    layer6_outputs(3049) <= a and not b;
    layer6_outputs(3050) <= b and not a;
    layer6_outputs(3051) <= '0';
    layer6_outputs(3052) <= b and not a;
    layer6_outputs(3053) <= not a;
    layer6_outputs(3054) <= not a;
    layer6_outputs(3055) <= b;
    layer6_outputs(3056) <= not (a and b);
    layer6_outputs(3057) <= not a;
    layer6_outputs(3058) <= a;
    layer6_outputs(3059) <= not b;
    layer6_outputs(3060) <= not a;
    layer6_outputs(3061) <= not b;
    layer6_outputs(3062) <= b;
    layer6_outputs(3063) <= not a or b;
    layer6_outputs(3064) <= not b;
    layer6_outputs(3065) <= not (a and b);
    layer6_outputs(3066) <= a and not b;
    layer6_outputs(3067) <= not b;
    layer6_outputs(3068) <= a xor b;
    layer6_outputs(3069) <= b;
    layer6_outputs(3070) <= not b;
    layer6_outputs(3071) <= a and not b;
    layer6_outputs(3072) <= not (a or b);
    layer6_outputs(3073) <= a or b;
    layer6_outputs(3074) <= b and not a;
    layer6_outputs(3075) <= not (a xor b);
    layer6_outputs(3076) <= a;
    layer6_outputs(3077) <= not (a or b);
    layer6_outputs(3078) <= not (a or b);
    layer6_outputs(3079) <= not (a xor b);
    layer6_outputs(3080) <= a or b;
    layer6_outputs(3081) <= not a;
    layer6_outputs(3082) <= not b;
    layer6_outputs(3083) <= '0';
    layer6_outputs(3084) <= not a;
    layer6_outputs(3085) <= b and not a;
    layer6_outputs(3086) <= not a;
    layer6_outputs(3087) <= b and not a;
    layer6_outputs(3088) <= not a;
    layer6_outputs(3089) <= not (a xor b);
    layer6_outputs(3090) <= not (a and b);
    layer6_outputs(3091) <= not b;
    layer6_outputs(3092) <= not (a xor b);
    layer6_outputs(3093) <= not (a or b);
    layer6_outputs(3094) <= a and not b;
    layer6_outputs(3095) <= b and not a;
    layer6_outputs(3096) <= a or b;
    layer6_outputs(3097) <= b;
    layer6_outputs(3098) <= a;
    layer6_outputs(3099) <= a xor b;
    layer6_outputs(3100) <= not (a or b);
    layer6_outputs(3101) <= a;
    layer6_outputs(3102) <= a and b;
    layer6_outputs(3103) <= a;
    layer6_outputs(3104) <= not a;
    layer6_outputs(3105) <= a;
    layer6_outputs(3106) <= a or b;
    layer6_outputs(3107) <= not a;
    layer6_outputs(3108) <= not a or b;
    layer6_outputs(3109) <= not b;
    layer6_outputs(3110) <= a and b;
    layer6_outputs(3111) <= b;
    layer6_outputs(3112) <= b;
    layer6_outputs(3113) <= not (a and b);
    layer6_outputs(3114) <= b and not a;
    layer6_outputs(3115) <= not a;
    layer6_outputs(3116) <= not b;
    layer6_outputs(3117) <= not b;
    layer6_outputs(3118) <= a xor b;
    layer6_outputs(3119) <= a xor b;
    layer6_outputs(3120) <= not b or a;
    layer6_outputs(3121) <= not (a xor b);
    layer6_outputs(3122) <= a or b;
    layer6_outputs(3123) <= not (a or b);
    layer6_outputs(3124) <= b and not a;
    layer6_outputs(3125) <= not a;
    layer6_outputs(3126) <= not (a or b);
    layer6_outputs(3127) <= not a or b;
    layer6_outputs(3128) <= b and not a;
    layer6_outputs(3129) <= not a or b;
    layer6_outputs(3130) <= not a or b;
    layer6_outputs(3131) <= not a or b;
    layer6_outputs(3132) <= a xor b;
    layer6_outputs(3133) <= b;
    layer6_outputs(3134) <= not a or b;
    layer6_outputs(3135) <= not b;
    layer6_outputs(3136) <= not (a and b);
    layer6_outputs(3137) <= not b;
    layer6_outputs(3138) <= a or b;
    layer6_outputs(3139) <= a;
    layer6_outputs(3140) <= not a;
    layer6_outputs(3141) <= b and not a;
    layer6_outputs(3142) <= not b or a;
    layer6_outputs(3143) <= a;
    layer6_outputs(3144) <= a xor b;
    layer6_outputs(3145) <= a and b;
    layer6_outputs(3146) <= not b;
    layer6_outputs(3147) <= b and not a;
    layer6_outputs(3148) <= not a;
    layer6_outputs(3149) <= not (a and b);
    layer6_outputs(3150) <= not a;
    layer6_outputs(3151) <= '1';
    layer6_outputs(3152) <= not (a xor b);
    layer6_outputs(3153) <= not b;
    layer6_outputs(3154) <= '0';
    layer6_outputs(3155) <= b;
    layer6_outputs(3156) <= not b or a;
    layer6_outputs(3157) <= a;
    layer6_outputs(3158) <= b;
    layer6_outputs(3159) <= a;
    layer6_outputs(3160) <= b and not a;
    layer6_outputs(3161) <= not b or a;
    layer6_outputs(3162) <= not a or b;
    layer6_outputs(3163) <= not (a or b);
    layer6_outputs(3164) <= not a;
    layer6_outputs(3165) <= b and not a;
    layer6_outputs(3166) <= not b;
    layer6_outputs(3167) <= not (a and b);
    layer6_outputs(3168) <= not b or a;
    layer6_outputs(3169) <= not a or b;
    layer6_outputs(3170) <= not (a xor b);
    layer6_outputs(3171) <= a or b;
    layer6_outputs(3172) <= not b;
    layer6_outputs(3173) <= not (a or b);
    layer6_outputs(3174) <= '0';
    layer6_outputs(3175) <= not b;
    layer6_outputs(3176) <= a and b;
    layer6_outputs(3177) <= a;
    layer6_outputs(3178) <= not a;
    layer6_outputs(3179) <= not (a or b);
    layer6_outputs(3180) <= b;
    layer6_outputs(3181) <= not b;
    layer6_outputs(3182) <= not b;
    layer6_outputs(3183) <= not a or b;
    layer6_outputs(3184) <= a or b;
    layer6_outputs(3185) <= a and not b;
    layer6_outputs(3186) <= not b;
    layer6_outputs(3187) <= not a;
    layer6_outputs(3188) <= not b;
    layer6_outputs(3189) <= a;
    layer6_outputs(3190) <= a;
    layer6_outputs(3191) <= a and not b;
    layer6_outputs(3192) <= a and not b;
    layer6_outputs(3193) <= b and not a;
    layer6_outputs(3194) <= not (a xor b);
    layer6_outputs(3195) <= not a;
    layer6_outputs(3196) <= not b or a;
    layer6_outputs(3197) <= b;
    layer6_outputs(3198) <= a or b;
    layer6_outputs(3199) <= not (a xor b);
    layer6_outputs(3200) <= not b or a;
    layer6_outputs(3201) <= a and b;
    layer6_outputs(3202) <= not b;
    layer6_outputs(3203) <= a xor b;
    layer6_outputs(3204) <= a xor b;
    layer6_outputs(3205) <= not (a or b);
    layer6_outputs(3206) <= not b;
    layer6_outputs(3207) <= a;
    layer6_outputs(3208) <= not a;
    layer6_outputs(3209) <= not (a or b);
    layer6_outputs(3210) <= not (a or b);
    layer6_outputs(3211) <= b;
    layer6_outputs(3212) <= not b or a;
    layer6_outputs(3213) <= not (a or b);
    layer6_outputs(3214) <= a or b;
    layer6_outputs(3215) <= b;
    layer6_outputs(3216) <= not a;
    layer6_outputs(3217) <= '0';
    layer6_outputs(3218) <= b;
    layer6_outputs(3219) <= b;
    layer6_outputs(3220) <= not (a and b);
    layer6_outputs(3221) <= b;
    layer6_outputs(3222) <= not b;
    layer6_outputs(3223) <= not (a or b);
    layer6_outputs(3224) <= a;
    layer6_outputs(3225) <= a or b;
    layer6_outputs(3226) <= not a;
    layer6_outputs(3227) <= not (a and b);
    layer6_outputs(3228) <= not a or b;
    layer6_outputs(3229) <= a and b;
    layer6_outputs(3230) <= not a or b;
    layer6_outputs(3231) <= a xor b;
    layer6_outputs(3232) <= not a;
    layer6_outputs(3233) <= not a or b;
    layer6_outputs(3234) <= a and not b;
    layer6_outputs(3235) <= b and not a;
    layer6_outputs(3236) <= b;
    layer6_outputs(3237) <= not a;
    layer6_outputs(3238) <= not (a and b);
    layer6_outputs(3239) <= b and not a;
    layer6_outputs(3240) <= not a;
    layer6_outputs(3241) <= a and b;
    layer6_outputs(3242) <= not b;
    layer6_outputs(3243) <= not b or a;
    layer6_outputs(3244) <= not (a xor b);
    layer6_outputs(3245) <= a or b;
    layer6_outputs(3246) <= a;
    layer6_outputs(3247) <= not b or a;
    layer6_outputs(3248) <= a or b;
    layer6_outputs(3249) <= a;
    layer6_outputs(3250) <= not b;
    layer6_outputs(3251) <= b;
    layer6_outputs(3252) <= not (a xor b);
    layer6_outputs(3253) <= a;
    layer6_outputs(3254) <= not (a or b);
    layer6_outputs(3255) <= a and b;
    layer6_outputs(3256) <= b and not a;
    layer6_outputs(3257) <= not (a xor b);
    layer6_outputs(3258) <= not (a or b);
    layer6_outputs(3259) <= not (a xor b);
    layer6_outputs(3260) <= a;
    layer6_outputs(3261) <= a or b;
    layer6_outputs(3262) <= not b;
    layer6_outputs(3263) <= a xor b;
    layer6_outputs(3264) <= a;
    layer6_outputs(3265) <= a or b;
    layer6_outputs(3266) <= not a or b;
    layer6_outputs(3267) <= a and b;
    layer6_outputs(3268) <= not a;
    layer6_outputs(3269) <= b;
    layer6_outputs(3270) <= not b;
    layer6_outputs(3271) <= not (a or b);
    layer6_outputs(3272) <= not b or a;
    layer6_outputs(3273) <= not b or a;
    layer6_outputs(3274) <= b and not a;
    layer6_outputs(3275) <= not a;
    layer6_outputs(3276) <= b and not a;
    layer6_outputs(3277) <= not (a xor b);
    layer6_outputs(3278) <= a and b;
    layer6_outputs(3279) <= a;
    layer6_outputs(3280) <= a;
    layer6_outputs(3281) <= not b or a;
    layer6_outputs(3282) <= b;
    layer6_outputs(3283) <= b;
    layer6_outputs(3284) <= a;
    layer6_outputs(3285) <= not a;
    layer6_outputs(3286) <= not (a xor b);
    layer6_outputs(3287) <= b;
    layer6_outputs(3288) <= b;
    layer6_outputs(3289) <= a xor b;
    layer6_outputs(3290) <= not b;
    layer6_outputs(3291) <= not (a or b);
    layer6_outputs(3292) <= a;
    layer6_outputs(3293) <= b and not a;
    layer6_outputs(3294) <= not a or b;
    layer6_outputs(3295) <= not (a xor b);
    layer6_outputs(3296) <= a and b;
    layer6_outputs(3297) <= a;
    layer6_outputs(3298) <= a;
    layer6_outputs(3299) <= not b;
    layer6_outputs(3300) <= a xor b;
    layer6_outputs(3301) <= not (a and b);
    layer6_outputs(3302) <= a or b;
    layer6_outputs(3303) <= not b or a;
    layer6_outputs(3304) <= b;
    layer6_outputs(3305) <= not b or a;
    layer6_outputs(3306) <= not a;
    layer6_outputs(3307) <= a;
    layer6_outputs(3308) <= '0';
    layer6_outputs(3309) <= a;
    layer6_outputs(3310) <= a or b;
    layer6_outputs(3311) <= a;
    layer6_outputs(3312) <= not b;
    layer6_outputs(3313) <= b;
    layer6_outputs(3314) <= not b;
    layer6_outputs(3315) <= '1';
    layer6_outputs(3316) <= a and b;
    layer6_outputs(3317) <= not b;
    layer6_outputs(3318) <= a or b;
    layer6_outputs(3319) <= a;
    layer6_outputs(3320) <= not a;
    layer6_outputs(3321) <= a;
    layer6_outputs(3322) <= not b or a;
    layer6_outputs(3323) <= not a or b;
    layer6_outputs(3324) <= b;
    layer6_outputs(3325) <= not b or a;
    layer6_outputs(3326) <= a;
    layer6_outputs(3327) <= not b;
    layer6_outputs(3328) <= b;
    layer6_outputs(3329) <= a and b;
    layer6_outputs(3330) <= a and not b;
    layer6_outputs(3331) <= b;
    layer6_outputs(3332) <= not a;
    layer6_outputs(3333) <= not (a and b);
    layer6_outputs(3334) <= not (a xor b);
    layer6_outputs(3335) <= not a;
    layer6_outputs(3336) <= not b or a;
    layer6_outputs(3337) <= b;
    layer6_outputs(3338) <= not (a or b);
    layer6_outputs(3339) <= a and b;
    layer6_outputs(3340) <= not a;
    layer6_outputs(3341) <= b;
    layer6_outputs(3342) <= a xor b;
    layer6_outputs(3343) <= not a or b;
    layer6_outputs(3344) <= not a;
    layer6_outputs(3345) <= a or b;
    layer6_outputs(3346) <= not (a xor b);
    layer6_outputs(3347) <= not b;
    layer6_outputs(3348) <= b;
    layer6_outputs(3349) <= a;
    layer6_outputs(3350) <= a or b;
    layer6_outputs(3351) <= a or b;
    layer6_outputs(3352) <= a and not b;
    layer6_outputs(3353) <= '0';
    layer6_outputs(3354) <= b;
    layer6_outputs(3355) <= not (a or b);
    layer6_outputs(3356) <= a;
    layer6_outputs(3357) <= a;
    layer6_outputs(3358) <= a or b;
    layer6_outputs(3359) <= a;
    layer6_outputs(3360) <= not a or b;
    layer6_outputs(3361) <= not (a and b);
    layer6_outputs(3362) <= not (a or b);
    layer6_outputs(3363) <= not b;
    layer6_outputs(3364) <= '1';
    layer6_outputs(3365) <= a xor b;
    layer6_outputs(3366) <= not a;
    layer6_outputs(3367) <= not b or a;
    layer6_outputs(3368) <= not (a or b);
    layer6_outputs(3369) <= not b;
    layer6_outputs(3370) <= b and not a;
    layer6_outputs(3371) <= '0';
    layer6_outputs(3372) <= a and b;
    layer6_outputs(3373) <= a;
    layer6_outputs(3374) <= a;
    layer6_outputs(3375) <= not b;
    layer6_outputs(3376) <= not a;
    layer6_outputs(3377) <= not b;
    layer6_outputs(3378) <= not b;
    layer6_outputs(3379) <= not b;
    layer6_outputs(3380) <= b and not a;
    layer6_outputs(3381) <= not b;
    layer6_outputs(3382) <= a;
    layer6_outputs(3383) <= b;
    layer6_outputs(3384) <= a xor b;
    layer6_outputs(3385) <= b;
    layer6_outputs(3386) <= a and b;
    layer6_outputs(3387) <= not a;
    layer6_outputs(3388) <= not a;
    layer6_outputs(3389) <= a;
    layer6_outputs(3390) <= not (a xor b);
    layer6_outputs(3391) <= a and not b;
    layer6_outputs(3392) <= not (a and b);
    layer6_outputs(3393) <= a;
    layer6_outputs(3394) <= b and not a;
    layer6_outputs(3395) <= not (a xor b);
    layer6_outputs(3396) <= '1';
    layer6_outputs(3397) <= a or b;
    layer6_outputs(3398) <= not b;
    layer6_outputs(3399) <= not a or b;
    layer6_outputs(3400) <= not b;
    layer6_outputs(3401) <= a or b;
    layer6_outputs(3402) <= a;
    layer6_outputs(3403) <= b and not a;
    layer6_outputs(3404) <= not (a and b);
    layer6_outputs(3405) <= not b;
    layer6_outputs(3406) <= not (a or b);
    layer6_outputs(3407) <= a xor b;
    layer6_outputs(3408) <= not b;
    layer6_outputs(3409) <= b and not a;
    layer6_outputs(3410) <= not a or b;
    layer6_outputs(3411) <= '0';
    layer6_outputs(3412) <= not (a and b);
    layer6_outputs(3413) <= b;
    layer6_outputs(3414) <= '1';
    layer6_outputs(3415) <= a;
    layer6_outputs(3416) <= a;
    layer6_outputs(3417) <= b;
    layer6_outputs(3418) <= b;
    layer6_outputs(3419) <= b and not a;
    layer6_outputs(3420) <= '1';
    layer6_outputs(3421) <= not a;
    layer6_outputs(3422) <= b and not a;
    layer6_outputs(3423) <= b;
    layer6_outputs(3424) <= a;
    layer6_outputs(3425) <= not a or b;
    layer6_outputs(3426) <= not (a xor b);
    layer6_outputs(3427) <= not a;
    layer6_outputs(3428) <= a or b;
    layer6_outputs(3429) <= not b;
    layer6_outputs(3430) <= not (a or b);
    layer6_outputs(3431) <= not b;
    layer6_outputs(3432) <= b;
    layer6_outputs(3433) <= not b;
    layer6_outputs(3434) <= a;
    layer6_outputs(3435) <= a xor b;
    layer6_outputs(3436) <= a;
    layer6_outputs(3437) <= a and not b;
    layer6_outputs(3438) <= not b or a;
    layer6_outputs(3439) <= a;
    layer6_outputs(3440) <= b;
    layer6_outputs(3441) <= not a or b;
    layer6_outputs(3442) <= not a;
    layer6_outputs(3443) <= b;
    layer6_outputs(3444) <= b;
    layer6_outputs(3445) <= not b;
    layer6_outputs(3446) <= not (a and b);
    layer6_outputs(3447) <= a or b;
    layer6_outputs(3448) <= not (a or b);
    layer6_outputs(3449) <= not b;
    layer6_outputs(3450) <= not b;
    layer6_outputs(3451) <= b and not a;
    layer6_outputs(3452) <= a;
    layer6_outputs(3453) <= a and b;
    layer6_outputs(3454) <= a and b;
    layer6_outputs(3455) <= a;
    layer6_outputs(3456) <= a xor b;
    layer6_outputs(3457) <= not a;
    layer6_outputs(3458) <= b;
    layer6_outputs(3459) <= not a or b;
    layer6_outputs(3460) <= '1';
    layer6_outputs(3461) <= not a;
    layer6_outputs(3462) <= not a or b;
    layer6_outputs(3463) <= a;
    layer6_outputs(3464) <= b;
    layer6_outputs(3465) <= b;
    layer6_outputs(3466) <= a and not b;
    layer6_outputs(3467) <= a or b;
    layer6_outputs(3468) <= not a;
    layer6_outputs(3469) <= not a;
    layer6_outputs(3470) <= not (a or b);
    layer6_outputs(3471) <= not b;
    layer6_outputs(3472) <= '0';
    layer6_outputs(3473) <= not a or b;
    layer6_outputs(3474) <= b and not a;
    layer6_outputs(3475) <= not a;
    layer6_outputs(3476) <= not b;
    layer6_outputs(3477) <= not a;
    layer6_outputs(3478) <= a and not b;
    layer6_outputs(3479) <= a and not b;
    layer6_outputs(3480) <= b;
    layer6_outputs(3481) <= not a;
    layer6_outputs(3482) <= not (a and b);
    layer6_outputs(3483) <= b and not a;
    layer6_outputs(3484) <= not (a and b);
    layer6_outputs(3485) <= not b;
    layer6_outputs(3486) <= b;
    layer6_outputs(3487) <= b;
    layer6_outputs(3488) <= not a;
    layer6_outputs(3489) <= a and b;
    layer6_outputs(3490) <= a and b;
    layer6_outputs(3491) <= b and not a;
    layer6_outputs(3492) <= not a or b;
    layer6_outputs(3493) <= a xor b;
    layer6_outputs(3494) <= b and not a;
    layer6_outputs(3495) <= a;
    layer6_outputs(3496) <= b and not a;
    layer6_outputs(3497) <= not a;
    layer6_outputs(3498) <= not (a or b);
    layer6_outputs(3499) <= a xor b;
    layer6_outputs(3500) <= not (a or b);
    layer6_outputs(3501) <= not b;
    layer6_outputs(3502) <= a xor b;
    layer6_outputs(3503) <= b and not a;
    layer6_outputs(3504) <= not a;
    layer6_outputs(3505) <= a or b;
    layer6_outputs(3506) <= b;
    layer6_outputs(3507) <= not b;
    layer6_outputs(3508) <= not a;
    layer6_outputs(3509) <= b;
    layer6_outputs(3510) <= not b;
    layer6_outputs(3511) <= not (a xor b);
    layer6_outputs(3512) <= not b or a;
    layer6_outputs(3513) <= a;
    layer6_outputs(3514) <= '1';
    layer6_outputs(3515) <= not b;
    layer6_outputs(3516) <= not (a xor b);
    layer6_outputs(3517) <= a xor b;
    layer6_outputs(3518) <= a;
    layer6_outputs(3519) <= not (a xor b);
    layer6_outputs(3520) <= a;
    layer6_outputs(3521) <= b;
    layer6_outputs(3522) <= not b;
    layer6_outputs(3523) <= not a;
    layer6_outputs(3524) <= a;
    layer6_outputs(3525) <= b and not a;
    layer6_outputs(3526) <= a or b;
    layer6_outputs(3527) <= not (a xor b);
    layer6_outputs(3528) <= a and not b;
    layer6_outputs(3529) <= not a or b;
    layer6_outputs(3530) <= a or b;
    layer6_outputs(3531) <= a;
    layer6_outputs(3532) <= not (a or b);
    layer6_outputs(3533) <= '1';
    layer6_outputs(3534) <= not (a and b);
    layer6_outputs(3535) <= not (a and b);
    layer6_outputs(3536) <= not b;
    layer6_outputs(3537) <= not b or a;
    layer6_outputs(3538) <= not a;
    layer6_outputs(3539) <= not b;
    layer6_outputs(3540) <= b and not a;
    layer6_outputs(3541) <= not a or b;
    layer6_outputs(3542) <= a or b;
    layer6_outputs(3543) <= a;
    layer6_outputs(3544) <= a;
    layer6_outputs(3545) <= not a;
    layer6_outputs(3546) <= not (a xor b);
    layer6_outputs(3547) <= not a;
    layer6_outputs(3548) <= b and not a;
    layer6_outputs(3549) <= not b;
    layer6_outputs(3550) <= a;
    layer6_outputs(3551) <= not a;
    layer6_outputs(3552) <= not a;
    layer6_outputs(3553) <= a xor b;
    layer6_outputs(3554) <= b;
    layer6_outputs(3555) <= not b;
    layer6_outputs(3556) <= a and not b;
    layer6_outputs(3557) <= not b or a;
    layer6_outputs(3558) <= a and b;
    layer6_outputs(3559) <= a or b;
    layer6_outputs(3560) <= not a;
    layer6_outputs(3561) <= not b or a;
    layer6_outputs(3562) <= not (a or b);
    layer6_outputs(3563) <= b;
    layer6_outputs(3564) <= a;
    layer6_outputs(3565) <= a xor b;
    layer6_outputs(3566) <= not b;
    layer6_outputs(3567) <= a or b;
    layer6_outputs(3568) <= b;
    layer6_outputs(3569) <= a xor b;
    layer6_outputs(3570) <= not a or b;
    layer6_outputs(3571) <= not b or a;
    layer6_outputs(3572) <= b;
    layer6_outputs(3573) <= not b;
    layer6_outputs(3574) <= not (a or b);
    layer6_outputs(3575) <= not (a or b);
    layer6_outputs(3576) <= b;
    layer6_outputs(3577) <= not (a or b);
    layer6_outputs(3578) <= not b;
    layer6_outputs(3579) <= not a;
    layer6_outputs(3580) <= a;
    layer6_outputs(3581) <= a and b;
    layer6_outputs(3582) <= a and b;
    layer6_outputs(3583) <= not a;
    layer6_outputs(3584) <= b and not a;
    layer6_outputs(3585) <= a and not b;
    layer6_outputs(3586) <= not a;
    layer6_outputs(3587) <= not a or b;
    layer6_outputs(3588) <= not (a and b);
    layer6_outputs(3589) <= not b;
    layer6_outputs(3590) <= not b;
    layer6_outputs(3591) <= not (a or b);
    layer6_outputs(3592) <= not a;
    layer6_outputs(3593) <= a xor b;
    layer6_outputs(3594) <= b and not a;
    layer6_outputs(3595) <= not b;
    layer6_outputs(3596) <= a and not b;
    layer6_outputs(3597) <= a xor b;
    layer6_outputs(3598) <= not (a or b);
    layer6_outputs(3599) <= not a;
    layer6_outputs(3600) <= '0';
    layer6_outputs(3601) <= not b;
    layer6_outputs(3602) <= '1';
    layer6_outputs(3603) <= not a;
    layer6_outputs(3604) <= b;
    layer6_outputs(3605) <= not b;
    layer6_outputs(3606) <= b and not a;
    layer6_outputs(3607) <= a and b;
    layer6_outputs(3608) <= not b or a;
    layer6_outputs(3609) <= not (a or b);
    layer6_outputs(3610) <= b and not a;
    layer6_outputs(3611) <= b;
    layer6_outputs(3612) <= b;
    layer6_outputs(3613) <= not (a xor b);
    layer6_outputs(3614) <= not (a or b);
    layer6_outputs(3615) <= not b or a;
    layer6_outputs(3616) <= b;
    layer6_outputs(3617) <= a and not b;
    layer6_outputs(3618) <= not a;
    layer6_outputs(3619) <= not (a xor b);
    layer6_outputs(3620) <= not a;
    layer6_outputs(3621) <= not a or b;
    layer6_outputs(3622) <= not b;
    layer6_outputs(3623) <= a and not b;
    layer6_outputs(3624) <= a;
    layer6_outputs(3625) <= a xor b;
    layer6_outputs(3626) <= a xor b;
    layer6_outputs(3627) <= not (a xor b);
    layer6_outputs(3628) <= '0';
    layer6_outputs(3629) <= a and b;
    layer6_outputs(3630) <= not b;
    layer6_outputs(3631) <= not (a and b);
    layer6_outputs(3632) <= not b;
    layer6_outputs(3633) <= a xor b;
    layer6_outputs(3634) <= b;
    layer6_outputs(3635) <= b;
    layer6_outputs(3636) <= not b;
    layer6_outputs(3637) <= a;
    layer6_outputs(3638) <= a;
    layer6_outputs(3639) <= not (a and b);
    layer6_outputs(3640) <= a xor b;
    layer6_outputs(3641) <= not (a and b);
    layer6_outputs(3642) <= not b;
    layer6_outputs(3643) <= not a or b;
    layer6_outputs(3644) <= not a;
    layer6_outputs(3645) <= not b;
    layer6_outputs(3646) <= not b;
    layer6_outputs(3647) <= a and b;
    layer6_outputs(3648) <= not b;
    layer6_outputs(3649) <= b;
    layer6_outputs(3650) <= a and b;
    layer6_outputs(3651) <= a and not b;
    layer6_outputs(3652) <= not b;
    layer6_outputs(3653) <= not a or b;
    layer6_outputs(3654) <= not a;
    layer6_outputs(3655) <= b;
    layer6_outputs(3656) <= a and not b;
    layer6_outputs(3657) <= not a or b;
    layer6_outputs(3658) <= not a;
    layer6_outputs(3659) <= not a;
    layer6_outputs(3660) <= not b;
    layer6_outputs(3661) <= b;
    layer6_outputs(3662) <= not a or b;
    layer6_outputs(3663) <= b;
    layer6_outputs(3664) <= not b;
    layer6_outputs(3665) <= not b;
    layer6_outputs(3666) <= not b;
    layer6_outputs(3667) <= not (a and b);
    layer6_outputs(3668) <= a or b;
    layer6_outputs(3669) <= not b or a;
    layer6_outputs(3670) <= not a or b;
    layer6_outputs(3671) <= not a or b;
    layer6_outputs(3672) <= not a;
    layer6_outputs(3673) <= b and not a;
    layer6_outputs(3674) <= not b;
    layer6_outputs(3675) <= a and not b;
    layer6_outputs(3676) <= not (a or b);
    layer6_outputs(3677) <= b and not a;
    layer6_outputs(3678) <= not (a xor b);
    layer6_outputs(3679) <= b;
    layer6_outputs(3680) <= a;
    layer6_outputs(3681) <= b and not a;
    layer6_outputs(3682) <= a;
    layer6_outputs(3683) <= not (a or b);
    layer6_outputs(3684) <= not b;
    layer6_outputs(3685) <= '1';
    layer6_outputs(3686) <= not (a xor b);
    layer6_outputs(3687) <= a;
    layer6_outputs(3688) <= not a or b;
    layer6_outputs(3689) <= b;
    layer6_outputs(3690) <= b;
    layer6_outputs(3691) <= b and not a;
    layer6_outputs(3692) <= a;
    layer6_outputs(3693) <= a and not b;
    layer6_outputs(3694) <= not b or a;
    layer6_outputs(3695) <= b;
    layer6_outputs(3696) <= a and not b;
    layer6_outputs(3697) <= not (a and b);
    layer6_outputs(3698) <= not a;
    layer6_outputs(3699) <= a;
    layer6_outputs(3700) <= not b or a;
    layer6_outputs(3701) <= a and not b;
    layer6_outputs(3702) <= not b;
    layer6_outputs(3703) <= not b;
    layer6_outputs(3704) <= not (a xor b);
    layer6_outputs(3705) <= a;
    layer6_outputs(3706) <= not b;
    layer6_outputs(3707) <= a;
    layer6_outputs(3708) <= not (a xor b);
    layer6_outputs(3709) <= not a or b;
    layer6_outputs(3710) <= not b;
    layer6_outputs(3711) <= a or b;
    layer6_outputs(3712) <= not (a xor b);
    layer6_outputs(3713) <= not a or b;
    layer6_outputs(3714) <= not b;
    layer6_outputs(3715) <= a;
    layer6_outputs(3716) <= b;
    layer6_outputs(3717) <= not (a xor b);
    layer6_outputs(3718) <= not (a or b);
    layer6_outputs(3719) <= not b;
    layer6_outputs(3720) <= a;
    layer6_outputs(3721) <= a;
    layer6_outputs(3722) <= not a;
    layer6_outputs(3723) <= not (a or b);
    layer6_outputs(3724) <= not (a or b);
    layer6_outputs(3725) <= a;
    layer6_outputs(3726) <= b and not a;
    layer6_outputs(3727) <= a and not b;
    layer6_outputs(3728) <= a xor b;
    layer6_outputs(3729) <= '0';
    layer6_outputs(3730) <= not a;
    layer6_outputs(3731) <= not b or a;
    layer6_outputs(3732) <= b;
    layer6_outputs(3733) <= a;
    layer6_outputs(3734) <= b;
    layer6_outputs(3735) <= '0';
    layer6_outputs(3736) <= not a;
    layer6_outputs(3737) <= a;
    layer6_outputs(3738) <= a;
    layer6_outputs(3739) <= a or b;
    layer6_outputs(3740) <= b;
    layer6_outputs(3741) <= a and not b;
    layer6_outputs(3742) <= not b;
    layer6_outputs(3743) <= a and b;
    layer6_outputs(3744) <= '0';
    layer6_outputs(3745) <= not b or a;
    layer6_outputs(3746) <= a and not b;
    layer6_outputs(3747) <= a;
    layer6_outputs(3748) <= '1';
    layer6_outputs(3749) <= not a;
    layer6_outputs(3750) <= b and not a;
    layer6_outputs(3751) <= not b;
    layer6_outputs(3752) <= b;
    layer6_outputs(3753) <= not b;
    layer6_outputs(3754) <= a or b;
    layer6_outputs(3755) <= '1';
    layer6_outputs(3756) <= b;
    layer6_outputs(3757) <= not (a xor b);
    layer6_outputs(3758) <= not (a xor b);
    layer6_outputs(3759) <= a or b;
    layer6_outputs(3760) <= not b;
    layer6_outputs(3761) <= b;
    layer6_outputs(3762) <= a;
    layer6_outputs(3763) <= not a or b;
    layer6_outputs(3764) <= not (a or b);
    layer6_outputs(3765) <= not (a xor b);
    layer6_outputs(3766) <= '0';
    layer6_outputs(3767) <= b;
    layer6_outputs(3768) <= a and not b;
    layer6_outputs(3769) <= not (a xor b);
    layer6_outputs(3770) <= b;
    layer6_outputs(3771) <= not b or a;
    layer6_outputs(3772) <= not (a and b);
    layer6_outputs(3773) <= a and b;
    layer6_outputs(3774) <= not b;
    layer6_outputs(3775) <= b;
    layer6_outputs(3776) <= a;
    layer6_outputs(3777) <= a and not b;
    layer6_outputs(3778) <= not b;
    layer6_outputs(3779) <= not b;
    layer6_outputs(3780) <= a xor b;
    layer6_outputs(3781) <= '1';
    layer6_outputs(3782) <= b;
    layer6_outputs(3783) <= a;
    layer6_outputs(3784) <= not b;
    layer6_outputs(3785) <= not a or b;
    layer6_outputs(3786) <= not b or a;
    layer6_outputs(3787) <= b;
    layer6_outputs(3788) <= a xor b;
    layer6_outputs(3789) <= a xor b;
    layer6_outputs(3790) <= a and b;
    layer6_outputs(3791) <= a;
    layer6_outputs(3792) <= a xor b;
    layer6_outputs(3793) <= a;
    layer6_outputs(3794) <= not a;
    layer6_outputs(3795) <= not b;
    layer6_outputs(3796) <= not (a or b);
    layer6_outputs(3797) <= '1';
    layer6_outputs(3798) <= not b;
    layer6_outputs(3799) <= not b or a;
    layer6_outputs(3800) <= not a or b;
    layer6_outputs(3801) <= not a or b;
    layer6_outputs(3802) <= not (a and b);
    layer6_outputs(3803) <= a;
    layer6_outputs(3804) <= not b or a;
    layer6_outputs(3805) <= a and b;
    layer6_outputs(3806) <= not b;
    layer6_outputs(3807) <= a;
    layer6_outputs(3808) <= '0';
    layer6_outputs(3809) <= not (a and b);
    layer6_outputs(3810) <= a and not b;
    layer6_outputs(3811) <= a;
    layer6_outputs(3812) <= not a or b;
    layer6_outputs(3813) <= a and not b;
    layer6_outputs(3814) <= not (a and b);
    layer6_outputs(3815) <= not b or a;
    layer6_outputs(3816) <= not b or a;
    layer6_outputs(3817) <= a;
    layer6_outputs(3818) <= a;
    layer6_outputs(3819) <= not (a xor b);
    layer6_outputs(3820) <= a and not b;
    layer6_outputs(3821) <= not (a and b);
    layer6_outputs(3822) <= b;
    layer6_outputs(3823) <= '1';
    layer6_outputs(3824) <= not a;
    layer6_outputs(3825) <= a;
    layer6_outputs(3826) <= not b or a;
    layer6_outputs(3827) <= '0';
    layer6_outputs(3828) <= not b;
    layer6_outputs(3829) <= a or b;
    layer6_outputs(3830) <= a and b;
    layer6_outputs(3831) <= '0';
    layer6_outputs(3832) <= not a or b;
    layer6_outputs(3833) <= a and not b;
    layer6_outputs(3834) <= a and not b;
    layer6_outputs(3835) <= '1';
    layer6_outputs(3836) <= '1';
    layer6_outputs(3837) <= a and b;
    layer6_outputs(3838) <= not (a xor b);
    layer6_outputs(3839) <= not a;
    layer6_outputs(3840) <= a;
    layer6_outputs(3841) <= not a;
    layer6_outputs(3842) <= not (a and b);
    layer6_outputs(3843) <= not a or b;
    layer6_outputs(3844) <= not a;
    layer6_outputs(3845) <= a and b;
    layer6_outputs(3846) <= not b;
    layer6_outputs(3847) <= not a;
    layer6_outputs(3848) <= not b;
    layer6_outputs(3849) <= a or b;
    layer6_outputs(3850) <= a xor b;
    layer6_outputs(3851) <= a and b;
    layer6_outputs(3852) <= not (a and b);
    layer6_outputs(3853) <= not b or a;
    layer6_outputs(3854) <= a;
    layer6_outputs(3855) <= not a;
    layer6_outputs(3856) <= not (a and b);
    layer6_outputs(3857) <= a and b;
    layer6_outputs(3858) <= a and not b;
    layer6_outputs(3859) <= a;
    layer6_outputs(3860) <= a;
    layer6_outputs(3861) <= not b or a;
    layer6_outputs(3862) <= not (a or b);
    layer6_outputs(3863) <= not a;
    layer6_outputs(3864) <= not (a or b);
    layer6_outputs(3865) <= not (a and b);
    layer6_outputs(3866) <= not b;
    layer6_outputs(3867) <= not a or b;
    layer6_outputs(3868) <= not b;
    layer6_outputs(3869) <= a;
    layer6_outputs(3870) <= a;
    layer6_outputs(3871) <= not a;
    layer6_outputs(3872) <= not (a and b);
    layer6_outputs(3873) <= not (a and b);
    layer6_outputs(3874) <= not a;
    layer6_outputs(3875) <= not b;
    layer6_outputs(3876) <= a and not b;
    layer6_outputs(3877) <= not (a and b);
    layer6_outputs(3878) <= not (a and b);
    layer6_outputs(3879) <= a xor b;
    layer6_outputs(3880) <= a and b;
    layer6_outputs(3881) <= not (a or b);
    layer6_outputs(3882) <= a and b;
    layer6_outputs(3883) <= not a;
    layer6_outputs(3884) <= a;
    layer6_outputs(3885) <= not (a and b);
    layer6_outputs(3886) <= b and not a;
    layer6_outputs(3887) <= b;
    layer6_outputs(3888) <= not (a xor b);
    layer6_outputs(3889) <= '0';
    layer6_outputs(3890) <= not b;
    layer6_outputs(3891) <= a;
    layer6_outputs(3892) <= a;
    layer6_outputs(3893) <= not b;
    layer6_outputs(3894) <= a or b;
    layer6_outputs(3895) <= not a;
    layer6_outputs(3896) <= a or b;
    layer6_outputs(3897) <= a xor b;
    layer6_outputs(3898) <= a;
    layer6_outputs(3899) <= not (a or b);
    layer6_outputs(3900) <= not (a xor b);
    layer6_outputs(3901) <= not a or b;
    layer6_outputs(3902) <= not b;
    layer6_outputs(3903) <= b;
    layer6_outputs(3904) <= not (a xor b);
    layer6_outputs(3905) <= not (a xor b);
    layer6_outputs(3906) <= not a or b;
    layer6_outputs(3907) <= not a;
    layer6_outputs(3908) <= not (a and b);
    layer6_outputs(3909) <= not b;
    layer6_outputs(3910) <= b;
    layer6_outputs(3911) <= not (a or b);
    layer6_outputs(3912) <= not b;
    layer6_outputs(3913) <= not a;
    layer6_outputs(3914) <= not a;
    layer6_outputs(3915) <= not b;
    layer6_outputs(3916) <= a;
    layer6_outputs(3917) <= a or b;
    layer6_outputs(3918) <= not a or b;
    layer6_outputs(3919) <= not b;
    layer6_outputs(3920) <= not (a or b);
    layer6_outputs(3921) <= not b or a;
    layer6_outputs(3922) <= not a;
    layer6_outputs(3923) <= b;
    layer6_outputs(3924) <= b and not a;
    layer6_outputs(3925) <= a and not b;
    layer6_outputs(3926) <= b;
    layer6_outputs(3927) <= a;
    layer6_outputs(3928) <= not a;
    layer6_outputs(3929) <= not b;
    layer6_outputs(3930) <= a and not b;
    layer6_outputs(3931) <= not a;
    layer6_outputs(3932) <= a and not b;
    layer6_outputs(3933) <= not a;
    layer6_outputs(3934) <= not a;
    layer6_outputs(3935) <= a or b;
    layer6_outputs(3936) <= a and b;
    layer6_outputs(3937) <= a or b;
    layer6_outputs(3938) <= '1';
    layer6_outputs(3939) <= b;
    layer6_outputs(3940) <= not (a or b);
    layer6_outputs(3941) <= not b;
    layer6_outputs(3942) <= not a;
    layer6_outputs(3943) <= not (a or b);
    layer6_outputs(3944) <= not (a and b);
    layer6_outputs(3945) <= not (a or b);
    layer6_outputs(3946) <= not a or b;
    layer6_outputs(3947) <= not b or a;
    layer6_outputs(3948) <= not a;
    layer6_outputs(3949) <= a and b;
    layer6_outputs(3950) <= a;
    layer6_outputs(3951) <= not a or b;
    layer6_outputs(3952) <= not a or b;
    layer6_outputs(3953) <= a and b;
    layer6_outputs(3954) <= not b or a;
    layer6_outputs(3955) <= not b;
    layer6_outputs(3956) <= not (a and b);
    layer6_outputs(3957) <= not a;
    layer6_outputs(3958) <= not a;
    layer6_outputs(3959) <= not (a and b);
    layer6_outputs(3960) <= not a;
    layer6_outputs(3961) <= not b;
    layer6_outputs(3962) <= a;
    layer6_outputs(3963) <= b;
    layer6_outputs(3964) <= not a or b;
    layer6_outputs(3965) <= not b;
    layer6_outputs(3966) <= not (a xor b);
    layer6_outputs(3967) <= a xor b;
    layer6_outputs(3968) <= not a;
    layer6_outputs(3969) <= not (a and b);
    layer6_outputs(3970) <= not (a xor b);
    layer6_outputs(3971) <= not (a xor b);
    layer6_outputs(3972) <= not b or a;
    layer6_outputs(3973) <= not a;
    layer6_outputs(3974) <= a or b;
    layer6_outputs(3975) <= a;
    layer6_outputs(3976) <= not b or a;
    layer6_outputs(3977) <= not b;
    layer6_outputs(3978) <= a;
    layer6_outputs(3979) <= not b;
    layer6_outputs(3980) <= not b;
    layer6_outputs(3981) <= a;
    layer6_outputs(3982) <= not b;
    layer6_outputs(3983) <= not a;
    layer6_outputs(3984) <= b;
    layer6_outputs(3985) <= b and not a;
    layer6_outputs(3986) <= not a;
    layer6_outputs(3987) <= a;
    layer6_outputs(3988) <= not a;
    layer6_outputs(3989) <= a or b;
    layer6_outputs(3990) <= not b;
    layer6_outputs(3991) <= not a;
    layer6_outputs(3992) <= b and not a;
    layer6_outputs(3993) <= a and not b;
    layer6_outputs(3994) <= a or b;
    layer6_outputs(3995) <= b;
    layer6_outputs(3996) <= not (a xor b);
    layer6_outputs(3997) <= a and b;
    layer6_outputs(3998) <= a and b;
    layer6_outputs(3999) <= '1';
    layer6_outputs(4000) <= a;
    layer6_outputs(4001) <= b and not a;
    layer6_outputs(4002) <= a;
    layer6_outputs(4003) <= a xor b;
    layer6_outputs(4004) <= a xor b;
    layer6_outputs(4005) <= b and not a;
    layer6_outputs(4006) <= not (a and b);
    layer6_outputs(4007) <= not a;
    layer6_outputs(4008) <= a;
    layer6_outputs(4009) <= '0';
    layer6_outputs(4010) <= a and b;
    layer6_outputs(4011) <= a or b;
    layer6_outputs(4012) <= b;
    layer6_outputs(4013) <= not b or a;
    layer6_outputs(4014) <= b;
    layer6_outputs(4015) <= not b;
    layer6_outputs(4016) <= not (a and b);
    layer6_outputs(4017) <= a;
    layer6_outputs(4018) <= a or b;
    layer6_outputs(4019) <= not b or a;
    layer6_outputs(4020) <= not (a or b);
    layer6_outputs(4021) <= not (a or b);
    layer6_outputs(4022) <= a and b;
    layer6_outputs(4023) <= b and not a;
    layer6_outputs(4024) <= b and not a;
    layer6_outputs(4025) <= b and not a;
    layer6_outputs(4026) <= not (a and b);
    layer6_outputs(4027) <= b;
    layer6_outputs(4028) <= b and not a;
    layer6_outputs(4029) <= b;
    layer6_outputs(4030) <= b and not a;
    layer6_outputs(4031) <= a;
    layer6_outputs(4032) <= a or b;
    layer6_outputs(4033) <= not (a or b);
    layer6_outputs(4034) <= not a;
    layer6_outputs(4035) <= a and b;
    layer6_outputs(4036) <= b;
    layer6_outputs(4037) <= a or b;
    layer6_outputs(4038) <= a or b;
    layer6_outputs(4039) <= b;
    layer6_outputs(4040) <= not b;
    layer6_outputs(4041) <= a;
    layer6_outputs(4042) <= not a;
    layer6_outputs(4043) <= a or b;
    layer6_outputs(4044) <= not (a and b);
    layer6_outputs(4045) <= a and not b;
    layer6_outputs(4046) <= not a or b;
    layer6_outputs(4047) <= not (a xor b);
    layer6_outputs(4048) <= b;
    layer6_outputs(4049) <= b;
    layer6_outputs(4050) <= b;
    layer6_outputs(4051) <= b and not a;
    layer6_outputs(4052) <= not a or b;
    layer6_outputs(4053) <= a and b;
    layer6_outputs(4054) <= not b;
    layer6_outputs(4055) <= not b;
    layer6_outputs(4056) <= not a;
    layer6_outputs(4057) <= a;
    layer6_outputs(4058) <= not (a xor b);
    layer6_outputs(4059) <= not (a or b);
    layer6_outputs(4060) <= a or b;
    layer6_outputs(4061) <= not (a and b);
    layer6_outputs(4062) <= a;
    layer6_outputs(4063) <= not (a and b);
    layer6_outputs(4064) <= not (a and b);
    layer6_outputs(4065) <= a xor b;
    layer6_outputs(4066) <= not a;
    layer6_outputs(4067) <= a and b;
    layer6_outputs(4068) <= not a or b;
    layer6_outputs(4069) <= a xor b;
    layer6_outputs(4070) <= b;
    layer6_outputs(4071) <= a and b;
    layer6_outputs(4072) <= a;
    layer6_outputs(4073) <= a xor b;
    layer6_outputs(4074) <= not (a xor b);
    layer6_outputs(4075) <= a xor b;
    layer6_outputs(4076) <= a and not b;
    layer6_outputs(4077) <= '1';
    layer6_outputs(4078) <= b;
    layer6_outputs(4079) <= a or b;
    layer6_outputs(4080) <= b and not a;
    layer6_outputs(4081) <= a;
    layer6_outputs(4082) <= b;
    layer6_outputs(4083) <= not b or a;
    layer6_outputs(4084) <= a;
    layer6_outputs(4085) <= a;
    layer6_outputs(4086) <= b and not a;
    layer6_outputs(4087) <= a xor b;
    layer6_outputs(4088) <= not a;
    layer6_outputs(4089) <= b and not a;
    layer6_outputs(4090) <= b and not a;
    layer6_outputs(4091) <= not b or a;
    layer6_outputs(4092) <= a;
    layer6_outputs(4093) <= not a;
    layer6_outputs(4094) <= a and b;
    layer6_outputs(4095) <= not a or b;
    layer6_outputs(4096) <= not b;
    layer6_outputs(4097) <= b;
    layer6_outputs(4098) <= not b or a;
    layer6_outputs(4099) <= '1';
    layer6_outputs(4100) <= '1';
    layer6_outputs(4101) <= not a;
    layer6_outputs(4102) <= a;
    layer6_outputs(4103) <= b;
    layer6_outputs(4104) <= not (a and b);
    layer6_outputs(4105) <= not (a xor b);
    layer6_outputs(4106) <= not b or a;
    layer6_outputs(4107) <= not b or a;
    layer6_outputs(4108) <= b and not a;
    layer6_outputs(4109) <= not (a xor b);
    layer6_outputs(4110) <= a;
    layer6_outputs(4111) <= not (a xor b);
    layer6_outputs(4112) <= not a;
    layer6_outputs(4113) <= not (a and b);
    layer6_outputs(4114) <= not (a xor b);
    layer6_outputs(4115) <= not b or a;
    layer6_outputs(4116) <= not a;
    layer6_outputs(4117) <= a;
    layer6_outputs(4118) <= not a;
    layer6_outputs(4119) <= not b or a;
    layer6_outputs(4120) <= a;
    layer6_outputs(4121) <= not a;
    layer6_outputs(4122) <= not (a and b);
    layer6_outputs(4123) <= a;
    layer6_outputs(4124) <= a xor b;
    layer6_outputs(4125) <= '1';
    layer6_outputs(4126) <= not (a xor b);
    layer6_outputs(4127) <= a and b;
    layer6_outputs(4128) <= not (a and b);
    layer6_outputs(4129) <= b;
    layer6_outputs(4130) <= not a;
    layer6_outputs(4131) <= not b or a;
    layer6_outputs(4132) <= a;
    layer6_outputs(4133) <= not (a or b);
    layer6_outputs(4134) <= a and not b;
    layer6_outputs(4135) <= not (a and b);
    layer6_outputs(4136) <= a or b;
    layer6_outputs(4137) <= not (a and b);
    layer6_outputs(4138) <= a and b;
    layer6_outputs(4139) <= not (a and b);
    layer6_outputs(4140) <= a or b;
    layer6_outputs(4141) <= a;
    layer6_outputs(4142) <= not (a and b);
    layer6_outputs(4143) <= a and b;
    layer6_outputs(4144) <= a xor b;
    layer6_outputs(4145) <= not b or a;
    layer6_outputs(4146) <= not a or b;
    layer6_outputs(4147) <= b and not a;
    layer6_outputs(4148) <= a;
    layer6_outputs(4149) <= a;
    layer6_outputs(4150) <= not b;
    layer6_outputs(4151) <= not b or a;
    layer6_outputs(4152) <= a or b;
    layer6_outputs(4153) <= '1';
    layer6_outputs(4154) <= a and b;
    layer6_outputs(4155) <= a;
    layer6_outputs(4156) <= not a;
    layer6_outputs(4157) <= b;
    layer6_outputs(4158) <= a or b;
    layer6_outputs(4159) <= a and b;
    layer6_outputs(4160) <= a and not b;
    layer6_outputs(4161) <= not a;
    layer6_outputs(4162) <= not a;
    layer6_outputs(4163) <= a and b;
    layer6_outputs(4164) <= a;
    layer6_outputs(4165) <= not (a xor b);
    layer6_outputs(4166) <= a xor b;
    layer6_outputs(4167) <= not b;
    layer6_outputs(4168) <= not (a and b);
    layer6_outputs(4169) <= b and not a;
    layer6_outputs(4170) <= b;
    layer6_outputs(4171) <= not (a or b);
    layer6_outputs(4172) <= not (a or b);
    layer6_outputs(4173) <= not b or a;
    layer6_outputs(4174) <= not a or b;
    layer6_outputs(4175) <= not a;
    layer6_outputs(4176) <= '1';
    layer6_outputs(4177) <= a and b;
    layer6_outputs(4178) <= not (a xor b);
    layer6_outputs(4179) <= b and not a;
    layer6_outputs(4180) <= not a;
    layer6_outputs(4181) <= not b or a;
    layer6_outputs(4182) <= not a;
    layer6_outputs(4183) <= not a;
    layer6_outputs(4184) <= b and not a;
    layer6_outputs(4185) <= a and not b;
    layer6_outputs(4186) <= a;
    layer6_outputs(4187) <= a xor b;
    layer6_outputs(4188) <= not a;
    layer6_outputs(4189) <= not (a or b);
    layer6_outputs(4190) <= not (a or b);
    layer6_outputs(4191) <= not b;
    layer6_outputs(4192) <= not a;
    layer6_outputs(4193) <= '1';
    layer6_outputs(4194) <= a xor b;
    layer6_outputs(4195) <= not b or a;
    layer6_outputs(4196) <= not (a or b);
    layer6_outputs(4197) <= not a;
    layer6_outputs(4198) <= not a;
    layer6_outputs(4199) <= a xor b;
    layer6_outputs(4200) <= b;
    layer6_outputs(4201) <= a or b;
    layer6_outputs(4202) <= b;
    layer6_outputs(4203) <= a or b;
    layer6_outputs(4204) <= not (a xor b);
    layer6_outputs(4205) <= a and b;
    layer6_outputs(4206) <= not b;
    layer6_outputs(4207) <= not a;
    layer6_outputs(4208) <= not a;
    layer6_outputs(4209) <= '0';
    layer6_outputs(4210) <= not (a or b);
    layer6_outputs(4211) <= not b or a;
    layer6_outputs(4212) <= a;
    layer6_outputs(4213) <= b;
    layer6_outputs(4214) <= not (a or b);
    layer6_outputs(4215) <= not b or a;
    layer6_outputs(4216) <= not b;
    layer6_outputs(4217) <= not a or b;
    layer6_outputs(4218) <= not a;
    layer6_outputs(4219) <= a and b;
    layer6_outputs(4220) <= a and b;
    layer6_outputs(4221) <= '0';
    layer6_outputs(4222) <= not b;
    layer6_outputs(4223) <= not a or b;
    layer6_outputs(4224) <= not (a or b);
    layer6_outputs(4225) <= not a;
    layer6_outputs(4226) <= b and not a;
    layer6_outputs(4227) <= not b;
    layer6_outputs(4228) <= a and not b;
    layer6_outputs(4229) <= a;
    layer6_outputs(4230) <= not (a xor b);
    layer6_outputs(4231) <= b and not a;
    layer6_outputs(4232) <= b and not a;
    layer6_outputs(4233) <= not b;
    layer6_outputs(4234) <= not (a or b);
    layer6_outputs(4235) <= a;
    layer6_outputs(4236) <= '0';
    layer6_outputs(4237) <= a and not b;
    layer6_outputs(4238) <= b;
    layer6_outputs(4239) <= a and b;
    layer6_outputs(4240) <= not b;
    layer6_outputs(4241) <= not (a xor b);
    layer6_outputs(4242) <= a;
    layer6_outputs(4243) <= b;
    layer6_outputs(4244) <= a;
    layer6_outputs(4245) <= not a;
    layer6_outputs(4246) <= a and not b;
    layer6_outputs(4247) <= not b;
    layer6_outputs(4248) <= not b or a;
    layer6_outputs(4249) <= not a;
    layer6_outputs(4250) <= b;
    layer6_outputs(4251) <= a or b;
    layer6_outputs(4252) <= not b or a;
    layer6_outputs(4253) <= a and not b;
    layer6_outputs(4254) <= a;
    layer6_outputs(4255) <= b;
    layer6_outputs(4256) <= not a;
    layer6_outputs(4257) <= not b;
    layer6_outputs(4258) <= a xor b;
    layer6_outputs(4259) <= not b;
    layer6_outputs(4260) <= not b or a;
    layer6_outputs(4261) <= not a or b;
    layer6_outputs(4262) <= a xor b;
    layer6_outputs(4263) <= a;
    layer6_outputs(4264) <= b;
    layer6_outputs(4265) <= not (a xor b);
    layer6_outputs(4266) <= not b or a;
    layer6_outputs(4267) <= a xor b;
    layer6_outputs(4268) <= a;
    layer6_outputs(4269) <= not (a xor b);
    layer6_outputs(4270) <= a;
    layer6_outputs(4271) <= not (a or b);
    layer6_outputs(4272) <= a or b;
    layer6_outputs(4273) <= not b or a;
    layer6_outputs(4274) <= b;
    layer6_outputs(4275) <= not b;
    layer6_outputs(4276) <= a and not b;
    layer6_outputs(4277) <= a;
    layer6_outputs(4278) <= a or b;
    layer6_outputs(4279) <= b;
    layer6_outputs(4280) <= a or b;
    layer6_outputs(4281) <= a and b;
    layer6_outputs(4282) <= b;
    layer6_outputs(4283) <= not a;
    layer6_outputs(4284) <= not (a or b);
    layer6_outputs(4285) <= a or b;
    layer6_outputs(4286) <= a or b;
    layer6_outputs(4287) <= not b;
    layer6_outputs(4288) <= b;
    layer6_outputs(4289) <= not a;
    layer6_outputs(4290) <= not a or b;
    layer6_outputs(4291) <= not a;
    layer6_outputs(4292) <= b;
    layer6_outputs(4293) <= not b;
    layer6_outputs(4294) <= not b or a;
    layer6_outputs(4295) <= a or b;
    layer6_outputs(4296) <= a or b;
    layer6_outputs(4297) <= a and not b;
    layer6_outputs(4298) <= b;
    layer6_outputs(4299) <= a and not b;
    layer6_outputs(4300) <= not a;
    layer6_outputs(4301) <= '0';
    layer6_outputs(4302) <= a;
    layer6_outputs(4303) <= a;
    layer6_outputs(4304) <= not b;
    layer6_outputs(4305) <= a and not b;
    layer6_outputs(4306) <= a and b;
    layer6_outputs(4307) <= b;
    layer6_outputs(4308) <= not a;
    layer6_outputs(4309) <= b and not a;
    layer6_outputs(4310) <= not b or a;
    layer6_outputs(4311) <= not a or b;
    layer6_outputs(4312) <= b;
    layer6_outputs(4313) <= not a;
    layer6_outputs(4314) <= a or b;
    layer6_outputs(4315) <= b and not a;
    layer6_outputs(4316) <= a or b;
    layer6_outputs(4317) <= not a;
    layer6_outputs(4318) <= b and not a;
    layer6_outputs(4319) <= '0';
    layer6_outputs(4320) <= a or b;
    layer6_outputs(4321) <= a;
    layer6_outputs(4322) <= not (a and b);
    layer6_outputs(4323) <= a and not b;
    layer6_outputs(4324) <= a and not b;
    layer6_outputs(4325) <= a xor b;
    layer6_outputs(4326) <= not b or a;
    layer6_outputs(4327) <= not (a or b);
    layer6_outputs(4328) <= b and not a;
    layer6_outputs(4329) <= not (a or b);
    layer6_outputs(4330) <= not a;
    layer6_outputs(4331) <= a;
    layer6_outputs(4332) <= a and not b;
    layer6_outputs(4333) <= not (a xor b);
    layer6_outputs(4334) <= b;
    layer6_outputs(4335) <= a xor b;
    layer6_outputs(4336) <= not a;
    layer6_outputs(4337) <= not b;
    layer6_outputs(4338) <= not a or b;
    layer6_outputs(4339) <= not b or a;
    layer6_outputs(4340) <= not a or b;
    layer6_outputs(4341) <= b and not a;
    layer6_outputs(4342) <= not b;
    layer6_outputs(4343) <= b;
    layer6_outputs(4344) <= not a;
    layer6_outputs(4345) <= not a;
    layer6_outputs(4346) <= b;
    layer6_outputs(4347) <= not b or a;
    layer6_outputs(4348) <= a and not b;
    layer6_outputs(4349) <= '1';
    layer6_outputs(4350) <= not b;
    layer6_outputs(4351) <= not a or b;
    layer6_outputs(4352) <= not a or b;
    layer6_outputs(4353) <= b;
    layer6_outputs(4354) <= not (a xor b);
    layer6_outputs(4355) <= a and not b;
    layer6_outputs(4356) <= b;
    layer6_outputs(4357) <= a or b;
    layer6_outputs(4358) <= not b;
    layer6_outputs(4359) <= not a;
    layer6_outputs(4360) <= not (a or b);
    layer6_outputs(4361) <= not a;
    layer6_outputs(4362) <= a;
    layer6_outputs(4363) <= a or b;
    layer6_outputs(4364) <= a and not b;
    layer6_outputs(4365) <= not b or a;
    layer6_outputs(4366) <= not a or b;
    layer6_outputs(4367) <= not b;
    layer6_outputs(4368) <= b;
    layer6_outputs(4369) <= b;
    layer6_outputs(4370) <= a;
    layer6_outputs(4371) <= b;
    layer6_outputs(4372) <= not (a or b);
    layer6_outputs(4373) <= not (a or b);
    layer6_outputs(4374) <= a and not b;
    layer6_outputs(4375) <= not a or b;
    layer6_outputs(4376) <= a;
    layer6_outputs(4377) <= b;
    layer6_outputs(4378) <= b;
    layer6_outputs(4379) <= a;
    layer6_outputs(4380) <= not b;
    layer6_outputs(4381) <= a;
    layer6_outputs(4382) <= a and not b;
    layer6_outputs(4383) <= b;
    layer6_outputs(4384) <= a;
    layer6_outputs(4385) <= b;
    layer6_outputs(4386) <= a;
    layer6_outputs(4387) <= a;
    layer6_outputs(4388) <= not b;
    layer6_outputs(4389) <= not a or b;
    layer6_outputs(4390) <= not a;
    layer6_outputs(4391) <= b and not a;
    layer6_outputs(4392) <= a;
    layer6_outputs(4393) <= b;
    layer6_outputs(4394) <= not b;
    layer6_outputs(4395) <= not (a or b);
    layer6_outputs(4396) <= a;
    layer6_outputs(4397) <= not b;
    layer6_outputs(4398) <= a or b;
    layer6_outputs(4399) <= a;
    layer6_outputs(4400) <= not a;
    layer6_outputs(4401) <= a and b;
    layer6_outputs(4402) <= b;
    layer6_outputs(4403) <= not (a and b);
    layer6_outputs(4404) <= a;
    layer6_outputs(4405) <= b;
    layer6_outputs(4406) <= not (a and b);
    layer6_outputs(4407) <= not (a or b);
    layer6_outputs(4408) <= a xor b;
    layer6_outputs(4409) <= a;
    layer6_outputs(4410) <= not (a or b);
    layer6_outputs(4411) <= a and not b;
    layer6_outputs(4412) <= b;
    layer6_outputs(4413) <= a;
    layer6_outputs(4414) <= a or b;
    layer6_outputs(4415) <= a and b;
    layer6_outputs(4416) <= a xor b;
    layer6_outputs(4417) <= not (a xor b);
    layer6_outputs(4418) <= not (a xor b);
    layer6_outputs(4419) <= not a;
    layer6_outputs(4420) <= not b;
    layer6_outputs(4421) <= not (a xor b);
    layer6_outputs(4422) <= b;
    layer6_outputs(4423) <= a;
    layer6_outputs(4424) <= not b;
    layer6_outputs(4425) <= not (a or b);
    layer6_outputs(4426) <= not (a xor b);
    layer6_outputs(4427) <= not b or a;
    layer6_outputs(4428) <= not (a or b);
    layer6_outputs(4429) <= a;
    layer6_outputs(4430) <= not b or a;
    layer6_outputs(4431) <= '0';
    layer6_outputs(4432) <= not b;
    layer6_outputs(4433) <= a;
    layer6_outputs(4434) <= not a;
    layer6_outputs(4435) <= a;
    layer6_outputs(4436) <= not a;
    layer6_outputs(4437) <= a or b;
    layer6_outputs(4438) <= not (a and b);
    layer6_outputs(4439) <= not a;
    layer6_outputs(4440) <= a or b;
    layer6_outputs(4441) <= a xor b;
    layer6_outputs(4442) <= not b;
    layer6_outputs(4443) <= a and b;
    layer6_outputs(4444) <= not (a or b);
    layer6_outputs(4445) <= a;
    layer6_outputs(4446) <= not b;
    layer6_outputs(4447) <= a xor b;
    layer6_outputs(4448) <= a and b;
    layer6_outputs(4449) <= not (a and b);
    layer6_outputs(4450) <= not (a and b);
    layer6_outputs(4451) <= a and not b;
    layer6_outputs(4452) <= a xor b;
    layer6_outputs(4453) <= a xor b;
    layer6_outputs(4454) <= not (a and b);
    layer6_outputs(4455) <= a and b;
    layer6_outputs(4456) <= b;
    layer6_outputs(4457) <= not b or a;
    layer6_outputs(4458) <= not (a xor b);
    layer6_outputs(4459) <= not (a xor b);
    layer6_outputs(4460) <= a and not b;
    layer6_outputs(4461) <= b;
    layer6_outputs(4462) <= not b or a;
    layer6_outputs(4463) <= not a or b;
    layer6_outputs(4464) <= not (a and b);
    layer6_outputs(4465) <= a xor b;
    layer6_outputs(4466) <= b;
    layer6_outputs(4467) <= b and not a;
    layer6_outputs(4468) <= not b;
    layer6_outputs(4469) <= b;
    layer6_outputs(4470) <= a and b;
    layer6_outputs(4471) <= not (a or b);
    layer6_outputs(4472) <= not (a and b);
    layer6_outputs(4473) <= not b or a;
    layer6_outputs(4474) <= not a;
    layer6_outputs(4475) <= not a or b;
    layer6_outputs(4476) <= not (a xor b);
    layer6_outputs(4477) <= a xor b;
    layer6_outputs(4478) <= not a;
    layer6_outputs(4479) <= a xor b;
    layer6_outputs(4480) <= not a;
    layer6_outputs(4481) <= not b or a;
    layer6_outputs(4482) <= not a or b;
    layer6_outputs(4483) <= a and not b;
    layer6_outputs(4484) <= a or b;
    layer6_outputs(4485) <= not a;
    layer6_outputs(4486) <= b;
    layer6_outputs(4487) <= not b or a;
    layer6_outputs(4488) <= a;
    layer6_outputs(4489) <= a xor b;
    layer6_outputs(4490) <= not b;
    layer6_outputs(4491) <= not a or b;
    layer6_outputs(4492) <= b;
    layer6_outputs(4493) <= a and not b;
    layer6_outputs(4494) <= a;
    layer6_outputs(4495) <= a;
    layer6_outputs(4496) <= a xor b;
    layer6_outputs(4497) <= a;
    layer6_outputs(4498) <= not b;
    layer6_outputs(4499) <= a or b;
    layer6_outputs(4500) <= not b;
    layer6_outputs(4501) <= b;
    layer6_outputs(4502) <= a xor b;
    layer6_outputs(4503) <= not b or a;
    layer6_outputs(4504) <= a;
    layer6_outputs(4505) <= not (a or b);
    layer6_outputs(4506) <= a and not b;
    layer6_outputs(4507) <= not b;
    layer6_outputs(4508) <= not (a and b);
    layer6_outputs(4509) <= not b;
    layer6_outputs(4510) <= b;
    layer6_outputs(4511) <= a and b;
    layer6_outputs(4512) <= a and not b;
    layer6_outputs(4513) <= not a or b;
    layer6_outputs(4514) <= not (a and b);
    layer6_outputs(4515) <= not b;
    layer6_outputs(4516) <= a;
    layer6_outputs(4517) <= not a;
    layer6_outputs(4518) <= not a;
    layer6_outputs(4519) <= b and not a;
    layer6_outputs(4520) <= not (a and b);
    layer6_outputs(4521) <= a and not b;
    layer6_outputs(4522) <= not a or b;
    layer6_outputs(4523) <= b;
    layer6_outputs(4524) <= not b;
    layer6_outputs(4525) <= not b or a;
    layer6_outputs(4526) <= a or b;
    layer6_outputs(4527) <= a and not b;
    layer6_outputs(4528) <= b and not a;
    layer6_outputs(4529) <= a;
    layer6_outputs(4530) <= not (a and b);
    layer6_outputs(4531) <= not a or b;
    layer6_outputs(4532) <= not b;
    layer6_outputs(4533) <= a or b;
    layer6_outputs(4534) <= not a or b;
    layer6_outputs(4535) <= not (a xor b);
    layer6_outputs(4536) <= not a or b;
    layer6_outputs(4537) <= not a;
    layer6_outputs(4538) <= a;
    layer6_outputs(4539) <= b;
    layer6_outputs(4540) <= not a;
    layer6_outputs(4541) <= not a;
    layer6_outputs(4542) <= a or b;
    layer6_outputs(4543) <= not (a or b);
    layer6_outputs(4544) <= not a;
    layer6_outputs(4545) <= not a or b;
    layer6_outputs(4546) <= not b;
    layer6_outputs(4547) <= a and not b;
    layer6_outputs(4548) <= not a;
    layer6_outputs(4549) <= a xor b;
    layer6_outputs(4550) <= not b;
    layer6_outputs(4551) <= not b or a;
    layer6_outputs(4552) <= b;
    layer6_outputs(4553) <= a or b;
    layer6_outputs(4554) <= not b or a;
    layer6_outputs(4555) <= a;
    layer6_outputs(4556) <= not a;
    layer6_outputs(4557) <= '0';
    layer6_outputs(4558) <= a;
    layer6_outputs(4559) <= not (a and b);
    layer6_outputs(4560) <= a or b;
    layer6_outputs(4561) <= a xor b;
    layer6_outputs(4562) <= not (a xor b);
    layer6_outputs(4563) <= not a or b;
    layer6_outputs(4564) <= b;
    layer6_outputs(4565) <= '1';
    layer6_outputs(4566) <= not a or b;
    layer6_outputs(4567) <= a;
    layer6_outputs(4568) <= not a;
    layer6_outputs(4569) <= not a;
    layer6_outputs(4570) <= not a;
    layer6_outputs(4571) <= not b;
    layer6_outputs(4572) <= b;
    layer6_outputs(4573) <= b;
    layer6_outputs(4574) <= not a;
    layer6_outputs(4575) <= a;
    layer6_outputs(4576) <= b;
    layer6_outputs(4577) <= not (a xor b);
    layer6_outputs(4578) <= not a;
    layer6_outputs(4579) <= a and b;
    layer6_outputs(4580) <= a;
    layer6_outputs(4581) <= a xor b;
    layer6_outputs(4582) <= not (a or b);
    layer6_outputs(4583) <= not (a or b);
    layer6_outputs(4584) <= not b;
    layer6_outputs(4585) <= not (a or b);
    layer6_outputs(4586) <= a and b;
    layer6_outputs(4587) <= not a;
    layer6_outputs(4588) <= not b;
    layer6_outputs(4589) <= b;
    layer6_outputs(4590) <= not (a or b);
    layer6_outputs(4591) <= a and b;
    layer6_outputs(4592) <= b and not a;
    layer6_outputs(4593) <= b;
    layer6_outputs(4594) <= a and not b;
    layer6_outputs(4595) <= b and not a;
    layer6_outputs(4596) <= not a;
    layer6_outputs(4597) <= not b;
    layer6_outputs(4598) <= not a or b;
    layer6_outputs(4599) <= a and not b;
    layer6_outputs(4600) <= b;
    layer6_outputs(4601) <= b;
    layer6_outputs(4602) <= a and not b;
    layer6_outputs(4603) <= not (a xor b);
    layer6_outputs(4604) <= b;
    layer6_outputs(4605) <= b and not a;
    layer6_outputs(4606) <= a or b;
    layer6_outputs(4607) <= not a or b;
    layer6_outputs(4608) <= not a or b;
    layer6_outputs(4609) <= a and not b;
    layer6_outputs(4610) <= a and not b;
    layer6_outputs(4611) <= not b;
    layer6_outputs(4612) <= b and not a;
    layer6_outputs(4613) <= not a or b;
    layer6_outputs(4614) <= b and not a;
    layer6_outputs(4615) <= b;
    layer6_outputs(4616) <= not (a or b);
    layer6_outputs(4617) <= a xor b;
    layer6_outputs(4618) <= not a or b;
    layer6_outputs(4619) <= a xor b;
    layer6_outputs(4620) <= a and b;
    layer6_outputs(4621) <= b;
    layer6_outputs(4622) <= a xor b;
    layer6_outputs(4623) <= not a;
    layer6_outputs(4624) <= '1';
    layer6_outputs(4625) <= not (a and b);
    layer6_outputs(4626) <= not b or a;
    layer6_outputs(4627) <= not (a or b);
    layer6_outputs(4628) <= a;
    layer6_outputs(4629) <= not a;
    layer6_outputs(4630) <= b;
    layer6_outputs(4631) <= not (a and b);
    layer6_outputs(4632) <= a and b;
    layer6_outputs(4633) <= not a or b;
    layer6_outputs(4634) <= b;
    layer6_outputs(4635) <= a;
    layer6_outputs(4636) <= a and not b;
    layer6_outputs(4637) <= a;
    layer6_outputs(4638) <= not b;
    layer6_outputs(4639) <= a or b;
    layer6_outputs(4640) <= not b;
    layer6_outputs(4641) <= a;
    layer6_outputs(4642) <= not (a and b);
    layer6_outputs(4643) <= not b or a;
    layer6_outputs(4644) <= b and not a;
    layer6_outputs(4645) <= a or b;
    layer6_outputs(4646) <= a and b;
    layer6_outputs(4647) <= not a;
    layer6_outputs(4648) <= not (a or b);
    layer6_outputs(4649) <= not b or a;
    layer6_outputs(4650) <= not (a xor b);
    layer6_outputs(4651) <= not (a xor b);
    layer6_outputs(4652) <= a xor b;
    layer6_outputs(4653) <= '1';
    layer6_outputs(4654) <= not (a xor b);
    layer6_outputs(4655) <= not (a xor b);
    layer6_outputs(4656) <= not b;
    layer6_outputs(4657) <= not (a xor b);
    layer6_outputs(4658) <= a and not b;
    layer6_outputs(4659) <= not b or a;
    layer6_outputs(4660) <= '0';
    layer6_outputs(4661) <= not (a or b);
    layer6_outputs(4662) <= b;
    layer6_outputs(4663) <= a xor b;
    layer6_outputs(4664) <= not b or a;
    layer6_outputs(4665) <= a or b;
    layer6_outputs(4666) <= not (a or b);
    layer6_outputs(4667) <= not a;
    layer6_outputs(4668) <= a;
    layer6_outputs(4669) <= not a;
    layer6_outputs(4670) <= not (a or b);
    layer6_outputs(4671) <= not a;
    layer6_outputs(4672) <= not (a xor b);
    layer6_outputs(4673) <= a and b;
    layer6_outputs(4674) <= a;
    layer6_outputs(4675) <= not a or b;
    layer6_outputs(4676) <= b and not a;
    layer6_outputs(4677) <= not (a and b);
    layer6_outputs(4678) <= not a;
    layer6_outputs(4679) <= b and not a;
    layer6_outputs(4680) <= not (a xor b);
    layer6_outputs(4681) <= not b;
    layer6_outputs(4682) <= a and not b;
    layer6_outputs(4683) <= not (a xor b);
    layer6_outputs(4684) <= a and b;
    layer6_outputs(4685) <= b;
    layer6_outputs(4686) <= b and not a;
    layer6_outputs(4687) <= a;
    layer6_outputs(4688) <= not b or a;
    layer6_outputs(4689) <= not b;
    layer6_outputs(4690) <= b;
    layer6_outputs(4691) <= not a;
    layer6_outputs(4692) <= a;
    layer6_outputs(4693) <= b;
    layer6_outputs(4694) <= not b or a;
    layer6_outputs(4695) <= a;
    layer6_outputs(4696) <= b and not a;
    layer6_outputs(4697) <= not a or b;
    layer6_outputs(4698) <= not b or a;
    layer6_outputs(4699) <= a and not b;
    layer6_outputs(4700) <= a and b;
    layer6_outputs(4701) <= a;
    layer6_outputs(4702) <= not b;
    layer6_outputs(4703) <= a xor b;
    layer6_outputs(4704) <= a;
    layer6_outputs(4705) <= a;
    layer6_outputs(4706) <= not (a and b);
    layer6_outputs(4707) <= a;
    layer6_outputs(4708) <= not b;
    layer6_outputs(4709) <= not b;
    layer6_outputs(4710) <= not (a xor b);
    layer6_outputs(4711) <= not (a or b);
    layer6_outputs(4712) <= '0';
    layer6_outputs(4713) <= b and not a;
    layer6_outputs(4714) <= not b or a;
    layer6_outputs(4715) <= not a;
    layer6_outputs(4716) <= not (a or b);
    layer6_outputs(4717) <= not b or a;
    layer6_outputs(4718) <= b;
    layer6_outputs(4719) <= '1';
    layer6_outputs(4720) <= a and not b;
    layer6_outputs(4721) <= not a;
    layer6_outputs(4722) <= not a;
    layer6_outputs(4723) <= not a;
    layer6_outputs(4724) <= a and not b;
    layer6_outputs(4725) <= not a;
    layer6_outputs(4726) <= not b or a;
    layer6_outputs(4727) <= '0';
    layer6_outputs(4728) <= a;
    layer6_outputs(4729) <= a and not b;
    layer6_outputs(4730) <= not (a and b);
    layer6_outputs(4731) <= not (a or b);
    layer6_outputs(4732) <= b;
    layer6_outputs(4733) <= not b;
    layer6_outputs(4734) <= b;
    layer6_outputs(4735) <= b;
    layer6_outputs(4736) <= a and not b;
    layer6_outputs(4737) <= not a or b;
    layer6_outputs(4738) <= a;
    layer6_outputs(4739) <= a;
    layer6_outputs(4740) <= a;
    layer6_outputs(4741) <= a xor b;
    layer6_outputs(4742) <= a;
    layer6_outputs(4743) <= b;
    layer6_outputs(4744) <= a and b;
    layer6_outputs(4745) <= not b or a;
    layer6_outputs(4746) <= b;
    layer6_outputs(4747) <= b;
    layer6_outputs(4748) <= a;
    layer6_outputs(4749) <= not b;
    layer6_outputs(4750) <= a or b;
    layer6_outputs(4751) <= not b or a;
    layer6_outputs(4752) <= not a or b;
    layer6_outputs(4753) <= not b;
    layer6_outputs(4754) <= not b;
    layer6_outputs(4755) <= '1';
    layer6_outputs(4756) <= a;
    layer6_outputs(4757) <= a;
    layer6_outputs(4758) <= not b;
    layer6_outputs(4759) <= b;
    layer6_outputs(4760) <= not (a xor b);
    layer6_outputs(4761) <= not b or a;
    layer6_outputs(4762) <= a xor b;
    layer6_outputs(4763) <= not (a xor b);
    layer6_outputs(4764) <= a or b;
    layer6_outputs(4765) <= a xor b;
    layer6_outputs(4766) <= not a;
    layer6_outputs(4767) <= not b;
    layer6_outputs(4768) <= a and not b;
    layer6_outputs(4769) <= not a or b;
    layer6_outputs(4770) <= not a or b;
    layer6_outputs(4771) <= a;
    layer6_outputs(4772) <= a and not b;
    layer6_outputs(4773) <= a xor b;
    layer6_outputs(4774) <= b;
    layer6_outputs(4775) <= '1';
    layer6_outputs(4776) <= not (a or b);
    layer6_outputs(4777) <= not a;
    layer6_outputs(4778) <= b and not a;
    layer6_outputs(4779) <= a;
    layer6_outputs(4780) <= a and not b;
    layer6_outputs(4781) <= b;
    layer6_outputs(4782) <= not (a or b);
    layer6_outputs(4783) <= b;
    layer6_outputs(4784) <= b and not a;
    layer6_outputs(4785) <= not (a xor b);
    layer6_outputs(4786) <= not a;
    layer6_outputs(4787) <= not (a and b);
    layer6_outputs(4788) <= not b;
    layer6_outputs(4789) <= a or b;
    layer6_outputs(4790) <= not a or b;
    layer6_outputs(4791) <= a and not b;
    layer6_outputs(4792) <= b and not a;
    layer6_outputs(4793) <= a and b;
    layer6_outputs(4794) <= a or b;
    layer6_outputs(4795) <= a and not b;
    layer6_outputs(4796) <= not (a or b);
    layer6_outputs(4797) <= not b;
    layer6_outputs(4798) <= a and not b;
    layer6_outputs(4799) <= not a;
    layer6_outputs(4800) <= b;
    layer6_outputs(4801) <= not a or b;
    layer6_outputs(4802) <= b;
    layer6_outputs(4803) <= not (a or b);
    layer6_outputs(4804) <= a xor b;
    layer6_outputs(4805) <= not b;
    layer6_outputs(4806) <= not (a xor b);
    layer6_outputs(4807) <= not a or b;
    layer6_outputs(4808) <= not b;
    layer6_outputs(4809) <= a xor b;
    layer6_outputs(4810) <= a and b;
    layer6_outputs(4811) <= a and b;
    layer6_outputs(4812) <= not b;
    layer6_outputs(4813) <= b;
    layer6_outputs(4814) <= not a;
    layer6_outputs(4815) <= not (a or b);
    layer6_outputs(4816) <= a;
    layer6_outputs(4817) <= not (a xor b);
    layer6_outputs(4818) <= not a;
    layer6_outputs(4819) <= a or b;
    layer6_outputs(4820) <= not b or a;
    layer6_outputs(4821) <= not (a and b);
    layer6_outputs(4822) <= not b;
    layer6_outputs(4823) <= a and not b;
    layer6_outputs(4824) <= not a;
    layer6_outputs(4825) <= b;
    layer6_outputs(4826) <= b and not a;
    layer6_outputs(4827) <= not a;
    layer6_outputs(4828) <= not (a or b);
    layer6_outputs(4829) <= b;
    layer6_outputs(4830) <= not a or b;
    layer6_outputs(4831) <= not a;
    layer6_outputs(4832) <= not b or a;
    layer6_outputs(4833) <= not a;
    layer6_outputs(4834) <= not b;
    layer6_outputs(4835) <= b and not a;
    layer6_outputs(4836) <= b and not a;
    layer6_outputs(4837) <= a;
    layer6_outputs(4838) <= not (a xor b);
    layer6_outputs(4839) <= a xor b;
    layer6_outputs(4840) <= a and b;
    layer6_outputs(4841) <= not (a xor b);
    layer6_outputs(4842) <= not a;
    layer6_outputs(4843) <= not a;
    layer6_outputs(4844) <= '0';
    layer6_outputs(4845) <= a;
    layer6_outputs(4846) <= not (a or b);
    layer6_outputs(4847) <= a or b;
    layer6_outputs(4848) <= a or b;
    layer6_outputs(4849) <= a and b;
    layer6_outputs(4850) <= not (a or b);
    layer6_outputs(4851) <= not (a or b);
    layer6_outputs(4852) <= b;
    layer6_outputs(4853) <= not (a xor b);
    layer6_outputs(4854) <= b;
    layer6_outputs(4855) <= b;
    layer6_outputs(4856) <= a;
    layer6_outputs(4857) <= '1';
    layer6_outputs(4858) <= a xor b;
    layer6_outputs(4859) <= not a;
    layer6_outputs(4860) <= not a or b;
    layer6_outputs(4861) <= not a;
    layer6_outputs(4862) <= a;
    layer6_outputs(4863) <= b and not a;
    layer6_outputs(4864) <= b;
    layer6_outputs(4865) <= b;
    layer6_outputs(4866) <= not (a xor b);
    layer6_outputs(4867) <= a and b;
    layer6_outputs(4868) <= not a;
    layer6_outputs(4869) <= not (a xor b);
    layer6_outputs(4870) <= b and not a;
    layer6_outputs(4871) <= not (a xor b);
    layer6_outputs(4872) <= b and not a;
    layer6_outputs(4873) <= b and not a;
    layer6_outputs(4874) <= b;
    layer6_outputs(4875) <= not a;
    layer6_outputs(4876) <= a;
    layer6_outputs(4877) <= not b;
    layer6_outputs(4878) <= not (a and b);
    layer6_outputs(4879) <= not b;
    layer6_outputs(4880) <= not b;
    layer6_outputs(4881) <= a;
    layer6_outputs(4882) <= not b;
    layer6_outputs(4883) <= not b;
    layer6_outputs(4884) <= b;
    layer6_outputs(4885) <= not a;
    layer6_outputs(4886) <= a and not b;
    layer6_outputs(4887) <= not a;
    layer6_outputs(4888) <= b;
    layer6_outputs(4889) <= not a;
    layer6_outputs(4890) <= a and not b;
    layer6_outputs(4891) <= a xor b;
    layer6_outputs(4892) <= not (a or b);
    layer6_outputs(4893) <= a xor b;
    layer6_outputs(4894) <= b;
    layer6_outputs(4895) <= a or b;
    layer6_outputs(4896) <= not b;
    layer6_outputs(4897) <= b and not a;
    layer6_outputs(4898) <= not b;
    layer6_outputs(4899) <= not b;
    layer6_outputs(4900) <= not b or a;
    layer6_outputs(4901) <= not b;
    layer6_outputs(4902) <= not (a and b);
    layer6_outputs(4903) <= not b;
    layer6_outputs(4904) <= a or b;
    layer6_outputs(4905) <= a xor b;
    layer6_outputs(4906) <= b;
    layer6_outputs(4907) <= not a;
    layer6_outputs(4908) <= b;
    layer6_outputs(4909) <= a xor b;
    layer6_outputs(4910) <= not a or b;
    layer6_outputs(4911) <= not b;
    layer6_outputs(4912) <= a and b;
    layer6_outputs(4913) <= not b or a;
    layer6_outputs(4914) <= b;
    layer6_outputs(4915) <= not a;
    layer6_outputs(4916) <= a and b;
    layer6_outputs(4917) <= '0';
    layer6_outputs(4918) <= not a;
    layer6_outputs(4919) <= not a or b;
    layer6_outputs(4920) <= b;
    layer6_outputs(4921) <= not a;
    layer6_outputs(4922) <= a;
    layer6_outputs(4923) <= b and not a;
    layer6_outputs(4924) <= b;
    layer6_outputs(4925) <= a;
    layer6_outputs(4926) <= a;
    layer6_outputs(4927) <= not b;
    layer6_outputs(4928) <= b and not a;
    layer6_outputs(4929) <= b;
    layer6_outputs(4930) <= not b or a;
    layer6_outputs(4931) <= a and b;
    layer6_outputs(4932) <= b;
    layer6_outputs(4933) <= not b;
    layer6_outputs(4934) <= b and not a;
    layer6_outputs(4935) <= a xor b;
    layer6_outputs(4936) <= not b;
    layer6_outputs(4937) <= a;
    layer6_outputs(4938) <= a and b;
    layer6_outputs(4939) <= not b or a;
    layer6_outputs(4940) <= not a or b;
    layer6_outputs(4941) <= not (a or b);
    layer6_outputs(4942) <= not b;
    layer6_outputs(4943) <= a;
    layer6_outputs(4944) <= not (a and b);
    layer6_outputs(4945) <= not a or b;
    layer6_outputs(4946) <= b;
    layer6_outputs(4947) <= not b or a;
    layer6_outputs(4948) <= a and b;
    layer6_outputs(4949) <= a;
    layer6_outputs(4950) <= not (a or b);
    layer6_outputs(4951) <= a xor b;
    layer6_outputs(4952) <= a;
    layer6_outputs(4953) <= not b;
    layer6_outputs(4954) <= a xor b;
    layer6_outputs(4955) <= not (a xor b);
    layer6_outputs(4956) <= a;
    layer6_outputs(4957) <= not (a or b);
    layer6_outputs(4958) <= not a;
    layer6_outputs(4959) <= b;
    layer6_outputs(4960) <= a;
    layer6_outputs(4961) <= '0';
    layer6_outputs(4962) <= '1';
    layer6_outputs(4963) <= a and b;
    layer6_outputs(4964) <= not a or b;
    layer6_outputs(4965) <= not b;
    layer6_outputs(4966) <= not a or b;
    layer6_outputs(4967) <= a and b;
    layer6_outputs(4968) <= a and b;
    layer6_outputs(4969) <= a and not b;
    layer6_outputs(4970) <= a and b;
    layer6_outputs(4971) <= a and not b;
    layer6_outputs(4972) <= not (a or b);
    layer6_outputs(4973) <= a or b;
    layer6_outputs(4974) <= a;
    layer6_outputs(4975) <= not b or a;
    layer6_outputs(4976) <= not (a and b);
    layer6_outputs(4977) <= a or b;
    layer6_outputs(4978) <= b;
    layer6_outputs(4979) <= a;
    layer6_outputs(4980) <= not a;
    layer6_outputs(4981) <= a or b;
    layer6_outputs(4982) <= a or b;
    layer6_outputs(4983) <= b;
    layer6_outputs(4984) <= not b or a;
    layer6_outputs(4985) <= a;
    layer6_outputs(4986) <= a xor b;
    layer6_outputs(4987) <= b and not a;
    layer6_outputs(4988) <= not (a or b);
    layer6_outputs(4989) <= a;
    layer6_outputs(4990) <= not b;
    layer6_outputs(4991) <= a and not b;
    layer6_outputs(4992) <= a and b;
    layer6_outputs(4993) <= a;
    layer6_outputs(4994) <= not a or b;
    layer6_outputs(4995) <= not a;
    layer6_outputs(4996) <= not (a and b);
    layer6_outputs(4997) <= not (a and b);
    layer6_outputs(4998) <= a and b;
    layer6_outputs(4999) <= not b or a;
    layer6_outputs(5000) <= a and not b;
    layer6_outputs(5001) <= a and b;
    layer6_outputs(5002) <= a;
    layer6_outputs(5003) <= a;
    layer6_outputs(5004) <= a or b;
    layer6_outputs(5005) <= not b or a;
    layer6_outputs(5006) <= b and not a;
    layer6_outputs(5007) <= a xor b;
    layer6_outputs(5008) <= a and not b;
    layer6_outputs(5009) <= not (a or b);
    layer6_outputs(5010) <= not a or b;
    layer6_outputs(5011) <= a;
    layer6_outputs(5012) <= a;
    layer6_outputs(5013) <= b;
    layer6_outputs(5014) <= b;
    layer6_outputs(5015) <= not (a and b);
    layer6_outputs(5016) <= b and not a;
    layer6_outputs(5017) <= a;
    layer6_outputs(5018) <= a xor b;
    layer6_outputs(5019) <= b;
    layer6_outputs(5020) <= a;
    layer6_outputs(5021) <= b;
    layer6_outputs(5022) <= not (a or b);
    layer6_outputs(5023) <= not (a or b);
    layer6_outputs(5024) <= a;
    layer6_outputs(5025) <= not a or b;
    layer6_outputs(5026) <= not (a xor b);
    layer6_outputs(5027) <= not a;
    layer6_outputs(5028) <= a;
    layer6_outputs(5029) <= a and b;
    layer6_outputs(5030) <= a or b;
    layer6_outputs(5031) <= not (a and b);
    layer6_outputs(5032) <= not a;
    layer6_outputs(5033) <= b;
    layer6_outputs(5034) <= a;
    layer6_outputs(5035) <= not a;
    layer6_outputs(5036) <= not (a and b);
    layer6_outputs(5037) <= not b;
    layer6_outputs(5038) <= a and not b;
    layer6_outputs(5039) <= not b;
    layer6_outputs(5040) <= not a;
    layer6_outputs(5041) <= a and b;
    layer6_outputs(5042) <= not (a and b);
    layer6_outputs(5043) <= not a;
    layer6_outputs(5044) <= not b;
    layer6_outputs(5045) <= a;
    layer6_outputs(5046) <= not b;
    layer6_outputs(5047) <= not (a xor b);
    layer6_outputs(5048) <= not b or a;
    layer6_outputs(5049) <= a;
    layer6_outputs(5050) <= b;
    layer6_outputs(5051) <= not (a or b);
    layer6_outputs(5052) <= not (a or b);
    layer6_outputs(5053) <= not (a or b);
    layer6_outputs(5054) <= a and b;
    layer6_outputs(5055) <= a;
    layer6_outputs(5056) <= not b;
    layer6_outputs(5057) <= a and not b;
    layer6_outputs(5058) <= not a;
    layer6_outputs(5059) <= not b or a;
    layer6_outputs(5060) <= not a or b;
    layer6_outputs(5061) <= b and not a;
    layer6_outputs(5062) <= a xor b;
    layer6_outputs(5063) <= not (a xor b);
    layer6_outputs(5064) <= a and not b;
    layer6_outputs(5065) <= '1';
    layer6_outputs(5066) <= not (a and b);
    layer6_outputs(5067) <= a;
    layer6_outputs(5068) <= a;
    layer6_outputs(5069) <= not (a or b);
    layer6_outputs(5070) <= b;
    layer6_outputs(5071) <= a and b;
    layer6_outputs(5072) <= not b;
    layer6_outputs(5073) <= a xor b;
    layer6_outputs(5074) <= not b or a;
    layer6_outputs(5075) <= not b;
    layer6_outputs(5076) <= not a or b;
    layer6_outputs(5077) <= not a or b;
    layer6_outputs(5078) <= not (a xor b);
    layer6_outputs(5079) <= a xor b;
    layer6_outputs(5080) <= not a;
    layer6_outputs(5081) <= a or b;
    layer6_outputs(5082) <= a xor b;
    layer6_outputs(5083) <= a;
    layer6_outputs(5084) <= a and not b;
    layer6_outputs(5085) <= not a or b;
    layer6_outputs(5086) <= not a;
    layer6_outputs(5087) <= b;
    layer6_outputs(5088) <= a;
    layer6_outputs(5089) <= not a;
    layer6_outputs(5090) <= b;
    layer6_outputs(5091) <= not a or b;
    layer6_outputs(5092) <= a xor b;
    layer6_outputs(5093) <= a or b;
    layer6_outputs(5094) <= not a;
    layer6_outputs(5095) <= not (a or b);
    layer6_outputs(5096) <= not (a and b);
    layer6_outputs(5097) <= a xor b;
    layer6_outputs(5098) <= a and b;
    layer6_outputs(5099) <= not a;
    layer6_outputs(5100) <= a and b;
    layer6_outputs(5101) <= not a or b;
    layer6_outputs(5102) <= b;
    layer6_outputs(5103) <= not a;
    layer6_outputs(5104) <= not (a and b);
    layer6_outputs(5105) <= not (a xor b);
    layer6_outputs(5106) <= not (a xor b);
    layer6_outputs(5107) <= b;
    layer6_outputs(5108) <= not a;
    layer6_outputs(5109) <= not a;
    layer6_outputs(5110) <= a;
    layer6_outputs(5111) <= a or b;
    layer6_outputs(5112) <= not b or a;
    layer6_outputs(5113) <= b and not a;
    layer6_outputs(5114) <= not b;
    layer6_outputs(5115) <= a and b;
    layer6_outputs(5116) <= b and not a;
    layer6_outputs(5117) <= not (a or b);
    layer6_outputs(5118) <= not a;
    layer6_outputs(5119) <= a;
    layer7_outputs(0) <= not (a xor b);
    layer7_outputs(1) <= not a or b;
    layer7_outputs(2) <= a and not b;
    layer7_outputs(3) <= a and b;
    layer7_outputs(4) <= not a;
    layer7_outputs(5) <= not (a or b);
    layer7_outputs(6) <= b;
    layer7_outputs(7) <= a and b;
    layer7_outputs(8) <= not (a or b);
    layer7_outputs(9) <= not (a and b);
    layer7_outputs(10) <= not b;
    layer7_outputs(11) <= a or b;
    layer7_outputs(12) <= b and not a;
    layer7_outputs(13) <= not a;
    layer7_outputs(14) <= a xor b;
    layer7_outputs(15) <= not b;
    layer7_outputs(16) <= not b or a;
    layer7_outputs(17) <= a or b;
    layer7_outputs(18) <= a and b;
    layer7_outputs(19) <= '1';
    layer7_outputs(20) <= a or b;
    layer7_outputs(21) <= not a;
    layer7_outputs(22) <= not b;
    layer7_outputs(23) <= not a;
    layer7_outputs(24) <= not a;
    layer7_outputs(25) <= not b;
    layer7_outputs(26) <= not b;
    layer7_outputs(27) <= '0';
    layer7_outputs(28) <= not b;
    layer7_outputs(29) <= a xor b;
    layer7_outputs(30) <= not (a xor b);
    layer7_outputs(31) <= b;
    layer7_outputs(32) <= not b;
    layer7_outputs(33) <= a xor b;
    layer7_outputs(34) <= a and not b;
    layer7_outputs(35) <= a xor b;
    layer7_outputs(36) <= a and b;
    layer7_outputs(37) <= not (a and b);
    layer7_outputs(38) <= not (a or b);
    layer7_outputs(39) <= b;
    layer7_outputs(40) <= not a;
    layer7_outputs(41) <= not b or a;
    layer7_outputs(42) <= b and not a;
    layer7_outputs(43) <= not a or b;
    layer7_outputs(44) <= a and b;
    layer7_outputs(45) <= a or b;
    layer7_outputs(46) <= not a;
    layer7_outputs(47) <= not (a and b);
    layer7_outputs(48) <= not a or b;
    layer7_outputs(49) <= a xor b;
    layer7_outputs(50) <= b and not a;
    layer7_outputs(51) <= not (a or b);
    layer7_outputs(52) <= not b or a;
    layer7_outputs(53) <= not b;
    layer7_outputs(54) <= not (a or b);
    layer7_outputs(55) <= a;
    layer7_outputs(56) <= not b;
    layer7_outputs(57) <= not a;
    layer7_outputs(58) <= a and b;
    layer7_outputs(59) <= b;
    layer7_outputs(60) <= not a;
    layer7_outputs(61) <= not a;
    layer7_outputs(62) <= a;
    layer7_outputs(63) <= b;
    layer7_outputs(64) <= a and b;
    layer7_outputs(65) <= not a;
    layer7_outputs(66) <= not (a xor b);
    layer7_outputs(67) <= b and not a;
    layer7_outputs(68) <= a;
    layer7_outputs(69) <= not b;
    layer7_outputs(70) <= not b;
    layer7_outputs(71) <= not (a and b);
    layer7_outputs(72) <= not a;
    layer7_outputs(73) <= a;
    layer7_outputs(74) <= b;
    layer7_outputs(75) <= b and not a;
    layer7_outputs(76) <= not b;
    layer7_outputs(77) <= not a;
    layer7_outputs(78) <= not a;
    layer7_outputs(79) <= not b;
    layer7_outputs(80) <= a;
    layer7_outputs(81) <= not a or b;
    layer7_outputs(82) <= not (a and b);
    layer7_outputs(83) <= a or b;
    layer7_outputs(84) <= '0';
    layer7_outputs(85) <= not (a or b);
    layer7_outputs(86) <= not b;
    layer7_outputs(87) <= a xor b;
    layer7_outputs(88) <= not a;
    layer7_outputs(89) <= a or b;
    layer7_outputs(90) <= a;
    layer7_outputs(91) <= a and b;
    layer7_outputs(92) <= not (a xor b);
    layer7_outputs(93) <= not b;
    layer7_outputs(94) <= a and not b;
    layer7_outputs(95) <= not (a or b);
    layer7_outputs(96) <= not a;
    layer7_outputs(97) <= not a;
    layer7_outputs(98) <= b and not a;
    layer7_outputs(99) <= a and b;
    layer7_outputs(100) <= b;
    layer7_outputs(101) <= not b or a;
    layer7_outputs(102) <= a xor b;
    layer7_outputs(103) <= not a;
    layer7_outputs(104) <= a xor b;
    layer7_outputs(105) <= b;
    layer7_outputs(106) <= not b;
    layer7_outputs(107) <= b;
    layer7_outputs(108) <= not (a xor b);
    layer7_outputs(109) <= not a or b;
    layer7_outputs(110) <= a and not b;
    layer7_outputs(111) <= a xor b;
    layer7_outputs(112) <= not b or a;
    layer7_outputs(113) <= not a;
    layer7_outputs(114) <= '1';
    layer7_outputs(115) <= not a;
    layer7_outputs(116) <= not a;
    layer7_outputs(117) <= not (a xor b);
    layer7_outputs(118) <= not a or b;
    layer7_outputs(119) <= a xor b;
    layer7_outputs(120) <= not (a or b);
    layer7_outputs(121) <= not (a and b);
    layer7_outputs(122) <= a;
    layer7_outputs(123) <= a or b;
    layer7_outputs(124) <= not a;
    layer7_outputs(125) <= not b;
    layer7_outputs(126) <= b and not a;
    layer7_outputs(127) <= a xor b;
    layer7_outputs(128) <= not b;
    layer7_outputs(129) <= not b or a;
    layer7_outputs(130) <= a and not b;
    layer7_outputs(131) <= b and not a;
    layer7_outputs(132) <= b;
    layer7_outputs(133) <= not a or b;
    layer7_outputs(134) <= a xor b;
    layer7_outputs(135) <= not b;
    layer7_outputs(136) <= a xor b;
    layer7_outputs(137) <= not (a xor b);
    layer7_outputs(138) <= b and not a;
    layer7_outputs(139) <= a;
    layer7_outputs(140) <= a;
    layer7_outputs(141) <= not b or a;
    layer7_outputs(142) <= b;
    layer7_outputs(143) <= not (a xor b);
    layer7_outputs(144) <= not b or a;
    layer7_outputs(145) <= b;
    layer7_outputs(146) <= not a or b;
    layer7_outputs(147) <= not b or a;
    layer7_outputs(148) <= not (a xor b);
    layer7_outputs(149) <= not (a and b);
    layer7_outputs(150) <= not b;
    layer7_outputs(151) <= not b or a;
    layer7_outputs(152) <= a and not b;
    layer7_outputs(153) <= a;
    layer7_outputs(154) <= not b;
    layer7_outputs(155) <= not (a xor b);
    layer7_outputs(156) <= a;
    layer7_outputs(157) <= not (a xor b);
    layer7_outputs(158) <= not b;
    layer7_outputs(159) <= b;
    layer7_outputs(160) <= a and b;
    layer7_outputs(161) <= b;
    layer7_outputs(162) <= not b or a;
    layer7_outputs(163) <= not (a or b);
    layer7_outputs(164) <= not a or b;
    layer7_outputs(165) <= not b;
    layer7_outputs(166) <= b;
    layer7_outputs(167) <= a;
    layer7_outputs(168) <= a or b;
    layer7_outputs(169) <= not (a or b);
    layer7_outputs(170) <= a and not b;
    layer7_outputs(171) <= not a;
    layer7_outputs(172) <= a;
    layer7_outputs(173) <= not (a xor b);
    layer7_outputs(174) <= not b;
    layer7_outputs(175) <= not b;
    layer7_outputs(176) <= not (a xor b);
    layer7_outputs(177) <= not a or b;
    layer7_outputs(178) <= b;
    layer7_outputs(179) <= a;
    layer7_outputs(180) <= b;
    layer7_outputs(181) <= a;
    layer7_outputs(182) <= a or b;
    layer7_outputs(183) <= not a;
    layer7_outputs(184) <= a or b;
    layer7_outputs(185) <= not (a and b);
    layer7_outputs(186) <= not (a or b);
    layer7_outputs(187) <= not (a xor b);
    layer7_outputs(188) <= not a;
    layer7_outputs(189) <= a;
    layer7_outputs(190) <= a xor b;
    layer7_outputs(191) <= not b;
    layer7_outputs(192) <= not a or b;
    layer7_outputs(193) <= a or b;
    layer7_outputs(194) <= b;
    layer7_outputs(195) <= a;
    layer7_outputs(196) <= not b or a;
    layer7_outputs(197) <= not a;
    layer7_outputs(198) <= a;
    layer7_outputs(199) <= not a or b;
    layer7_outputs(200) <= b and not a;
    layer7_outputs(201) <= not b;
    layer7_outputs(202) <= a;
    layer7_outputs(203) <= a and b;
    layer7_outputs(204) <= not a or b;
    layer7_outputs(205) <= b;
    layer7_outputs(206) <= not (a or b);
    layer7_outputs(207) <= b;
    layer7_outputs(208) <= not b;
    layer7_outputs(209) <= not a;
    layer7_outputs(210) <= a and b;
    layer7_outputs(211) <= not b;
    layer7_outputs(212) <= not (a xor b);
    layer7_outputs(213) <= b;
    layer7_outputs(214) <= b and not a;
    layer7_outputs(215) <= '0';
    layer7_outputs(216) <= not b or a;
    layer7_outputs(217) <= not a;
    layer7_outputs(218) <= not a or b;
    layer7_outputs(219) <= not (a or b);
    layer7_outputs(220) <= '0';
    layer7_outputs(221) <= a xor b;
    layer7_outputs(222) <= a or b;
    layer7_outputs(223) <= not (a or b);
    layer7_outputs(224) <= b;
    layer7_outputs(225) <= not (a and b);
    layer7_outputs(226) <= not (a xor b);
    layer7_outputs(227) <= not (a or b);
    layer7_outputs(228) <= a or b;
    layer7_outputs(229) <= not a;
    layer7_outputs(230) <= not a;
    layer7_outputs(231) <= a or b;
    layer7_outputs(232) <= a and not b;
    layer7_outputs(233) <= not b;
    layer7_outputs(234) <= a and not b;
    layer7_outputs(235) <= not b or a;
    layer7_outputs(236) <= a and b;
    layer7_outputs(237) <= a and not b;
    layer7_outputs(238) <= not a;
    layer7_outputs(239) <= not (a or b);
    layer7_outputs(240) <= a and not b;
    layer7_outputs(241) <= not b or a;
    layer7_outputs(242) <= not (a and b);
    layer7_outputs(243) <= b;
    layer7_outputs(244) <= a xor b;
    layer7_outputs(245) <= not a;
    layer7_outputs(246) <= a or b;
    layer7_outputs(247) <= a and not b;
    layer7_outputs(248) <= a and b;
    layer7_outputs(249) <= not a;
    layer7_outputs(250) <= not b;
    layer7_outputs(251) <= b and not a;
    layer7_outputs(252) <= not a;
    layer7_outputs(253) <= not a;
    layer7_outputs(254) <= not a or b;
    layer7_outputs(255) <= a;
    layer7_outputs(256) <= not b;
    layer7_outputs(257) <= not b;
    layer7_outputs(258) <= not b;
    layer7_outputs(259) <= not (a and b);
    layer7_outputs(260) <= not b;
    layer7_outputs(261) <= not b;
    layer7_outputs(262) <= not a or b;
    layer7_outputs(263) <= a;
    layer7_outputs(264) <= not (a and b);
    layer7_outputs(265) <= not b;
    layer7_outputs(266) <= not (a or b);
    layer7_outputs(267) <= not b;
    layer7_outputs(268) <= not b;
    layer7_outputs(269) <= a xor b;
    layer7_outputs(270) <= a;
    layer7_outputs(271) <= b;
    layer7_outputs(272) <= a or b;
    layer7_outputs(273) <= not (a or b);
    layer7_outputs(274) <= a;
    layer7_outputs(275) <= a and b;
    layer7_outputs(276) <= not b;
    layer7_outputs(277) <= a;
    layer7_outputs(278) <= a xor b;
    layer7_outputs(279) <= a and b;
    layer7_outputs(280) <= a;
    layer7_outputs(281) <= not b or a;
    layer7_outputs(282) <= a and b;
    layer7_outputs(283) <= not (a xor b);
    layer7_outputs(284) <= not (a and b);
    layer7_outputs(285) <= '0';
    layer7_outputs(286) <= a and not b;
    layer7_outputs(287) <= a;
    layer7_outputs(288) <= b;
    layer7_outputs(289) <= a or b;
    layer7_outputs(290) <= not (a xor b);
    layer7_outputs(291) <= a;
    layer7_outputs(292) <= not b;
    layer7_outputs(293) <= a xor b;
    layer7_outputs(294) <= a and not b;
    layer7_outputs(295) <= a or b;
    layer7_outputs(296) <= a and not b;
    layer7_outputs(297) <= a xor b;
    layer7_outputs(298) <= a xor b;
    layer7_outputs(299) <= a;
    layer7_outputs(300) <= not (a or b);
    layer7_outputs(301) <= a and b;
    layer7_outputs(302) <= b;
    layer7_outputs(303) <= not (a or b);
    layer7_outputs(304) <= not a;
    layer7_outputs(305) <= not b;
    layer7_outputs(306) <= a;
    layer7_outputs(307) <= not a or b;
    layer7_outputs(308) <= not (a and b);
    layer7_outputs(309) <= b;
    layer7_outputs(310) <= not b;
    layer7_outputs(311) <= a;
    layer7_outputs(312) <= not b;
    layer7_outputs(313) <= not a;
    layer7_outputs(314) <= not a;
    layer7_outputs(315) <= not a or b;
    layer7_outputs(316) <= not a or b;
    layer7_outputs(317) <= not b;
    layer7_outputs(318) <= not (a and b);
    layer7_outputs(319) <= a;
    layer7_outputs(320) <= not b;
    layer7_outputs(321) <= a;
    layer7_outputs(322) <= not (a or b);
    layer7_outputs(323) <= not b;
    layer7_outputs(324) <= b and not a;
    layer7_outputs(325) <= not (a and b);
    layer7_outputs(326) <= a xor b;
    layer7_outputs(327) <= not (a xor b);
    layer7_outputs(328) <= not a;
    layer7_outputs(329) <= a xor b;
    layer7_outputs(330) <= a xor b;
    layer7_outputs(331) <= not a;
    layer7_outputs(332) <= not a;
    layer7_outputs(333) <= not (a or b);
    layer7_outputs(334) <= not b;
    layer7_outputs(335) <= not b;
    layer7_outputs(336) <= not a;
    layer7_outputs(337) <= not (a or b);
    layer7_outputs(338) <= b;
    layer7_outputs(339) <= b;
    layer7_outputs(340) <= not a;
    layer7_outputs(341) <= b;
    layer7_outputs(342) <= not (a or b);
    layer7_outputs(343) <= a;
    layer7_outputs(344) <= not b;
    layer7_outputs(345) <= b;
    layer7_outputs(346) <= a xor b;
    layer7_outputs(347) <= not b;
    layer7_outputs(348) <= not b;
    layer7_outputs(349) <= not a;
    layer7_outputs(350) <= not a;
    layer7_outputs(351) <= '1';
    layer7_outputs(352) <= not a or b;
    layer7_outputs(353) <= not a;
    layer7_outputs(354) <= a;
    layer7_outputs(355) <= not (a and b);
    layer7_outputs(356) <= not (a or b);
    layer7_outputs(357) <= b and not a;
    layer7_outputs(358) <= not a or b;
    layer7_outputs(359) <= a xor b;
    layer7_outputs(360) <= a;
    layer7_outputs(361) <= not a;
    layer7_outputs(362) <= b;
    layer7_outputs(363) <= not (a or b);
    layer7_outputs(364) <= not a;
    layer7_outputs(365) <= a or b;
    layer7_outputs(366) <= not b or a;
    layer7_outputs(367) <= a and not b;
    layer7_outputs(368) <= not a;
    layer7_outputs(369) <= a and b;
    layer7_outputs(370) <= not a;
    layer7_outputs(371) <= not (a xor b);
    layer7_outputs(372) <= not (a xor b);
    layer7_outputs(373) <= not (a or b);
    layer7_outputs(374) <= b;
    layer7_outputs(375) <= a and b;
    layer7_outputs(376) <= not (a or b);
    layer7_outputs(377) <= b;
    layer7_outputs(378) <= a;
    layer7_outputs(379) <= '1';
    layer7_outputs(380) <= not (a and b);
    layer7_outputs(381) <= not b;
    layer7_outputs(382) <= a and b;
    layer7_outputs(383) <= a;
    layer7_outputs(384) <= a;
    layer7_outputs(385) <= b;
    layer7_outputs(386) <= b;
    layer7_outputs(387) <= not b;
    layer7_outputs(388) <= not (a xor b);
    layer7_outputs(389) <= not a;
    layer7_outputs(390) <= a xor b;
    layer7_outputs(391) <= not b or a;
    layer7_outputs(392) <= a;
    layer7_outputs(393) <= not (a xor b);
    layer7_outputs(394) <= not (a xor b);
    layer7_outputs(395) <= a;
    layer7_outputs(396) <= '0';
    layer7_outputs(397) <= not (a and b);
    layer7_outputs(398) <= not b;
    layer7_outputs(399) <= b and not a;
    layer7_outputs(400) <= not a;
    layer7_outputs(401) <= not a or b;
    layer7_outputs(402) <= a xor b;
    layer7_outputs(403) <= not (a and b);
    layer7_outputs(404) <= not a;
    layer7_outputs(405) <= not a;
    layer7_outputs(406) <= a;
    layer7_outputs(407) <= b and not a;
    layer7_outputs(408) <= a or b;
    layer7_outputs(409) <= not (a xor b);
    layer7_outputs(410) <= b;
    layer7_outputs(411) <= a xor b;
    layer7_outputs(412) <= not (a or b);
    layer7_outputs(413) <= '1';
    layer7_outputs(414) <= not a or b;
    layer7_outputs(415) <= a and not b;
    layer7_outputs(416) <= a xor b;
    layer7_outputs(417) <= b;
    layer7_outputs(418) <= a;
    layer7_outputs(419) <= not (a and b);
    layer7_outputs(420) <= not (a and b);
    layer7_outputs(421) <= a xor b;
    layer7_outputs(422) <= not b;
    layer7_outputs(423) <= not (a or b);
    layer7_outputs(424) <= a;
    layer7_outputs(425) <= a xor b;
    layer7_outputs(426) <= a xor b;
    layer7_outputs(427) <= not (a xor b);
    layer7_outputs(428) <= b and not a;
    layer7_outputs(429) <= b and not a;
    layer7_outputs(430) <= not b or a;
    layer7_outputs(431) <= not (a xor b);
    layer7_outputs(432) <= not a;
    layer7_outputs(433) <= a xor b;
    layer7_outputs(434) <= not b;
    layer7_outputs(435) <= not (a or b);
    layer7_outputs(436) <= b;
    layer7_outputs(437) <= not b;
    layer7_outputs(438) <= b and not a;
    layer7_outputs(439) <= not a;
    layer7_outputs(440) <= a and not b;
    layer7_outputs(441) <= a xor b;
    layer7_outputs(442) <= a;
    layer7_outputs(443) <= a;
    layer7_outputs(444) <= not a;
    layer7_outputs(445) <= not a or b;
    layer7_outputs(446) <= a;
    layer7_outputs(447) <= not (a or b);
    layer7_outputs(448) <= a;
    layer7_outputs(449) <= a;
    layer7_outputs(450) <= not (a xor b);
    layer7_outputs(451) <= not a;
    layer7_outputs(452) <= a xor b;
    layer7_outputs(453) <= not a;
    layer7_outputs(454) <= a;
    layer7_outputs(455) <= b;
    layer7_outputs(456) <= not (a xor b);
    layer7_outputs(457) <= not b;
    layer7_outputs(458) <= a or b;
    layer7_outputs(459) <= not b;
    layer7_outputs(460) <= b;
    layer7_outputs(461) <= not a or b;
    layer7_outputs(462) <= not b;
    layer7_outputs(463) <= a xor b;
    layer7_outputs(464) <= not (a or b);
    layer7_outputs(465) <= not b;
    layer7_outputs(466) <= b;
    layer7_outputs(467) <= b;
    layer7_outputs(468) <= not b;
    layer7_outputs(469) <= a;
    layer7_outputs(470) <= not b;
    layer7_outputs(471) <= '1';
    layer7_outputs(472) <= not (a xor b);
    layer7_outputs(473) <= a;
    layer7_outputs(474) <= a or b;
    layer7_outputs(475) <= a;
    layer7_outputs(476) <= a and b;
    layer7_outputs(477) <= not b;
    layer7_outputs(478) <= not (a xor b);
    layer7_outputs(479) <= not (a or b);
    layer7_outputs(480) <= not (a xor b);
    layer7_outputs(481) <= not b or a;
    layer7_outputs(482) <= b;
    layer7_outputs(483) <= not b;
    layer7_outputs(484) <= not b;
    layer7_outputs(485) <= a and not b;
    layer7_outputs(486) <= not b;
    layer7_outputs(487) <= not a;
    layer7_outputs(488) <= not b or a;
    layer7_outputs(489) <= not b or a;
    layer7_outputs(490) <= b;
    layer7_outputs(491) <= not b;
    layer7_outputs(492) <= not a or b;
    layer7_outputs(493) <= not b or a;
    layer7_outputs(494) <= a and b;
    layer7_outputs(495) <= not b;
    layer7_outputs(496) <= a;
    layer7_outputs(497) <= b;
    layer7_outputs(498) <= not b;
    layer7_outputs(499) <= b;
    layer7_outputs(500) <= not (a xor b);
    layer7_outputs(501) <= not a;
    layer7_outputs(502) <= b;
    layer7_outputs(503) <= b;
    layer7_outputs(504) <= not (a or b);
    layer7_outputs(505) <= a or b;
    layer7_outputs(506) <= not (a xor b);
    layer7_outputs(507) <= a;
    layer7_outputs(508) <= a xor b;
    layer7_outputs(509) <= a or b;
    layer7_outputs(510) <= a and b;
    layer7_outputs(511) <= a;
    layer7_outputs(512) <= a;
    layer7_outputs(513) <= a xor b;
    layer7_outputs(514) <= b;
    layer7_outputs(515) <= b;
    layer7_outputs(516) <= b and not a;
    layer7_outputs(517) <= not (a xor b);
    layer7_outputs(518) <= b;
    layer7_outputs(519) <= not b or a;
    layer7_outputs(520) <= not a or b;
    layer7_outputs(521) <= a xor b;
    layer7_outputs(522) <= not (a or b);
    layer7_outputs(523) <= b and not a;
    layer7_outputs(524) <= a or b;
    layer7_outputs(525) <= a and not b;
    layer7_outputs(526) <= not a or b;
    layer7_outputs(527) <= a;
    layer7_outputs(528) <= a xor b;
    layer7_outputs(529) <= a or b;
    layer7_outputs(530) <= a;
    layer7_outputs(531) <= b;
    layer7_outputs(532) <= b;
    layer7_outputs(533) <= not (a or b);
    layer7_outputs(534) <= a or b;
    layer7_outputs(535) <= a;
    layer7_outputs(536) <= b and not a;
    layer7_outputs(537) <= not (a xor b);
    layer7_outputs(538) <= b;
    layer7_outputs(539) <= not a;
    layer7_outputs(540) <= not (a and b);
    layer7_outputs(541) <= not b;
    layer7_outputs(542) <= a xor b;
    layer7_outputs(543) <= a;
    layer7_outputs(544) <= b;
    layer7_outputs(545) <= b and not a;
    layer7_outputs(546) <= not b;
    layer7_outputs(547) <= a;
    layer7_outputs(548) <= a xor b;
    layer7_outputs(549) <= b;
    layer7_outputs(550) <= b and not a;
    layer7_outputs(551) <= '0';
    layer7_outputs(552) <= a and b;
    layer7_outputs(553) <= a or b;
    layer7_outputs(554) <= a;
    layer7_outputs(555) <= '1';
    layer7_outputs(556) <= not a;
    layer7_outputs(557) <= b;
    layer7_outputs(558) <= a;
    layer7_outputs(559) <= a;
    layer7_outputs(560) <= not a;
    layer7_outputs(561) <= not a or b;
    layer7_outputs(562) <= a;
    layer7_outputs(563) <= a;
    layer7_outputs(564) <= a or b;
    layer7_outputs(565) <= b;
    layer7_outputs(566) <= a and not b;
    layer7_outputs(567) <= a and not b;
    layer7_outputs(568) <= '1';
    layer7_outputs(569) <= not (a and b);
    layer7_outputs(570) <= not (a xor b);
    layer7_outputs(571) <= b;
    layer7_outputs(572) <= a;
    layer7_outputs(573) <= a and b;
    layer7_outputs(574) <= not b;
    layer7_outputs(575) <= a and b;
    layer7_outputs(576) <= not (a and b);
    layer7_outputs(577) <= a;
    layer7_outputs(578) <= not (a and b);
    layer7_outputs(579) <= a and b;
    layer7_outputs(580) <= a xor b;
    layer7_outputs(581) <= not (a xor b);
    layer7_outputs(582) <= not (a or b);
    layer7_outputs(583) <= not a;
    layer7_outputs(584) <= b;
    layer7_outputs(585) <= not a;
    layer7_outputs(586) <= a or b;
    layer7_outputs(587) <= a and not b;
    layer7_outputs(588) <= b and not a;
    layer7_outputs(589) <= a xor b;
    layer7_outputs(590) <= not (a and b);
    layer7_outputs(591) <= not b or a;
    layer7_outputs(592) <= a;
    layer7_outputs(593) <= a;
    layer7_outputs(594) <= not (a xor b);
    layer7_outputs(595) <= a or b;
    layer7_outputs(596) <= not b;
    layer7_outputs(597) <= '0';
    layer7_outputs(598) <= not b;
    layer7_outputs(599) <= not b or a;
    layer7_outputs(600) <= not b;
    layer7_outputs(601) <= not b;
    layer7_outputs(602) <= a or b;
    layer7_outputs(603) <= not b;
    layer7_outputs(604) <= a xor b;
    layer7_outputs(605) <= a;
    layer7_outputs(606) <= not a;
    layer7_outputs(607) <= a and not b;
    layer7_outputs(608) <= not a or b;
    layer7_outputs(609) <= '1';
    layer7_outputs(610) <= not b;
    layer7_outputs(611) <= b and not a;
    layer7_outputs(612) <= b;
    layer7_outputs(613) <= a xor b;
    layer7_outputs(614) <= not a;
    layer7_outputs(615) <= not b;
    layer7_outputs(616) <= a;
    layer7_outputs(617) <= not b or a;
    layer7_outputs(618) <= not b;
    layer7_outputs(619) <= b;
    layer7_outputs(620) <= b;
    layer7_outputs(621) <= not a;
    layer7_outputs(622) <= b;
    layer7_outputs(623) <= not (a and b);
    layer7_outputs(624) <= not a or b;
    layer7_outputs(625) <= a and not b;
    layer7_outputs(626) <= '1';
    layer7_outputs(627) <= b;
    layer7_outputs(628) <= a xor b;
    layer7_outputs(629) <= b;
    layer7_outputs(630) <= a;
    layer7_outputs(631) <= not b;
    layer7_outputs(632) <= not (a and b);
    layer7_outputs(633) <= not (a and b);
    layer7_outputs(634) <= a or b;
    layer7_outputs(635) <= b;
    layer7_outputs(636) <= a and b;
    layer7_outputs(637) <= not a;
    layer7_outputs(638) <= not (a or b);
    layer7_outputs(639) <= b and not a;
    layer7_outputs(640) <= b;
    layer7_outputs(641) <= not (a xor b);
    layer7_outputs(642) <= not a or b;
    layer7_outputs(643) <= not (a xor b);
    layer7_outputs(644) <= b;
    layer7_outputs(645) <= a xor b;
    layer7_outputs(646) <= b and not a;
    layer7_outputs(647) <= a xor b;
    layer7_outputs(648) <= a xor b;
    layer7_outputs(649) <= a and b;
    layer7_outputs(650) <= not a;
    layer7_outputs(651) <= a and b;
    layer7_outputs(652) <= not b or a;
    layer7_outputs(653) <= a or b;
    layer7_outputs(654) <= not (a xor b);
    layer7_outputs(655) <= a and b;
    layer7_outputs(656) <= not b;
    layer7_outputs(657) <= not (a xor b);
    layer7_outputs(658) <= not (a xor b);
    layer7_outputs(659) <= not a;
    layer7_outputs(660) <= not (a xor b);
    layer7_outputs(661) <= a or b;
    layer7_outputs(662) <= not a;
    layer7_outputs(663) <= b;
    layer7_outputs(664) <= a and not b;
    layer7_outputs(665) <= not b;
    layer7_outputs(666) <= b;
    layer7_outputs(667) <= a;
    layer7_outputs(668) <= a;
    layer7_outputs(669) <= not b or a;
    layer7_outputs(670) <= a or b;
    layer7_outputs(671) <= a;
    layer7_outputs(672) <= not a;
    layer7_outputs(673) <= a and not b;
    layer7_outputs(674) <= not b;
    layer7_outputs(675) <= not (a and b);
    layer7_outputs(676) <= a or b;
    layer7_outputs(677) <= a or b;
    layer7_outputs(678) <= a and not b;
    layer7_outputs(679) <= not (a xor b);
    layer7_outputs(680) <= a;
    layer7_outputs(681) <= a xor b;
    layer7_outputs(682) <= b and not a;
    layer7_outputs(683) <= not b;
    layer7_outputs(684) <= a;
    layer7_outputs(685) <= a and b;
    layer7_outputs(686) <= a and b;
    layer7_outputs(687) <= a xor b;
    layer7_outputs(688) <= not b;
    layer7_outputs(689) <= b;
    layer7_outputs(690) <= not a;
    layer7_outputs(691) <= not a or b;
    layer7_outputs(692) <= not (a or b);
    layer7_outputs(693) <= not a;
    layer7_outputs(694) <= not a or b;
    layer7_outputs(695) <= not b;
    layer7_outputs(696) <= a and b;
    layer7_outputs(697) <= not (a xor b);
    layer7_outputs(698) <= b;
    layer7_outputs(699) <= a and b;
    layer7_outputs(700) <= a and not b;
    layer7_outputs(701) <= a xor b;
    layer7_outputs(702) <= a;
    layer7_outputs(703) <= not (a xor b);
    layer7_outputs(704) <= a and not b;
    layer7_outputs(705) <= a and not b;
    layer7_outputs(706) <= a or b;
    layer7_outputs(707) <= a and not b;
    layer7_outputs(708) <= a;
    layer7_outputs(709) <= a xor b;
    layer7_outputs(710) <= not (a or b);
    layer7_outputs(711) <= a xor b;
    layer7_outputs(712) <= a;
    layer7_outputs(713) <= not b;
    layer7_outputs(714) <= not (a xor b);
    layer7_outputs(715) <= not a;
    layer7_outputs(716) <= not (a or b);
    layer7_outputs(717) <= a xor b;
    layer7_outputs(718) <= not a;
    layer7_outputs(719) <= not a;
    layer7_outputs(720) <= not b;
    layer7_outputs(721) <= not a;
    layer7_outputs(722) <= a xor b;
    layer7_outputs(723) <= a and not b;
    layer7_outputs(724) <= a xor b;
    layer7_outputs(725) <= not a;
    layer7_outputs(726) <= a xor b;
    layer7_outputs(727) <= b;
    layer7_outputs(728) <= not (a xor b);
    layer7_outputs(729) <= a;
    layer7_outputs(730) <= b;
    layer7_outputs(731) <= not (a or b);
    layer7_outputs(732) <= not b or a;
    layer7_outputs(733) <= a and not b;
    layer7_outputs(734) <= not (a xor b);
    layer7_outputs(735) <= a and not b;
    layer7_outputs(736) <= b;
    layer7_outputs(737) <= a and not b;
    layer7_outputs(738) <= not b;
    layer7_outputs(739) <= a;
    layer7_outputs(740) <= not (a or b);
    layer7_outputs(741) <= not (a and b);
    layer7_outputs(742) <= not a;
    layer7_outputs(743) <= a;
    layer7_outputs(744) <= not b;
    layer7_outputs(745) <= a and b;
    layer7_outputs(746) <= not a or b;
    layer7_outputs(747) <= not b or a;
    layer7_outputs(748) <= not a;
    layer7_outputs(749) <= not a or b;
    layer7_outputs(750) <= '0';
    layer7_outputs(751) <= b;
    layer7_outputs(752) <= not (a xor b);
    layer7_outputs(753) <= not a or b;
    layer7_outputs(754) <= not b;
    layer7_outputs(755) <= a xor b;
    layer7_outputs(756) <= not b;
    layer7_outputs(757) <= not b or a;
    layer7_outputs(758) <= a and b;
    layer7_outputs(759) <= not a or b;
    layer7_outputs(760) <= not b or a;
    layer7_outputs(761) <= not a;
    layer7_outputs(762) <= not (a xor b);
    layer7_outputs(763) <= not b or a;
    layer7_outputs(764) <= a or b;
    layer7_outputs(765) <= not (a or b);
    layer7_outputs(766) <= not a;
    layer7_outputs(767) <= not b or a;
    layer7_outputs(768) <= b;
    layer7_outputs(769) <= a;
    layer7_outputs(770) <= '1';
    layer7_outputs(771) <= '1';
    layer7_outputs(772) <= not a;
    layer7_outputs(773) <= '1';
    layer7_outputs(774) <= b;
    layer7_outputs(775) <= a;
    layer7_outputs(776) <= a xor b;
    layer7_outputs(777) <= not b;
    layer7_outputs(778) <= a;
    layer7_outputs(779) <= not (a or b);
    layer7_outputs(780) <= a;
    layer7_outputs(781) <= not a;
    layer7_outputs(782) <= not a;
    layer7_outputs(783) <= not b;
    layer7_outputs(784) <= not (a xor b);
    layer7_outputs(785) <= a xor b;
    layer7_outputs(786) <= a or b;
    layer7_outputs(787) <= a and b;
    layer7_outputs(788) <= a;
    layer7_outputs(789) <= a and not b;
    layer7_outputs(790) <= b;
    layer7_outputs(791) <= b;
    layer7_outputs(792) <= b;
    layer7_outputs(793) <= a;
    layer7_outputs(794) <= not b;
    layer7_outputs(795) <= '0';
    layer7_outputs(796) <= not (a or b);
    layer7_outputs(797) <= a;
    layer7_outputs(798) <= a and not b;
    layer7_outputs(799) <= a or b;
    layer7_outputs(800) <= a;
    layer7_outputs(801) <= not a;
    layer7_outputs(802) <= not (a or b);
    layer7_outputs(803) <= not a;
    layer7_outputs(804) <= not a;
    layer7_outputs(805) <= a and b;
    layer7_outputs(806) <= b;
    layer7_outputs(807) <= a and b;
    layer7_outputs(808) <= not b;
    layer7_outputs(809) <= a or b;
    layer7_outputs(810) <= not b or a;
    layer7_outputs(811) <= not (a xor b);
    layer7_outputs(812) <= not b or a;
    layer7_outputs(813) <= not a;
    layer7_outputs(814) <= not (a xor b);
    layer7_outputs(815) <= a;
    layer7_outputs(816) <= not a;
    layer7_outputs(817) <= a and not b;
    layer7_outputs(818) <= b;
    layer7_outputs(819) <= b;
    layer7_outputs(820) <= b;
    layer7_outputs(821) <= not (a and b);
    layer7_outputs(822) <= a or b;
    layer7_outputs(823) <= not a;
    layer7_outputs(824) <= a;
    layer7_outputs(825) <= not a;
    layer7_outputs(826) <= not b;
    layer7_outputs(827) <= a xor b;
    layer7_outputs(828) <= b;
    layer7_outputs(829) <= a xor b;
    layer7_outputs(830) <= not a or b;
    layer7_outputs(831) <= not b;
    layer7_outputs(832) <= not (a xor b);
    layer7_outputs(833) <= a and b;
    layer7_outputs(834) <= b;
    layer7_outputs(835) <= a;
    layer7_outputs(836) <= a and b;
    layer7_outputs(837) <= a;
    layer7_outputs(838) <= not (a and b);
    layer7_outputs(839) <= not (a xor b);
    layer7_outputs(840) <= not (a xor b);
    layer7_outputs(841) <= not b;
    layer7_outputs(842) <= a and b;
    layer7_outputs(843) <= a and not b;
    layer7_outputs(844) <= a;
    layer7_outputs(845) <= not (a and b);
    layer7_outputs(846) <= b;
    layer7_outputs(847) <= a;
    layer7_outputs(848) <= not b or a;
    layer7_outputs(849) <= b and not a;
    layer7_outputs(850) <= not b;
    layer7_outputs(851) <= a xor b;
    layer7_outputs(852) <= not (a xor b);
    layer7_outputs(853) <= a;
    layer7_outputs(854) <= a xor b;
    layer7_outputs(855) <= not b or a;
    layer7_outputs(856) <= a;
    layer7_outputs(857) <= a xor b;
    layer7_outputs(858) <= not (a and b);
    layer7_outputs(859) <= b and not a;
    layer7_outputs(860) <= a and not b;
    layer7_outputs(861) <= not b or a;
    layer7_outputs(862) <= a xor b;
    layer7_outputs(863) <= a or b;
    layer7_outputs(864) <= not b;
    layer7_outputs(865) <= not a;
    layer7_outputs(866) <= a and not b;
    layer7_outputs(867) <= a;
    layer7_outputs(868) <= a or b;
    layer7_outputs(869) <= not b or a;
    layer7_outputs(870) <= a and not b;
    layer7_outputs(871) <= not b;
    layer7_outputs(872) <= not a;
    layer7_outputs(873) <= a;
    layer7_outputs(874) <= not (a and b);
    layer7_outputs(875) <= b;
    layer7_outputs(876) <= '1';
    layer7_outputs(877) <= not (a or b);
    layer7_outputs(878) <= a;
    layer7_outputs(879) <= a;
    layer7_outputs(880) <= a and b;
    layer7_outputs(881) <= not b;
    layer7_outputs(882) <= not b or a;
    layer7_outputs(883) <= a;
    layer7_outputs(884) <= not a;
    layer7_outputs(885) <= not (a xor b);
    layer7_outputs(886) <= not a;
    layer7_outputs(887) <= a and not b;
    layer7_outputs(888) <= not b;
    layer7_outputs(889) <= a or b;
    layer7_outputs(890) <= a xor b;
    layer7_outputs(891) <= b;
    layer7_outputs(892) <= not b;
    layer7_outputs(893) <= b;
    layer7_outputs(894) <= not a or b;
    layer7_outputs(895) <= not b;
    layer7_outputs(896) <= a and b;
    layer7_outputs(897) <= a or b;
    layer7_outputs(898) <= a and b;
    layer7_outputs(899) <= not b;
    layer7_outputs(900) <= a;
    layer7_outputs(901) <= not b;
    layer7_outputs(902) <= a;
    layer7_outputs(903) <= a and not b;
    layer7_outputs(904) <= a and b;
    layer7_outputs(905) <= not (a xor b);
    layer7_outputs(906) <= a and not b;
    layer7_outputs(907) <= not (a or b);
    layer7_outputs(908) <= not (a xor b);
    layer7_outputs(909) <= a xor b;
    layer7_outputs(910) <= '0';
    layer7_outputs(911) <= a and not b;
    layer7_outputs(912) <= not a or b;
    layer7_outputs(913) <= '0';
    layer7_outputs(914) <= a;
    layer7_outputs(915) <= not a;
    layer7_outputs(916) <= a and not b;
    layer7_outputs(917) <= a;
    layer7_outputs(918) <= a and b;
    layer7_outputs(919) <= not (a or b);
    layer7_outputs(920) <= not b or a;
    layer7_outputs(921) <= not b;
    layer7_outputs(922) <= a xor b;
    layer7_outputs(923) <= b;
    layer7_outputs(924) <= not b;
    layer7_outputs(925) <= b;
    layer7_outputs(926) <= not (a xor b);
    layer7_outputs(927) <= b;
    layer7_outputs(928) <= not (a or b);
    layer7_outputs(929) <= not b;
    layer7_outputs(930) <= not a;
    layer7_outputs(931) <= not b or a;
    layer7_outputs(932) <= b and not a;
    layer7_outputs(933) <= not (a or b);
    layer7_outputs(934) <= not b;
    layer7_outputs(935) <= not (a xor b);
    layer7_outputs(936) <= a or b;
    layer7_outputs(937) <= a xor b;
    layer7_outputs(938) <= a xor b;
    layer7_outputs(939) <= a or b;
    layer7_outputs(940) <= not b;
    layer7_outputs(941) <= not a;
    layer7_outputs(942) <= b;
    layer7_outputs(943) <= not (a and b);
    layer7_outputs(944) <= a xor b;
    layer7_outputs(945) <= a and b;
    layer7_outputs(946) <= a and b;
    layer7_outputs(947) <= b;
    layer7_outputs(948) <= b and not a;
    layer7_outputs(949) <= not a;
    layer7_outputs(950) <= not a;
    layer7_outputs(951) <= b and not a;
    layer7_outputs(952) <= a and not b;
    layer7_outputs(953) <= not (a xor b);
    layer7_outputs(954) <= b;
    layer7_outputs(955) <= a and not b;
    layer7_outputs(956) <= not b or a;
    layer7_outputs(957) <= not (a and b);
    layer7_outputs(958) <= not a;
    layer7_outputs(959) <= '1';
    layer7_outputs(960) <= a and b;
    layer7_outputs(961) <= a and b;
    layer7_outputs(962) <= a;
    layer7_outputs(963) <= b and not a;
    layer7_outputs(964) <= a;
    layer7_outputs(965) <= a;
    layer7_outputs(966) <= not b;
    layer7_outputs(967) <= a;
    layer7_outputs(968) <= not a;
    layer7_outputs(969) <= b;
    layer7_outputs(970) <= a;
    layer7_outputs(971) <= not (a and b);
    layer7_outputs(972) <= not (a xor b);
    layer7_outputs(973) <= a xor b;
    layer7_outputs(974) <= not a;
    layer7_outputs(975) <= not b;
    layer7_outputs(976) <= a or b;
    layer7_outputs(977) <= not b;
    layer7_outputs(978) <= not b;
    layer7_outputs(979) <= not b;
    layer7_outputs(980) <= not a;
    layer7_outputs(981) <= not (a xor b);
    layer7_outputs(982) <= a xor b;
    layer7_outputs(983) <= a;
    layer7_outputs(984) <= not b;
    layer7_outputs(985) <= not b;
    layer7_outputs(986) <= a and not b;
    layer7_outputs(987) <= not (a xor b);
    layer7_outputs(988) <= not b;
    layer7_outputs(989) <= b;
    layer7_outputs(990) <= not a;
    layer7_outputs(991) <= b;
    layer7_outputs(992) <= a;
    layer7_outputs(993) <= a;
    layer7_outputs(994) <= not (a or b);
    layer7_outputs(995) <= not b or a;
    layer7_outputs(996) <= not b;
    layer7_outputs(997) <= not (a or b);
    layer7_outputs(998) <= not b;
    layer7_outputs(999) <= not (a or b);
    layer7_outputs(1000) <= a;
    layer7_outputs(1001) <= not b;
    layer7_outputs(1002) <= not (a or b);
    layer7_outputs(1003) <= a and not b;
    layer7_outputs(1004) <= not a;
    layer7_outputs(1005) <= not b;
    layer7_outputs(1006) <= not b or a;
    layer7_outputs(1007) <= not a;
    layer7_outputs(1008) <= not b;
    layer7_outputs(1009) <= not a or b;
    layer7_outputs(1010) <= b;
    layer7_outputs(1011) <= b and not a;
    layer7_outputs(1012) <= a;
    layer7_outputs(1013) <= a and b;
    layer7_outputs(1014) <= not (a xor b);
    layer7_outputs(1015) <= not (a and b);
    layer7_outputs(1016) <= not a;
    layer7_outputs(1017) <= not a;
    layer7_outputs(1018) <= b and not a;
    layer7_outputs(1019) <= a;
    layer7_outputs(1020) <= not b;
    layer7_outputs(1021) <= not b;
    layer7_outputs(1022) <= a xor b;
    layer7_outputs(1023) <= b;
    layer7_outputs(1024) <= a or b;
    layer7_outputs(1025) <= a;
    layer7_outputs(1026) <= b;
    layer7_outputs(1027) <= not b;
    layer7_outputs(1028) <= b;
    layer7_outputs(1029) <= not (a xor b);
    layer7_outputs(1030) <= a;
    layer7_outputs(1031) <= not (a xor b);
    layer7_outputs(1032) <= a and not b;
    layer7_outputs(1033) <= b;
    layer7_outputs(1034) <= a;
    layer7_outputs(1035) <= not (a xor b);
    layer7_outputs(1036) <= a xor b;
    layer7_outputs(1037) <= not a or b;
    layer7_outputs(1038) <= '1';
    layer7_outputs(1039) <= not b;
    layer7_outputs(1040) <= not a;
    layer7_outputs(1041) <= not b;
    layer7_outputs(1042) <= not (a or b);
    layer7_outputs(1043) <= b;
    layer7_outputs(1044) <= a and not b;
    layer7_outputs(1045) <= b;
    layer7_outputs(1046) <= not (a and b);
    layer7_outputs(1047) <= not (a or b);
    layer7_outputs(1048) <= b;
    layer7_outputs(1049) <= not a;
    layer7_outputs(1050) <= not a;
    layer7_outputs(1051) <= not a;
    layer7_outputs(1052) <= '1';
    layer7_outputs(1053) <= not b or a;
    layer7_outputs(1054) <= not (a and b);
    layer7_outputs(1055) <= b;
    layer7_outputs(1056) <= not b;
    layer7_outputs(1057) <= a or b;
    layer7_outputs(1058) <= a;
    layer7_outputs(1059) <= b and not a;
    layer7_outputs(1060) <= b and not a;
    layer7_outputs(1061) <= not (a and b);
    layer7_outputs(1062) <= b;
    layer7_outputs(1063) <= b;
    layer7_outputs(1064) <= a and not b;
    layer7_outputs(1065) <= not a or b;
    layer7_outputs(1066) <= '1';
    layer7_outputs(1067) <= a;
    layer7_outputs(1068) <= a;
    layer7_outputs(1069) <= a xor b;
    layer7_outputs(1070) <= not b;
    layer7_outputs(1071) <= not (a xor b);
    layer7_outputs(1072) <= a xor b;
    layer7_outputs(1073) <= '1';
    layer7_outputs(1074) <= b;
    layer7_outputs(1075) <= not (a and b);
    layer7_outputs(1076) <= a;
    layer7_outputs(1077) <= not (a or b);
    layer7_outputs(1078) <= b;
    layer7_outputs(1079) <= not b;
    layer7_outputs(1080) <= not b;
    layer7_outputs(1081) <= not a or b;
    layer7_outputs(1082) <= a or b;
    layer7_outputs(1083) <= b;
    layer7_outputs(1084) <= a xor b;
    layer7_outputs(1085) <= '0';
    layer7_outputs(1086) <= b and not a;
    layer7_outputs(1087) <= '1';
    layer7_outputs(1088) <= b;
    layer7_outputs(1089) <= not b;
    layer7_outputs(1090) <= b;
    layer7_outputs(1091) <= a;
    layer7_outputs(1092) <= a;
    layer7_outputs(1093) <= a xor b;
    layer7_outputs(1094) <= not a;
    layer7_outputs(1095) <= a xor b;
    layer7_outputs(1096) <= not a;
    layer7_outputs(1097) <= a;
    layer7_outputs(1098) <= not (a and b);
    layer7_outputs(1099) <= a xor b;
    layer7_outputs(1100) <= not (a xor b);
    layer7_outputs(1101) <= a and not b;
    layer7_outputs(1102) <= a and b;
    layer7_outputs(1103) <= b and not a;
    layer7_outputs(1104) <= b and not a;
    layer7_outputs(1105) <= not b;
    layer7_outputs(1106) <= not (a and b);
    layer7_outputs(1107) <= a;
    layer7_outputs(1108) <= a and b;
    layer7_outputs(1109) <= '1';
    layer7_outputs(1110) <= a;
    layer7_outputs(1111) <= a or b;
    layer7_outputs(1112) <= a;
    layer7_outputs(1113) <= b and not a;
    layer7_outputs(1114) <= a;
    layer7_outputs(1115) <= b;
    layer7_outputs(1116) <= not a;
    layer7_outputs(1117) <= not b;
    layer7_outputs(1118) <= a;
    layer7_outputs(1119) <= not b;
    layer7_outputs(1120) <= b;
    layer7_outputs(1121) <= not a;
    layer7_outputs(1122) <= b;
    layer7_outputs(1123) <= not a;
    layer7_outputs(1124) <= b and not a;
    layer7_outputs(1125) <= b;
    layer7_outputs(1126) <= a xor b;
    layer7_outputs(1127) <= not a or b;
    layer7_outputs(1128) <= a and b;
    layer7_outputs(1129) <= a;
    layer7_outputs(1130) <= not a;
    layer7_outputs(1131) <= not (a or b);
    layer7_outputs(1132) <= not a;
    layer7_outputs(1133) <= not (a or b);
    layer7_outputs(1134) <= a xor b;
    layer7_outputs(1135) <= b;
    layer7_outputs(1136) <= not (a xor b);
    layer7_outputs(1137) <= a and not b;
    layer7_outputs(1138) <= a;
    layer7_outputs(1139) <= a and b;
    layer7_outputs(1140) <= a;
    layer7_outputs(1141) <= a;
    layer7_outputs(1142) <= a;
    layer7_outputs(1143) <= not (a and b);
    layer7_outputs(1144) <= not b;
    layer7_outputs(1145) <= not (a xor b);
    layer7_outputs(1146) <= a and b;
    layer7_outputs(1147) <= not a or b;
    layer7_outputs(1148) <= not (a and b);
    layer7_outputs(1149) <= not (a or b);
    layer7_outputs(1150) <= b;
    layer7_outputs(1151) <= a and b;
    layer7_outputs(1152) <= a xor b;
    layer7_outputs(1153) <= not (a xor b);
    layer7_outputs(1154) <= a xor b;
    layer7_outputs(1155) <= a and not b;
    layer7_outputs(1156) <= a xor b;
    layer7_outputs(1157) <= not a;
    layer7_outputs(1158) <= a xor b;
    layer7_outputs(1159) <= b;
    layer7_outputs(1160) <= b;
    layer7_outputs(1161) <= a and not b;
    layer7_outputs(1162) <= not a or b;
    layer7_outputs(1163) <= not a;
    layer7_outputs(1164) <= a and b;
    layer7_outputs(1165) <= not (a and b);
    layer7_outputs(1166) <= not a;
    layer7_outputs(1167) <= not (a or b);
    layer7_outputs(1168) <= a;
    layer7_outputs(1169) <= not (a xor b);
    layer7_outputs(1170) <= not b or a;
    layer7_outputs(1171) <= not b;
    layer7_outputs(1172) <= not b;
    layer7_outputs(1173) <= a or b;
    layer7_outputs(1174) <= not a;
    layer7_outputs(1175) <= not (a xor b);
    layer7_outputs(1176) <= not a;
    layer7_outputs(1177) <= not b or a;
    layer7_outputs(1178) <= not a or b;
    layer7_outputs(1179) <= not b;
    layer7_outputs(1180) <= not (a or b);
    layer7_outputs(1181) <= a;
    layer7_outputs(1182) <= a;
    layer7_outputs(1183) <= not b or a;
    layer7_outputs(1184) <= not b;
    layer7_outputs(1185) <= not (a xor b);
    layer7_outputs(1186) <= not a;
    layer7_outputs(1187) <= not a or b;
    layer7_outputs(1188) <= a or b;
    layer7_outputs(1189) <= not b;
    layer7_outputs(1190) <= not (a or b);
    layer7_outputs(1191) <= a;
    layer7_outputs(1192) <= not b;
    layer7_outputs(1193) <= not b or a;
    layer7_outputs(1194) <= not a or b;
    layer7_outputs(1195) <= not (a xor b);
    layer7_outputs(1196) <= not a;
    layer7_outputs(1197) <= a xor b;
    layer7_outputs(1198) <= not b;
    layer7_outputs(1199) <= a and b;
    layer7_outputs(1200) <= a;
    layer7_outputs(1201) <= a xor b;
    layer7_outputs(1202) <= b;
    layer7_outputs(1203) <= a;
    layer7_outputs(1204) <= a and not b;
    layer7_outputs(1205) <= not (a or b);
    layer7_outputs(1206) <= not b;
    layer7_outputs(1207) <= not (a xor b);
    layer7_outputs(1208) <= not a;
    layer7_outputs(1209) <= b;
    layer7_outputs(1210) <= not (a or b);
    layer7_outputs(1211) <= a xor b;
    layer7_outputs(1212) <= not b or a;
    layer7_outputs(1213) <= not a;
    layer7_outputs(1214) <= not b or a;
    layer7_outputs(1215) <= not b;
    layer7_outputs(1216) <= b;
    layer7_outputs(1217) <= not b or a;
    layer7_outputs(1218) <= b;
    layer7_outputs(1219) <= not a;
    layer7_outputs(1220) <= b and not a;
    layer7_outputs(1221) <= a or b;
    layer7_outputs(1222) <= b and not a;
    layer7_outputs(1223) <= a xor b;
    layer7_outputs(1224) <= a;
    layer7_outputs(1225) <= not a;
    layer7_outputs(1226) <= a xor b;
    layer7_outputs(1227) <= not a;
    layer7_outputs(1228) <= b;
    layer7_outputs(1229) <= not b;
    layer7_outputs(1230) <= not b;
    layer7_outputs(1231) <= not b;
    layer7_outputs(1232) <= not b;
    layer7_outputs(1233) <= not (a and b);
    layer7_outputs(1234) <= b and not a;
    layer7_outputs(1235) <= not (a or b);
    layer7_outputs(1236) <= not a;
    layer7_outputs(1237) <= not (a xor b);
    layer7_outputs(1238) <= a;
    layer7_outputs(1239) <= a or b;
    layer7_outputs(1240) <= not (a or b);
    layer7_outputs(1241) <= not (a and b);
    layer7_outputs(1242) <= b and not a;
    layer7_outputs(1243) <= b;
    layer7_outputs(1244) <= not b;
    layer7_outputs(1245) <= not b;
    layer7_outputs(1246) <= a or b;
    layer7_outputs(1247) <= not b;
    layer7_outputs(1248) <= a xor b;
    layer7_outputs(1249) <= not b;
    layer7_outputs(1250) <= not b or a;
    layer7_outputs(1251) <= not (a and b);
    layer7_outputs(1252) <= not b;
    layer7_outputs(1253) <= not a;
    layer7_outputs(1254) <= a;
    layer7_outputs(1255) <= a and b;
    layer7_outputs(1256) <= a and not b;
    layer7_outputs(1257) <= a or b;
    layer7_outputs(1258) <= not a;
    layer7_outputs(1259) <= a and not b;
    layer7_outputs(1260) <= not b;
    layer7_outputs(1261) <= a xor b;
    layer7_outputs(1262) <= b;
    layer7_outputs(1263) <= b;
    layer7_outputs(1264) <= b;
    layer7_outputs(1265) <= not b;
    layer7_outputs(1266) <= b;
    layer7_outputs(1267) <= b;
    layer7_outputs(1268) <= not (a or b);
    layer7_outputs(1269) <= not b or a;
    layer7_outputs(1270) <= '0';
    layer7_outputs(1271) <= a;
    layer7_outputs(1272) <= a and not b;
    layer7_outputs(1273) <= b;
    layer7_outputs(1274) <= not b or a;
    layer7_outputs(1275) <= not (a and b);
    layer7_outputs(1276) <= not b;
    layer7_outputs(1277) <= b;
    layer7_outputs(1278) <= not b;
    layer7_outputs(1279) <= not (a xor b);
    layer7_outputs(1280) <= not a;
    layer7_outputs(1281) <= not b;
    layer7_outputs(1282) <= not (a xor b);
    layer7_outputs(1283) <= not a or b;
    layer7_outputs(1284) <= a or b;
    layer7_outputs(1285) <= not (a and b);
    layer7_outputs(1286) <= not a or b;
    layer7_outputs(1287) <= not a or b;
    layer7_outputs(1288) <= a and not b;
    layer7_outputs(1289) <= a xor b;
    layer7_outputs(1290) <= a;
    layer7_outputs(1291) <= a;
    layer7_outputs(1292) <= not a;
    layer7_outputs(1293) <= not b;
    layer7_outputs(1294) <= not a;
    layer7_outputs(1295) <= not a;
    layer7_outputs(1296) <= a;
    layer7_outputs(1297) <= a and b;
    layer7_outputs(1298) <= not b;
    layer7_outputs(1299) <= not b;
    layer7_outputs(1300) <= not (a or b);
    layer7_outputs(1301) <= b;
    layer7_outputs(1302) <= a xor b;
    layer7_outputs(1303) <= a;
    layer7_outputs(1304) <= not (a xor b);
    layer7_outputs(1305) <= not b or a;
    layer7_outputs(1306) <= not (a xor b);
    layer7_outputs(1307) <= not b;
    layer7_outputs(1308) <= a;
    layer7_outputs(1309) <= a and not b;
    layer7_outputs(1310) <= not b or a;
    layer7_outputs(1311) <= b;
    layer7_outputs(1312) <= a;
    layer7_outputs(1313) <= not (a and b);
    layer7_outputs(1314) <= not (a xor b);
    layer7_outputs(1315) <= not b or a;
    layer7_outputs(1316) <= not a;
    layer7_outputs(1317) <= a or b;
    layer7_outputs(1318) <= not (a or b);
    layer7_outputs(1319) <= a;
    layer7_outputs(1320) <= not a or b;
    layer7_outputs(1321) <= not a;
    layer7_outputs(1322) <= a xor b;
    layer7_outputs(1323) <= a and not b;
    layer7_outputs(1324) <= not (a and b);
    layer7_outputs(1325) <= not (a or b);
    layer7_outputs(1326) <= b;
    layer7_outputs(1327) <= not b or a;
    layer7_outputs(1328) <= not (a or b);
    layer7_outputs(1329) <= not (a and b);
    layer7_outputs(1330) <= a and b;
    layer7_outputs(1331) <= b and not a;
    layer7_outputs(1332) <= a and b;
    layer7_outputs(1333) <= not a;
    layer7_outputs(1334) <= a xor b;
    layer7_outputs(1335) <= a;
    layer7_outputs(1336) <= a xor b;
    layer7_outputs(1337) <= not (a xor b);
    layer7_outputs(1338) <= not a;
    layer7_outputs(1339) <= not a;
    layer7_outputs(1340) <= not a;
    layer7_outputs(1341) <= a;
    layer7_outputs(1342) <= b;
    layer7_outputs(1343) <= b;
    layer7_outputs(1344) <= not (a or b);
    layer7_outputs(1345) <= not b or a;
    layer7_outputs(1346) <= not b;
    layer7_outputs(1347) <= not a;
    layer7_outputs(1348) <= a or b;
    layer7_outputs(1349) <= b;
    layer7_outputs(1350) <= not b;
    layer7_outputs(1351) <= not b;
    layer7_outputs(1352) <= not a;
    layer7_outputs(1353) <= a;
    layer7_outputs(1354) <= not a or b;
    layer7_outputs(1355) <= not (a xor b);
    layer7_outputs(1356) <= not a;
    layer7_outputs(1357) <= a and not b;
    layer7_outputs(1358) <= not b or a;
    layer7_outputs(1359) <= a;
    layer7_outputs(1360) <= not (a xor b);
    layer7_outputs(1361) <= a or b;
    layer7_outputs(1362) <= b;
    layer7_outputs(1363) <= not b;
    layer7_outputs(1364) <= b and not a;
    layer7_outputs(1365) <= a and not b;
    layer7_outputs(1366) <= not (a and b);
    layer7_outputs(1367) <= not b or a;
    layer7_outputs(1368) <= not (a or b);
    layer7_outputs(1369) <= a;
    layer7_outputs(1370) <= b;
    layer7_outputs(1371) <= b;
    layer7_outputs(1372) <= a or b;
    layer7_outputs(1373) <= a xor b;
    layer7_outputs(1374) <= not a;
    layer7_outputs(1375) <= a and b;
    layer7_outputs(1376) <= b;
    layer7_outputs(1377) <= not b or a;
    layer7_outputs(1378) <= not b;
    layer7_outputs(1379) <= b and not a;
    layer7_outputs(1380) <= a and not b;
    layer7_outputs(1381) <= not (a and b);
    layer7_outputs(1382) <= a xor b;
    layer7_outputs(1383) <= a;
    layer7_outputs(1384) <= not b or a;
    layer7_outputs(1385) <= a or b;
    layer7_outputs(1386) <= not b or a;
    layer7_outputs(1387) <= b and not a;
    layer7_outputs(1388) <= not b or a;
    layer7_outputs(1389) <= b;
    layer7_outputs(1390) <= a;
    layer7_outputs(1391) <= not (a xor b);
    layer7_outputs(1392) <= not b;
    layer7_outputs(1393) <= b;
    layer7_outputs(1394) <= a;
    layer7_outputs(1395) <= a and b;
    layer7_outputs(1396) <= a or b;
    layer7_outputs(1397) <= not (a and b);
    layer7_outputs(1398) <= a and not b;
    layer7_outputs(1399) <= not (a xor b);
    layer7_outputs(1400) <= b;
    layer7_outputs(1401) <= not b;
    layer7_outputs(1402) <= not (a xor b);
    layer7_outputs(1403) <= not (a and b);
    layer7_outputs(1404) <= not (a or b);
    layer7_outputs(1405) <= a xor b;
    layer7_outputs(1406) <= b and not a;
    layer7_outputs(1407) <= a;
    layer7_outputs(1408) <= a;
    layer7_outputs(1409) <= not b or a;
    layer7_outputs(1410) <= not a or b;
    layer7_outputs(1411) <= not (a and b);
    layer7_outputs(1412) <= not b;
    layer7_outputs(1413) <= b and not a;
    layer7_outputs(1414) <= a;
    layer7_outputs(1415) <= not (a xor b);
    layer7_outputs(1416) <= not (a xor b);
    layer7_outputs(1417) <= a xor b;
    layer7_outputs(1418) <= a;
    layer7_outputs(1419) <= a or b;
    layer7_outputs(1420) <= not (a xor b);
    layer7_outputs(1421) <= not (a and b);
    layer7_outputs(1422) <= not (a xor b);
    layer7_outputs(1423) <= not a or b;
    layer7_outputs(1424) <= not (a or b);
    layer7_outputs(1425) <= '0';
    layer7_outputs(1426) <= not b;
    layer7_outputs(1427) <= not a;
    layer7_outputs(1428) <= a xor b;
    layer7_outputs(1429) <= a xor b;
    layer7_outputs(1430) <= b and not a;
    layer7_outputs(1431) <= not b;
    layer7_outputs(1432) <= a xor b;
    layer7_outputs(1433) <= a and b;
    layer7_outputs(1434) <= not (a xor b);
    layer7_outputs(1435) <= b;
    layer7_outputs(1436) <= not a;
    layer7_outputs(1437) <= not b;
    layer7_outputs(1438) <= a;
    layer7_outputs(1439) <= a;
    layer7_outputs(1440) <= b and not a;
    layer7_outputs(1441) <= not a;
    layer7_outputs(1442) <= not b;
    layer7_outputs(1443) <= not (a xor b);
    layer7_outputs(1444) <= a and not b;
    layer7_outputs(1445) <= not a;
    layer7_outputs(1446) <= '0';
    layer7_outputs(1447) <= a xor b;
    layer7_outputs(1448) <= a;
    layer7_outputs(1449) <= not a;
    layer7_outputs(1450) <= not b;
    layer7_outputs(1451) <= a;
    layer7_outputs(1452) <= a xor b;
    layer7_outputs(1453) <= not a;
    layer7_outputs(1454) <= a and not b;
    layer7_outputs(1455) <= not b;
    layer7_outputs(1456) <= not a;
    layer7_outputs(1457) <= a xor b;
    layer7_outputs(1458) <= b;
    layer7_outputs(1459) <= a and b;
    layer7_outputs(1460) <= b;
    layer7_outputs(1461) <= b and not a;
    layer7_outputs(1462) <= not a;
    layer7_outputs(1463) <= not a;
    layer7_outputs(1464) <= a xor b;
    layer7_outputs(1465) <= b;
    layer7_outputs(1466) <= a or b;
    layer7_outputs(1467) <= b;
    layer7_outputs(1468) <= a;
    layer7_outputs(1469) <= not b;
    layer7_outputs(1470) <= not b or a;
    layer7_outputs(1471) <= not b;
    layer7_outputs(1472) <= not (a xor b);
    layer7_outputs(1473) <= not b;
    layer7_outputs(1474) <= b and not a;
    layer7_outputs(1475) <= not b;
    layer7_outputs(1476) <= not b;
    layer7_outputs(1477) <= not (a and b);
    layer7_outputs(1478) <= b;
    layer7_outputs(1479) <= not b or a;
    layer7_outputs(1480) <= not (a xor b);
    layer7_outputs(1481) <= not (a xor b);
    layer7_outputs(1482) <= not b;
    layer7_outputs(1483) <= not (a xor b);
    layer7_outputs(1484) <= a xor b;
    layer7_outputs(1485) <= not b or a;
    layer7_outputs(1486) <= a or b;
    layer7_outputs(1487) <= b;
    layer7_outputs(1488) <= not b;
    layer7_outputs(1489) <= a xor b;
    layer7_outputs(1490) <= not b;
    layer7_outputs(1491) <= a;
    layer7_outputs(1492) <= not b;
    layer7_outputs(1493) <= b;
    layer7_outputs(1494) <= not a;
    layer7_outputs(1495) <= a or b;
    layer7_outputs(1496) <= a;
    layer7_outputs(1497) <= not (a xor b);
    layer7_outputs(1498) <= not (a or b);
    layer7_outputs(1499) <= b;
    layer7_outputs(1500) <= not (a and b);
    layer7_outputs(1501) <= b;
    layer7_outputs(1502) <= b;
    layer7_outputs(1503) <= b;
    layer7_outputs(1504) <= not a or b;
    layer7_outputs(1505) <= b;
    layer7_outputs(1506) <= a xor b;
    layer7_outputs(1507) <= b;
    layer7_outputs(1508) <= not (a xor b);
    layer7_outputs(1509) <= not b;
    layer7_outputs(1510) <= not b;
    layer7_outputs(1511) <= b;
    layer7_outputs(1512) <= a or b;
    layer7_outputs(1513) <= not b;
    layer7_outputs(1514) <= not a;
    layer7_outputs(1515) <= not (a and b);
    layer7_outputs(1516) <= a;
    layer7_outputs(1517) <= a xor b;
    layer7_outputs(1518) <= a;
    layer7_outputs(1519) <= not (a or b);
    layer7_outputs(1520) <= a xor b;
    layer7_outputs(1521) <= not a or b;
    layer7_outputs(1522) <= a;
    layer7_outputs(1523) <= a xor b;
    layer7_outputs(1524) <= a;
    layer7_outputs(1525) <= not (a and b);
    layer7_outputs(1526) <= not (a xor b);
    layer7_outputs(1527) <= a;
    layer7_outputs(1528) <= not b;
    layer7_outputs(1529) <= not (a xor b);
    layer7_outputs(1530) <= a;
    layer7_outputs(1531) <= not (a xor b);
    layer7_outputs(1532) <= not (a xor b);
    layer7_outputs(1533) <= b;
    layer7_outputs(1534) <= not (a and b);
    layer7_outputs(1535) <= not b;
    layer7_outputs(1536) <= not (a xor b);
    layer7_outputs(1537) <= not b or a;
    layer7_outputs(1538) <= b;
    layer7_outputs(1539) <= not b;
    layer7_outputs(1540) <= a and not b;
    layer7_outputs(1541) <= a or b;
    layer7_outputs(1542) <= not a;
    layer7_outputs(1543) <= not b;
    layer7_outputs(1544) <= a and b;
    layer7_outputs(1545) <= not b or a;
    layer7_outputs(1546) <= a xor b;
    layer7_outputs(1547) <= a xor b;
    layer7_outputs(1548) <= not b;
    layer7_outputs(1549) <= not b or a;
    layer7_outputs(1550) <= b;
    layer7_outputs(1551) <= a;
    layer7_outputs(1552) <= b;
    layer7_outputs(1553) <= a and not b;
    layer7_outputs(1554) <= b;
    layer7_outputs(1555) <= not a;
    layer7_outputs(1556) <= not (a or b);
    layer7_outputs(1557) <= b and not a;
    layer7_outputs(1558) <= not (a and b);
    layer7_outputs(1559) <= not (a xor b);
    layer7_outputs(1560) <= not (a xor b);
    layer7_outputs(1561) <= not b;
    layer7_outputs(1562) <= not a;
    layer7_outputs(1563) <= a xor b;
    layer7_outputs(1564) <= not a;
    layer7_outputs(1565) <= not b;
    layer7_outputs(1566) <= a;
    layer7_outputs(1567) <= b;
    layer7_outputs(1568) <= not b or a;
    layer7_outputs(1569) <= not b or a;
    layer7_outputs(1570) <= a;
    layer7_outputs(1571) <= not b or a;
    layer7_outputs(1572) <= not b or a;
    layer7_outputs(1573) <= a or b;
    layer7_outputs(1574) <= not b;
    layer7_outputs(1575) <= a;
    layer7_outputs(1576) <= a and not b;
    layer7_outputs(1577) <= a;
    layer7_outputs(1578) <= not a or b;
    layer7_outputs(1579) <= b;
    layer7_outputs(1580) <= b;
    layer7_outputs(1581) <= b;
    layer7_outputs(1582) <= a;
    layer7_outputs(1583) <= not b;
    layer7_outputs(1584) <= a;
    layer7_outputs(1585) <= not b;
    layer7_outputs(1586) <= a xor b;
    layer7_outputs(1587) <= '1';
    layer7_outputs(1588) <= not b;
    layer7_outputs(1589) <= b and not a;
    layer7_outputs(1590) <= not (a xor b);
    layer7_outputs(1591) <= a;
    layer7_outputs(1592) <= b;
    layer7_outputs(1593) <= not (a and b);
    layer7_outputs(1594) <= b;
    layer7_outputs(1595) <= not b;
    layer7_outputs(1596) <= a and not b;
    layer7_outputs(1597) <= a and b;
    layer7_outputs(1598) <= not (a xor b);
    layer7_outputs(1599) <= not b;
    layer7_outputs(1600) <= not b or a;
    layer7_outputs(1601) <= not (a and b);
    layer7_outputs(1602) <= not (a and b);
    layer7_outputs(1603) <= b;
    layer7_outputs(1604) <= a;
    layer7_outputs(1605) <= not (a xor b);
    layer7_outputs(1606) <= not (a and b);
    layer7_outputs(1607) <= b;
    layer7_outputs(1608) <= not a;
    layer7_outputs(1609) <= b;
    layer7_outputs(1610) <= not b or a;
    layer7_outputs(1611) <= b;
    layer7_outputs(1612) <= not a;
    layer7_outputs(1613) <= a;
    layer7_outputs(1614) <= a and b;
    layer7_outputs(1615) <= b;
    layer7_outputs(1616) <= a;
    layer7_outputs(1617) <= '1';
    layer7_outputs(1618) <= not a or b;
    layer7_outputs(1619) <= a xor b;
    layer7_outputs(1620) <= not a;
    layer7_outputs(1621) <= not (a xor b);
    layer7_outputs(1622) <= not b or a;
    layer7_outputs(1623) <= not a;
    layer7_outputs(1624) <= b and not a;
    layer7_outputs(1625) <= not b;
    layer7_outputs(1626) <= not (a xor b);
    layer7_outputs(1627) <= not (a xor b);
    layer7_outputs(1628) <= a;
    layer7_outputs(1629) <= not b;
    layer7_outputs(1630) <= not b;
    layer7_outputs(1631) <= not b;
    layer7_outputs(1632) <= not a or b;
    layer7_outputs(1633) <= a and b;
    layer7_outputs(1634) <= a or b;
    layer7_outputs(1635) <= b;
    layer7_outputs(1636) <= not a;
    layer7_outputs(1637) <= not a;
    layer7_outputs(1638) <= a;
    layer7_outputs(1639) <= b and not a;
    layer7_outputs(1640) <= not (a or b);
    layer7_outputs(1641) <= not b;
    layer7_outputs(1642) <= not b;
    layer7_outputs(1643) <= b;
    layer7_outputs(1644) <= a and b;
    layer7_outputs(1645) <= not (a xor b);
    layer7_outputs(1646) <= not (a and b);
    layer7_outputs(1647) <= not a;
    layer7_outputs(1648) <= not (a xor b);
    layer7_outputs(1649) <= not b or a;
    layer7_outputs(1650) <= not b;
    layer7_outputs(1651) <= a;
    layer7_outputs(1652) <= b;
    layer7_outputs(1653) <= not a;
    layer7_outputs(1654) <= b;
    layer7_outputs(1655) <= not a;
    layer7_outputs(1656) <= a xor b;
    layer7_outputs(1657) <= a and not b;
    layer7_outputs(1658) <= '1';
    layer7_outputs(1659) <= a;
    layer7_outputs(1660) <= not (a or b);
    layer7_outputs(1661) <= not (a xor b);
    layer7_outputs(1662) <= not (a xor b);
    layer7_outputs(1663) <= a;
    layer7_outputs(1664) <= a or b;
    layer7_outputs(1665) <= a or b;
    layer7_outputs(1666) <= not (a and b);
    layer7_outputs(1667) <= not b;
    layer7_outputs(1668) <= not (a or b);
    layer7_outputs(1669) <= a and b;
    layer7_outputs(1670) <= not (a xor b);
    layer7_outputs(1671) <= not (a xor b);
    layer7_outputs(1672) <= a xor b;
    layer7_outputs(1673) <= not b;
    layer7_outputs(1674) <= b;
    layer7_outputs(1675) <= not a;
    layer7_outputs(1676) <= not (a xor b);
    layer7_outputs(1677) <= not a;
    layer7_outputs(1678) <= a and not b;
    layer7_outputs(1679) <= not (a xor b);
    layer7_outputs(1680) <= not a;
    layer7_outputs(1681) <= not b or a;
    layer7_outputs(1682) <= not (a or b);
    layer7_outputs(1683) <= b;
    layer7_outputs(1684) <= not a or b;
    layer7_outputs(1685) <= b;
    layer7_outputs(1686) <= not (a or b);
    layer7_outputs(1687) <= not (a or b);
    layer7_outputs(1688) <= not (a or b);
    layer7_outputs(1689) <= a xor b;
    layer7_outputs(1690) <= not (a or b);
    layer7_outputs(1691) <= not a;
    layer7_outputs(1692) <= b;
    layer7_outputs(1693) <= a or b;
    layer7_outputs(1694) <= not a;
    layer7_outputs(1695) <= b;
    layer7_outputs(1696) <= not (a and b);
    layer7_outputs(1697) <= a;
    layer7_outputs(1698) <= a;
    layer7_outputs(1699) <= not b or a;
    layer7_outputs(1700) <= not b;
    layer7_outputs(1701) <= not b or a;
    layer7_outputs(1702) <= b and not a;
    layer7_outputs(1703) <= not a;
    layer7_outputs(1704) <= not a;
    layer7_outputs(1705) <= not b or a;
    layer7_outputs(1706) <= not a or b;
    layer7_outputs(1707) <= a and not b;
    layer7_outputs(1708) <= not a;
    layer7_outputs(1709) <= a;
    layer7_outputs(1710) <= not (a xor b);
    layer7_outputs(1711) <= b;
    layer7_outputs(1712) <= a or b;
    layer7_outputs(1713) <= not (a xor b);
    layer7_outputs(1714) <= a;
    layer7_outputs(1715) <= not a;
    layer7_outputs(1716) <= b;
    layer7_outputs(1717) <= not (a and b);
    layer7_outputs(1718) <= not a;
    layer7_outputs(1719) <= not a;
    layer7_outputs(1720) <= not b or a;
    layer7_outputs(1721) <= not (a xor b);
    layer7_outputs(1722) <= a;
    layer7_outputs(1723) <= not b or a;
    layer7_outputs(1724) <= a and b;
    layer7_outputs(1725) <= a xor b;
    layer7_outputs(1726) <= not a;
    layer7_outputs(1727) <= a;
    layer7_outputs(1728) <= a and b;
    layer7_outputs(1729) <= not a;
    layer7_outputs(1730) <= not a;
    layer7_outputs(1731) <= a;
    layer7_outputs(1732) <= not a or b;
    layer7_outputs(1733) <= a xor b;
    layer7_outputs(1734) <= not b;
    layer7_outputs(1735) <= b;
    layer7_outputs(1736) <= not (a or b);
    layer7_outputs(1737) <= not a or b;
    layer7_outputs(1738) <= a and b;
    layer7_outputs(1739) <= not a or b;
    layer7_outputs(1740) <= not a;
    layer7_outputs(1741) <= b and not a;
    layer7_outputs(1742) <= not (a xor b);
    layer7_outputs(1743) <= not b or a;
    layer7_outputs(1744) <= b;
    layer7_outputs(1745) <= not a;
    layer7_outputs(1746) <= a;
    layer7_outputs(1747) <= not b;
    layer7_outputs(1748) <= not b;
    layer7_outputs(1749) <= a or b;
    layer7_outputs(1750) <= a xor b;
    layer7_outputs(1751) <= a xor b;
    layer7_outputs(1752) <= not (a xor b);
    layer7_outputs(1753) <= a;
    layer7_outputs(1754) <= a and b;
    layer7_outputs(1755) <= a xor b;
    layer7_outputs(1756) <= b;
    layer7_outputs(1757) <= a xor b;
    layer7_outputs(1758) <= a;
    layer7_outputs(1759) <= not (a xor b);
    layer7_outputs(1760) <= not a;
    layer7_outputs(1761) <= b;
    layer7_outputs(1762) <= not (a or b);
    layer7_outputs(1763) <= not b;
    layer7_outputs(1764) <= not (a or b);
    layer7_outputs(1765) <= not a;
    layer7_outputs(1766) <= a and not b;
    layer7_outputs(1767) <= not b;
    layer7_outputs(1768) <= not (a xor b);
    layer7_outputs(1769) <= a or b;
    layer7_outputs(1770) <= not b;
    layer7_outputs(1771) <= b;
    layer7_outputs(1772) <= not b;
    layer7_outputs(1773) <= a and not b;
    layer7_outputs(1774) <= not a;
    layer7_outputs(1775) <= not (a xor b);
    layer7_outputs(1776) <= not b or a;
    layer7_outputs(1777) <= not a;
    layer7_outputs(1778) <= b;
    layer7_outputs(1779) <= not (a xor b);
    layer7_outputs(1780) <= b;
    layer7_outputs(1781) <= a or b;
    layer7_outputs(1782) <= b;
    layer7_outputs(1783) <= a xor b;
    layer7_outputs(1784) <= not a or b;
    layer7_outputs(1785) <= a and not b;
    layer7_outputs(1786) <= a;
    layer7_outputs(1787) <= a;
    layer7_outputs(1788) <= not b;
    layer7_outputs(1789) <= not (a xor b);
    layer7_outputs(1790) <= a xor b;
    layer7_outputs(1791) <= b;
    layer7_outputs(1792) <= b;
    layer7_outputs(1793) <= a and not b;
    layer7_outputs(1794) <= a xor b;
    layer7_outputs(1795) <= not a;
    layer7_outputs(1796) <= not (a and b);
    layer7_outputs(1797) <= not (a xor b);
    layer7_outputs(1798) <= not (a and b);
    layer7_outputs(1799) <= not (a xor b);
    layer7_outputs(1800) <= b;
    layer7_outputs(1801) <= b;
    layer7_outputs(1802) <= not b;
    layer7_outputs(1803) <= not (a or b);
    layer7_outputs(1804) <= a;
    layer7_outputs(1805) <= a;
    layer7_outputs(1806) <= not a;
    layer7_outputs(1807) <= not b;
    layer7_outputs(1808) <= a and not b;
    layer7_outputs(1809) <= b and not a;
    layer7_outputs(1810) <= a xor b;
    layer7_outputs(1811) <= a or b;
    layer7_outputs(1812) <= not (a xor b);
    layer7_outputs(1813) <= a;
    layer7_outputs(1814) <= a and not b;
    layer7_outputs(1815) <= a or b;
    layer7_outputs(1816) <= not b;
    layer7_outputs(1817) <= a xor b;
    layer7_outputs(1818) <= a and not b;
    layer7_outputs(1819) <= a xor b;
    layer7_outputs(1820) <= not (a or b);
    layer7_outputs(1821) <= b and not a;
    layer7_outputs(1822) <= not (a and b);
    layer7_outputs(1823) <= not b;
    layer7_outputs(1824) <= a xor b;
    layer7_outputs(1825) <= not b;
    layer7_outputs(1826) <= not a or b;
    layer7_outputs(1827) <= not a;
    layer7_outputs(1828) <= not a;
    layer7_outputs(1829) <= a xor b;
    layer7_outputs(1830) <= a and b;
    layer7_outputs(1831) <= a;
    layer7_outputs(1832) <= a or b;
    layer7_outputs(1833) <= not a;
    layer7_outputs(1834) <= a;
    layer7_outputs(1835) <= not (a and b);
    layer7_outputs(1836) <= a and b;
    layer7_outputs(1837) <= not a;
    layer7_outputs(1838) <= not (a or b);
    layer7_outputs(1839) <= a xor b;
    layer7_outputs(1840) <= b and not a;
    layer7_outputs(1841) <= a and not b;
    layer7_outputs(1842) <= a and b;
    layer7_outputs(1843) <= not b;
    layer7_outputs(1844) <= b and not a;
    layer7_outputs(1845) <= b;
    layer7_outputs(1846) <= b;
    layer7_outputs(1847) <= a and not b;
    layer7_outputs(1848) <= a or b;
    layer7_outputs(1849) <= not a;
    layer7_outputs(1850) <= not a;
    layer7_outputs(1851) <= b;
    layer7_outputs(1852) <= b;
    layer7_outputs(1853) <= a and not b;
    layer7_outputs(1854) <= '0';
    layer7_outputs(1855) <= not (a or b);
    layer7_outputs(1856) <= b and not a;
    layer7_outputs(1857) <= a xor b;
    layer7_outputs(1858) <= not a;
    layer7_outputs(1859) <= not a;
    layer7_outputs(1860) <= not b;
    layer7_outputs(1861) <= not (a and b);
    layer7_outputs(1862) <= not a or b;
    layer7_outputs(1863) <= not (a xor b);
    layer7_outputs(1864) <= a xor b;
    layer7_outputs(1865) <= b;
    layer7_outputs(1866) <= not (a and b);
    layer7_outputs(1867) <= not b;
    layer7_outputs(1868) <= a;
    layer7_outputs(1869) <= a and not b;
    layer7_outputs(1870) <= not (a xor b);
    layer7_outputs(1871) <= not b;
    layer7_outputs(1872) <= not a;
    layer7_outputs(1873) <= a;
    layer7_outputs(1874) <= not (a xor b);
    layer7_outputs(1875) <= a;
    layer7_outputs(1876) <= a or b;
    layer7_outputs(1877) <= not a;
    layer7_outputs(1878) <= not a;
    layer7_outputs(1879) <= b;
    layer7_outputs(1880) <= a and not b;
    layer7_outputs(1881) <= not a;
    layer7_outputs(1882) <= b;
    layer7_outputs(1883) <= a or b;
    layer7_outputs(1884) <= not (a xor b);
    layer7_outputs(1885) <= a;
    layer7_outputs(1886) <= not (a xor b);
    layer7_outputs(1887) <= '1';
    layer7_outputs(1888) <= not (a and b);
    layer7_outputs(1889) <= not a;
    layer7_outputs(1890) <= a and b;
    layer7_outputs(1891) <= b;
    layer7_outputs(1892) <= a and b;
    layer7_outputs(1893) <= a and b;
    layer7_outputs(1894) <= a;
    layer7_outputs(1895) <= a xor b;
    layer7_outputs(1896) <= b;
    layer7_outputs(1897) <= not (a and b);
    layer7_outputs(1898) <= not (a or b);
    layer7_outputs(1899) <= b and not a;
    layer7_outputs(1900) <= b;
    layer7_outputs(1901) <= b and not a;
    layer7_outputs(1902) <= a;
    layer7_outputs(1903) <= not (a and b);
    layer7_outputs(1904) <= b;
    layer7_outputs(1905) <= a;
    layer7_outputs(1906) <= a xor b;
    layer7_outputs(1907) <= b and not a;
    layer7_outputs(1908) <= not (a xor b);
    layer7_outputs(1909) <= b and not a;
    layer7_outputs(1910) <= not (a xor b);
    layer7_outputs(1911) <= a xor b;
    layer7_outputs(1912) <= not a or b;
    layer7_outputs(1913) <= not a or b;
    layer7_outputs(1914) <= not b;
    layer7_outputs(1915) <= a;
    layer7_outputs(1916) <= not (a and b);
    layer7_outputs(1917) <= not (a xor b);
    layer7_outputs(1918) <= not a;
    layer7_outputs(1919) <= not (a xor b);
    layer7_outputs(1920) <= not (a xor b);
    layer7_outputs(1921) <= a and b;
    layer7_outputs(1922) <= b;
    layer7_outputs(1923) <= a xor b;
    layer7_outputs(1924) <= not (a and b);
    layer7_outputs(1925) <= not a or b;
    layer7_outputs(1926) <= not a;
    layer7_outputs(1927) <= a and not b;
    layer7_outputs(1928) <= a;
    layer7_outputs(1929) <= not (a and b);
    layer7_outputs(1930) <= not b;
    layer7_outputs(1931) <= not (a or b);
    layer7_outputs(1932) <= a and b;
    layer7_outputs(1933) <= a;
    layer7_outputs(1934) <= not a;
    layer7_outputs(1935) <= not (a xor b);
    layer7_outputs(1936) <= '1';
    layer7_outputs(1937) <= a and b;
    layer7_outputs(1938) <= not a;
    layer7_outputs(1939) <= not b or a;
    layer7_outputs(1940) <= a or b;
    layer7_outputs(1941) <= not a;
    layer7_outputs(1942) <= a xor b;
    layer7_outputs(1943) <= b;
    layer7_outputs(1944) <= not b or a;
    layer7_outputs(1945) <= a and b;
    layer7_outputs(1946) <= not (a xor b);
    layer7_outputs(1947) <= not (a xor b);
    layer7_outputs(1948) <= not (a and b);
    layer7_outputs(1949) <= not (a or b);
    layer7_outputs(1950) <= a and b;
    layer7_outputs(1951) <= a;
    layer7_outputs(1952) <= b;
    layer7_outputs(1953) <= not (a or b);
    layer7_outputs(1954) <= b and not a;
    layer7_outputs(1955) <= a;
    layer7_outputs(1956) <= a xor b;
    layer7_outputs(1957) <= not (a xor b);
    layer7_outputs(1958) <= not a;
    layer7_outputs(1959) <= '0';
    layer7_outputs(1960) <= b;
    layer7_outputs(1961) <= not a;
    layer7_outputs(1962) <= not a;
    layer7_outputs(1963) <= a or b;
    layer7_outputs(1964) <= not b;
    layer7_outputs(1965) <= b;
    layer7_outputs(1966) <= not (a and b);
    layer7_outputs(1967) <= not a;
    layer7_outputs(1968) <= not (a or b);
    layer7_outputs(1969) <= not a;
    layer7_outputs(1970) <= not b;
    layer7_outputs(1971) <= a and not b;
    layer7_outputs(1972) <= b;
    layer7_outputs(1973) <= a;
    layer7_outputs(1974) <= not (a xor b);
    layer7_outputs(1975) <= a;
    layer7_outputs(1976) <= not b;
    layer7_outputs(1977) <= not b or a;
    layer7_outputs(1978) <= not (a and b);
    layer7_outputs(1979) <= a and not b;
    layer7_outputs(1980) <= a or b;
    layer7_outputs(1981) <= a xor b;
    layer7_outputs(1982) <= a;
    layer7_outputs(1983) <= not a;
    layer7_outputs(1984) <= a and not b;
    layer7_outputs(1985) <= '1';
    layer7_outputs(1986) <= b;
    layer7_outputs(1987) <= b;
    layer7_outputs(1988) <= b;
    layer7_outputs(1989) <= a;
    layer7_outputs(1990) <= a and b;
    layer7_outputs(1991) <= a;
    layer7_outputs(1992) <= b;
    layer7_outputs(1993) <= b;
    layer7_outputs(1994) <= a and not b;
    layer7_outputs(1995) <= not (a or b);
    layer7_outputs(1996) <= a and not b;
    layer7_outputs(1997) <= not b;
    layer7_outputs(1998) <= a;
    layer7_outputs(1999) <= not a;
    layer7_outputs(2000) <= a and not b;
    layer7_outputs(2001) <= a;
    layer7_outputs(2002) <= not (a and b);
    layer7_outputs(2003) <= not (a or b);
    layer7_outputs(2004) <= '0';
    layer7_outputs(2005) <= a or b;
    layer7_outputs(2006) <= not a or b;
    layer7_outputs(2007) <= a;
    layer7_outputs(2008) <= not b;
    layer7_outputs(2009) <= not (a and b);
    layer7_outputs(2010) <= a;
    layer7_outputs(2011) <= not a or b;
    layer7_outputs(2012) <= '0';
    layer7_outputs(2013) <= not b;
    layer7_outputs(2014) <= not (a and b);
    layer7_outputs(2015) <= not b;
    layer7_outputs(2016) <= a;
    layer7_outputs(2017) <= b;
    layer7_outputs(2018) <= not (a or b);
    layer7_outputs(2019) <= b;
    layer7_outputs(2020) <= not b;
    layer7_outputs(2021) <= a;
    layer7_outputs(2022) <= a xor b;
    layer7_outputs(2023) <= a and not b;
    layer7_outputs(2024) <= b;
    layer7_outputs(2025) <= a xor b;
    layer7_outputs(2026) <= a xor b;
    layer7_outputs(2027) <= b;
    layer7_outputs(2028) <= not a;
    layer7_outputs(2029) <= not a;
    layer7_outputs(2030) <= a;
    layer7_outputs(2031) <= a;
    layer7_outputs(2032) <= not a;
    layer7_outputs(2033) <= not a;
    layer7_outputs(2034) <= not (a xor b);
    layer7_outputs(2035) <= '0';
    layer7_outputs(2036) <= not a;
    layer7_outputs(2037) <= a xor b;
    layer7_outputs(2038) <= not a;
    layer7_outputs(2039) <= a and b;
    layer7_outputs(2040) <= not b;
    layer7_outputs(2041) <= b and not a;
    layer7_outputs(2042) <= not a;
    layer7_outputs(2043) <= b;
    layer7_outputs(2044) <= a or b;
    layer7_outputs(2045) <= not a;
    layer7_outputs(2046) <= not b or a;
    layer7_outputs(2047) <= a and not b;
    layer7_outputs(2048) <= a xor b;
    layer7_outputs(2049) <= not (a or b);
    layer7_outputs(2050) <= not a;
    layer7_outputs(2051) <= a xor b;
    layer7_outputs(2052) <= not a;
    layer7_outputs(2053) <= not b;
    layer7_outputs(2054) <= b;
    layer7_outputs(2055) <= a;
    layer7_outputs(2056) <= not a or b;
    layer7_outputs(2057) <= not b or a;
    layer7_outputs(2058) <= a and not b;
    layer7_outputs(2059) <= a xor b;
    layer7_outputs(2060) <= not (a xor b);
    layer7_outputs(2061) <= not b;
    layer7_outputs(2062) <= a and b;
    layer7_outputs(2063) <= not b;
    layer7_outputs(2064) <= a;
    layer7_outputs(2065) <= not b;
    layer7_outputs(2066) <= not (a xor b);
    layer7_outputs(2067) <= a and not b;
    layer7_outputs(2068) <= a or b;
    layer7_outputs(2069) <= a and b;
    layer7_outputs(2070) <= not b;
    layer7_outputs(2071) <= a;
    layer7_outputs(2072) <= b;
    layer7_outputs(2073) <= not (a xor b);
    layer7_outputs(2074) <= b;
    layer7_outputs(2075) <= not (a xor b);
    layer7_outputs(2076) <= b;
    layer7_outputs(2077) <= not b;
    layer7_outputs(2078) <= not (a and b);
    layer7_outputs(2079) <= not (a or b);
    layer7_outputs(2080) <= a and b;
    layer7_outputs(2081) <= not b;
    layer7_outputs(2082) <= b;
    layer7_outputs(2083) <= '0';
    layer7_outputs(2084) <= not b;
    layer7_outputs(2085) <= not b;
    layer7_outputs(2086) <= b;
    layer7_outputs(2087) <= not (a or b);
    layer7_outputs(2088) <= not a or b;
    layer7_outputs(2089) <= b and not a;
    layer7_outputs(2090) <= a xor b;
    layer7_outputs(2091) <= a and b;
    layer7_outputs(2092) <= a xor b;
    layer7_outputs(2093) <= a;
    layer7_outputs(2094) <= a xor b;
    layer7_outputs(2095) <= not (a or b);
    layer7_outputs(2096) <= b;
    layer7_outputs(2097) <= not (a and b);
    layer7_outputs(2098) <= a and not b;
    layer7_outputs(2099) <= not a or b;
    layer7_outputs(2100) <= b;
    layer7_outputs(2101) <= a or b;
    layer7_outputs(2102) <= not b;
    layer7_outputs(2103) <= not (a and b);
    layer7_outputs(2104) <= a;
    layer7_outputs(2105) <= not b or a;
    layer7_outputs(2106) <= a;
    layer7_outputs(2107) <= b;
    layer7_outputs(2108) <= b;
    layer7_outputs(2109) <= not a or b;
    layer7_outputs(2110) <= a xor b;
    layer7_outputs(2111) <= not a;
    layer7_outputs(2112) <= not b;
    layer7_outputs(2113) <= b and not a;
    layer7_outputs(2114) <= b;
    layer7_outputs(2115) <= b;
    layer7_outputs(2116) <= a;
    layer7_outputs(2117) <= not a or b;
    layer7_outputs(2118) <= a;
    layer7_outputs(2119) <= not a;
    layer7_outputs(2120) <= not a;
    layer7_outputs(2121) <= not (a xor b);
    layer7_outputs(2122) <= a xor b;
    layer7_outputs(2123) <= '1';
    layer7_outputs(2124) <= not a or b;
    layer7_outputs(2125) <= not b or a;
    layer7_outputs(2126) <= not a;
    layer7_outputs(2127) <= a;
    layer7_outputs(2128) <= not a or b;
    layer7_outputs(2129) <= b;
    layer7_outputs(2130) <= not b;
    layer7_outputs(2131) <= not a;
    layer7_outputs(2132) <= not b or a;
    layer7_outputs(2133) <= not (a or b);
    layer7_outputs(2134) <= a and not b;
    layer7_outputs(2135) <= not (a or b);
    layer7_outputs(2136) <= not (a and b);
    layer7_outputs(2137) <= not b;
    layer7_outputs(2138) <= a;
    layer7_outputs(2139) <= not a;
    layer7_outputs(2140) <= a xor b;
    layer7_outputs(2141) <= not (a or b);
    layer7_outputs(2142) <= b;
    layer7_outputs(2143) <= a and not b;
    layer7_outputs(2144) <= b and not a;
    layer7_outputs(2145) <= a or b;
    layer7_outputs(2146) <= a xor b;
    layer7_outputs(2147) <= a and not b;
    layer7_outputs(2148) <= b;
    layer7_outputs(2149) <= not (a xor b);
    layer7_outputs(2150) <= a and not b;
    layer7_outputs(2151) <= not b;
    layer7_outputs(2152) <= b;
    layer7_outputs(2153) <= not a;
    layer7_outputs(2154) <= not b or a;
    layer7_outputs(2155) <= a;
    layer7_outputs(2156) <= not (a xor b);
    layer7_outputs(2157) <= b and not a;
    layer7_outputs(2158) <= a;
    layer7_outputs(2159) <= not (a or b);
    layer7_outputs(2160) <= b;
    layer7_outputs(2161) <= not b;
    layer7_outputs(2162) <= not b;
    layer7_outputs(2163) <= a and b;
    layer7_outputs(2164) <= a xor b;
    layer7_outputs(2165) <= '0';
    layer7_outputs(2166) <= not (a xor b);
    layer7_outputs(2167) <= not b;
    layer7_outputs(2168) <= not b;
    layer7_outputs(2169) <= a;
    layer7_outputs(2170) <= not a;
    layer7_outputs(2171) <= a and not b;
    layer7_outputs(2172) <= not b;
    layer7_outputs(2173) <= not b;
    layer7_outputs(2174) <= not a or b;
    layer7_outputs(2175) <= a or b;
    layer7_outputs(2176) <= not a;
    layer7_outputs(2177) <= not a;
    layer7_outputs(2178) <= not b or a;
    layer7_outputs(2179) <= a;
    layer7_outputs(2180) <= not b;
    layer7_outputs(2181) <= a and b;
    layer7_outputs(2182) <= not a;
    layer7_outputs(2183) <= a or b;
    layer7_outputs(2184) <= a or b;
    layer7_outputs(2185) <= not a;
    layer7_outputs(2186) <= b;
    layer7_outputs(2187) <= b;
    layer7_outputs(2188) <= not a;
    layer7_outputs(2189) <= a;
    layer7_outputs(2190) <= not b;
    layer7_outputs(2191) <= not b;
    layer7_outputs(2192) <= not a;
    layer7_outputs(2193) <= a and b;
    layer7_outputs(2194) <= not a;
    layer7_outputs(2195) <= not (a and b);
    layer7_outputs(2196) <= not b or a;
    layer7_outputs(2197) <= not (a or b);
    layer7_outputs(2198) <= a;
    layer7_outputs(2199) <= a;
    layer7_outputs(2200) <= a or b;
    layer7_outputs(2201) <= b;
    layer7_outputs(2202) <= b and not a;
    layer7_outputs(2203) <= not b;
    layer7_outputs(2204) <= not b;
    layer7_outputs(2205) <= a xor b;
    layer7_outputs(2206) <= not (a xor b);
    layer7_outputs(2207) <= a or b;
    layer7_outputs(2208) <= not a;
    layer7_outputs(2209) <= a;
    layer7_outputs(2210) <= not a;
    layer7_outputs(2211) <= not (a and b);
    layer7_outputs(2212) <= not (a xor b);
    layer7_outputs(2213) <= not (a and b);
    layer7_outputs(2214) <= not (a xor b);
    layer7_outputs(2215) <= not (a xor b);
    layer7_outputs(2216) <= not a;
    layer7_outputs(2217) <= a;
    layer7_outputs(2218) <= not b;
    layer7_outputs(2219) <= not b or a;
    layer7_outputs(2220) <= a;
    layer7_outputs(2221) <= not a;
    layer7_outputs(2222) <= not (a xor b);
    layer7_outputs(2223) <= not (a and b);
    layer7_outputs(2224) <= a xor b;
    layer7_outputs(2225) <= not a;
    layer7_outputs(2226) <= not a;
    layer7_outputs(2227) <= '0';
    layer7_outputs(2228) <= a and b;
    layer7_outputs(2229) <= a and not b;
    layer7_outputs(2230) <= b;
    layer7_outputs(2231) <= not (a or b);
    layer7_outputs(2232) <= a;
    layer7_outputs(2233) <= not b;
    layer7_outputs(2234) <= b;
    layer7_outputs(2235) <= a and b;
    layer7_outputs(2236) <= a xor b;
    layer7_outputs(2237) <= a;
    layer7_outputs(2238) <= a;
    layer7_outputs(2239) <= b;
    layer7_outputs(2240) <= not (a and b);
    layer7_outputs(2241) <= not a;
    layer7_outputs(2242) <= not (a and b);
    layer7_outputs(2243) <= a xor b;
    layer7_outputs(2244) <= a or b;
    layer7_outputs(2245) <= not (a and b);
    layer7_outputs(2246) <= not a;
    layer7_outputs(2247) <= not (a and b);
    layer7_outputs(2248) <= not a;
    layer7_outputs(2249) <= not a;
    layer7_outputs(2250) <= a or b;
    layer7_outputs(2251) <= not (a or b);
    layer7_outputs(2252) <= not b;
    layer7_outputs(2253) <= a and b;
    layer7_outputs(2254) <= b;
    layer7_outputs(2255) <= not a or b;
    layer7_outputs(2256) <= a;
    layer7_outputs(2257) <= a;
    layer7_outputs(2258) <= a;
    layer7_outputs(2259) <= not b or a;
    layer7_outputs(2260) <= not b;
    layer7_outputs(2261) <= a and not b;
    layer7_outputs(2262) <= not a or b;
    layer7_outputs(2263) <= a and b;
    layer7_outputs(2264) <= a and not b;
    layer7_outputs(2265) <= '1';
    layer7_outputs(2266) <= not b;
    layer7_outputs(2267) <= b;
    layer7_outputs(2268) <= not (a xor b);
    layer7_outputs(2269) <= not b;
    layer7_outputs(2270) <= not a or b;
    layer7_outputs(2271) <= a xor b;
    layer7_outputs(2272) <= b and not a;
    layer7_outputs(2273) <= not b;
    layer7_outputs(2274) <= not b or a;
    layer7_outputs(2275) <= not b or a;
    layer7_outputs(2276) <= not a or b;
    layer7_outputs(2277) <= not (a and b);
    layer7_outputs(2278) <= a;
    layer7_outputs(2279) <= not a;
    layer7_outputs(2280) <= not a or b;
    layer7_outputs(2281) <= b;
    layer7_outputs(2282) <= b;
    layer7_outputs(2283) <= not (a xor b);
    layer7_outputs(2284) <= b;
    layer7_outputs(2285) <= not (a and b);
    layer7_outputs(2286) <= not a;
    layer7_outputs(2287) <= not (a and b);
    layer7_outputs(2288) <= a xor b;
    layer7_outputs(2289) <= b;
    layer7_outputs(2290) <= not a or b;
    layer7_outputs(2291) <= not (a and b);
    layer7_outputs(2292) <= '1';
    layer7_outputs(2293) <= a;
    layer7_outputs(2294) <= a and not b;
    layer7_outputs(2295) <= not (a or b);
    layer7_outputs(2296) <= a;
    layer7_outputs(2297) <= not (a and b);
    layer7_outputs(2298) <= not a;
    layer7_outputs(2299) <= not (a or b);
    layer7_outputs(2300) <= a xor b;
    layer7_outputs(2301) <= b;
    layer7_outputs(2302) <= a xor b;
    layer7_outputs(2303) <= b;
    layer7_outputs(2304) <= a and b;
    layer7_outputs(2305) <= not a;
    layer7_outputs(2306) <= a and b;
    layer7_outputs(2307) <= a and not b;
    layer7_outputs(2308) <= not (a and b);
    layer7_outputs(2309) <= a xor b;
    layer7_outputs(2310) <= not a;
    layer7_outputs(2311) <= a;
    layer7_outputs(2312) <= b and not a;
    layer7_outputs(2313) <= a and b;
    layer7_outputs(2314) <= a;
    layer7_outputs(2315) <= a and b;
    layer7_outputs(2316) <= not a;
    layer7_outputs(2317) <= b;
    layer7_outputs(2318) <= not (a xor b);
    layer7_outputs(2319) <= a;
    layer7_outputs(2320) <= not a or b;
    layer7_outputs(2321) <= not b;
    layer7_outputs(2322) <= not b;
    layer7_outputs(2323) <= a;
    layer7_outputs(2324) <= not a or b;
    layer7_outputs(2325) <= not (a xor b);
    layer7_outputs(2326) <= b and not a;
    layer7_outputs(2327) <= a and not b;
    layer7_outputs(2328) <= not b or a;
    layer7_outputs(2329) <= b and not a;
    layer7_outputs(2330) <= not a;
    layer7_outputs(2331) <= not (a xor b);
    layer7_outputs(2332) <= not (a or b);
    layer7_outputs(2333) <= not b;
    layer7_outputs(2334) <= not a;
    layer7_outputs(2335) <= not b;
    layer7_outputs(2336) <= not b;
    layer7_outputs(2337) <= not a;
    layer7_outputs(2338) <= not b or a;
    layer7_outputs(2339) <= '1';
    layer7_outputs(2340) <= not (a or b);
    layer7_outputs(2341) <= not (a or b);
    layer7_outputs(2342) <= not a or b;
    layer7_outputs(2343) <= a;
    layer7_outputs(2344) <= b;
    layer7_outputs(2345) <= not (a xor b);
    layer7_outputs(2346) <= not (a and b);
    layer7_outputs(2347) <= a xor b;
    layer7_outputs(2348) <= a and not b;
    layer7_outputs(2349) <= not b or a;
    layer7_outputs(2350) <= b and not a;
    layer7_outputs(2351) <= a;
    layer7_outputs(2352) <= not b;
    layer7_outputs(2353) <= a and b;
    layer7_outputs(2354) <= a xor b;
    layer7_outputs(2355) <= not b or a;
    layer7_outputs(2356) <= not b or a;
    layer7_outputs(2357) <= not a;
    layer7_outputs(2358) <= b;
    layer7_outputs(2359) <= not (a and b);
    layer7_outputs(2360) <= a or b;
    layer7_outputs(2361) <= a or b;
    layer7_outputs(2362) <= not a;
    layer7_outputs(2363) <= a and not b;
    layer7_outputs(2364) <= a;
    layer7_outputs(2365) <= not (a or b);
    layer7_outputs(2366) <= not b;
    layer7_outputs(2367) <= b;
    layer7_outputs(2368) <= a;
    layer7_outputs(2369) <= not (a and b);
    layer7_outputs(2370) <= a xor b;
    layer7_outputs(2371) <= not b or a;
    layer7_outputs(2372) <= b and not a;
    layer7_outputs(2373) <= a xor b;
    layer7_outputs(2374) <= not b;
    layer7_outputs(2375) <= not (a xor b);
    layer7_outputs(2376) <= a;
    layer7_outputs(2377) <= a and b;
    layer7_outputs(2378) <= a or b;
    layer7_outputs(2379) <= not b;
    layer7_outputs(2380) <= a or b;
    layer7_outputs(2381) <= not b;
    layer7_outputs(2382) <= a;
    layer7_outputs(2383) <= not b;
    layer7_outputs(2384) <= not (a and b);
    layer7_outputs(2385) <= not (a xor b);
    layer7_outputs(2386) <= not b;
    layer7_outputs(2387) <= b;
    layer7_outputs(2388) <= a and b;
    layer7_outputs(2389) <= b and not a;
    layer7_outputs(2390) <= a;
    layer7_outputs(2391) <= a xor b;
    layer7_outputs(2392) <= a;
    layer7_outputs(2393) <= not (a or b);
    layer7_outputs(2394) <= b;
    layer7_outputs(2395) <= not a;
    layer7_outputs(2396) <= a xor b;
    layer7_outputs(2397) <= a and not b;
    layer7_outputs(2398) <= not (a or b);
    layer7_outputs(2399) <= not a or b;
    layer7_outputs(2400) <= a xor b;
    layer7_outputs(2401) <= a;
    layer7_outputs(2402) <= a;
    layer7_outputs(2403) <= a;
    layer7_outputs(2404) <= a or b;
    layer7_outputs(2405) <= b;
    layer7_outputs(2406) <= a xor b;
    layer7_outputs(2407) <= a and not b;
    layer7_outputs(2408) <= not a or b;
    layer7_outputs(2409) <= not b or a;
    layer7_outputs(2410) <= a;
    layer7_outputs(2411) <= a;
    layer7_outputs(2412) <= not a;
    layer7_outputs(2413) <= a or b;
    layer7_outputs(2414) <= a;
    layer7_outputs(2415) <= not b or a;
    layer7_outputs(2416) <= a xor b;
    layer7_outputs(2417) <= b;
    layer7_outputs(2418) <= a;
    layer7_outputs(2419) <= b;
    layer7_outputs(2420) <= b;
    layer7_outputs(2421) <= b;
    layer7_outputs(2422) <= a and not b;
    layer7_outputs(2423) <= b and not a;
    layer7_outputs(2424) <= a or b;
    layer7_outputs(2425) <= b;
    layer7_outputs(2426) <= a and b;
    layer7_outputs(2427) <= not (a xor b);
    layer7_outputs(2428) <= a xor b;
    layer7_outputs(2429) <= not (a and b);
    layer7_outputs(2430) <= not (a and b);
    layer7_outputs(2431) <= not (a xor b);
    layer7_outputs(2432) <= a and not b;
    layer7_outputs(2433) <= a xor b;
    layer7_outputs(2434) <= a;
    layer7_outputs(2435) <= not a;
    layer7_outputs(2436) <= a;
    layer7_outputs(2437) <= not (a or b);
    layer7_outputs(2438) <= a xor b;
    layer7_outputs(2439) <= b;
    layer7_outputs(2440) <= a xor b;
    layer7_outputs(2441) <= not b;
    layer7_outputs(2442) <= not a or b;
    layer7_outputs(2443) <= b;
    layer7_outputs(2444) <= not (a and b);
    layer7_outputs(2445) <= not b;
    layer7_outputs(2446) <= a;
    layer7_outputs(2447) <= a and not b;
    layer7_outputs(2448) <= a;
    layer7_outputs(2449) <= a;
    layer7_outputs(2450) <= b;
    layer7_outputs(2451) <= a and not b;
    layer7_outputs(2452) <= not b;
    layer7_outputs(2453) <= b;
    layer7_outputs(2454) <= not (a and b);
    layer7_outputs(2455) <= a;
    layer7_outputs(2456) <= not (a or b);
    layer7_outputs(2457) <= not (a or b);
    layer7_outputs(2458) <= a and b;
    layer7_outputs(2459) <= not (a xor b);
    layer7_outputs(2460) <= b and not a;
    layer7_outputs(2461) <= a and not b;
    layer7_outputs(2462) <= a;
    layer7_outputs(2463) <= not (a xor b);
    layer7_outputs(2464) <= not b;
    layer7_outputs(2465) <= a and not b;
    layer7_outputs(2466) <= not (a and b);
    layer7_outputs(2467) <= b and not a;
    layer7_outputs(2468) <= b;
    layer7_outputs(2469) <= not b or a;
    layer7_outputs(2470) <= a and not b;
    layer7_outputs(2471) <= not a;
    layer7_outputs(2472) <= a xor b;
    layer7_outputs(2473) <= a;
    layer7_outputs(2474) <= b;
    layer7_outputs(2475) <= b;
    layer7_outputs(2476) <= not a;
    layer7_outputs(2477) <= b;
    layer7_outputs(2478) <= b;
    layer7_outputs(2479) <= not a;
    layer7_outputs(2480) <= a xor b;
    layer7_outputs(2481) <= a;
    layer7_outputs(2482) <= b;
    layer7_outputs(2483) <= not b;
    layer7_outputs(2484) <= not b;
    layer7_outputs(2485) <= b;
    layer7_outputs(2486) <= not (a and b);
    layer7_outputs(2487) <= not (a and b);
    layer7_outputs(2488) <= not b or a;
    layer7_outputs(2489) <= not b;
    layer7_outputs(2490) <= not a;
    layer7_outputs(2491) <= not a;
    layer7_outputs(2492) <= a and b;
    layer7_outputs(2493) <= a and b;
    layer7_outputs(2494) <= not b;
    layer7_outputs(2495) <= not (a xor b);
    layer7_outputs(2496) <= a;
    layer7_outputs(2497) <= a xor b;
    layer7_outputs(2498) <= a and not b;
    layer7_outputs(2499) <= b;
    layer7_outputs(2500) <= not (a and b);
    layer7_outputs(2501) <= not (a and b);
    layer7_outputs(2502) <= a or b;
    layer7_outputs(2503) <= a and b;
    layer7_outputs(2504) <= not b or a;
    layer7_outputs(2505) <= not b;
    layer7_outputs(2506) <= a and not b;
    layer7_outputs(2507) <= not b or a;
    layer7_outputs(2508) <= a and not b;
    layer7_outputs(2509) <= b and not a;
    layer7_outputs(2510) <= not (a and b);
    layer7_outputs(2511) <= not (a xor b);
    layer7_outputs(2512) <= b;
    layer7_outputs(2513) <= b;
    layer7_outputs(2514) <= a;
    layer7_outputs(2515) <= not b;
    layer7_outputs(2516) <= b;
    layer7_outputs(2517) <= b and not a;
    layer7_outputs(2518) <= not (a or b);
    layer7_outputs(2519) <= not a;
    layer7_outputs(2520) <= a xor b;
    layer7_outputs(2521) <= not b or a;
    layer7_outputs(2522) <= a;
    layer7_outputs(2523) <= b;
    layer7_outputs(2524) <= a;
    layer7_outputs(2525) <= b;
    layer7_outputs(2526) <= a and not b;
    layer7_outputs(2527) <= b;
    layer7_outputs(2528) <= not (a and b);
    layer7_outputs(2529) <= not a or b;
    layer7_outputs(2530) <= b and not a;
    layer7_outputs(2531) <= not (a and b);
    layer7_outputs(2532) <= not a or b;
    layer7_outputs(2533) <= a xor b;
    layer7_outputs(2534) <= b and not a;
    layer7_outputs(2535) <= b;
    layer7_outputs(2536) <= not a or b;
    layer7_outputs(2537) <= not b;
    layer7_outputs(2538) <= b;
    layer7_outputs(2539) <= a xor b;
    layer7_outputs(2540) <= '1';
    layer7_outputs(2541) <= a xor b;
    layer7_outputs(2542) <= '0';
    layer7_outputs(2543) <= a or b;
    layer7_outputs(2544) <= not (a or b);
    layer7_outputs(2545) <= b;
    layer7_outputs(2546) <= a;
    layer7_outputs(2547) <= not b or a;
    layer7_outputs(2548) <= not a;
    layer7_outputs(2549) <= b;
    layer7_outputs(2550) <= not b or a;
    layer7_outputs(2551) <= not b;
    layer7_outputs(2552) <= a and not b;
    layer7_outputs(2553) <= not (a and b);
    layer7_outputs(2554) <= b;
    layer7_outputs(2555) <= a or b;
    layer7_outputs(2556) <= a and not b;
    layer7_outputs(2557) <= not b or a;
    layer7_outputs(2558) <= b;
    layer7_outputs(2559) <= not b;
    layer7_outputs(2560) <= not (a xor b);
    layer7_outputs(2561) <= not (a or b);
    layer7_outputs(2562) <= a and b;
    layer7_outputs(2563) <= a;
    layer7_outputs(2564) <= not b;
    layer7_outputs(2565) <= a and not b;
    layer7_outputs(2566) <= not b;
    layer7_outputs(2567) <= a and not b;
    layer7_outputs(2568) <= not b;
    layer7_outputs(2569) <= a;
    layer7_outputs(2570) <= a or b;
    layer7_outputs(2571) <= not b;
    layer7_outputs(2572) <= a and b;
    layer7_outputs(2573) <= not (a and b);
    layer7_outputs(2574) <= a or b;
    layer7_outputs(2575) <= a and b;
    layer7_outputs(2576) <= b;
    layer7_outputs(2577) <= b;
    layer7_outputs(2578) <= not (a xor b);
    layer7_outputs(2579) <= not a;
    layer7_outputs(2580) <= a or b;
    layer7_outputs(2581) <= not b or a;
    layer7_outputs(2582) <= not a;
    layer7_outputs(2583) <= a or b;
    layer7_outputs(2584) <= a or b;
    layer7_outputs(2585) <= b;
    layer7_outputs(2586) <= a xor b;
    layer7_outputs(2587) <= not a;
    layer7_outputs(2588) <= not a;
    layer7_outputs(2589) <= not b;
    layer7_outputs(2590) <= b;
    layer7_outputs(2591) <= a;
    layer7_outputs(2592) <= not (a and b);
    layer7_outputs(2593) <= not (a or b);
    layer7_outputs(2594) <= '0';
    layer7_outputs(2595) <= not a or b;
    layer7_outputs(2596) <= a or b;
    layer7_outputs(2597) <= not b or a;
    layer7_outputs(2598) <= not a;
    layer7_outputs(2599) <= a xor b;
    layer7_outputs(2600) <= a xor b;
    layer7_outputs(2601) <= a or b;
    layer7_outputs(2602) <= a xor b;
    layer7_outputs(2603) <= not (a xor b);
    layer7_outputs(2604) <= not (a or b);
    layer7_outputs(2605) <= not b;
    layer7_outputs(2606) <= '0';
    layer7_outputs(2607) <= a;
    layer7_outputs(2608) <= b;
    layer7_outputs(2609) <= not a;
    layer7_outputs(2610) <= not a;
    layer7_outputs(2611) <= a and b;
    layer7_outputs(2612) <= a xor b;
    layer7_outputs(2613) <= a xor b;
    layer7_outputs(2614) <= not (a xor b);
    layer7_outputs(2615) <= not b;
    layer7_outputs(2616) <= b;
    layer7_outputs(2617) <= '0';
    layer7_outputs(2618) <= '0';
    layer7_outputs(2619) <= not a or b;
    layer7_outputs(2620) <= b and not a;
    layer7_outputs(2621) <= not b;
    layer7_outputs(2622) <= not (a or b);
    layer7_outputs(2623) <= b;
    layer7_outputs(2624) <= a or b;
    layer7_outputs(2625) <= b;
    layer7_outputs(2626) <= b and not a;
    layer7_outputs(2627) <= not b;
    layer7_outputs(2628) <= b;
    layer7_outputs(2629) <= not b;
    layer7_outputs(2630) <= not (a and b);
    layer7_outputs(2631) <= '1';
    layer7_outputs(2632) <= a xor b;
    layer7_outputs(2633) <= a or b;
    layer7_outputs(2634) <= b and not a;
    layer7_outputs(2635) <= a and not b;
    layer7_outputs(2636) <= not (a and b);
    layer7_outputs(2637) <= b;
    layer7_outputs(2638) <= a;
    layer7_outputs(2639) <= b;
    layer7_outputs(2640) <= a;
    layer7_outputs(2641) <= b;
    layer7_outputs(2642) <= a or b;
    layer7_outputs(2643) <= a or b;
    layer7_outputs(2644) <= a;
    layer7_outputs(2645) <= not b or a;
    layer7_outputs(2646) <= a and not b;
    layer7_outputs(2647) <= a and not b;
    layer7_outputs(2648) <= b;
    layer7_outputs(2649) <= a xor b;
    layer7_outputs(2650) <= not b;
    layer7_outputs(2651) <= not b;
    layer7_outputs(2652) <= not a;
    layer7_outputs(2653) <= not a;
    layer7_outputs(2654) <= a xor b;
    layer7_outputs(2655) <= b;
    layer7_outputs(2656) <= not b or a;
    layer7_outputs(2657) <= a xor b;
    layer7_outputs(2658) <= not a;
    layer7_outputs(2659) <= b;
    layer7_outputs(2660) <= b;
    layer7_outputs(2661) <= not a;
    layer7_outputs(2662) <= a or b;
    layer7_outputs(2663) <= a or b;
    layer7_outputs(2664) <= not (a xor b);
    layer7_outputs(2665) <= a and b;
    layer7_outputs(2666) <= b;
    layer7_outputs(2667) <= not a;
    layer7_outputs(2668) <= not (a xor b);
    layer7_outputs(2669) <= not b;
    layer7_outputs(2670) <= not a;
    layer7_outputs(2671) <= not b;
    layer7_outputs(2672) <= not a;
    layer7_outputs(2673) <= not b or a;
    layer7_outputs(2674) <= not a;
    layer7_outputs(2675) <= not (a and b);
    layer7_outputs(2676) <= a xor b;
    layer7_outputs(2677) <= a and b;
    layer7_outputs(2678) <= a and not b;
    layer7_outputs(2679) <= not (a xor b);
    layer7_outputs(2680) <= b and not a;
    layer7_outputs(2681) <= a;
    layer7_outputs(2682) <= a xor b;
    layer7_outputs(2683) <= b;
    layer7_outputs(2684) <= not b or a;
    layer7_outputs(2685) <= not b;
    layer7_outputs(2686) <= a and not b;
    layer7_outputs(2687) <= a;
    layer7_outputs(2688) <= a;
    layer7_outputs(2689) <= not b or a;
    layer7_outputs(2690) <= not a;
    layer7_outputs(2691) <= a xor b;
    layer7_outputs(2692) <= not a or b;
    layer7_outputs(2693) <= a and b;
    layer7_outputs(2694) <= '1';
    layer7_outputs(2695) <= b;
    layer7_outputs(2696) <= not (a xor b);
    layer7_outputs(2697) <= b;
    layer7_outputs(2698) <= a and not b;
    layer7_outputs(2699) <= not a or b;
    layer7_outputs(2700) <= not (a or b);
    layer7_outputs(2701) <= b;
    layer7_outputs(2702) <= not b;
    layer7_outputs(2703) <= a;
    layer7_outputs(2704) <= not b or a;
    layer7_outputs(2705) <= a and not b;
    layer7_outputs(2706) <= a;
    layer7_outputs(2707) <= b;
    layer7_outputs(2708) <= a and b;
    layer7_outputs(2709) <= b;
    layer7_outputs(2710) <= a;
    layer7_outputs(2711) <= b;
    layer7_outputs(2712) <= b and not a;
    layer7_outputs(2713) <= not b;
    layer7_outputs(2714) <= not (a xor b);
    layer7_outputs(2715) <= a xor b;
    layer7_outputs(2716) <= not (a or b);
    layer7_outputs(2717) <= not (a and b);
    layer7_outputs(2718) <= a;
    layer7_outputs(2719) <= '0';
    layer7_outputs(2720) <= not b;
    layer7_outputs(2721) <= not a or b;
    layer7_outputs(2722) <= not (a xor b);
    layer7_outputs(2723) <= a;
    layer7_outputs(2724) <= not b or a;
    layer7_outputs(2725) <= not (a and b);
    layer7_outputs(2726) <= not b or a;
    layer7_outputs(2727) <= b and not a;
    layer7_outputs(2728) <= not b;
    layer7_outputs(2729) <= a;
    layer7_outputs(2730) <= not b;
    layer7_outputs(2731) <= not a;
    layer7_outputs(2732) <= a;
    layer7_outputs(2733) <= a;
    layer7_outputs(2734) <= '0';
    layer7_outputs(2735) <= a;
    layer7_outputs(2736) <= not b;
    layer7_outputs(2737) <= not (a xor b);
    layer7_outputs(2738) <= a or b;
    layer7_outputs(2739) <= not b;
    layer7_outputs(2740) <= not b;
    layer7_outputs(2741) <= not b;
    layer7_outputs(2742) <= a;
    layer7_outputs(2743) <= not (a or b);
    layer7_outputs(2744) <= b;
    layer7_outputs(2745) <= a and b;
    layer7_outputs(2746) <= not (a xor b);
    layer7_outputs(2747) <= b;
    layer7_outputs(2748) <= not b;
    layer7_outputs(2749) <= a or b;
    layer7_outputs(2750) <= not (a or b);
    layer7_outputs(2751) <= '1';
    layer7_outputs(2752) <= a or b;
    layer7_outputs(2753) <= '1';
    layer7_outputs(2754) <= a and not b;
    layer7_outputs(2755) <= a and not b;
    layer7_outputs(2756) <= b and not a;
    layer7_outputs(2757) <= not a;
    layer7_outputs(2758) <= not (a or b);
    layer7_outputs(2759) <= b;
    layer7_outputs(2760) <= a and not b;
    layer7_outputs(2761) <= a xor b;
    layer7_outputs(2762) <= b;
    layer7_outputs(2763) <= a xor b;
    layer7_outputs(2764) <= b and not a;
    layer7_outputs(2765) <= not a;
    layer7_outputs(2766) <= a;
    layer7_outputs(2767) <= b;
    layer7_outputs(2768) <= b;
    layer7_outputs(2769) <= a and b;
    layer7_outputs(2770) <= a xor b;
    layer7_outputs(2771) <= a and not b;
    layer7_outputs(2772) <= a;
    layer7_outputs(2773) <= a;
    layer7_outputs(2774) <= a;
    layer7_outputs(2775) <= b and not a;
    layer7_outputs(2776) <= not (a xor b);
    layer7_outputs(2777) <= b and not a;
    layer7_outputs(2778) <= a xor b;
    layer7_outputs(2779) <= a and b;
    layer7_outputs(2780) <= not b;
    layer7_outputs(2781) <= not a or b;
    layer7_outputs(2782) <= a and not b;
    layer7_outputs(2783) <= b;
    layer7_outputs(2784) <= a;
    layer7_outputs(2785) <= '1';
    layer7_outputs(2786) <= b;
    layer7_outputs(2787) <= not a or b;
    layer7_outputs(2788) <= a;
    layer7_outputs(2789) <= b;
    layer7_outputs(2790) <= a xor b;
    layer7_outputs(2791) <= not a or b;
    layer7_outputs(2792) <= b and not a;
    layer7_outputs(2793) <= b and not a;
    layer7_outputs(2794) <= a and not b;
    layer7_outputs(2795) <= not b;
    layer7_outputs(2796) <= not b or a;
    layer7_outputs(2797) <= not (a or b);
    layer7_outputs(2798) <= not a or b;
    layer7_outputs(2799) <= b;
    layer7_outputs(2800) <= not (a xor b);
    layer7_outputs(2801) <= not (a xor b);
    layer7_outputs(2802) <= not b;
    layer7_outputs(2803) <= not b;
    layer7_outputs(2804) <= not (a or b);
    layer7_outputs(2805) <= not (a xor b);
    layer7_outputs(2806) <= not a;
    layer7_outputs(2807) <= not a;
    layer7_outputs(2808) <= b and not a;
    layer7_outputs(2809) <= not b or a;
    layer7_outputs(2810) <= not a or b;
    layer7_outputs(2811) <= b;
    layer7_outputs(2812) <= not (a xor b);
    layer7_outputs(2813) <= b;
    layer7_outputs(2814) <= not b or a;
    layer7_outputs(2815) <= a;
    layer7_outputs(2816) <= not (a and b);
    layer7_outputs(2817) <= not a or b;
    layer7_outputs(2818) <= not a;
    layer7_outputs(2819) <= a;
    layer7_outputs(2820) <= not a or b;
    layer7_outputs(2821) <= a;
    layer7_outputs(2822) <= a or b;
    layer7_outputs(2823) <= b;
    layer7_outputs(2824) <= not (a and b);
    layer7_outputs(2825) <= not b;
    layer7_outputs(2826) <= not (a xor b);
    layer7_outputs(2827) <= a and not b;
    layer7_outputs(2828) <= b;
    layer7_outputs(2829) <= not a or b;
    layer7_outputs(2830) <= a xor b;
    layer7_outputs(2831) <= '1';
    layer7_outputs(2832) <= b;
    layer7_outputs(2833) <= a and not b;
    layer7_outputs(2834) <= not (a and b);
    layer7_outputs(2835) <= not (a or b);
    layer7_outputs(2836) <= a;
    layer7_outputs(2837) <= not b;
    layer7_outputs(2838) <= not b or a;
    layer7_outputs(2839) <= not (a and b);
    layer7_outputs(2840) <= not a;
    layer7_outputs(2841) <= not b;
    layer7_outputs(2842) <= not b;
    layer7_outputs(2843) <= a;
    layer7_outputs(2844) <= a;
    layer7_outputs(2845) <= not (a xor b);
    layer7_outputs(2846) <= not b;
    layer7_outputs(2847) <= not a;
    layer7_outputs(2848) <= a;
    layer7_outputs(2849) <= not (a xor b);
    layer7_outputs(2850) <= a xor b;
    layer7_outputs(2851) <= not (a or b);
    layer7_outputs(2852) <= a;
    layer7_outputs(2853) <= not (a xor b);
    layer7_outputs(2854) <= b;
    layer7_outputs(2855) <= not (a and b);
    layer7_outputs(2856) <= b;
    layer7_outputs(2857) <= not b;
    layer7_outputs(2858) <= a and b;
    layer7_outputs(2859) <= a and not b;
    layer7_outputs(2860) <= not (a and b);
    layer7_outputs(2861) <= not (a and b);
    layer7_outputs(2862) <= not b;
    layer7_outputs(2863) <= a xor b;
    layer7_outputs(2864) <= a or b;
    layer7_outputs(2865) <= a;
    layer7_outputs(2866) <= a and not b;
    layer7_outputs(2867) <= not a or b;
    layer7_outputs(2868) <= b;
    layer7_outputs(2869) <= b;
    layer7_outputs(2870) <= not (a or b);
    layer7_outputs(2871) <= not a;
    layer7_outputs(2872) <= a;
    layer7_outputs(2873) <= not b;
    layer7_outputs(2874) <= not a;
    layer7_outputs(2875) <= not b;
    layer7_outputs(2876) <= b;
    layer7_outputs(2877) <= a and b;
    layer7_outputs(2878) <= not a;
    layer7_outputs(2879) <= b;
    layer7_outputs(2880) <= '1';
    layer7_outputs(2881) <= a;
    layer7_outputs(2882) <= not a or b;
    layer7_outputs(2883) <= not (a and b);
    layer7_outputs(2884) <= a xor b;
    layer7_outputs(2885) <= not b;
    layer7_outputs(2886) <= not b or a;
    layer7_outputs(2887) <= b;
    layer7_outputs(2888) <= not (a and b);
    layer7_outputs(2889) <= not (a xor b);
    layer7_outputs(2890) <= a or b;
    layer7_outputs(2891) <= not (a and b);
    layer7_outputs(2892) <= not a;
    layer7_outputs(2893) <= b and not a;
    layer7_outputs(2894) <= b;
    layer7_outputs(2895) <= not b or a;
    layer7_outputs(2896) <= not (a xor b);
    layer7_outputs(2897) <= not a;
    layer7_outputs(2898) <= a;
    layer7_outputs(2899) <= not (a or b);
    layer7_outputs(2900) <= a xor b;
    layer7_outputs(2901) <= b and not a;
    layer7_outputs(2902) <= a or b;
    layer7_outputs(2903) <= not b;
    layer7_outputs(2904) <= a xor b;
    layer7_outputs(2905) <= not (a and b);
    layer7_outputs(2906) <= a;
    layer7_outputs(2907) <= not (a xor b);
    layer7_outputs(2908) <= not (a xor b);
    layer7_outputs(2909) <= a or b;
    layer7_outputs(2910) <= not a;
    layer7_outputs(2911) <= b;
    layer7_outputs(2912) <= not a;
    layer7_outputs(2913) <= '1';
    layer7_outputs(2914) <= not b;
    layer7_outputs(2915) <= not a;
    layer7_outputs(2916) <= a xor b;
    layer7_outputs(2917) <= not a or b;
    layer7_outputs(2918) <= not b;
    layer7_outputs(2919) <= not a;
    layer7_outputs(2920) <= not a;
    layer7_outputs(2921) <= b;
    layer7_outputs(2922) <= not b or a;
    layer7_outputs(2923) <= a xor b;
    layer7_outputs(2924) <= not (a xor b);
    layer7_outputs(2925) <= not b;
    layer7_outputs(2926) <= a xor b;
    layer7_outputs(2927) <= not a;
    layer7_outputs(2928) <= a;
    layer7_outputs(2929) <= b;
    layer7_outputs(2930) <= a and not b;
    layer7_outputs(2931) <= '1';
    layer7_outputs(2932) <= a and b;
    layer7_outputs(2933) <= not (a or b);
    layer7_outputs(2934) <= b;
    layer7_outputs(2935) <= b;
    layer7_outputs(2936) <= '1';
    layer7_outputs(2937) <= a xor b;
    layer7_outputs(2938) <= a;
    layer7_outputs(2939) <= a and not b;
    layer7_outputs(2940) <= not b;
    layer7_outputs(2941) <= not (a or b);
    layer7_outputs(2942) <= a;
    layer7_outputs(2943) <= b and not a;
    layer7_outputs(2944) <= not (a xor b);
    layer7_outputs(2945) <= a or b;
    layer7_outputs(2946) <= a and not b;
    layer7_outputs(2947) <= b;
    layer7_outputs(2948) <= a;
    layer7_outputs(2949) <= not (a and b);
    layer7_outputs(2950) <= b;
    layer7_outputs(2951) <= not a;
    layer7_outputs(2952) <= not (a and b);
    layer7_outputs(2953) <= not b or a;
    layer7_outputs(2954) <= not a or b;
    layer7_outputs(2955) <= b and not a;
    layer7_outputs(2956) <= b and not a;
    layer7_outputs(2957) <= a xor b;
    layer7_outputs(2958) <= not b;
    layer7_outputs(2959) <= a or b;
    layer7_outputs(2960) <= a and b;
    layer7_outputs(2961) <= b and not a;
    layer7_outputs(2962) <= not a or b;
    layer7_outputs(2963) <= '1';
    layer7_outputs(2964) <= '1';
    layer7_outputs(2965) <= b;
    layer7_outputs(2966) <= not a or b;
    layer7_outputs(2967) <= a and b;
    layer7_outputs(2968) <= not a;
    layer7_outputs(2969) <= not a;
    layer7_outputs(2970) <= '0';
    layer7_outputs(2971) <= b and not a;
    layer7_outputs(2972) <= not b;
    layer7_outputs(2973) <= a or b;
    layer7_outputs(2974) <= not b;
    layer7_outputs(2975) <= not (a xor b);
    layer7_outputs(2976) <= not b;
    layer7_outputs(2977) <= a;
    layer7_outputs(2978) <= a;
    layer7_outputs(2979) <= a;
    layer7_outputs(2980) <= not (a or b);
    layer7_outputs(2981) <= not b;
    layer7_outputs(2982) <= not a or b;
    layer7_outputs(2983) <= not (a xor b);
    layer7_outputs(2984) <= not b;
    layer7_outputs(2985) <= not a;
    layer7_outputs(2986) <= a and b;
    layer7_outputs(2987) <= not b or a;
    layer7_outputs(2988) <= not b;
    layer7_outputs(2989) <= not a;
    layer7_outputs(2990) <= not a;
    layer7_outputs(2991) <= a and b;
    layer7_outputs(2992) <= a and b;
    layer7_outputs(2993) <= not b;
    layer7_outputs(2994) <= b and not a;
    layer7_outputs(2995) <= a;
    layer7_outputs(2996) <= a;
    layer7_outputs(2997) <= b and not a;
    layer7_outputs(2998) <= not (a or b);
    layer7_outputs(2999) <= not a;
    layer7_outputs(3000) <= not b or a;
    layer7_outputs(3001) <= not b or a;
    layer7_outputs(3002) <= not a;
    layer7_outputs(3003) <= a or b;
    layer7_outputs(3004) <= not (a xor b);
    layer7_outputs(3005) <= not b or a;
    layer7_outputs(3006) <= not b;
    layer7_outputs(3007) <= '0';
    layer7_outputs(3008) <= a and not b;
    layer7_outputs(3009) <= not (a or b);
    layer7_outputs(3010) <= not a or b;
    layer7_outputs(3011) <= b and not a;
    layer7_outputs(3012) <= a and not b;
    layer7_outputs(3013) <= not a;
    layer7_outputs(3014) <= b;
    layer7_outputs(3015) <= not a;
    layer7_outputs(3016) <= a and b;
    layer7_outputs(3017) <= not b;
    layer7_outputs(3018) <= not (a xor b);
    layer7_outputs(3019) <= a;
    layer7_outputs(3020) <= not (a or b);
    layer7_outputs(3021) <= b;
    layer7_outputs(3022) <= a and not b;
    layer7_outputs(3023) <= not b;
    layer7_outputs(3024) <= b and not a;
    layer7_outputs(3025) <= not b;
    layer7_outputs(3026) <= a xor b;
    layer7_outputs(3027) <= not a;
    layer7_outputs(3028) <= not (a and b);
    layer7_outputs(3029) <= not a or b;
    layer7_outputs(3030) <= a xor b;
    layer7_outputs(3031) <= a and not b;
    layer7_outputs(3032) <= a xor b;
    layer7_outputs(3033) <= a xor b;
    layer7_outputs(3034) <= not (a or b);
    layer7_outputs(3035) <= not (a or b);
    layer7_outputs(3036) <= not (a xor b);
    layer7_outputs(3037) <= b;
    layer7_outputs(3038) <= a and not b;
    layer7_outputs(3039) <= a and b;
    layer7_outputs(3040) <= not (a xor b);
    layer7_outputs(3041) <= a and b;
    layer7_outputs(3042) <= not b;
    layer7_outputs(3043) <= a and b;
    layer7_outputs(3044) <= a and not b;
    layer7_outputs(3045) <= a and b;
    layer7_outputs(3046) <= a xor b;
    layer7_outputs(3047) <= not (a and b);
    layer7_outputs(3048) <= not (a or b);
    layer7_outputs(3049) <= a;
    layer7_outputs(3050) <= not a or b;
    layer7_outputs(3051) <= b;
    layer7_outputs(3052) <= not a or b;
    layer7_outputs(3053) <= not (a and b);
    layer7_outputs(3054) <= a;
    layer7_outputs(3055) <= not b or a;
    layer7_outputs(3056) <= '0';
    layer7_outputs(3057) <= not b or a;
    layer7_outputs(3058) <= not b;
    layer7_outputs(3059) <= a or b;
    layer7_outputs(3060) <= a or b;
    layer7_outputs(3061) <= a;
    layer7_outputs(3062) <= not a or b;
    layer7_outputs(3063) <= a;
    layer7_outputs(3064) <= not a;
    layer7_outputs(3065) <= not (a xor b);
    layer7_outputs(3066) <= b and not a;
    layer7_outputs(3067) <= not a;
    layer7_outputs(3068) <= not b or a;
    layer7_outputs(3069) <= a and not b;
    layer7_outputs(3070) <= a and not b;
    layer7_outputs(3071) <= b;
    layer7_outputs(3072) <= '1';
    layer7_outputs(3073) <= a and not b;
    layer7_outputs(3074) <= not a;
    layer7_outputs(3075) <= not a;
    layer7_outputs(3076) <= not (a xor b);
    layer7_outputs(3077) <= b;
    layer7_outputs(3078) <= not a or b;
    layer7_outputs(3079) <= not a;
    layer7_outputs(3080) <= not a;
    layer7_outputs(3081) <= not (a or b);
    layer7_outputs(3082) <= a;
    layer7_outputs(3083) <= not (a xor b);
    layer7_outputs(3084) <= not b or a;
    layer7_outputs(3085) <= a;
    layer7_outputs(3086) <= not a or b;
    layer7_outputs(3087) <= '1';
    layer7_outputs(3088) <= not a or b;
    layer7_outputs(3089) <= a and b;
    layer7_outputs(3090) <= b;
    layer7_outputs(3091) <= a and not b;
    layer7_outputs(3092) <= a and b;
    layer7_outputs(3093) <= not (a xor b);
    layer7_outputs(3094) <= not a or b;
    layer7_outputs(3095) <= not a or b;
    layer7_outputs(3096) <= not (a or b);
    layer7_outputs(3097) <= a xor b;
    layer7_outputs(3098) <= not b;
    layer7_outputs(3099) <= a;
    layer7_outputs(3100) <= not a;
    layer7_outputs(3101) <= a or b;
    layer7_outputs(3102) <= a xor b;
    layer7_outputs(3103) <= not a;
    layer7_outputs(3104) <= not (a xor b);
    layer7_outputs(3105) <= a and not b;
    layer7_outputs(3106) <= '0';
    layer7_outputs(3107) <= b;
    layer7_outputs(3108) <= a or b;
    layer7_outputs(3109) <= a and not b;
    layer7_outputs(3110) <= a xor b;
    layer7_outputs(3111) <= b;
    layer7_outputs(3112) <= not (a or b);
    layer7_outputs(3113) <= not b;
    layer7_outputs(3114) <= not b;
    layer7_outputs(3115) <= not a;
    layer7_outputs(3116) <= '0';
    layer7_outputs(3117) <= a and b;
    layer7_outputs(3118) <= a;
    layer7_outputs(3119) <= b and not a;
    layer7_outputs(3120) <= b and not a;
    layer7_outputs(3121) <= a;
    layer7_outputs(3122) <= not (a or b);
    layer7_outputs(3123) <= not (a xor b);
    layer7_outputs(3124) <= not b;
    layer7_outputs(3125) <= not (a xor b);
    layer7_outputs(3126) <= not a;
    layer7_outputs(3127) <= a;
    layer7_outputs(3128) <= not a or b;
    layer7_outputs(3129) <= b and not a;
    layer7_outputs(3130) <= a xor b;
    layer7_outputs(3131) <= a and b;
    layer7_outputs(3132) <= not b;
    layer7_outputs(3133) <= a and b;
    layer7_outputs(3134) <= not a;
    layer7_outputs(3135) <= not (a xor b);
    layer7_outputs(3136) <= a;
    layer7_outputs(3137) <= a or b;
    layer7_outputs(3138) <= a and not b;
    layer7_outputs(3139) <= a and b;
    layer7_outputs(3140) <= b and not a;
    layer7_outputs(3141) <= not (a or b);
    layer7_outputs(3142) <= not (a and b);
    layer7_outputs(3143) <= a;
    layer7_outputs(3144) <= b;
    layer7_outputs(3145) <= a xor b;
    layer7_outputs(3146) <= a;
    layer7_outputs(3147) <= a xor b;
    layer7_outputs(3148) <= not b;
    layer7_outputs(3149) <= not (a xor b);
    layer7_outputs(3150) <= not b;
    layer7_outputs(3151) <= not a;
    layer7_outputs(3152) <= a;
    layer7_outputs(3153) <= a and b;
    layer7_outputs(3154) <= a or b;
    layer7_outputs(3155) <= not a or b;
    layer7_outputs(3156) <= a or b;
    layer7_outputs(3157) <= not a;
    layer7_outputs(3158) <= a xor b;
    layer7_outputs(3159) <= a and not b;
    layer7_outputs(3160) <= not b;
    layer7_outputs(3161) <= b;
    layer7_outputs(3162) <= not (a or b);
    layer7_outputs(3163) <= a and b;
    layer7_outputs(3164) <= a;
    layer7_outputs(3165) <= not a or b;
    layer7_outputs(3166) <= b;
    layer7_outputs(3167) <= not b;
    layer7_outputs(3168) <= '0';
    layer7_outputs(3169) <= not (a and b);
    layer7_outputs(3170) <= not b;
    layer7_outputs(3171) <= a xor b;
    layer7_outputs(3172) <= a or b;
    layer7_outputs(3173) <= not a;
    layer7_outputs(3174) <= a xor b;
    layer7_outputs(3175) <= a;
    layer7_outputs(3176) <= b;
    layer7_outputs(3177) <= not (a or b);
    layer7_outputs(3178) <= a;
    layer7_outputs(3179) <= '0';
    layer7_outputs(3180) <= a;
    layer7_outputs(3181) <= not b;
    layer7_outputs(3182) <= not a or b;
    layer7_outputs(3183) <= not (a xor b);
    layer7_outputs(3184) <= a;
    layer7_outputs(3185) <= a xor b;
    layer7_outputs(3186) <= not (a or b);
    layer7_outputs(3187) <= a or b;
    layer7_outputs(3188) <= a and b;
    layer7_outputs(3189) <= a and not b;
    layer7_outputs(3190) <= b and not a;
    layer7_outputs(3191) <= not b or a;
    layer7_outputs(3192) <= a;
    layer7_outputs(3193) <= a;
    layer7_outputs(3194) <= b;
    layer7_outputs(3195) <= not a;
    layer7_outputs(3196) <= a;
    layer7_outputs(3197) <= not (a xor b);
    layer7_outputs(3198) <= a or b;
    layer7_outputs(3199) <= b;
    layer7_outputs(3200) <= b;
    layer7_outputs(3201) <= a xor b;
    layer7_outputs(3202) <= not b or a;
    layer7_outputs(3203) <= not a;
    layer7_outputs(3204) <= not (a xor b);
    layer7_outputs(3205) <= a and not b;
    layer7_outputs(3206) <= not a or b;
    layer7_outputs(3207) <= b and not a;
    layer7_outputs(3208) <= not b;
    layer7_outputs(3209) <= not (a xor b);
    layer7_outputs(3210) <= a xor b;
    layer7_outputs(3211) <= not (a or b);
    layer7_outputs(3212) <= not b;
    layer7_outputs(3213) <= not (a xor b);
    layer7_outputs(3214) <= b and not a;
    layer7_outputs(3215) <= b;
    layer7_outputs(3216) <= not b or a;
    layer7_outputs(3217) <= '1';
    layer7_outputs(3218) <= not a;
    layer7_outputs(3219) <= a and not b;
    layer7_outputs(3220) <= not (a and b);
    layer7_outputs(3221) <= not (a or b);
    layer7_outputs(3222) <= a xor b;
    layer7_outputs(3223) <= not b;
    layer7_outputs(3224) <= not (a or b);
    layer7_outputs(3225) <= a;
    layer7_outputs(3226) <= b;
    layer7_outputs(3227) <= not (a or b);
    layer7_outputs(3228) <= a;
    layer7_outputs(3229) <= not (a or b);
    layer7_outputs(3230) <= '0';
    layer7_outputs(3231) <= not a or b;
    layer7_outputs(3232) <= a and b;
    layer7_outputs(3233) <= not (a and b);
    layer7_outputs(3234) <= b;
    layer7_outputs(3235) <= a;
    layer7_outputs(3236) <= a or b;
    layer7_outputs(3237) <= b;
    layer7_outputs(3238) <= not (a or b);
    layer7_outputs(3239) <= '1';
    layer7_outputs(3240) <= a;
    layer7_outputs(3241) <= b;
    layer7_outputs(3242) <= not (a xor b);
    layer7_outputs(3243) <= b;
    layer7_outputs(3244) <= not (a or b);
    layer7_outputs(3245) <= b;
    layer7_outputs(3246) <= not b;
    layer7_outputs(3247) <= a and not b;
    layer7_outputs(3248) <= b and not a;
    layer7_outputs(3249) <= not b or a;
    layer7_outputs(3250) <= a xor b;
    layer7_outputs(3251) <= b;
    layer7_outputs(3252) <= not a;
    layer7_outputs(3253) <= a and not b;
    layer7_outputs(3254) <= not a;
    layer7_outputs(3255) <= not (a or b);
    layer7_outputs(3256) <= not b;
    layer7_outputs(3257) <= a and b;
    layer7_outputs(3258) <= a and b;
    layer7_outputs(3259) <= a;
    layer7_outputs(3260) <= a xor b;
    layer7_outputs(3261) <= a;
    layer7_outputs(3262) <= b and not a;
    layer7_outputs(3263) <= not (a xor b);
    layer7_outputs(3264) <= not (a and b);
    layer7_outputs(3265) <= not a;
    layer7_outputs(3266) <= a and not b;
    layer7_outputs(3267) <= not (a xor b);
    layer7_outputs(3268) <= a;
    layer7_outputs(3269) <= a xor b;
    layer7_outputs(3270) <= b and not a;
    layer7_outputs(3271) <= a xor b;
    layer7_outputs(3272) <= a xor b;
    layer7_outputs(3273) <= a;
    layer7_outputs(3274) <= not a;
    layer7_outputs(3275) <= b;
    layer7_outputs(3276) <= a and b;
    layer7_outputs(3277) <= not (a or b);
    layer7_outputs(3278) <= not (a or b);
    layer7_outputs(3279) <= not a or b;
    layer7_outputs(3280) <= a;
    layer7_outputs(3281) <= not (a xor b);
    layer7_outputs(3282) <= not b;
    layer7_outputs(3283) <= not b;
    layer7_outputs(3284) <= not b or a;
    layer7_outputs(3285) <= not b;
    layer7_outputs(3286) <= not b or a;
    layer7_outputs(3287) <= not a;
    layer7_outputs(3288) <= not a;
    layer7_outputs(3289) <= a;
    layer7_outputs(3290) <= not b;
    layer7_outputs(3291) <= a xor b;
    layer7_outputs(3292) <= not (a xor b);
    layer7_outputs(3293) <= not b;
    layer7_outputs(3294) <= not (a and b);
    layer7_outputs(3295) <= a or b;
    layer7_outputs(3296) <= a xor b;
    layer7_outputs(3297) <= b;
    layer7_outputs(3298) <= a or b;
    layer7_outputs(3299) <= not b or a;
    layer7_outputs(3300) <= not b or a;
    layer7_outputs(3301) <= a;
    layer7_outputs(3302) <= b;
    layer7_outputs(3303) <= not (a xor b);
    layer7_outputs(3304) <= not a;
    layer7_outputs(3305) <= not (a or b);
    layer7_outputs(3306) <= not a;
    layer7_outputs(3307) <= a;
    layer7_outputs(3308) <= not (a or b);
    layer7_outputs(3309) <= a or b;
    layer7_outputs(3310) <= a;
    layer7_outputs(3311) <= not b;
    layer7_outputs(3312) <= not a;
    layer7_outputs(3313) <= not b or a;
    layer7_outputs(3314) <= not b;
    layer7_outputs(3315) <= not b;
    layer7_outputs(3316) <= a;
    layer7_outputs(3317) <= a;
    layer7_outputs(3318) <= not (a or b);
    layer7_outputs(3319) <= not b or a;
    layer7_outputs(3320) <= b;
    layer7_outputs(3321) <= not (a and b);
    layer7_outputs(3322) <= not b;
    layer7_outputs(3323) <= not (a xor b);
    layer7_outputs(3324) <= a;
    layer7_outputs(3325) <= not b;
    layer7_outputs(3326) <= not b;
    layer7_outputs(3327) <= b;
    layer7_outputs(3328) <= not a;
    layer7_outputs(3329) <= a xor b;
    layer7_outputs(3330) <= a;
    layer7_outputs(3331) <= a xor b;
    layer7_outputs(3332) <= not a;
    layer7_outputs(3333) <= '1';
    layer7_outputs(3334) <= a or b;
    layer7_outputs(3335) <= not a or b;
    layer7_outputs(3336) <= a;
    layer7_outputs(3337) <= a xor b;
    layer7_outputs(3338) <= a and b;
    layer7_outputs(3339) <= b;
    layer7_outputs(3340) <= b;
    layer7_outputs(3341) <= b;
    layer7_outputs(3342) <= not (a and b);
    layer7_outputs(3343) <= a and b;
    layer7_outputs(3344) <= not b;
    layer7_outputs(3345) <= a xor b;
    layer7_outputs(3346) <= b and not a;
    layer7_outputs(3347) <= not a;
    layer7_outputs(3348) <= not (a and b);
    layer7_outputs(3349) <= not b;
    layer7_outputs(3350) <= not a or b;
    layer7_outputs(3351) <= not (a or b);
    layer7_outputs(3352) <= not b;
    layer7_outputs(3353) <= not a;
    layer7_outputs(3354) <= b and not a;
    layer7_outputs(3355) <= a;
    layer7_outputs(3356) <= not b;
    layer7_outputs(3357) <= not b or a;
    layer7_outputs(3358) <= a and b;
    layer7_outputs(3359) <= not a;
    layer7_outputs(3360) <= a and not b;
    layer7_outputs(3361) <= a;
    layer7_outputs(3362) <= b;
    layer7_outputs(3363) <= a xor b;
    layer7_outputs(3364) <= not b;
    layer7_outputs(3365) <= not b;
    layer7_outputs(3366) <= not a;
    layer7_outputs(3367) <= not a;
    layer7_outputs(3368) <= a or b;
    layer7_outputs(3369) <= a and not b;
    layer7_outputs(3370) <= a xor b;
    layer7_outputs(3371) <= b and not a;
    layer7_outputs(3372) <= a;
    layer7_outputs(3373) <= not b or a;
    layer7_outputs(3374) <= a and b;
    layer7_outputs(3375) <= b;
    layer7_outputs(3376) <= a;
    layer7_outputs(3377) <= b;
    layer7_outputs(3378) <= not b;
    layer7_outputs(3379) <= a;
    layer7_outputs(3380) <= not (a or b);
    layer7_outputs(3381) <= not b;
    layer7_outputs(3382) <= a;
    layer7_outputs(3383) <= b;
    layer7_outputs(3384) <= b;
    layer7_outputs(3385) <= not (a or b);
    layer7_outputs(3386) <= a;
    layer7_outputs(3387) <= a and b;
    layer7_outputs(3388) <= a;
    layer7_outputs(3389) <= a xor b;
    layer7_outputs(3390) <= a;
    layer7_outputs(3391) <= not (a and b);
    layer7_outputs(3392) <= not (a and b);
    layer7_outputs(3393) <= not b;
    layer7_outputs(3394) <= a;
    layer7_outputs(3395) <= not (a or b);
    layer7_outputs(3396) <= not b;
    layer7_outputs(3397) <= not a or b;
    layer7_outputs(3398) <= b;
    layer7_outputs(3399) <= not b;
    layer7_outputs(3400) <= not b;
    layer7_outputs(3401) <= a;
    layer7_outputs(3402) <= not b;
    layer7_outputs(3403) <= not b or a;
    layer7_outputs(3404) <= not a;
    layer7_outputs(3405) <= a and not b;
    layer7_outputs(3406) <= a and b;
    layer7_outputs(3407) <= a;
    layer7_outputs(3408) <= b and not a;
    layer7_outputs(3409) <= not (a or b);
    layer7_outputs(3410) <= a and b;
    layer7_outputs(3411) <= a;
    layer7_outputs(3412) <= a xor b;
    layer7_outputs(3413) <= a and b;
    layer7_outputs(3414) <= not a;
    layer7_outputs(3415) <= '1';
    layer7_outputs(3416) <= b;
    layer7_outputs(3417) <= a and b;
    layer7_outputs(3418) <= a;
    layer7_outputs(3419) <= a;
    layer7_outputs(3420) <= b;
    layer7_outputs(3421) <= not (a and b);
    layer7_outputs(3422) <= not b;
    layer7_outputs(3423) <= a and not b;
    layer7_outputs(3424) <= not a;
    layer7_outputs(3425) <= b;
    layer7_outputs(3426) <= not b;
    layer7_outputs(3427) <= b and not a;
    layer7_outputs(3428) <= not a or b;
    layer7_outputs(3429) <= b and not a;
    layer7_outputs(3430) <= a xor b;
    layer7_outputs(3431) <= not b;
    layer7_outputs(3432) <= not a;
    layer7_outputs(3433) <= not a;
    layer7_outputs(3434) <= b;
    layer7_outputs(3435) <= not a or b;
    layer7_outputs(3436) <= not (a and b);
    layer7_outputs(3437) <= a;
    layer7_outputs(3438) <= a;
    layer7_outputs(3439) <= b and not a;
    layer7_outputs(3440) <= a xor b;
    layer7_outputs(3441) <= a and not b;
    layer7_outputs(3442) <= a xor b;
    layer7_outputs(3443) <= a and not b;
    layer7_outputs(3444) <= not a or b;
    layer7_outputs(3445) <= a;
    layer7_outputs(3446) <= not (a xor b);
    layer7_outputs(3447) <= b;
    layer7_outputs(3448) <= not (a or b);
    layer7_outputs(3449) <= not a or b;
    layer7_outputs(3450) <= a;
    layer7_outputs(3451) <= not a;
    layer7_outputs(3452) <= a xor b;
    layer7_outputs(3453) <= not (a or b);
    layer7_outputs(3454) <= not b;
    layer7_outputs(3455) <= a;
    layer7_outputs(3456) <= b and not a;
    layer7_outputs(3457) <= not (a xor b);
    layer7_outputs(3458) <= a;
    layer7_outputs(3459) <= not b or a;
    layer7_outputs(3460) <= not a;
    layer7_outputs(3461) <= not b;
    layer7_outputs(3462) <= not (a and b);
    layer7_outputs(3463) <= b;
    layer7_outputs(3464) <= '0';
    layer7_outputs(3465) <= b;
    layer7_outputs(3466) <= not (a and b);
    layer7_outputs(3467) <= a;
    layer7_outputs(3468) <= b;
    layer7_outputs(3469) <= not a or b;
    layer7_outputs(3470) <= not (a xor b);
    layer7_outputs(3471) <= a;
    layer7_outputs(3472) <= a or b;
    layer7_outputs(3473) <= a and b;
    layer7_outputs(3474) <= not (a or b);
    layer7_outputs(3475) <= a;
    layer7_outputs(3476) <= not a or b;
    layer7_outputs(3477) <= not b;
    layer7_outputs(3478) <= a;
    layer7_outputs(3479) <= not b;
    layer7_outputs(3480) <= not (a or b);
    layer7_outputs(3481) <= not a;
    layer7_outputs(3482) <= not a;
    layer7_outputs(3483) <= a xor b;
    layer7_outputs(3484) <= not (a xor b);
    layer7_outputs(3485) <= b and not a;
    layer7_outputs(3486) <= a or b;
    layer7_outputs(3487) <= not (a and b);
    layer7_outputs(3488) <= a;
    layer7_outputs(3489) <= a;
    layer7_outputs(3490) <= not (a xor b);
    layer7_outputs(3491) <= a xor b;
    layer7_outputs(3492) <= a xor b;
    layer7_outputs(3493) <= b and not a;
    layer7_outputs(3494) <= a xor b;
    layer7_outputs(3495) <= not (a xor b);
    layer7_outputs(3496) <= b and not a;
    layer7_outputs(3497) <= not a;
    layer7_outputs(3498) <= not (a and b);
    layer7_outputs(3499) <= not (a and b);
    layer7_outputs(3500) <= a xor b;
    layer7_outputs(3501) <= b and not a;
    layer7_outputs(3502) <= not (a xor b);
    layer7_outputs(3503) <= not (a xor b);
    layer7_outputs(3504) <= a and not b;
    layer7_outputs(3505) <= not a or b;
    layer7_outputs(3506) <= a and not b;
    layer7_outputs(3507) <= b;
    layer7_outputs(3508) <= not a;
    layer7_outputs(3509) <= a xor b;
    layer7_outputs(3510) <= not a or b;
    layer7_outputs(3511) <= a xor b;
    layer7_outputs(3512) <= not (a xor b);
    layer7_outputs(3513) <= '0';
    layer7_outputs(3514) <= a xor b;
    layer7_outputs(3515) <= not (a xor b);
    layer7_outputs(3516) <= not b;
    layer7_outputs(3517) <= b;
    layer7_outputs(3518) <= a;
    layer7_outputs(3519) <= b and not a;
    layer7_outputs(3520) <= not (a and b);
    layer7_outputs(3521) <= b and not a;
    layer7_outputs(3522) <= not (a xor b);
    layer7_outputs(3523) <= a;
    layer7_outputs(3524) <= b;
    layer7_outputs(3525) <= a;
    layer7_outputs(3526) <= b and not a;
    layer7_outputs(3527) <= not (a and b);
    layer7_outputs(3528) <= not b;
    layer7_outputs(3529) <= a;
    layer7_outputs(3530) <= not a;
    layer7_outputs(3531) <= not (a or b);
    layer7_outputs(3532) <= '1';
    layer7_outputs(3533) <= b;
    layer7_outputs(3534) <= a or b;
    layer7_outputs(3535) <= b;
    layer7_outputs(3536) <= not (a xor b);
    layer7_outputs(3537) <= not a;
    layer7_outputs(3538) <= a and not b;
    layer7_outputs(3539) <= b and not a;
    layer7_outputs(3540) <= not (a and b);
    layer7_outputs(3541) <= b;
    layer7_outputs(3542) <= a and not b;
    layer7_outputs(3543) <= a and b;
    layer7_outputs(3544) <= a;
    layer7_outputs(3545) <= b and not a;
    layer7_outputs(3546) <= a;
    layer7_outputs(3547) <= b and not a;
    layer7_outputs(3548) <= not a or b;
    layer7_outputs(3549) <= not b or a;
    layer7_outputs(3550) <= not a;
    layer7_outputs(3551) <= not (a or b);
    layer7_outputs(3552) <= not b or a;
    layer7_outputs(3553) <= not b;
    layer7_outputs(3554) <= '1';
    layer7_outputs(3555) <= b;
    layer7_outputs(3556) <= not b or a;
    layer7_outputs(3557) <= not b;
    layer7_outputs(3558) <= a;
    layer7_outputs(3559) <= not (a and b);
    layer7_outputs(3560) <= a xor b;
    layer7_outputs(3561) <= not (a xor b);
    layer7_outputs(3562) <= b;
    layer7_outputs(3563) <= not a;
    layer7_outputs(3564) <= b;
    layer7_outputs(3565) <= b and not a;
    layer7_outputs(3566) <= not b or a;
    layer7_outputs(3567) <= not a;
    layer7_outputs(3568) <= not (a and b);
    layer7_outputs(3569) <= b and not a;
    layer7_outputs(3570) <= not (a xor b);
    layer7_outputs(3571) <= a and b;
    layer7_outputs(3572) <= a and not b;
    layer7_outputs(3573) <= a;
    layer7_outputs(3574) <= not b;
    layer7_outputs(3575) <= a;
    layer7_outputs(3576) <= not b or a;
    layer7_outputs(3577) <= b;
    layer7_outputs(3578) <= not a;
    layer7_outputs(3579) <= not (a or b);
    layer7_outputs(3580) <= not (a xor b);
    layer7_outputs(3581) <= b;
    layer7_outputs(3582) <= b;
    layer7_outputs(3583) <= not (a or b);
    layer7_outputs(3584) <= a and b;
    layer7_outputs(3585) <= not b;
    layer7_outputs(3586) <= a;
    layer7_outputs(3587) <= not a or b;
    layer7_outputs(3588) <= b and not a;
    layer7_outputs(3589) <= not a;
    layer7_outputs(3590) <= a and b;
    layer7_outputs(3591) <= not (a xor b);
    layer7_outputs(3592) <= not b;
    layer7_outputs(3593) <= b;
    layer7_outputs(3594) <= not b;
    layer7_outputs(3595) <= not a;
    layer7_outputs(3596) <= not b;
    layer7_outputs(3597) <= a and b;
    layer7_outputs(3598) <= not a;
    layer7_outputs(3599) <= not (a or b);
    layer7_outputs(3600) <= not b;
    layer7_outputs(3601) <= not a or b;
    layer7_outputs(3602) <= not (a or b);
    layer7_outputs(3603) <= not a;
    layer7_outputs(3604) <= not a;
    layer7_outputs(3605) <= b and not a;
    layer7_outputs(3606) <= not a;
    layer7_outputs(3607) <= a;
    layer7_outputs(3608) <= a xor b;
    layer7_outputs(3609) <= not b;
    layer7_outputs(3610) <= a or b;
    layer7_outputs(3611) <= a or b;
    layer7_outputs(3612) <= not b;
    layer7_outputs(3613) <= b and not a;
    layer7_outputs(3614) <= a;
    layer7_outputs(3615) <= not a;
    layer7_outputs(3616) <= not b;
    layer7_outputs(3617) <= a and b;
    layer7_outputs(3618) <= not a;
    layer7_outputs(3619) <= a;
    layer7_outputs(3620) <= not (a and b);
    layer7_outputs(3621) <= a;
    layer7_outputs(3622) <= not b;
    layer7_outputs(3623) <= not a;
    layer7_outputs(3624) <= not (a xor b);
    layer7_outputs(3625) <= not (a and b);
    layer7_outputs(3626) <= a;
    layer7_outputs(3627) <= a and not b;
    layer7_outputs(3628) <= b;
    layer7_outputs(3629) <= a;
    layer7_outputs(3630) <= not (a xor b);
    layer7_outputs(3631) <= a xor b;
    layer7_outputs(3632) <= not a;
    layer7_outputs(3633) <= a or b;
    layer7_outputs(3634) <= not (a xor b);
    layer7_outputs(3635) <= a xor b;
    layer7_outputs(3636) <= not a or b;
    layer7_outputs(3637) <= a;
    layer7_outputs(3638) <= not a;
    layer7_outputs(3639) <= b;
    layer7_outputs(3640) <= not a or b;
    layer7_outputs(3641) <= a;
    layer7_outputs(3642) <= b;
    layer7_outputs(3643) <= a;
    layer7_outputs(3644) <= a or b;
    layer7_outputs(3645) <= a xor b;
    layer7_outputs(3646) <= a and b;
    layer7_outputs(3647) <= not a or b;
    layer7_outputs(3648) <= not a or b;
    layer7_outputs(3649) <= not b or a;
    layer7_outputs(3650) <= not (a xor b);
    layer7_outputs(3651) <= not a or b;
    layer7_outputs(3652) <= a and not b;
    layer7_outputs(3653) <= not b or a;
    layer7_outputs(3654) <= b;
    layer7_outputs(3655) <= a and b;
    layer7_outputs(3656) <= not (a or b);
    layer7_outputs(3657) <= b;
    layer7_outputs(3658) <= not b;
    layer7_outputs(3659) <= not b or a;
    layer7_outputs(3660) <= b;
    layer7_outputs(3661) <= a;
    layer7_outputs(3662) <= not a or b;
    layer7_outputs(3663) <= a or b;
    layer7_outputs(3664) <= not (a or b);
    layer7_outputs(3665) <= a or b;
    layer7_outputs(3666) <= not (a or b);
    layer7_outputs(3667) <= a xor b;
    layer7_outputs(3668) <= not b or a;
    layer7_outputs(3669) <= b;
    layer7_outputs(3670) <= a or b;
    layer7_outputs(3671) <= a and not b;
    layer7_outputs(3672) <= not a;
    layer7_outputs(3673) <= a;
    layer7_outputs(3674) <= a;
    layer7_outputs(3675) <= a xor b;
    layer7_outputs(3676) <= a xor b;
    layer7_outputs(3677) <= a;
    layer7_outputs(3678) <= not a;
    layer7_outputs(3679) <= '0';
    layer7_outputs(3680) <= a or b;
    layer7_outputs(3681) <= not b;
    layer7_outputs(3682) <= not (a xor b);
    layer7_outputs(3683) <= not a or b;
    layer7_outputs(3684) <= a and b;
    layer7_outputs(3685) <= b;
    layer7_outputs(3686) <= a;
    layer7_outputs(3687) <= not b;
    layer7_outputs(3688) <= '1';
    layer7_outputs(3689) <= not (a xor b);
    layer7_outputs(3690) <= not (a or b);
    layer7_outputs(3691) <= not b;
    layer7_outputs(3692) <= b;
    layer7_outputs(3693) <= not b;
    layer7_outputs(3694) <= a and b;
    layer7_outputs(3695) <= a;
    layer7_outputs(3696) <= not (a or b);
    layer7_outputs(3697) <= a and not b;
    layer7_outputs(3698) <= not b;
    layer7_outputs(3699) <= a xor b;
    layer7_outputs(3700) <= not b;
    layer7_outputs(3701) <= not b;
    layer7_outputs(3702) <= a;
    layer7_outputs(3703) <= a and b;
    layer7_outputs(3704) <= not (a and b);
    layer7_outputs(3705) <= '0';
    layer7_outputs(3706) <= b and not a;
    layer7_outputs(3707) <= not b;
    layer7_outputs(3708) <= a or b;
    layer7_outputs(3709) <= not a or b;
    layer7_outputs(3710) <= a and not b;
    layer7_outputs(3711) <= b and not a;
    layer7_outputs(3712) <= a or b;
    layer7_outputs(3713) <= a or b;
    layer7_outputs(3714) <= not b;
    layer7_outputs(3715) <= not b;
    layer7_outputs(3716) <= a xor b;
    layer7_outputs(3717) <= not a;
    layer7_outputs(3718) <= not a;
    layer7_outputs(3719) <= not a;
    layer7_outputs(3720) <= not b;
    layer7_outputs(3721) <= not b or a;
    layer7_outputs(3722) <= not a or b;
    layer7_outputs(3723) <= a and not b;
    layer7_outputs(3724) <= a and not b;
    layer7_outputs(3725) <= '1';
    layer7_outputs(3726) <= not a;
    layer7_outputs(3727) <= a and b;
    layer7_outputs(3728) <= a or b;
    layer7_outputs(3729) <= a;
    layer7_outputs(3730) <= not a;
    layer7_outputs(3731) <= not a or b;
    layer7_outputs(3732) <= not a;
    layer7_outputs(3733) <= not b;
    layer7_outputs(3734) <= a;
    layer7_outputs(3735) <= a and b;
    layer7_outputs(3736) <= not a or b;
    layer7_outputs(3737) <= a;
    layer7_outputs(3738) <= not a;
    layer7_outputs(3739) <= not b;
    layer7_outputs(3740) <= not a;
    layer7_outputs(3741) <= a xor b;
    layer7_outputs(3742) <= b;
    layer7_outputs(3743) <= not (a or b);
    layer7_outputs(3744) <= not b or a;
    layer7_outputs(3745) <= not a or b;
    layer7_outputs(3746) <= not b;
    layer7_outputs(3747) <= b;
    layer7_outputs(3748) <= a;
    layer7_outputs(3749) <= b;
    layer7_outputs(3750) <= not a;
    layer7_outputs(3751) <= a or b;
    layer7_outputs(3752) <= '1';
    layer7_outputs(3753) <= a and not b;
    layer7_outputs(3754) <= a and not b;
    layer7_outputs(3755) <= b;
    layer7_outputs(3756) <= a;
    layer7_outputs(3757) <= a and b;
    layer7_outputs(3758) <= a and not b;
    layer7_outputs(3759) <= not b or a;
    layer7_outputs(3760) <= b;
    layer7_outputs(3761) <= b;
    layer7_outputs(3762) <= b;
    layer7_outputs(3763) <= not b or a;
    layer7_outputs(3764) <= not b;
    layer7_outputs(3765) <= a and not b;
    layer7_outputs(3766) <= not (a and b);
    layer7_outputs(3767) <= not b;
    layer7_outputs(3768) <= not (a or b);
    layer7_outputs(3769) <= not a;
    layer7_outputs(3770) <= a xor b;
    layer7_outputs(3771) <= b;
    layer7_outputs(3772) <= not a;
    layer7_outputs(3773) <= a;
    layer7_outputs(3774) <= b;
    layer7_outputs(3775) <= not b or a;
    layer7_outputs(3776) <= not a;
    layer7_outputs(3777) <= not a;
    layer7_outputs(3778) <= b;
    layer7_outputs(3779) <= b;
    layer7_outputs(3780) <= a and not b;
    layer7_outputs(3781) <= not a;
    layer7_outputs(3782) <= b;
    layer7_outputs(3783) <= b;
    layer7_outputs(3784) <= not (a or b);
    layer7_outputs(3785) <= not b;
    layer7_outputs(3786) <= not (a or b);
    layer7_outputs(3787) <= a xor b;
    layer7_outputs(3788) <= a xor b;
    layer7_outputs(3789) <= not b or a;
    layer7_outputs(3790) <= not b;
    layer7_outputs(3791) <= a and b;
    layer7_outputs(3792) <= not b or a;
    layer7_outputs(3793) <= not b;
    layer7_outputs(3794) <= a;
    layer7_outputs(3795) <= a;
    layer7_outputs(3796) <= a;
    layer7_outputs(3797) <= not (a or b);
    layer7_outputs(3798) <= not a;
    layer7_outputs(3799) <= a xor b;
    layer7_outputs(3800) <= not a;
    layer7_outputs(3801) <= a and not b;
    layer7_outputs(3802) <= not (a and b);
    layer7_outputs(3803) <= a xor b;
    layer7_outputs(3804) <= not b or a;
    layer7_outputs(3805) <= not b;
    layer7_outputs(3806) <= not b;
    layer7_outputs(3807) <= a;
    layer7_outputs(3808) <= not (a or b);
    layer7_outputs(3809) <= a;
    layer7_outputs(3810) <= not a or b;
    layer7_outputs(3811) <= b and not a;
    layer7_outputs(3812) <= a;
    layer7_outputs(3813) <= not b or a;
    layer7_outputs(3814) <= '0';
    layer7_outputs(3815) <= a xor b;
    layer7_outputs(3816) <= not a;
    layer7_outputs(3817) <= a and not b;
    layer7_outputs(3818) <= a xor b;
    layer7_outputs(3819) <= a xor b;
    layer7_outputs(3820) <= not b;
    layer7_outputs(3821) <= b;
    layer7_outputs(3822) <= a and b;
    layer7_outputs(3823) <= a xor b;
    layer7_outputs(3824) <= not (a or b);
    layer7_outputs(3825) <= not b;
    layer7_outputs(3826) <= b and not a;
    layer7_outputs(3827) <= a xor b;
    layer7_outputs(3828) <= not b or a;
    layer7_outputs(3829) <= a;
    layer7_outputs(3830) <= b;
    layer7_outputs(3831) <= a;
    layer7_outputs(3832) <= not a or b;
    layer7_outputs(3833) <= a xor b;
    layer7_outputs(3834) <= not (a and b);
    layer7_outputs(3835) <= a or b;
    layer7_outputs(3836) <= '0';
    layer7_outputs(3837) <= a;
    layer7_outputs(3838) <= a;
    layer7_outputs(3839) <= a or b;
    layer7_outputs(3840) <= b;
    layer7_outputs(3841) <= not (a or b);
    layer7_outputs(3842) <= b;
    layer7_outputs(3843) <= not (a xor b);
    layer7_outputs(3844) <= a;
    layer7_outputs(3845) <= not a or b;
    layer7_outputs(3846) <= a or b;
    layer7_outputs(3847) <= b and not a;
    layer7_outputs(3848) <= a xor b;
    layer7_outputs(3849) <= not a;
    layer7_outputs(3850) <= not b or a;
    layer7_outputs(3851) <= not a;
    layer7_outputs(3852) <= a or b;
    layer7_outputs(3853) <= not (a or b);
    layer7_outputs(3854) <= a and b;
    layer7_outputs(3855) <= not a;
    layer7_outputs(3856) <= a;
    layer7_outputs(3857) <= a or b;
    layer7_outputs(3858) <= a;
    layer7_outputs(3859) <= b;
    layer7_outputs(3860) <= a;
    layer7_outputs(3861) <= b;
    layer7_outputs(3862) <= not b;
    layer7_outputs(3863) <= not b or a;
    layer7_outputs(3864) <= '0';
    layer7_outputs(3865) <= a or b;
    layer7_outputs(3866) <= b;
    layer7_outputs(3867) <= a;
    layer7_outputs(3868) <= not (a and b);
    layer7_outputs(3869) <= not (a and b);
    layer7_outputs(3870) <= not (a and b);
    layer7_outputs(3871) <= a and not b;
    layer7_outputs(3872) <= not a;
    layer7_outputs(3873) <= not a or b;
    layer7_outputs(3874) <= not b;
    layer7_outputs(3875) <= not b;
    layer7_outputs(3876) <= not b or a;
    layer7_outputs(3877) <= a;
    layer7_outputs(3878) <= b;
    layer7_outputs(3879) <= b;
    layer7_outputs(3880) <= not b;
    layer7_outputs(3881) <= b and not a;
    layer7_outputs(3882) <= not b or a;
    layer7_outputs(3883) <= not (a and b);
    layer7_outputs(3884) <= not a;
    layer7_outputs(3885) <= a;
    layer7_outputs(3886) <= not (a xor b);
    layer7_outputs(3887) <= a;
    layer7_outputs(3888) <= a xor b;
    layer7_outputs(3889) <= a;
    layer7_outputs(3890) <= '0';
    layer7_outputs(3891) <= not (a xor b);
    layer7_outputs(3892) <= not b;
    layer7_outputs(3893) <= not a or b;
    layer7_outputs(3894) <= a or b;
    layer7_outputs(3895) <= not (a and b);
    layer7_outputs(3896) <= b;
    layer7_outputs(3897) <= b;
    layer7_outputs(3898) <= not b;
    layer7_outputs(3899) <= b;
    layer7_outputs(3900) <= not (a or b);
    layer7_outputs(3901) <= a xor b;
    layer7_outputs(3902) <= not a;
    layer7_outputs(3903) <= not a;
    layer7_outputs(3904) <= a and not b;
    layer7_outputs(3905) <= a or b;
    layer7_outputs(3906) <= not (a xor b);
    layer7_outputs(3907) <= not a or b;
    layer7_outputs(3908) <= a and not b;
    layer7_outputs(3909) <= a;
    layer7_outputs(3910) <= a or b;
    layer7_outputs(3911) <= a or b;
    layer7_outputs(3912) <= not b;
    layer7_outputs(3913) <= a;
    layer7_outputs(3914) <= b and not a;
    layer7_outputs(3915) <= a or b;
    layer7_outputs(3916) <= not b or a;
    layer7_outputs(3917) <= not (a and b);
    layer7_outputs(3918) <= not a;
    layer7_outputs(3919) <= a xor b;
    layer7_outputs(3920) <= not a;
    layer7_outputs(3921) <= a and not b;
    layer7_outputs(3922) <= a and not b;
    layer7_outputs(3923) <= not (a xor b);
    layer7_outputs(3924) <= '0';
    layer7_outputs(3925) <= not (a and b);
    layer7_outputs(3926) <= b and not a;
    layer7_outputs(3927) <= not b;
    layer7_outputs(3928) <= not a;
    layer7_outputs(3929) <= b and not a;
    layer7_outputs(3930) <= not a;
    layer7_outputs(3931) <= b and not a;
    layer7_outputs(3932) <= not a;
    layer7_outputs(3933) <= a;
    layer7_outputs(3934) <= a and not b;
    layer7_outputs(3935) <= not a;
    layer7_outputs(3936) <= not (a xor b);
    layer7_outputs(3937) <= a xor b;
    layer7_outputs(3938) <= not (a xor b);
    layer7_outputs(3939) <= b;
    layer7_outputs(3940) <= not a;
    layer7_outputs(3941) <= not b;
    layer7_outputs(3942) <= not b;
    layer7_outputs(3943) <= not b or a;
    layer7_outputs(3944) <= not (a and b);
    layer7_outputs(3945) <= a xor b;
    layer7_outputs(3946) <= not b;
    layer7_outputs(3947) <= not a;
    layer7_outputs(3948) <= not b;
    layer7_outputs(3949) <= a and not b;
    layer7_outputs(3950) <= not a;
    layer7_outputs(3951) <= a and b;
    layer7_outputs(3952) <= not a;
    layer7_outputs(3953) <= not b;
    layer7_outputs(3954) <= a xor b;
    layer7_outputs(3955) <= b;
    layer7_outputs(3956) <= a;
    layer7_outputs(3957) <= not (a and b);
    layer7_outputs(3958) <= not b or a;
    layer7_outputs(3959) <= not b;
    layer7_outputs(3960) <= not (a xor b);
    layer7_outputs(3961) <= a xor b;
    layer7_outputs(3962) <= b;
    layer7_outputs(3963) <= not (a or b);
    layer7_outputs(3964) <= a;
    layer7_outputs(3965) <= not (a xor b);
    layer7_outputs(3966) <= b and not a;
    layer7_outputs(3967) <= a and not b;
    layer7_outputs(3968) <= not (a xor b);
    layer7_outputs(3969) <= not b;
    layer7_outputs(3970) <= a and b;
    layer7_outputs(3971) <= not (a or b);
    layer7_outputs(3972) <= b;
    layer7_outputs(3973) <= b;
    layer7_outputs(3974) <= not b;
    layer7_outputs(3975) <= a;
    layer7_outputs(3976) <= a;
    layer7_outputs(3977) <= not (a or b);
    layer7_outputs(3978) <= not a or b;
    layer7_outputs(3979) <= a;
    layer7_outputs(3980) <= a and b;
    layer7_outputs(3981) <= not b;
    layer7_outputs(3982) <= not (a or b);
    layer7_outputs(3983) <= a;
    layer7_outputs(3984) <= not b;
    layer7_outputs(3985) <= not b or a;
    layer7_outputs(3986) <= not b;
    layer7_outputs(3987) <= b;
    layer7_outputs(3988) <= a and not b;
    layer7_outputs(3989) <= not (a xor b);
    layer7_outputs(3990) <= not (a xor b);
    layer7_outputs(3991) <= a xor b;
    layer7_outputs(3992) <= a;
    layer7_outputs(3993) <= not (a or b);
    layer7_outputs(3994) <= b;
    layer7_outputs(3995) <= '0';
    layer7_outputs(3996) <= not a;
    layer7_outputs(3997) <= not (a or b);
    layer7_outputs(3998) <= b;
    layer7_outputs(3999) <= not (a and b);
    layer7_outputs(4000) <= a;
    layer7_outputs(4001) <= not b;
    layer7_outputs(4002) <= b;
    layer7_outputs(4003) <= not b;
    layer7_outputs(4004) <= a;
    layer7_outputs(4005) <= b;
    layer7_outputs(4006) <= not (a xor b);
    layer7_outputs(4007) <= not b or a;
    layer7_outputs(4008) <= a or b;
    layer7_outputs(4009) <= a xor b;
    layer7_outputs(4010) <= a;
    layer7_outputs(4011) <= not a or b;
    layer7_outputs(4012) <= a xor b;
    layer7_outputs(4013) <= a and not b;
    layer7_outputs(4014) <= not (a or b);
    layer7_outputs(4015) <= a;
    layer7_outputs(4016) <= not (a xor b);
    layer7_outputs(4017) <= a or b;
    layer7_outputs(4018) <= b and not a;
    layer7_outputs(4019) <= not (a or b);
    layer7_outputs(4020) <= not (a xor b);
    layer7_outputs(4021) <= not b;
    layer7_outputs(4022) <= not (a xor b);
    layer7_outputs(4023) <= b;
    layer7_outputs(4024) <= not (a and b);
    layer7_outputs(4025) <= a;
    layer7_outputs(4026) <= a and not b;
    layer7_outputs(4027) <= not b;
    layer7_outputs(4028) <= a and b;
    layer7_outputs(4029) <= not a;
    layer7_outputs(4030) <= b and not a;
    layer7_outputs(4031) <= a;
    layer7_outputs(4032) <= b;
    layer7_outputs(4033) <= a and not b;
    layer7_outputs(4034) <= a;
    layer7_outputs(4035) <= a xor b;
    layer7_outputs(4036) <= not (a and b);
    layer7_outputs(4037) <= b;
    layer7_outputs(4038) <= a;
    layer7_outputs(4039) <= not (a xor b);
    layer7_outputs(4040) <= b and not a;
    layer7_outputs(4041) <= a xor b;
    layer7_outputs(4042) <= not b;
    layer7_outputs(4043) <= not a or b;
    layer7_outputs(4044) <= a and b;
    layer7_outputs(4045) <= b and not a;
    layer7_outputs(4046) <= b;
    layer7_outputs(4047) <= not (a and b);
    layer7_outputs(4048) <= a;
    layer7_outputs(4049) <= b and not a;
    layer7_outputs(4050) <= not (a or b);
    layer7_outputs(4051) <= a and not b;
    layer7_outputs(4052) <= not a or b;
    layer7_outputs(4053) <= not b or a;
    layer7_outputs(4054) <= b;
    layer7_outputs(4055) <= a xor b;
    layer7_outputs(4056) <= b;
    layer7_outputs(4057) <= a xor b;
    layer7_outputs(4058) <= not (a or b);
    layer7_outputs(4059) <= not b or a;
    layer7_outputs(4060) <= b;
    layer7_outputs(4061) <= not a or b;
    layer7_outputs(4062) <= a xor b;
    layer7_outputs(4063) <= a xor b;
    layer7_outputs(4064) <= a;
    layer7_outputs(4065) <= a xor b;
    layer7_outputs(4066) <= b;
    layer7_outputs(4067) <= b;
    layer7_outputs(4068) <= a and b;
    layer7_outputs(4069) <= not (a xor b);
    layer7_outputs(4070) <= a and b;
    layer7_outputs(4071) <= not (a xor b);
    layer7_outputs(4072) <= not a;
    layer7_outputs(4073) <= not a;
    layer7_outputs(4074) <= not b;
    layer7_outputs(4075) <= a and b;
    layer7_outputs(4076) <= not b or a;
    layer7_outputs(4077) <= b and not a;
    layer7_outputs(4078) <= '0';
    layer7_outputs(4079) <= a and b;
    layer7_outputs(4080) <= b and not a;
    layer7_outputs(4081) <= b;
    layer7_outputs(4082) <= not a;
    layer7_outputs(4083) <= not a or b;
    layer7_outputs(4084) <= not b or a;
    layer7_outputs(4085) <= not a;
    layer7_outputs(4086) <= a and b;
    layer7_outputs(4087) <= b and not a;
    layer7_outputs(4088) <= a;
    layer7_outputs(4089) <= not b;
    layer7_outputs(4090) <= not b;
    layer7_outputs(4091) <= not a;
    layer7_outputs(4092) <= a and b;
    layer7_outputs(4093) <= not a;
    layer7_outputs(4094) <= not a or b;
    layer7_outputs(4095) <= not b;
    layer7_outputs(4096) <= not b;
    layer7_outputs(4097) <= b and not a;
    layer7_outputs(4098) <= not (a xor b);
    layer7_outputs(4099) <= not (a or b);
    layer7_outputs(4100) <= not b or a;
    layer7_outputs(4101) <= b;
    layer7_outputs(4102) <= not b;
    layer7_outputs(4103) <= not b;
    layer7_outputs(4104) <= not b or a;
    layer7_outputs(4105) <= b;
    layer7_outputs(4106) <= a or b;
    layer7_outputs(4107) <= a;
    layer7_outputs(4108) <= b;
    layer7_outputs(4109) <= a;
    layer7_outputs(4110) <= a and b;
    layer7_outputs(4111) <= '0';
    layer7_outputs(4112) <= not b or a;
    layer7_outputs(4113) <= a and not b;
    layer7_outputs(4114) <= not b;
    layer7_outputs(4115) <= not b;
    layer7_outputs(4116) <= a;
    layer7_outputs(4117) <= not a or b;
    layer7_outputs(4118) <= not b;
    layer7_outputs(4119) <= a xor b;
    layer7_outputs(4120) <= not (a xor b);
    layer7_outputs(4121) <= a;
    layer7_outputs(4122) <= not a;
    layer7_outputs(4123) <= a or b;
    layer7_outputs(4124) <= not (a and b);
    layer7_outputs(4125) <= a xor b;
    layer7_outputs(4126) <= not (a and b);
    layer7_outputs(4127) <= not a;
    layer7_outputs(4128) <= b;
    layer7_outputs(4129) <= a;
    layer7_outputs(4130) <= not a or b;
    layer7_outputs(4131) <= a or b;
    layer7_outputs(4132) <= b;
    layer7_outputs(4133) <= '1';
    layer7_outputs(4134) <= a xor b;
    layer7_outputs(4135) <= not a;
    layer7_outputs(4136) <= '1';
    layer7_outputs(4137) <= not (a xor b);
    layer7_outputs(4138) <= not (a and b);
    layer7_outputs(4139) <= a xor b;
    layer7_outputs(4140) <= not a;
    layer7_outputs(4141) <= a xor b;
    layer7_outputs(4142) <= a xor b;
    layer7_outputs(4143) <= a xor b;
    layer7_outputs(4144) <= a;
    layer7_outputs(4145) <= not a;
    layer7_outputs(4146) <= not b;
    layer7_outputs(4147) <= b and not a;
    layer7_outputs(4148) <= not (a xor b);
    layer7_outputs(4149) <= not (a xor b);
    layer7_outputs(4150) <= a and not b;
    layer7_outputs(4151) <= b and not a;
    layer7_outputs(4152) <= a and not b;
    layer7_outputs(4153) <= not (a or b);
    layer7_outputs(4154) <= not a;
    layer7_outputs(4155) <= a and not b;
    layer7_outputs(4156) <= b;
    layer7_outputs(4157) <= not a;
    layer7_outputs(4158) <= not b or a;
    layer7_outputs(4159) <= b;
    layer7_outputs(4160) <= not (a and b);
    layer7_outputs(4161) <= b;
    layer7_outputs(4162) <= not b or a;
    layer7_outputs(4163) <= a xor b;
    layer7_outputs(4164) <= not (a xor b);
    layer7_outputs(4165) <= a xor b;
    layer7_outputs(4166) <= b;
    layer7_outputs(4167) <= a and not b;
    layer7_outputs(4168) <= a and b;
    layer7_outputs(4169) <= not (a xor b);
    layer7_outputs(4170) <= not (a xor b);
    layer7_outputs(4171) <= a xor b;
    layer7_outputs(4172) <= not (a xor b);
    layer7_outputs(4173) <= not a;
    layer7_outputs(4174) <= b;
    layer7_outputs(4175) <= a;
    layer7_outputs(4176) <= not a;
    layer7_outputs(4177) <= not a;
    layer7_outputs(4178) <= b;
    layer7_outputs(4179) <= b;
    layer7_outputs(4180) <= b;
    layer7_outputs(4181) <= not (a or b);
    layer7_outputs(4182) <= a and b;
    layer7_outputs(4183) <= not a;
    layer7_outputs(4184) <= not (a or b);
    layer7_outputs(4185) <= not a;
    layer7_outputs(4186) <= not a;
    layer7_outputs(4187) <= a xor b;
    layer7_outputs(4188) <= b;
    layer7_outputs(4189) <= not a;
    layer7_outputs(4190) <= not b;
    layer7_outputs(4191) <= not a;
    layer7_outputs(4192) <= a or b;
    layer7_outputs(4193) <= b;
    layer7_outputs(4194) <= a or b;
    layer7_outputs(4195) <= not (a and b);
    layer7_outputs(4196) <= a and not b;
    layer7_outputs(4197) <= not b;
    layer7_outputs(4198) <= not a or b;
    layer7_outputs(4199) <= not (a xor b);
    layer7_outputs(4200) <= not b or a;
    layer7_outputs(4201) <= not b or a;
    layer7_outputs(4202) <= a xor b;
    layer7_outputs(4203) <= a xor b;
    layer7_outputs(4204) <= a and not b;
    layer7_outputs(4205) <= a or b;
    layer7_outputs(4206) <= a xor b;
    layer7_outputs(4207) <= not b;
    layer7_outputs(4208) <= not a;
    layer7_outputs(4209) <= b and not a;
    layer7_outputs(4210) <= not b or a;
    layer7_outputs(4211) <= not (a and b);
    layer7_outputs(4212) <= not b;
    layer7_outputs(4213) <= b and not a;
    layer7_outputs(4214) <= not a;
    layer7_outputs(4215) <= not (a or b);
    layer7_outputs(4216) <= a;
    layer7_outputs(4217) <= b;
    layer7_outputs(4218) <= a and not b;
    layer7_outputs(4219) <= not b;
    layer7_outputs(4220) <= a xor b;
    layer7_outputs(4221) <= not a;
    layer7_outputs(4222) <= not b;
    layer7_outputs(4223) <= not a;
    layer7_outputs(4224) <= not (a and b);
    layer7_outputs(4225) <= not b;
    layer7_outputs(4226) <= not a;
    layer7_outputs(4227) <= b;
    layer7_outputs(4228) <= not (a xor b);
    layer7_outputs(4229) <= a and not b;
    layer7_outputs(4230) <= a and b;
    layer7_outputs(4231) <= a;
    layer7_outputs(4232) <= a xor b;
    layer7_outputs(4233) <= b;
    layer7_outputs(4234) <= not (a or b);
    layer7_outputs(4235) <= not a;
    layer7_outputs(4236) <= not b;
    layer7_outputs(4237) <= not (a xor b);
    layer7_outputs(4238) <= not b or a;
    layer7_outputs(4239) <= a xor b;
    layer7_outputs(4240) <= not (a or b);
    layer7_outputs(4241) <= not a;
    layer7_outputs(4242) <= not b;
    layer7_outputs(4243) <= a or b;
    layer7_outputs(4244) <= not (a and b);
    layer7_outputs(4245) <= b;
    layer7_outputs(4246) <= a xor b;
    layer7_outputs(4247) <= not a;
    layer7_outputs(4248) <= not a;
    layer7_outputs(4249) <= not (a xor b);
    layer7_outputs(4250) <= not (a xor b);
    layer7_outputs(4251) <= not b;
    layer7_outputs(4252) <= b and not a;
    layer7_outputs(4253) <= a;
    layer7_outputs(4254) <= a;
    layer7_outputs(4255) <= a;
    layer7_outputs(4256) <= a xor b;
    layer7_outputs(4257) <= not a;
    layer7_outputs(4258) <= not a;
    layer7_outputs(4259) <= a and b;
    layer7_outputs(4260) <= not a;
    layer7_outputs(4261) <= not a;
    layer7_outputs(4262) <= b and not a;
    layer7_outputs(4263) <= not (a xor b);
    layer7_outputs(4264) <= a and b;
    layer7_outputs(4265) <= not a;
    layer7_outputs(4266) <= not b;
    layer7_outputs(4267) <= not (a or b);
    layer7_outputs(4268) <= a xor b;
    layer7_outputs(4269) <= a or b;
    layer7_outputs(4270) <= a;
    layer7_outputs(4271) <= a;
    layer7_outputs(4272) <= not (a or b);
    layer7_outputs(4273) <= a;
    layer7_outputs(4274) <= b;
    layer7_outputs(4275) <= not b;
    layer7_outputs(4276) <= not a;
    layer7_outputs(4277) <= a;
    layer7_outputs(4278) <= not (a xor b);
    layer7_outputs(4279) <= not b or a;
    layer7_outputs(4280) <= not (a and b);
    layer7_outputs(4281) <= not (a xor b);
    layer7_outputs(4282) <= not a;
    layer7_outputs(4283) <= not a;
    layer7_outputs(4284) <= a;
    layer7_outputs(4285) <= a xor b;
    layer7_outputs(4286) <= not b;
    layer7_outputs(4287) <= a;
    layer7_outputs(4288) <= not b or a;
    layer7_outputs(4289) <= a;
    layer7_outputs(4290) <= b;
    layer7_outputs(4291) <= a;
    layer7_outputs(4292) <= a or b;
    layer7_outputs(4293) <= not a;
    layer7_outputs(4294) <= not b;
    layer7_outputs(4295) <= a xor b;
    layer7_outputs(4296) <= not b;
    layer7_outputs(4297) <= a;
    layer7_outputs(4298) <= b;
    layer7_outputs(4299) <= a and b;
    layer7_outputs(4300) <= not a or b;
    layer7_outputs(4301) <= not (a xor b);
    layer7_outputs(4302) <= not a;
    layer7_outputs(4303) <= not (a xor b);
    layer7_outputs(4304) <= not a;
    layer7_outputs(4305) <= '1';
    layer7_outputs(4306) <= a or b;
    layer7_outputs(4307) <= b and not a;
    layer7_outputs(4308) <= not b;
    layer7_outputs(4309) <= a;
    layer7_outputs(4310) <= not b or a;
    layer7_outputs(4311) <= not a;
    layer7_outputs(4312) <= a xor b;
    layer7_outputs(4313) <= a xor b;
    layer7_outputs(4314) <= a or b;
    layer7_outputs(4315) <= not b or a;
    layer7_outputs(4316) <= not b;
    layer7_outputs(4317) <= a and not b;
    layer7_outputs(4318) <= b;
    layer7_outputs(4319) <= not (a and b);
    layer7_outputs(4320) <= a;
    layer7_outputs(4321) <= a;
    layer7_outputs(4322) <= a or b;
    layer7_outputs(4323) <= a or b;
    layer7_outputs(4324) <= not b;
    layer7_outputs(4325) <= a xor b;
    layer7_outputs(4326) <= b and not a;
    layer7_outputs(4327) <= not b;
    layer7_outputs(4328) <= not b;
    layer7_outputs(4329) <= not a;
    layer7_outputs(4330) <= not a or b;
    layer7_outputs(4331) <= b;
    layer7_outputs(4332) <= a and not b;
    layer7_outputs(4333) <= not a;
    layer7_outputs(4334) <= not b;
    layer7_outputs(4335) <= not (a xor b);
    layer7_outputs(4336) <= not (a xor b);
    layer7_outputs(4337) <= not (a or b);
    layer7_outputs(4338) <= a and not b;
    layer7_outputs(4339) <= not b;
    layer7_outputs(4340) <= b;
    layer7_outputs(4341) <= a xor b;
    layer7_outputs(4342) <= b;
    layer7_outputs(4343) <= not (a or b);
    layer7_outputs(4344) <= a xor b;
    layer7_outputs(4345) <= b;
    layer7_outputs(4346) <= b and not a;
    layer7_outputs(4347) <= not a;
    layer7_outputs(4348) <= not (a and b);
    layer7_outputs(4349) <= not (a and b);
    layer7_outputs(4350) <= not b or a;
    layer7_outputs(4351) <= not a or b;
    layer7_outputs(4352) <= not b or a;
    layer7_outputs(4353) <= not (a and b);
    layer7_outputs(4354) <= b;
    layer7_outputs(4355) <= not a;
    layer7_outputs(4356) <= a;
    layer7_outputs(4357) <= a;
    layer7_outputs(4358) <= not b;
    layer7_outputs(4359) <= not b;
    layer7_outputs(4360) <= not b;
    layer7_outputs(4361) <= not b;
    layer7_outputs(4362) <= not a;
    layer7_outputs(4363) <= not (a or b);
    layer7_outputs(4364) <= a and not b;
    layer7_outputs(4365) <= a and b;
    layer7_outputs(4366) <= not (a and b);
    layer7_outputs(4367) <= not b;
    layer7_outputs(4368) <= not (a and b);
    layer7_outputs(4369) <= not (a or b);
    layer7_outputs(4370) <= not b;
    layer7_outputs(4371) <= a xor b;
    layer7_outputs(4372) <= not b or a;
    layer7_outputs(4373) <= not (a xor b);
    layer7_outputs(4374) <= b;
    layer7_outputs(4375) <= not a;
    layer7_outputs(4376) <= not a;
    layer7_outputs(4377) <= not (a or b);
    layer7_outputs(4378) <= not (a and b);
    layer7_outputs(4379) <= a or b;
    layer7_outputs(4380) <= b and not a;
    layer7_outputs(4381) <= not b or a;
    layer7_outputs(4382) <= not a;
    layer7_outputs(4383) <= not (a and b);
    layer7_outputs(4384) <= b;
    layer7_outputs(4385) <= not (a or b);
    layer7_outputs(4386) <= not a;
    layer7_outputs(4387) <= a and not b;
    layer7_outputs(4388) <= a and b;
    layer7_outputs(4389) <= not (a xor b);
    layer7_outputs(4390) <= a or b;
    layer7_outputs(4391) <= not (a xor b);
    layer7_outputs(4392) <= b;
    layer7_outputs(4393) <= not b;
    layer7_outputs(4394) <= a and b;
    layer7_outputs(4395) <= not a;
    layer7_outputs(4396) <= a or b;
    layer7_outputs(4397) <= not a or b;
    layer7_outputs(4398) <= not (a or b);
    layer7_outputs(4399) <= '1';
    layer7_outputs(4400) <= not (a and b);
    layer7_outputs(4401) <= not (a xor b);
    layer7_outputs(4402) <= '1';
    layer7_outputs(4403) <= a;
    layer7_outputs(4404) <= a xor b;
    layer7_outputs(4405) <= not b;
    layer7_outputs(4406) <= not b;
    layer7_outputs(4407) <= b and not a;
    layer7_outputs(4408) <= a xor b;
    layer7_outputs(4409) <= a or b;
    layer7_outputs(4410) <= not a or b;
    layer7_outputs(4411) <= not (a and b);
    layer7_outputs(4412) <= '0';
    layer7_outputs(4413) <= not a or b;
    layer7_outputs(4414) <= b and not a;
    layer7_outputs(4415) <= not (a or b);
    layer7_outputs(4416) <= not a or b;
    layer7_outputs(4417) <= b and not a;
    layer7_outputs(4418) <= a xor b;
    layer7_outputs(4419) <= '0';
    layer7_outputs(4420) <= a;
    layer7_outputs(4421) <= a;
    layer7_outputs(4422) <= a and not b;
    layer7_outputs(4423) <= not (a or b);
    layer7_outputs(4424) <= not b;
    layer7_outputs(4425) <= a;
    layer7_outputs(4426) <= a;
    layer7_outputs(4427) <= a;
    layer7_outputs(4428) <= not b;
    layer7_outputs(4429) <= not a;
    layer7_outputs(4430) <= a and b;
    layer7_outputs(4431) <= a;
    layer7_outputs(4432) <= b and not a;
    layer7_outputs(4433) <= not (a and b);
    layer7_outputs(4434) <= a or b;
    layer7_outputs(4435) <= not (a xor b);
    layer7_outputs(4436) <= not a;
    layer7_outputs(4437) <= b;
    layer7_outputs(4438) <= not (a or b);
    layer7_outputs(4439) <= not a;
    layer7_outputs(4440) <= not b;
    layer7_outputs(4441) <= a;
    layer7_outputs(4442) <= b and not a;
    layer7_outputs(4443) <= not (a or b);
    layer7_outputs(4444) <= b;
    layer7_outputs(4445) <= not b;
    layer7_outputs(4446) <= not b or a;
    layer7_outputs(4447) <= not b;
    layer7_outputs(4448) <= b and not a;
    layer7_outputs(4449) <= not (a or b);
    layer7_outputs(4450) <= b;
    layer7_outputs(4451) <= not b or a;
    layer7_outputs(4452) <= a;
    layer7_outputs(4453) <= b;
    layer7_outputs(4454) <= a xor b;
    layer7_outputs(4455) <= not (a or b);
    layer7_outputs(4456) <= a and b;
    layer7_outputs(4457) <= b and not a;
    layer7_outputs(4458) <= not (a xor b);
    layer7_outputs(4459) <= '1';
    layer7_outputs(4460) <= b;
    layer7_outputs(4461) <= not (a or b);
    layer7_outputs(4462) <= a and b;
    layer7_outputs(4463) <= b;
    layer7_outputs(4464) <= not (a and b);
    layer7_outputs(4465) <= a or b;
    layer7_outputs(4466) <= a or b;
    layer7_outputs(4467) <= a;
    layer7_outputs(4468) <= b;
    layer7_outputs(4469) <= not a or b;
    layer7_outputs(4470) <= not b;
    layer7_outputs(4471) <= not b or a;
    layer7_outputs(4472) <= not a;
    layer7_outputs(4473) <= not a;
    layer7_outputs(4474) <= a;
    layer7_outputs(4475) <= not (a xor b);
    layer7_outputs(4476) <= not a or b;
    layer7_outputs(4477) <= a;
    layer7_outputs(4478) <= not a or b;
    layer7_outputs(4479) <= b and not a;
    layer7_outputs(4480) <= b and not a;
    layer7_outputs(4481) <= not b or a;
    layer7_outputs(4482) <= not b;
    layer7_outputs(4483) <= not (a xor b);
    layer7_outputs(4484) <= not a;
    layer7_outputs(4485) <= a and b;
    layer7_outputs(4486) <= a;
    layer7_outputs(4487) <= not b;
    layer7_outputs(4488) <= not a;
    layer7_outputs(4489) <= not b;
    layer7_outputs(4490) <= b;
    layer7_outputs(4491) <= a and not b;
    layer7_outputs(4492) <= a xor b;
    layer7_outputs(4493) <= not (a and b);
    layer7_outputs(4494) <= not b or a;
    layer7_outputs(4495) <= not a;
    layer7_outputs(4496) <= not a or b;
    layer7_outputs(4497) <= not b;
    layer7_outputs(4498) <= a xor b;
    layer7_outputs(4499) <= not a;
    layer7_outputs(4500) <= a;
    layer7_outputs(4501) <= not a;
    layer7_outputs(4502) <= not a;
    layer7_outputs(4503) <= not b or a;
    layer7_outputs(4504) <= a or b;
    layer7_outputs(4505) <= a or b;
    layer7_outputs(4506) <= b and not a;
    layer7_outputs(4507) <= a;
    layer7_outputs(4508) <= not (a and b);
    layer7_outputs(4509) <= a and not b;
    layer7_outputs(4510) <= not (a xor b);
    layer7_outputs(4511) <= not (a or b);
    layer7_outputs(4512) <= a and not b;
    layer7_outputs(4513) <= a;
    layer7_outputs(4514) <= a xor b;
    layer7_outputs(4515) <= not (a or b);
    layer7_outputs(4516) <= b;
    layer7_outputs(4517) <= b;
    layer7_outputs(4518) <= b;
    layer7_outputs(4519) <= a and b;
    layer7_outputs(4520) <= not b;
    layer7_outputs(4521) <= b and not a;
    layer7_outputs(4522) <= not a or b;
    layer7_outputs(4523) <= a;
    layer7_outputs(4524) <= a or b;
    layer7_outputs(4525) <= b and not a;
    layer7_outputs(4526) <= not (a and b);
    layer7_outputs(4527) <= a and not b;
    layer7_outputs(4528) <= not b;
    layer7_outputs(4529) <= not (a xor b);
    layer7_outputs(4530) <= a xor b;
    layer7_outputs(4531) <= a and not b;
    layer7_outputs(4532) <= not b or a;
    layer7_outputs(4533) <= not a;
    layer7_outputs(4534) <= a and not b;
    layer7_outputs(4535) <= not a;
    layer7_outputs(4536) <= not (a xor b);
    layer7_outputs(4537) <= not a or b;
    layer7_outputs(4538) <= not b or a;
    layer7_outputs(4539) <= not a or b;
    layer7_outputs(4540) <= b and not a;
    layer7_outputs(4541) <= not b;
    layer7_outputs(4542) <= not (a and b);
    layer7_outputs(4543) <= not (a and b);
    layer7_outputs(4544) <= not b;
    layer7_outputs(4545) <= a;
    layer7_outputs(4546) <= a and not b;
    layer7_outputs(4547) <= not b or a;
    layer7_outputs(4548) <= a;
    layer7_outputs(4549) <= not (a and b);
    layer7_outputs(4550) <= not (a xor b);
    layer7_outputs(4551) <= b;
    layer7_outputs(4552) <= b;
    layer7_outputs(4553) <= b;
    layer7_outputs(4554) <= not b;
    layer7_outputs(4555) <= b;
    layer7_outputs(4556) <= a xor b;
    layer7_outputs(4557) <= b and not a;
    layer7_outputs(4558) <= a;
    layer7_outputs(4559) <= not (a or b);
    layer7_outputs(4560) <= not b;
    layer7_outputs(4561) <= not (a xor b);
    layer7_outputs(4562) <= b and not a;
    layer7_outputs(4563) <= not a;
    layer7_outputs(4564) <= a;
    layer7_outputs(4565) <= b and not a;
    layer7_outputs(4566) <= not a or b;
    layer7_outputs(4567) <= b and not a;
    layer7_outputs(4568) <= not b;
    layer7_outputs(4569) <= not b;
    layer7_outputs(4570) <= not a;
    layer7_outputs(4571) <= a;
    layer7_outputs(4572) <= b;
    layer7_outputs(4573) <= not a;
    layer7_outputs(4574) <= not b;
    layer7_outputs(4575) <= not a or b;
    layer7_outputs(4576) <= b;
    layer7_outputs(4577) <= a or b;
    layer7_outputs(4578) <= b;
    layer7_outputs(4579) <= not (a or b);
    layer7_outputs(4580) <= a;
    layer7_outputs(4581) <= b and not a;
    layer7_outputs(4582) <= not a or b;
    layer7_outputs(4583) <= not a or b;
    layer7_outputs(4584) <= a xor b;
    layer7_outputs(4585) <= not b;
    layer7_outputs(4586) <= a xor b;
    layer7_outputs(4587) <= a xor b;
    layer7_outputs(4588) <= not b;
    layer7_outputs(4589) <= a xor b;
    layer7_outputs(4590) <= a;
    layer7_outputs(4591) <= not b;
    layer7_outputs(4592) <= not b;
    layer7_outputs(4593) <= not (a or b);
    layer7_outputs(4594) <= not b;
    layer7_outputs(4595) <= a or b;
    layer7_outputs(4596) <= a or b;
    layer7_outputs(4597) <= a xor b;
    layer7_outputs(4598) <= not a;
    layer7_outputs(4599) <= not (a xor b);
    layer7_outputs(4600) <= not (a xor b);
    layer7_outputs(4601) <= b;
    layer7_outputs(4602) <= not b;
    layer7_outputs(4603) <= not b or a;
    layer7_outputs(4604) <= b;
    layer7_outputs(4605) <= not (a xor b);
    layer7_outputs(4606) <= not a;
    layer7_outputs(4607) <= not b or a;
    layer7_outputs(4608) <= '1';
    layer7_outputs(4609) <= not b or a;
    layer7_outputs(4610) <= a xor b;
    layer7_outputs(4611) <= not (a xor b);
    layer7_outputs(4612) <= not (a or b);
    layer7_outputs(4613) <= not (a and b);
    layer7_outputs(4614) <= b;
    layer7_outputs(4615) <= not (a xor b);
    layer7_outputs(4616) <= '0';
    layer7_outputs(4617) <= not b or a;
    layer7_outputs(4618) <= b;
    layer7_outputs(4619) <= a and not b;
    layer7_outputs(4620) <= not b;
    layer7_outputs(4621) <= not (a xor b);
    layer7_outputs(4622) <= a;
    layer7_outputs(4623) <= not b;
    layer7_outputs(4624) <= not (a and b);
    layer7_outputs(4625) <= a and not b;
    layer7_outputs(4626) <= a or b;
    layer7_outputs(4627) <= not b;
    layer7_outputs(4628) <= '0';
    layer7_outputs(4629) <= not (a and b);
    layer7_outputs(4630) <= a xor b;
    layer7_outputs(4631) <= not b;
    layer7_outputs(4632) <= a;
    layer7_outputs(4633) <= not (a and b);
    layer7_outputs(4634) <= b and not a;
    layer7_outputs(4635) <= not b or a;
    layer7_outputs(4636) <= a;
    layer7_outputs(4637) <= a and not b;
    layer7_outputs(4638) <= b;
    layer7_outputs(4639) <= not a;
    layer7_outputs(4640) <= not b;
    layer7_outputs(4641) <= a;
    layer7_outputs(4642) <= not (a xor b);
    layer7_outputs(4643) <= a xor b;
    layer7_outputs(4644) <= b and not a;
    layer7_outputs(4645) <= b;
    layer7_outputs(4646) <= b;
    layer7_outputs(4647) <= not b;
    layer7_outputs(4648) <= not b;
    layer7_outputs(4649) <= not a or b;
    layer7_outputs(4650) <= not a;
    layer7_outputs(4651) <= a;
    layer7_outputs(4652) <= a xor b;
    layer7_outputs(4653) <= a;
    layer7_outputs(4654) <= b and not a;
    layer7_outputs(4655) <= not b or a;
    layer7_outputs(4656) <= b and not a;
    layer7_outputs(4657) <= a or b;
    layer7_outputs(4658) <= a or b;
    layer7_outputs(4659) <= not b;
    layer7_outputs(4660) <= not a;
    layer7_outputs(4661) <= not b or a;
    layer7_outputs(4662) <= a and b;
    layer7_outputs(4663) <= not a or b;
    layer7_outputs(4664) <= not b;
    layer7_outputs(4665) <= a;
    layer7_outputs(4666) <= not a;
    layer7_outputs(4667) <= not b;
    layer7_outputs(4668) <= b and not a;
    layer7_outputs(4669) <= a or b;
    layer7_outputs(4670) <= b;
    layer7_outputs(4671) <= a xor b;
    layer7_outputs(4672) <= not a;
    layer7_outputs(4673) <= b and not a;
    layer7_outputs(4674) <= not a or b;
    layer7_outputs(4675) <= a or b;
    layer7_outputs(4676) <= not a;
    layer7_outputs(4677) <= b and not a;
    layer7_outputs(4678) <= a xor b;
    layer7_outputs(4679) <= a and b;
    layer7_outputs(4680) <= a;
    layer7_outputs(4681) <= a or b;
    layer7_outputs(4682) <= not (a xor b);
    layer7_outputs(4683) <= a;
    layer7_outputs(4684) <= not (a xor b);
    layer7_outputs(4685) <= not (a or b);
    layer7_outputs(4686) <= not b;
    layer7_outputs(4687) <= a;
    layer7_outputs(4688) <= not b;
    layer7_outputs(4689) <= not a;
    layer7_outputs(4690) <= a;
    layer7_outputs(4691) <= a xor b;
    layer7_outputs(4692) <= not (a or b);
    layer7_outputs(4693) <= not a;
    layer7_outputs(4694) <= b;
    layer7_outputs(4695) <= not b or a;
    layer7_outputs(4696) <= not b;
    layer7_outputs(4697) <= '1';
    layer7_outputs(4698) <= b and not a;
    layer7_outputs(4699) <= b and not a;
    layer7_outputs(4700) <= b;
    layer7_outputs(4701) <= a and not b;
    layer7_outputs(4702) <= a;
    layer7_outputs(4703) <= b;
    layer7_outputs(4704) <= a;
    layer7_outputs(4705) <= not b;
    layer7_outputs(4706) <= not b;
    layer7_outputs(4707) <= b;
    layer7_outputs(4708) <= not a;
    layer7_outputs(4709) <= a;
    layer7_outputs(4710) <= a or b;
    layer7_outputs(4711) <= not (a xor b);
    layer7_outputs(4712) <= not a or b;
    layer7_outputs(4713) <= a and b;
    layer7_outputs(4714) <= b and not a;
    layer7_outputs(4715) <= not a or b;
    layer7_outputs(4716) <= not (a and b);
    layer7_outputs(4717) <= b and not a;
    layer7_outputs(4718) <= a xor b;
    layer7_outputs(4719) <= not (a and b);
    layer7_outputs(4720) <= not (a xor b);
    layer7_outputs(4721) <= b and not a;
    layer7_outputs(4722) <= not (a or b);
    layer7_outputs(4723) <= a;
    layer7_outputs(4724) <= not b;
    layer7_outputs(4725) <= a;
    layer7_outputs(4726) <= not a;
    layer7_outputs(4727) <= a and not b;
    layer7_outputs(4728) <= not a or b;
    layer7_outputs(4729) <= not b;
    layer7_outputs(4730) <= not a;
    layer7_outputs(4731) <= a and b;
    layer7_outputs(4732) <= not a;
    layer7_outputs(4733) <= not b;
    layer7_outputs(4734) <= a;
    layer7_outputs(4735) <= not (a or b);
    layer7_outputs(4736) <= a;
    layer7_outputs(4737) <= not (a xor b);
    layer7_outputs(4738) <= not a or b;
    layer7_outputs(4739) <= not b;
    layer7_outputs(4740) <= not b;
    layer7_outputs(4741) <= not (a xor b);
    layer7_outputs(4742) <= not (a or b);
    layer7_outputs(4743) <= a xor b;
    layer7_outputs(4744) <= not a;
    layer7_outputs(4745) <= a;
    layer7_outputs(4746) <= a;
    layer7_outputs(4747) <= '1';
    layer7_outputs(4748) <= not (a and b);
    layer7_outputs(4749) <= not (a xor b);
    layer7_outputs(4750) <= not a;
    layer7_outputs(4751) <= a and not b;
    layer7_outputs(4752) <= a and not b;
    layer7_outputs(4753) <= a and b;
    layer7_outputs(4754) <= not b or a;
    layer7_outputs(4755) <= not a;
    layer7_outputs(4756) <= not (a xor b);
    layer7_outputs(4757) <= a or b;
    layer7_outputs(4758) <= '0';
    layer7_outputs(4759) <= a xor b;
    layer7_outputs(4760) <= not a;
    layer7_outputs(4761) <= b;
    layer7_outputs(4762) <= b and not a;
    layer7_outputs(4763) <= not a or b;
    layer7_outputs(4764) <= not b or a;
    layer7_outputs(4765) <= a;
    layer7_outputs(4766) <= not b;
    layer7_outputs(4767) <= b and not a;
    layer7_outputs(4768) <= a xor b;
    layer7_outputs(4769) <= b;
    layer7_outputs(4770) <= not (a and b);
    layer7_outputs(4771) <= not b;
    layer7_outputs(4772) <= not b or a;
    layer7_outputs(4773) <= a;
    layer7_outputs(4774) <= not a or b;
    layer7_outputs(4775) <= not (a and b);
    layer7_outputs(4776) <= a xor b;
    layer7_outputs(4777) <= a xor b;
    layer7_outputs(4778) <= not a;
    layer7_outputs(4779) <= b;
    layer7_outputs(4780) <= not b;
    layer7_outputs(4781) <= b and not a;
    layer7_outputs(4782) <= b;
    layer7_outputs(4783) <= not b;
    layer7_outputs(4784) <= b;
    layer7_outputs(4785) <= not a or b;
    layer7_outputs(4786) <= b and not a;
    layer7_outputs(4787) <= a or b;
    layer7_outputs(4788) <= not a;
    layer7_outputs(4789) <= not a;
    layer7_outputs(4790) <= b;
    layer7_outputs(4791) <= a;
    layer7_outputs(4792) <= a and not b;
    layer7_outputs(4793) <= not b;
    layer7_outputs(4794) <= '0';
    layer7_outputs(4795) <= a and b;
    layer7_outputs(4796) <= not a;
    layer7_outputs(4797) <= not b;
    layer7_outputs(4798) <= a and b;
    layer7_outputs(4799) <= not b;
    layer7_outputs(4800) <= not (a or b);
    layer7_outputs(4801) <= '0';
    layer7_outputs(4802) <= not (a xor b);
    layer7_outputs(4803) <= not (a or b);
    layer7_outputs(4804) <= a and b;
    layer7_outputs(4805) <= a;
    layer7_outputs(4806) <= not (a xor b);
    layer7_outputs(4807) <= b;
    layer7_outputs(4808) <= b;
    layer7_outputs(4809) <= a xor b;
    layer7_outputs(4810) <= not (a or b);
    layer7_outputs(4811) <= not b;
    layer7_outputs(4812) <= a and not b;
    layer7_outputs(4813) <= not a;
    layer7_outputs(4814) <= a and b;
    layer7_outputs(4815) <= b and not a;
    layer7_outputs(4816) <= b;
    layer7_outputs(4817) <= not (a xor b);
    layer7_outputs(4818) <= a;
    layer7_outputs(4819) <= a and not b;
    layer7_outputs(4820) <= not b or a;
    layer7_outputs(4821) <= a;
    layer7_outputs(4822) <= b;
    layer7_outputs(4823) <= b;
    layer7_outputs(4824) <= a and b;
    layer7_outputs(4825) <= '1';
    layer7_outputs(4826) <= a and b;
    layer7_outputs(4827) <= not b;
    layer7_outputs(4828) <= a and b;
    layer7_outputs(4829) <= a;
    layer7_outputs(4830) <= b and not a;
    layer7_outputs(4831) <= not b;
    layer7_outputs(4832) <= not b;
    layer7_outputs(4833) <= a and not b;
    layer7_outputs(4834) <= not b;
    layer7_outputs(4835) <= not (a xor b);
    layer7_outputs(4836) <= b and not a;
    layer7_outputs(4837) <= b;
    layer7_outputs(4838) <= '1';
    layer7_outputs(4839) <= not (a and b);
    layer7_outputs(4840) <= not (a xor b);
    layer7_outputs(4841) <= b;
    layer7_outputs(4842) <= not (a xor b);
    layer7_outputs(4843) <= a;
    layer7_outputs(4844) <= b and not a;
    layer7_outputs(4845) <= not a or b;
    layer7_outputs(4846) <= a;
    layer7_outputs(4847) <= not (a xor b);
    layer7_outputs(4848) <= b;
    layer7_outputs(4849) <= a;
    layer7_outputs(4850) <= not a;
    layer7_outputs(4851) <= a or b;
    layer7_outputs(4852) <= b;
    layer7_outputs(4853) <= a and not b;
    layer7_outputs(4854) <= a or b;
    layer7_outputs(4855) <= not a;
    layer7_outputs(4856) <= not (a and b);
    layer7_outputs(4857) <= not a;
    layer7_outputs(4858) <= not b;
    layer7_outputs(4859) <= a;
    layer7_outputs(4860) <= a xor b;
    layer7_outputs(4861) <= b;
    layer7_outputs(4862) <= not b;
    layer7_outputs(4863) <= not b;
    layer7_outputs(4864) <= '0';
    layer7_outputs(4865) <= a or b;
    layer7_outputs(4866) <= a xor b;
    layer7_outputs(4867) <= not b or a;
    layer7_outputs(4868) <= a;
    layer7_outputs(4869) <= not a;
    layer7_outputs(4870) <= not b or a;
    layer7_outputs(4871) <= not (a xor b);
    layer7_outputs(4872) <= not a;
    layer7_outputs(4873) <= a or b;
    layer7_outputs(4874) <= b;
    layer7_outputs(4875) <= a or b;
    layer7_outputs(4876) <= not a;
    layer7_outputs(4877) <= not a or b;
    layer7_outputs(4878) <= not (a xor b);
    layer7_outputs(4879) <= not b;
    layer7_outputs(4880) <= a;
    layer7_outputs(4881) <= not (a xor b);
    layer7_outputs(4882) <= not a;
    layer7_outputs(4883) <= not a;
    layer7_outputs(4884) <= not (a xor b);
    layer7_outputs(4885) <= not b or a;
    layer7_outputs(4886) <= not a;
    layer7_outputs(4887) <= not (a and b);
    layer7_outputs(4888) <= not a;
    layer7_outputs(4889) <= not (a xor b);
    layer7_outputs(4890) <= b and not a;
    layer7_outputs(4891) <= not b;
    layer7_outputs(4892) <= a xor b;
    layer7_outputs(4893) <= not b or a;
    layer7_outputs(4894) <= a;
    layer7_outputs(4895) <= a and b;
    layer7_outputs(4896) <= a;
    layer7_outputs(4897) <= b;
    layer7_outputs(4898) <= b;
    layer7_outputs(4899) <= not a;
    layer7_outputs(4900) <= b;
    layer7_outputs(4901) <= not b;
    layer7_outputs(4902) <= not b;
    layer7_outputs(4903) <= a and b;
    layer7_outputs(4904) <= a or b;
    layer7_outputs(4905) <= not a;
    layer7_outputs(4906) <= a xor b;
    layer7_outputs(4907) <= a and not b;
    layer7_outputs(4908) <= a;
    layer7_outputs(4909) <= a and b;
    layer7_outputs(4910) <= a xor b;
    layer7_outputs(4911) <= a xor b;
    layer7_outputs(4912) <= a or b;
    layer7_outputs(4913) <= not a;
    layer7_outputs(4914) <= not a;
    layer7_outputs(4915) <= a or b;
    layer7_outputs(4916) <= b;
    layer7_outputs(4917) <= not (a or b);
    layer7_outputs(4918) <= a xor b;
    layer7_outputs(4919) <= not (a xor b);
    layer7_outputs(4920) <= a and not b;
    layer7_outputs(4921) <= b and not a;
    layer7_outputs(4922) <= a and not b;
    layer7_outputs(4923) <= not (a xor b);
    layer7_outputs(4924) <= '1';
    layer7_outputs(4925) <= b;
    layer7_outputs(4926) <= b;
    layer7_outputs(4927) <= not b;
    layer7_outputs(4928) <= not b;
    layer7_outputs(4929) <= a and b;
    layer7_outputs(4930) <= b and not a;
    layer7_outputs(4931) <= b;
    layer7_outputs(4932) <= not b or a;
    layer7_outputs(4933) <= a;
    layer7_outputs(4934) <= not (a xor b);
    layer7_outputs(4935) <= not a;
    layer7_outputs(4936) <= not b or a;
    layer7_outputs(4937) <= b;
    layer7_outputs(4938) <= not a or b;
    layer7_outputs(4939) <= a xor b;
    layer7_outputs(4940) <= not (a or b);
    layer7_outputs(4941) <= b and not a;
    layer7_outputs(4942) <= a;
    layer7_outputs(4943) <= b and not a;
    layer7_outputs(4944) <= not b;
    layer7_outputs(4945) <= a;
    layer7_outputs(4946) <= not b;
    layer7_outputs(4947) <= not b;
    layer7_outputs(4948) <= a;
    layer7_outputs(4949) <= not b;
    layer7_outputs(4950) <= a and not b;
    layer7_outputs(4951) <= not (a xor b);
    layer7_outputs(4952) <= a xor b;
    layer7_outputs(4953) <= not (a or b);
    layer7_outputs(4954) <= not (a or b);
    layer7_outputs(4955) <= a and b;
    layer7_outputs(4956) <= not (a and b);
    layer7_outputs(4957) <= a and not b;
    layer7_outputs(4958) <= a or b;
    layer7_outputs(4959) <= a;
    layer7_outputs(4960) <= not a or b;
    layer7_outputs(4961) <= not (a and b);
    layer7_outputs(4962) <= b;
    layer7_outputs(4963) <= a and not b;
    layer7_outputs(4964) <= b and not a;
    layer7_outputs(4965) <= not (a xor b);
    layer7_outputs(4966) <= not a;
    layer7_outputs(4967) <= a;
    layer7_outputs(4968) <= not (a xor b);
    layer7_outputs(4969) <= '1';
    layer7_outputs(4970) <= a;
    layer7_outputs(4971) <= b;
    layer7_outputs(4972) <= not a or b;
    layer7_outputs(4973) <= not (a and b);
    layer7_outputs(4974) <= not b;
    layer7_outputs(4975) <= a and not b;
    layer7_outputs(4976) <= not (a xor b);
    layer7_outputs(4977) <= '1';
    layer7_outputs(4978) <= not a;
    layer7_outputs(4979) <= b and not a;
    layer7_outputs(4980) <= a or b;
    layer7_outputs(4981) <= a xor b;
    layer7_outputs(4982) <= not a or b;
    layer7_outputs(4983) <= not a or b;
    layer7_outputs(4984) <= not a;
    layer7_outputs(4985) <= '0';
    layer7_outputs(4986) <= a or b;
    layer7_outputs(4987) <= not (a or b);
    layer7_outputs(4988) <= a;
    layer7_outputs(4989) <= not a;
    layer7_outputs(4990) <= b;
    layer7_outputs(4991) <= not (a xor b);
    layer7_outputs(4992) <= a;
    layer7_outputs(4993) <= b and not a;
    layer7_outputs(4994) <= not (a xor b);
    layer7_outputs(4995) <= not a or b;
    layer7_outputs(4996) <= a;
    layer7_outputs(4997) <= b;
    layer7_outputs(4998) <= a;
    layer7_outputs(4999) <= b and not a;
    layer7_outputs(5000) <= b;
    layer7_outputs(5001) <= not b;
    layer7_outputs(5002) <= not a or b;
    layer7_outputs(5003) <= b;
    layer7_outputs(5004) <= b;
    layer7_outputs(5005) <= a and b;
    layer7_outputs(5006) <= a xor b;
    layer7_outputs(5007) <= a;
    layer7_outputs(5008) <= not a;
    layer7_outputs(5009) <= b;
    layer7_outputs(5010) <= a xor b;
    layer7_outputs(5011) <= a or b;
    layer7_outputs(5012) <= a and b;
    layer7_outputs(5013) <= not b;
    layer7_outputs(5014) <= a and b;
    layer7_outputs(5015) <= a;
    layer7_outputs(5016) <= not b;
    layer7_outputs(5017) <= a xor b;
    layer7_outputs(5018) <= a;
    layer7_outputs(5019) <= a xor b;
    layer7_outputs(5020) <= not b;
    layer7_outputs(5021) <= a xor b;
    layer7_outputs(5022) <= b;
    layer7_outputs(5023) <= a and not b;
    layer7_outputs(5024) <= b;
    layer7_outputs(5025) <= b;
    layer7_outputs(5026) <= not a or b;
    layer7_outputs(5027) <= not b;
    layer7_outputs(5028) <= not b;
    layer7_outputs(5029) <= a and not b;
    layer7_outputs(5030) <= not (a or b);
    layer7_outputs(5031) <= not a or b;
    layer7_outputs(5032) <= not (a or b);
    layer7_outputs(5033) <= not b or a;
    layer7_outputs(5034) <= b;
    layer7_outputs(5035) <= a or b;
    layer7_outputs(5036) <= b;
    layer7_outputs(5037) <= a;
    layer7_outputs(5038) <= b and not a;
    layer7_outputs(5039) <= not (a or b);
    layer7_outputs(5040) <= a;
    layer7_outputs(5041) <= not b;
    layer7_outputs(5042) <= not a;
    layer7_outputs(5043) <= b;
    layer7_outputs(5044) <= not (a or b);
    layer7_outputs(5045) <= b;
    layer7_outputs(5046) <= a xor b;
    layer7_outputs(5047) <= not (a xor b);
    layer7_outputs(5048) <= b and not a;
    layer7_outputs(5049) <= not a or b;
    layer7_outputs(5050) <= not a;
    layer7_outputs(5051) <= not b;
    layer7_outputs(5052) <= a and not b;
    layer7_outputs(5053) <= not a or b;
    layer7_outputs(5054) <= not b;
    layer7_outputs(5055) <= not a or b;
    layer7_outputs(5056) <= not a;
    layer7_outputs(5057) <= not b;
    layer7_outputs(5058) <= a and b;
    layer7_outputs(5059) <= not (a and b);
    layer7_outputs(5060) <= not b or a;
    layer7_outputs(5061) <= a xor b;
    layer7_outputs(5062) <= not (a or b);
    layer7_outputs(5063) <= a xor b;
    layer7_outputs(5064) <= a;
    layer7_outputs(5065) <= not a;
    layer7_outputs(5066) <= b;
    layer7_outputs(5067) <= not b or a;
    layer7_outputs(5068) <= not b;
    layer7_outputs(5069) <= b and not a;
    layer7_outputs(5070) <= not a;
    layer7_outputs(5071) <= not (a xor b);
    layer7_outputs(5072) <= a;
    layer7_outputs(5073) <= not a;
    layer7_outputs(5074) <= not b;
    layer7_outputs(5075) <= not a;
    layer7_outputs(5076) <= a and not b;
    layer7_outputs(5077) <= b;
    layer7_outputs(5078) <= b;
    layer7_outputs(5079) <= not a;
    layer7_outputs(5080) <= a;
    layer7_outputs(5081) <= not (a and b);
    layer7_outputs(5082) <= not a;
    layer7_outputs(5083) <= a and not b;
    layer7_outputs(5084) <= b and not a;
    layer7_outputs(5085) <= a;
    layer7_outputs(5086) <= not b;
    layer7_outputs(5087) <= not a or b;
    layer7_outputs(5088) <= not b;
    layer7_outputs(5089) <= not a;
    layer7_outputs(5090) <= not b;
    layer7_outputs(5091) <= not a or b;
    layer7_outputs(5092) <= a and b;
    layer7_outputs(5093) <= a;
    layer7_outputs(5094) <= not (a xor b);
    layer7_outputs(5095) <= b;
    layer7_outputs(5096) <= not (a xor b);
    layer7_outputs(5097) <= not (a xor b);
    layer7_outputs(5098) <= a;
    layer7_outputs(5099) <= not (a and b);
    layer7_outputs(5100) <= a;
    layer7_outputs(5101) <= not b;
    layer7_outputs(5102) <= a;
    layer7_outputs(5103) <= b;
    layer7_outputs(5104) <= a xor b;
    layer7_outputs(5105) <= a;
    layer7_outputs(5106) <= not b;
    layer7_outputs(5107) <= a and b;
    layer7_outputs(5108) <= b;
    layer7_outputs(5109) <= not (a xor b);
    layer7_outputs(5110) <= a and not b;
    layer7_outputs(5111) <= not b or a;
    layer7_outputs(5112) <= b and not a;
    layer7_outputs(5113) <= not a or b;
    layer7_outputs(5114) <= a;
    layer7_outputs(5115) <= not a or b;
    layer7_outputs(5116) <= not a;
    layer7_outputs(5117) <= a and b;
    layer7_outputs(5118) <= b and not a;
    layer7_outputs(5119) <= b and not a;
    layer8_outputs(0) <= a or b;
    layer8_outputs(1) <= not b;
    layer8_outputs(2) <= a or b;
    layer8_outputs(3) <= not (a xor b);
    layer8_outputs(4) <= b and not a;
    layer8_outputs(5) <= a;
    layer8_outputs(6) <= b;
    layer8_outputs(7) <= not a;
    layer8_outputs(8) <= not (a and b);
    layer8_outputs(9) <= not a;
    layer8_outputs(10) <= a xor b;
    layer8_outputs(11) <= a;
    layer8_outputs(12) <= not a;
    layer8_outputs(13) <= a and not b;
    layer8_outputs(14) <= b;
    layer8_outputs(15) <= b;
    layer8_outputs(16) <= not b;
    layer8_outputs(17) <= a;
    layer8_outputs(18) <= not a or b;
    layer8_outputs(19) <= not (a or b);
    layer8_outputs(20) <= not (a xor b);
    layer8_outputs(21) <= a and not b;
    layer8_outputs(22) <= b;
    layer8_outputs(23) <= not b or a;
    layer8_outputs(24) <= a xor b;
    layer8_outputs(25) <= a;
    layer8_outputs(26) <= not a;
    layer8_outputs(27) <= a or b;
    layer8_outputs(28) <= not a;
    layer8_outputs(29) <= not a or b;
    layer8_outputs(30) <= b;
    layer8_outputs(31) <= not (a xor b);
    layer8_outputs(32) <= b;
    layer8_outputs(33) <= not (a xor b);
    layer8_outputs(34) <= '0';
    layer8_outputs(35) <= b;
    layer8_outputs(36) <= a and not b;
    layer8_outputs(37) <= not a or b;
    layer8_outputs(38) <= a;
    layer8_outputs(39) <= not b;
    layer8_outputs(40) <= not (a xor b);
    layer8_outputs(41) <= b;
    layer8_outputs(42) <= b;
    layer8_outputs(43) <= not (a or b);
    layer8_outputs(44) <= a;
    layer8_outputs(45) <= not (a and b);
    layer8_outputs(46) <= a xor b;
    layer8_outputs(47) <= not a;
    layer8_outputs(48) <= not b;
    layer8_outputs(49) <= a or b;
    layer8_outputs(50) <= not b;
    layer8_outputs(51) <= a;
    layer8_outputs(52) <= a xor b;
    layer8_outputs(53) <= not (a and b);
    layer8_outputs(54) <= a;
    layer8_outputs(55) <= not (a or b);
    layer8_outputs(56) <= not a;
    layer8_outputs(57) <= a;
    layer8_outputs(58) <= not a or b;
    layer8_outputs(59) <= a xor b;
    layer8_outputs(60) <= b;
    layer8_outputs(61) <= not (a xor b);
    layer8_outputs(62) <= not a;
    layer8_outputs(63) <= b;
    layer8_outputs(64) <= a xor b;
    layer8_outputs(65) <= a xor b;
    layer8_outputs(66) <= not (a xor b);
    layer8_outputs(67) <= a xor b;
    layer8_outputs(68) <= b and not a;
    layer8_outputs(69) <= not (a and b);
    layer8_outputs(70) <= a or b;
    layer8_outputs(71) <= not (a or b);
    layer8_outputs(72) <= not b or a;
    layer8_outputs(73) <= a or b;
    layer8_outputs(74) <= a xor b;
    layer8_outputs(75) <= not a or b;
    layer8_outputs(76) <= a;
    layer8_outputs(77) <= a;
    layer8_outputs(78) <= not a;
    layer8_outputs(79) <= a or b;
    layer8_outputs(80) <= not a;
    layer8_outputs(81) <= a and not b;
    layer8_outputs(82) <= b;
    layer8_outputs(83) <= a and b;
    layer8_outputs(84) <= not (a and b);
    layer8_outputs(85) <= a and b;
    layer8_outputs(86) <= a and b;
    layer8_outputs(87) <= not (a or b);
    layer8_outputs(88) <= not (a xor b);
    layer8_outputs(89) <= not (a xor b);
    layer8_outputs(90) <= a or b;
    layer8_outputs(91) <= b;
    layer8_outputs(92) <= not b;
    layer8_outputs(93) <= not b;
    layer8_outputs(94) <= not a;
    layer8_outputs(95) <= a xor b;
    layer8_outputs(96) <= not (a xor b);
    layer8_outputs(97) <= not (a and b);
    layer8_outputs(98) <= not b or a;
    layer8_outputs(99) <= '1';
    layer8_outputs(100) <= not a;
    layer8_outputs(101) <= not (a and b);
    layer8_outputs(102) <= a xor b;
    layer8_outputs(103) <= a and not b;
    layer8_outputs(104) <= a;
    layer8_outputs(105) <= a or b;
    layer8_outputs(106) <= a and not b;
    layer8_outputs(107) <= a;
    layer8_outputs(108) <= a and not b;
    layer8_outputs(109) <= a xor b;
    layer8_outputs(110) <= '0';
    layer8_outputs(111) <= not (a xor b);
    layer8_outputs(112) <= b;
    layer8_outputs(113) <= a and b;
    layer8_outputs(114) <= a xor b;
    layer8_outputs(115) <= a and not b;
    layer8_outputs(116) <= not b;
    layer8_outputs(117) <= not (a xor b);
    layer8_outputs(118) <= b;
    layer8_outputs(119) <= a xor b;
    layer8_outputs(120) <= not a;
    layer8_outputs(121) <= a xor b;
    layer8_outputs(122) <= not a;
    layer8_outputs(123) <= b and not a;
    layer8_outputs(124) <= not (a xor b);
    layer8_outputs(125) <= not a or b;
    layer8_outputs(126) <= a and b;
    layer8_outputs(127) <= not a;
    layer8_outputs(128) <= a;
    layer8_outputs(129) <= a xor b;
    layer8_outputs(130) <= '1';
    layer8_outputs(131) <= not a;
    layer8_outputs(132) <= not (a xor b);
    layer8_outputs(133) <= b;
    layer8_outputs(134) <= a xor b;
    layer8_outputs(135) <= b;
    layer8_outputs(136) <= a and b;
    layer8_outputs(137) <= b;
    layer8_outputs(138) <= b and not a;
    layer8_outputs(139) <= b;
    layer8_outputs(140) <= b;
    layer8_outputs(141) <= a xor b;
    layer8_outputs(142) <= b;
    layer8_outputs(143) <= not b;
    layer8_outputs(144) <= not (a xor b);
    layer8_outputs(145) <= a;
    layer8_outputs(146) <= a;
    layer8_outputs(147) <= a xor b;
    layer8_outputs(148) <= a and not b;
    layer8_outputs(149) <= a;
    layer8_outputs(150) <= not b or a;
    layer8_outputs(151) <= not a or b;
    layer8_outputs(152) <= not (a xor b);
    layer8_outputs(153) <= b and not a;
    layer8_outputs(154) <= b;
    layer8_outputs(155) <= a;
    layer8_outputs(156) <= not b or a;
    layer8_outputs(157) <= not a;
    layer8_outputs(158) <= not b;
    layer8_outputs(159) <= b;
    layer8_outputs(160) <= a;
    layer8_outputs(161) <= not b;
    layer8_outputs(162) <= not b;
    layer8_outputs(163) <= '0';
    layer8_outputs(164) <= not (a xor b);
    layer8_outputs(165) <= b;
    layer8_outputs(166) <= not a;
    layer8_outputs(167) <= a or b;
    layer8_outputs(168) <= a and b;
    layer8_outputs(169) <= a and not b;
    layer8_outputs(170) <= not (a and b);
    layer8_outputs(171) <= not a;
    layer8_outputs(172) <= a and b;
    layer8_outputs(173) <= b;
    layer8_outputs(174) <= a and not b;
    layer8_outputs(175) <= a xor b;
    layer8_outputs(176) <= not (a xor b);
    layer8_outputs(177) <= not a;
    layer8_outputs(178) <= a;
    layer8_outputs(179) <= '1';
    layer8_outputs(180) <= not (a xor b);
    layer8_outputs(181) <= not (a xor b);
    layer8_outputs(182) <= not b;
    layer8_outputs(183) <= a and not b;
    layer8_outputs(184) <= b and not a;
    layer8_outputs(185) <= a;
    layer8_outputs(186) <= not (a or b);
    layer8_outputs(187) <= not (a xor b);
    layer8_outputs(188) <= not (a and b);
    layer8_outputs(189) <= not a;
    layer8_outputs(190) <= not (a or b);
    layer8_outputs(191) <= b;
    layer8_outputs(192) <= b;
    layer8_outputs(193) <= b and not a;
    layer8_outputs(194) <= b;
    layer8_outputs(195) <= not (a xor b);
    layer8_outputs(196) <= not b or a;
    layer8_outputs(197) <= b;
    layer8_outputs(198) <= not b;
    layer8_outputs(199) <= a and b;
    layer8_outputs(200) <= b;
    layer8_outputs(201) <= not b;
    layer8_outputs(202) <= a and not b;
    layer8_outputs(203) <= not (a xor b);
    layer8_outputs(204) <= a and not b;
    layer8_outputs(205) <= b and not a;
    layer8_outputs(206) <= not (a xor b);
    layer8_outputs(207) <= not (a xor b);
    layer8_outputs(208) <= not (a xor b);
    layer8_outputs(209) <= not b;
    layer8_outputs(210) <= a xor b;
    layer8_outputs(211) <= not a or b;
    layer8_outputs(212) <= not a or b;
    layer8_outputs(213) <= not b or a;
    layer8_outputs(214) <= not a;
    layer8_outputs(215) <= a;
    layer8_outputs(216) <= not (a xor b);
    layer8_outputs(217) <= not b;
    layer8_outputs(218) <= a xor b;
    layer8_outputs(219) <= a;
    layer8_outputs(220) <= not a;
    layer8_outputs(221) <= not b or a;
    layer8_outputs(222) <= not (a xor b);
    layer8_outputs(223) <= not b;
    layer8_outputs(224) <= a;
    layer8_outputs(225) <= a;
    layer8_outputs(226) <= not a;
    layer8_outputs(227) <= a and not b;
    layer8_outputs(228) <= b;
    layer8_outputs(229) <= a;
    layer8_outputs(230) <= a;
    layer8_outputs(231) <= a or b;
    layer8_outputs(232) <= not a;
    layer8_outputs(233) <= not b;
    layer8_outputs(234) <= not (a and b);
    layer8_outputs(235) <= b;
    layer8_outputs(236) <= a and b;
    layer8_outputs(237) <= not b;
    layer8_outputs(238) <= not (a or b);
    layer8_outputs(239) <= not a;
    layer8_outputs(240) <= a and b;
    layer8_outputs(241) <= b;
    layer8_outputs(242) <= a;
    layer8_outputs(243) <= not b or a;
    layer8_outputs(244) <= not (a xor b);
    layer8_outputs(245) <= not (a or b);
    layer8_outputs(246) <= a and not b;
    layer8_outputs(247) <= a xor b;
    layer8_outputs(248) <= not (a xor b);
    layer8_outputs(249) <= a and not b;
    layer8_outputs(250) <= b;
    layer8_outputs(251) <= not b or a;
    layer8_outputs(252) <= b;
    layer8_outputs(253) <= not b;
    layer8_outputs(254) <= b and not a;
    layer8_outputs(255) <= not (a and b);
    layer8_outputs(256) <= a;
    layer8_outputs(257) <= a;
    layer8_outputs(258) <= b;
    layer8_outputs(259) <= not b;
    layer8_outputs(260) <= not (a or b);
    layer8_outputs(261) <= a or b;
    layer8_outputs(262) <= b and not a;
    layer8_outputs(263) <= a and b;
    layer8_outputs(264) <= a xor b;
    layer8_outputs(265) <= not (a xor b);
    layer8_outputs(266) <= not a or b;
    layer8_outputs(267) <= not a or b;
    layer8_outputs(268) <= b and not a;
    layer8_outputs(269) <= not (a xor b);
    layer8_outputs(270) <= not a;
    layer8_outputs(271) <= b and not a;
    layer8_outputs(272) <= not a;
    layer8_outputs(273) <= b;
    layer8_outputs(274) <= not b or a;
    layer8_outputs(275) <= not b;
    layer8_outputs(276) <= not b;
    layer8_outputs(277) <= a or b;
    layer8_outputs(278) <= not b;
    layer8_outputs(279) <= not b;
    layer8_outputs(280) <= a;
    layer8_outputs(281) <= not a;
    layer8_outputs(282) <= not (a and b);
    layer8_outputs(283) <= a;
    layer8_outputs(284) <= a and b;
    layer8_outputs(285) <= not (a and b);
    layer8_outputs(286) <= not (a xor b);
    layer8_outputs(287) <= a;
    layer8_outputs(288) <= not (a xor b);
    layer8_outputs(289) <= a or b;
    layer8_outputs(290) <= a and not b;
    layer8_outputs(291) <= a or b;
    layer8_outputs(292) <= not b;
    layer8_outputs(293) <= not b;
    layer8_outputs(294) <= b;
    layer8_outputs(295) <= a and b;
    layer8_outputs(296) <= not a;
    layer8_outputs(297) <= b;
    layer8_outputs(298) <= not (a and b);
    layer8_outputs(299) <= a xor b;
    layer8_outputs(300) <= a or b;
    layer8_outputs(301) <= not b;
    layer8_outputs(302) <= a;
    layer8_outputs(303) <= a xor b;
    layer8_outputs(304) <= a and b;
    layer8_outputs(305) <= a;
    layer8_outputs(306) <= '0';
    layer8_outputs(307) <= not a;
    layer8_outputs(308) <= a or b;
    layer8_outputs(309) <= a and b;
    layer8_outputs(310) <= b;
    layer8_outputs(311) <= not (a xor b);
    layer8_outputs(312) <= not a or b;
    layer8_outputs(313) <= a xor b;
    layer8_outputs(314) <= not a;
    layer8_outputs(315) <= not (a or b);
    layer8_outputs(316) <= not (a or b);
    layer8_outputs(317) <= not (a xor b);
    layer8_outputs(318) <= a xor b;
    layer8_outputs(319) <= a or b;
    layer8_outputs(320) <= b and not a;
    layer8_outputs(321) <= a;
    layer8_outputs(322) <= not (a xor b);
    layer8_outputs(323) <= a xor b;
    layer8_outputs(324) <= not a;
    layer8_outputs(325) <= a xor b;
    layer8_outputs(326) <= a xor b;
    layer8_outputs(327) <= a;
    layer8_outputs(328) <= not a;
    layer8_outputs(329) <= a;
    layer8_outputs(330) <= not a or b;
    layer8_outputs(331) <= not a;
    layer8_outputs(332) <= not (a xor b);
    layer8_outputs(333) <= not a;
    layer8_outputs(334) <= a or b;
    layer8_outputs(335) <= a xor b;
    layer8_outputs(336) <= not b;
    layer8_outputs(337) <= b and not a;
    layer8_outputs(338) <= a xor b;
    layer8_outputs(339) <= a xor b;
    layer8_outputs(340) <= not (a or b);
    layer8_outputs(341) <= b and not a;
    layer8_outputs(342) <= not a or b;
    layer8_outputs(343) <= not b;
    layer8_outputs(344) <= not (a or b);
    layer8_outputs(345) <= not (a xor b);
    layer8_outputs(346) <= a xor b;
    layer8_outputs(347) <= not (a xor b);
    layer8_outputs(348) <= a xor b;
    layer8_outputs(349) <= not (a xor b);
    layer8_outputs(350) <= a or b;
    layer8_outputs(351) <= a;
    layer8_outputs(352) <= a xor b;
    layer8_outputs(353) <= a and b;
    layer8_outputs(354) <= not (a xor b);
    layer8_outputs(355) <= not b;
    layer8_outputs(356) <= not b;
    layer8_outputs(357) <= a xor b;
    layer8_outputs(358) <= not (a or b);
    layer8_outputs(359) <= a;
    layer8_outputs(360) <= a xor b;
    layer8_outputs(361) <= not b;
    layer8_outputs(362) <= b and not a;
    layer8_outputs(363) <= not (a xor b);
    layer8_outputs(364) <= not b;
    layer8_outputs(365) <= b and not a;
    layer8_outputs(366) <= b;
    layer8_outputs(367) <= not b;
    layer8_outputs(368) <= a xor b;
    layer8_outputs(369) <= a xor b;
    layer8_outputs(370) <= a;
    layer8_outputs(371) <= a and not b;
    layer8_outputs(372) <= a;
    layer8_outputs(373) <= a xor b;
    layer8_outputs(374) <= not (a xor b);
    layer8_outputs(375) <= not (a or b);
    layer8_outputs(376) <= '0';
    layer8_outputs(377) <= a and b;
    layer8_outputs(378) <= a;
    layer8_outputs(379) <= a xor b;
    layer8_outputs(380) <= not b;
    layer8_outputs(381) <= b and not a;
    layer8_outputs(382) <= a;
    layer8_outputs(383) <= not a;
    layer8_outputs(384) <= a xor b;
    layer8_outputs(385) <= a or b;
    layer8_outputs(386) <= b;
    layer8_outputs(387) <= a or b;
    layer8_outputs(388) <= not a;
    layer8_outputs(389) <= a xor b;
    layer8_outputs(390) <= not (a xor b);
    layer8_outputs(391) <= not a or b;
    layer8_outputs(392) <= a;
    layer8_outputs(393) <= not (a or b);
    layer8_outputs(394) <= not (a xor b);
    layer8_outputs(395) <= not b;
    layer8_outputs(396) <= not b;
    layer8_outputs(397) <= not a;
    layer8_outputs(398) <= not b;
    layer8_outputs(399) <= a and not b;
    layer8_outputs(400) <= a xor b;
    layer8_outputs(401) <= not b;
    layer8_outputs(402) <= b;
    layer8_outputs(403) <= a xor b;
    layer8_outputs(404) <= not a or b;
    layer8_outputs(405) <= b;
    layer8_outputs(406) <= a and b;
    layer8_outputs(407) <= b;
    layer8_outputs(408) <= b;
    layer8_outputs(409) <= not (a and b);
    layer8_outputs(410) <= a;
    layer8_outputs(411) <= not b;
    layer8_outputs(412) <= not b or a;
    layer8_outputs(413) <= a and b;
    layer8_outputs(414) <= not (a or b);
    layer8_outputs(415) <= not (a xor b);
    layer8_outputs(416) <= not (a xor b);
    layer8_outputs(417) <= a;
    layer8_outputs(418) <= not (a or b);
    layer8_outputs(419) <= a;
    layer8_outputs(420) <= b and not a;
    layer8_outputs(421) <= not b or a;
    layer8_outputs(422) <= not (a xor b);
    layer8_outputs(423) <= a or b;
    layer8_outputs(424) <= not a;
    layer8_outputs(425) <= a xor b;
    layer8_outputs(426) <= a;
    layer8_outputs(427) <= not b;
    layer8_outputs(428) <= a and b;
    layer8_outputs(429) <= not b;
    layer8_outputs(430) <= not (a xor b);
    layer8_outputs(431) <= not (a xor b);
    layer8_outputs(432) <= b and not a;
    layer8_outputs(433) <= not (a xor b);
    layer8_outputs(434) <= a;
    layer8_outputs(435) <= a xor b;
    layer8_outputs(436) <= not a or b;
    layer8_outputs(437) <= b and not a;
    layer8_outputs(438) <= a;
    layer8_outputs(439) <= not b;
    layer8_outputs(440) <= not b;
    layer8_outputs(441) <= not a;
    layer8_outputs(442) <= a xor b;
    layer8_outputs(443) <= a xor b;
    layer8_outputs(444) <= not (a xor b);
    layer8_outputs(445) <= a xor b;
    layer8_outputs(446) <= not (a xor b);
    layer8_outputs(447) <= not b or a;
    layer8_outputs(448) <= b and not a;
    layer8_outputs(449) <= not a;
    layer8_outputs(450) <= a xor b;
    layer8_outputs(451) <= b;
    layer8_outputs(452) <= not (a and b);
    layer8_outputs(453) <= b and not a;
    layer8_outputs(454) <= b;
    layer8_outputs(455) <= not (a or b);
    layer8_outputs(456) <= a xor b;
    layer8_outputs(457) <= not a;
    layer8_outputs(458) <= a and not b;
    layer8_outputs(459) <= a;
    layer8_outputs(460) <= a xor b;
    layer8_outputs(461) <= a and not b;
    layer8_outputs(462) <= not b;
    layer8_outputs(463) <= b;
    layer8_outputs(464) <= not (a xor b);
    layer8_outputs(465) <= not b;
    layer8_outputs(466) <= not a;
    layer8_outputs(467) <= not (a and b);
    layer8_outputs(468) <= not (a xor b);
    layer8_outputs(469) <= a xor b;
    layer8_outputs(470) <= not a;
    layer8_outputs(471) <= a xor b;
    layer8_outputs(472) <= b;
    layer8_outputs(473) <= '1';
    layer8_outputs(474) <= a and b;
    layer8_outputs(475) <= not (a xor b);
    layer8_outputs(476) <= '1';
    layer8_outputs(477) <= not a;
    layer8_outputs(478) <= b;
    layer8_outputs(479) <= b;
    layer8_outputs(480) <= not (a xor b);
    layer8_outputs(481) <= a xor b;
    layer8_outputs(482) <= a;
    layer8_outputs(483) <= not a;
    layer8_outputs(484) <= not a or b;
    layer8_outputs(485) <= not a;
    layer8_outputs(486) <= a;
    layer8_outputs(487) <= a and b;
    layer8_outputs(488) <= b;
    layer8_outputs(489) <= not b;
    layer8_outputs(490) <= b and not a;
    layer8_outputs(491) <= not a;
    layer8_outputs(492) <= not (a xor b);
    layer8_outputs(493) <= not b or a;
    layer8_outputs(494) <= a or b;
    layer8_outputs(495) <= a xor b;
    layer8_outputs(496) <= not a or b;
    layer8_outputs(497) <= a;
    layer8_outputs(498) <= a or b;
    layer8_outputs(499) <= not b;
    layer8_outputs(500) <= not a;
    layer8_outputs(501) <= a;
    layer8_outputs(502) <= a and not b;
    layer8_outputs(503) <= a;
    layer8_outputs(504) <= a;
    layer8_outputs(505) <= a and b;
    layer8_outputs(506) <= not b;
    layer8_outputs(507) <= not (a xor b);
    layer8_outputs(508) <= not b;
    layer8_outputs(509) <= not a;
    layer8_outputs(510) <= not a or b;
    layer8_outputs(511) <= not (a or b);
    layer8_outputs(512) <= a;
    layer8_outputs(513) <= a xor b;
    layer8_outputs(514) <= b and not a;
    layer8_outputs(515) <= not (a or b);
    layer8_outputs(516) <= not b or a;
    layer8_outputs(517) <= a xor b;
    layer8_outputs(518) <= not b or a;
    layer8_outputs(519) <= b;
    layer8_outputs(520) <= b;
    layer8_outputs(521) <= a;
    layer8_outputs(522) <= a xor b;
    layer8_outputs(523) <= not b;
    layer8_outputs(524) <= a;
    layer8_outputs(525) <= a xor b;
    layer8_outputs(526) <= not (a xor b);
    layer8_outputs(527) <= not (a xor b);
    layer8_outputs(528) <= not b;
    layer8_outputs(529) <= a xor b;
    layer8_outputs(530) <= a;
    layer8_outputs(531) <= a;
    layer8_outputs(532) <= a or b;
    layer8_outputs(533) <= a;
    layer8_outputs(534) <= not a;
    layer8_outputs(535) <= not b or a;
    layer8_outputs(536) <= not b;
    layer8_outputs(537) <= a;
    layer8_outputs(538) <= not a or b;
    layer8_outputs(539) <= a;
    layer8_outputs(540) <= a xor b;
    layer8_outputs(541) <= a;
    layer8_outputs(542) <= not b or a;
    layer8_outputs(543) <= a xor b;
    layer8_outputs(544) <= not a;
    layer8_outputs(545) <= a;
    layer8_outputs(546) <= not a;
    layer8_outputs(547) <= a xor b;
    layer8_outputs(548) <= not (a xor b);
    layer8_outputs(549) <= not b;
    layer8_outputs(550) <= b and not a;
    layer8_outputs(551) <= not a;
    layer8_outputs(552) <= b;
    layer8_outputs(553) <= not a;
    layer8_outputs(554) <= b;
    layer8_outputs(555) <= not b;
    layer8_outputs(556) <= not (a or b);
    layer8_outputs(557) <= not (a and b);
    layer8_outputs(558) <= not a or b;
    layer8_outputs(559) <= not a;
    layer8_outputs(560) <= not b;
    layer8_outputs(561) <= a or b;
    layer8_outputs(562) <= not (a xor b);
    layer8_outputs(563) <= not a;
    layer8_outputs(564) <= a or b;
    layer8_outputs(565) <= a and b;
    layer8_outputs(566) <= a xor b;
    layer8_outputs(567) <= a;
    layer8_outputs(568) <= a and not b;
    layer8_outputs(569) <= a and b;
    layer8_outputs(570) <= b;
    layer8_outputs(571) <= not a;
    layer8_outputs(572) <= not a;
    layer8_outputs(573) <= '0';
    layer8_outputs(574) <= not a;
    layer8_outputs(575) <= a xor b;
    layer8_outputs(576) <= a xor b;
    layer8_outputs(577) <= a and not b;
    layer8_outputs(578) <= b;
    layer8_outputs(579) <= a xor b;
    layer8_outputs(580) <= not b or a;
    layer8_outputs(581) <= not (a and b);
    layer8_outputs(582) <= not a;
    layer8_outputs(583) <= a xor b;
    layer8_outputs(584) <= '1';
    layer8_outputs(585) <= b;
    layer8_outputs(586) <= a;
    layer8_outputs(587) <= not (a or b);
    layer8_outputs(588) <= b and not a;
    layer8_outputs(589) <= not (a xor b);
    layer8_outputs(590) <= a;
    layer8_outputs(591) <= not a or b;
    layer8_outputs(592) <= a and not b;
    layer8_outputs(593) <= b and not a;
    layer8_outputs(594) <= b and not a;
    layer8_outputs(595) <= a or b;
    layer8_outputs(596) <= not (a or b);
    layer8_outputs(597) <= not b;
    layer8_outputs(598) <= not b or a;
    layer8_outputs(599) <= b and not a;
    layer8_outputs(600) <= not (a xor b);
    layer8_outputs(601) <= not a;
    layer8_outputs(602) <= not b;
    layer8_outputs(603) <= a xor b;
    layer8_outputs(604) <= a xor b;
    layer8_outputs(605) <= a and not b;
    layer8_outputs(606) <= a;
    layer8_outputs(607) <= a and not b;
    layer8_outputs(608) <= a;
    layer8_outputs(609) <= not b or a;
    layer8_outputs(610) <= not b;
    layer8_outputs(611) <= not a;
    layer8_outputs(612) <= b and not a;
    layer8_outputs(613) <= not a;
    layer8_outputs(614) <= b;
    layer8_outputs(615) <= a xor b;
    layer8_outputs(616) <= a and not b;
    layer8_outputs(617) <= b;
    layer8_outputs(618) <= b and not a;
    layer8_outputs(619) <= not (a or b);
    layer8_outputs(620) <= not b;
    layer8_outputs(621) <= b;
    layer8_outputs(622) <= not a;
    layer8_outputs(623) <= not b;
    layer8_outputs(624) <= not (a xor b);
    layer8_outputs(625) <= not b or a;
    layer8_outputs(626) <= b and not a;
    layer8_outputs(627) <= a or b;
    layer8_outputs(628) <= not a;
    layer8_outputs(629) <= a;
    layer8_outputs(630) <= not b;
    layer8_outputs(631) <= not (a xor b);
    layer8_outputs(632) <= b and not a;
    layer8_outputs(633) <= a;
    layer8_outputs(634) <= a xor b;
    layer8_outputs(635) <= a xor b;
    layer8_outputs(636) <= a and not b;
    layer8_outputs(637) <= not a;
    layer8_outputs(638) <= a and b;
    layer8_outputs(639) <= not a;
    layer8_outputs(640) <= not a;
    layer8_outputs(641) <= not a;
    layer8_outputs(642) <= not (a and b);
    layer8_outputs(643) <= not b;
    layer8_outputs(644) <= not a or b;
    layer8_outputs(645) <= not a;
    layer8_outputs(646) <= not b or a;
    layer8_outputs(647) <= not (a xor b);
    layer8_outputs(648) <= a or b;
    layer8_outputs(649) <= a or b;
    layer8_outputs(650) <= not a;
    layer8_outputs(651) <= not b or a;
    layer8_outputs(652) <= not (a and b);
    layer8_outputs(653) <= not b;
    layer8_outputs(654) <= not a;
    layer8_outputs(655) <= not b;
    layer8_outputs(656) <= not b;
    layer8_outputs(657) <= '1';
    layer8_outputs(658) <= not b;
    layer8_outputs(659) <= not (a xor b);
    layer8_outputs(660) <= a;
    layer8_outputs(661) <= a;
    layer8_outputs(662) <= a or b;
    layer8_outputs(663) <= a xor b;
    layer8_outputs(664) <= a and not b;
    layer8_outputs(665) <= not (a xor b);
    layer8_outputs(666) <= not b;
    layer8_outputs(667) <= not b;
    layer8_outputs(668) <= not (a xor b);
    layer8_outputs(669) <= not b;
    layer8_outputs(670) <= not a;
    layer8_outputs(671) <= b;
    layer8_outputs(672) <= b;
    layer8_outputs(673) <= a xor b;
    layer8_outputs(674) <= not (a xor b);
    layer8_outputs(675) <= a xor b;
    layer8_outputs(676) <= a and not b;
    layer8_outputs(677) <= a and b;
    layer8_outputs(678) <= not a;
    layer8_outputs(679) <= not b;
    layer8_outputs(680) <= not a;
    layer8_outputs(681) <= b;
    layer8_outputs(682) <= a xor b;
    layer8_outputs(683) <= not a;
    layer8_outputs(684) <= a;
    layer8_outputs(685) <= b;
    layer8_outputs(686) <= a;
    layer8_outputs(687) <= not (a and b);
    layer8_outputs(688) <= a xor b;
    layer8_outputs(689) <= a xor b;
    layer8_outputs(690) <= a or b;
    layer8_outputs(691) <= b;
    layer8_outputs(692) <= not a;
    layer8_outputs(693) <= a xor b;
    layer8_outputs(694) <= not (a xor b);
    layer8_outputs(695) <= not a;
    layer8_outputs(696) <= not a;
    layer8_outputs(697) <= a;
    layer8_outputs(698) <= a or b;
    layer8_outputs(699) <= a xor b;
    layer8_outputs(700) <= a xor b;
    layer8_outputs(701) <= not (a xor b);
    layer8_outputs(702) <= not (a or b);
    layer8_outputs(703) <= b;
    layer8_outputs(704) <= b;
    layer8_outputs(705) <= a xor b;
    layer8_outputs(706) <= a and not b;
    layer8_outputs(707) <= not a;
    layer8_outputs(708) <= not (a or b);
    layer8_outputs(709) <= not (a xor b);
    layer8_outputs(710) <= b;
    layer8_outputs(711) <= not b or a;
    layer8_outputs(712) <= a;
    layer8_outputs(713) <= not (a xor b);
    layer8_outputs(714) <= not (a or b);
    layer8_outputs(715) <= a;
    layer8_outputs(716) <= not a;
    layer8_outputs(717) <= not b;
    layer8_outputs(718) <= a;
    layer8_outputs(719) <= b;
    layer8_outputs(720) <= a or b;
    layer8_outputs(721) <= a xor b;
    layer8_outputs(722) <= not a or b;
    layer8_outputs(723) <= a and not b;
    layer8_outputs(724) <= not (a or b);
    layer8_outputs(725) <= a;
    layer8_outputs(726) <= b;
    layer8_outputs(727) <= b and not a;
    layer8_outputs(728) <= a xor b;
    layer8_outputs(729) <= not a;
    layer8_outputs(730) <= not (a or b);
    layer8_outputs(731) <= a;
    layer8_outputs(732) <= b;
    layer8_outputs(733) <= a or b;
    layer8_outputs(734) <= a;
    layer8_outputs(735) <= a or b;
    layer8_outputs(736) <= not b;
    layer8_outputs(737) <= not (a xor b);
    layer8_outputs(738) <= a;
    layer8_outputs(739) <= a xor b;
    layer8_outputs(740) <= a;
    layer8_outputs(741) <= not (a xor b);
    layer8_outputs(742) <= a xor b;
    layer8_outputs(743) <= not b or a;
    layer8_outputs(744) <= a;
    layer8_outputs(745) <= not b;
    layer8_outputs(746) <= a;
    layer8_outputs(747) <= not b;
    layer8_outputs(748) <= a xor b;
    layer8_outputs(749) <= a;
    layer8_outputs(750) <= a;
    layer8_outputs(751) <= a or b;
    layer8_outputs(752) <= not (a xor b);
    layer8_outputs(753) <= a;
    layer8_outputs(754) <= b;
    layer8_outputs(755) <= a and b;
    layer8_outputs(756) <= b;
    layer8_outputs(757) <= not b;
    layer8_outputs(758) <= not (a or b);
    layer8_outputs(759) <= not (a xor b);
    layer8_outputs(760) <= a xor b;
    layer8_outputs(761) <= b;
    layer8_outputs(762) <= not (a xor b);
    layer8_outputs(763) <= b;
    layer8_outputs(764) <= b;
    layer8_outputs(765) <= a or b;
    layer8_outputs(766) <= a or b;
    layer8_outputs(767) <= not a;
    layer8_outputs(768) <= a;
    layer8_outputs(769) <= a;
    layer8_outputs(770) <= not (a and b);
    layer8_outputs(771) <= not a;
    layer8_outputs(772) <= a xor b;
    layer8_outputs(773) <= not b;
    layer8_outputs(774) <= not b;
    layer8_outputs(775) <= not b;
    layer8_outputs(776) <= '1';
    layer8_outputs(777) <= not (a or b);
    layer8_outputs(778) <= a;
    layer8_outputs(779) <= a xor b;
    layer8_outputs(780) <= not (a or b);
    layer8_outputs(781) <= b;
    layer8_outputs(782) <= not a;
    layer8_outputs(783) <= not a;
    layer8_outputs(784) <= a and b;
    layer8_outputs(785) <= not a;
    layer8_outputs(786) <= a and not b;
    layer8_outputs(787) <= not (a xor b);
    layer8_outputs(788) <= not b;
    layer8_outputs(789) <= not b;
    layer8_outputs(790) <= b;
    layer8_outputs(791) <= a;
    layer8_outputs(792) <= not (a xor b);
    layer8_outputs(793) <= not a or b;
    layer8_outputs(794) <= a;
    layer8_outputs(795) <= not a;
    layer8_outputs(796) <= not (a xor b);
    layer8_outputs(797) <= not b;
    layer8_outputs(798) <= not (a or b);
    layer8_outputs(799) <= not a;
    layer8_outputs(800) <= b and not a;
    layer8_outputs(801) <= not a;
    layer8_outputs(802) <= a or b;
    layer8_outputs(803) <= a xor b;
    layer8_outputs(804) <= not b;
    layer8_outputs(805) <= not (a xor b);
    layer8_outputs(806) <= b;
    layer8_outputs(807) <= a and not b;
    layer8_outputs(808) <= not a;
    layer8_outputs(809) <= a xor b;
    layer8_outputs(810) <= not b;
    layer8_outputs(811) <= not b or a;
    layer8_outputs(812) <= not a;
    layer8_outputs(813) <= b;
    layer8_outputs(814) <= a and not b;
    layer8_outputs(815) <= a or b;
    layer8_outputs(816) <= not b;
    layer8_outputs(817) <= not a;
    layer8_outputs(818) <= a xor b;
    layer8_outputs(819) <= b and not a;
    layer8_outputs(820) <= not (a xor b);
    layer8_outputs(821) <= b;
    layer8_outputs(822) <= not b;
    layer8_outputs(823) <= not (a xor b);
    layer8_outputs(824) <= a and b;
    layer8_outputs(825) <= a and b;
    layer8_outputs(826) <= not a;
    layer8_outputs(827) <= not (a xor b);
    layer8_outputs(828) <= not (a xor b);
    layer8_outputs(829) <= not a;
    layer8_outputs(830) <= a xor b;
    layer8_outputs(831) <= not (a or b);
    layer8_outputs(832) <= not (a xor b);
    layer8_outputs(833) <= a;
    layer8_outputs(834) <= a;
    layer8_outputs(835) <= a and b;
    layer8_outputs(836) <= a or b;
    layer8_outputs(837) <= not (a xor b);
    layer8_outputs(838) <= a xor b;
    layer8_outputs(839) <= b;
    layer8_outputs(840) <= a and not b;
    layer8_outputs(841) <= a;
    layer8_outputs(842) <= not (a xor b);
    layer8_outputs(843) <= a and b;
    layer8_outputs(844) <= a xor b;
    layer8_outputs(845) <= not b;
    layer8_outputs(846) <= not a;
    layer8_outputs(847) <= not a;
    layer8_outputs(848) <= a and b;
    layer8_outputs(849) <= not b or a;
    layer8_outputs(850) <= b;
    layer8_outputs(851) <= a xor b;
    layer8_outputs(852) <= not b or a;
    layer8_outputs(853) <= not (a xor b);
    layer8_outputs(854) <= a;
    layer8_outputs(855) <= b and not a;
    layer8_outputs(856) <= a;
    layer8_outputs(857) <= not b;
    layer8_outputs(858) <= a xor b;
    layer8_outputs(859) <= a;
    layer8_outputs(860) <= not a;
    layer8_outputs(861) <= a and not b;
    layer8_outputs(862) <= a;
    layer8_outputs(863) <= a and b;
    layer8_outputs(864) <= a xor b;
    layer8_outputs(865) <= not (a xor b);
    layer8_outputs(866) <= a and b;
    layer8_outputs(867) <= b;
    layer8_outputs(868) <= a xor b;
    layer8_outputs(869) <= b;
    layer8_outputs(870) <= not b or a;
    layer8_outputs(871) <= not (a and b);
    layer8_outputs(872) <= a xor b;
    layer8_outputs(873) <= '1';
    layer8_outputs(874) <= not a;
    layer8_outputs(875) <= a;
    layer8_outputs(876) <= a xor b;
    layer8_outputs(877) <= b;
    layer8_outputs(878) <= a and b;
    layer8_outputs(879) <= not b;
    layer8_outputs(880) <= a xor b;
    layer8_outputs(881) <= a and b;
    layer8_outputs(882) <= not a or b;
    layer8_outputs(883) <= not (a and b);
    layer8_outputs(884) <= not (a and b);
    layer8_outputs(885) <= a or b;
    layer8_outputs(886) <= b and not a;
    layer8_outputs(887) <= not a;
    layer8_outputs(888) <= not (a and b);
    layer8_outputs(889) <= a;
    layer8_outputs(890) <= a xor b;
    layer8_outputs(891) <= a or b;
    layer8_outputs(892) <= b;
    layer8_outputs(893) <= not b;
    layer8_outputs(894) <= not (a xor b);
    layer8_outputs(895) <= not (a xor b);
    layer8_outputs(896) <= b;
    layer8_outputs(897) <= not a or b;
    layer8_outputs(898) <= a and not b;
    layer8_outputs(899) <= a or b;
    layer8_outputs(900) <= b;
    layer8_outputs(901) <= a;
    layer8_outputs(902) <= a;
    layer8_outputs(903) <= not (a and b);
    layer8_outputs(904) <= not (a and b);
    layer8_outputs(905) <= b;
    layer8_outputs(906) <= not a;
    layer8_outputs(907) <= b;
    layer8_outputs(908) <= a or b;
    layer8_outputs(909) <= a and not b;
    layer8_outputs(910) <= not a;
    layer8_outputs(911) <= not (a xor b);
    layer8_outputs(912) <= a;
    layer8_outputs(913) <= not (a xor b);
    layer8_outputs(914) <= b and not a;
    layer8_outputs(915) <= not a;
    layer8_outputs(916) <= a and b;
    layer8_outputs(917) <= not (a xor b);
    layer8_outputs(918) <= a;
    layer8_outputs(919) <= a;
    layer8_outputs(920) <= not (a and b);
    layer8_outputs(921) <= b;
    layer8_outputs(922) <= a;
    layer8_outputs(923) <= a and not b;
    layer8_outputs(924) <= a;
    layer8_outputs(925) <= b;
    layer8_outputs(926) <= a and b;
    layer8_outputs(927) <= a and not b;
    layer8_outputs(928) <= a;
    layer8_outputs(929) <= a and b;
    layer8_outputs(930) <= not b;
    layer8_outputs(931) <= not (a xor b);
    layer8_outputs(932) <= not b;
    layer8_outputs(933) <= not a or b;
    layer8_outputs(934) <= not (a xor b);
    layer8_outputs(935) <= not a or b;
    layer8_outputs(936) <= a xor b;
    layer8_outputs(937) <= not b or a;
    layer8_outputs(938) <= not a;
    layer8_outputs(939) <= not a;
    layer8_outputs(940) <= a xor b;
    layer8_outputs(941) <= not b;
    layer8_outputs(942) <= not a;
    layer8_outputs(943) <= a xor b;
    layer8_outputs(944) <= not b;
    layer8_outputs(945) <= a and not b;
    layer8_outputs(946) <= a xor b;
    layer8_outputs(947) <= not (a or b);
    layer8_outputs(948) <= b and not a;
    layer8_outputs(949) <= b;
    layer8_outputs(950) <= a;
    layer8_outputs(951) <= b;
    layer8_outputs(952) <= not b or a;
    layer8_outputs(953) <= not (a xor b);
    layer8_outputs(954) <= not (a and b);
    layer8_outputs(955) <= not b;
    layer8_outputs(956) <= b;
    layer8_outputs(957) <= not a;
    layer8_outputs(958) <= a xor b;
    layer8_outputs(959) <= not (a xor b);
    layer8_outputs(960) <= a xor b;
    layer8_outputs(961) <= not b;
    layer8_outputs(962) <= not (a xor b);
    layer8_outputs(963) <= a;
    layer8_outputs(964) <= not (a and b);
    layer8_outputs(965) <= a xor b;
    layer8_outputs(966) <= not a;
    layer8_outputs(967) <= a xor b;
    layer8_outputs(968) <= not (a xor b);
    layer8_outputs(969) <= a;
    layer8_outputs(970) <= a;
    layer8_outputs(971) <= a;
    layer8_outputs(972) <= a;
    layer8_outputs(973) <= a and not b;
    layer8_outputs(974) <= not a;
    layer8_outputs(975) <= not (a or b);
    layer8_outputs(976) <= not a;
    layer8_outputs(977) <= not b;
    layer8_outputs(978) <= a and not b;
    layer8_outputs(979) <= b;
    layer8_outputs(980) <= b and not a;
    layer8_outputs(981) <= not a or b;
    layer8_outputs(982) <= a and b;
    layer8_outputs(983) <= not (a and b);
    layer8_outputs(984) <= not a or b;
    layer8_outputs(985) <= a xor b;
    layer8_outputs(986) <= not (a and b);
    layer8_outputs(987) <= b and not a;
    layer8_outputs(988) <= not (a xor b);
    layer8_outputs(989) <= not a;
    layer8_outputs(990) <= not a or b;
    layer8_outputs(991) <= not b;
    layer8_outputs(992) <= a or b;
    layer8_outputs(993) <= b;
    layer8_outputs(994) <= b;
    layer8_outputs(995) <= not b or a;
    layer8_outputs(996) <= a and not b;
    layer8_outputs(997) <= b;
    layer8_outputs(998) <= a xor b;
    layer8_outputs(999) <= not b;
    layer8_outputs(1000) <= b;
    layer8_outputs(1001) <= not (a and b);
    layer8_outputs(1002) <= not b or a;
    layer8_outputs(1003) <= a xor b;
    layer8_outputs(1004) <= not b or a;
    layer8_outputs(1005) <= b and not a;
    layer8_outputs(1006) <= not (a or b);
    layer8_outputs(1007) <= not a;
    layer8_outputs(1008) <= not a or b;
    layer8_outputs(1009) <= not (a and b);
    layer8_outputs(1010) <= not b or a;
    layer8_outputs(1011) <= not b;
    layer8_outputs(1012) <= '1';
    layer8_outputs(1013) <= a;
    layer8_outputs(1014) <= not b;
    layer8_outputs(1015) <= b;
    layer8_outputs(1016) <= b;
    layer8_outputs(1017) <= a xor b;
    layer8_outputs(1018) <= '1';
    layer8_outputs(1019) <= not a;
    layer8_outputs(1020) <= not b;
    layer8_outputs(1021) <= a;
    layer8_outputs(1022) <= a and not b;
    layer8_outputs(1023) <= not (a and b);
    layer8_outputs(1024) <= not a or b;
    layer8_outputs(1025) <= a and b;
    layer8_outputs(1026) <= not (a xor b);
    layer8_outputs(1027) <= not a;
    layer8_outputs(1028) <= not a;
    layer8_outputs(1029) <= not (a xor b);
    layer8_outputs(1030) <= a;
    layer8_outputs(1031) <= not a or b;
    layer8_outputs(1032) <= not (a xor b);
    layer8_outputs(1033) <= not a;
    layer8_outputs(1034) <= not a or b;
    layer8_outputs(1035) <= a xor b;
    layer8_outputs(1036) <= b;
    layer8_outputs(1037) <= a or b;
    layer8_outputs(1038) <= b;
    layer8_outputs(1039) <= not b;
    layer8_outputs(1040) <= a;
    layer8_outputs(1041) <= not (a and b);
    layer8_outputs(1042) <= a;
    layer8_outputs(1043) <= not a;
    layer8_outputs(1044) <= a;
    layer8_outputs(1045) <= not a;
    layer8_outputs(1046) <= not a;
    layer8_outputs(1047) <= a;
    layer8_outputs(1048) <= not b or a;
    layer8_outputs(1049) <= not b;
    layer8_outputs(1050) <= not a;
    layer8_outputs(1051) <= not (a xor b);
    layer8_outputs(1052) <= a;
    layer8_outputs(1053) <= b;
    layer8_outputs(1054) <= not (a and b);
    layer8_outputs(1055) <= a;
    layer8_outputs(1056) <= b;
    layer8_outputs(1057) <= not a;
    layer8_outputs(1058) <= a and b;
    layer8_outputs(1059) <= a and b;
    layer8_outputs(1060) <= a and not b;
    layer8_outputs(1061) <= '0';
    layer8_outputs(1062) <= a or b;
    layer8_outputs(1063) <= a and not b;
    layer8_outputs(1064) <= a;
    layer8_outputs(1065) <= b;
    layer8_outputs(1066) <= a xor b;
    layer8_outputs(1067) <= not a;
    layer8_outputs(1068) <= not a or b;
    layer8_outputs(1069) <= not (a or b);
    layer8_outputs(1070) <= b;
    layer8_outputs(1071) <= a xor b;
    layer8_outputs(1072) <= b;
    layer8_outputs(1073) <= not a;
    layer8_outputs(1074) <= b;
    layer8_outputs(1075) <= a and not b;
    layer8_outputs(1076) <= a or b;
    layer8_outputs(1077) <= not (a xor b);
    layer8_outputs(1078) <= not (a xor b);
    layer8_outputs(1079) <= a xor b;
    layer8_outputs(1080) <= not b;
    layer8_outputs(1081) <= b;
    layer8_outputs(1082) <= a xor b;
    layer8_outputs(1083) <= a;
    layer8_outputs(1084) <= not b;
    layer8_outputs(1085) <= not b or a;
    layer8_outputs(1086) <= a xor b;
    layer8_outputs(1087) <= a xor b;
    layer8_outputs(1088) <= b;
    layer8_outputs(1089) <= not (a or b);
    layer8_outputs(1090) <= not b or a;
    layer8_outputs(1091) <= not a;
    layer8_outputs(1092) <= not a;
    layer8_outputs(1093) <= a xor b;
    layer8_outputs(1094) <= b;
    layer8_outputs(1095) <= a;
    layer8_outputs(1096) <= not (a and b);
    layer8_outputs(1097) <= not b or a;
    layer8_outputs(1098) <= not a;
    layer8_outputs(1099) <= not (a xor b);
    layer8_outputs(1100) <= a;
    layer8_outputs(1101) <= not (a xor b);
    layer8_outputs(1102) <= not b;
    layer8_outputs(1103) <= a or b;
    layer8_outputs(1104) <= not b or a;
    layer8_outputs(1105) <= not b;
    layer8_outputs(1106) <= not a;
    layer8_outputs(1107) <= a xor b;
    layer8_outputs(1108) <= not b or a;
    layer8_outputs(1109) <= b;
    layer8_outputs(1110) <= a and not b;
    layer8_outputs(1111) <= a xor b;
    layer8_outputs(1112) <= b;
    layer8_outputs(1113) <= a or b;
    layer8_outputs(1114) <= not b or a;
    layer8_outputs(1115) <= not (a xor b);
    layer8_outputs(1116) <= not (a or b);
    layer8_outputs(1117) <= not (a or b);
    layer8_outputs(1118) <= not (a and b);
    layer8_outputs(1119) <= a and b;
    layer8_outputs(1120) <= a xor b;
    layer8_outputs(1121) <= a or b;
    layer8_outputs(1122) <= not a;
    layer8_outputs(1123) <= not b or a;
    layer8_outputs(1124) <= not (a and b);
    layer8_outputs(1125) <= b and not a;
    layer8_outputs(1126) <= b;
    layer8_outputs(1127) <= b and not a;
    layer8_outputs(1128) <= a;
    layer8_outputs(1129) <= b;
    layer8_outputs(1130) <= a xor b;
    layer8_outputs(1131) <= a and not b;
    layer8_outputs(1132) <= a;
    layer8_outputs(1133) <= b;
    layer8_outputs(1134) <= a xor b;
    layer8_outputs(1135) <= a xor b;
    layer8_outputs(1136) <= b;
    layer8_outputs(1137) <= b;
    layer8_outputs(1138) <= not b;
    layer8_outputs(1139) <= a;
    layer8_outputs(1140) <= a;
    layer8_outputs(1141) <= not b or a;
    layer8_outputs(1142) <= not a;
    layer8_outputs(1143) <= not (a or b);
    layer8_outputs(1144) <= not b;
    layer8_outputs(1145) <= a and b;
    layer8_outputs(1146) <= b;
    layer8_outputs(1147) <= a xor b;
    layer8_outputs(1148) <= a xor b;
    layer8_outputs(1149) <= b and not a;
    layer8_outputs(1150) <= not a;
    layer8_outputs(1151) <= not b;
    layer8_outputs(1152) <= a;
    layer8_outputs(1153) <= a or b;
    layer8_outputs(1154) <= not a;
    layer8_outputs(1155) <= not b;
    layer8_outputs(1156) <= not a or b;
    layer8_outputs(1157) <= a;
    layer8_outputs(1158) <= not a or b;
    layer8_outputs(1159) <= b;
    layer8_outputs(1160) <= a xor b;
    layer8_outputs(1161) <= not b or a;
    layer8_outputs(1162) <= a;
    layer8_outputs(1163) <= a;
    layer8_outputs(1164) <= a or b;
    layer8_outputs(1165) <= a and not b;
    layer8_outputs(1166) <= b;
    layer8_outputs(1167) <= not b;
    layer8_outputs(1168) <= not (a or b);
    layer8_outputs(1169) <= b;
    layer8_outputs(1170) <= b;
    layer8_outputs(1171) <= a xor b;
    layer8_outputs(1172) <= not (a xor b);
    layer8_outputs(1173) <= b;
    layer8_outputs(1174) <= not a or b;
    layer8_outputs(1175) <= b;
    layer8_outputs(1176) <= a and not b;
    layer8_outputs(1177) <= not b;
    layer8_outputs(1178) <= b;
    layer8_outputs(1179) <= a xor b;
    layer8_outputs(1180) <= b;
    layer8_outputs(1181) <= not b or a;
    layer8_outputs(1182) <= not a or b;
    layer8_outputs(1183) <= a xor b;
    layer8_outputs(1184) <= b;
    layer8_outputs(1185) <= a and b;
    layer8_outputs(1186) <= not a;
    layer8_outputs(1187) <= not a;
    layer8_outputs(1188) <= '0';
    layer8_outputs(1189) <= a xor b;
    layer8_outputs(1190) <= not b;
    layer8_outputs(1191) <= b;
    layer8_outputs(1192) <= b;
    layer8_outputs(1193) <= a and b;
    layer8_outputs(1194) <= not (a and b);
    layer8_outputs(1195) <= not b;
    layer8_outputs(1196) <= not b;
    layer8_outputs(1197) <= a and b;
    layer8_outputs(1198) <= a;
    layer8_outputs(1199) <= not b;
    layer8_outputs(1200) <= not (a xor b);
    layer8_outputs(1201) <= b;
    layer8_outputs(1202) <= b;
    layer8_outputs(1203) <= not (a and b);
    layer8_outputs(1204) <= not (a xor b);
    layer8_outputs(1205) <= b;
    layer8_outputs(1206) <= not (a xor b);
    layer8_outputs(1207) <= a;
    layer8_outputs(1208) <= a;
    layer8_outputs(1209) <= a xor b;
    layer8_outputs(1210) <= not (a and b);
    layer8_outputs(1211) <= a xor b;
    layer8_outputs(1212) <= not a;
    layer8_outputs(1213) <= b;
    layer8_outputs(1214) <= a or b;
    layer8_outputs(1215) <= not (a and b);
    layer8_outputs(1216) <= not b;
    layer8_outputs(1217) <= a and b;
    layer8_outputs(1218) <= not a;
    layer8_outputs(1219) <= not (a xor b);
    layer8_outputs(1220) <= a;
    layer8_outputs(1221) <= a;
    layer8_outputs(1222) <= b;
    layer8_outputs(1223) <= a and not b;
    layer8_outputs(1224) <= a xor b;
    layer8_outputs(1225) <= a and b;
    layer8_outputs(1226) <= not b;
    layer8_outputs(1227) <= '1';
    layer8_outputs(1228) <= not b;
    layer8_outputs(1229) <= '0';
    layer8_outputs(1230) <= not b or a;
    layer8_outputs(1231) <= '1';
    layer8_outputs(1232) <= b;
    layer8_outputs(1233) <= a;
    layer8_outputs(1234) <= a and not b;
    layer8_outputs(1235) <= not a or b;
    layer8_outputs(1236) <= b;
    layer8_outputs(1237) <= not (a or b);
    layer8_outputs(1238) <= b;
    layer8_outputs(1239) <= b and not a;
    layer8_outputs(1240) <= not a or b;
    layer8_outputs(1241) <= not (a xor b);
    layer8_outputs(1242) <= a and not b;
    layer8_outputs(1243) <= not a;
    layer8_outputs(1244) <= not (a xor b);
    layer8_outputs(1245) <= not a;
    layer8_outputs(1246) <= not b;
    layer8_outputs(1247) <= not a;
    layer8_outputs(1248) <= not b;
    layer8_outputs(1249) <= not b;
    layer8_outputs(1250) <= a xor b;
    layer8_outputs(1251) <= not (a xor b);
    layer8_outputs(1252) <= not (a xor b);
    layer8_outputs(1253) <= not (a or b);
    layer8_outputs(1254) <= not (a or b);
    layer8_outputs(1255) <= not a;
    layer8_outputs(1256) <= a;
    layer8_outputs(1257) <= b;
    layer8_outputs(1258) <= b;
    layer8_outputs(1259) <= a and b;
    layer8_outputs(1260) <= b;
    layer8_outputs(1261) <= b;
    layer8_outputs(1262) <= a xor b;
    layer8_outputs(1263) <= not (a and b);
    layer8_outputs(1264) <= b;
    layer8_outputs(1265) <= a and not b;
    layer8_outputs(1266) <= not (a and b);
    layer8_outputs(1267) <= '1';
    layer8_outputs(1268) <= not a;
    layer8_outputs(1269) <= a and not b;
    layer8_outputs(1270) <= a;
    layer8_outputs(1271) <= a and b;
    layer8_outputs(1272) <= b;
    layer8_outputs(1273) <= not b;
    layer8_outputs(1274) <= a xor b;
    layer8_outputs(1275) <= a and not b;
    layer8_outputs(1276) <= not b;
    layer8_outputs(1277) <= b;
    layer8_outputs(1278) <= not (a xor b);
    layer8_outputs(1279) <= not (a xor b);
    layer8_outputs(1280) <= not b;
    layer8_outputs(1281) <= not a or b;
    layer8_outputs(1282) <= b and not a;
    layer8_outputs(1283) <= not a;
    layer8_outputs(1284) <= a xor b;
    layer8_outputs(1285) <= not a;
    layer8_outputs(1286) <= b;
    layer8_outputs(1287) <= a;
    layer8_outputs(1288) <= not a;
    layer8_outputs(1289) <= a;
    layer8_outputs(1290) <= not (a and b);
    layer8_outputs(1291) <= a xor b;
    layer8_outputs(1292) <= not (a xor b);
    layer8_outputs(1293) <= not (a and b);
    layer8_outputs(1294) <= not b;
    layer8_outputs(1295) <= not a;
    layer8_outputs(1296) <= not b;
    layer8_outputs(1297) <= a xor b;
    layer8_outputs(1298) <= not (a or b);
    layer8_outputs(1299) <= a;
    layer8_outputs(1300) <= not (a or b);
    layer8_outputs(1301) <= not (a and b);
    layer8_outputs(1302) <= not (a or b);
    layer8_outputs(1303) <= not (a or b);
    layer8_outputs(1304) <= '0';
    layer8_outputs(1305) <= a and b;
    layer8_outputs(1306) <= not (a xor b);
    layer8_outputs(1307) <= b;
    layer8_outputs(1308) <= b and not a;
    layer8_outputs(1309) <= not b;
    layer8_outputs(1310) <= not (a xor b);
    layer8_outputs(1311) <= not (a xor b);
    layer8_outputs(1312) <= not a or b;
    layer8_outputs(1313) <= a;
    layer8_outputs(1314) <= not b;
    layer8_outputs(1315) <= a or b;
    layer8_outputs(1316) <= b and not a;
    layer8_outputs(1317) <= not b or a;
    layer8_outputs(1318) <= b;
    layer8_outputs(1319) <= a xor b;
    layer8_outputs(1320) <= not b or a;
    layer8_outputs(1321) <= a;
    layer8_outputs(1322) <= not (a xor b);
    layer8_outputs(1323) <= a;
    layer8_outputs(1324) <= not (a or b);
    layer8_outputs(1325) <= not a;
    layer8_outputs(1326) <= not (a and b);
    layer8_outputs(1327) <= not a;
    layer8_outputs(1328) <= not b;
    layer8_outputs(1329) <= a xor b;
    layer8_outputs(1330) <= not b;
    layer8_outputs(1331) <= a;
    layer8_outputs(1332) <= a and not b;
    layer8_outputs(1333) <= '1';
    layer8_outputs(1334) <= b;
    layer8_outputs(1335) <= not b;
    layer8_outputs(1336) <= a xor b;
    layer8_outputs(1337) <= not (a and b);
    layer8_outputs(1338) <= a and not b;
    layer8_outputs(1339) <= not a;
    layer8_outputs(1340) <= not (a or b);
    layer8_outputs(1341) <= not b;
    layer8_outputs(1342) <= not (a and b);
    layer8_outputs(1343) <= a and not b;
    layer8_outputs(1344) <= a and b;
    layer8_outputs(1345) <= not b;
    layer8_outputs(1346) <= '1';
    layer8_outputs(1347) <= not a;
    layer8_outputs(1348) <= not a or b;
    layer8_outputs(1349) <= not b;
    layer8_outputs(1350) <= not (a xor b);
    layer8_outputs(1351) <= not (a xor b);
    layer8_outputs(1352) <= not a;
    layer8_outputs(1353) <= a xor b;
    layer8_outputs(1354) <= not a or b;
    layer8_outputs(1355) <= a;
    layer8_outputs(1356) <= b;
    layer8_outputs(1357) <= a xor b;
    layer8_outputs(1358) <= not a;
    layer8_outputs(1359) <= a xor b;
    layer8_outputs(1360) <= a or b;
    layer8_outputs(1361) <= not b;
    layer8_outputs(1362) <= not b;
    layer8_outputs(1363) <= a and not b;
    layer8_outputs(1364) <= not (a xor b);
    layer8_outputs(1365) <= a or b;
    layer8_outputs(1366) <= a;
    layer8_outputs(1367) <= a and not b;
    layer8_outputs(1368) <= not (a xor b);
    layer8_outputs(1369) <= a;
    layer8_outputs(1370) <= not a or b;
    layer8_outputs(1371) <= not a;
    layer8_outputs(1372) <= b;
    layer8_outputs(1373) <= b and not a;
    layer8_outputs(1374) <= not a;
    layer8_outputs(1375) <= not a;
    layer8_outputs(1376) <= b and not a;
    layer8_outputs(1377) <= a;
    layer8_outputs(1378) <= not a;
    layer8_outputs(1379) <= a;
    layer8_outputs(1380) <= b;
    layer8_outputs(1381) <= a;
    layer8_outputs(1382) <= a and not b;
    layer8_outputs(1383) <= not a;
    layer8_outputs(1384) <= a xor b;
    layer8_outputs(1385) <= a;
    layer8_outputs(1386) <= a and b;
    layer8_outputs(1387) <= not b;
    layer8_outputs(1388) <= not (a and b);
    layer8_outputs(1389) <= '0';
    layer8_outputs(1390) <= not b or a;
    layer8_outputs(1391) <= b;
    layer8_outputs(1392) <= a xor b;
    layer8_outputs(1393) <= not a;
    layer8_outputs(1394) <= not (a or b);
    layer8_outputs(1395) <= not a or b;
    layer8_outputs(1396) <= a and b;
    layer8_outputs(1397) <= not (a xor b);
    layer8_outputs(1398) <= b;
    layer8_outputs(1399) <= b;
    layer8_outputs(1400) <= b;
    layer8_outputs(1401) <= not a;
    layer8_outputs(1402) <= not b;
    layer8_outputs(1403) <= a xor b;
    layer8_outputs(1404) <= not b;
    layer8_outputs(1405) <= a and not b;
    layer8_outputs(1406) <= not (a xor b);
    layer8_outputs(1407) <= b;
    layer8_outputs(1408) <= '1';
    layer8_outputs(1409) <= b and not a;
    layer8_outputs(1410) <= b and not a;
    layer8_outputs(1411) <= not b;
    layer8_outputs(1412) <= a xor b;
    layer8_outputs(1413) <= not b;
    layer8_outputs(1414) <= a;
    layer8_outputs(1415) <= not a;
    layer8_outputs(1416) <= a or b;
    layer8_outputs(1417) <= a xor b;
    layer8_outputs(1418) <= b;
    layer8_outputs(1419) <= a xor b;
    layer8_outputs(1420) <= a and not b;
    layer8_outputs(1421) <= a xor b;
    layer8_outputs(1422) <= not (a and b);
    layer8_outputs(1423) <= a;
    layer8_outputs(1424) <= not b or a;
    layer8_outputs(1425) <= not a;
    layer8_outputs(1426) <= not a;
    layer8_outputs(1427) <= not a;
    layer8_outputs(1428) <= not (a and b);
    layer8_outputs(1429) <= a and b;
    layer8_outputs(1430) <= not b;
    layer8_outputs(1431) <= not a;
    layer8_outputs(1432) <= not (a xor b);
    layer8_outputs(1433) <= not a;
    layer8_outputs(1434) <= not (a and b);
    layer8_outputs(1435) <= b;
    layer8_outputs(1436) <= a;
    layer8_outputs(1437) <= not b;
    layer8_outputs(1438) <= a xor b;
    layer8_outputs(1439) <= not (a xor b);
    layer8_outputs(1440) <= not a;
    layer8_outputs(1441) <= a xor b;
    layer8_outputs(1442) <= a;
    layer8_outputs(1443) <= a or b;
    layer8_outputs(1444) <= a xor b;
    layer8_outputs(1445) <= a and b;
    layer8_outputs(1446) <= b and not a;
    layer8_outputs(1447) <= not (a and b);
    layer8_outputs(1448) <= not (a xor b);
    layer8_outputs(1449) <= a xor b;
    layer8_outputs(1450) <= a xor b;
    layer8_outputs(1451) <= b;
    layer8_outputs(1452) <= not b;
    layer8_outputs(1453) <= not b;
    layer8_outputs(1454) <= not a;
    layer8_outputs(1455) <= a;
    layer8_outputs(1456) <= a and b;
    layer8_outputs(1457) <= not a or b;
    layer8_outputs(1458) <= not a;
    layer8_outputs(1459) <= not a;
    layer8_outputs(1460) <= b and not a;
    layer8_outputs(1461) <= not (a or b);
    layer8_outputs(1462) <= a xor b;
    layer8_outputs(1463) <= not b or a;
    layer8_outputs(1464) <= not b or a;
    layer8_outputs(1465) <= not b;
    layer8_outputs(1466) <= not (a xor b);
    layer8_outputs(1467) <= not (a xor b);
    layer8_outputs(1468) <= not (a or b);
    layer8_outputs(1469) <= not b;
    layer8_outputs(1470) <= not (a or b);
    layer8_outputs(1471) <= not a;
    layer8_outputs(1472) <= b and not a;
    layer8_outputs(1473) <= not b;
    layer8_outputs(1474) <= a;
    layer8_outputs(1475) <= a xor b;
    layer8_outputs(1476) <= not (a xor b);
    layer8_outputs(1477) <= not b or a;
    layer8_outputs(1478) <= not b;
    layer8_outputs(1479) <= a;
    layer8_outputs(1480) <= not (a xor b);
    layer8_outputs(1481) <= not (a xor b);
    layer8_outputs(1482) <= not b;
    layer8_outputs(1483) <= not b;
    layer8_outputs(1484) <= not (a and b);
    layer8_outputs(1485) <= not (a or b);
    layer8_outputs(1486) <= b;
    layer8_outputs(1487) <= not a;
    layer8_outputs(1488) <= b;
    layer8_outputs(1489) <= b;
    layer8_outputs(1490) <= a xor b;
    layer8_outputs(1491) <= a;
    layer8_outputs(1492) <= a xor b;
    layer8_outputs(1493) <= a and not b;
    layer8_outputs(1494) <= not a;
    layer8_outputs(1495) <= b;
    layer8_outputs(1496) <= b;
    layer8_outputs(1497) <= a xor b;
    layer8_outputs(1498) <= not a;
    layer8_outputs(1499) <= not a;
    layer8_outputs(1500) <= not b or a;
    layer8_outputs(1501) <= not a;
    layer8_outputs(1502) <= not (a xor b);
    layer8_outputs(1503) <= not b;
    layer8_outputs(1504) <= b;
    layer8_outputs(1505) <= b and not a;
    layer8_outputs(1506) <= a xor b;
    layer8_outputs(1507) <= b;
    layer8_outputs(1508) <= b;
    layer8_outputs(1509) <= not a;
    layer8_outputs(1510) <= not b;
    layer8_outputs(1511) <= b;
    layer8_outputs(1512) <= b;
    layer8_outputs(1513) <= a and b;
    layer8_outputs(1514) <= not b;
    layer8_outputs(1515) <= not a or b;
    layer8_outputs(1516) <= not a;
    layer8_outputs(1517) <= not (a xor b);
    layer8_outputs(1518) <= not (a or b);
    layer8_outputs(1519) <= a;
    layer8_outputs(1520) <= not (a xor b);
    layer8_outputs(1521) <= not a;
    layer8_outputs(1522) <= not a;
    layer8_outputs(1523) <= a and not b;
    layer8_outputs(1524) <= not (a xor b);
    layer8_outputs(1525) <= a xor b;
    layer8_outputs(1526) <= not a;
    layer8_outputs(1527) <= a and not b;
    layer8_outputs(1528) <= a and not b;
    layer8_outputs(1529) <= not (a or b);
    layer8_outputs(1530) <= a xor b;
    layer8_outputs(1531) <= not (a and b);
    layer8_outputs(1532) <= a;
    layer8_outputs(1533) <= not (a and b);
    layer8_outputs(1534) <= a and b;
    layer8_outputs(1535) <= b;
    layer8_outputs(1536) <= a or b;
    layer8_outputs(1537) <= b;
    layer8_outputs(1538) <= a;
    layer8_outputs(1539) <= not (a and b);
    layer8_outputs(1540) <= b and not a;
    layer8_outputs(1541) <= not a or b;
    layer8_outputs(1542) <= a;
    layer8_outputs(1543) <= not b;
    layer8_outputs(1544) <= a;
    layer8_outputs(1545) <= a and not b;
    layer8_outputs(1546) <= not (a xor b);
    layer8_outputs(1547) <= not b;
    layer8_outputs(1548) <= a;
    layer8_outputs(1549) <= not b or a;
    layer8_outputs(1550) <= a;
    layer8_outputs(1551) <= a xor b;
    layer8_outputs(1552) <= not a;
    layer8_outputs(1553) <= not a;
    layer8_outputs(1554) <= a xor b;
    layer8_outputs(1555) <= not a;
    layer8_outputs(1556) <= b and not a;
    layer8_outputs(1557) <= not (a xor b);
    layer8_outputs(1558) <= not (a xor b);
    layer8_outputs(1559) <= a xor b;
    layer8_outputs(1560) <= b;
    layer8_outputs(1561) <= b;
    layer8_outputs(1562) <= not (a xor b);
    layer8_outputs(1563) <= not b;
    layer8_outputs(1564) <= not (a or b);
    layer8_outputs(1565) <= not a or b;
    layer8_outputs(1566) <= not (a xor b);
    layer8_outputs(1567) <= not b;
    layer8_outputs(1568) <= b and not a;
    layer8_outputs(1569) <= not b;
    layer8_outputs(1570) <= not a;
    layer8_outputs(1571) <= a xor b;
    layer8_outputs(1572) <= a xor b;
    layer8_outputs(1573) <= not (a xor b);
    layer8_outputs(1574) <= not (a xor b);
    layer8_outputs(1575) <= not b;
    layer8_outputs(1576) <= not a or b;
    layer8_outputs(1577) <= a xor b;
    layer8_outputs(1578) <= b and not a;
    layer8_outputs(1579) <= b;
    layer8_outputs(1580) <= not (a xor b);
    layer8_outputs(1581) <= not b or a;
    layer8_outputs(1582) <= not a;
    layer8_outputs(1583) <= not a;
    layer8_outputs(1584) <= not (a or b);
    layer8_outputs(1585) <= not (a xor b);
    layer8_outputs(1586) <= a or b;
    layer8_outputs(1587) <= a and b;
    layer8_outputs(1588) <= a xor b;
    layer8_outputs(1589) <= a and b;
    layer8_outputs(1590) <= not b or a;
    layer8_outputs(1591) <= not (a xor b);
    layer8_outputs(1592) <= a xor b;
    layer8_outputs(1593) <= not (a xor b);
    layer8_outputs(1594) <= a xor b;
    layer8_outputs(1595) <= not b or a;
    layer8_outputs(1596) <= a;
    layer8_outputs(1597) <= b;
    layer8_outputs(1598) <= b;
    layer8_outputs(1599) <= not a;
    layer8_outputs(1600) <= not b;
    layer8_outputs(1601) <= not b or a;
    layer8_outputs(1602) <= a;
    layer8_outputs(1603) <= a;
    layer8_outputs(1604) <= b and not a;
    layer8_outputs(1605) <= a or b;
    layer8_outputs(1606) <= not a;
    layer8_outputs(1607) <= a;
    layer8_outputs(1608) <= b;
    layer8_outputs(1609) <= not a;
    layer8_outputs(1610) <= not a;
    layer8_outputs(1611) <= not a;
    layer8_outputs(1612) <= not a;
    layer8_outputs(1613) <= a and not b;
    layer8_outputs(1614) <= not b or a;
    layer8_outputs(1615) <= not (a or b);
    layer8_outputs(1616) <= not (a or b);
    layer8_outputs(1617) <= not a or b;
    layer8_outputs(1618) <= b;
    layer8_outputs(1619) <= a or b;
    layer8_outputs(1620) <= a xor b;
    layer8_outputs(1621) <= not b;
    layer8_outputs(1622) <= b and not a;
    layer8_outputs(1623) <= not b;
    layer8_outputs(1624) <= not b;
    layer8_outputs(1625) <= a;
    layer8_outputs(1626) <= b;
    layer8_outputs(1627) <= not (a xor b);
    layer8_outputs(1628) <= a or b;
    layer8_outputs(1629) <= not b;
    layer8_outputs(1630) <= a xor b;
    layer8_outputs(1631) <= not a or b;
    layer8_outputs(1632) <= a;
    layer8_outputs(1633) <= not b or a;
    layer8_outputs(1634) <= not b;
    layer8_outputs(1635) <= not b or a;
    layer8_outputs(1636) <= not a;
    layer8_outputs(1637) <= not (a and b);
    layer8_outputs(1638) <= a or b;
    layer8_outputs(1639) <= b and not a;
    layer8_outputs(1640) <= a or b;
    layer8_outputs(1641) <= not b;
    layer8_outputs(1642) <= not (a or b);
    layer8_outputs(1643) <= not a;
    layer8_outputs(1644) <= a and not b;
    layer8_outputs(1645) <= a xor b;
    layer8_outputs(1646) <= not a;
    layer8_outputs(1647) <= not a;
    layer8_outputs(1648) <= not (a xor b);
    layer8_outputs(1649) <= a;
    layer8_outputs(1650) <= not a;
    layer8_outputs(1651) <= b;
    layer8_outputs(1652) <= not (a or b);
    layer8_outputs(1653) <= not (a xor b);
    layer8_outputs(1654) <= a xor b;
    layer8_outputs(1655) <= a;
    layer8_outputs(1656) <= not (a xor b);
    layer8_outputs(1657) <= not b;
    layer8_outputs(1658) <= b and not a;
    layer8_outputs(1659) <= a;
    layer8_outputs(1660) <= a;
    layer8_outputs(1661) <= a and b;
    layer8_outputs(1662) <= not (a or b);
    layer8_outputs(1663) <= not (a and b);
    layer8_outputs(1664) <= a and not b;
    layer8_outputs(1665) <= a xor b;
    layer8_outputs(1666) <= not a or b;
    layer8_outputs(1667) <= not a;
    layer8_outputs(1668) <= a;
    layer8_outputs(1669) <= not b;
    layer8_outputs(1670) <= not (a or b);
    layer8_outputs(1671) <= b and not a;
    layer8_outputs(1672) <= '0';
    layer8_outputs(1673) <= not b;
    layer8_outputs(1674) <= a or b;
    layer8_outputs(1675) <= a xor b;
    layer8_outputs(1676) <= a;
    layer8_outputs(1677) <= '1';
    layer8_outputs(1678) <= not (a xor b);
    layer8_outputs(1679) <= a xor b;
    layer8_outputs(1680) <= a xor b;
    layer8_outputs(1681) <= a and not b;
    layer8_outputs(1682) <= a and not b;
    layer8_outputs(1683) <= a and not b;
    layer8_outputs(1684) <= b;
    layer8_outputs(1685) <= not b;
    layer8_outputs(1686) <= a or b;
    layer8_outputs(1687) <= not b;
    layer8_outputs(1688) <= a and b;
    layer8_outputs(1689) <= not a or b;
    layer8_outputs(1690) <= not b;
    layer8_outputs(1691) <= not (a xor b);
    layer8_outputs(1692) <= a and b;
    layer8_outputs(1693) <= a and b;
    layer8_outputs(1694) <= not b or a;
    layer8_outputs(1695) <= not (a xor b);
    layer8_outputs(1696) <= not (a xor b);
    layer8_outputs(1697) <= not (a xor b);
    layer8_outputs(1698) <= a or b;
    layer8_outputs(1699) <= a xor b;
    layer8_outputs(1700) <= b;
    layer8_outputs(1701) <= b;
    layer8_outputs(1702) <= not (a xor b);
    layer8_outputs(1703) <= not (a xor b);
    layer8_outputs(1704) <= not (a or b);
    layer8_outputs(1705) <= not (a xor b);
    layer8_outputs(1706) <= a;
    layer8_outputs(1707) <= b;
    layer8_outputs(1708) <= not b or a;
    layer8_outputs(1709) <= not (a and b);
    layer8_outputs(1710) <= a and not b;
    layer8_outputs(1711) <= a and b;
    layer8_outputs(1712) <= not a;
    layer8_outputs(1713) <= not a;
    layer8_outputs(1714) <= b;
    layer8_outputs(1715) <= not a;
    layer8_outputs(1716) <= b;
    layer8_outputs(1717) <= not (a xor b);
    layer8_outputs(1718) <= not (a xor b);
    layer8_outputs(1719) <= not a or b;
    layer8_outputs(1720) <= b;
    layer8_outputs(1721) <= not (a xor b);
    layer8_outputs(1722) <= a xor b;
    layer8_outputs(1723) <= a and not b;
    layer8_outputs(1724) <= not (a or b);
    layer8_outputs(1725) <= not a or b;
    layer8_outputs(1726) <= b;
    layer8_outputs(1727) <= b;
    layer8_outputs(1728) <= b and not a;
    layer8_outputs(1729) <= not (a xor b);
    layer8_outputs(1730) <= not (a or b);
    layer8_outputs(1731) <= a xor b;
    layer8_outputs(1732) <= '1';
    layer8_outputs(1733) <= not (a xor b);
    layer8_outputs(1734) <= a and b;
    layer8_outputs(1735) <= b;
    layer8_outputs(1736) <= a;
    layer8_outputs(1737) <= not (a and b);
    layer8_outputs(1738) <= not (a or b);
    layer8_outputs(1739) <= not b;
    layer8_outputs(1740) <= not b;
    layer8_outputs(1741) <= not b;
    layer8_outputs(1742) <= a xor b;
    layer8_outputs(1743) <= a;
    layer8_outputs(1744) <= a xor b;
    layer8_outputs(1745) <= not b;
    layer8_outputs(1746) <= a xor b;
    layer8_outputs(1747) <= not (a xor b);
    layer8_outputs(1748) <= b;
    layer8_outputs(1749) <= b and not a;
    layer8_outputs(1750) <= '1';
    layer8_outputs(1751) <= a;
    layer8_outputs(1752) <= not (a or b);
    layer8_outputs(1753) <= b and not a;
    layer8_outputs(1754) <= not b;
    layer8_outputs(1755) <= not (a or b);
    layer8_outputs(1756) <= not a;
    layer8_outputs(1757) <= a;
    layer8_outputs(1758) <= not (a and b);
    layer8_outputs(1759) <= a;
    layer8_outputs(1760) <= not b;
    layer8_outputs(1761) <= a;
    layer8_outputs(1762) <= not b;
    layer8_outputs(1763) <= not (a and b);
    layer8_outputs(1764) <= a xor b;
    layer8_outputs(1765) <= not a;
    layer8_outputs(1766) <= not a or b;
    layer8_outputs(1767) <= not (a xor b);
    layer8_outputs(1768) <= not (a xor b);
    layer8_outputs(1769) <= b;
    layer8_outputs(1770) <= not (a or b);
    layer8_outputs(1771) <= not (a and b);
    layer8_outputs(1772) <= a;
    layer8_outputs(1773) <= a;
    layer8_outputs(1774) <= b and not a;
    layer8_outputs(1775) <= a xor b;
    layer8_outputs(1776) <= b and not a;
    layer8_outputs(1777) <= a;
    layer8_outputs(1778) <= not b or a;
    layer8_outputs(1779) <= a and b;
    layer8_outputs(1780) <= not (a and b);
    layer8_outputs(1781) <= not b;
    layer8_outputs(1782) <= not a;
    layer8_outputs(1783) <= b and not a;
    layer8_outputs(1784) <= not (a and b);
    layer8_outputs(1785) <= not (a or b);
    layer8_outputs(1786) <= not (a xor b);
    layer8_outputs(1787) <= not (a or b);
    layer8_outputs(1788) <= not (a or b);
    layer8_outputs(1789) <= not b;
    layer8_outputs(1790) <= not b;
    layer8_outputs(1791) <= '1';
    layer8_outputs(1792) <= not (a or b);
    layer8_outputs(1793) <= not (a or b);
    layer8_outputs(1794) <= a and b;
    layer8_outputs(1795) <= not a;
    layer8_outputs(1796) <= a and b;
    layer8_outputs(1797) <= a;
    layer8_outputs(1798) <= not b or a;
    layer8_outputs(1799) <= not a;
    layer8_outputs(1800) <= not b or a;
    layer8_outputs(1801) <= not b;
    layer8_outputs(1802) <= a and not b;
    layer8_outputs(1803) <= not (a xor b);
    layer8_outputs(1804) <= a and b;
    layer8_outputs(1805) <= a xor b;
    layer8_outputs(1806) <= a and not b;
    layer8_outputs(1807) <= not a;
    layer8_outputs(1808) <= a;
    layer8_outputs(1809) <= a xor b;
    layer8_outputs(1810) <= a;
    layer8_outputs(1811) <= not a or b;
    layer8_outputs(1812) <= b;
    layer8_outputs(1813) <= a and b;
    layer8_outputs(1814) <= not (a and b);
    layer8_outputs(1815) <= not a or b;
    layer8_outputs(1816) <= b;
    layer8_outputs(1817) <= b;
    layer8_outputs(1818) <= not (a xor b);
    layer8_outputs(1819) <= b;
    layer8_outputs(1820) <= b;
    layer8_outputs(1821) <= not b;
    layer8_outputs(1822) <= a;
    layer8_outputs(1823) <= b and not a;
    layer8_outputs(1824) <= b;
    layer8_outputs(1825) <= a;
    layer8_outputs(1826) <= b;
    layer8_outputs(1827) <= not b;
    layer8_outputs(1828) <= a and not b;
    layer8_outputs(1829) <= a xor b;
    layer8_outputs(1830) <= a xor b;
    layer8_outputs(1831) <= a;
    layer8_outputs(1832) <= a and not b;
    layer8_outputs(1833) <= not b;
    layer8_outputs(1834) <= not (a and b);
    layer8_outputs(1835) <= not (a xor b);
    layer8_outputs(1836) <= a xor b;
    layer8_outputs(1837) <= a and b;
    layer8_outputs(1838) <= a;
    layer8_outputs(1839) <= not a;
    layer8_outputs(1840) <= a;
    layer8_outputs(1841) <= a;
    layer8_outputs(1842) <= b;
    layer8_outputs(1843) <= not (a xor b);
    layer8_outputs(1844) <= not (a xor b);
    layer8_outputs(1845) <= not (a xor b);
    layer8_outputs(1846) <= not (a xor b);
    layer8_outputs(1847) <= b and not a;
    layer8_outputs(1848) <= not b;
    layer8_outputs(1849) <= b and not a;
    layer8_outputs(1850) <= not a;
    layer8_outputs(1851) <= not a;
    layer8_outputs(1852) <= not (a or b);
    layer8_outputs(1853) <= a;
    layer8_outputs(1854) <= a and b;
    layer8_outputs(1855) <= not (a xor b);
    layer8_outputs(1856) <= a xor b;
    layer8_outputs(1857) <= a xor b;
    layer8_outputs(1858) <= a or b;
    layer8_outputs(1859) <= a or b;
    layer8_outputs(1860) <= a or b;
    layer8_outputs(1861) <= not (a xor b);
    layer8_outputs(1862) <= not a or b;
    layer8_outputs(1863) <= b;
    layer8_outputs(1864) <= a or b;
    layer8_outputs(1865) <= not a;
    layer8_outputs(1866) <= not a or b;
    layer8_outputs(1867) <= b;
    layer8_outputs(1868) <= not b;
    layer8_outputs(1869) <= not a;
    layer8_outputs(1870) <= not a;
    layer8_outputs(1871) <= b and not a;
    layer8_outputs(1872) <= '1';
    layer8_outputs(1873) <= a and b;
    layer8_outputs(1874) <= not a or b;
    layer8_outputs(1875) <= a and b;
    layer8_outputs(1876) <= not b or a;
    layer8_outputs(1877) <= not (a or b);
    layer8_outputs(1878) <= a;
    layer8_outputs(1879) <= a xor b;
    layer8_outputs(1880) <= a and not b;
    layer8_outputs(1881) <= a;
    layer8_outputs(1882) <= a;
    layer8_outputs(1883) <= not (a xor b);
    layer8_outputs(1884) <= a and not b;
    layer8_outputs(1885) <= b and not a;
    layer8_outputs(1886) <= b;
    layer8_outputs(1887) <= not b or a;
    layer8_outputs(1888) <= b;
    layer8_outputs(1889) <= not b;
    layer8_outputs(1890) <= a;
    layer8_outputs(1891) <= not b or a;
    layer8_outputs(1892) <= a and not b;
    layer8_outputs(1893) <= a and not b;
    layer8_outputs(1894) <= a;
    layer8_outputs(1895) <= b and not a;
    layer8_outputs(1896) <= a;
    layer8_outputs(1897) <= not b;
    layer8_outputs(1898) <= a xor b;
    layer8_outputs(1899) <= not a or b;
    layer8_outputs(1900) <= not a;
    layer8_outputs(1901) <= b;
    layer8_outputs(1902) <= b;
    layer8_outputs(1903) <= not b or a;
    layer8_outputs(1904) <= a;
    layer8_outputs(1905) <= a xor b;
    layer8_outputs(1906) <= a;
    layer8_outputs(1907) <= b;
    layer8_outputs(1908) <= not (a xor b);
    layer8_outputs(1909) <= not b;
    layer8_outputs(1910) <= a;
    layer8_outputs(1911) <= a;
    layer8_outputs(1912) <= not (a xor b);
    layer8_outputs(1913) <= not (a and b);
    layer8_outputs(1914) <= a;
    layer8_outputs(1915) <= not (a xor b);
    layer8_outputs(1916) <= not a;
    layer8_outputs(1917) <= b and not a;
    layer8_outputs(1918) <= a xor b;
    layer8_outputs(1919) <= not b;
    layer8_outputs(1920) <= a;
    layer8_outputs(1921) <= b;
    layer8_outputs(1922) <= a and b;
    layer8_outputs(1923) <= b;
    layer8_outputs(1924) <= b and not a;
    layer8_outputs(1925) <= not (a or b);
    layer8_outputs(1926) <= not a;
    layer8_outputs(1927) <= not b;
    layer8_outputs(1928) <= not b;
    layer8_outputs(1929) <= a;
    layer8_outputs(1930) <= not b;
    layer8_outputs(1931) <= not (a and b);
    layer8_outputs(1932) <= not b;
    layer8_outputs(1933) <= not b;
    layer8_outputs(1934) <= not (a and b);
    layer8_outputs(1935) <= b and not a;
    layer8_outputs(1936) <= a and b;
    layer8_outputs(1937) <= not b or a;
    layer8_outputs(1938) <= a;
    layer8_outputs(1939) <= not (a xor b);
    layer8_outputs(1940) <= not b;
    layer8_outputs(1941) <= not (a xor b);
    layer8_outputs(1942) <= a xor b;
    layer8_outputs(1943) <= not a or b;
    layer8_outputs(1944) <= not (a or b);
    layer8_outputs(1945) <= not a;
    layer8_outputs(1946) <= not b;
    layer8_outputs(1947) <= not a or b;
    layer8_outputs(1948) <= a xor b;
    layer8_outputs(1949) <= not a;
    layer8_outputs(1950) <= a xor b;
    layer8_outputs(1951) <= a;
    layer8_outputs(1952) <= not (a and b);
    layer8_outputs(1953) <= not a or b;
    layer8_outputs(1954) <= not b or a;
    layer8_outputs(1955) <= not (a and b);
    layer8_outputs(1956) <= a xor b;
    layer8_outputs(1957) <= not b;
    layer8_outputs(1958) <= a xor b;
    layer8_outputs(1959) <= not a or b;
    layer8_outputs(1960) <= a or b;
    layer8_outputs(1961) <= a or b;
    layer8_outputs(1962) <= not b or a;
    layer8_outputs(1963) <= a and b;
    layer8_outputs(1964) <= b and not a;
    layer8_outputs(1965) <= a;
    layer8_outputs(1966) <= not (a or b);
    layer8_outputs(1967) <= a;
    layer8_outputs(1968) <= a and not b;
    layer8_outputs(1969) <= not b or a;
    layer8_outputs(1970) <= not a or b;
    layer8_outputs(1971) <= a or b;
    layer8_outputs(1972) <= not (a xor b);
    layer8_outputs(1973) <= a;
    layer8_outputs(1974) <= not b or a;
    layer8_outputs(1975) <= a or b;
    layer8_outputs(1976) <= a and b;
    layer8_outputs(1977) <= not a or b;
    layer8_outputs(1978) <= a and not b;
    layer8_outputs(1979) <= not b;
    layer8_outputs(1980) <= not b or a;
    layer8_outputs(1981) <= a xor b;
    layer8_outputs(1982) <= a;
    layer8_outputs(1983) <= not b;
    layer8_outputs(1984) <= not (a or b);
    layer8_outputs(1985) <= b;
    layer8_outputs(1986) <= not (a and b);
    layer8_outputs(1987) <= not (a xor b);
    layer8_outputs(1988) <= not a;
    layer8_outputs(1989) <= a xor b;
    layer8_outputs(1990) <= not (a xor b);
    layer8_outputs(1991) <= not a or b;
    layer8_outputs(1992) <= not (a or b);
    layer8_outputs(1993) <= not (a xor b);
    layer8_outputs(1994) <= a and not b;
    layer8_outputs(1995) <= not a;
    layer8_outputs(1996) <= a;
    layer8_outputs(1997) <= not a;
    layer8_outputs(1998) <= a and b;
    layer8_outputs(1999) <= not b;
    layer8_outputs(2000) <= b and not a;
    layer8_outputs(2001) <= not b;
    layer8_outputs(2002) <= not b or a;
    layer8_outputs(2003) <= not a;
    layer8_outputs(2004) <= not (a and b);
    layer8_outputs(2005) <= not b;
    layer8_outputs(2006) <= a xor b;
    layer8_outputs(2007) <= not b;
    layer8_outputs(2008) <= a;
    layer8_outputs(2009) <= a and not b;
    layer8_outputs(2010) <= b;
    layer8_outputs(2011) <= a;
    layer8_outputs(2012) <= a;
    layer8_outputs(2013) <= not a;
    layer8_outputs(2014) <= not b or a;
    layer8_outputs(2015) <= a and b;
    layer8_outputs(2016) <= not a or b;
    layer8_outputs(2017) <= not (a and b);
    layer8_outputs(2018) <= not (a or b);
    layer8_outputs(2019) <= not a;
    layer8_outputs(2020) <= a xor b;
    layer8_outputs(2021) <= not (a xor b);
    layer8_outputs(2022) <= not (a and b);
    layer8_outputs(2023) <= b;
    layer8_outputs(2024) <= a and b;
    layer8_outputs(2025) <= a xor b;
    layer8_outputs(2026) <= not a or b;
    layer8_outputs(2027) <= '1';
    layer8_outputs(2028) <= not b;
    layer8_outputs(2029) <= not (a xor b);
    layer8_outputs(2030) <= a and not b;
    layer8_outputs(2031) <= not (a xor b);
    layer8_outputs(2032) <= not b;
    layer8_outputs(2033) <= not b;
    layer8_outputs(2034) <= a and b;
    layer8_outputs(2035) <= not (a and b);
    layer8_outputs(2036) <= a xor b;
    layer8_outputs(2037) <= a xor b;
    layer8_outputs(2038) <= a xor b;
    layer8_outputs(2039) <= not (a xor b);
    layer8_outputs(2040) <= a xor b;
    layer8_outputs(2041) <= not b;
    layer8_outputs(2042) <= b;
    layer8_outputs(2043) <= not a;
    layer8_outputs(2044) <= b and not a;
    layer8_outputs(2045) <= a and not b;
    layer8_outputs(2046) <= not (a or b);
    layer8_outputs(2047) <= a;
    layer8_outputs(2048) <= b and not a;
    layer8_outputs(2049) <= not (a and b);
    layer8_outputs(2050) <= not (a or b);
    layer8_outputs(2051) <= a and not b;
    layer8_outputs(2052) <= a and b;
    layer8_outputs(2053) <= not a;
    layer8_outputs(2054) <= a and not b;
    layer8_outputs(2055) <= not b;
    layer8_outputs(2056) <= a;
    layer8_outputs(2057) <= not (a xor b);
    layer8_outputs(2058) <= not b;
    layer8_outputs(2059) <= b and not a;
    layer8_outputs(2060) <= b and not a;
    layer8_outputs(2061) <= not a;
    layer8_outputs(2062) <= b and not a;
    layer8_outputs(2063) <= not (a xor b);
    layer8_outputs(2064) <= b;
    layer8_outputs(2065) <= a;
    layer8_outputs(2066) <= a;
    layer8_outputs(2067) <= b;
    layer8_outputs(2068) <= not a or b;
    layer8_outputs(2069) <= b and not a;
    layer8_outputs(2070) <= a and b;
    layer8_outputs(2071) <= not (a and b);
    layer8_outputs(2072) <= not (a xor b);
    layer8_outputs(2073) <= '1';
    layer8_outputs(2074) <= a xor b;
    layer8_outputs(2075) <= not b;
    layer8_outputs(2076) <= a xor b;
    layer8_outputs(2077) <= a and not b;
    layer8_outputs(2078) <= a and not b;
    layer8_outputs(2079) <= not a;
    layer8_outputs(2080) <= b;
    layer8_outputs(2081) <= not (a or b);
    layer8_outputs(2082) <= not (a and b);
    layer8_outputs(2083) <= a or b;
    layer8_outputs(2084) <= not a;
    layer8_outputs(2085) <= a and b;
    layer8_outputs(2086) <= not (a xor b);
    layer8_outputs(2087) <= b and not a;
    layer8_outputs(2088) <= not a or b;
    layer8_outputs(2089) <= not (a xor b);
    layer8_outputs(2090) <= not (a xor b);
    layer8_outputs(2091) <= not (a and b);
    layer8_outputs(2092) <= not b;
    layer8_outputs(2093) <= not (a xor b);
    layer8_outputs(2094) <= b;
    layer8_outputs(2095) <= b;
    layer8_outputs(2096) <= not b or a;
    layer8_outputs(2097) <= a or b;
    layer8_outputs(2098) <= not (a or b);
    layer8_outputs(2099) <= b;
    layer8_outputs(2100) <= a xor b;
    layer8_outputs(2101) <= a;
    layer8_outputs(2102) <= a;
    layer8_outputs(2103) <= not a or b;
    layer8_outputs(2104) <= a and b;
    layer8_outputs(2105) <= a;
    layer8_outputs(2106) <= a;
    layer8_outputs(2107) <= not a;
    layer8_outputs(2108) <= not a;
    layer8_outputs(2109) <= not a;
    layer8_outputs(2110) <= not a;
    layer8_outputs(2111) <= a;
    layer8_outputs(2112) <= not b or a;
    layer8_outputs(2113) <= not (a xor b);
    layer8_outputs(2114) <= a and not b;
    layer8_outputs(2115) <= b and not a;
    layer8_outputs(2116) <= b;
    layer8_outputs(2117) <= b;
    layer8_outputs(2118) <= not a;
    layer8_outputs(2119) <= not b;
    layer8_outputs(2120) <= a xor b;
    layer8_outputs(2121) <= not a or b;
    layer8_outputs(2122) <= not a;
    layer8_outputs(2123) <= b and not a;
    layer8_outputs(2124) <= not a;
    layer8_outputs(2125) <= not a or b;
    layer8_outputs(2126) <= a or b;
    layer8_outputs(2127) <= not b or a;
    layer8_outputs(2128) <= not a;
    layer8_outputs(2129) <= not (a and b);
    layer8_outputs(2130) <= not b;
    layer8_outputs(2131) <= a xor b;
    layer8_outputs(2132) <= not a or b;
    layer8_outputs(2133) <= a;
    layer8_outputs(2134) <= a;
    layer8_outputs(2135) <= b;
    layer8_outputs(2136) <= not (a or b);
    layer8_outputs(2137) <= a or b;
    layer8_outputs(2138) <= a;
    layer8_outputs(2139) <= a;
    layer8_outputs(2140) <= not b or a;
    layer8_outputs(2141) <= b;
    layer8_outputs(2142) <= b and not a;
    layer8_outputs(2143) <= a and not b;
    layer8_outputs(2144) <= not a;
    layer8_outputs(2145) <= not (a and b);
    layer8_outputs(2146) <= a and not b;
    layer8_outputs(2147) <= b and not a;
    layer8_outputs(2148) <= b;
    layer8_outputs(2149) <= not b;
    layer8_outputs(2150) <= a xor b;
    layer8_outputs(2151) <= not a;
    layer8_outputs(2152) <= not a;
    layer8_outputs(2153) <= b and not a;
    layer8_outputs(2154) <= not b or a;
    layer8_outputs(2155) <= a or b;
    layer8_outputs(2156) <= not (a xor b);
    layer8_outputs(2157) <= not (a and b);
    layer8_outputs(2158) <= b;
    layer8_outputs(2159) <= a xor b;
    layer8_outputs(2160) <= b and not a;
    layer8_outputs(2161) <= b;
    layer8_outputs(2162) <= a;
    layer8_outputs(2163) <= b;
    layer8_outputs(2164) <= not a or b;
    layer8_outputs(2165) <= a;
    layer8_outputs(2166) <= a xor b;
    layer8_outputs(2167) <= not a or b;
    layer8_outputs(2168) <= not b;
    layer8_outputs(2169) <= not b or a;
    layer8_outputs(2170) <= b;
    layer8_outputs(2171) <= not (a xor b);
    layer8_outputs(2172) <= a;
    layer8_outputs(2173) <= not (a xor b);
    layer8_outputs(2174) <= not b;
    layer8_outputs(2175) <= not b;
    layer8_outputs(2176) <= not b;
    layer8_outputs(2177) <= a and b;
    layer8_outputs(2178) <= not (a and b);
    layer8_outputs(2179) <= not b;
    layer8_outputs(2180) <= not (a xor b);
    layer8_outputs(2181) <= not a;
    layer8_outputs(2182) <= not (a or b);
    layer8_outputs(2183) <= b;
    layer8_outputs(2184) <= not b or a;
    layer8_outputs(2185) <= not a;
    layer8_outputs(2186) <= b and not a;
    layer8_outputs(2187) <= b and not a;
    layer8_outputs(2188) <= a and not b;
    layer8_outputs(2189) <= not b;
    layer8_outputs(2190) <= not (a xor b);
    layer8_outputs(2191) <= not b;
    layer8_outputs(2192) <= not (a or b);
    layer8_outputs(2193) <= not b or a;
    layer8_outputs(2194) <= not (a or b);
    layer8_outputs(2195) <= not (a xor b);
    layer8_outputs(2196) <= b and not a;
    layer8_outputs(2197) <= a or b;
    layer8_outputs(2198) <= not (a and b);
    layer8_outputs(2199) <= not (a xor b);
    layer8_outputs(2200) <= not (a or b);
    layer8_outputs(2201) <= b;
    layer8_outputs(2202) <= b;
    layer8_outputs(2203) <= a;
    layer8_outputs(2204) <= a;
    layer8_outputs(2205) <= not b or a;
    layer8_outputs(2206) <= not a;
    layer8_outputs(2207) <= not b;
    layer8_outputs(2208) <= a;
    layer8_outputs(2209) <= b;
    layer8_outputs(2210) <= b and not a;
    layer8_outputs(2211) <= not b;
    layer8_outputs(2212) <= a xor b;
    layer8_outputs(2213) <= a;
    layer8_outputs(2214) <= not b;
    layer8_outputs(2215) <= not b;
    layer8_outputs(2216) <= b;
    layer8_outputs(2217) <= a and b;
    layer8_outputs(2218) <= not (a xor b);
    layer8_outputs(2219) <= not b;
    layer8_outputs(2220) <= not (a or b);
    layer8_outputs(2221) <= a xor b;
    layer8_outputs(2222) <= not b;
    layer8_outputs(2223) <= not b or a;
    layer8_outputs(2224) <= not b or a;
    layer8_outputs(2225) <= not b;
    layer8_outputs(2226) <= b and not a;
    layer8_outputs(2227) <= a and not b;
    layer8_outputs(2228) <= b;
    layer8_outputs(2229) <= a;
    layer8_outputs(2230) <= a and b;
    layer8_outputs(2231) <= not b;
    layer8_outputs(2232) <= b;
    layer8_outputs(2233) <= a;
    layer8_outputs(2234) <= a xor b;
    layer8_outputs(2235) <= not a;
    layer8_outputs(2236) <= not (a xor b);
    layer8_outputs(2237) <= not b;
    layer8_outputs(2238) <= a and not b;
    layer8_outputs(2239) <= not (a or b);
    layer8_outputs(2240) <= not a;
    layer8_outputs(2241) <= b;
    layer8_outputs(2242) <= not (a xor b);
    layer8_outputs(2243) <= not b or a;
    layer8_outputs(2244) <= a xor b;
    layer8_outputs(2245) <= not b;
    layer8_outputs(2246) <= a;
    layer8_outputs(2247) <= a xor b;
    layer8_outputs(2248) <= not (a xor b);
    layer8_outputs(2249) <= a and b;
    layer8_outputs(2250) <= a xor b;
    layer8_outputs(2251) <= a and b;
    layer8_outputs(2252) <= a;
    layer8_outputs(2253) <= a;
    layer8_outputs(2254) <= not a;
    layer8_outputs(2255) <= not a;
    layer8_outputs(2256) <= not b;
    layer8_outputs(2257) <= b;
    layer8_outputs(2258) <= not a;
    layer8_outputs(2259) <= not a or b;
    layer8_outputs(2260) <= not b;
    layer8_outputs(2261) <= a;
    layer8_outputs(2262) <= not a;
    layer8_outputs(2263) <= not (a or b);
    layer8_outputs(2264) <= a xor b;
    layer8_outputs(2265) <= not (a and b);
    layer8_outputs(2266) <= not (a xor b);
    layer8_outputs(2267) <= not b;
    layer8_outputs(2268) <= b;
    layer8_outputs(2269) <= not a or b;
    layer8_outputs(2270) <= a;
    layer8_outputs(2271) <= b;
    layer8_outputs(2272) <= not (a or b);
    layer8_outputs(2273) <= not b;
    layer8_outputs(2274) <= a xor b;
    layer8_outputs(2275) <= b;
    layer8_outputs(2276) <= a xor b;
    layer8_outputs(2277) <= not a;
    layer8_outputs(2278) <= not (a or b);
    layer8_outputs(2279) <= not (a and b);
    layer8_outputs(2280) <= not a or b;
    layer8_outputs(2281) <= not a or b;
    layer8_outputs(2282) <= not a or b;
    layer8_outputs(2283) <= not b;
    layer8_outputs(2284) <= a and b;
    layer8_outputs(2285) <= not (a and b);
    layer8_outputs(2286) <= a;
    layer8_outputs(2287) <= not a;
    layer8_outputs(2288) <= not (a xor b);
    layer8_outputs(2289) <= not (a xor b);
    layer8_outputs(2290) <= not (a xor b);
    layer8_outputs(2291) <= a or b;
    layer8_outputs(2292) <= not b;
    layer8_outputs(2293) <= not b;
    layer8_outputs(2294) <= b and not a;
    layer8_outputs(2295) <= not a or b;
    layer8_outputs(2296) <= a and not b;
    layer8_outputs(2297) <= '0';
    layer8_outputs(2298) <= a;
    layer8_outputs(2299) <= not a;
    layer8_outputs(2300) <= not (a xor b);
    layer8_outputs(2301) <= not (a or b);
    layer8_outputs(2302) <= not b;
    layer8_outputs(2303) <= not (a and b);
    layer8_outputs(2304) <= not b;
    layer8_outputs(2305) <= a or b;
    layer8_outputs(2306) <= a xor b;
    layer8_outputs(2307) <= not b;
    layer8_outputs(2308) <= a xor b;
    layer8_outputs(2309) <= a xor b;
    layer8_outputs(2310) <= not (a xor b);
    layer8_outputs(2311) <= b;
    layer8_outputs(2312) <= a;
    layer8_outputs(2313) <= b;
    layer8_outputs(2314) <= not b or a;
    layer8_outputs(2315) <= b;
    layer8_outputs(2316) <= b;
    layer8_outputs(2317) <= not b or a;
    layer8_outputs(2318) <= not a;
    layer8_outputs(2319) <= not (a xor b);
    layer8_outputs(2320) <= a xor b;
    layer8_outputs(2321) <= a xor b;
    layer8_outputs(2322) <= not a;
    layer8_outputs(2323) <= not (a xor b);
    layer8_outputs(2324) <= not b;
    layer8_outputs(2325) <= a or b;
    layer8_outputs(2326) <= a;
    layer8_outputs(2327) <= not b;
    layer8_outputs(2328) <= not a;
    layer8_outputs(2329) <= b and not a;
    layer8_outputs(2330) <= b;
    layer8_outputs(2331) <= not (a xor b);
    layer8_outputs(2332) <= not b;
    layer8_outputs(2333) <= b;
    layer8_outputs(2334) <= not a;
    layer8_outputs(2335) <= not (a and b);
    layer8_outputs(2336) <= not (a or b);
    layer8_outputs(2337) <= a and not b;
    layer8_outputs(2338) <= b;
    layer8_outputs(2339) <= a or b;
    layer8_outputs(2340) <= not b or a;
    layer8_outputs(2341) <= not b;
    layer8_outputs(2342) <= not (a and b);
    layer8_outputs(2343) <= not (a or b);
    layer8_outputs(2344) <= a xor b;
    layer8_outputs(2345) <= a xor b;
    layer8_outputs(2346) <= a;
    layer8_outputs(2347) <= not (a or b);
    layer8_outputs(2348) <= b;
    layer8_outputs(2349) <= not b;
    layer8_outputs(2350) <= b;
    layer8_outputs(2351) <= a or b;
    layer8_outputs(2352) <= not a or b;
    layer8_outputs(2353) <= not a;
    layer8_outputs(2354) <= b;
    layer8_outputs(2355) <= a or b;
    layer8_outputs(2356) <= b;
    layer8_outputs(2357) <= b and not a;
    layer8_outputs(2358) <= a xor b;
    layer8_outputs(2359) <= not a;
    layer8_outputs(2360) <= not (a xor b);
    layer8_outputs(2361) <= not (a xor b);
    layer8_outputs(2362) <= not b;
    layer8_outputs(2363) <= a xor b;
    layer8_outputs(2364) <= not b or a;
    layer8_outputs(2365) <= not (a xor b);
    layer8_outputs(2366) <= not a or b;
    layer8_outputs(2367) <= a;
    layer8_outputs(2368) <= b;
    layer8_outputs(2369) <= '0';
    layer8_outputs(2370) <= not (a xor b);
    layer8_outputs(2371) <= b and not a;
    layer8_outputs(2372) <= not a;
    layer8_outputs(2373) <= a xor b;
    layer8_outputs(2374) <= not a;
    layer8_outputs(2375) <= not a or b;
    layer8_outputs(2376) <= not (a xor b);
    layer8_outputs(2377) <= not a;
    layer8_outputs(2378) <= a xor b;
    layer8_outputs(2379) <= not a;
    layer8_outputs(2380) <= a xor b;
    layer8_outputs(2381) <= not b;
    layer8_outputs(2382) <= not a;
    layer8_outputs(2383) <= not b;
    layer8_outputs(2384) <= not b;
    layer8_outputs(2385) <= a xor b;
    layer8_outputs(2386) <= a or b;
    layer8_outputs(2387) <= a and b;
    layer8_outputs(2388) <= a or b;
    layer8_outputs(2389) <= b;
    layer8_outputs(2390) <= a or b;
    layer8_outputs(2391) <= a and b;
    layer8_outputs(2392) <= a;
    layer8_outputs(2393) <= a;
    layer8_outputs(2394) <= a and not b;
    layer8_outputs(2395) <= not b;
    layer8_outputs(2396) <= not a;
    layer8_outputs(2397) <= a xor b;
    layer8_outputs(2398) <= not b;
    layer8_outputs(2399) <= a;
    layer8_outputs(2400) <= b;
    layer8_outputs(2401) <= a and not b;
    layer8_outputs(2402) <= not b;
    layer8_outputs(2403) <= a xor b;
    layer8_outputs(2404) <= a;
    layer8_outputs(2405) <= a xor b;
    layer8_outputs(2406) <= a xor b;
    layer8_outputs(2407) <= not (a or b);
    layer8_outputs(2408) <= a or b;
    layer8_outputs(2409) <= a and not b;
    layer8_outputs(2410) <= not a or b;
    layer8_outputs(2411) <= b;
    layer8_outputs(2412) <= not a or b;
    layer8_outputs(2413) <= a and not b;
    layer8_outputs(2414) <= a and not b;
    layer8_outputs(2415) <= a or b;
    layer8_outputs(2416) <= b;
    layer8_outputs(2417) <= not (a and b);
    layer8_outputs(2418) <= not b;
    layer8_outputs(2419) <= not b;
    layer8_outputs(2420) <= not a;
    layer8_outputs(2421) <= b;
    layer8_outputs(2422) <= not b;
    layer8_outputs(2423) <= not (a xor b);
    layer8_outputs(2424) <= not (a xor b);
    layer8_outputs(2425) <= not b;
    layer8_outputs(2426) <= a xor b;
    layer8_outputs(2427) <= not b;
    layer8_outputs(2428) <= a and b;
    layer8_outputs(2429) <= not b;
    layer8_outputs(2430) <= not (a or b);
    layer8_outputs(2431) <= a or b;
    layer8_outputs(2432) <= not b or a;
    layer8_outputs(2433) <= not a or b;
    layer8_outputs(2434) <= b;
    layer8_outputs(2435) <= not (a and b);
    layer8_outputs(2436) <= a xor b;
    layer8_outputs(2437) <= a;
    layer8_outputs(2438) <= a and b;
    layer8_outputs(2439) <= a or b;
    layer8_outputs(2440) <= a xor b;
    layer8_outputs(2441) <= b;
    layer8_outputs(2442) <= b;
    layer8_outputs(2443) <= not b;
    layer8_outputs(2444) <= not b or a;
    layer8_outputs(2445) <= not b;
    layer8_outputs(2446) <= a xor b;
    layer8_outputs(2447) <= a xor b;
    layer8_outputs(2448) <= not (a xor b);
    layer8_outputs(2449) <= b;
    layer8_outputs(2450) <= a or b;
    layer8_outputs(2451) <= b;
    layer8_outputs(2452) <= not b;
    layer8_outputs(2453) <= not b;
    layer8_outputs(2454) <= a and not b;
    layer8_outputs(2455) <= not b;
    layer8_outputs(2456) <= a xor b;
    layer8_outputs(2457) <= not (a and b);
    layer8_outputs(2458) <= not (a xor b);
    layer8_outputs(2459) <= not (a or b);
    layer8_outputs(2460) <= not a;
    layer8_outputs(2461) <= b and not a;
    layer8_outputs(2462) <= a and not b;
    layer8_outputs(2463) <= not b or a;
    layer8_outputs(2464) <= not b;
    layer8_outputs(2465) <= not b;
    layer8_outputs(2466) <= a or b;
    layer8_outputs(2467) <= a;
    layer8_outputs(2468) <= b;
    layer8_outputs(2469) <= not (a and b);
    layer8_outputs(2470) <= a and not b;
    layer8_outputs(2471) <= b and not a;
    layer8_outputs(2472) <= a xor b;
    layer8_outputs(2473) <= b and not a;
    layer8_outputs(2474) <= a and not b;
    layer8_outputs(2475) <= not a;
    layer8_outputs(2476) <= not (a xor b);
    layer8_outputs(2477) <= b;
    layer8_outputs(2478) <= a and b;
    layer8_outputs(2479) <= a;
    layer8_outputs(2480) <= not (a or b);
    layer8_outputs(2481) <= b;
    layer8_outputs(2482) <= not (a and b);
    layer8_outputs(2483) <= b;
    layer8_outputs(2484) <= b;
    layer8_outputs(2485) <= a;
    layer8_outputs(2486) <= not (a and b);
    layer8_outputs(2487) <= a;
    layer8_outputs(2488) <= a and not b;
    layer8_outputs(2489) <= a xor b;
    layer8_outputs(2490) <= not b;
    layer8_outputs(2491) <= not b;
    layer8_outputs(2492) <= not a or b;
    layer8_outputs(2493) <= a xor b;
    layer8_outputs(2494) <= not a;
    layer8_outputs(2495) <= b and not a;
    layer8_outputs(2496) <= a;
    layer8_outputs(2497) <= not b;
    layer8_outputs(2498) <= a and b;
    layer8_outputs(2499) <= b and not a;
    layer8_outputs(2500) <= not (a or b);
    layer8_outputs(2501) <= a xor b;
    layer8_outputs(2502) <= not (a or b);
    layer8_outputs(2503) <= a;
    layer8_outputs(2504) <= not b;
    layer8_outputs(2505) <= not (a xor b);
    layer8_outputs(2506) <= b and not a;
    layer8_outputs(2507) <= not a or b;
    layer8_outputs(2508) <= not (a and b);
    layer8_outputs(2509) <= not a;
    layer8_outputs(2510) <= a;
    layer8_outputs(2511) <= b;
    layer8_outputs(2512) <= not a;
    layer8_outputs(2513) <= a xor b;
    layer8_outputs(2514) <= b;
    layer8_outputs(2515) <= not (a and b);
    layer8_outputs(2516) <= not (a or b);
    layer8_outputs(2517) <= not b;
    layer8_outputs(2518) <= not b or a;
    layer8_outputs(2519) <= not a;
    layer8_outputs(2520) <= not (a and b);
    layer8_outputs(2521) <= b;
    layer8_outputs(2522) <= '1';
    layer8_outputs(2523) <= not a;
    layer8_outputs(2524) <= b;
    layer8_outputs(2525) <= a or b;
    layer8_outputs(2526) <= '1';
    layer8_outputs(2527) <= not (a xor b);
    layer8_outputs(2528) <= not a or b;
    layer8_outputs(2529) <= not a;
    layer8_outputs(2530) <= not b;
    layer8_outputs(2531) <= b;
    layer8_outputs(2532) <= not a;
    layer8_outputs(2533) <= b;
    layer8_outputs(2534) <= not a;
    layer8_outputs(2535) <= not b;
    layer8_outputs(2536) <= not a;
    layer8_outputs(2537) <= '0';
    layer8_outputs(2538) <= not b or a;
    layer8_outputs(2539) <= b;
    layer8_outputs(2540) <= b;
    layer8_outputs(2541) <= b;
    layer8_outputs(2542) <= not b or a;
    layer8_outputs(2543) <= not b;
    layer8_outputs(2544) <= not b or a;
    layer8_outputs(2545) <= not (a and b);
    layer8_outputs(2546) <= not a;
    layer8_outputs(2547) <= not (a xor b);
    layer8_outputs(2548) <= a;
    layer8_outputs(2549) <= a and b;
    layer8_outputs(2550) <= not b;
    layer8_outputs(2551) <= not b;
    layer8_outputs(2552) <= not a;
    layer8_outputs(2553) <= not (a and b);
    layer8_outputs(2554) <= not b;
    layer8_outputs(2555) <= a;
    layer8_outputs(2556) <= b and not a;
    layer8_outputs(2557) <= b;
    layer8_outputs(2558) <= not (a xor b);
    layer8_outputs(2559) <= a xor b;
    layer8_outputs(2560) <= a and not b;
    layer8_outputs(2561) <= a;
    layer8_outputs(2562) <= not (a and b);
    layer8_outputs(2563) <= b;
    layer8_outputs(2564) <= a and not b;
    layer8_outputs(2565) <= a xor b;
    layer8_outputs(2566) <= a;
    layer8_outputs(2567) <= not a;
    layer8_outputs(2568) <= not (a xor b);
    layer8_outputs(2569) <= a;
    layer8_outputs(2570) <= not a;
    layer8_outputs(2571) <= not b;
    layer8_outputs(2572) <= not b or a;
    layer8_outputs(2573) <= not (a xor b);
    layer8_outputs(2574) <= b;
    layer8_outputs(2575) <= not (a xor b);
    layer8_outputs(2576) <= b and not a;
    layer8_outputs(2577) <= not (a and b);
    layer8_outputs(2578) <= not b or a;
    layer8_outputs(2579) <= a xor b;
    layer8_outputs(2580) <= a or b;
    layer8_outputs(2581) <= a xor b;
    layer8_outputs(2582) <= a xor b;
    layer8_outputs(2583) <= not a;
    layer8_outputs(2584) <= not b;
    layer8_outputs(2585) <= a;
    layer8_outputs(2586) <= b and not a;
    layer8_outputs(2587) <= a xor b;
    layer8_outputs(2588) <= b;
    layer8_outputs(2589) <= b;
    layer8_outputs(2590) <= not (a xor b);
    layer8_outputs(2591) <= not b;
    layer8_outputs(2592) <= a or b;
    layer8_outputs(2593) <= not b or a;
    layer8_outputs(2594) <= not b;
    layer8_outputs(2595) <= a or b;
    layer8_outputs(2596) <= a or b;
    layer8_outputs(2597) <= '1';
    layer8_outputs(2598) <= '1';
    layer8_outputs(2599) <= b and not a;
    layer8_outputs(2600) <= b and not a;
    layer8_outputs(2601) <= b;
    layer8_outputs(2602) <= a;
    layer8_outputs(2603) <= b and not a;
    layer8_outputs(2604) <= a;
    layer8_outputs(2605) <= a or b;
    layer8_outputs(2606) <= a;
    layer8_outputs(2607) <= not (a and b);
    layer8_outputs(2608) <= not a or b;
    layer8_outputs(2609) <= not b;
    layer8_outputs(2610) <= not b;
    layer8_outputs(2611) <= not (a xor b);
    layer8_outputs(2612) <= a or b;
    layer8_outputs(2613) <= b;
    layer8_outputs(2614) <= not b or a;
    layer8_outputs(2615) <= not (a xor b);
    layer8_outputs(2616) <= a;
    layer8_outputs(2617) <= not a;
    layer8_outputs(2618) <= b;
    layer8_outputs(2619) <= a xor b;
    layer8_outputs(2620) <= not (a xor b);
    layer8_outputs(2621) <= not a or b;
    layer8_outputs(2622) <= a;
    layer8_outputs(2623) <= a and b;
    layer8_outputs(2624) <= b;
    layer8_outputs(2625) <= not (a xor b);
    layer8_outputs(2626) <= a;
    layer8_outputs(2627) <= a;
    layer8_outputs(2628) <= not a;
    layer8_outputs(2629) <= a;
    layer8_outputs(2630) <= not b;
    layer8_outputs(2631) <= not (a xor b);
    layer8_outputs(2632) <= a xor b;
    layer8_outputs(2633) <= b and not a;
    layer8_outputs(2634) <= a xor b;
    layer8_outputs(2635) <= not b or a;
    layer8_outputs(2636) <= a and not b;
    layer8_outputs(2637) <= not (a and b);
    layer8_outputs(2638) <= not (a xor b);
    layer8_outputs(2639) <= a xor b;
    layer8_outputs(2640) <= b;
    layer8_outputs(2641) <= a xor b;
    layer8_outputs(2642) <= not (a xor b);
    layer8_outputs(2643) <= a xor b;
    layer8_outputs(2644) <= not (a and b);
    layer8_outputs(2645) <= not (a and b);
    layer8_outputs(2646) <= a or b;
    layer8_outputs(2647) <= b;
    layer8_outputs(2648) <= not b;
    layer8_outputs(2649) <= not b or a;
    layer8_outputs(2650) <= not b;
    layer8_outputs(2651) <= b;
    layer8_outputs(2652) <= not (a xor b);
    layer8_outputs(2653) <= a and b;
    layer8_outputs(2654) <= a;
    layer8_outputs(2655) <= not a;
    layer8_outputs(2656) <= not (a xor b);
    layer8_outputs(2657) <= a and b;
    layer8_outputs(2658) <= b;
    layer8_outputs(2659) <= not b;
    layer8_outputs(2660) <= not b;
    layer8_outputs(2661) <= not b;
    layer8_outputs(2662) <= not a or b;
    layer8_outputs(2663) <= a and b;
    layer8_outputs(2664) <= a;
    layer8_outputs(2665) <= not (a xor b);
    layer8_outputs(2666) <= not b or a;
    layer8_outputs(2667) <= not b or a;
    layer8_outputs(2668) <= not a;
    layer8_outputs(2669) <= not (a or b);
    layer8_outputs(2670) <= not a;
    layer8_outputs(2671) <= not (a and b);
    layer8_outputs(2672) <= not a;
    layer8_outputs(2673) <= not b;
    layer8_outputs(2674) <= a;
    layer8_outputs(2675) <= not a;
    layer8_outputs(2676) <= not (a xor b);
    layer8_outputs(2677) <= b;
    layer8_outputs(2678) <= b and not a;
    layer8_outputs(2679) <= not a or b;
    layer8_outputs(2680) <= not (a xor b);
    layer8_outputs(2681) <= b;
    layer8_outputs(2682) <= not (a xor b);
    layer8_outputs(2683) <= not a;
    layer8_outputs(2684) <= not b or a;
    layer8_outputs(2685) <= not (a and b);
    layer8_outputs(2686) <= b and not a;
    layer8_outputs(2687) <= not (a xor b);
    layer8_outputs(2688) <= a;
    layer8_outputs(2689) <= b;
    layer8_outputs(2690) <= a and b;
    layer8_outputs(2691) <= b;
    layer8_outputs(2692) <= not b;
    layer8_outputs(2693) <= b;
    layer8_outputs(2694) <= b;
    layer8_outputs(2695) <= not b or a;
    layer8_outputs(2696) <= not (a xor b);
    layer8_outputs(2697) <= a and not b;
    layer8_outputs(2698) <= a;
    layer8_outputs(2699) <= not (a or b);
    layer8_outputs(2700) <= a;
    layer8_outputs(2701) <= a xor b;
    layer8_outputs(2702) <= a xor b;
    layer8_outputs(2703) <= not (a and b);
    layer8_outputs(2704) <= a;
    layer8_outputs(2705) <= a and b;
    layer8_outputs(2706) <= not b;
    layer8_outputs(2707) <= b;
    layer8_outputs(2708) <= a xor b;
    layer8_outputs(2709) <= not (a xor b);
    layer8_outputs(2710) <= b and not a;
    layer8_outputs(2711) <= a;
    layer8_outputs(2712) <= '0';
    layer8_outputs(2713) <= not (a xor b);
    layer8_outputs(2714) <= not b or a;
    layer8_outputs(2715) <= a;
    layer8_outputs(2716) <= not b;
    layer8_outputs(2717) <= b;
    layer8_outputs(2718) <= a and not b;
    layer8_outputs(2719) <= b;
    layer8_outputs(2720) <= a;
    layer8_outputs(2721) <= not b;
    layer8_outputs(2722) <= not (a and b);
    layer8_outputs(2723) <= a and b;
    layer8_outputs(2724) <= not (a and b);
    layer8_outputs(2725) <= a xor b;
    layer8_outputs(2726) <= not a or b;
    layer8_outputs(2727) <= not a;
    layer8_outputs(2728) <= not a;
    layer8_outputs(2729) <= a and b;
    layer8_outputs(2730) <= not a or b;
    layer8_outputs(2731) <= a;
    layer8_outputs(2732) <= a xor b;
    layer8_outputs(2733) <= not (a and b);
    layer8_outputs(2734) <= a or b;
    layer8_outputs(2735) <= not (a or b);
    layer8_outputs(2736) <= not (a or b);
    layer8_outputs(2737) <= a xor b;
    layer8_outputs(2738) <= a and not b;
    layer8_outputs(2739) <= not b;
    layer8_outputs(2740) <= a or b;
    layer8_outputs(2741) <= a;
    layer8_outputs(2742) <= a;
    layer8_outputs(2743) <= not b;
    layer8_outputs(2744) <= a;
    layer8_outputs(2745) <= not (a xor b);
    layer8_outputs(2746) <= a;
    layer8_outputs(2747) <= not (a and b);
    layer8_outputs(2748) <= a xor b;
    layer8_outputs(2749) <= a or b;
    layer8_outputs(2750) <= not (a xor b);
    layer8_outputs(2751) <= a or b;
    layer8_outputs(2752) <= b;
    layer8_outputs(2753) <= not b;
    layer8_outputs(2754) <= b;
    layer8_outputs(2755) <= not (a xor b);
    layer8_outputs(2756) <= not b or a;
    layer8_outputs(2757) <= not (a xor b);
    layer8_outputs(2758) <= a xor b;
    layer8_outputs(2759) <= not b;
    layer8_outputs(2760) <= a;
    layer8_outputs(2761) <= b;
    layer8_outputs(2762) <= a xor b;
    layer8_outputs(2763) <= a and not b;
    layer8_outputs(2764) <= b;
    layer8_outputs(2765) <= not (a xor b);
    layer8_outputs(2766) <= a;
    layer8_outputs(2767) <= not b;
    layer8_outputs(2768) <= not b;
    layer8_outputs(2769) <= not (a or b);
    layer8_outputs(2770) <= not (a xor b);
    layer8_outputs(2771) <= b;
    layer8_outputs(2772) <= not (a and b);
    layer8_outputs(2773) <= a xor b;
    layer8_outputs(2774) <= a and not b;
    layer8_outputs(2775) <= not (a and b);
    layer8_outputs(2776) <= not (a xor b);
    layer8_outputs(2777) <= b and not a;
    layer8_outputs(2778) <= b and not a;
    layer8_outputs(2779) <= a and b;
    layer8_outputs(2780) <= a;
    layer8_outputs(2781) <= a;
    layer8_outputs(2782) <= '0';
    layer8_outputs(2783) <= a;
    layer8_outputs(2784) <= b;
    layer8_outputs(2785) <= not a;
    layer8_outputs(2786) <= a xor b;
    layer8_outputs(2787) <= b;
    layer8_outputs(2788) <= not a or b;
    layer8_outputs(2789) <= not a;
    layer8_outputs(2790) <= not b;
    layer8_outputs(2791) <= not (a xor b);
    layer8_outputs(2792) <= a;
    layer8_outputs(2793) <= not (a or b);
    layer8_outputs(2794) <= not (a or b);
    layer8_outputs(2795) <= a and not b;
    layer8_outputs(2796) <= not a;
    layer8_outputs(2797) <= a xor b;
    layer8_outputs(2798) <= not (a or b);
    layer8_outputs(2799) <= not (a xor b);
    layer8_outputs(2800) <= not a;
    layer8_outputs(2801) <= b;
    layer8_outputs(2802) <= a;
    layer8_outputs(2803) <= a or b;
    layer8_outputs(2804) <= not a or b;
    layer8_outputs(2805) <= a or b;
    layer8_outputs(2806) <= not b;
    layer8_outputs(2807) <= not (a xor b);
    layer8_outputs(2808) <= not (a and b);
    layer8_outputs(2809) <= b and not a;
    layer8_outputs(2810) <= not b;
    layer8_outputs(2811) <= b;
    layer8_outputs(2812) <= not (a and b);
    layer8_outputs(2813) <= not (a xor b);
    layer8_outputs(2814) <= a xor b;
    layer8_outputs(2815) <= not b or a;
    layer8_outputs(2816) <= not (a xor b);
    layer8_outputs(2817) <= not (a xor b);
    layer8_outputs(2818) <= a and b;
    layer8_outputs(2819) <= not b;
    layer8_outputs(2820) <= a;
    layer8_outputs(2821) <= a xor b;
    layer8_outputs(2822) <= not (a xor b);
    layer8_outputs(2823) <= a or b;
    layer8_outputs(2824) <= not (a and b);
    layer8_outputs(2825) <= not a;
    layer8_outputs(2826) <= b and not a;
    layer8_outputs(2827) <= a xor b;
    layer8_outputs(2828) <= not a;
    layer8_outputs(2829) <= not (a xor b);
    layer8_outputs(2830) <= not a;
    layer8_outputs(2831) <= not a or b;
    layer8_outputs(2832) <= not b;
    layer8_outputs(2833) <= not b;
    layer8_outputs(2834) <= not (a xor b);
    layer8_outputs(2835) <= not (a and b);
    layer8_outputs(2836) <= not (a and b);
    layer8_outputs(2837) <= b and not a;
    layer8_outputs(2838) <= b and not a;
    layer8_outputs(2839) <= not a;
    layer8_outputs(2840) <= a;
    layer8_outputs(2841) <= a xor b;
    layer8_outputs(2842) <= b;
    layer8_outputs(2843) <= not a;
    layer8_outputs(2844) <= not b or a;
    layer8_outputs(2845) <= not (a or b);
    layer8_outputs(2846) <= not (a and b);
    layer8_outputs(2847) <= not (a xor b);
    layer8_outputs(2848) <= not b;
    layer8_outputs(2849) <= a;
    layer8_outputs(2850) <= b;
    layer8_outputs(2851) <= not b;
    layer8_outputs(2852) <= a;
    layer8_outputs(2853) <= not (a and b);
    layer8_outputs(2854) <= a;
    layer8_outputs(2855) <= a xor b;
    layer8_outputs(2856) <= b;
    layer8_outputs(2857) <= not (a or b);
    layer8_outputs(2858) <= a;
    layer8_outputs(2859) <= not (a and b);
    layer8_outputs(2860) <= not a;
    layer8_outputs(2861) <= not (a and b);
    layer8_outputs(2862) <= a and not b;
    layer8_outputs(2863) <= not a;
    layer8_outputs(2864) <= not a or b;
    layer8_outputs(2865) <= b and not a;
    layer8_outputs(2866) <= b;
    layer8_outputs(2867) <= a xor b;
    layer8_outputs(2868) <= a xor b;
    layer8_outputs(2869) <= a xor b;
    layer8_outputs(2870) <= not b;
    layer8_outputs(2871) <= a xor b;
    layer8_outputs(2872) <= not (a xor b);
    layer8_outputs(2873) <= b and not a;
    layer8_outputs(2874) <= not a;
    layer8_outputs(2875) <= a;
    layer8_outputs(2876) <= b and not a;
    layer8_outputs(2877) <= not a;
    layer8_outputs(2878) <= a xor b;
    layer8_outputs(2879) <= b and not a;
    layer8_outputs(2880) <= a or b;
    layer8_outputs(2881) <= b and not a;
    layer8_outputs(2882) <= b;
    layer8_outputs(2883) <= not b;
    layer8_outputs(2884) <= not (a xor b);
    layer8_outputs(2885) <= not b;
    layer8_outputs(2886) <= a;
    layer8_outputs(2887) <= not b or a;
    layer8_outputs(2888) <= a and b;
    layer8_outputs(2889) <= a;
    layer8_outputs(2890) <= not a;
    layer8_outputs(2891) <= not (a xor b);
    layer8_outputs(2892) <= not (a xor b);
    layer8_outputs(2893) <= not (a xor b);
    layer8_outputs(2894) <= b;
    layer8_outputs(2895) <= not b;
    layer8_outputs(2896) <= a;
    layer8_outputs(2897) <= '0';
    layer8_outputs(2898) <= a;
    layer8_outputs(2899) <= not a;
    layer8_outputs(2900) <= not b;
    layer8_outputs(2901) <= not (a xor b);
    layer8_outputs(2902) <= not a;
    layer8_outputs(2903) <= not (a xor b);
    layer8_outputs(2904) <= not b or a;
    layer8_outputs(2905) <= a xor b;
    layer8_outputs(2906) <= not (a or b);
    layer8_outputs(2907) <= '0';
    layer8_outputs(2908) <= a xor b;
    layer8_outputs(2909) <= a;
    layer8_outputs(2910) <= not (a xor b);
    layer8_outputs(2911) <= not a;
    layer8_outputs(2912) <= not a;
    layer8_outputs(2913) <= a;
    layer8_outputs(2914) <= not a;
    layer8_outputs(2915) <= b;
    layer8_outputs(2916) <= not a;
    layer8_outputs(2917) <= a;
    layer8_outputs(2918) <= not b or a;
    layer8_outputs(2919) <= b;
    layer8_outputs(2920) <= b;
    layer8_outputs(2921) <= not a;
    layer8_outputs(2922) <= a xor b;
    layer8_outputs(2923) <= b;
    layer8_outputs(2924) <= not b;
    layer8_outputs(2925) <= a;
    layer8_outputs(2926) <= a xor b;
    layer8_outputs(2927) <= b;
    layer8_outputs(2928) <= a xor b;
    layer8_outputs(2929) <= a xor b;
    layer8_outputs(2930) <= a;
    layer8_outputs(2931) <= not (a and b);
    layer8_outputs(2932) <= not (a or b);
    layer8_outputs(2933) <= a;
    layer8_outputs(2934) <= not (a xor b);
    layer8_outputs(2935) <= b;
    layer8_outputs(2936) <= b;
    layer8_outputs(2937) <= not b or a;
    layer8_outputs(2938) <= a xor b;
    layer8_outputs(2939) <= not a;
    layer8_outputs(2940) <= a and b;
    layer8_outputs(2941) <= a and not b;
    layer8_outputs(2942) <= b and not a;
    layer8_outputs(2943) <= b and not a;
    layer8_outputs(2944) <= b;
    layer8_outputs(2945) <= a and not b;
    layer8_outputs(2946) <= b;
    layer8_outputs(2947) <= a xor b;
    layer8_outputs(2948) <= a xor b;
    layer8_outputs(2949) <= a and b;
    layer8_outputs(2950) <= a;
    layer8_outputs(2951) <= b and not a;
    layer8_outputs(2952) <= not (a xor b);
    layer8_outputs(2953) <= a;
    layer8_outputs(2954) <= not b;
    layer8_outputs(2955) <= not (a and b);
    layer8_outputs(2956) <= not b or a;
    layer8_outputs(2957) <= a and b;
    layer8_outputs(2958) <= a;
    layer8_outputs(2959) <= not b or a;
    layer8_outputs(2960) <= b;
    layer8_outputs(2961) <= a or b;
    layer8_outputs(2962) <= not a;
    layer8_outputs(2963) <= a or b;
    layer8_outputs(2964) <= a;
    layer8_outputs(2965) <= not b;
    layer8_outputs(2966) <= not a;
    layer8_outputs(2967) <= not b or a;
    layer8_outputs(2968) <= a xor b;
    layer8_outputs(2969) <= a;
    layer8_outputs(2970) <= a;
    layer8_outputs(2971) <= b;
    layer8_outputs(2972) <= not b;
    layer8_outputs(2973) <= not b;
    layer8_outputs(2974) <= not (a and b);
    layer8_outputs(2975) <= not b or a;
    layer8_outputs(2976) <= a;
    layer8_outputs(2977) <= a or b;
    layer8_outputs(2978) <= b;
    layer8_outputs(2979) <= not a or b;
    layer8_outputs(2980) <= a and b;
    layer8_outputs(2981) <= not a;
    layer8_outputs(2982) <= a;
    layer8_outputs(2983) <= not a or b;
    layer8_outputs(2984) <= not a;
    layer8_outputs(2985) <= a xor b;
    layer8_outputs(2986) <= not a;
    layer8_outputs(2987) <= b;
    layer8_outputs(2988) <= not a;
    layer8_outputs(2989) <= not a;
    layer8_outputs(2990) <= not a;
    layer8_outputs(2991) <= b;
    layer8_outputs(2992) <= b and not a;
    layer8_outputs(2993) <= a and not b;
    layer8_outputs(2994) <= not b;
    layer8_outputs(2995) <= a xor b;
    layer8_outputs(2996) <= not b;
    layer8_outputs(2997) <= not (a xor b);
    layer8_outputs(2998) <= not b or a;
    layer8_outputs(2999) <= not a or b;
    layer8_outputs(3000) <= not (a or b);
    layer8_outputs(3001) <= b;
    layer8_outputs(3002) <= not (a or b);
    layer8_outputs(3003) <= not b;
    layer8_outputs(3004) <= a xor b;
    layer8_outputs(3005) <= b;
    layer8_outputs(3006) <= b;
    layer8_outputs(3007) <= a xor b;
    layer8_outputs(3008) <= a;
    layer8_outputs(3009) <= not (a and b);
    layer8_outputs(3010) <= not (a or b);
    layer8_outputs(3011) <= not b;
    layer8_outputs(3012) <= b;
    layer8_outputs(3013) <= b;
    layer8_outputs(3014) <= not (a xor b);
    layer8_outputs(3015) <= b;
    layer8_outputs(3016) <= b;
    layer8_outputs(3017) <= not (a xor b);
    layer8_outputs(3018) <= a;
    layer8_outputs(3019) <= not a or b;
    layer8_outputs(3020) <= '1';
    layer8_outputs(3021) <= not b;
    layer8_outputs(3022) <= not b;
    layer8_outputs(3023) <= not a;
    layer8_outputs(3024) <= not (a or b);
    layer8_outputs(3025) <= a xor b;
    layer8_outputs(3026) <= b;
    layer8_outputs(3027) <= not b or a;
    layer8_outputs(3028) <= not b;
    layer8_outputs(3029) <= not (a and b);
    layer8_outputs(3030) <= b;
    layer8_outputs(3031) <= not b;
    layer8_outputs(3032) <= a;
    layer8_outputs(3033) <= not b;
    layer8_outputs(3034) <= not b;
    layer8_outputs(3035) <= not b or a;
    layer8_outputs(3036) <= not (a and b);
    layer8_outputs(3037) <= not b or a;
    layer8_outputs(3038) <= not (a xor b);
    layer8_outputs(3039) <= a and b;
    layer8_outputs(3040) <= a and b;
    layer8_outputs(3041) <= not (a xor b);
    layer8_outputs(3042) <= not (a xor b);
    layer8_outputs(3043) <= a;
    layer8_outputs(3044) <= b;
    layer8_outputs(3045) <= b;
    layer8_outputs(3046) <= a;
    layer8_outputs(3047) <= not b;
    layer8_outputs(3048) <= a xor b;
    layer8_outputs(3049) <= b;
    layer8_outputs(3050) <= not (a xor b);
    layer8_outputs(3051) <= not b;
    layer8_outputs(3052) <= not a;
    layer8_outputs(3053) <= a or b;
    layer8_outputs(3054) <= a;
    layer8_outputs(3055) <= a xor b;
    layer8_outputs(3056) <= not (a and b);
    layer8_outputs(3057) <= not (a or b);
    layer8_outputs(3058) <= not a;
    layer8_outputs(3059) <= a or b;
    layer8_outputs(3060) <= a xor b;
    layer8_outputs(3061) <= not (a xor b);
    layer8_outputs(3062) <= a or b;
    layer8_outputs(3063) <= a xor b;
    layer8_outputs(3064) <= a;
    layer8_outputs(3065) <= not a;
    layer8_outputs(3066) <= not b;
    layer8_outputs(3067) <= a xor b;
    layer8_outputs(3068) <= a;
    layer8_outputs(3069) <= a;
    layer8_outputs(3070) <= a xor b;
    layer8_outputs(3071) <= a xor b;
    layer8_outputs(3072) <= not b;
    layer8_outputs(3073) <= not (a xor b);
    layer8_outputs(3074) <= not b;
    layer8_outputs(3075) <= not b or a;
    layer8_outputs(3076) <= not b;
    layer8_outputs(3077) <= a and not b;
    layer8_outputs(3078) <= b;
    layer8_outputs(3079) <= a or b;
    layer8_outputs(3080) <= not a;
    layer8_outputs(3081) <= not b;
    layer8_outputs(3082) <= a;
    layer8_outputs(3083) <= not (a and b);
    layer8_outputs(3084) <= a;
    layer8_outputs(3085) <= not (a and b);
    layer8_outputs(3086) <= not b or a;
    layer8_outputs(3087) <= not b;
    layer8_outputs(3088) <= b;
    layer8_outputs(3089) <= b;
    layer8_outputs(3090) <= not (a or b);
    layer8_outputs(3091) <= not (a and b);
    layer8_outputs(3092) <= not b;
    layer8_outputs(3093) <= a xor b;
    layer8_outputs(3094) <= a and not b;
    layer8_outputs(3095) <= b and not a;
    layer8_outputs(3096) <= not a;
    layer8_outputs(3097) <= b;
    layer8_outputs(3098) <= not (a and b);
    layer8_outputs(3099) <= a and b;
    layer8_outputs(3100) <= not b;
    layer8_outputs(3101) <= b;
    layer8_outputs(3102) <= a xor b;
    layer8_outputs(3103) <= a xor b;
    layer8_outputs(3104) <= a xor b;
    layer8_outputs(3105) <= a xor b;
    layer8_outputs(3106) <= not (a or b);
    layer8_outputs(3107) <= a or b;
    layer8_outputs(3108) <= a;
    layer8_outputs(3109) <= not (a xor b);
    layer8_outputs(3110) <= a xor b;
    layer8_outputs(3111) <= a xor b;
    layer8_outputs(3112) <= not a;
    layer8_outputs(3113) <= a;
    layer8_outputs(3114) <= not b;
    layer8_outputs(3115) <= b;
    layer8_outputs(3116) <= a;
    layer8_outputs(3117) <= not a or b;
    layer8_outputs(3118) <= a or b;
    layer8_outputs(3119) <= not b;
    layer8_outputs(3120) <= not (a and b);
    layer8_outputs(3121) <= not b;
    layer8_outputs(3122) <= a and b;
    layer8_outputs(3123) <= not (a or b);
    layer8_outputs(3124) <= not (a xor b);
    layer8_outputs(3125) <= b and not a;
    layer8_outputs(3126) <= not a;
    layer8_outputs(3127) <= a and b;
    layer8_outputs(3128) <= b;
    layer8_outputs(3129) <= not a;
    layer8_outputs(3130) <= not a;
    layer8_outputs(3131) <= a and b;
    layer8_outputs(3132) <= b;
    layer8_outputs(3133) <= a;
    layer8_outputs(3134) <= not (a xor b);
    layer8_outputs(3135) <= not b or a;
    layer8_outputs(3136) <= not b;
    layer8_outputs(3137) <= a;
    layer8_outputs(3138) <= not b;
    layer8_outputs(3139) <= b;
    layer8_outputs(3140) <= not a;
    layer8_outputs(3141) <= not (a and b);
    layer8_outputs(3142) <= a or b;
    layer8_outputs(3143) <= not b;
    layer8_outputs(3144) <= not a or b;
    layer8_outputs(3145) <= a xor b;
    layer8_outputs(3146) <= not a;
    layer8_outputs(3147) <= a xor b;
    layer8_outputs(3148) <= b;
    layer8_outputs(3149) <= not a or b;
    layer8_outputs(3150) <= not b;
    layer8_outputs(3151) <= not a or b;
    layer8_outputs(3152) <= not (a and b);
    layer8_outputs(3153) <= not b;
    layer8_outputs(3154) <= not (a xor b);
    layer8_outputs(3155) <= b;
    layer8_outputs(3156) <= a and b;
    layer8_outputs(3157) <= not b;
    layer8_outputs(3158) <= a;
    layer8_outputs(3159) <= a and not b;
    layer8_outputs(3160) <= a and b;
    layer8_outputs(3161) <= b;
    layer8_outputs(3162) <= a xor b;
    layer8_outputs(3163) <= a;
    layer8_outputs(3164) <= b;
    layer8_outputs(3165) <= a and b;
    layer8_outputs(3166) <= not a or b;
    layer8_outputs(3167) <= not b;
    layer8_outputs(3168) <= b;
    layer8_outputs(3169) <= b;
    layer8_outputs(3170) <= a;
    layer8_outputs(3171) <= a;
    layer8_outputs(3172) <= not (a xor b);
    layer8_outputs(3173) <= a;
    layer8_outputs(3174) <= b;
    layer8_outputs(3175) <= not b;
    layer8_outputs(3176) <= not a;
    layer8_outputs(3177) <= b;
    layer8_outputs(3178) <= not a or b;
    layer8_outputs(3179) <= not b;
    layer8_outputs(3180) <= a or b;
    layer8_outputs(3181) <= a or b;
    layer8_outputs(3182) <= not a;
    layer8_outputs(3183) <= a xor b;
    layer8_outputs(3184) <= a and b;
    layer8_outputs(3185) <= not b;
    layer8_outputs(3186) <= a xor b;
    layer8_outputs(3187) <= not b;
    layer8_outputs(3188) <= a xor b;
    layer8_outputs(3189) <= not b or a;
    layer8_outputs(3190) <= not b;
    layer8_outputs(3191) <= a;
    layer8_outputs(3192) <= not b;
    layer8_outputs(3193) <= a;
    layer8_outputs(3194) <= a and not b;
    layer8_outputs(3195) <= not a;
    layer8_outputs(3196) <= not a or b;
    layer8_outputs(3197) <= not b;
    layer8_outputs(3198) <= not (a and b);
    layer8_outputs(3199) <= a;
    layer8_outputs(3200) <= a xor b;
    layer8_outputs(3201) <= not b;
    layer8_outputs(3202) <= not a;
    layer8_outputs(3203) <= not a or b;
    layer8_outputs(3204) <= b;
    layer8_outputs(3205) <= not (a and b);
    layer8_outputs(3206) <= a;
    layer8_outputs(3207) <= not (a xor b);
    layer8_outputs(3208) <= a;
    layer8_outputs(3209) <= a;
    layer8_outputs(3210) <= not (a xor b);
    layer8_outputs(3211) <= not a;
    layer8_outputs(3212) <= not b;
    layer8_outputs(3213) <= not b;
    layer8_outputs(3214) <= not (a or b);
    layer8_outputs(3215) <= a and not b;
    layer8_outputs(3216) <= not a;
    layer8_outputs(3217) <= not b;
    layer8_outputs(3218) <= a;
    layer8_outputs(3219) <= b and not a;
    layer8_outputs(3220) <= not b or a;
    layer8_outputs(3221) <= a xor b;
    layer8_outputs(3222) <= not b or a;
    layer8_outputs(3223) <= a and b;
    layer8_outputs(3224) <= not a;
    layer8_outputs(3225) <= a or b;
    layer8_outputs(3226) <= a or b;
    layer8_outputs(3227) <= a xor b;
    layer8_outputs(3228) <= not b;
    layer8_outputs(3229) <= not a;
    layer8_outputs(3230) <= not (a xor b);
    layer8_outputs(3231) <= a;
    layer8_outputs(3232) <= not b;
    layer8_outputs(3233) <= not (a xor b);
    layer8_outputs(3234) <= not b or a;
    layer8_outputs(3235) <= b;
    layer8_outputs(3236) <= not (a and b);
    layer8_outputs(3237) <= a;
    layer8_outputs(3238) <= not b;
    layer8_outputs(3239) <= b and not a;
    layer8_outputs(3240) <= not b;
    layer8_outputs(3241) <= not a or b;
    layer8_outputs(3242) <= not b;
    layer8_outputs(3243) <= not a or b;
    layer8_outputs(3244) <= not (a xor b);
    layer8_outputs(3245) <= b;
    layer8_outputs(3246) <= not (a and b);
    layer8_outputs(3247) <= b;
    layer8_outputs(3248) <= a xor b;
    layer8_outputs(3249) <= a and not b;
    layer8_outputs(3250) <= not b or a;
    layer8_outputs(3251) <= not (a or b);
    layer8_outputs(3252) <= a and b;
    layer8_outputs(3253) <= not (a and b);
    layer8_outputs(3254) <= not (a or b);
    layer8_outputs(3255) <= not b or a;
    layer8_outputs(3256) <= b and not a;
    layer8_outputs(3257) <= a and not b;
    layer8_outputs(3258) <= a xor b;
    layer8_outputs(3259) <= a;
    layer8_outputs(3260) <= not a;
    layer8_outputs(3261) <= not b or a;
    layer8_outputs(3262) <= not a;
    layer8_outputs(3263) <= a;
    layer8_outputs(3264) <= b;
    layer8_outputs(3265) <= not (a xor b);
    layer8_outputs(3266) <= not a;
    layer8_outputs(3267) <= b;
    layer8_outputs(3268) <= not (a xor b);
    layer8_outputs(3269) <= not b or a;
    layer8_outputs(3270) <= a xor b;
    layer8_outputs(3271) <= a;
    layer8_outputs(3272) <= not b or a;
    layer8_outputs(3273) <= b and not a;
    layer8_outputs(3274) <= not b;
    layer8_outputs(3275) <= not a;
    layer8_outputs(3276) <= a xor b;
    layer8_outputs(3277) <= not b or a;
    layer8_outputs(3278) <= a;
    layer8_outputs(3279) <= not a;
    layer8_outputs(3280) <= b and not a;
    layer8_outputs(3281) <= not b;
    layer8_outputs(3282) <= a and b;
    layer8_outputs(3283) <= not (a xor b);
    layer8_outputs(3284) <= not a;
    layer8_outputs(3285) <= not b;
    layer8_outputs(3286) <= not (a xor b);
    layer8_outputs(3287) <= a xor b;
    layer8_outputs(3288) <= a;
    layer8_outputs(3289) <= not a;
    layer8_outputs(3290) <= not b or a;
    layer8_outputs(3291) <= a;
    layer8_outputs(3292) <= not a;
    layer8_outputs(3293) <= a;
    layer8_outputs(3294) <= a;
    layer8_outputs(3295) <= a or b;
    layer8_outputs(3296) <= a;
    layer8_outputs(3297) <= not b;
    layer8_outputs(3298) <= a or b;
    layer8_outputs(3299) <= a and not b;
    layer8_outputs(3300) <= a;
    layer8_outputs(3301) <= not (a and b);
    layer8_outputs(3302) <= a;
    layer8_outputs(3303) <= not (a xor b);
    layer8_outputs(3304) <= b;
    layer8_outputs(3305) <= b;
    layer8_outputs(3306) <= a or b;
    layer8_outputs(3307) <= not (a and b);
    layer8_outputs(3308) <= b;
    layer8_outputs(3309) <= a and not b;
    layer8_outputs(3310) <= a and b;
    layer8_outputs(3311) <= a;
    layer8_outputs(3312) <= a xor b;
    layer8_outputs(3313) <= not (a xor b);
    layer8_outputs(3314) <= not a;
    layer8_outputs(3315) <= not b;
    layer8_outputs(3316) <= not a;
    layer8_outputs(3317) <= not (a xor b);
    layer8_outputs(3318) <= a and b;
    layer8_outputs(3319) <= not (a xor b);
    layer8_outputs(3320) <= b;
    layer8_outputs(3321) <= a xor b;
    layer8_outputs(3322) <= b;
    layer8_outputs(3323) <= '0';
    layer8_outputs(3324) <= b and not a;
    layer8_outputs(3325) <= not (a xor b);
    layer8_outputs(3326) <= not (a xor b);
    layer8_outputs(3327) <= a;
    layer8_outputs(3328) <= a and b;
    layer8_outputs(3329) <= not a;
    layer8_outputs(3330) <= not a;
    layer8_outputs(3331) <= not b;
    layer8_outputs(3332) <= b and not a;
    layer8_outputs(3333) <= not b;
    layer8_outputs(3334) <= b;
    layer8_outputs(3335) <= not (a and b);
    layer8_outputs(3336) <= not b;
    layer8_outputs(3337) <= a or b;
    layer8_outputs(3338) <= a and not b;
    layer8_outputs(3339) <= not b or a;
    layer8_outputs(3340) <= not a;
    layer8_outputs(3341) <= not a;
    layer8_outputs(3342) <= b and not a;
    layer8_outputs(3343) <= b;
    layer8_outputs(3344) <= not a;
    layer8_outputs(3345) <= a and b;
    layer8_outputs(3346) <= a xor b;
    layer8_outputs(3347) <= not (a or b);
    layer8_outputs(3348) <= not b;
    layer8_outputs(3349) <= a;
    layer8_outputs(3350) <= not a or b;
    layer8_outputs(3351) <= not a or b;
    layer8_outputs(3352) <= not a;
    layer8_outputs(3353) <= not a;
    layer8_outputs(3354) <= a or b;
    layer8_outputs(3355) <= a and b;
    layer8_outputs(3356) <= b;
    layer8_outputs(3357) <= not b or a;
    layer8_outputs(3358) <= not a;
    layer8_outputs(3359) <= not a;
    layer8_outputs(3360) <= a;
    layer8_outputs(3361) <= not (a or b);
    layer8_outputs(3362) <= b;
    layer8_outputs(3363) <= not (a xor b);
    layer8_outputs(3364) <= not b or a;
    layer8_outputs(3365) <= a xor b;
    layer8_outputs(3366) <= a xor b;
    layer8_outputs(3367) <= not b;
    layer8_outputs(3368) <= a or b;
    layer8_outputs(3369) <= not a or b;
    layer8_outputs(3370) <= a;
    layer8_outputs(3371) <= not b or a;
    layer8_outputs(3372) <= not a;
    layer8_outputs(3373) <= b;
    layer8_outputs(3374) <= not (a and b);
    layer8_outputs(3375) <= not a;
    layer8_outputs(3376) <= not (a and b);
    layer8_outputs(3377) <= b;
    layer8_outputs(3378) <= a xor b;
    layer8_outputs(3379) <= not a;
    layer8_outputs(3380) <= a;
    layer8_outputs(3381) <= not (a xor b);
    layer8_outputs(3382) <= not b;
    layer8_outputs(3383) <= not (a xor b);
    layer8_outputs(3384) <= b and not a;
    layer8_outputs(3385) <= not (a and b);
    layer8_outputs(3386) <= not a;
    layer8_outputs(3387) <= not b;
    layer8_outputs(3388) <= not a;
    layer8_outputs(3389) <= not (a xor b);
    layer8_outputs(3390) <= not a;
    layer8_outputs(3391) <= a;
    layer8_outputs(3392) <= b;
    layer8_outputs(3393) <= not a;
    layer8_outputs(3394) <= a xor b;
    layer8_outputs(3395) <= not (a or b);
    layer8_outputs(3396) <= not b;
    layer8_outputs(3397) <= a xor b;
    layer8_outputs(3398) <= not (a xor b);
    layer8_outputs(3399) <= not (a or b);
    layer8_outputs(3400) <= not b;
    layer8_outputs(3401) <= b;
    layer8_outputs(3402) <= not b;
    layer8_outputs(3403) <= a xor b;
    layer8_outputs(3404) <= a and b;
    layer8_outputs(3405) <= not a;
    layer8_outputs(3406) <= not b or a;
    layer8_outputs(3407) <= not b or a;
    layer8_outputs(3408) <= not b;
    layer8_outputs(3409) <= not (a xor b);
    layer8_outputs(3410) <= not a or b;
    layer8_outputs(3411) <= a;
    layer8_outputs(3412) <= b;
    layer8_outputs(3413) <= not (a xor b);
    layer8_outputs(3414) <= not a;
    layer8_outputs(3415) <= not b or a;
    layer8_outputs(3416) <= a xor b;
    layer8_outputs(3417) <= b;
    layer8_outputs(3418) <= b and not a;
    layer8_outputs(3419) <= '0';
    layer8_outputs(3420) <= not a;
    layer8_outputs(3421) <= b;
    layer8_outputs(3422) <= not a or b;
    layer8_outputs(3423) <= not b;
    layer8_outputs(3424) <= a;
    layer8_outputs(3425) <= a and b;
    layer8_outputs(3426) <= not a;
    layer8_outputs(3427) <= not (a and b);
    layer8_outputs(3428) <= not b;
    layer8_outputs(3429) <= not b;
    layer8_outputs(3430) <= not b;
    layer8_outputs(3431) <= b;
    layer8_outputs(3432) <= a or b;
    layer8_outputs(3433) <= a and b;
    layer8_outputs(3434) <= not b or a;
    layer8_outputs(3435) <= not a;
    layer8_outputs(3436) <= a;
    layer8_outputs(3437) <= not b;
    layer8_outputs(3438) <= not (a or b);
    layer8_outputs(3439) <= b;
    layer8_outputs(3440) <= not (a xor b);
    layer8_outputs(3441) <= not b;
    layer8_outputs(3442) <= not b;
    layer8_outputs(3443) <= b and not a;
    layer8_outputs(3444) <= b;
    layer8_outputs(3445) <= a xor b;
    layer8_outputs(3446) <= a xor b;
    layer8_outputs(3447) <= b and not a;
    layer8_outputs(3448) <= not b or a;
    layer8_outputs(3449) <= not b;
    layer8_outputs(3450) <= b and not a;
    layer8_outputs(3451) <= not b;
    layer8_outputs(3452) <= a;
    layer8_outputs(3453) <= a xor b;
    layer8_outputs(3454) <= b and not a;
    layer8_outputs(3455) <= not b;
    layer8_outputs(3456) <= not (a xor b);
    layer8_outputs(3457) <= a;
    layer8_outputs(3458) <= not (a or b);
    layer8_outputs(3459) <= a xor b;
    layer8_outputs(3460) <= not (a or b);
    layer8_outputs(3461) <= not (a or b);
    layer8_outputs(3462) <= not a;
    layer8_outputs(3463) <= a;
    layer8_outputs(3464) <= not a;
    layer8_outputs(3465) <= a;
    layer8_outputs(3466) <= not b or a;
    layer8_outputs(3467) <= b;
    layer8_outputs(3468) <= not a;
    layer8_outputs(3469) <= not (a xor b);
    layer8_outputs(3470) <= a and b;
    layer8_outputs(3471) <= a;
    layer8_outputs(3472) <= not (a or b);
    layer8_outputs(3473) <= b;
    layer8_outputs(3474) <= b;
    layer8_outputs(3475) <= not a;
    layer8_outputs(3476) <= not a;
    layer8_outputs(3477) <= a or b;
    layer8_outputs(3478) <= a;
    layer8_outputs(3479) <= a;
    layer8_outputs(3480) <= a and not b;
    layer8_outputs(3481) <= not (a and b);
    layer8_outputs(3482) <= a;
    layer8_outputs(3483) <= not b;
    layer8_outputs(3484) <= a and b;
    layer8_outputs(3485) <= a;
    layer8_outputs(3486) <= a xor b;
    layer8_outputs(3487) <= not b or a;
    layer8_outputs(3488) <= not b or a;
    layer8_outputs(3489) <= not a or b;
    layer8_outputs(3490) <= not b;
    layer8_outputs(3491) <= a and not b;
    layer8_outputs(3492) <= a and not b;
    layer8_outputs(3493) <= not (a and b);
    layer8_outputs(3494) <= not b;
    layer8_outputs(3495) <= not b or a;
    layer8_outputs(3496) <= a;
    layer8_outputs(3497) <= a and b;
    layer8_outputs(3498) <= b;
    layer8_outputs(3499) <= a or b;
    layer8_outputs(3500) <= a and not b;
    layer8_outputs(3501) <= a or b;
    layer8_outputs(3502) <= not b or a;
    layer8_outputs(3503) <= not b or a;
    layer8_outputs(3504) <= b;
    layer8_outputs(3505) <= a;
    layer8_outputs(3506) <= a;
    layer8_outputs(3507) <= a xor b;
    layer8_outputs(3508) <= b;
    layer8_outputs(3509) <= a xor b;
    layer8_outputs(3510) <= a or b;
    layer8_outputs(3511) <= a xor b;
    layer8_outputs(3512) <= not a;
    layer8_outputs(3513) <= a;
    layer8_outputs(3514) <= a;
    layer8_outputs(3515) <= a;
    layer8_outputs(3516) <= b;
    layer8_outputs(3517) <= not b or a;
    layer8_outputs(3518) <= not (a and b);
    layer8_outputs(3519) <= not b;
    layer8_outputs(3520) <= b;
    layer8_outputs(3521) <= b;
    layer8_outputs(3522) <= a xor b;
    layer8_outputs(3523) <= not (a and b);
    layer8_outputs(3524) <= '1';
    layer8_outputs(3525) <= not (a and b);
    layer8_outputs(3526) <= not (a and b);
    layer8_outputs(3527) <= b;
    layer8_outputs(3528) <= not (a xor b);
    layer8_outputs(3529) <= not (a or b);
    layer8_outputs(3530) <= not a or b;
    layer8_outputs(3531) <= not a;
    layer8_outputs(3532) <= not a;
    layer8_outputs(3533) <= not a or b;
    layer8_outputs(3534) <= b;
    layer8_outputs(3535) <= a or b;
    layer8_outputs(3536) <= b and not a;
    layer8_outputs(3537) <= b;
    layer8_outputs(3538) <= a;
    layer8_outputs(3539) <= not a;
    layer8_outputs(3540) <= a xor b;
    layer8_outputs(3541) <= a xor b;
    layer8_outputs(3542) <= not b;
    layer8_outputs(3543) <= not (a xor b);
    layer8_outputs(3544) <= b and not a;
    layer8_outputs(3545) <= a;
    layer8_outputs(3546) <= not (a xor b);
    layer8_outputs(3547) <= not (a xor b);
    layer8_outputs(3548) <= a and b;
    layer8_outputs(3549) <= not (a and b);
    layer8_outputs(3550) <= not (a or b);
    layer8_outputs(3551) <= not (a and b);
    layer8_outputs(3552) <= not (a xor b);
    layer8_outputs(3553) <= not b;
    layer8_outputs(3554) <= not (a xor b);
    layer8_outputs(3555) <= not (a xor b);
    layer8_outputs(3556) <= a and not b;
    layer8_outputs(3557) <= b;
    layer8_outputs(3558) <= not b;
    layer8_outputs(3559) <= not a or b;
    layer8_outputs(3560) <= a;
    layer8_outputs(3561) <= a or b;
    layer8_outputs(3562) <= a and b;
    layer8_outputs(3563) <= not b or a;
    layer8_outputs(3564) <= not b or a;
    layer8_outputs(3565) <= not b;
    layer8_outputs(3566) <= not b;
    layer8_outputs(3567) <= b;
    layer8_outputs(3568) <= a and b;
    layer8_outputs(3569) <= a or b;
    layer8_outputs(3570) <= not b;
    layer8_outputs(3571) <= not b;
    layer8_outputs(3572) <= b;
    layer8_outputs(3573) <= b;
    layer8_outputs(3574) <= b;
    layer8_outputs(3575) <= a or b;
    layer8_outputs(3576) <= not a;
    layer8_outputs(3577) <= not b;
    layer8_outputs(3578) <= b and not a;
    layer8_outputs(3579) <= not (a xor b);
    layer8_outputs(3580) <= a xor b;
    layer8_outputs(3581) <= not b;
    layer8_outputs(3582) <= a xor b;
    layer8_outputs(3583) <= not (a and b);
    layer8_outputs(3584) <= not (a and b);
    layer8_outputs(3585) <= b;
    layer8_outputs(3586) <= b;
    layer8_outputs(3587) <= not b or a;
    layer8_outputs(3588) <= b and not a;
    layer8_outputs(3589) <= not b;
    layer8_outputs(3590) <= not b;
    layer8_outputs(3591) <= not b;
    layer8_outputs(3592) <= not (a or b);
    layer8_outputs(3593) <= not (a and b);
    layer8_outputs(3594) <= not (a and b);
    layer8_outputs(3595) <= b;
    layer8_outputs(3596) <= not a;
    layer8_outputs(3597) <= a;
    layer8_outputs(3598) <= b;
    layer8_outputs(3599) <= b and not a;
    layer8_outputs(3600) <= not b;
    layer8_outputs(3601) <= b and not a;
    layer8_outputs(3602) <= not b;
    layer8_outputs(3603) <= a or b;
    layer8_outputs(3604) <= not (a xor b);
    layer8_outputs(3605) <= not b;
    layer8_outputs(3606) <= not b;
    layer8_outputs(3607) <= b and not a;
    layer8_outputs(3608) <= not a or b;
    layer8_outputs(3609) <= not b;
    layer8_outputs(3610) <= not b;
    layer8_outputs(3611) <= a;
    layer8_outputs(3612) <= b and not a;
    layer8_outputs(3613) <= b;
    layer8_outputs(3614) <= b;
    layer8_outputs(3615) <= not (a or b);
    layer8_outputs(3616) <= not a or b;
    layer8_outputs(3617) <= not b;
    layer8_outputs(3618) <= '0';
    layer8_outputs(3619) <= a and b;
    layer8_outputs(3620) <= not a or b;
    layer8_outputs(3621) <= b;
    layer8_outputs(3622) <= not (a xor b);
    layer8_outputs(3623) <= not b;
    layer8_outputs(3624) <= not (a or b);
    layer8_outputs(3625) <= a and b;
    layer8_outputs(3626) <= a xor b;
    layer8_outputs(3627) <= '1';
    layer8_outputs(3628) <= not b or a;
    layer8_outputs(3629) <= b and not a;
    layer8_outputs(3630) <= not b;
    layer8_outputs(3631) <= b and not a;
    layer8_outputs(3632) <= a;
    layer8_outputs(3633) <= not (a and b);
    layer8_outputs(3634) <= a;
    layer8_outputs(3635) <= not b;
    layer8_outputs(3636) <= b and not a;
    layer8_outputs(3637) <= a;
    layer8_outputs(3638) <= a and not b;
    layer8_outputs(3639) <= not b;
    layer8_outputs(3640) <= not a;
    layer8_outputs(3641) <= b;
    layer8_outputs(3642) <= not (a and b);
    layer8_outputs(3643) <= not (a and b);
    layer8_outputs(3644) <= not a;
    layer8_outputs(3645) <= not b;
    layer8_outputs(3646) <= a and not b;
    layer8_outputs(3647) <= a;
    layer8_outputs(3648) <= not b;
    layer8_outputs(3649) <= not b;
    layer8_outputs(3650) <= a or b;
    layer8_outputs(3651) <= b;
    layer8_outputs(3652) <= a xor b;
    layer8_outputs(3653) <= not b;
    layer8_outputs(3654) <= a;
    layer8_outputs(3655) <= a xor b;
    layer8_outputs(3656) <= not a;
    layer8_outputs(3657) <= b and not a;
    layer8_outputs(3658) <= a;
    layer8_outputs(3659) <= a and b;
    layer8_outputs(3660) <= not (a xor b);
    layer8_outputs(3661) <= a xor b;
    layer8_outputs(3662) <= b;
    layer8_outputs(3663) <= b and not a;
    layer8_outputs(3664) <= a xor b;
    layer8_outputs(3665) <= not b or a;
    layer8_outputs(3666) <= not a;
    layer8_outputs(3667) <= a and not b;
    layer8_outputs(3668) <= b;
    layer8_outputs(3669) <= not (a xor b);
    layer8_outputs(3670) <= a or b;
    layer8_outputs(3671) <= not b;
    layer8_outputs(3672) <= a;
    layer8_outputs(3673) <= a;
    layer8_outputs(3674) <= a and b;
    layer8_outputs(3675) <= '0';
    layer8_outputs(3676) <= not a or b;
    layer8_outputs(3677) <= not b;
    layer8_outputs(3678) <= b;
    layer8_outputs(3679) <= a;
    layer8_outputs(3680) <= a xor b;
    layer8_outputs(3681) <= not b;
    layer8_outputs(3682) <= not a or b;
    layer8_outputs(3683) <= a or b;
    layer8_outputs(3684) <= b and not a;
    layer8_outputs(3685) <= not (a or b);
    layer8_outputs(3686) <= not b or a;
    layer8_outputs(3687) <= a and b;
    layer8_outputs(3688) <= b;
    layer8_outputs(3689) <= a and not b;
    layer8_outputs(3690) <= not a;
    layer8_outputs(3691) <= a;
    layer8_outputs(3692) <= a xor b;
    layer8_outputs(3693) <= b;
    layer8_outputs(3694) <= not b or a;
    layer8_outputs(3695) <= not (a xor b);
    layer8_outputs(3696) <= not a;
    layer8_outputs(3697) <= not a;
    layer8_outputs(3698) <= not (a and b);
    layer8_outputs(3699) <= not b or a;
    layer8_outputs(3700) <= a xor b;
    layer8_outputs(3701) <= b;
    layer8_outputs(3702) <= not b;
    layer8_outputs(3703) <= a or b;
    layer8_outputs(3704) <= a or b;
    layer8_outputs(3705) <= not a or b;
    layer8_outputs(3706) <= not (a xor b);
    layer8_outputs(3707) <= a and b;
    layer8_outputs(3708) <= b and not a;
    layer8_outputs(3709) <= not (a and b);
    layer8_outputs(3710) <= not b;
    layer8_outputs(3711) <= a;
    layer8_outputs(3712) <= not b;
    layer8_outputs(3713) <= not a;
    layer8_outputs(3714) <= not b or a;
    layer8_outputs(3715) <= a and not b;
    layer8_outputs(3716) <= a and not b;
    layer8_outputs(3717) <= not b;
    layer8_outputs(3718) <= not a;
    layer8_outputs(3719) <= a and not b;
    layer8_outputs(3720) <= not (a xor b);
    layer8_outputs(3721) <= b;
    layer8_outputs(3722) <= not a or b;
    layer8_outputs(3723) <= a xor b;
    layer8_outputs(3724) <= b and not a;
    layer8_outputs(3725) <= a xor b;
    layer8_outputs(3726) <= not b or a;
    layer8_outputs(3727) <= b;
    layer8_outputs(3728) <= not (a xor b);
    layer8_outputs(3729) <= b and not a;
    layer8_outputs(3730) <= not (a and b);
    layer8_outputs(3731) <= b;
    layer8_outputs(3732) <= not a;
    layer8_outputs(3733) <= a xor b;
    layer8_outputs(3734) <= not (a xor b);
    layer8_outputs(3735) <= not a;
    layer8_outputs(3736) <= b;
    layer8_outputs(3737) <= not b;
    layer8_outputs(3738) <= b;
    layer8_outputs(3739) <= a or b;
    layer8_outputs(3740) <= not b;
    layer8_outputs(3741) <= not a;
    layer8_outputs(3742) <= not a;
    layer8_outputs(3743) <= not a or b;
    layer8_outputs(3744) <= b;
    layer8_outputs(3745) <= a xor b;
    layer8_outputs(3746) <= a and not b;
    layer8_outputs(3747) <= not (a and b);
    layer8_outputs(3748) <= not (a xor b);
    layer8_outputs(3749) <= b;
    layer8_outputs(3750) <= a xor b;
    layer8_outputs(3751) <= a and b;
    layer8_outputs(3752) <= not (a xor b);
    layer8_outputs(3753) <= not a or b;
    layer8_outputs(3754) <= not (a xor b);
    layer8_outputs(3755) <= a and b;
    layer8_outputs(3756) <= not (a xor b);
    layer8_outputs(3757) <= not (a xor b);
    layer8_outputs(3758) <= a xor b;
    layer8_outputs(3759) <= b and not a;
    layer8_outputs(3760) <= a and not b;
    layer8_outputs(3761) <= a;
    layer8_outputs(3762) <= not a;
    layer8_outputs(3763) <= not (a xor b);
    layer8_outputs(3764) <= not b;
    layer8_outputs(3765) <= not b or a;
    layer8_outputs(3766) <= b;
    layer8_outputs(3767) <= not (a xor b);
    layer8_outputs(3768) <= not b;
    layer8_outputs(3769) <= a xor b;
    layer8_outputs(3770) <= not (a and b);
    layer8_outputs(3771) <= a or b;
    layer8_outputs(3772) <= not b;
    layer8_outputs(3773) <= a and not b;
    layer8_outputs(3774) <= not a;
    layer8_outputs(3775) <= not a;
    layer8_outputs(3776) <= not a;
    layer8_outputs(3777) <= a and not b;
    layer8_outputs(3778) <= not (a and b);
    layer8_outputs(3779) <= not (a and b);
    layer8_outputs(3780) <= not (a xor b);
    layer8_outputs(3781) <= not (a xor b);
    layer8_outputs(3782) <= not b;
    layer8_outputs(3783) <= b;
    layer8_outputs(3784) <= not a;
    layer8_outputs(3785) <= b;
    layer8_outputs(3786) <= b;
    layer8_outputs(3787) <= b;
    layer8_outputs(3788) <= a or b;
    layer8_outputs(3789) <= a and b;
    layer8_outputs(3790) <= not b;
    layer8_outputs(3791) <= a and not b;
    layer8_outputs(3792) <= a and b;
    layer8_outputs(3793) <= a;
    layer8_outputs(3794) <= not (a or b);
    layer8_outputs(3795) <= not (a or b);
    layer8_outputs(3796) <= not a;
    layer8_outputs(3797) <= a;
    layer8_outputs(3798) <= b;
    layer8_outputs(3799) <= a and not b;
    layer8_outputs(3800) <= b and not a;
    layer8_outputs(3801) <= not a or b;
    layer8_outputs(3802) <= not (a xor b);
    layer8_outputs(3803) <= a xor b;
    layer8_outputs(3804) <= not a;
    layer8_outputs(3805) <= a or b;
    layer8_outputs(3806) <= b;
    layer8_outputs(3807) <= not (a and b);
    layer8_outputs(3808) <= a and b;
    layer8_outputs(3809) <= b;
    layer8_outputs(3810) <= not b;
    layer8_outputs(3811) <= not (a xor b);
    layer8_outputs(3812) <= b;
    layer8_outputs(3813) <= a xor b;
    layer8_outputs(3814) <= not b;
    layer8_outputs(3815) <= not (a xor b);
    layer8_outputs(3816) <= not b;
    layer8_outputs(3817) <= b;
    layer8_outputs(3818) <= not b;
    layer8_outputs(3819) <= a xor b;
    layer8_outputs(3820) <= not (a or b);
    layer8_outputs(3821) <= not b or a;
    layer8_outputs(3822) <= not (a and b);
    layer8_outputs(3823) <= a;
    layer8_outputs(3824) <= a and b;
    layer8_outputs(3825) <= a xor b;
    layer8_outputs(3826) <= not a;
    layer8_outputs(3827) <= not a;
    layer8_outputs(3828) <= a and b;
    layer8_outputs(3829) <= not b;
    layer8_outputs(3830) <= not b;
    layer8_outputs(3831) <= '0';
    layer8_outputs(3832) <= b;
    layer8_outputs(3833) <= a;
    layer8_outputs(3834) <= a or b;
    layer8_outputs(3835) <= a and b;
    layer8_outputs(3836) <= not a;
    layer8_outputs(3837) <= not a;
    layer8_outputs(3838) <= not a;
    layer8_outputs(3839) <= not b or a;
    layer8_outputs(3840) <= not (a xor b);
    layer8_outputs(3841) <= not (a xor b);
    layer8_outputs(3842) <= not a;
    layer8_outputs(3843) <= a;
    layer8_outputs(3844) <= not (a or b);
    layer8_outputs(3845) <= a and not b;
    layer8_outputs(3846) <= a;
    layer8_outputs(3847) <= not (a xor b);
    layer8_outputs(3848) <= b and not a;
    layer8_outputs(3849) <= not a or b;
    layer8_outputs(3850) <= not (a xor b);
    layer8_outputs(3851) <= a xor b;
    layer8_outputs(3852) <= not (a or b);
    layer8_outputs(3853) <= a and b;
    layer8_outputs(3854) <= not a or b;
    layer8_outputs(3855) <= not (a xor b);
    layer8_outputs(3856) <= a and b;
    layer8_outputs(3857) <= a or b;
    layer8_outputs(3858) <= not a;
    layer8_outputs(3859) <= a and b;
    layer8_outputs(3860) <= not (a xor b);
    layer8_outputs(3861) <= a and not b;
    layer8_outputs(3862) <= b;
    layer8_outputs(3863) <= not a;
    layer8_outputs(3864) <= a;
    layer8_outputs(3865) <= a or b;
    layer8_outputs(3866) <= b;
    layer8_outputs(3867) <= a xor b;
    layer8_outputs(3868) <= b;
    layer8_outputs(3869) <= a;
    layer8_outputs(3870) <= not (a xor b);
    layer8_outputs(3871) <= not b or a;
    layer8_outputs(3872) <= a or b;
    layer8_outputs(3873) <= a xor b;
    layer8_outputs(3874) <= not a;
    layer8_outputs(3875) <= not a;
    layer8_outputs(3876) <= a and not b;
    layer8_outputs(3877) <= not (a or b);
    layer8_outputs(3878) <= not b;
    layer8_outputs(3879) <= not a;
    layer8_outputs(3880) <= not a or b;
    layer8_outputs(3881) <= not a;
    layer8_outputs(3882) <= a;
    layer8_outputs(3883) <= a and b;
    layer8_outputs(3884) <= a or b;
    layer8_outputs(3885) <= not (a xor b);
    layer8_outputs(3886) <= not b or a;
    layer8_outputs(3887) <= not (a xor b);
    layer8_outputs(3888) <= b;
    layer8_outputs(3889) <= not a or b;
    layer8_outputs(3890) <= not b;
    layer8_outputs(3891) <= not b;
    layer8_outputs(3892) <= b;
    layer8_outputs(3893) <= a or b;
    layer8_outputs(3894) <= a xor b;
    layer8_outputs(3895) <= not (a xor b);
    layer8_outputs(3896) <= not (a xor b);
    layer8_outputs(3897) <= a or b;
    layer8_outputs(3898) <= not b;
    layer8_outputs(3899) <= not b;
    layer8_outputs(3900) <= not (a xor b);
    layer8_outputs(3901) <= not a;
    layer8_outputs(3902) <= not a;
    layer8_outputs(3903) <= not (a xor b);
    layer8_outputs(3904) <= not (a xor b);
    layer8_outputs(3905) <= not (a and b);
    layer8_outputs(3906) <= not b or a;
    layer8_outputs(3907) <= b and not a;
    layer8_outputs(3908) <= a;
    layer8_outputs(3909) <= a or b;
    layer8_outputs(3910) <= not (a or b);
    layer8_outputs(3911) <= not b;
    layer8_outputs(3912) <= not b;
    layer8_outputs(3913) <= not a or b;
    layer8_outputs(3914) <= not (a xor b);
    layer8_outputs(3915) <= b and not a;
    layer8_outputs(3916) <= not (a xor b);
    layer8_outputs(3917) <= a xor b;
    layer8_outputs(3918) <= a;
    layer8_outputs(3919) <= not b;
    layer8_outputs(3920) <= b;
    layer8_outputs(3921) <= not (a xor b);
    layer8_outputs(3922) <= b;
    layer8_outputs(3923) <= a xor b;
    layer8_outputs(3924) <= not (a xor b);
    layer8_outputs(3925) <= a xor b;
    layer8_outputs(3926) <= not b;
    layer8_outputs(3927) <= b;
    layer8_outputs(3928) <= not (a xor b);
    layer8_outputs(3929) <= not (a xor b);
    layer8_outputs(3930) <= not a;
    layer8_outputs(3931) <= a xor b;
    layer8_outputs(3932) <= a;
    layer8_outputs(3933) <= not b;
    layer8_outputs(3934) <= not a or b;
    layer8_outputs(3935) <= a and b;
    layer8_outputs(3936) <= a xor b;
    layer8_outputs(3937) <= not a;
    layer8_outputs(3938) <= b and not a;
    layer8_outputs(3939) <= b and not a;
    layer8_outputs(3940) <= a;
    layer8_outputs(3941) <= a xor b;
    layer8_outputs(3942) <= b and not a;
    layer8_outputs(3943) <= not (a or b);
    layer8_outputs(3944) <= not a;
    layer8_outputs(3945) <= a;
    layer8_outputs(3946) <= a and b;
    layer8_outputs(3947) <= b;
    layer8_outputs(3948) <= a;
    layer8_outputs(3949) <= not b or a;
    layer8_outputs(3950) <= not (a and b);
    layer8_outputs(3951) <= not b;
    layer8_outputs(3952) <= not a;
    layer8_outputs(3953) <= not b or a;
    layer8_outputs(3954) <= a xor b;
    layer8_outputs(3955) <= a xor b;
    layer8_outputs(3956) <= not (a and b);
    layer8_outputs(3957) <= b;
    layer8_outputs(3958) <= b;
    layer8_outputs(3959) <= not b;
    layer8_outputs(3960) <= a xor b;
    layer8_outputs(3961) <= not a;
    layer8_outputs(3962) <= not b;
    layer8_outputs(3963) <= not b;
    layer8_outputs(3964) <= not b;
    layer8_outputs(3965) <= not b;
    layer8_outputs(3966) <= a and not b;
    layer8_outputs(3967) <= a and not b;
    layer8_outputs(3968) <= not a or b;
    layer8_outputs(3969) <= not a or b;
    layer8_outputs(3970) <= a and not b;
    layer8_outputs(3971) <= a xor b;
    layer8_outputs(3972) <= a;
    layer8_outputs(3973) <= not b;
    layer8_outputs(3974) <= a or b;
    layer8_outputs(3975) <= a and b;
    layer8_outputs(3976) <= b and not a;
    layer8_outputs(3977) <= a;
    layer8_outputs(3978) <= a and not b;
    layer8_outputs(3979) <= not (a and b);
    layer8_outputs(3980) <= not b or a;
    layer8_outputs(3981) <= a xor b;
    layer8_outputs(3982) <= b;
    layer8_outputs(3983) <= not (a xor b);
    layer8_outputs(3984) <= a xor b;
    layer8_outputs(3985) <= not (a xor b);
    layer8_outputs(3986) <= a;
    layer8_outputs(3987) <= b and not a;
    layer8_outputs(3988) <= not a;
    layer8_outputs(3989) <= not b;
    layer8_outputs(3990) <= a xor b;
    layer8_outputs(3991) <= a xor b;
    layer8_outputs(3992) <= b;
    layer8_outputs(3993) <= a or b;
    layer8_outputs(3994) <= not (a xor b);
    layer8_outputs(3995) <= b;
    layer8_outputs(3996) <= a or b;
    layer8_outputs(3997) <= a xor b;
    layer8_outputs(3998) <= a and not b;
    layer8_outputs(3999) <= '1';
    layer8_outputs(4000) <= not a;
    layer8_outputs(4001) <= a and b;
    layer8_outputs(4002) <= a;
    layer8_outputs(4003) <= not (a xor b);
    layer8_outputs(4004) <= not b or a;
    layer8_outputs(4005) <= not b;
    layer8_outputs(4006) <= not a;
    layer8_outputs(4007) <= not a;
    layer8_outputs(4008) <= not b;
    layer8_outputs(4009) <= b;
    layer8_outputs(4010) <= not b or a;
    layer8_outputs(4011) <= b;
    layer8_outputs(4012) <= a xor b;
    layer8_outputs(4013) <= not b;
    layer8_outputs(4014) <= a xor b;
    layer8_outputs(4015) <= b;
    layer8_outputs(4016) <= a;
    layer8_outputs(4017) <= not a or b;
    layer8_outputs(4018) <= not a;
    layer8_outputs(4019) <= not a;
    layer8_outputs(4020) <= a or b;
    layer8_outputs(4021) <= a xor b;
    layer8_outputs(4022) <= b;
    layer8_outputs(4023) <= a;
    layer8_outputs(4024) <= a xor b;
    layer8_outputs(4025) <= not (a xor b);
    layer8_outputs(4026) <= b;
    layer8_outputs(4027) <= '0';
    layer8_outputs(4028) <= not (a xor b);
    layer8_outputs(4029) <= not (a xor b);
    layer8_outputs(4030) <= b;
    layer8_outputs(4031) <= not (a xor b);
    layer8_outputs(4032) <= a;
    layer8_outputs(4033) <= not (a or b);
    layer8_outputs(4034) <= a;
    layer8_outputs(4035) <= not (a and b);
    layer8_outputs(4036) <= a xor b;
    layer8_outputs(4037) <= not (a or b);
    layer8_outputs(4038) <= not a;
    layer8_outputs(4039) <= not a;
    layer8_outputs(4040) <= a xor b;
    layer8_outputs(4041) <= a;
    layer8_outputs(4042) <= not (a xor b);
    layer8_outputs(4043) <= a xor b;
    layer8_outputs(4044) <= a;
    layer8_outputs(4045) <= a;
    layer8_outputs(4046) <= not b;
    layer8_outputs(4047) <= a;
    layer8_outputs(4048) <= not a;
    layer8_outputs(4049) <= a;
    layer8_outputs(4050) <= not b;
    layer8_outputs(4051) <= not (a and b);
    layer8_outputs(4052) <= not b;
    layer8_outputs(4053) <= not b;
    layer8_outputs(4054) <= not (a xor b);
    layer8_outputs(4055) <= a xor b;
    layer8_outputs(4056) <= b;
    layer8_outputs(4057) <= not a or b;
    layer8_outputs(4058) <= b and not a;
    layer8_outputs(4059) <= not b or a;
    layer8_outputs(4060) <= a xor b;
    layer8_outputs(4061) <= not a or b;
    layer8_outputs(4062) <= b;
    layer8_outputs(4063) <= a and not b;
    layer8_outputs(4064) <= a;
    layer8_outputs(4065) <= a xor b;
    layer8_outputs(4066) <= not b;
    layer8_outputs(4067) <= b;
    layer8_outputs(4068) <= not a;
    layer8_outputs(4069) <= b;
    layer8_outputs(4070) <= not b;
    layer8_outputs(4071) <= not (a xor b);
    layer8_outputs(4072) <= not (a or b);
    layer8_outputs(4073) <= not b;
    layer8_outputs(4074) <= '0';
    layer8_outputs(4075) <= a xor b;
    layer8_outputs(4076) <= not a;
    layer8_outputs(4077) <= b;
    layer8_outputs(4078) <= not (a or b);
    layer8_outputs(4079) <= a xor b;
    layer8_outputs(4080) <= a;
    layer8_outputs(4081) <= not (a xor b);
    layer8_outputs(4082) <= a xor b;
    layer8_outputs(4083) <= a and not b;
    layer8_outputs(4084) <= not a or b;
    layer8_outputs(4085) <= not b;
    layer8_outputs(4086) <= b and not a;
    layer8_outputs(4087) <= not (a and b);
    layer8_outputs(4088) <= not (a and b);
    layer8_outputs(4089) <= a xor b;
    layer8_outputs(4090) <= not (a and b);
    layer8_outputs(4091) <= not b or a;
    layer8_outputs(4092) <= not a;
    layer8_outputs(4093) <= b;
    layer8_outputs(4094) <= a;
    layer8_outputs(4095) <= not (a xor b);
    layer8_outputs(4096) <= a and b;
    layer8_outputs(4097) <= a;
    layer8_outputs(4098) <= not a;
    layer8_outputs(4099) <= not b;
    layer8_outputs(4100) <= b;
    layer8_outputs(4101) <= not a;
    layer8_outputs(4102) <= b;
    layer8_outputs(4103) <= not b;
    layer8_outputs(4104) <= b;
    layer8_outputs(4105) <= not a or b;
    layer8_outputs(4106) <= not a;
    layer8_outputs(4107) <= not b;
    layer8_outputs(4108) <= a xor b;
    layer8_outputs(4109) <= a and b;
    layer8_outputs(4110) <= not b or a;
    layer8_outputs(4111) <= not a;
    layer8_outputs(4112) <= b and not a;
    layer8_outputs(4113) <= b;
    layer8_outputs(4114) <= b and not a;
    layer8_outputs(4115) <= a xor b;
    layer8_outputs(4116) <= not a;
    layer8_outputs(4117) <= b;
    layer8_outputs(4118) <= a and b;
    layer8_outputs(4119) <= not a;
    layer8_outputs(4120) <= b;
    layer8_outputs(4121) <= a xor b;
    layer8_outputs(4122) <= '0';
    layer8_outputs(4123) <= not a;
    layer8_outputs(4124) <= not a or b;
    layer8_outputs(4125) <= not (a xor b);
    layer8_outputs(4126) <= a xor b;
    layer8_outputs(4127) <= b;
    layer8_outputs(4128) <= not a or b;
    layer8_outputs(4129) <= not a;
    layer8_outputs(4130) <= not b;
    layer8_outputs(4131) <= a and b;
    layer8_outputs(4132) <= a and not b;
    layer8_outputs(4133) <= a;
    layer8_outputs(4134) <= not b or a;
    layer8_outputs(4135) <= not b;
    layer8_outputs(4136) <= a and b;
    layer8_outputs(4137) <= b;
    layer8_outputs(4138) <= not b or a;
    layer8_outputs(4139) <= a and not b;
    layer8_outputs(4140) <= not (a or b);
    layer8_outputs(4141) <= not a;
    layer8_outputs(4142) <= a;
    layer8_outputs(4143) <= a and not b;
    layer8_outputs(4144) <= not (a or b);
    layer8_outputs(4145) <= not b or a;
    layer8_outputs(4146) <= a and b;
    layer8_outputs(4147) <= not a;
    layer8_outputs(4148) <= not b;
    layer8_outputs(4149) <= not (a and b);
    layer8_outputs(4150) <= b;
    layer8_outputs(4151) <= not (a xor b);
    layer8_outputs(4152) <= b;
    layer8_outputs(4153) <= b and not a;
    layer8_outputs(4154) <= not a;
    layer8_outputs(4155) <= a;
    layer8_outputs(4156) <= not b;
    layer8_outputs(4157) <= not (a xor b);
    layer8_outputs(4158) <= not (a xor b);
    layer8_outputs(4159) <= a;
    layer8_outputs(4160) <= a;
    layer8_outputs(4161) <= a xor b;
    layer8_outputs(4162) <= a;
    layer8_outputs(4163) <= a;
    layer8_outputs(4164) <= not a;
    layer8_outputs(4165) <= not b;
    layer8_outputs(4166) <= b and not a;
    layer8_outputs(4167) <= a and not b;
    layer8_outputs(4168) <= not a;
    layer8_outputs(4169) <= not (a xor b);
    layer8_outputs(4170) <= a and b;
    layer8_outputs(4171) <= a xor b;
    layer8_outputs(4172) <= a;
    layer8_outputs(4173) <= a;
    layer8_outputs(4174) <= not (a and b);
    layer8_outputs(4175) <= a;
    layer8_outputs(4176) <= not b;
    layer8_outputs(4177) <= a;
    layer8_outputs(4178) <= a;
    layer8_outputs(4179) <= not a;
    layer8_outputs(4180) <= a and b;
    layer8_outputs(4181) <= a xor b;
    layer8_outputs(4182) <= not a;
    layer8_outputs(4183) <= b and not a;
    layer8_outputs(4184) <= not b;
    layer8_outputs(4185) <= not (a and b);
    layer8_outputs(4186) <= not (a or b);
    layer8_outputs(4187) <= not b;
    layer8_outputs(4188) <= b;
    layer8_outputs(4189) <= a and b;
    layer8_outputs(4190) <= a xor b;
    layer8_outputs(4191) <= not (a or b);
    layer8_outputs(4192) <= not b;
    layer8_outputs(4193) <= not b or a;
    layer8_outputs(4194) <= not (a xor b);
    layer8_outputs(4195) <= not b or a;
    layer8_outputs(4196) <= a and not b;
    layer8_outputs(4197) <= not a or b;
    layer8_outputs(4198) <= a xor b;
    layer8_outputs(4199) <= not (a or b);
    layer8_outputs(4200) <= a or b;
    layer8_outputs(4201) <= not (a xor b);
    layer8_outputs(4202) <= not b;
    layer8_outputs(4203) <= a and not b;
    layer8_outputs(4204) <= not b;
    layer8_outputs(4205) <= not (a xor b);
    layer8_outputs(4206) <= a xor b;
    layer8_outputs(4207) <= b;
    layer8_outputs(4208) <= a;
    layer8_outputs(4209) <= b;
    layer8_outputs(4210) <= not (a xor b);
    layer8_outputs(4211) <= not (a xor b);
    layer8_outputs(4212) <= b;
    layer8_outputs(4213) <= a;
    layer8_outputs(4214) <= b and not a;
    layer8_outputs(4215) <= a or b;
    layer8_outputs(4216) <= a;
    layer8_outputs(4217) <= b;
    layer8_outputs(4218) <= not b;
    layer8_outputs(4219) <= a and not b;
    layer8_outputs(4220) <= a and b;
    layer8_outputs(4221) <= not (a xor b);
    layer8_outputs(4222) <= not (a xor b);
    layer8_outputs(4223) <= a xor b;
    layer8_outputs(4224) <= not (a and b);
    layer8_outputs(4225) <= a;
    layer8_outputs(4226) <= not (a xor b);
    layer8_outputs(4227) <= not a or b;
    layer8_outputs(4228) <= not (a or b);
    layer8_outputs(4229) <= not (a and b);
    layer8_outputs(4230) <= a xor b;
    layer8_outputs(4231) <= not a or b;
    layer8_outputs(4232) <= a xor b;
    layer8_outputs(4233) <= b;
    layer8_outputs(4234) <= b and not a;
    layer8_outputs(4235) <= a xor b;
    layer8_outputs(4236) <= not (a xor b);
    layer8_outputs(4237) <= not (a xor b);
    layer8_outputs(4238) <= a and b;
    layer8_outputs(4239) <= not a;
    layer8_outputs(4240) <= not a or b;
    layer8_outputs(4241) <= not b;
    layer8_outputs(4242) <= b;
    layer8_outputs(4243) <= b;
    layer8_outputs(4244) <= not b;
    layer8_outputs(4245) <= not a or b;
    layer8_outputs(4246) <= a;
    layer8_outputs(4247) <= not b;
    layer8_outputs(4248) <= not b;
    layer8_outputs(4249) <= b;
    layer8_outputs(4250) <= not a;
    layer8_outputs(4251) <= not a or b;
    layer8_outputs(4252) <= not a;
    layer8_outputs(4253) <= not b;
    layer8_outputs(4254) <= not b;
    layer8_outputs(4255) <= b and not a;
    layer8_outputs(4256) <= a or b;
    layer8_outputs(4257) <= b and not a;
    layer8_outputs(4258) <= not b;
    layer8_outputs(4259) <= b;
    layer8_outputs(4260) <= a and not b;
    layer8_outputs(4261) <= not (a xor b);
    layer8_outputs(4262) <= a;
    layer8_outputs(4263) <= a and not b;
    layer8_outputs(4264) <= not a or b;
    layer8_outputs(4265) <= not a;
    layer8_outputs(4266) <= a and not b;
    layer8_outputs(4267) <= b and not a;
    layer8_outputs(4268) <= not (a xor b);
    layer8_outputs(4269) <= a xor b;
    layer8_outputs(4270) <= not a;
    layer8_outputs(4271) <= a xor b;
    layer8_outputs(4272) <= not (a xor b);
    layer8_outputs(4273) <= not a or b;
    layer8_outputs(4274) <= a;
    layer8_outputs(4275) <= '1';
    layer8_outputs(4276) <= b;
    layer8_outputs(4277) <= a and b;
    layer8_outputs(4278) <= not (a and b);
    layer8_outputs(4279) <= a and not b;
    layer8_outputs(4280) <= not a;
    layer8_outputs(4281) <= not (a or b);
    layer8_outputs(4282) <= not (a or b);
    layer8_outputs(4283) <= a xor b;
    layer8_outputs(4284) <= not (a xor b);
    layer8_outputs(4285) <= not (a xor b);
    layer8_outputs(4286) <= not (a or b);
    layer8_outputs(4287) <= a;
    layer8_outputs(4288) <= b;
    layer8_outputs(4289) <= not b;
    layer8_outputs(4290) <= a or b;
    layer8_outputs(4291) <= b;
    layer8_outputs(4292) <= not b or a;
    layer8_outputs(4293) <= a or b;
    layer8_outputs(4294) <= a xor b;
    layer8_outputs(4295) <= a;
    layer8_outputs(4296) <= not a;
    layer8_outputs(4297) <= b and not a;
    layer8_outputs(4298) <= not b;
    layer8_outputs(4299) <= '1';
    layer8_outputs(4300) <= not a or b;
    layer8_outputs(4301) <= a or b;
    layer8_outputs(4302) <= a and b;
    layer8_outputs(4303) <= b;
    layer8_outputs(4304) <= not a;
    layer8_outputs(4305) <= not (a xor b);
    layer8_outputs(4306) <= not (a and b);
    layer8_outputs(4307) <= a xor b;
    layer8_outputs(4308) <= a and b;
    layer8_outputs(4309) <= b;
    layer8_outputs(4310) <= not a;
    layer8_outputs(4311) <= a;
    layer8_outputs(4312) <= b;
    layer8_outputs(4313) <= not a or b;
    layer8_outputs(4314) <= not (a xor b);
    layer8_outputs(4315) <= a;
    layer8_outputs(4316) <= a xor b;
    layer8_outputs(4317) <= a xor b;
    layer8_outputs(4318) <= a;
    layer8_outputs(4319) <= a and not b;
    layer8_outputs(4320) <= b;
    layer8_outputs(4321) <= not b or a;
    layer8_outputs(4322) <= not b;
    layer8_outputs(4323) <= not b or a;
    layer8_outputs(4324) <= not a;
    layer8_outputs(4325) <= b;
    layer8_outputs(4326) <= not a;
    layer8_outputs(4327) <= b and not a;
    layer8_outputs(4328) <= not (a xor b);
    layer8_outputs(4329) <= not a;
    layer8_outputs(4330) <= not (a xor b);
    layer8_outputs(4331) <= not b or a;
    layer8_outputs(4332) <= b;
    layer8_outputs(4333) <= a xor b;
    layer8_outputs(4334) <= a;
    layer8_outputs(4335) <= a and not b;
    layer8_outputs(4336) <= b and not a;
    layer8_outputs(4337) <= b;
    layer8_outputs(4338) <= a and b;
    layer8_outputs(4339) <= a xor b;
    layer8_outputs(4340) <= a;
    layer8_outputs(4341) <= a and b;
    layer8_outputs(4342) <= b;
    layer8_outputs(4343) <= a xor b;
    layer8_outputs(4344) <= a or b;
    layer8_outputs(4345) <= not a;
    layer8_outputs(4346) <= not (a xor b);
    layer8_outputs(4347) <= a;
    layer8_outputs(4348) <= b;
    layer8_outputs(4349) <= a or b;
    layer8_outputs(4350) <= a xor b;
    layer8_outputs(4351) <= not (a xor b);
    layer8_outputs(4352) <= not (a or b);
    layer8_outputs(4353) <= not (a and b);
    layer8_outputs(4354) <= a xor b;
    layer8_outputs(4355) <= not b;
    layer8_outputs(4356) <= not a;
    layer8_outputs(4357) <= a xor b;
    layer8_outputs(4358) <= not (a and b);
    layer8_outputs(4359) <= not b;
    layer8_outputs(4360) <= b;
    layer8_outputs(4361) <= not a or b;
    layer8_outputs(4362) <= a;
    layer8_outputs(4363) <= not b;
    layer8_outputs(4364) <= not (a xor b);
    layer8_outputs(4365) <= a or b;
    layer8_outputs(4366) <= not b;
    layer8_outputs(4367) <= not a;
    layer8_outputs(4368) <= a;
    layer8_outputs(4369) <= b and not a;
    layer8_outputs(4370) <= a and not b;
    layer8_outputs(4371) <= a xor b;
    layer8_outputs(4372) <= b and not a;
    layer8_outputs(4373) <= a xor b;
    layer8_outputs(4374) <= not (a or b);
    layer8_outputs(4375) <= a;
    layer8_outputs(4376) <= not (a or b);
    layer8_outputs(4377) <= not b or a;
    layer8_outputs(4378) <= a and b;
    layer8_outputs(4379) <= a xor b;
    layer8_outputs(4380) <= a;
    layer8_outputs(4381) <= a or b;
    layer8_outputs(4382) <= not a;
    layer8_outputs(4383) <= not a;
    layer8_outputs(4384) <= not (a and b);
    layer8_outputs(4385) <= b and not a;
    layer8_outputs(4386) <= a;
    layer8_outputs(4387) <= a xor b;
    layer8_outputs(4388) <= not (a xor b);
    layer8_outputs(4389) <= not (a xor b);
    layer8_outputs(4390) <= '1';
    layer8_outputs(4391) <= a xor b;
    layer8_outputs(4392) <= a xor b;
    layer8_outputs(4393) <= not (a xor b);
    layer8_outputs(4394) <= not (a xor b);
    layer8_outputs(4395) <= not (a xor b);
    layer8_outputs(4396) <= b;
    layer8_outputs(4397) <= a and b;
    layer8_outputs(4398) <= a and b;
    layer8_outputs(4399) <= b;
    layer8_outputs(4400) <= not b;
    layer8_outputs(4401) <= b;
    layer8_outputs(4402) <= a;
    layer8_outputs(4403) <= not a or b;
    layer8_outputs(4404) <= a and not b;
    layer8_outputs(4405) <= a and b;
    layer8_outputs(4406) <= b;
    layer8_outputs(4407) <= b;
    layer8_outputs(4408) <= a xor b;
    layer8_outputs(4409) <= b and not a;
    layer8_outputs(4410) <= not b;
    layer8_outputs(4411) <= not b;
    layer8_outputs(4412) <= not b;
    layer8_outputs(4413) <= not (a and b);
    layer8_outputs(4414) <= a;
    layer8_outputs(4415) <= b;
    layer8_outputs(4416) <= not a;
    layer8_outputs(4417) <= a xor b;
    layer8_outputs(4418) <= not b;
    layer8_outputs(4419) <= a;
    layer8_outputs(4420) <= a xor b;
    layer8_outputs(4421) <= a xor b;
    layer8_outputs(4422) <= not a;
    layer8_outputs(4423) <= b and not a;
    layer8_outputs(4424) <= not (a xor b);
    layer8_outputs(4425) <= a;
    layer8_outputs(4426) <= b;
    layer8_outputs(4427) <= not (a or b);
    layer8_outputs(4428) <= not (a and b);
    layer8_outputs(4429) <= a;
    layer8_outputs(4430) <= a xor b;
    layer8_outputs(4431) <= not (a xor b);
    layer8_outputs(4432) <= b and not a;
    layer8_outputs(4433) <= a;
    layer8_outputs(4434) <= not (a or b);
    layer8_outputs(4435) <= a;
    layer8_outputs(4436) <= not (a and b);
    layer8_outputs(4437) <= a xor b;
    layer8_outputs(4438) <= a and b;
    layer8_outputs(4439) <= a;
    layer8_outputs(4440) <= not a;
    layer8_outputs(4441) <= b;
    layer8_outputs(4442) <= a;
    layer8_outputs(4443) <= not a or b;
    layer8_outputs(4444) <= a and not b;
    layer8_outputs(4445) <= not a;
    layer8_outputs(4446) <= a xor b;
    layer8_outputs(4447) <= a;
    layer8_outputs(4448) <= b;
    layer8_outputs(4449) <= b;
    layer8_outputs(4450) <= not a;
    layer8_outputs(4451) <= a xor b;
    layer8_outputs(4452) <= a;
    layer8_outputs(4453) <= not b;
    layer8_outputs(4454) <= b;
    layer8_outputs(4455) <= not (a and b);
    layer8_outputs(4456) <= a or b;
    layer8_outputs(4457) <= a xor b;
    layer8_outputs(4458) <= not a;
    layer8_outputs(4459) <= not (a and b);
    layer8_outputs(4460) <= not a;
    layer8_outputs(4461) <= not (a and b);
    layer8_outputs(4462) <= not a or b;
    layer8_outputs(4463) <= not a;
    layer8_outputs(4464) <= a;
    layer8_outputs(4465) <= b and not a;
    layer8_outputs(4466) <= not (a xor b);
    layer8_outputs(4467) <= b;
    layer8_outputs(4468) <= b;
    layer8_outputs(4469) <= not b;
    layer8_outputs(4470) <= not (a xor b);
    layer8_outputs(4471) <= not a or b;
    layer8_outputs(4472) <= b;
    layer8_outputs(4473) <= b;
    layer8_outputs(4474) <= a and not b;
    layer8_outputs(4475) <= a;
    layer8_outputs(4476) <= b;
    layer8_outputs(4477) <= not (a or b);
    layer8_outputs(4478) <= a xor b;
    layer8_outputs(4479) <= a and not b;
    layer8_outputs(4480) <= b;
    layer8_outputs(4481) <= a and b;
    layer8_outputs(4482) <= not b;
    layer8_outputs(4483) <= a xor b;
    layer8_outputs(4484) <= not (a xor b);
    layer8_outputs(4485) <= a xor b;
    layer8_outputs(4486) <= not b;
    layer8_outputs(4487) <= a and b;
    layer8_outputs(4488) <= a xor b;
    layer8_outputs(4489) <= a and b;
    layer8_outputs(4490) <= a xor b;
    layer8_outputs(4491) <= a and not b;
    layer8_outputs(4492) <= not b;
    layer8_outputs(4493) <= a and b;
    layer8_outputs(4494) <= a xor b;
    layer8_outputs(4495) <= not a;
    layer8_outputs(4496) <= not a;
    layer8_outputs(4497) <= not a or b;
    layer8_outputs(4498) <= not (a and b);
    layer8_outputs(4499) <= b;
    layer8_outputs(4500) <= not b;
    layer8_outputs(4501) <= a xor b;
    layer8_outputs(4502) <= a;
    layer8_outputs(4503) <= not b;
    layer8_outputs(4504) <= a and b;
    layer8_outputs(4505) <= not (a xor b);
    layer8_outputs(4506) <= not a;
    layer8_outputs(4507) <= not b;
    layer8_outputs(4508) <= not b;
    layer8_outputs(4509) <= not a or b;
    layer8_outputs(4510) <= not b;
    layer8_outputs(4511) <= not a;
    layer8_outputs(4512) <= a xor b;
    layer8_outputs(4513) <= a xor b;
    layer8_outputs(4514) <= a xor b;
    layer8_outputs(4515) <= not b;
    layer8_outputs(4516) <= b;
    layer8_outputs(4517) <= not b or a;
    layer8_outputs(4518) <= a and not b;
    layer8_outputs(4519) <= a;
    layer8_outputs(4520) <= a xor b;
    layer8_outputs(4521) <= not b;
    layer8_outputs(4522) <= a;
    layer8_outputs(4523) <= b;
    layer8_outputs(4524) <= a and not b;
    layer8_outputs(4525) <= a xor b;
    layer8_outputs(4526) <= not (a xor b);
    layer8_outputs(4527) <= not b;
    layer8_outputs(4528) <= not (a xor b);
    layer8_outputs(4529) <= a;
    layer8_outputs(4530) <= a;
    layer8_outputs(4531) <= not (a xor b);
    layer8_outputs(4532) <= a;
    layer8_outputs(4533) <= not a or b;
    layer8_outputs(4534) <= not (a xor b);
    layer8_outputs(4535) <= not (a xor b);
    layer8_outputs(4536) <= b;
    layer8_outputs(4537) <= not (a xor b);
    layer8_outputs(4538) <= a;
    layer8_outputs(4539) <= not a;
    layer8_outputs(4540) <= a;
    layer8_outputs(4541) <= not (a or b);
    layer8_outputs(4542) <= b;
    layer8_outputs(4543) <= not a;
    layer8_outputs(4544) <= a or b;
    layer8_outputs(4545) <= b;
    layer8_outputs(4546) <= not a;
    layer8_outputs(4547) <= not (a xor b);
    layer8_outputs(4548) <= a xor b;
    layer8_outputs(4549) <= not a;
    layer8_outputs(4550) <= not b;
    layer8_outputs(4551) <= a;
    layer8_outputs(4552) <= not a;
    layer8_outputs(4553) <= not b;
    layer8_outputs(4554) <= a xor b;
    layer8_outputs(4555) <= a;
    layer8_outputs(4556) <= not (a xor b);
    layer8_outputs(4557) <= b and not a;
    layer8_outputs(4558) <= not a;
    layer8_outputs(4559) <= a xor b;
    layer8_outputs(4560) <= b;
    layer8_outputs(4561) <= not (a and b);
    layer8_outputs(4562) <= a and b;
    layer8_outputs(4563) <= not b;
    layer8_outputs(4564) <= not a;
    layer8_outputs(4565) <= not b or a;
    layer8_outputs(4566) <= a xor b;
    layer8_outputs(4567) <= a xor b;
    layer8_outputs(4568) <= not b;
    layer8_outputs(4569) <= not (a xor b);
    layer8_outputs(4570) <= b;
    layer8_outputs(4571) <= a;
    layer8_outputs(4572) <= not (a or b);
    layer8_outputs(4573) <= not b;
    layer8_outputs(4574) <= not (a xor b);
    layer8_outputs(4575) <= not a;
    layer8_outputs(4576) <= b;
    layer8_outputs(4577) <= not (a and b);
    layer8_outputs(4578) <= not (a xor b);
    layer8_outputs(4579) <= not a;
    layer8_outputs(4580) <= b;
    layer8_outputs(4581) <= not (a xor b);
    layer8_outputs(4582) <= a;
    layer8_outputs(4583) <= not (a or b);
    layer8_outputs(4584) <= a;
    layer8_outputs(4585) <= not (a xor b);
    layer8_outputs(4586) <= not b or a;
    layer8_outputs(4587) <= a and not b;
    layer8_outputs(4588) <= not (a xor b);
    layer8_outputs(4589) <= b and not a;
    layer8_outputs(4590) <= '1';
    layer8_outputs(4591) <= a and not b;
    layer8_outputs(4592) <= a xor b;
    layer8_outputs(4593) <= not b;
    layer8_outputs(4594) <= not (a or b);
    layer8_outputs(4595) <= a and b;
    layer8_outputs(4596) <= a or b;
    layer8_outputs(4597) <= not b;
    layer8_outputs(4598) <= not (a and b);
    layer8_outputs(4599) <= not b;
    layer8_outputs(4600) <= not (a and b);
    layer8_outputs(4601) <= not (a or b);
    layer8_outputs(4602) <= not (a xor b);
    layer8_outputs(4603) <= a and not b;
    layer8_outputs(4604) <= not (a or b);
    layer8_outputs(4605) <= not (a xor b);
    layer8_outputs(4606) <= a xor b;
    layer8_outputs(4607) <= a xor b;
    layer8_outputs(4608) <= b;
    layer8_outputs(4609) <= not (a xor b);
    layer8_outputs(4610) <= not a;
    layer8_outputs(4611) <= not a;
    layer8_outputs(4612) <= not a;
    layer8_outputs(4613) <= a;
    layer8_outputs(4614) <= not a;
    layer8_outputs(4615) <= not b;
    layer8_outputs(4616) <= not a or b;
    layer8_outputs(4617) <= not a;
    layer8_outputs(4618) <= b and not a;
    layer8_outputs(4619) <= not b or a;
    layer8_outputs(4620) <= not a or b;
    layer8_outputs(4621) <= not b;
    layer8_outputs(4622) <= not b;
    layer8_outputs(4623) <= a xor b;
    layer8_outputs(4624) <= a;
    layer8_outputs(4625) <= a;
    layer8_outputs(4626) <= not (a or b);
    layer8_outputs(4627) <= b;
    layer8_outputs(4628) <= not b;
    layer8_outputs(4629) <= a xor b;
    layer8_outputs(4630) <= a;
    layer8_outputs(4631) <= b;
    layer8_outputs(4632) <= not a;
    layer8_outputs(4633) <= not a;
    layer8_outputs(4634) <= b;
    layer8_outputs(4635) <= not b;
    layer8_outputs(4636) <= not (a xor b);
    layer8_outputs(4637) <= not a;
    layer8_outputs(4638) <= not a;
    layer8_outputs(4639) <= not (a xor b);
    layer8_outputs(4640) <= not (a xor b);
    layer8_outputs(4641) <= a xor b;
    layer8_outputs(4642) <= b and not a;
    layer8_outputs(4643) <= not a;
    layer8_outputs(4644) <= a;
    layer8_outputs(4645) <= a;
    layer8_outputs(4646) <= a and b;
    layer8_outputs(4647) <= a xor b;
    layer8_outputs(4648) <= a;
    layer8_outputs(4649) <= a;
    layer8_outputs(4650) <= not a;
    layer8_outputs(4651) <= b and not a;
    layer8_outputs(4652) <= b;
    layer8_outputs(4653) <= not a;
    layer8_outputs(4654) <= not a;
    layer8_outputs(4655) <= '0';
    layer8_outputs(4656) <= a and b;
    layer8_outputs(4657) <= b;
    layer8_outputs(4658) <= a and not b;
    layer8_outputs(4659) <= b;
    layer8_outputs(4660) <= not a;
    layer8_outputs(4661) <= b and not a;
    layer8_outputs(4662) <= not b;
    layer8_outputs(4663) <= a and not b;
    layer8_outputs(4664) <= b and not a;
    layer8_outputs(4665) <= a xor b;
    layer8_outputs(4666) <= a and b;
    layer8_outputs(4667) <= a and b;
    layer8_outputs(4668) <= not b;
    layer8_outputs(4669) <= a;
    layer8_outputs(4670) <= a xor b;
    layer8_outputs(4671) <= not (a xor b);
    layer8_outputs(4672) <= not b;
    layer8_outputs(4673) <= not b;
    layer8_outputs(4674) <= not b;
    layer8_outputs(4675) <= not b;
    layer8_outputs(4676) <= not b;
    layer8_outputs(4677) <= not (a and b);
    layer8_outputs(4678) <= a;
    layer8_outputs(4679) <= not b or a;
    layer8_outputs(4680) <= a xor b;
    layer8_outputs(4681) <= not a;
    layer8_outputs(4682) <= a and b;
    layer8_outputs(4683) <= a xor b;
    layer8_outputs(4684) <= not (a xor b);
    layer8_outputs(4685) <= a;
    layer8_outputs(4686) <= not a or b;
    layer8_outputs(4687) <= a xor b;
    layer8_outputs(4688) <= a or b;
    layer8_outputs(4689) <= b;
    layer8_outputs(4690) <= not (a and b);
    layer8_outputs(4691) <= a and b;
    layer8_outputs(4692) <= not (a xor b);
    layer8_outputs(4693) <= a and not b;
    layer8_outputs(4694) <= not a;
    layer8_outputs(4695) <= not (a xor b);
    layer8_outputs(4696) <= b and not a;
    layer8_outputs(4697) <= a and not b;
    layer8_outputs(4698) <= a xor b;
    layer8_outputs(4699) <= b;
    layer8_outputs(4700) <= not (a xor b);
    layer8_outputs(4701) <= not (a xor b);
    layer8_outputs(4702) <= b;
    layer8_outputs(4703) <= not a;
    layer8_outputs(4704) <= a xor b;
    layer8_outputs(4705) <= a xor b;
    layer8_outputs(4706) <= a or b;
    layer8_outputs(4707) <= not b;
    layer8_outputs(4708) <= a xor b;
    layer8_outputs(4709) <= a;
    layer8_outputs(4710) <= b;
    layer8_outputs(4711) <= a;
    layer8_outputs(4712) <= not a or b;
    layer8_outputs(4713) <= a xor b;
    layer8_outputs(4714) <= not a;
    layer8_outputs(4715) <= not (a or b);
    layer8_outputs(4716) <= not (a and b);
    layer8_outputs(4717) <= b and not a;
    layer8_outputs(4718) <= not (a or b);
    layer8_outputs(4719) <= a or b;
    layer8_outputs(4720) <= not (a xor b);
    layer8_outputs(4721) <= not a or b;
    layer8_outputs(4722) <= a;
    layer8_outputs(4723) <= b;
    layer8_outputs(4724) <= not (a and b);
    layer8_outputs(4725) <= a;
    layer8_outputs(4726) <= not a;
    layer8_outputs(4727) <= not (a or b);
    layer8_outputs(4728) <= not b;
    layer8_outputs(4729) <= b;
    layer8_outputs(4730) <= a or b;
    layer8_outputs(4731) <= a;
    layer8_outputs(4732) <= not b or a;
    layer8_outputs(4733) <= not (a xor b);
    layer8_outputs(4734) <= not (a or b);
    layer8_outputs(4735) <= a xor b;
    layer8_outputs(4736) <= not (a or b);
    layer8_outputs(4737) <= b;
    layer8_outputs(4738) <= not a;
    layer8_outputs(4739) <= not b;
    layer8_outputs(4740) <= not b;
    layer8_outputs(4741) <= a xor b;
    layer8_outputs(4742) <= not b;
    layer8_outputs(4743) <= not b;
    layer8_outputs(4744) <= a and not b;
    layer8_outputs(4745) <= not b;
    layer8_outputs(4746) <= b;
    layer8_outputs(4747) <= not (a and b);
    layer8_outputs(4748) <= not a;
    layer8_outputs(4749) <= not b or a;
    layer8_outputs(4750) <= not b;
    layer8_outputs(4751) <= not (a xor b);
    layer8_outputs(4752) <= b and not a;
    layer8_outputs(4753) <= not a;
    layer8_outputs(4754) <= not b;
    layer8_outputs(4755) <= a xor b;
    layer8_outputs(4756) <= not a;
    layer8_outputs(4757) <= a xor b;
    layer8_outputs(4758) <= not (a and b);
    layer8_outputs(4759) <= not a or b;
    layer8_outputs(4760) <= a;
    layer8_outputs(4761) <= not a;
    layer8_outputs(4762) <= a xor b;
    layer8_outputs(4763) <= a;
    layer8_outputs(4764) <= b and not a;
    layer8_outputs(4765) <= not a;
    layer8_outputs(4766) <= not (a or b);
    layer8_outputs(4767) <= b and not a;
    layer8_outputs(4768) <= not (a xor b);
    layer8_outputs(4769) <= not (a xor b);
    layer8_outputs(4770) <= a xor b;
    layer8_outputs(4771) <= b;
    layer8_outputs(4772) <= a;
    layer8_outputs(4773) <= a;
    layer8_outputs(4774) <= not (a and b);
    layer8_outputs(4775) <= not (a or b);
    layer8_outputs(4776) <= not b;
    layer8_outputs(4777) <= not b or a;
    layer8_outputs(4778) <= a or b;
    layer8_outputs(4779) <= not a;
    layer8_outputs(4780) <= not (a xor b);
    layer8_outputs(4781) <= b;
    layer8_outputs(4782) <= not (a xor b);
    layer8_outputs(4783) <= not b;
    layer8_outputs(4784) <= not b;
    layer8_outputs(4785) <= not (a or b);
    layer8_outputs(4786) <= not a;
    layer8_outputs(4787) <= not b;
    layer8_outputs(4788) <= not (a or b);
    layer8_outputs(4789) <= a or b;
    layer8_outputs(4790) <= b and not a;
    layer8_outputs(4791) <= a or b;
    layer8_outputs(4792) <= a and b;
    layer8_outputs(4793) <= a and b;
    layer8_outputs(4794) <= b;
    layer8_outputs(4795) <= b;
    layer8_outputs(4796) <= b;
    layer8_outputs(4797) <= a and not b;
    layer8_outputs(4798) <= not a or b;
    layer8_outputs(4799) <= b;
    layer8_outputs(4800) <= not b;
    layer8_outputs(4801) <= b;
    layer8_outputs(4802) <= '1';
    layer8_outputs(4803) <= a;
    layer8_outputs(4804) <= a xor b;
    layer8_outputs(4805) <= a;
    layer8_outputs(4806) <= a xor b;
    layer8_outputs(4807) <= a;
    layer8_outputs(4808) <= not a;
    layer8_outputs(4809) <= not b;
    layer8_outputs(4810) <= not a or b;
    layer8_outputs(4811) <= not (a or b);
    layer8_outputs(4812) <= not b;
    layer8_outputs(4813) <= a;
    layer8_outputs(4814) <= not b;
    layer8_outputs(4815) <= a or b;
    layer8_outputs(4816) <= a xor b;
    layer8_outputs(4817) <= not (a and b);
    layer8_outputs(4818) <= not a;
    layer8_outputs(4819) <= a xor b;
    layer8_outputs(4820) <= not a;
    layer8_outputs(4821) <= b;
    layer8_outputs(4822) <= not (a or b);
    layer8_outputs(4823) <= not b;
    layer8_outputs(4824) <= b;
    layer8_outputs(4825) <= not b;
    layer8_outputs(4826) <= a;
    layer8_outputs(4827) <= not (a xor b);
    layer8_outputs(4828) <= a;
    layer8_outputs(4829) <= a xor b;
    layer8_outputs(4830) <= b;
    layer8_outputs(4831) <= b;
    layer8_outputs(4832) <= a xor b;
    layer8_outputs(4833) <= not (a xor b);
    layer8_outputs(4834) <= a;
    layer8_outputs(4835) <= a;
    layer8_outputs(4836) <= not a;
    layer8_outputs(4837) <= not (a and b);
    layer8_outputs(4838) <= a and not b;
    layer8_outputs(4839) <= not b or a;
    layer8_outputs(4840) <= a and b;
    layer8_outputs(4841) <= a;
    layer8_outputs(4842) <= not b;
    layer8_outputs(4843) <= a;
    layer8_outputs(4844) <= a and not b;
    layer8_outputs(4845) <= not (a xor b);
    layer8_outputs(4846) <= a;
    layer8_outputs(4847) <= a xor b;
    layer8_outputs(4848) <= not a;
    layer8_outputs(4849) <= not b;
    layer8_outputs(4850) <= a;
    layer8_outputs(4851) <= not (a xor b);
    layer8_outputs(4852) <= a xor b;
    layer8_outputs(4853) <= b;
    layer8_outputs(4854) <= not (a xor b);
    layer8_outputs(4855) <= a xor b;
    layer8_outputs(4856) <= b;
    layer8_outputs(4857) <= not a;
    layer8_outputs(4858) <= a xor b;
    layer8_outputs(4859) <= b and not a;
    layer8_outputs(4860) <= b;
    layer8_outputs(4861) <= a or b;
    layer8_outputs(4862) <= a and not b;
    layer8_outputs(4863) <= not b;
    layer8_outputs(4864) <= b;
    layer8_outputs(4865) <= not (a or b);
    layer8_outputs(4866) <= not b;
    layer8_outputs(4867) <= b;
    layer8_outputs(4868) <= a and not b;
    layer8_outputs(4869) <= b;
    layer8_outputs(4870) <= not b;
    layer8_outputs(4871) <= a or b;
    layer8_outputs(4872) <= not a;
    layer8_outputs(4873) <= not (a and b);
    layer8_outputs(4874) <= a and not b;
    layer8_outputs(4875) <= b;
    layer8_outputs(4876) <= not a or b;
    layer8_outputs(4877) <= not a;
    layer8_outputs(4878) <= a and not b;
    layer8_outputs(4879) <= not b or a;
    layer8_outputs(4880) <= not (a and b);
    layer8_outputs(4881) <= b;
    layer8_outputs(4882) <= not a or b;
    layer8_outputs(4883) <= a;
    layer8_outputs(4884) <= a and b;
    layer8_outputs(4885) <= a xor b;
    layer8_outputs(4886) <= not b;
    layer8_outputs(4887) <= not (a xor b);
    layer8_outputs(4888) <= a;
    layer8_outputs(4889) <= a;
    layer8_outputs(4890) <= a;
    layer8_outputs(4891) <= not a;
    layer8_outputs(4892) <= not (a xor b);
    layer8_outputs(4893) <= not a;
    layer8_outputs(4894) <= a;
    layer8_outputs(4895) <= a and not b;
    layer8_outputs(4896) <= not (a and b);
    layer8_outputs(4897) <= a or b;
    layer8_outputs(4898) <= not b;
    layer8_outputs(4899) <= b and not a;
    layer8_outputs(4900) <= not b;
    layer8_outputs(4901) <= a;
    layer8_outputs(4902) <= a;
    layer8_outputs(4903) <= not a;
    layer8_outputs(4904) <= not (a xor b);
    layer8_outputs(4905) <= a xor b;
    layer8_outputs(4906) <= a or b;
    layer8_outputs(4907) <= not (a xor b);
    layer8_outputs(4908) <= not (a xor b);
    layer8_outputs(4909) <= a;
    layer8_outputs(4910) <= not b;
    layer8_outputs(4911) <= not (a or b);
    layer8_outputs(4912) <= not a;
    layer8_outputs(4913) <= not a or b;
    layer8_outputs(4914) <= not a or b;
    layer8_outputs(4915) <= b;
    layer8_outputs(4916) <= not (a and b);
    layer8_outputs(4917) <= not (a xor b);
    layer8_outputs(4918) <= a;
    layer8_outputs(4919) <= b;
    layer8_outputs(4920) <= a xor b;
    layer8_outputs(4921) <= b;
    layer8_outputs(4922) <= not b;
    layer8_outputs(4923) <= b;
    layer8_outputs(4924) <= a and b;
    layer8_outputs(4925) <= not b;
    layer8_outputs(4926) <= a xor b;
    layer8_outputs(4927) <= b;
    layer8_outputs(4928) <= b;
    layer8_outputs(4929) <= a or b;
    layer8_outputs(4930) <= not a;
    layer8_outputs(4931) <= '1';
    layer8_outputs(4932) <= a and b;
    layer8_outputs(4933) <= b;
    layer8_outputs(4934) <= a;
    layer8_outputs(4935) <= not (a and b);
    layer8_outputs(4936) <= a xor b;
    layer8_outputs(4937) <= not b;
    layer8_outputs(4938) <= not b;
    layer8_outputs(4939) <= not b;
    layer8_outputs(4940) <= a;
    layer8_outputs(4941) <= a xor b;
    layer8_outputs(4942) <= not a or b;
    layer8_outputs(4943) <= a and b;
    layer8_outputs(4944) <= a and b;
    layer8_outputs(4945) <= a;
    layer8_outputs(4946) <= a and b;
    layer8_outputs(4947) <= not a or b;
    layer8_outputs(4948) <= not a;
    layer8_outputs(4949) <= b;
    layer8_outputs(4950) <= a xor b;
    layer8_outputs(4951) <= a xor b;
    layer8_outputs(4952) <= a xor b;
    layer8_outputs(4953) <= a xor b;
    layer8_outputs(4954) <= a xor b;
    layer8_outputs(4955) <= not (a and b);
    layer8_outputs(4956) <= not (a xor b);
    layer8_outputs(4957) <= not (a and b);
    layer8_outputs(4958) <= a and not b;
    layer8_outputs(4959) <= a and not b;
    layer8_outputs(4960) <= a or b;
    layer8_outputs(4961) <= a;
    layer8_outputs(4962) <= a xor b;
    layer8_outputs(4963) <= a xor b;
    layer8_outputs(4964) <= not (a or b);
    layer8_outputs(4965) <= not a;
    layer8_outputs(4966) <= not (a and b);
    layer8_outputs(4967) <= not b;
    layer8_outputs(4968) <= b and not a;
    layer8_outputs(4969) <= a and not b;
    layer8_outputs(4970) <= not (a xor b);
    layer8_outputs(4971) <= a;
    layer8_outputs(4972) <= not (a or b);
    layer8_outputs(4973) <= not a or b;
    layer8_outputs(4974) <= not a;
    layer8_outputs(4975) <= b;
    layer8_outputs(4976) <= b;
    layer8_outputs(4977) <= not b;
    layer8_outputs(4978) <= b and not a;
    layer8_outputs(4979) <= not (a or b);
    layer8_outputs(4980) <= b;
    layer8_outputs(4981) <= not b;
    layer8_outputs(4982) <= not a;
    layer8_outputs(4983) <= not b;
    layer8_outputs(4984) <= a xor b;
    layer8_outputs(4985) <= not a or b;
    layer8_outputs(4986) <= not b or a;
    layer8_outputs(4987) <= not b or a;
    layer8_outputs(4988) <= not a;
    layer8_outputs(4989) <= a xor b;
    layer8_outputs(4990) <= not b;
    layer8_outputs(4991) <= a or b;
    layer8_outputs(4992) <= not (a or b);
    layer8_outputs(4993) <= not b;
    layer8_outputs(4994) <= not a;
    layer8_outputs(4995) <= a and not b;
    layer8_outputs(4996) <= not b or a;
    layer8_outputs(4997) <= not (a xor b);
    layer8_outputs(4998) <= not (a xor b);
    layer8_outputs(4999) <= not b;
    layer8_outputs(5000) <= b;
    layer8_outputs(5001) <= b and not a;
    layer8_outputs(5002) <= b and not a;
    layer8_outputs(5003) <= a or b;
    layer8_outputs(5004) <= not (a and b);
    layer8_outputs(5005) <= not a;
    layer8_outputs(5006) <= b;
    layer8_outputs(5007) <= a or b;
    layer8_outputs(5008) <= a and not b;
    layer8_outputs(5009) <= a or b;
    layer8_outputs(5010) <= not b;
    layer8_outputs(5011) <= not (a xor b);
    layer8_outputs(5012) <= a and not b;
    layer8_outputs(5013) <= not b or a;
    layer8_outputs(5014) <= not b or a;
    layer8_outputs(5015) <= not (a xor b);
    layer8_outputs(5016) <= a and b;
    layer8_outputs(5017) <= not a;
    layer8_outputs(5018) <= a or b;
    layer8_outputs(5019) <= a xor b;
    layer8_outputs(5020) <= not a;
    layer8_outputs(5021) <= b;
    layer8_outputs(5022) <= a;
    layer8_outputs(5023) <= not a;
    layer8_outputs(5024) <= a;
    layer8_outputs(5025) <= b;
    layer8_outputs(5026) <= b;
    layer8_outputs(5027) <= a xor b;
    layer8_outputs(5028) <= a and b;
    layer8_outputs(5029) <= not a or b;
    layer8_outputs(5030) <= a;
    layer8_outputs(5031) <= not b or a;
    layer8_outputs(5032) <= not b;
    layer8_outputs(5033) <= b;
    layer8_outputs(5034) <= not a;
    layer8_outputs(5035) <= a and not b;
    layer8_outputs(5036) <= a;
    layer8_outputs(5037) <= not (a or b);
    layer8_outputs(5038) <= not (a xor b);
    layer8_outputs(5039) <= a and not b;
    layer8_outputs(5040) <= not a;
    layer8_outputs(5041) <= a xor b;
    layer8_outputs(5042) <= not a or b;
    layer8_outputs(5043) <= not a;
    layer8_outputs(5044) <= not (a xor b);
    layer8_outputs(5045) <= a and b;
    layer8_outputs(5046) <= not a;
    layer8_outputs(5047) <= not (a xor b);
    layer8_outputs(5048) <= not (a xor b);
    layer8_outputs(5049) <= a xor b;
    layer8_outputs(5050) <= not (a xor b);
    layer8_outputs(5051) <= a xor b;
    layer8_outputs(5052) <= a and b;
    layer8_outputs(5053) <= a;
    layer8_outputs(5054) <= not (a xor b);
    layer8_outputs(5055) <= b;
    layer8_outputs(5056) <= not a;
    layer8_outputs(5057) <= not a;
    layer8_outputs(5058) <= a;
    layer8_outputs(5059) <= not b or a;
    layer8_outputs(5060) <= not b;
    layer8_outputs(5061) <= not (a xor b);
    layer8_outputs(5062) <= b;
    layer8_outputs(5063) <= not a or b;
    layer8_outputs(5064) <= not b;
    layer8_outputs(5065) <= a;
    layer8_outputs(5066) <= a and not b;
    layer8_outputs(5067) <= b;
    layer8_outputs(5068) <= b;
    layer8_outputs(5069) <= a;
    layer8_outputs(5070) <= not (a and b);
    layer8_outputs(5071) <= not (a xor b);
    layer8_outputs(5072) <= b and not a;
    layer8_outputs(5073) <= a and not b;
    layer8_outputs(5074) <= b;
    layer8_outputs(5075) <= a xor b;
    layer8_outputs(5076) <= b;
    layer8_outputs(5077) <= not a;
    layer8_outputs(5078) <= a or b;
    layer8_outputs(5079) <= a and b;
    layer8_outputs(5080) <= not (a and b);
    layer8_outputs(5081) <= a or b;
    layer8_outputs(5082) <= not (a xor b);
    layer8_outputs(5083) <= not b or a;
    layer8_outputs(5084) <= b and not a;
    layer8_outputs(5085) <= not (a and b);
    layer8_outputs(5086) <= not b;
    layer8_outputs(5087) <= not (a xor b);
    layer8_outputs(5088) <= not (a and b);
    layer8_outputs(5089) <= not (a xor b);
    layer8_outputs(5090) <= not (a xor b);
    layer8_outputs(5091) <= a and b;
    layer8_outputs(5092) <= b and not a;
    layer8_outputs(5093) <= not (a and b);
    layer8_outputs(5094) <= not b;
    layer8_outputs(5095) <= not b;
    layer8_outputs(5096) <= not b;
    layer8_outputs(5097) <= not b;
    layer8_outputs(5098) <= not (a and b);
    layer8_outputs(5099) <= not b;
    layer8_outputs(5100) <= not b;
    layer8_outputs(5101) <= not b or a;
    layer8_outputs(5102) <= b;
    layer8_outputs(5103) <= a and b;
    layer8_outputs(5104) <= a;
    layer8_outputs(5105) <= not (a or b);
    layer8_outputs(5106) <= not b;
    layer8_outputs(5107) <= not (a or b);
    layer8_outputs(5108) <= not a;
    layer8_outputs(5109) <= a and not b;
    layer8_outputs(5110) <= not (a xor b);
    layer8_outputs(5111) <= not a;
    layer8_outputs(5112) <= '0';
    layer8_outputs(5113) <= not b or a;
    layer8_outputs(5114) <= not b;
    layer8_outputs(5115) <= a xor b;
    layer8_outputs(5116) <= b;
    layer8_outputs(5117) <= a xor b;
    layer8_outputs(5118) <= b and not a;
    layer8_outputs(5119) <= a;
    outputs(0) <= a;
    outputs(1) <= a xor b;
    outputs(2) <= b and not a;
    outputs(3) <= a;
    outputs(4) <= not (a and b);
    outputs(5) <= not (a xor b);
    outputs(6) <= b;
    outputs(7) <= a;
    outputs(8) <= b;
    outputs(9) <= a;
    outputs(10) <= a;
    outputs(11) <= b;
    outputs(12) <= a and not b;
    outputs(13) <= not a;
    outputs(14) <= a and not b;
    outputs(15) <= a;
    outputs(16) <= not (a or b);
    outputs(17) <= not (a or b);
    outputs(18) <= not b;
    outputs(19) <= not a;
    outputs(20) <= a;
    outputs(21) <= not a;
    outputs(22) <= not (a and b);
    outputs(23) <= a xor b;
    outputs(24) <= not (a or b);
    outputs(25) <= b;
    outputs(26) <= not (a xor b);
    outputs(27) <= a and b;
    outputs(28) <= a;
    outputs(29) <= not b;
    outputs(30) <= not a;
    outputs(31) <= a xor b;
    outputs(32) <= a xor b;
    outputs(33) <= a;
    outputs(34) <= a xor b;
    outputs(35) <= not b;
    outputs(36) <= a;
    outputs(37) <= a;
    outputs(38) <= not (a xor b);
    outputs(39) <= b;
    outputs(40) <= not (a xor b);
    outputs(41) <= not a;
    outputs(42) <= not (a xor b);
    outputs(43) <= not b or a;
    outputs(44) <= not (a xor b);
    outputs(45) <= b;
    outputs(46) <= not b;
    outputs(47) <= b and not a;
    outputs(48) <= a;
    outputs(49) <= a;
    outputs(50) <= not a;
    outputs(51) <= not b;
    outputs(52) <= not a;
    outputs(53) <= not a;
    outputs(54) <= not a;
    outputs(55) <= not (a or b);
    outputs(56) <= a xor b;
    outputs(57) <= a;
    outputs(58) <= not a;
    outputs(59) <= a;
    outputs(60) <= a and not b;
    outputs(61) <= a and b;
    outputs(62) <= a;
    outputs(63) <= not (a or b);
    outputs(64) <= not (a xor b);
    outputs(65) <= b;
    outputs(66) <= a;
    outputs(67) <= not a;
    outputs(68) <= not b;
    outputs(69) <= a and not b;
    outputs(70) <= a and b;
    outputs(71) <= not a;
    outputs(72) <= a and not b;
    outputs(73) <= not a;
    outputs(74) <= not b or a;
    outputs(75) <= a;
    outputs(76) <= b;
    outputs(77) <= not b;
    outputs(78) <= not b;
    outputs(79) <= a xor b;
    outputs(80) <= a and not b;
    outputs(81) <= not b;
    outputs(82) <= b and not a;
    outputs(83) <= not (a or b);
    outputs(84) <= not b;
    outputs(85) <= not a;
    outputs(86) <= a and not b;
    outputs(87) <= a xor b;
    outputs(88) <= not (a xor b);
    outputs(89) <= not a;
    outputs(90) <= b;
    outputs(91) <= not b;
    outputs(92) <= a and not b;
    outputs(93) <= b;
    outputs(94) <= a;
    outputs(95) <= a or b;
    outputs(96) <= not b;
    outputs(97) <= b and not a;
    outputs(98) <= not (a xor b);
    outputs(99) <= not a;
    outputs(100) <= not b;
    outputs(101) <= b;
    outputs(102) <= not a;
    outputs(103) <= a and not b;
    outputs(104) <= b;
    outputs(105) <= not b;
    outputs(106) <= b;
    outputs(107) <= a and not b;
    outputs(108) <= a and b;
    outputs(109) <= not b;
    outputs(110) <= b;
    outputs(111) <= a;
    outputs(112) <= b and not a;
    outputs(113) <= not (a or b);
    outputs(114) <= not a;
    outputs(115) <= a and not b;
    outputs(116) <= a xor b;
    outputs(117) <= not b;
    outputs(118) <= a and b;
    outputs(119) <= not (a xor b);
    outputs(120) <= not b;
    outputs(121) <= a and not b;
    outputs(122) <= a;
    outputs(123) <= not a;
    outputs(124) <= not a;
    outputs(125) <= b;
    outputs(126) <= not a;
    outputs(127) <= not b;
    outputs(128) <= b and not a;
    outputs(129) <= a xor b;
    outputs(130) <= not b;
    outputs(131) <= b and not a;
    outputs(132) <= a and not b;
    outputs(133) <= b;
    outputs(134) <= not (a xor b);
    outputs(135) <= not (a xor b);
    outputs(136) <= a or b;
    outputs(137) <= a;
    outputs(138) <= not (a or b);
    outputs(139) <= a and not b;
    outputs(140) <= not a;
    outputs(141) <= not (a xor b);
    outputs(142) <= a xor b;
    outputs(143) <= b;
    outputs(144) <= a;
    outputs(145) <= b;
    outputs(146) <= not (a xor b);
    outputs(147) <= not a;
    outputs(148) <= not (a xor b);
    outputs(149) <= a xor b;
    outputs(150) <= a and b;
    outputs(151) <= a and b;
    outputs(152) <= not b;
    outputs(153) <= not b;
    outputs(154) <= not a;
    outputs(155) <= a;
    outputs(156) <= b;
    outputs(157) <= b;
    outputs(158) <= not b;
    outputs(159) <= not (a xor b);
    outputs(160) <= a and not b;
    outputs(161) <= not b or a;
    outputs(162) <= not a;
    outputs(163) <= b;
    outputs(164) <= not b;
    outputs(165) <= not a;
    outputs(166) <= b;
    outputs(167) <= not a;
    outputs(168) <= a xor b;
    outputs(169) <= not (a xor b);
    outputs(170) <= not b;
    outputs(171) <= b;
    outputs(172) <= not a;
    outputs(173) <= not b;
    outputs(174) <= a xor b;
    outputs(175) <= a and b;
    outputs(176) <= not (a and b);
    outputs(177) <= a or b;
    outputs(178) <= a xor b;
    outputs(179) <= b;
    outputs(180) <= b;
    outputs(181) <= not a;
    outputs(182) <= not a;
    outputs(183) <= not a;
    outputs(184) <= not b;
    outputs(185) <= a and b;
    outputs(186) <= a and not b;
    outputs(187) <= b and not a;
    outputs(188) <= not a;
    outputs(189) <= a or b;
    outputs(190) <= not a;
    outputs(191) <= a;
    outputs(192) <= not a;
    outputs(193) <= b;
    outputs(194) <= a and b;
    outputs(195) <= a;
    outputs(196) <= b;
    outputs(197) <= not (a or b);
    outputs(198) <= b;
    outputs(199) <= b;
    outputs(200) <= a xor b;
    outputs(201) <= not a or b;
    outputs(202) <= a;
    outputs(203) <= a and not b;
    outputs(204) <= not (a or b);
    outputs(205) <= not (a xor b);
    outputs(206) <= a or b;
    outputs(207) <= not b or a;
    outputs(208) <= a and b;
    outputs(209) <= not (a xor b);
    outputs(210) <= not a;
    outputs(211) <= a and not b;
    outputs(212) <= not (a xor b);
    outputs(213) <= b and not a;
    outputs(214) <= not (a xor b);
    outputs(215) <= not a;
    outputs(216) <= not a;
    outputs(217) <= not b or a;
    outputs(218) <= not a;
    outputs(219) <= a;
    outputs(220) <= not a;
    outputs(221) <= a and not b;
    outputs(222) <= a or b;
    outputs(223) <= b;
    outputs(224) <= a;
    outputs(225) <= not b;
    outputs(226) <= a;
    outputs(227) <= not a;
    outputs(228) <= a;
    outputs(229) <= not (a or b);
    outputs(230) <= not b;
    outputs(231) <= not b;
    outputs(232) <= not a;
    outputs(233) <= b and not a;
    outputs(234) <= not a;
    outputs(235) <= not a;
    outputs(236) <= not b;
    outputs(237) <= a;
    outputs(238) <= b;
    outputs(239) <= not (a and b);
    outputs(240) <= not b;
    outputs(241) <= not (a and b);
    outputs(242) <= not a;
    outputs(243) <= not (a or b);
    outputs(244) <= not a;
    outputs(245) <= not a;
    outputs(246) <= a and b;
    outputs(247) <= not b;
    outputs(248) <= a and b;
    outputs(249) <= a and not b;
    outputs(250) <= a and not b;
    outputs(251) <= b and not a;
    outputs(252) <= a xor b;
    outputs(253) <= a xor b;
    outputs(254) <= not (a xor b);
    outputs(255) <= a xor b;
    outputs(256) <= not b or a;
    outputs(257) <= a;
    outputs(258) <= not (a xor b);
    outputs(259) <= not (a xor b);
    outputs(260) <= not a;
    outputs(261) <= not (a xor b);
    outputs(262) <= not (a xor b);
    outputs(263) <= not b;
    outputs(264) <= a;
    outputs(265) <= not a;
    outputs(266) <= a or b;
    outputs(267) <= b and not a;
    outputs(268) <= a and not b;
    outputs(269) <= b;
    outputs(270) <= not b;
    outputs(271) <= b;
    outputs(272) <= a;
    outputs(273) <= b;
    outputs(274) <= a;
    outputs(275) <= a;
    outputs(276) <= a xor b;
    outputs(277) <= not (a or b);
    outputs(278) <= a;
    outputs(279) <= not b;
    outputs(280) <= not (a xor b);
    outputs(281) <= b;
    outputs(282) <= b;
    outputs(283) <= not (a xor b);
    outputs(284) <= not b;
    outputs(285) <= a;
    outputs(286) <= b;
    outputs(287) <= a and not b;
    outputs(288) <= not (a or b);
    outputs(289) <= a xor b;
    outputs(290) <= not b;
    outputs(291) <= not a;
    outputs(292) <= not b;
    outputs(293) <= a and not b;
    outputs(294) <= not b;
    outputs(295) <= not (a or b);
    outputs(296) <= not b;
    outputs(297) <= a xor b;
    outputs(298) <= a;
    outputs(299) <= not (a xor b);
    outputs(300) <= a;
    outputs(301) <= a;
    outputs(302) <= not b;
    outputs(303) <= a and b;
    outputs(304) <= not b;
    outputs(305) <= a;
    outputs(306) <= not b;
    outputs(307) <= not (a and b);
    outputs(308) <= not a;
    outputs(309) <= a or b;
    outputs(310) <= not (a xor b);
    outputs(311) <= b;
    outputs(312) <= a and b;
    outputs(313) <= a and b;
    outputs(314) <= a xor b;
    outputs(315) <= a and b;
    outputs(316) <= not b;
    outputs(317) <= a;
    outputs(318) <= not a;
    outputs(319) <= a;
    outputs(320) <= not (a xor b);
    outputs(321) <= a and not b;
    outputs(322) <= b;
    outputs(323) <= a;
    outputs(324) <= not a;
    outputs(325) <= not b;
    outputs(326) <= a and not b;
    outputs(327) <= not (a or b);
    outputs(328) <= a and not b;
    outputs(329) <= b;
    outputs(330) <= not (a and b);
    outputs(331) <= not b;
    outputs(332) <= not a;
    outputs(333) <= b;
    outputs(334) <= not b;
    outputs(335) <= not a;
    outputs(336) <= a and not b;
    outputs(337) <= not a;
    outputs(338) <= not (a and b);
    outputs(339) <= a xor b;
    outputs(340) <= a and not b;
    outputs(341) <= not b;
    outputs(342) <= a and b;
    outputs(343) <= b;
    outputs(344) <= not (a xor b);
    outputs(345) <= a xor b;
    outputs(346) <= b;
    outputs(347) <= a;
    outputs(348) <= a and b;
    outputs(349) <= b;
    outputs(350) <= not a;
    outputs(351) <= a xor b;
    outputs(352) <= b;
    outputs(353) <= b and not a;
    outputs(354) <= not a;
    outputs(355) <= a and not b;
    outputs(356) <= not (a or b);
    outputs(357) <= a xor b;
    outputs(358) <= a;
    outputs(359) <= a xor b;
    outputs(360) <= not (a xor b);
    outputs(361) <= a and not b;
    outputs(362) <= b and not a;
    outputs(363) <= a and b;
    outputs(364) <= not a or b;
    outputs(365) <= not a;
    outputs(366) <= not b;
    outputs(367) <= not (a xor b);
    outputs(368) <= not b;
    outputs(369) <= b;
    outputs(370) <= a;
    outputs(371) <= b and not a;
    outputs(372) <= a and not b;
    outputs(373) <= a;
    outputs(374) <= not b;
    outputs(375) <= not (a or b);
    outputs(376) <= a xor b;
    outputs(377) <= a xor b;
    outputs(378) <= not (a or b);
    outputs(379) <= a;
    outputs(380) <= a and b;
    outputs(381) <= not a;
    outputs(382) <= b;
    outputs(383) <= not (a or b);
    outputs(384) <= not (a and b);
    outputs(385) <= a and b;
    outputs(386) <= not b;
    outputs(387) <= b;
    outputs(388) <= b;
    outputs(389) <= a xor b;
    outputs(390) <= not a;
    outputs(391) <= not b;
    outputs(392) <= not (a xor b);
    outputs(393) <= a;
    outputs(394) <= b;
    outputs(395) <= not (a xor b);
    outputs(396) <= not a;
    outputs(397) <= not b;
    outputs(398) <= a;
    outputs(399) <= not a;
    outputs(400) <= a and not b;
    outputs(401) <= not a;
    outputs(402) <= a xor b;
    outputs(403) <= a;
    outputs(404) <= a;
    outputs(405) <= a and not b;
    outputs(406) <= a xor b;
    outputs(407) <= b;
    outputs(408) <= a;
    outputs(409) <= a;
    outputs(410) <= b and not a;
    outputs(411) <= not (a xor b);
    outputs(412) <= a and not b;
    outputs(413) <= b;
    outputs(414) <= a and not b;
    outputs(415) <= a xor b;
    outputs(416) <= not (a xor b);
    outputs(417) <= not a or b;
    outputs(418) <= not (a and b);
    outputs(419) <= not (a or b);
    outputs(420) <= not (a xor b);
    outputs(421) <= a;
    outputs(422) <= a xor b;
    outputs(423) <= not (a and b);
    outputs(424) <= not a or b;
    outputs(425) <= not a;
    outputs(426) <= b and not a;
    outputs(427) <= a and b;
    outputs(428) <= a and b;
    outputs(429) <= a xor b;
    outputs(430) <= a;
    outputs(431) <= not (a and b);
    outputs(432) <= a;
    outputs(433) <= a and not b;
    outputs(434) <= a and not b;
    outputs(435) <= a xor b;
    outputs(436) <= not a;
    outputs(437) <= not (a xor b);
    outputs(438) <= not (a xor b);
    outputs(439) <= a xor b;
    outputs(440) <= not a;
    outputs(441) <= not a;
    outputs(442) <= not a;
    outputs(443) <= b;
    outputs(444) <= b;
    outputs(445) <= b;
    outputs(446) <= a;
    outputs(447) <= a and not b;
    outputs(448) <= not (a and b);
    outputs(449) <= not b;
    outputs(450) <= not (a or b);
    outputs(451) <= not a;
    outputs(452) <= not b;
    outputs(453) <= not a;
    outputs(454) <= a;
    outputs(455) <= not b;
    outputs(456) <= not (a xor b);
    outputs(457) <= not (a or b);
    outputs(458) <= not a;
    outputs(459) <= b and not a;
    outputs(460) <= b;
    outputs(461) <= not b;
    outputs(462) <= a xor b;
    outputs(463) <= not b or a;
    outputs(464) <= b;
    outputs(465) <= not a;
    outputs(466) <= not (a or b);
    outputs(467) <= not (a or b);
    outputs(468) <= b and not a;
    outputs(469) <= b;
    outputs(470) <= not (a xor b);
    outputs(471) <= a xor b;
    outputs(472) <= a xor b;
    outputs(473) <= not a;
    outputs(474) <= not b or a;
    outputs(475) <= not a;
    outputs(476) <= a;
    outputs(477) <= a and b;
    outputs(478) <= b and not a;
    outputs(479) <= a;
    outputs(480) <= not b or a;
    outputs(481) <= a;
    outputs(482) <= not a;
    outputs(483) <= a xor b;
    outputs(484) <= a xor b;
    outputs(485) <= b;
    outputs(486) <= not b;
    outputs(487) <= a and b;
    outputs(488) <= not b;
    outputs(489) <= not a;
    outputs(490) <= not (a xor b);
    outputs(491) <= not (a and b);
    outputs(492) <= b;
    outputs(493) <= not (a xor b);
    outputs(494) <= a and b;
    outputs(495) <= a;
    outputs(496) <= not b;
    outputs(497) <= b;
    outputs(498) <= b;
    outputs(499) <= not b;
    outputs(500) <= b and not a;
    outputs(501) <= b;
    outputs(502) <= a xor b;
    outputs(503) <= a and b;
    outputs(504) <= not (a xor b);
    outputs(505) <= b;
    outputs(506) <= not a;
    outputs(507) <= not b;
    outputs(508) <= b;
    outputs(509) <= b;
    outputs(510) <= b and not a;
    outputs(511) <= a xor b;
    outputs(512) <= not (a xor b);
    outputs(513) <= a;
    outputs(514) <= b and not a;
    outputs(515) <= b;
    outputs(516) <= not b;
    outputs(517) <= b;
    outputs(518) <= not (a and b);
    outputs(519) <= not b;
    outputs(520) <= not (a or b);
    outputs(521) <= not a;
    outputs(522) <= b;
    outputs(523) <= a and not b;
    outputs(524) <= a and not b;
    outputs(525) <= not b;
    outputs(526) <= not a;
    outputs(527) <= not b;
    outputs(528) <= a xor b;
    outputs(529) <= not (a xor b);
    outputs(530) <= not (a or b);
    outputs(531) <= not b;
    outputs(532) <= not b;
    outputs(533) <= a and not b;
    outputs(534) <= a;
    outputs(535) <= not (a xor b);
    outputs(536) <= a and not b;
    outputs(537) <= not a;
    outputs(538) <= not (a or b);
    outputs(539) <= b;
    outputs(540) <= a;
    outputs(541) <= a and b;
    outputs(542) <= a xor b;
    outputs(543) <= not b;
    outputs(544) <= b and not a;
    outputs(545) <= not (a or b);
    outputs(546) <= a and not b;
    outputs(547) <= a xor b;
    outputs(548) <= not a;
    outputs(549) <= '0';
    outputs(550) <= not a;
    outputs(551) <= not a;
    outputs(552) <= a xor b;
    outputs(553) <= a and b;
    outputs(554) <= not (a xor b);
    outputs(555) <= a;
    outputs(556) <= a xor b;
    outputs(557) <= not (a or b);
    outputs(558) <= not (a or b);
    outputs(559) <= b and not a;
    outputs(560) <= a xor b;
    outputs(561) <= not (a or b);
    outputs(562) <= b;
    outputs(563) <= b and not a;
    outputs(564) <= a and b;
    outputs(565) <= b;
    outputs(566) <= b and not a;
    outputs(567) <= not (a or b);
    outputs(568) <= not (a xor b);
    outputs(569) <= a xor b;
    outputs(570) <= a xor b;
    outputs(571) <= a;
    outputs(572) <= not b;
    outputs(573) <= not (a and b);
    outputs(574) <= a xor b;
    outputs(575) <= not b;
    outputs(576) <= b;
    outputs(577) <= b;
    outputs(578) <= not a;
    outputs(579) <= not a;
    outputs(580) <= a and b;
    outputs(581) <= a;
    outputs(582) <= not a;
    outputs(583) <= b;
    outputs(584) <= not b;
    outputs(585) <= not a;
    outputs(586) <= not a;
    outputs(587) <= a xor b;
    outputs(588) <= a xor b;
    outputs(589) <= b;
    outputs(590) <= not (a or b);
    outputs(591) <= b;
    outputs(592) <= a;
    outputs(593) <= not b;
    outputs(594) <= a xor b;
    outputs(595) <= not a;
    outputs(596) <= b and not a;
    outputs(597) <= b;
    outputs(598) <= not (a xor b);
    outputs(599) <= a or b;
    outputs(600) <= a and b;
    outputs(601) <= not a;
    outputs(602) <= a;
    outputs(603) <= b;
    outputs(604) <= not (a or b);
    outputs(605) <= b;
    outputs(606) <= a and b;
    outputs(607) <= not a or b;
    outputs(608) <= not b;
    outputs(609) <= not b;
    outputs(610) <= not (a xor b);
    outputs(611) <= a xor b;
    outputs(612) <= not (a or b);
    outputs(613) <= a and not b;
    outputs(614) <= a;
    outputs(615) <= a xor b;
    outputs(616) <= a and b;
    outputs(617) <= a xor b;
    outputs(618) <= b;
    outputs(619) <= not a;
    outputs(620) <= not b;
    outputs(621) <= not (a xor b);
    outputs(622) <= a and b;
    outputs(623) <= b;
    outputs(624) <= a and b;
    outputs(625) <= b;
    outputs(626) <= not (a or b);
    outputs(627) <= not a;
    outputs(628) <= a;
    outputs(629) <= not (a and b);
    outputs(630) <= a and b;
    outputs(631) <= b and not a;
    outputs(632) <= b;
    outputs(633) <= not (a xor b);
    outputs(634) <= b and not a;
    outputs(635) <= not a;
    outputs(636) <= not (a or b);
    outputs(637) <= b and not a;
    outputs(638) <= a and b;
    outputs(639) <= not b;
    outputs(640) <= b;
    outputs(641) <= b and not a;
    outputs(642) <= b and not a;
    outputs(643) <= not a;
    outputs(644) <= not (a xor b);
    outputs(645) <= a;
    outputs(646) <= b and not a;
    outputs(647) <= b and not a;
    outputs(648) <= not b;
    outputs(649) <= a xor b;
    outputs(650) <= a;
    outputs(651) <= not (a xor b);
    outputs(652) <= not a;
    outputs(653) <= not (a xor b);
    outputs(654) <= a xor b;
    outputs(655) <= a;
    outputs(656) <= a and not b;
    outputs(657) <= a xor b;
    outputs(658) <= a and not b;
    outputs(659) <= a xor b;
    outputs(660) <= a and not b;
    outputs(661) <= a xor b;
    outputs(662) <= not (a xor b);
    outputs(663) <= a xor b;
    outputs(664) <= not (a xor b);
    outputs(665) <= not b or a;
    outputs(666) <= not b;
    outputs(667) <= a xor b;
    outputs(668) <= not (a xor b);
    outputs(669) <= a and not b;
    outputs(670) <= b;
    outputs(671) <= a and not b;
    outputs(672) <= a and not b;
    outputs(673) <= b and not a;
    outputs(674) <= a and b;
    outputs(675) <= a;
    outputs(676) <= b;
    outputs(677) <= b and not a;
    outputs(678) <= not a;
    outputs(679) <= not (a xor b);
    outputs(680) <= a;
    outputs(681) <= b and not a;
    outputs(682) <= b;
    outputs(683) <= not a;
    outputs(684) <= not (a and b);
    outputs(685) <= b and not a;
    outputs(686) <= not b or a;
    outputs(687) <= not a;
    outputs(688) <= not b;
    outputs(689) <= a and b;
    outputs(690) <= not (a xor b);
    outputs(691) <= not b;
    outputs(692) <= a xor b;
    outputs(693) <= not a;
    outputs(694) <= not b;
    outputs(695) <= not (a xor b);
    outputs(696) <= a;
    outputs(697) <= b and not a;
    outputs(698) <= a;
    outputs(699) <= not b;
    outputs(700) <= a and not b;
    outputs(701) <= b and not a;
    outputs(702) <= not (a or b);
    outputs(703) <= a and b;
    outputs(704) <= not b;
    outputs(705) <= a and not b;
    outputs(706) <= a and not b;
    outputs(707) <= a and b;
    outputs(708) <= b;
    outputs(709) <= not (a xor b);
    outputs(710) <= a xor b;
    outputs(711) <= a and not b;
    outputs(712) <= a;
    outputs(713) <= b;
    outputs(714) <= not (a or b);
    outputs(715) <= not b or a;
    outputs(716) <= not (a or b);
    outputs(717) <= not (a or b);
    outputs(718) <= a xor b;
    outputs(719) <= not a;
    outputs(720) <= not (a xor b);
    outputs(721) <= a and b;
    outputs(722) <= a xor b;
    outputs(723) <= b;
    outputs(724) <= not b;
    outputs(725) <= not (a and b);
    outputs(726) <= a or b;
    outputs(727) <= a and b;
    outputs(728) <= a xor b;
    outputs(729) <= b;
    outputs(730) <= a and b;
    outputs(731) <= not b;
    outputs(732) <= a and b;
    outputs(733) <= a and b;
    outputs(734) <= a and b;
    outputs(735) <= a or b;
    outputs(736) <= b;
    outputs(737) <= a;
    outputs(738) <= not (a or b);
    outputs(739) <= a and b;
    outputs(740) <= not (a xor b);
    outputs(741) <= b;
    outputs(742) <= b and not a;
    outputs(743) <= a xor b;
    outputs(744) <= a and not b;
    outputs(745) <= not (a xor b);
    outputs(746) <= not (a or b);
    outputs(747) <= a and not b;
    outputs(748) <= not (a xor b);
    outputs(749) <= not a;
    outputs(750) <= not (a or b);
    outputs(751) <= a and not b;
    outputs(752) <= not b;
    outputs(753) <= a;
    outputs(754) <= b and not a;
    outputs(755) <= not (a or b);
    outputs(756) <= not b;
    outputs(757) <= not a;
    outputs(758) <= a xor b;
    outputs(759) <= a and b;
    outputs(760) <= a and b;
    outputs(761) <= a and not b;
    outputs(762) <= a and b;
    outputs(763) <= b and not a;
    outputs(764) <= a xor b;
    outputs(765) <= b and not a;
    outputs(766) <= a and b;
    outputs(767) <= not (a or b);
    outputs(768) <= b;
    outputs(769) <= not (a xor b);
    outputs(770) <= a and not b;
    outputs(771) <= not a;
    outputs(772) <= a and not b;
    outputs(773) <= not (a xor b);
    outputs(774) <= not b;
    outputs(775) <= not a;
    outputs(776) <= not a;
    outputs(777) <= a and not b;
    outputs(778) <= a xor b;
    outputs(779) <= not a;
    outputs(780) <= not (a and b);
    outputs(781) <= not a;
    outputs(782) <= not (a xor b);
    outputs(783) <= a xor b;
    outputs(784) <= a or b;
    outputs(785) <= a and not b;
    outputs(786) <= not b;
    outputs(787) <= b;
    outputs(788) <= a;
    outputs(789) <= not b;
    outputs(790) <= not (a xor b);
    outputs(791) <= a;
    outputs(792) <= not a;
    outputs(793) <= '0';
    outputs(794) <= b;
    outputs(795) <= a and not b;
    outputs(796) <= not (a xor b);
    outputs(797) <= not (a or b);
    outputs(798) <= a and b;
    outputs(799) <= a xor b;
    outputs(800) <= b;
    outputs(801) <= not (a xor b);
    outputs(802) <= not b;
    outputs(803) <= not (a xor b);
    outputs(804) <= not (a xor b);
    outputs(805) <= a and b;
    outputs(806) <= not b;
    outputs(807) <= b and not a;
    outputs(808) <= not (a xor b);
    outputs(809) <= b and not a;
    outputs(810) <= a;
    outputs(811) <= not b;
    outputs(812) <= not a;
    outputs(813) <= a xor b;
    outputs(814) <= not a;
    outputs(815) <= not (a or b);
    outputs(816) <= a;
    outputs(817) <= a and not b;
    outputs(818) <= not (a xor b);
    outputs(819) <= a and not b;
    outputs(820) <= b;
    outputs(821) <= not b;
    outputs(822) <= a and b;
    outputs(823) <= not a or b;
    outputs(824) <= b and not a;
    outputs(825) <= not a;
    outputs(826) <= b;
    outputs(827) <= not (a or b);
    outputs(828) <= not (a or b);
    outputs(829) <= not b;
    outputs(830) <= not a;
    outputs(831) <= a xor b;
    outputs(832) <= b and not a;
    outputs(833) <= a;
    outputs(834) <= not (a xor b);
    outputs(835) <= not a;
    outputs(836) <= a and not b;
    outputs(837) <= not (a or b);
    outputs(838) <= b;
    outputs(839) <= b;
    outputs(840) <= a and b;
    outputs(841) <= a or b;
    outputs(842) <= a xor b;
    outputs(843) <= a and b;
    outputs(844) <= b;
    outputs(845) <= b and not a;
    outputs(846) <= a and b;
    outputs(847) <= '0';
    outputs(848) <= a;
    outputs(849) <= b;
    outputs(850) <= not (a xor b);
    outputs(851) <= not (a or b);
    outputs(852) <= a xor b;
    outputs(853) <= not (a xor b);
    outputs(854) <= not b;
    outputs(855) <= a;
    outputs(856) <= a and b;
    outputs(857) <= a;
    outputs(858) <= b;
    outputs(859) <= not b;
    outputs(860) <= '0';
    outputs(861) <= not (a or b);
    outputs(862) <= a;
    outputs(863) <= not a;
    outputs(864) <= a;
    outputs(865) <= b;
    outputs(866) <= not (a xor b);
    outputs(867) <= a;
    outputs(868) <= a and not b;
    outputs(869) <= b;
    outputs(870) <= not (a or b);
    outputs(871) <= a and not b;
    outputs(872) <= not (a xor b);
    outputs(873) <= not b;
    outputs(874) <= not (a xor b);
    outputs(875) <= not (a or b);
    outputs(876) <= not (a or b);
    outputs(877) <= b and not a;
    outputs(878) <= not b;
    outputs(879) <= not a;
    outputs(880) <= a and not b;
    outputs(881) <= not b;
    outputs(882) <= a and not b;
    outputs(883) <= not (a xor b);
    outputs(884) <= a;
    outputs(885) <= a and b;
    outputs(886) <= a and not b;
    outputs(887) <= not b or a;
    outputs(888) <= '0';
    outputs(889) <= a xor b;
    outputs(890) <= not (a xor b);
    outputs(891) <= b and not a;
    outputs(892) <= a and b;
    outputs(893) <= not (a xor b);
    outputs(894) <= a and b;
    outputs(895) <= not a;
    outputs(896) <= not (a xor b);
    outputs(897) <= not (a xor b);
    outputs(898) <= not (a and b);
    outputs(899) <= a xor b;
    outputs(900) <= a;
    outputs(901) <= a xor b;
    outputs(902) <= a xor b;
    outputs(903) <= a and not b;
    outputs(904) <= a and not b;
    outputs(905) <= not b;
    outputs(906) <= a xor b;
    outputs(907) <= not (a xor b);
    outputs(908) <= not (a xor b);
    outputs(909) <= not (a xor b);
    outputs(910) <= b;
    outputs(911) <= not (a xor b);
    outputs(912) <= not a;
    outputs(913) <= not b;
    outputs(914) <= a;
    outputs(915) <= a and not b;
    outputs(916) <= not (a xor b);
    outputs(917) <= not b;
    outputs(918) <= b and not a;
    outputs(919) <= b;
    outputs(920) <= not b;
    outputs(921) <= a xor b;
    outputs(922) <= a;
    outputs(923) <= not b;
    outputs(924) <= a and b;
    outputs(925) <= a;
    outputs(926) <= a and not b;
    outputs(927) <= a and b;
    outputs(928) <= b;
    outputs(929) <= a and not b;
    outputs(930) <= a xor b;
    outputs(931) <= a;
    outputs(932) <= a and not b;
    outputs(933) <= not (a xor b);
    outputs(934) <= a;
    outputs(935) <= a xor b;
    outputs(936) <= not (a or b);
    outputs(937) <= a and b;
    outputs(938) <= b and not a;
    outputs(939) <= a xor b;
    outputs(940) <= not (a xor b);
    outputs(941) <= a xor b;
    outputs(942) <= a xor b;
    outputs(943) <= not a;
    outputs(944) <= a or b;
    outputs(945) <= a;
    outputs(946) <= a;
    outputs(947) <= b;
    outputs(948) <= not (a xor b);
    outputs(949) <= a xor b;
    outputs(950) <= a;
    outputs(951) <= a and not b;
    outputs(952) <= not (a or b);
    outputs(953) <= a;
    outputs(954) <= a and not b;
    outputs(955) <= not (a or b);
    outputs(956) <= not b;
    outputs(957) <= b and not a;
    outputs(958) <= a;
    outputs(959) <= not a;
    outputs(960) <= not a;
    outputs(961) <= a;
    outputs(962) <= not (a or b);
    outputs(963) <= a and not b;
    outputs(964) <= not (a xor b);
    outputs(965) <= a and not b;
    outputs(966) <= not (a xor b);
    outputs(967) <= not (a xor b);
    outputs(968) <= a and b;
    outputs(969) <= not (a or b);
    outputs(970) <= not b;
    outputs(971) <= not (a xor b);
    outputs(972) <= a;
    outputs(973) <= not b;
    outputs(974) <= a and b;
    outputs(975) <= not a;
    outputs(976) <= a xor b;
    outputs(977) <= b and not a;
    outputs(978) <= a and not b;
    outputs(979) <= not (a xor b);
    outputs(980) <= a and b;
    outputs(981) <= not (a or b);
    outputs(982) <= not b;
    outputs(983) <= not b;
    outputs(984) <= a or b;
    outputs(985) <= not a;
    outputs(986) <= b;
    outputs(987) <= a and not b;
    outputs(988) <= not a;
    outputs(989) <= a and b;
    outputs(990) <= a and not b;
    outputs(991) <= not b;
    outputs(992) <= a xor b;
    outputs(993) <= a;
    outputs(994) <= not b;
    outputs(995) <= not (a xor b);
    outputs(996) <= not a;
    outputs(997) <= not b;
    outputs(998) <= not b;
    outputs(999) <= b;
    outputs(1000) <= b;
    outputs(1001) <= a and not b;
    outputs(1002) <= not a;
    outputs(1003) <= a xor b;
    outputs(1004) <= a and not b;
    outputs(1005) <= a xor b;
    outputs(1006) <= b and not a;
    outputs(1007) <= '0';
    outputs(1008) <= not a;
    outputs(1009) <= a xor b;
    outputs(1010) <= b;
    outputs(1011) <= not b;
    outputs(1012) <= a xor b;
    outputs(1013) <= a;
    outputs(1014) <= b and not a;
    outputs(1015) <= not a;
    outputs(1016) <= not (a xor b);
    outputs(1017) <= a and not b;
    outputs(1018) <= not a;
    outputs(1019) <= a and b;
    outputs(1020) <= not (a xor b);
    outputs(1021) <= not (a xor b);
    outputs(1022) <= not b;
    outputs(1023) <= a xor b;
    outputs(1024) <= not (a xor b);
    outputs(1025) <= b;
    outputs(1026) <= b;
    outputs(1027) <= not a or b;
    outputs(1028) <= not b;
    outputs(1029) <= not b;
    outputs(1030) <= not (a xor b);
    outputs(1031) <= not a or b;
    outputs(1032) <= b and not a;
    outputs(1033) <= not (a xor b);
    outputs(1034) <= not b or a;
    outputs(1035) <= a xor b;
    outputs(1036) <= not b;
    outputs(1037) <= a;
    outputs(1038) <= not a;
    outputs(1039) <= a and b;
    outputs(1040) <= a and b;
    outputs(1041) <= b;
    outputs(1042) <= b;
    outputs(1043) <= b;
    outputs(1044) <= a;
    outputs(1045) <= b;
    outputs(1046) <= b;
    outputs(1047) <= not b;
    outputs(1048) <= a xor b;
    outputs(1049) <= not b;
    outputs(1050) <= a and b;
    outputs(1051) <= b and not a;
    outputs(1052) <= not (a xor b);
    outputs(1053) <= not (a and b);
    outputs(1054) <= not (a xor b);
    outputs(1055) <= not a;
    outputs(1056) <= not a;
    outputs(1057) <= b;
    outputs(1058) <= b;
    outputs(1059) <= a xor b;
    outputs(1060) <= not b or a;
    outputs(1061) <= b;
    outputs(1062) <= a xor b;
    outputs(1063) <= not b;
    outputs(1064) <= not a;
    outputs(1065) <= not b;
    outputs(1066) <= not (a xor b);
    outputs(1067) <= not (a xor b);
    outputs(1068) <= not b;
    outputs(1069) <= a;
    outputs(1070) <= a xor b;
    outputs(1071) <= not (a and b);
    outputs(1072) <= not (a xor b);
    outputs(1073) <= not b or a;
    outputs(1074) <= not b;
    outputs(1075) <= not (a or b);
    outputs(1076) <= a xor b;
    outputs(1077) <= not a;
    outputs(1078) <= b;
    outputs(1079) <= not a;
    outputs(1080) <= a;
    outputs(1081) <= not (a xor b);
    outputs(1082) <= not a or b;
    outputs(1083) <= a and not b;
    outputs(1084) <= not (a or b);
    outputs(1085) <= not b or a;
    outputs(1086) <= a and not b;
    outputs(1087) <= a and not b;
    outputs(1088) <= not (a xor b);
    outputs(1089) <= a or b;
    outputs(1090) <= not a;
    outputs(1091) <= b;
    outputs(1092) <= not b;
    outputs(1093) <= a xor b;
    outputs(1094) <= a and not b;
    outputs(1095) <= not (a xor b);
    outputs(1096) <= not b;
    outputs(1097) <= not b;
    outputs(1098) <= a and b;
    outputs(1099) <= not b;
    outputs(1100) <= not a;
    outputs(1101) <= not (a xor b);
    outputs(1102) <= a;
    outputs(1103) <= not a;
    outputs(1104) <= not a;
    outputs(1105) <= not (a or b);
    outputs(1106) <= a and not b;
    outputs(1107) <= a;
    outputs(1108) <= a and not b;
    outputs(1109) <= a;
    outputs(1110) <= a xor b;
    outputs(1111) <= not b;
    outputs(1112) <= b;
    outputs(1113) <= b;
    outputs(1114) <= not b;
    outputs(1115) <= not (a or b);
    outputs(1116) <= a;
    outputs(1117) <= a and not b;
    outputs(1118) <= not (a xor b);
    outputs(1119) <= b;
    outputs(1120) <= not a;
    outputs(1121) <= not a;
    outputs(1122) <= not b or a;
    outputs(1123) <= b;
    outputs(1124) <= not b;
    outputs(1125) <= a xor b;
    outputs(1126) <= a and not b;
    outputs(1127) <= not b;
    outputs(1128) <= a xor b;
    outputs(1129) <= not a or b;
    outputs(1130) <= b and not a;
    outputs(1131) <= not a;
    outputs(1132) <= a xor b;
    outputs(1133) <= a xor b;
    outputs(1134) <= a and not b;
    outputs(1135) <= a;
    outputs(1136) <= b and not a;
    outputs(1137) <= not (a xor b);
    outputs(1138) <= not b or a;
    outputs(1139) <= a;
    outputs(1140) <= a;
    outputs(1141) <= a xor b;
    outputs(1142) <= a xor b;
    outputs(1143) <= a and b;
    outputs(1144) <= not (a or b);
    outputs(1145) <= not (a xor b);
    outputs(1146) <= not (a or b);
    outputs(1147) <= not (a or b);
    outputs(1148) <= a;
    outputs(1149) <= not (a and b);
    outputs(1150) <= a and b;
    outputs(1151) <= a xor b;
    outputs(1152) <= b and not a;
    outputs(1153) <= a and b;
    outputs(1154) <= a xor b;
    outputs(1155) <= a;
    outputs(1156) <= a;
    outputs(1157) <= not b;
    outputs(1158) <= a;
    outputs(1159) <= not a;
    outputs(1160) <= not (a xor b);
    outputs(1161) <= a and not b;
    outputs(1162) <= a xor b;
    outputs(1163) <= not a;
    outputs(1164) <= not b;
    outputs(1165) <= a or b;
    outputs(1166) <= not b;
    outputs(1167) <= a;
    outputs(1168) <= not a;
    outputs(1169) <= a;
    outputs(1170) <= b;
    outputs(1171) <= not b;
    outputs(1172) <= not b;
    outputs(1173) <= not b;
    outputs(1174) <= b;
    outputs(1175) <= a xor b;
    outputs(1176) <= a xor b;
    outputs(1177) <= a or b;
    outputs(1178) <= not (a or b);
    outputs(1179) <= b;
    outputs(1180) <= not b;
    outputs(1181) <= a and b;
    outputs(1182) <= not a;
    outputs(1183) <= a xor b;
    outputs(1184) <= a xor b;
    outputs(1185) <= a;
    outputs(1186) <= b;
    outputs(1187) <= a and b;
    outputs(1188) <= b and not a;
    outputs(1189) <= a xor b;
    outputs(1190) <= b and not a;
    outputs(1191) <= not (a xor b);
    outputs(1192) <= not (a xor b);
    outputs(1193) <= not b or a;
    outputs(1194) <= a;
    outputs(1195) <= not a;
    outputs(1196) <= not a;
    outputs(1197) <= not a or b;
    outputs(1198) <= not (a xor b);
    outputs(1199) <= not (a xor b);
    outputs(1200) <= a xor b;
    outputs(1201) <= a xor b;
    outputs(1202) <= a and not b;
    outputs(1203) <= a xor b;
    outputs(1204) <= not (a xor b);
    outputs(1205) <= not (a xor b);
    outputs(1206) <= a xor b;
    outputs(1207) <= a and b;
    outputs(1208) <= a or b;
    outputs(1209) <= a and not b;
    outputs(1210) <= not (a xor b);
    outputs(1211) <= not b or a;
    outputs(1212) <= not (a xor b);
    outputs(1213) <= not (a xor b);
    outputs(1214) <= a and not b;
    outputs(1215) <= b;
    outputs(1216) <= a and not b;
    outputs(1217) <= not a;
    outputs(1218) <= a;
    outputs(1219) <= a;
    outputs(1220) <= not b;
    outputs(1221) <= a and not b;
    outputs(1222) <= not a;
    outputs(1223) <= b and not a;
    outputs(1224) <= not a;
    outputs(1225) <= b;
    outputs(1226) <= a;
    outputs(1227) <= a and b;
    outputs(1228) <= a and b;
    outputs(1229) <= a;
    outputs(1230) <= b;
    outputs(1231) <= not (a xor b);
    outputs(1232) <= a xor b;
    outputs(1233) <= not (a xor b);
    outputs(1234) <= a;
    outputs(1235) <= not a or b;
    outputs(1236) <= not b or a;
    outputs(1237) <= a;
    outputs(1238) <= not (a xor b);
    outputs(1239) <= a and b;
    outputs(1240) <= b;
    outputs(1241) <= a;
    outputs(1242) <= b and not a;
    outputs(1243) <= not a;
    outputs(1244) <= not b;
    outputs(1245) <= a xor b;
    outputs(1246) <= b;
    outputs(1247) <= not b;
    outputs(1248) <= not b;
    outputs(1249) <= not b;
    outputs(1250) <= b;
    outputs(1251) <= not a;
    outputs(1252) <= not b;
    outputs(1253) <= not (a and b);
    outputs(1254) <= a xor b;
    outputs(1255) <= a and not b;
    outputs(1256) <= a;
    outputs(1257) <= not (a xor b);
    outputs(1258) <= a xor b;
    outputs(1259) <= not (a and b);
    outputs(1260) <= not (a xor b);
    outputs(1261) <= not (a xor b);
    outputs(1262) <= not (a and b);
    outputs(1263) <= not b;
    outputs(1264) <= b;
    outputs(1265) <= a xor b;
    outputs(1266) <= not (a xor b);
    outputs(1267) <= not b;
    outputs(1268) <= not a;
    outputs(1269) <= a;
    outputs(1270) <= not (a or b);
    outputs(1271) <= b;
    outputs(1272) <= not a;
    outputs(1273) <= not (a and b);
    outputs(1274) <= a;
    outputs(1275) <= b and not a;
    outputs(1276) <= not (a and b);
    outputs(1277) <= not a;
    outputs(1278) <= not (a xor b);
    outputs(1279) <= a;
    outputs(1280) <= a and not b;
    outputs(1281) <= a or b;
    outputs(1282) <= a xor b;
    outputs(1283) <= a or b;
    outputs(1284) <= b;
    outputs(1285) <= not b;
    outputs(1286) <= a and b;
    outputs(1287) <= a xor b;
    outputs(1288) <= not a;
    outputs(1289) <= b;
    outputs(1290) <= not b;
    outputs(1291) <= not (a or b);
    outputs(1292) <= a;
    outputs(1293) <= a xor b;
    outputs(1294) <= not (a xor b);
    outputs(1295) <= not b;
    outputs(1296) <= a xor b;
    outputs(1297) <= not (a xor b);
    outputs(1298) <= not (a and b);
    outputs(1299) <= not b;
    outputs(1300) <= not (a xor b);
    outputs(1301) <= a and not b;
    outputs(1302) <= not b;
    outputs(1303) <= a xor b;
    outputs(1304) <= not (a or b);
    outputs(1305) <= not (a xor b);
    outputs(1306) <= a and b;
    outputs(1307) <= a and not b;
    outputs(1308) <= a;
    outputs(1309) <= not a;
    outputs(1310) <= not (a xor b);
    outputs(1311) <= a xor b;
    outputs(1312) <= a and not b;
    outputs(1313) <= a xor b;
    outputs(1314) <= not b or a;
    outputs(1315) <= b;
    outputs(1316) <= a and not b;
    outputs(1317) <= b;
    outputs(1318) <= a;
    outputs(1319) <= b;
    outputs(1320) <= not a or b;
    outputs(1321) <= not (a xor b);
    outputs(1322) <= not (a or b);
    outputs(1323) <= b;
    outputs(1324) <= a and b;
    outputs(1325) <= not (a xor b);
    outputs(1326) <= a xor b;
    outputs(1327) <= a xor b;
    outputs(1328) <= not b;
    outputs(1329) <= a;
    outputs(1330) <= a;
    outputs(1331) <= not a;
    outputs(1332) <= not a;
    outputs(1333) <= a xor b;
    outputs(1334) <= b;
    outputs(1335) <= a xor b;
    outputs(1336) <= not (a and b);
    outputs(1337) <= b;
    outputs(1338) <= a or b;
    outputs(1339) <= not a;
    outputs(1340) <= not a or b;
    outputs(1341) <= a or b;
    outputs(1342) <= a xor b;
    outputs(1343) <= not a or b;
    outputs(1344) <= not a;
    outputs(1345) <= a xor b;
    outputs(1346) <= not b or a;
    outputs(1347) <= not (a xor b);
    outputs(1348) <= b;
    outputs(1349) <= b;
    outputs(1350) <= a;
    outputs(1351) <= not a;
    outputs(1352) <= not b or a;
    outputs(1353) <= a;
    outputs(1354) <= a xor b;
    outputs(1355) <= a and not b;
    outputs(1356) <= not (a or b);
    outputs(1357) <= a;
    outputs(1358) <= b;
    outputs(1359) <= a or b;
    outputs(1360) <= a xor b;
    outputs(1361) <= not a;
    outputs(1362) <= b and not a;
    outputs(1363) <= b;
    outputs(1364) <= not a;
    outputs(1365) <= not (a or b);
    outputs(1366) <= not a;
    outputs(1367) <= a;
    outputs(1368) <= b;
    outputs(1369) <= b;
    outputs(1370) <= a or b;
    outputs(1371) <= b and not a;
    outputs(1372) <= a and b;
    outputs(1373) <= not b;
    outputs(1374) <= not b;
    outputs(1375) <= not b;
    outputs(1376) <= not (a xor b);
    outputs(1377) <= b;
    outputs(1378) <= a and b;
    outputs(1379) <= not a;
    outputs(1380) <= a xor b;
    outputs(1381) <= a and not b;
    outputs(1382) <= not b;
    outputs(1383) <= a;
    outputs(1384) <= a xor b;
    outputs(1385) <= a and b;
    outputs(1386) <= not b or a;
    outputs(1387) <= not (a and b);
    outputs(1388) <= not a;
    outputs(1389) <= a and not b;
    outputs(1390) <= not b;
    outputs(1391) <= not a;
    outputs(1392) <= a;
    outputs(1393) <= a xor b;
    outputs(1394) <= not a;
    outputs(1395) <= a or b;
    outputs(1396) <= a;
    outputs(1397) <= a and not b;
    outputs(1398) <= not a or b;
    outputs(1399) <= not (a xor b);
    outputs(1400) <= a xor b;
    outputs(1401) <= b and not a;
    outputs(1402) <= not (a xor b);
    outputs(1403) <= b;
    outputs(1404) <= b;
    outputs(1405) <= a and b;
    outputs(1406) <= not a;
    outputs(1407) <= a;
    outputs(1408) <= not b;
    outputs(1409) <= not a or b;
    outputs(1410) <= not a or b;
    outputs(1411) <= a or b;
    outputs(1412) <= b;
    outputs(1413) <= not a or b;
    outputs(1414) <= a;
    outputs(1415) <= b;
    outputs(1416) <= a;
    outputs(1417) <= not b;
    outputs(1418) <= a xor b;
    outputs(1419) <= b;
    outputs(1420) <= b;
    outputs(1421) <= not (a xor b);
    outputs(1422) <= a and b;
    outputs(1423) <= a and not b;
    outputs(1424) <= a xor b;
    outputs(1425) <= not (a and b);
    outputs(1426) <= a xor b;
    outputs(1427) <= not (a and b);
    outputs(1428) <= not a;
    outputs(1429) <= a;
    outputs(1430) <= a xor b;
    outputs(1431) <= not (a xor b);
    outputs(1432) <= not (a or b);
    outputs(1433) <= not (a xor b);
    outputs(1434) <= a and b;
    outputs(1435) <= a or b;
    outputs(1436) <= not (a xor b);
    outputs(1437) <= a xor b;
    outputs(1438) <= a;
    outputs(1439) <= not (a or b);
    outputs(1440) <= b and not a;
    outputs(1441) <= a;
    outputs(1442) <= b;
    outputs(1443) <= a xor b;
    outputs(1444) <= a;
    outputs(1445) <= a xor b;
    outputs(1446) <= a xor b;
    outputs(1447) <= not (a xor b);
    outputs(1448) <= not b;
    outputs(1449) <= not b;
    outputs(1450) <= not (a xor b);
    outputs(1451) <= a;
    outputs(1452) <= not b;
    outputs(1453) <= b and not a;
    outputs(1454) <= a and not b;
    outputs(1455) <= not a;
    outputs(1456) <= not (a and b);
    outputs(1457) <= not (a xor b);
    outputs(1458) <= a;
    outputs(1459) <= not (a xor b);
    outputs(1460) <= not b;
    outputs(1461) <= a and not b;
    outputs(1462) <= not a;
    outputs(1463) <= a;
    outputs(1464) <= a xor b;
    outputs(1465) <= a or b;
    outputs(1466) <= b;
    outputs(1467) <= a and b;
    outputs(1468) <= a xor b;
    outputs(1469) <= a xor b;
    outputs(1470) <= b and not a;
    outputs(1471) <= not b;
    outputs(1472) <= a;
    outputs(1473) <= a;
    outputs(1474) <= b;
    outputs(1475) <= a and not b;
    outputs(1476) <= not (a xor b);
    outputs(1477) <= not (a or b);
    outputs(1478) <= not (a or b);
    outputs(1479) <= b;
    outputs(1480) <= not b;
    outputs(1481) <= a and not b;
    outputs(1482) <= not a;
    outputs(1483) <= b and not a;
    outputs(1484) <= a xor b;
    outputs(1485) <= a;
    outputs(1486) <= not a;
    outputs(1487) <= not (a and b);
    outputs(1488) <= not b;
    outputs(1489) <= b;
    outputs(1490) <= not a;
    outputs(1491) <= a xor b;
    outputs(1492) <= a and not b;
    outputs(1493) <= not (a xor b);
    outputs(1494) <= not (a xor b);
    outputs(1495) <= not a;
    outputs(1496) <= not b;
    outputs(1497) <= not b;
    outputs(1498) <= a;
    outputs(1499) <= not (a xor b);
    outputs(1500) <= a and not b;
    outputs(1501) <= a and b;
    outputs(1502) <= a xor b;
    outputs(1503) <= a and not b;
    outputs(1504) <= a xor b;
    outputs(1505) <= b and not a;
    outputs(1506) <= not (a and b);
    outputs(1507) <= b;
    outputs(1508) <= not (a xor b);
    outputs(1509) <= a;
    outputs(1510) <= a and b;
    outputs(1511) <= not a;
    outputs(1512) <= b;
    outputs(1513) <= not (a or b);
    outputs(1514) <= a and not b;
    outputs(1515) <= not b;
    outputs(1516) <= not b;
    outputs(1517) <= a;
    outputs(1518) <= not a;
    outputs(1519) <= a;
    outputs(1520) <= b;
    outputs(1521) <= b;
    outputs(1522) <= a xor b;
    outputs(1523) <= not (a xor b);
    outputs(1524) <= a and not b;
    outputs(1525) <= not a;
    outputs(1526) <= a and b;
    outputs(1527) <= not (a xor b);
    outputs(1528) <= b;
    outputs(1529) <= not b or a;
    outputs(1530) <= a xor b;
    outputs(1531) <= b;
    outputs(1532) <= a xor b;
    outputs(1533) <= not b;
    outputs(1534) <= b;
    outputs(1535) <= not a;
    outputs(1536) <= a xor b;
    outputs(1537) <= not (a xor b);
    outputs(1538) <= a xor b;
    outputs(1539) <= a and b;
    outputs(1540) <= not b;
    outputs(1541) <= not (a or b);
    outputs(1542) <= a;
    outputs(1543) <= a;
    outputs(1544) <= not (a xor b);
    outputs(1545) <= not a;
    outputs(1546) <= b;
    outputs(1547) <= not a or b;
    outputs(1548) <= not (a or b);
    outputs(1549) <= not a;
    outputs(1550) <= a;
    outputs(1551) <= not (a and b);
    outputs(1552) <= b;
    outputs(1553) <= a xor b;
    outputs(1554) <= b and not a;
    outputs(1555) <= a;
    outputs(1556) <= b;
    outputs(1557) <= not (a or b);
    outputs(1558) <= a xor b;
    outputs(1559) <= b;
    outputs(1560) <= not b;
    outputs(1561) <= not (a or b);
    outputs(1562) <= a and b;
    outputs(1563) <= not b or a;
    outputs(1564) <= a and b;
    outputs(1565) <= b and not a;
    outputs(1566) <= b;
    outputs(1567) <= a xor b;
    outputs(1568) <= not (a xor b);
    outputs(1569) <= not (a or b);
    outputs(1570) <= not b or a;
    outputs(1571) <= not a;
    outputs(1572) <= a xor b;
    outputs(1573) <= not a;
    outputs(1574) <= b;
    outputs(1575) <= not (a or b);
    outputs(1576) <= b;
    outputs(1577) <= not (a or b);
    outputs(1578) <= not b or a;
    outputs(1579) <= not (a or b);
    outputs(1580) <= b and not a;
    outputs(1581) <= a xor b;
    outputs(1582) <= not a;
    outputs(1583) <= not (a and b);
    outputs(1584) <= b;
    outputs(1585) <= not (a xor b);
    outputs(1586) <= b;
    outputs(1587) <= not a;
    outputs(1588) <= not a;
    outputs(1589) <= not (a xor b);
    outputs(1590) <= a;
    outputs(1591) <= not a;
    outputs(1592) <= not (a or b);
    outputs(1593) <= not (a xor b);
    outputs(1594) <= not a;
    outputs(1595) <= a and b;
    outputs(1596) <= not b;
    outputs(1597) <= a and not b;
    outputs(1598) <= not b;
    outputs(1599) <= not (a or b);
    outputs(1600) <= not b;
    outputs(1601) <= not a;
    outputs(1602) <= a and not b;
    outputs(1603) <= not (a xor b);
    outputs(1604) <= a;
    outputs(1605) <= not b;
    outputs(1606) <= a;
    outputs(1607) <= not (a or b);
    outputs(1608) <= not b;
    outputs(1609) <= not b or a;
    outputs(1610) <= not a;
    outputs(1611) <= b and not a;
    outputs(1612) <= b and not a;
    outputs(1613) <= a xor b;
    outputs(1614) <= not a;
    outputs(1615) <= b and not a;
    outputs(1616) <= not b or a;
    outputs(1617) <= a;
    outputs(1618) <= not b;
    outputs(1619) <= not b;
    outputs(1620) <= b and not a;
    outputs(1621) <= not (a xor b);
    outputs(1622) <= not (a xor b);
    outputs(1623) <= a;
    outputs(1624) <= a and b;
    outputs(1625) <= not (a xor b);
    outputs(1626) <= not a or b;
    outputs(1627) <= b and not a;
    outputs(1628) <= b;
    outputs(1629) <= not b;
    outputs(1630) <= a xor b;
    outputs(1631) <= b and not a;
    outputs(1632) <= not b;
    outputs(1633) <= a;
    outputs(1634) <= not b or a;
    outputs(1635) <= not (a xor b);
    outputs(1636) <= not (a xor b);
    outputs(1637) <= not a;
    outputs(1638) <= not (a xor b);
    outputs(1639) <= not (a xor b);
    outputs(1640) <= a;
    outputs(1641) <= a;
    outputs(1642) <= a and not b;
    outputs(1643) <= a;
    outputs(1644) <= a and b;
    outputs(1645) <= a and b;
    outputs(1646) <= not a or b;
    outputs(1647) <= not (a xor b);
    outputs(1648) <= not (a xor b);
    outputs(1649) <= not (a or b);
    outputs(1650) <= a and b;
    outputs(1651) <= b;
    outputs(1652) <= a and b;
    outputs(1653) <= not a or b;
    outputs(1654) <= not (a or b);
    outputs(1655) <= not a;
    outputs(1656) <= not a;
    outputs(1657) <= a;
    outputs(1658) <= not b;
    outputs(1659) <= a;
    outputs(1660) <= b;
    outputs(1661) <= not b;
    outputs(1662) <= a;
    outputs(1663) <= a;
    outputs(1664) <= not b;
    outputs(1665) <= a;
    outputs(1666) <= b and not a;
    outputs(1667) <= not a;
    outputs(1668) <= not b;
    outputs(1669) <= not a;
    outputs(1670) <= b;
    outputs(1671) <= a and not b;
    outputs(1672) <= a xor b;
    outputs(1673) <= not (a xor b);
    outputs(1674) <= b;
    outputs(1675) <= not (a xor b);
    outputs(1676) <= b;
    outputs(1677) <= not a or b;
    outputs(1678) <= not (a xor b);
    outputs(1679) <= a and not b;
    outputs(1680) <= a and b;
    outputs(1681) <= not a or b;
    outputs(1682) <= not a;
    outputs(1683) <= b;
    outputs(1684) <= a;
    outputs(1685) <= b;
    outputs(1686) <= a;
    outputs(1687) <= not a;
    outputs(1688) <= not a;
    outputs(1689) <= a and not b;
    outputs(1690) <= not a or b;
    outputs(1691) <= a and not b;
    outputs(1692) <= b and not a;
    outputs(1693) <= a;
    outputs(1694) <= not a;
    outputs(1695) <= a xor b;
    outputs(1696) <= not a;
    outputs(1697) <= not a;
    outputs(1698) <= a;
    outputs(1699) <= not a;
    outputs(1700) <= not (a or b);
    outputs(1701) <= a and b;
    outputs(1702) <= a xor b;
    outputs(1703) <= not (a or b);
    outputs(1704) <= not (a or b);
    outputs(1705) <= a;
    outputs(1706) <= not b;
    outputs(1707) <= not b or a;
    outputs(1708) <= not a or b;
    outputs(1709) <= not (a and b);
    outputs(1710) <= a and not b;
    outputs(1711) <= a;
    outputs(1712) <= b;
    outputs(1713) <= b and not a;
    outputs(1714) <= a and not b;
    outputs(1715) <= a xor b;
    outputs(1716) <= a xor b;
    outputs(1717) <= b;
    outputs(1718) <= a and b;
    outputs(1719) <= b and not a;
    outputs(1720) <= not (a xor b);
    outputs(1721) <= b and not a;
    outputs(1722) <= a and b;
    outputs(1723) <= a and b;
    outputs(1724) <= not b;
    outputs(1725) <= not (a xor b);
    outputs(1726) <= not b;
    outputs(1727) <= a;
    outputs(1728) <= a xor b;
    outputs(1729) <= a and not b;
    outputs(1730) <= a or b;
    outputs(1731) <= a and not b;
    outputs(1732) <= a;
    outputs(1733) <= not a;
    outputs(1734) <= not (a xor b);
    outputs(1735) <= b;
    outputs(1736) <= a xor b;
    outputs(1737) <= a and b;
    outputs(1738) <= a;
    outputs(1739) <= a xor b;
    outputs(1740) <= not (a or b);
    outputs(1741) <= not b;
    outputs(1742) <= b;
    outputs(1743) <= a and b;
    outputs(1744) <= not b;
    outputs(1745) <= a;
    outputs(1746) <= a;
    outputs(1747) <= b;
    outputs(1748) <= a;
    outputs(1749) <= not a;
    outputs(1750) <= not b;
    outputs(1751) <= b and not a;
    outputs(1752) <= b and not a;
    outputs(1753) <= b and not a;
    outputs(1754) <= a and b;
    outputs(1755) <= a xor b;
    outputs(1756) <= b and not a;
    outputs(1757) <= a or b;
    outputs(1758) <= not a;
    outputs(1759) <= not a;
    outputs(1760) <= a xor b;
    outputs(1761) <= not (a xor b);
    outputs(1762) <= b and not a;
    outputs(1763) <= not a;
    outputs(1764) <= a xor b;
    outputs(1765) <= not a;
    outputs(1766) <= a;
    outputs(1767) <= a and not b;
    outputs(1768) <= not (a xor b);
    outputs(1769) <= b and not a;
    outputs(1770) <= not (a xor b);
    outputs(1771) <= a and not b;
    outputs(1772) <= b;
    outputs(1773) <= not (a or b);
    outputs(1774) <= not (a xor b);
    outputs(1775) <= not (a xor b);
    outputs(1776) <= b;
    outputs(1777) <= not a;
    outputs(1778) <= a and not b;
    outputs(1779) <= not b;
    outputs(1780) <= b;
    outputs(1781) <= a;
    outputs(1782) <= a xor b;
    outputs(1783) <= a xor b;
    outputs(1784) <= a xor b;
    outputs(1785) <= not a;
    outputs(1786) <= a xor b;
    outputs(1787) <= a;
    outputs(1788) <= a and b;
    outputs(1789) <= not b;
    outputs(1790) <= a xor b;
    outputs(1791) <= not a;
    outputs(1792) <= not (a or b);
    outputs(1793) <= a xor b;
    outputs(1794) <= not (a xor b);
    outputs(1795) <= a;
    outputs(1796) <= b and not a;
    outputs(1797) <= b;
    outputs(1798) <= b;
    outputs(1799) <= a;
    outputs(1800) <= not a;
    outputs(1801) <= a and b;
    outputs(1802) <= not (a xor b);
    outputs(1803) <= not a;
    outputs(1804) <= not a;
    outputs(1805) <= b;
    outputs(1806) <= a and b;
    outputs(1807) <= not a;
    outputs(1808) <= not b;
    outputs(1809) <= not (a xor b);
    outputs(1810) <= a or b;
    outputs(1811) <= not b or a;
    outputs(1812) <= b and not a;
    outputs(1813) <= b;
    outputs(1814) <= not b or a;
    outputs(1815) <= not (a xor b);
    outputs(1816) <= a xor b;
    outputs(1817) <= a xor b;
    outputs(1818) <= a and b;
    outputs(1819) <= not (a xor b);
    outputs(1820) <= b;
    outputs(1821) <= not (a or b);
    outputs(1822) <= not b or a;
    outputs(1823) <= not a;
    outputs(1824) <= not (a or b);
    outputs(1825) <= not (a and b);
    outputs(1826) <= not (a xor b);
    outputs(1827) <= a;
    outputs(1828) <= a;
    outputs(1829) <= b;
    outputs(1830) <= a;
    outputs(1831) <= b and not a;
    outputs(1832) <= not b;
    outputs(1833) <= a;
    outputs(1834) <= not a;
    outputs(1835) <= b;
    outputs(1836) <= a xor b;
    outputs(1837) <= not a;
    outputs(1838) <= b;
    outputs(1839) <= not b or a;
    outputs(1840) <= a xor b;
    outputs(1841) <= not (a xor b);
    outputs(1842) <= a;
    outputs(1843) <= not (a xor b);
    outputs(1844) <= not (a and b);
    outputs(1845) <= b;
    outputs(1846) <= a and not b;
    outputs(1847) <= a;
    outputs(1848) <= a;
    outputs(1849) <= b;
    outputs(1850) <= a or b;
    outputs(1851) <= a xor b;
    outputs(1852) <= a and b;
    outputs(1853) <= not b;
    outputs(1854) <= not (a xor b);
    outputs(1855) <= not (a xor b);
    outputs(1856) <= b;
    outputs(1857) <= a and b;
    outputs(1858) <= not a;
    outputs(1859) <= not b;
    outputs(1860) <= not a or b;
    outputs(1861) <= a or b;
    outputs(1862) <= a and not b;
    outputs(1863) <= a;
    outputs(1864) <= not a;
    outputs(1865) <= not b;
    outputs(1866) <= not (a or b);
    outputs(1867) <= a and b;
    outputs(1868) <= a and b;
    outputs(1869) <= not b;
    outputs(1870) <= a xor b;
    outputs(1871) <= not (a xor b);
    outputs(1872) <= b and not a;
    outputs(1873) <= a and b;
    outputs(1874) <= not a;
    outputs(1875) <= not (a xor b);
    outputs(1876) <= b and not a;
    outputs(1877) <= a xor b;
    outputs(1878) <= a and b;
    outputs(1879) <= not b;
    outputs(1880) <= a xor b;
    outputs(1881) <= not a or b;
    outputs(1882) <= not a;
    outputs(1883) <= a xor b;
    outputs(1884) <= b and not a;
    outputs(1885) <= not (a xor b);
    outputs(1886) <= a and not b;
    outputs(1887) <= not b;
    outputs(1888) <= a or b;
    outputs(1889) <= b;
    outputs(1890) <= a xor b;
    outputs(1891) <= a;
    outputs(1892) <= not a;
    outputs(1893) <= not (a or b);
    outputs(1894) <= a xor b;
    outputs(1895) <= not a;
    outputs(1896) <= b;
    outputs(1897) <= a and not b;
    outputs(1898) <= b;
    outputs(1899) <= a;
    outputs(1900) <= a and b;
    outputs(1901) <= not (a xor b);
    outputs(1902) <= not b;
    outputs(1903) <= not a;
    outputs(1904) <= not a;
    outputs(1905) <= a;
    outputs(1906) <= not a or b;
    outputs(1907) <= b and not a;
    outputs(1908) <= a;
    outputs(1909) <= a xor b;
    outputs(1910) <= not b;
    outputs(1911) <= b;
    outputs(1912) <= a or b;
    outputs(1913) <= not b;
    outputs(1914) <= not a;
    outputs(1915) <= b;
    outputs(1916) <= not (a and b);
    outputs(1917) <= a;
    outputs(1918) <= a;
    outputs(1919) <= not (a xor b);
    outputs(1920) <= not (a xor b);
    outputs(1921) <= not a;
    outputs(1922) <= a and not b;
    outputs(1923) <= not b or a;
    outputs(1924) <= a;
    outputs(1925) <= not (a xor b);
    outputs(1926) <= not a or b;
    outputs(1927) <= not (a xor b);
    outputs(1928) <= not b;
    outputs(1929) <= not b or a;
    outputs(1930) <= a xor b;
    outputs(1931) <= not b;
    outputs(1932) <= not b;
    outputs(1933) <= b;
    outputs(1934) <= a xor b;
    outputs(1935) <= b and not a;
    outputs(1936) <= b;
    outputs(1937) <= a and b;
    outputs(1938) <= a or b;
    outputs(1939) <= a;
    outputs(1940) <= b;
    outputs(1941) <= b;
    outputs(1942) <= not a;
    outputs(1943) <= not b;
    outputs(1944) <= a and b;
    outputs(1945) <= not (a xor b);
    outputs(1946) <= not a;
    outputs(1947) <= not (a xor b);
    outputs(1948) <= b;
    outputs(1949) <= a and not b;
    outputs(1950) <= b and not a;
    outputs(1951) <= b;
    outputs(1952) <= a;
    outputs(1953) <= not a;
    outputs(1954) <= a xor b;
    outputs(1955) <= a and b;
    outputs(1956) <= b;
    outputs(1957) <= a;
    outputs(1958) <= a xor b;
    outputs(1959) <= not a;
    outputs(1960) <= a and b;
    outputs(1961) <= a xor b;
    outputs(1962) <= a and not b;
    outputs(1963) <= not (a or b);
    outputs(1964) <= not b;
    outputs(1965) <= a and not b;
    outputs(1966) <= a;
    outputs(1967) <= not b;
    outputs(1968) <= not b;
    outputs(1969) <= not b;
    outputs(1970) <= not a or b;
    outputs(1971) <= b and not a;
    outputs(1972) <= not a;
    outputs(1973) <= not (a xor b);
    outputs(1974) <= a;
    outputs(1975) <= not (a or b);
    outputs(1976) <= a xor b;
    outputs(1977) <= a xor b;
    outputs(1978) <= a xor b;
    outputs(1979) <= b;
    outputs(1980) <= a xor b;
    outputs(1981) <= not a or b;
    outputs(1982) <= a or b;
    outputs(1983) <= a;
    outputs(1984) <= a and not b;
    outputs(1985) <= a xor b;
    outputs(1986) <= b;
    outputs(1987) <= not (a xor b);
    outputs(1988) <= not (a xor b);
    outputs(1989) <= a;
    outputs(1990) <= not a;
    outputs(1991) <= not (a and b);
    outputs(1992) <= a and not b;
    outputs(1993) <= a xor b;
    outputs(1994) <= not a;
    outputs(1995) <= not (a and b);
    outputs(1996) <= b;
    outputs(1997) <= a and b;
    outputs(1998) <= b and not a;
    outputs(1999) <= a and b;
    outputs(2000) <= a and b;
    outputs(2001) <= a and not b;
    outputs(2002) <= b;
    outputs(2003) <= a and b;
    outputs(2004) <= not b;
    outputs(2005) <= b;
    outputs(2006) <= a xor b;
    outputs(2007) <= b and not a;
    outputs(2008) <= b and not a;
    outputs(2009) <= a xor b;
    outputs(2010) <= a and b;
    outputs(2011) <= not (a xor b);
    outputs(2012) <= a;
    outputs(2013) <= not b or a;
    outputs(2014) <= a;
    outputs(2015) <= not (a xor b);
    outputs(2016) <= a xor b;
    outputs(2017) <= not (a xor b);
    outputs(2018) <= not b;
    outputs(2019) <= a;
    outputs(2020) <= not a;
    outputs(2021) <= not a;
    outputs(2022) <= not a;
    outputs(2023) <= a;
    outputs(2024) <= b;
    outputs(2025) <= not a;
    outputs(2026) <= not (a xor b);
    outputs(2027) <= a and not b;
    outputs(2028) <= not (a xor b);
    outputs(2029) <= not (a xor b);
    outputs(2030) <= a or b;
    outputs(2031) <= not b;
    outputs(2032) <= b;
    outputs(2033) <= not (a xor b);
    outputs(2034) <= a xor b;
    outputs(2035) <= a;
    outputs(2036) <= a or b;
    outputs(2037) <= not (a xor b);
    outputs(2038) <= b and not a;
    outputs(2039) <= not a;
    outputs(2040) <= not b or a;
    outputs(2041) <= a;
    outputs(2042) <= a;
    outputs(2043) <= not b;
    outputs(2044) <= not (a or b);
    outputs(2045) <= a;
    outputs(2046) <= not a;
    outputs(2047) <= not (a xor b);
    outputs(2048) <= b and not a;
    outputs(2049) <= not a;
    outputs(2050) <= not a or b;
    outputs(2051) <= a xor b;
    outputs(2052) <= a;
    outputs(2053) <= not b;
    outputs(2054) <= a and b;
    outputs(2055) <= a xor b;
    outputs(2056) <= b and not a;
    outputs(2057) <= not b;
    outputs(2058) <= not (a xor b);
    outputs(2059) <= a;
    outputs(2060) <= b and not a;
    outputs(2061) <= a xor b;
    outputs(2062) <= not (a xor b);
    outputs(2063) <= a xor b;
    outputs(2064) <= not a or b;
    outputs(2065) <= a xor b;
    outputs(2066) <= a xor b;
    outputs(2067) <= b;
    outputs(2068) <= a;
    outputs(2069) <= not (a xor b);
    outputs(2070) <= a and not b;
    outputs(2071) <= not (a xor b);
    outputs(2072) <= not b or a;
    outputs(2073) <= a;
    outputs(2074) <= not (a xor b);
    outputs(2075) <= a xor b;
    outputs(2076) <= not a;
    outputs(2077) <= a and b;
    outputs(2078) <= not b;
    outputs(2079) <= a;
    outputs(2080) <= not b;
    outputs(2081) <= a and not b;
    outputs(2082) <= not a;
    outputs(2083) <= not (a or b);
    outputs(2084) <= not (a or b);
    outputs(2085) <= a xor b;
    outputs(2086) <= b;
    outputs(2087) <= not b;
    outputs(2088) <= not (a or b);
    outputs(2089) <= not a;
    outputs(2090) <= not (a or b);
    outputs(2091) <= a;
    outputs(2092) <= not (a xor b);
    outputs(2093) <= not (a xor b);
    outputs(2094) <= not b;
    outputs(2095) <= b;
    outputs(2096) <= not a;
    outputs(2097) <= not (a xor b);
    outputs(2098) <= not a;
    outputs(2099) <= a and not b;
    outputs(2100) <= not b;
    outputs(2101) <= not (a or b);
    outputs(2102) <= a and not b;
    outputs(2103) <= not (a or b);
    outputs(2104) <= b;
    outputs(2105) <= not b;
    outputs(2106) <= not (a xor b);
    outputs(2107) <= not (a xor b);
    outputs(2108) <= a and not b;
    outputs(2109) <= b;
    outputs(2110) <= not b;
    outputs(2111) <= b;
    outputs(2112) <= not (a xor b);
    outputs(2113) <= b and not a;
    outputs(2114) <= b;
    outputs(2115) <= not a;
    outputs(2116) <= b;
    outputs(2117) <= a xor b;
    outputs(2118) <= not a;
    outputs(2119) <= b;
    outputs(2120) <= not b;
    outputs(2121) <= a xor b;
    outputs(2122) <= b;
    outputs(2123) <= not b;
    outputs(2124) <= b;
    outputs(2125) <= not (a and b);
    outputs(2126) <= not a or b;
    outputs(2127) <= a xor b;
    outputs(2128) <= not b;
    outputs(2129) <= not (a xor b);
    outputs(2130) <= a or b;
    outputs(2131) <= not (a xor b);
    outputs(2132) <= not (a and b);
    outputs(2133) <= b;
    outputs(2134) <= b;
    outputs(2135) <= not (a or b);
    outputs(2136) <= not (a and b);
    outputs(2137) <= not (a and b);
    outputs(2138) <= a xor b;
    outputs(2139) <= not a or b;
    outputs(2140) <= not b;
    outputs(2141) <= not a;
    outputs(2142) <= a xor b;
    outputs(2143) <= not b;
    outputs(2144) <= a or b;
    outputs(2145) <= not (a xor b);
    outputs(2146) <= b;
    outputs(2147) <= not a;
    outputs(2148) <= a;
    outputs(2149) <= not (a xor b);
    outputs(2150) <= a xor b;
    outputs(2151) <= not a;
    outputs(2152) <= not (a xor b);
    outputs(2153) <= b;
    outputs(2154) <= not b;
    outputs(2155) <= a and not b;
    outputs(2156) <= not a;
    outputs(2157) <= a and not b;
    outputs(2158) <= a;
    outputs(2159) <= not (a xor b);
    outputs(2160) <= a xor b;
    outputs(2161) <= a;
    outputs(2162) <= a;
    outputs(2163) <= a xor b;
    outputs(2164) <= not (a xor b);
    outputs(2165) <= not a;
    outputs(2166) <= a xor b;
    outputs(2167) <= a and b;
    outputs(2168) <= not (a xor b);
    outputs(2169) <= a xor b;
    outputs(2170) <= not (a or b);
    outputs(2171) <= not a;
    outputs(2172) <= b and not a;
    outputs(2173) <= not b;
    outputs(2174) <= a xor b;
    outputs(2175) <= a and not b;
    outputs(2176) <= b;
    outputs(2177) <= b;
    outputs(2178) <= a or b;
    outputs(2179) <= a or b;
    outputs(2180) <= not (a xor b);
    outputs(2181) <= not a;
    outputs(2182) <= a xor b;
    outputs(2183) <= a;
    outputs(2184) <= a;
    outputs(2185) <= a;
    outputs(2186) <= not (a xor b);
    outputs(2187) <= a;
    outputs(2188) <= not (a xor b);
    outputs(2189) <= not b;
    outputs(2190) <= a or b;
    outputs(2191) <= not (a xor b);
    outputs(2192) <= not b;
    outputs(2193) <= a xor b;
    outputs(2194) <= a and not b;
    outputs(2195) <= not (a xor b);
    outputs(2196) <= not b or a;
    outputs(2197) <= b and not a;
    outputs(2198) <= a;
    outputs(2199) <= b;
    outputs(2200) <= b;
    outputs(2201) <= not b;
    outputs(2202) <= not (a xor b);
    outputs(2203) <= b;
    outputs(2204) <= b and not a;
    outputs(2205) <= not (a xor b);
    outputs(2206) <= not a;
    outputs(2207) <= not (a xor b);
    outputs(2208) <= not (a xor b);
    outputs(2209) <= a;
    outputs(2210) <= b and not a;
    outputs(2211) <= a xor b;
    outputs(2212) <= b;
    outputs(2213) <= not a;
    outputs(2214) <= a and not b;
    outputs(2215) <= b;
    outputs(2216) <= a;
    outputs(2217) <= a;
    outputs(2218) <= b and not a;
    outputs(2219) <= b and not a;
    outputs(2220) <= not b;
    outputs(2221) <= a xor b;
    outputs(2222) <= b;
    outputs(2223) <= a xor b;
    outputs(2224) <= a xor b;
    outputs(2225) <= not (a xor b);
    outputs(2226) <= not b;
    outputs(2227) <= not (a xor b);
    outputs(2228) <= not b;
    outputs(2229) <= a xor b;
    outputs(2230) <= a xor b;
    outputs(2231) <= b;
    outputs(2232) <= not b;
    outputs(2233) <= not b;
    outputs(2234) <= not b;
    outputs(2235) <= not a;
    outputs(2236) <= b;
    outputs(2237) <= not (a xor b);
    outputs(2238) <= a or b;
    outputs(2239) <= not a;
    outputs(2240) <= b;
    outputs(2241) <= a xor b;
    outputs(2242) <= not b;
    outputs(2243) <= b;
    outputs(2244) <= a;
    outputs(2245) <= a and not b;
    outputs(2246) <= not b;
    outputs(2247) <= b and not a;
    outputs(2248) <= not (a xor b);
    outputs(2249) <= a;
    outputs(2250) <= a;
    outputs(2251) <= not b;
    outputs(2252) <= a;
    outputs(2253) <= not b or a;
    outputs(2254) <= a and not b;
    outputs(2255) <= not (a or b);
    outputs(2256) <= not (a xor b);
    outputs(2257) <= a;
    outputs(2258) <= a xor b;
    outputs(2259) <= not a;
    outputs(2260) <= a;
    outputs(2261) <= not (a or b);
    outputs(2262) <= a and not b;
    outputs(2263) <= a and not b;
    outputs(2264) <= not a;
    outputs(2265) <= not (a or b);
    outputs(2266) <= not a;
    outputs(2267) <= not b;
    outputs(2268) <= b and not a;
    outputs(2269) <= a;
    outputs(2270) <= not a;
    outputs(2271) <= not a;
    outputs(2272) <= not (a or b);
    outputs(2273) <= a and b;
    outputs(2274) <= not a;
    outputs(2275) <= not a;
    outputs(2276) <= not b;
    outputs(2277) <= a xor b;
    outputs(2278) <= b;
    outputs(2279) <= a xor b;
    outputs(2280) <= a and b;
    outputs(2281) <= not a;
    outputs(2282) <= not b or a;
    outputs(2283) <= a xor b;
    outputs(2284) <= not b;
    outputs(2285) <= a xor b;
    outputs(2286) <= not b;
    outputs(2287) <= not (a xor b);
    outputs(2288) <= b and not a;
    outputs(2289) <= b;
    outputs(2290) <= not b;
    outputs(2291) <= a;
    outputs(2292) <= not (a or b);
    outputs(2293) <= a;
    outputs(2294) <= not a;
    outputs(2295) <= a and b;
    outputs(2296) <= b;
    outputs(2297) <= not a;
    outputs(2298) <= a xor b;
    outputs(2299) <= a;
    outputs(2300) <= not (a xor b);
    outputs(2301) <= a and not b;
    outputs(2302) <= a;
    outputs(2303) <= not b;
    outputs(2304) <= b;
    outputs(2305) <= not a;
    outputs(2306) <= not (a xor b);
    outputs(2307) <= a or b;
    outputs(2308) <= not (a xor b);
    outputs(2309) <= b;
    outputs(2310) <= a;
    outputs(2311) <= not a;
    outputs(2312) <= a xor b;
    outputs(2313) <= not (a and b);
    outputs(2314) <= not (a or b);
    outputs(2315) <= not a or b;
    outputs(2316) <= b;
    outputs(2317) <= not (a xor b);
    outputs(2318) <= a;
    outputs(2319) <= not b;
    outputs(2320) <= a;
    outputs(2321) <= a;
    outputs(2322) <= not a;
    outputs(2323) <= a;
    outputs(2324) <= a;
    outputs(2325) <= b;
    outputs(2326) <= a xor b;
    outputs(2327) <= not b;
    outputs(2328) <= not a;
    outputs(2329) <= not b;
    outputs(2330) <= a;
    outputs(2331) <= not (a xor b);
    outputs(2332) <= a xor b;
    outputs(2333) <= a;
    outputs(2334) <= a xor b;
    outputs(2335) <= not a;
    outputs(2336) <= a and not b;
    outputs(2337) <= not (a or b);
    outputs(2338) <= a and b;
    outputs(2339) <= b;
    outputs(2340) <= not (a or b);
    outputs(2341) <= a xor b;
    outputs(2342) <= not (a xor b);
    outputs(2343) <= a and b;
    outputs(2344) <= a and not b;
    outputs(2345) <= not (a and b);
    outputs(2346) <= not (a xor b);
    outputs(2347) <= a xor b;
    outputs(2348) <= not b;
    outputs(2349) <= a;
    outputs(2350) <= not a;
    outputs(2351) <= b;
    outputs(2352) <= not a or b;
    outputs(2353) <= not b;
    outputs(2354) <= a;
    outputs(2355) <= b and not a;
    outputs(2356) <= a xor b;
    outputs(2357) <= a and b;
    outputs(2358) <= not b;
    outputs(2359) <= a and b;
    outputs(2360) <= not b;
    outputs(2361) <= b;
    outputs(2362) <= a xor b;
    outputs(2363) <= not (a or b);
    outputs(2364) <= not b or a;
    outputs(2365) <= not a;
    outputs(2366) <= not a;
    outputs(2367) <= not a;
    outputs(2368) <= not (a xor b);
    outputs(2369) <= not a;
    outputs(2370) <= not a;
    outputs(2371) <= not b;
    outputs(2372) <= a xor b;
    outputs(2373) <= not b;
    outputs(2374) <= not a;
    outputs(2375) <= a and b;
    outputs(2376) <= a xor b;
    outputs(2377) <= a xor b;
    outputs(2378) <= a or b;
    outputs(2379) <= not b;
    outputs(2380) <= b and not a;
    outputs(2381) <= not b or a;
    outputs(2382) <= a xor b;
    outputs(2383) <= not (a xor b);
    outputs(2384) <= b and not a;
    outputs(2385) <= not b;
    outputs(2386) <= not (a xor b);
    outputs(2387) <= a and b;
    outputs(2388) <= not a;
    outputs(2389) <= not (a xor b);
    outputs(2390) <= a xor b;
    outputs(2391) <= a;
    outputs(2392) <= not (a or b);
    outputs(2393) <= not (a xor b);
    outputs(2394) <= not b or a;
    outputs(2395) <= a;
    outputs(2396) <= a xor b;
    outputs(2397) <= a;
    outputs(2398) <= not (a or b);
    outputs(2399) <= not a;
    outputs(2400) <= not a or b;
    outputs(2401) <= a;
    outputs(2402) <= not a;
    outputs(2403) <= not b;
    outputs(2404) <= not (a xor b);
    outputs(2405) <= b and not a;
    outputs(2406) <= not a;
    outputs(2407) <= a;
    outputs(2408) <= not b;
    outputs(2409) <= b;
    outputs(2410) <= not b;
    outputs(2411) <= not (a xor b);
    outputs(2412) <= not b;
    outputs(2413) <= a;
    outputs(2414) <= b;
    outputs(2415) <= not b;
    outputs(2416) <= not a;
    outputs(2417) <= a and not b;
    outputs(2418) <= not a;
    outputs(2419) <= not a;
    outputs(2420) <= a and not b;
    outputs(2421) <= not (a or b);
    outputs(2422) <= not b;
    outputs(2423) <= a and b;
    outputs(2424) <= a;
    outputs(2425) <= not b;
    outputs(2426) <= a xor b;
    outputs(2427) <= a;
    outputs(2428) <= b and not a;
    outputs(2429) <= not (a xor b);
    outputs(2430) <= b;
    outputs(2431) <= a and not b;
    outputs(2432) <= not b;
    outputs(2433) <= b and not a;
    outputs(2434) <= not b;
    outputs(2435) <= a and b;
    outputs(2436) <= not (a xor b);
    outputs(2437) <= b;
    outputs(2438) <= not b;
    outputs(2439) <= not b;
    outputs(2440) <= a and b;
    outputs(2441) <= b;
    outputs(2442) <= b;
    outputs(2443) <= a;
    outputs(2444) <= a xor b;
    outputs(2445) <= a and b;
    outputs(2446) <= a or b;
    outputs(2447) <= not (a xor b);
    outputs(2448) <= not a;
    outputs(2449) <= a or b;
    outputs(2450) <= a and not b;
    outputs(2451) <= not b;
    outputs(2452) <= b;
    outputs(2453) <= a or b;
    outputs(2454) <= a xor b;
    outputs(2455) <= a and b;
    outputs(2456) <= a xor b;
    outputs(2457) <= a xor b;
    outputs(2458) <= not b;
    outputs(2459) <= a or b;
    outputs(2460) <= b and not a;
    outputs(2461) <= not a;
    outputs(2462) <= a and not b;
    outputs(2463) <= a xor b;
    outputs(2464) <= a and b;
    outputs(2465) <= not a;
    outputs(2466) <= not a or b;
    outputs(2467) <= not a;
    outputs(2468) <= not b;
    outputs(2469) <= a;
    outputs(2470) <= a xor b;
    outputs(2471) <= a xor b;
    outputs(2472) <= a xor b;
    outputs(2473) <= not a;
    outputs(2474) <= not (a xor b);
    outputs(2475) <= a xor b;
    outputs(2476) <= not b;
    outputs(2477) <= not a or b;
    outputs(2478) <= a;
    outputs(2479) <= a and not b;
    outputs(2480) <= b;
    outputs(2481) <= b;
    outputs(2482) <= not a;
    outputs(2483) <= not a;
    outputs(2484) <= a xor b;
    outputs(2485) <= b;
    outputs(2486) <= not a;
    outputs(2487) <= not a;
    outputs(2488) <= not a or b;
    outputs(2489) <= not a;
    outputs(2490) <= not a;
    outputs(2491) <= not a;
    outputs(2492) <= not a;
    outputs(2493) <= not a;
    outputs(2494) <= not (a xor b);
    outputs(2495) <= b;
    outputs(2496) <= not a;
    outputs(2497) <= not a;
    outputs(2498) <= a and not b;
    outputs(2499) <= not a;
    outputs(2500) <= not (a xor b);
    outputs(2501) <= not (a xor b);
    outputs(2502) <= not a;
    outputs(2503) <= a;
    outputs(2504) <= b;
    outputs(2505) <= not b;
    outputs(2506) <= not a;
    outputs(2507) <= b;
    outputs(2508) <= a xor b;
    outputs(2509) <= a xor b;
    outputs(2510) <= not a;
    outputs(2511) <= a xor b;
    outputs(2512) <= not a or b;
    outputs(2513) <= b and not a;
    outputs(2514) <= not (a or b);
    outputs(2515) <= b and not a;
    outputs(2516) <= a;
    outputs(2517) <= not b;
    outputs(2518) <= not (a or b);
    outputs(2519) <= a;
    outputs(2520) <= not (a or b);
    outputs(2521) <= a xor b;
    outputs(2522) <= a xor b;
    outputs(2523) <= a xor b;
    outputs(2524) <= not a or b;
    outputs(2525) <= a xor b;
    outputs(2526) <= not (a or b);
    outputs(2527) <= not a;
    outputs(2528) <= a xor b;
    outputs(2529) <= not a;
    outputs(2530) <= not b;
    outputs(2531) <= not (a or b);
    outputs(2532) <= a and b;
    outputs(2533) <= a;
    outputs(2534) <= b and not a;
    outputs(2535) <= a and not b;
    outputs(2536) <= not b;
    outputs(2537) <= not b;
    outputs(2538) <= not b;
    outputs(2539) <= not b;
    outputs(2540) <= not a;
    outputs(2541) <= b and not a;
    outputs(2542) <= not b;
    outputs(2543) <= not (a xor b);
    outputs(2544) <= not (a or b);
    outputs(2545) <= not a;
    outputs(2546) <= not b;
    outputs(2547) <= b and not a;
    outputs(2548) <= a;
    outputs(2549) <= not a;
    outputs(2550) <= a;
    outputs(2551) <= not b;
    outputs(2552) <= a xor b;
    outputs(2553) <= a and b;
    outputs(2554) <= not (a xor b);
    outputs(2555) <= a xor b;
    outputs(2556) <= not a;
    outputs(2557) <= a xor b;
    outputs(2558) <= a and not b;
    outputs(2559) <= a and b;
    outputs(2560) <= not a;
    outputs(2561) <= not (a xor b);
    outputs(2562) <= a;
    outputs(2563) <= not (a xor b);
    outputs(2564) <= a;
    outputs(2565) <= a;
    outputs(2566) <= not a;
    outputs(2567) <= b and not a;
    outputs(2568) <= a and b;
    outputs(2569) <= not a;
    outputs(2570) <= not (a or b);
    outputs(2571) <= not a;
    outputs(2572) <= a;
    outputs(2573) <= a xor b;
    outputs(2574) <= a;
    outputs(2575) <= not a or b;
    outputs(2576) <= not (a xor b);
    outputs(2577) <= not (a or b);
    outputs(2578) <= not (a and b);
    outputs(2579) <= not a;
    outputs(2580) <= a;
    outputs(2581) <= not (a xor b);
    outputs(2582) <= a;
    outputs(2583) <= not (a xor b);
    outputs(2584) <= not b;
    outputs(2585) <= not (a xor b);
    outputs(2586) <= not (a xor b);
    outputs(2587) <= a xor b;
    outputs(2588) <= not b;
    outputs(2589) <= a or b;
    outputs(2590) <= b;
    outputs(2591) <= b;
    outputs(2592) <= not b;
    outputs(2593) <= b;
    outputs(2594) <= not (a and b);
    outputs(2595) <= not b;
    outputs(2596) <= a and not b;
    outputs(2597) <= not (a xor b);
    outputs(2598) <= not b;
    outputs(2599) <= not (a and b);
    outputs(2600) <= a;
    outputs(2601) <= not b;
    outputs(2602) <= a;
    outputs(2603) <= not a;
    outputs(2604) <= a and b;
    outputs(2605) <= a xor b;
    outputs(2606) <= a;
    outputs(2607) <= not b or a;
    outputs(2608) <= a xor b;
    outputs(2609) <= not (a xor b);
    outputs(2610) <= a xor b;
    outputs(2611) <= a;
    outputs(2612) <= not b;
    outputs(2613) <= not b;
    outputs(2614) <= a xor b;
    outputs(2615) <= not (a xor b);
    outputs(2616) <= not a or b;
    outputs(2617) <= not (a xor b);
    outputs(2618) <= a;
    outputs(2619) <= not b;
    outputs(2620) <= not a;
    outputs(2621) <= not b;
    outputs(2622) <= not (a xor b);
    outputs(2623) <= not (a xor b);
    outputs(2624) <= b;
    outputs(2625) <= b and not a;
    outputs(2626) <= b;
    outputs(2627) <= not (a or b);
    outputs(2628) <= not (a xor b);
    outputs(2629) <= a and not b;
    outputs(2630) <= not (a xor b);
    outputs(2631) <= not (a xor b);
    outputs(2632) <= not (a xor b);
    outputs(2633) <= not (a or b);
    outputs(2634) <= a;
    outputs(2635) <= a;
    outputs(2636) <= not a;
    outputs(2637) <= a or b;
    outputs(2638) <= a xor b;
    outputs(2639) <= not (a xor b);
    outputs(2640) <= not a;
    outputs(2641) <= b;
    outputs(2642) <= not a;
    outputs(2643) <= a and not b;
    outputs(2644) <= not b;
    outputs(2645) <= not (a xor b);
    outputs(2646) <= not b;
    outputs(2647) <= a xor b;
    outputs(2648) <= not b;
    outputs(2649) <= a and not b;
    outputs(2650) <= not (a xor b);
    outputs(2651) <= a;
    outputs(2652) <= a and not b;
    outputs(2653) <= not a;
    outputs(2654) <= not a;
    outputs(2655) <= not a;
    outputs(2656) <= b and not a;
    outputs(2657) <= not a;
    outputs(2658) <= a;
    outputs(2659) <= not (a xor b);
    outputs(2660) <= not (a xor b);
    outputs(2661) <= not (a or b);
    outputs(2662) <= b;
    outputs(2663) <= b;
    outputs(2664) <= not (a xor b);
    outputs(2665) <= a;
    outputs(2666) <= b;
    outputs(2667) <= a and b;
    outputs(2668) <= b;
    outputs(2669) <= b;
    outputs(2670) <= b;
    outputs(2671) <= a xor b;
    outputs(2672) <= a xor b;
    outputs(2673) <= not a;
    outputs(2674) <= not a;
    outputs(2675) <= a;
    outputs(2676) <= a and b;
    outputs(2677) <= b;
    outputs(2678) <= not (a xor b);
    outputs(2679) <= not (a xor b);
    outputs(2680) <= b;
    outputs(2681) <= a xor b;
    outputs(2682) <= a;
    outputs(2683) <= b;
    outputs(2684) <= b and not a;
    outputs(2685) <= not a or b;
    outputs(2686) <= b;
    outputs(2687) <= a xor b;
    outputs(2688) <= a;
    outputs(2689) <= b and not a;
    outputs(2690) <= a;
    outputs(2691) <= not a;
    outputs(2692) <= not (a or b);
    outputs(2693) <= a xor b;
    outputs(2694) <= not (a xor b);
    outputs(2695) <= b;
    outputs(2696) <= a or b;
    outputs(2697) <= a and b;
    outputs(2698) <= a and b;
    outputs(2699) <= not a;
    outputs(2700) <= a;
    outputs(2701) <= not b;
    outputs(2702) <= a;
    outputs(2703) <= not (a xor b);
    outputs(2704) <= not (a xor b);
    outputs(2705) <= a;
    outputs(2706) <= b;
    outputs(2707) <= a;
    outputs(2708) <= a;
    outputs(2709) <= not b;
    outputs(2710) <= a xor b;
    outputs(2711) <= not (a and b);
    outputs(2712) <= not (a xor b);
    outputs(2713) <= b;
    outputs(2714) <= b and not a;
    outputs(2715) <= not b;
    outputs(2716) <= a xor b;
    outputs(2717) <= not (a xor b);
    outputs(2718) <= a xor b;
    outputs(2719) <= b and not a;
    outputs(2720) <= a xor b;
    outputs(2721) <= b;
    outputs(2722) <= not (a xor b);
    outputs(2723) <= not b;
    outputs(2724) <= not b;
    outputs(2725) <= not a;
    outputs(2726) <= not (a xor b);
    outputs(2727) <= not a;
    outputs(2728) <= a xor b;
    outputs(2729) <= not b;
    outputs(2730) <= a and b;
    outputs(2731) <= a;
    outputs(2732) <= not b;
    outputs(2733) <= a;
    outputs(2734) <= not a;
    outputs(2735) <= not b;
    outputs(2736) <= a;
    outputs(2737) <= not b;
    outputs(2738) <= a xor b;
    outputs(2739) <= not a;
    outputs(2740) <= a xor b;
    outputs(2741) <= not b;
    outputs(2742) <= not a;
    outputs(2743) <= not a or b;
    outputs(2744) <= not (a xor b);
    outputs(2745) <= not (a xor b);
    outputs(2746) <= not b;
    outputs(2747) <= a xor b;
    outputs(2748) <= not a;
    outputs(2749) <= not a;
    outputs(2750) <= not (a xor b);
    outputs(2751) <= not (a xor b);
    outputs(2752) <= not (a xor b);
    outputs(2753) <= a and b;
    outputs(2754) <= b;
    outputs(2755) <= not (a xor b);
    outputs(2756) <= not (a xor b);
    outputs(2757) <= not (a xor b);
    outputs(2758) <= b and not a;
    outputs(2759) <= not (a xor b);
    outputs(2760) <= not a;
    outputs(2761) <= b and not a;
    outputs(2762) <= a and b;
    outputs(2763) <= not (a xor b);
    outputs(2764) <= b and not a;
    outputs(2765) <= a;
    outputs(2766) <= a and not b;
    outputs(2767) <= a;
    outputs(2768) <= a;
    outputs(2769) <= not (a xor b);
    outputs(2770) <= a;
    outputs(2771) <= not a;
    outputs(2772) <= not (a xor b);
    outputs(2773) <= not (a xor b);
    outputs(2774) <= not b;
    outputs(2775) <= a and b;
    outputs(2776) <= a xor b;
    outputs(2777) <= not (a xor b);
    outputs(2778) <= b;
    outputs(2779) <= not (a xor b);
    outputs(2780) <= a and not b;
    outputs(2781) <= not (a xor b);
    outputs(2782) <= b and not a;
    outputs(2783) <= a and not b;
    outputs(2784) <= not (a xor b);
    outputs(2785) <= not (a or b);
    outputs(2786) <= a xor b;
    outputs(2787) <= b;
    outputs(2788) <= not (a xor b);
    outputs(2789) <= a and b;
    outputs(2790) <= a and b;
    outputs(2791) <= a and b;
    outputs(2792) <= a;
    outputs(2793) <= not b;
    outputs(2794) <= not a;
    outputs(2795) <= not b;
    outputs(2796) <= not a or b;
    outputs(2797) <= not a;
    outputs(2798) <= b;
    outputs(2799) <= not a;
    outputs(2800) <= a xor b;
    outputs(2801) <= not a;
    outputs(2802) <= not (a xor b);
    outputs(2803) <= a and not b;
    outputs(2804) <= b;
    outputs(2805) <= not a or b;
    outputs(2806) <= not b;
    outputs(2807) <= a xor b;
    outputs(2808) <= not b;
    outputs(2809) <= a;
    outputs(2810) <= a and b;
    outputs(2811) <= not b;
    outputs(2812) <= a;
    outputs(2813) <= a;
    outputs(2814) <= a;
    outputs(2815) <= b and not a;
    outputs(2816) <= a;
    outputs(2817) <= not b;
    outputs(2818) <= not a or b;
    outputs(2819) <= a xor b;
    outputs(2820) <= a;
    outputs(2821) <= not (a xor b);
    outputs(2822) <= not b;
    outputs(2823) <= a;
    outputs(2824) <= a xor b;
    outputs(2825) <= not (a xor b);
    outputs(2826) <= not (a xor b);
    outputs(2827) <= a xor b;
    outputs(2828) <= a xor b;
    outputs(2829) <= not b;
    outputs(2830) <= a xor b;
    outputs(2831) <= a xor b;
    outputs(2832) <= not a or b;
    outputs(2833) <= a and b;
    outputs(2834) <= a xor b;
    outputs(2835) <= not (a xor b);
    outputs(2836) <= not b;
    outputs(2837) <= a and not b;
    outputs(2838) <= a xor b;
    outputs(2839) <= not (a and b);
    outputs(2840) <= not (a and b);
    outputs(2841) <= not (a xor b);
    outputs(2842) <= b;
    outputs(2843) <= a and not b;
    outputs(2844) <= not (a xor b);
    outputs(2845) <= a;
    outputs(2846) <= a and not b;
    outputs(2847) <= not a;
    outputs(2848) <= not (a xor b);
    outputs(2849) <= not (a xor b);
    outputs(2850) <= not (a xor b);
    outputs(2851) <= not a;
    outputs(2852) <= b;
    outputs(2853) <= not (a or b);
    outputs(2854) <= not a or b;
    outputs(2855) <= a;
    outputs(2856) <= a xor b;
    outputs(2857) <= not a;
    outputs(2858) <= not (a xor b);
    outputs(2859) <= not b;
    outputs(2860) <= not b;
    outputs(2861) <= a xor b;
    outputs(2862) <= not b or a;
    outputs(2863) <= b;
    outputs(2864) <= not (a and b);
    outputs(2865) <= a;
    outputs(2866) <= not b;
    outputs(2867) <= not b;
    outputs(2868) <= b;
    outputs(2869) <= not b;
    outputs(2870) <= a xor b;
    outputs(2871) <= not b;
    outputs(2872) <= b;
    outputs(2873) <= not a;
    outputs(2874) <= not (a or b);
    outputs(2875) <= b;
    outputs(2876) <= not a or b;
    outputs(2877) <= not a;
    outputs(2878) <= not (a or b);
    outputs(2879) <= a and b;
    outputs(2880) <= not (a or b);
    outputs(2881) <= not (a or b);
    outputs(2882) <= a and b;
    outputs(2883) <= not (a xor b);
    outputs(2884) <= a;
    outputs(2885) <= a and b;
    outputs(2886) <= not a;
    outputs(2887) <= a xor b;
    outputs(2888) <= not b or a;
    outputs(2889) <= a xor b;
    outputs(2890) <= not b;
    outputs(2891) <= not b;
    outputs(2892) <= a;
    outputs(2893) <= not a;
    outputs(2894) <= a xor b;
    outputs(2895) <= not b;
    outputs(2896) <= b;
    outputs(2897) <= b and not a;
    outputs(2898) <= a and not b;
    outputs(2899) <= not (a or b);
    outputs(2900) <= not a;
    outputs(2901) <= not (a xor b);
    outputs(2902) <= not (a xor b);
    outputs(2903) <= b;
    outputs(2904) <= not b;
    outputs(2905) <= not b;
    outputs(2906) <= a xor b;
    outputs(2907) <= a xor b;
    outputs(2908) <= not (a xor b);
    outputs(2909) <= not (a xor b);
    outputs(2910) <= not a;
    outputs(2911) <= b;
    outputs(2912) <= b and not a;
    outputs(2913) <= not a;
    outputs(2914) <= not b;
    outputs(2915) <= b and not a;
    outputs(2916) <= a and not b;
    outputs(2917) <= a;
    outputs(2918) <= not a;
    outputs(2919) <= a xor b;
    outputs(2920) <= not a;
    outputs(2921) <= b;
    outputs(2922) <= not b;
    outputs(2923) <= a xor b;
    outputs(2924) <= not (a xor b);
    outputs(2925) <= not (a or b);
    outputs(2926) <= b;
    outputs(2927) <= not b;
    outputs(2928) <= not (a xor b);
    outputs(2929) <= b and not a;
    outputs(2930) <= a and b;
    outputs(2931) <= not (a xor b);
    outputs(2932) <= not a;
    outputs(2933) <= not (a xor b);
    outputs(2934) <= not a;
    outputs(2935) <= not (a xor b);
    outputs(2936) <= not b;
    outputs(2937) <= a xor b;
    outputs(2938) <= a;
    outputs(2939) <= a xor b;
    outputs(2940) <= b;
    outputs(2941) <= not a;
    outputs(2942) <= not b;
    outputs(2943) <= b;
    outputs(2944) <= a xor b;
    outputs(2945) <= not (a xor b);
    outputs(2946) <= b;
    outputs(2947) <= a;
    outputs(2948) <= not b;
    outputs(2949) <= not (a xor b);
    outputs(2950) <= not a;
    outputs(2951) <= not (a xor b);
    outputs(2952) <= not (a xor b);
    outputs(2953) <= not (a xor b);
    outputs(2954) <= not (a xor b);
    outputs(2955) <= b and not a;
    outputs(2956) <= a xor b;
    outputs(2957) <= a xor b;
    outputs(2958) <= not (a xor b);
    outputs(2959) <= a xor b;
    outputs(2960) <= not (a xor b);
    outputs(2961) <= not b;
    outputs(2962) <= a xor b;
    outputs(2963) <= a and b;
    outputs(2964) <= not (a and b);
    outputs(2965) <= not a;
    outputs(2966) <= not (a xor b);
    outputs(2967) <= a;
    outputs(2968) <= not b;
    outputs(2969) <= b;
    outputs(2970) <= not (a xor b);
    outputs(2971) <= a xor b;
    outputs(2972) <= not a;
    outputs(2973) <= a and not b;
    outputs(2974) <= b and not a;
    outputs(2975) <= a and not b;
    outputs(2976) <= not (a xor b);
    outputs(2977) <= not (a or b);
    outputs(2978) <= b and not a;
    outputs(2979) <= a and b;
    outputs(2980) <= a xor b;
    outputs(2981) <= b;
    outputs(2982) <= not a;
    outputs(2983) <= b;
    outputs(2984) <= not (a xor b);
    outputs(2985) <= not (a and b);
    outputs(2986) <= not b;
    outputs(2987) <= not (a or b);
    outputs(2988) <= not a or b;
    outputs(2989) <= a xor b;
    outputs(2990) <= b and not a;
    outputs(2991) <= b and not a;
    outputs(2992) <= not b;
    outputs(2993) <= a or b;
    outputs(2994) <= not a or b;
    outputs(2995) <= not a;
    outputs(2996) <= a;
    outputs(2997) <= not a;
    outputs(2998) <= a;
    outputs(2999) <= not b;
    outputs(3000) <= a xor b;
    outputs(3001) <= not a;
    outputs(3002) <= b;
    outputs(3003) <= a xor b;
    outputs(3004) <= a or b;
    outputs(3005) <= not b;
    outputs(3006) <= not (a xor b);
    outputs(3007) <= not (a or b);
    outputs(3008) <= b;
    outputs(3009) <= not (a or b);
    outputs(3010) <= a;
    outputs(3011) <= a xor b;
    outputs(3012) <= a xor b;
    outputs(3013) <= not b;
    outputs(3014) <= not b;
    outputs(3015) <= a xor b;
    outputs(3016) <= a xor b;
    outputs(3017) <= not b;
    outputs(3018) <= a xor b;
    outputs(3019) <= not (a or b);
    outputs(3020) <= not (a xor b);
    outputs(3021) <= not a;
    outputs(3022) <= not a or b;
    outputs(3023) <= not b;
    outputs(3024) <= not a;
    outputs(3025) <= a and not b;
    outputs(3026) <= not a or b;
    outputs(3027) <= a and b;
    outputs(3028) <= not (a or b);
    outputs(3029) <= a xor b;
    outputs(3030) <= not a;
    outputs(3031) <= a xor b;
    outputs(3032) <= a xor b;
    outputs(3033) <= a and not b;
    outputs(3034) <= b;
    outputs(3035) <= a xor b;
    outputs(3036) <= not (a xor b);
    outputs(3037) <= a xor b;
    outputs(3038) <= a;
    outputs(3039) <= a;
    outputs(3040) <= a;
    outputs(3041) <= a and b;
    outputs(3042) <= not (a xor b);
    outputs(3043) <= a;
    outputs(3044) <= a and not b;
    outputs(3045) <= a xor b;
    outputs(3046) <= a and b;
    outputs(3047) <= not a;
    outputs(3048) <= a;
    outputs(3049) <= not b or a;
    outputs(3050) <= b;
    outputs(3051) <= not (a xor b);
    outputs(3052) <= not b;
    outputs(3053) <= not a;
    outputs(3054) <= b and not a;
    outputs(3055) <= not b or a;
    outputs(3056) <= a and b;
    outputs(3057) <= b;
    outputs(3058) <= a xor b;
    outputs(3059) <= not (a xor b);
    outputs(3060) <= not b or a;
    outputs(3061) <= b;
    outputs(3062) <= not (a xor b);
    outputs(3063) <= not (a or b);
    outputs(3064) <= a;
    outputs(3065) <= not (a xor b);
    outputs(3066) <= b and not a;
    outputs(3067) <= not (a or b);
    outputs(3068) <= not b;
    outputs(3069) <= not b;
    outputs(3070) <= a and not b;
    outputs(3071) <= not b;
    outputs(3072) <= not (a or b);
    outputs(3073) <= a xor b;
    outputs(3074) <= not a or b;
    outputs(3075) <= a xor b;
    outputs(3076) <= a or b;
    outputs(3077) <= a;
    outputs(3078) <= a xor b;
    outputs(3079) <= a or b;
    outputs(3080) <= not a;
    outputs(3081) <= a;
    outputs(3082) <= not (a xor b);
    outputs(3083) <= not a;
    outputs(3084) <= a and b;
    outputs(3085) <= not a;
    outputs(3086) <= a xor b;
    outputs(3087) <= not b;
    outputs(3088) <= a or b;
    outputs(3089) <= not b;
    outputs(3090) <= not (a xor b);
    outputs(3091) <= a and not b;
    outputs(3092) <= a;
    outputs(3093) <= b and not a;
    outputs(3094) <= not (a or b);
    outputs(3095) <= not a;
    outputs(3096) <= not a;
    outputs(3097) <= not a;
    outputs(3098) <= a;
    outputs(3099) <= b;
    outputs(3100) <= not a or b;
    outputs(3101) <= not (a xor b);
    outputs(3102) <= not a;
    outputs(3103) <= not b;
    outputs(3104) <= not b;
    outputs(3105) <= not (a xor b);
    outputs(3106) <= a xor b;
    outputs(3107) <= not a;
    outputs(3108) <= not a or b;
    outputs(3109) <= not (a or b);
    outputs(3110) <= a and not b;
    outputs(3111) <= not (a xor b);
    outputs(3112) <= a xor b;
    outputs(3113) <= a;
    outputs(3114) <= a xor b;
    outputs(3115) <= b and not a;
    outputs(3116) <= not (a and b);
    outputs(3117) <= a;
    outputs(3118) <= not a or b;
    outputs(3119) <= not b;
    outputs(3120) <= not (a or b);
    outputs(3121) <= a or b;
    outputs(3122) <= b;
    outputs(3123) <= b;
    outputs(3124) <= a and not b;
    outputs(3125) <= b;
    outputs(3126) <= a;
    outputs(3127) <= not (a xor b);
    outputs(3128) <= not a;
    outputs(3129) <= b and not a;
    outputs(3130) <= a;
    outputs(3131) <= b;
    outputs(3132) <= not b;
    outputs(3133) <= a or b;
    outputs(3134) <= not b;
    outputs(3135) <= not a;
    outputs(3136) <= not (a or b);
    outputs(3137) <= not (a and b);
    outputs(3138) <= not a;
    outputs(3139) <= not a;
    outputs(3140) <= not b;
    outputs(3141) <= not a;
    outputs(3142) <= a and not b;
    outputs(3143) <= a xor b;
    outputs(3144) <= not b;
    outputs(3145) <= a;
    outputs(3146) <= b and not a;
    outputs(3147) <= a xor b;
    outputs(3148) <= not b;
    outputs(3149) <= not a;
    outputs(3150) <= not (a xor b);
    outputs(3151) <= not (a xor b);
    outputs(3152) <= a and not b;
    outputs(3153) <= a;
    outputs(3154) <= not a;
    outputs(3155) <= not a;
    outputs(3156) <= not (a or b);
    outputs(3157) <= b;
    outputs(3158) <= not a;
    outputs(3159) <= not (a xor b);
    outputs(3160) <= a xor b;
    outputs(3161) <= not (a xor b);
    outputs(3162) <= not a;
    outputs(3163) <= a or b;
    outputs(3164) <= not (a xor b);
    outputs(3165) <= a;
    outputs(3166) <= not b;
    outputs(3167) <= not a;
    outputs(3168) <= not a;
    outputs(3169) <= not b or a;
    outputs(3170) <= not (a xor b);
    outputs(3171) <= not a or b;
    outputs(3172) <= a;
    outputs(3173) <= not b;
    outputs(3174) <= a xor b;
    outputs(3175) <= a or b;
    outputs(3176) <= not b;
    outputs(3177) <= not b;
    outputs(3178) <= a;
    outputs(3179) <= a;
    outputs(3180) <= b;
    outputs(3181) <= a;
    outputs(3182) <= not b;
    outputs(3183) <= not (a and b);
    outputs(3184) <= not a;
    outputs(3185) <= a;
    outputs(3186) <= a xor b;
    outputs(3187) <= not (a and b);
    outputs(3188) <= a;
    outputs(3189) <= not (a and b);
    outputs(3190) <= a or b;
    outputs(3191) <= a xor b;
    outputs(3192) <= b;
    outputs(3193) <= b;
    outputs(3194) <= not b;
    outputs(3195) <= not b;
    outputs(3196) <= b;
    outputs(3197) <= b;
    outputs(3198) <= not (a and b);
    outputs(3199) <= not a;
    outputs(3200) <= b;
    outputs(3201) <= a;
    outputs(3202) <= not b;
    outputs(3203) <= a;
    outputs(3204) <= a;
    outputs(3205) <= not a;
    outputs(3206) <= not (a xor b);
    outputs(3207) <= b and not a;
    outputs(3208) <= a xor b;
    outputs(3209) <= not (a xor b);
    outputs(3210) <= not (a xor b);
    outputs(3211) <= not (a xor b);
    outputs(3212) <= a;
    outputs(3213) <= a or b;
    outputs(3214) <= a and b;
    outputs(3215) <= not (a xor b);
    outputs(3216) <= a xor b;
    outputs(3217) <= not b;
    outputs(3218) <= not a;
    outputs(3219) <= b;
    outputs(3220) <= not (a xor b);
    outputs(3221) <= a xor b;
    outputs(3222) <= not (a xor b);
    outputs(3223) <= not b or a;
    outputs(3224) <= b;
    outputs(3225) <= a and b;
    outputs(3226) <= not (a xor b);
    outputs(3227) <= not (a xor b);
    outputs(3228) <= not (a xor b);
    outputs(3229) <= not a;
    outputs(3230) <= a xor b;
    outputs(3231) <= not (a xor b);
    outputs(3232) <= not b;
    outputs(3233) <= a;
    outputs(3234) <= a xor b;
    outputs(3235) <= a xor b;
    outputs(3236) <= a or b;
    outputs(3237) <= not b;
    outputs(3238) <= not a;
    outputs(3239) <= b;
    outputs(3240) <= not a;
    outputs(3241) <= a and b;
    outputs(3242) <= not (a or b);
    outputs(3243) <= not (a xor b);
    outputs(3244) <= not (a xor b);
    outputs(3245) <= a xor b;
    outputs(3246) <= not a or b;
    outputs(3247) <= a xor b;
    outputs(3248) <= a;
    outputs(3249) <= not b;
    outputs(3250) <= a;
    outputs(3251) <= not a;
    outputs(3252) <= a or b;
    outputs(3253) <= not (a or b);
    outputs(3254) <= a xor b;
    outputs(3255) <= not (a xor b);
    outputs(3256) <= a and b;
    outputs(3257) <= a xor b;
    outputs(3258) <= a xor b;
    outputs(3259) <= a;
    outputs(3260) <= a;
    outputs(3261) <= a and b;
    outputs(3262) <= b;
    outputs(3263) <= b;
    outputs(3264) <= not a;
    outputs(3265) <= not b;
    outputs(3266) <= not a or b;
    outputs(3267) <= not b;
    outputs(3268) <= not a;
    outputs(3269) <= a;
    outputs(3270) <= not a;
    outputs(3271) <= not (a xor b);
    outputs(3272) <= a;
    outputs(3273) <= b and not a;
    outputs(3274) <= not a;
    outputs(3275) <= not (a xor b);
    outputs(3276) <= not a or b;
    outputs(3277) <= not (a xor b);
    outputs(3278) <= not (a xor b);
    outputs(3279) <= a;
    outputs(3280) <= b;
    outputs(3281) <= a and b;
    outputs(3282) <= not (a xor b);
    outputs(3283) <= not a;
    outputs(3284) <= a and b;
    outputs(3285) <= not (a xor b);
    outputs(3286) <= b;
    outputs(3287) <= b;
    outputs(3288) <= not a;
    outputs(3289) <= a xor b;
    outputs(3290) <= b;
    outputs(3291) <= not a;
    outputs(3292) <= not a;
    outputs(3293) <= not a;
    outputs(3294) <= a and not b;
    outputs(3295) <= b and not a;
    outputs(3296) <= b;
    outputs(3297) <= not (a or b);
    outputs(3298) <= not (a xor b);
    outputs(3299) <= a and not b;
    outputs(3300) <= a xor b;
    outputs(3301) <= not (a xor b);
    outputs(3302) <= a;
    outputs(3303) <= not b;
    outputs(3304) <= not a or b;
    outputs(3305) <= b;
    outputs(3306) <= b;
    outputs(3307) <= not a or b;
    outputs(3308) <= a;
    outputs(3309) <= not a;
    outputs(3310) <= not a or b;
    outputs(3311) <= not a or b;
    outputs(3312) <= not (a xor b);
    outputs(3313) <= a;
    outputs(3314) <= not b;
    outputs(3315) <= a xor b;
    outputs(3316) <= not b;
    outputs(3317) <= b and not a;
    outputs(3318) <= not (a xor b);
    outputs(3319) <= not (a xor b);
    outputs(3320) <= not (a xor b);
    outputs(3321) <= not a;
    outputs(3322) <= not a;
    outputs(3323) <= not a;
    outputs(3324) <= not a;
    outputs(3325) <= a;
    outputs(3326) <= a xor b;
    outputs(3327) <= not a;
    outputs(3328) <= b and not a;
    outputs(3329) <= not b;
    outputs(3330) <= a;
    outputs(3331) <= a xor b;
    outputs(3332) <= not b;
    outputs(3333) <= a xor b;
    outputs(3334) <= a and not b;
    outputs(3335) <= a or b;
    outputs(3336) <= not (a xor b);
    outputs(3337) <= not (a and b);
    outputs(3338) <= not (a or b);
    outputs(3339) <= a xor b;
    outputs(3340) <= b;
    outputs(3341) <= a;
    outputs(3342) <= not a;
    outputs(3343) <= a and not b;
    outputs(3344) <= a or b;
    outputs(3345) <= b;
    outputs(3346) <= not (a xor b);
    outputs(3347) <= a and b;
    outputs(3348) <= b and not a;
    outputs(3349) <= not (a or b);
    outputs(3350) <= a xor b;
    outputs(3351) <= not b;
    outputs(3352) <= a and b;
    outputs(3353) <= b;
    outputs(3354) <= a and b;
    outputs(3355) <= not a;
    outputs(3356) <= not (a xor b);
    outputs(3357) <= not b or a;
    outputs(3358) <= a;
    outputs(3359) <= not a;
    outputs(3360) <= not b;
    outputs(3361) <= a;
    outputs(3362) <= not b;
    outputs(3363) <= a;
    outputs(3364) <= not (a or b);
    outputs(3365) <= not (a xor b);
    outputs(3366) <= not a;
    outputs(3367) <= b;
    outputs(3368) <= not (a xor b);
    outputs(3369) <= b;
    outputs(3370) <= b;
    outputs(3371) <= a or b;
    outputs(3372) <= a and b;
    outputs(3373) <= not a;
    outputs(3374) <= a;
    outputs(3375) <= not b;
    outputs(3376) <= a;
    outputs(3377) <= not (a xor b);
    outputs(3378) <= b;
    outputs(3379) <= b and not a;
    outputs(3380) <= not a;
    outputs(3381) <= b;
    outputs(3382) <= a and not b;
    outputs(3383) <= b;
    outputs(3384) <= b;
    outputs(3385) <= b and not a;
    outputs(3386) <= a;
    outputs(3387) <= a;
    outputs(3388) <= b;
    outputs(3389) <= a xor b;
    outputs(3390) <= b;
    outputs(3391) <= b;
    outputs(3392) <= b;
    outputs(3393) <= not b;
    outputs(3394) <= not b;
    outputs(3395) <= not a;
    outputs(3396) <= not b or a;
    outputs(3397) <= a xor b;
    outputs(3398) <= not b;
    outputs(3399) <= not a;
    outputs(3400) <= not (a and b);
    outputs(3401) <= b;
    outputs(3402) <= a xor b;
    outputs(3403) <= a and not b;
    outputs(3404) <= not (a xor b);
    outputs(3405) <= not (a xor b);
    outputs(3406) <= not (a xor b);
    outputs(3407) <= a;
    outputs(3408) <= not (a xor b);
    outputs(3409) <= a and not b;
    outputs(3410) <= b;
    outputs(3411) <= a and not b;
    outputs(3412) <= a and b;
    outputs(3413) <= a and b;
    outputs(3414) <= b and not a;
    outputs(3415) <= a xor b;
    outputs(3416) <= not (a xor b);
    outputs(3417) <= not (a or b);
    outputs(3418) <= a and not b;
    outputs(3419) <= b;
    outputs(3420) <= not b;
    outputs(3421) <= a and b;
    outputs(3422) <= not (a xor b);
    outputs(3423) <= not b;
    outputs(3424) <= b;
    outputs(3425) <= not a;
    outputs(3426) <= a xor b;
    outputs(3427) <= a;
    outputs(3428) <= not b;
    outputs(3429) <= not (a xor b);
    outputs(3430) <= a and not b;
    outputs(3431) <= not b;
    outputs(3432) <= not a;
    outputs(3433) <= b;
    outputs(3434) <= not (a and b);
    outputs(3435) <= not a;
    outputs(3436) <= b;
    outputs(3437) <= not a;
    outputs(3438) <= not (a xor b);
    outputs(3439) <= not (a or b);
    outputs(3440) <= not a or b;
    outputs(3441) <= not b or a;
    outputs(3442) <= b and not a;
    outputs(3443) <= not b;
    outputs(3444) <= a;
    outputs(3445) <= b and not a;
    outputs(3446) <= a;
    outputs(3447) <= b;
    outputs(3448) <= b;
    outputs(3449) <= a;
    outputs(3450) <= not b;
    outputs(3451) <= a;
    outputs(3452) <= not b;
    outputs(3453) <= a;
    outputs(3454) <= not b;
    outputs(3455) <= not a;
    outputs(3456) <= not b;
    outputs(3457) <= b;
    outputs(3458) <= not a;
    outputs(3459) <= a and b;
    outputs(3460) <= not (a xor b);
    outputs(3461) <= not (a xor b);
    outputs(3462) <= a xor b;
    outputs(3463) <= not (a xor b);
    outputs(3464) <= a xor b;
    outputs(3465) <= a xor b;
    outputs(3466) <= not b;
    outputs(3467) <= b;
    outputs(3468) <= a;
    outputs(3469) <= not a or b;
    outputs(3470) <= a;
    outputs(3471) <= not b or a;
    outputs(3472) <= a xor b;
    outputs(3473) <= not b;
    outputs(3474) <= not a;
    outputs(3475) <= b;
    outputs(3476) <= a and b;
    outputs(3477) <= a and b;
    outputs(3478) <= b;
    outputs(3479) <= not a;
    outputs(3480) <= a and not b;
    outputs(3481) <= a;
    outputs(3482) <= a;
    outputs(3483) <= a;
    outputs(3484) <= not b;
    outputs(3485) <= not a;
    outputs(3486) <= not b;
    outputs(3487) <= not b;
    outputs(3488) <= a xor b;
    outputs(3489) <= not (a or b);
    outputs(3490) <= not (a xor b);
    outputs(3491) <= not b;
    outputs(3492) <= not (a xor b);
    outputs(3493) <= not (a and b);
    outputs(3494) <= not b;
    outputs(3495) <= a;
    outputs(3496) <= b;
    outputs(3497) <= a xor b;
    outputs(3498) <= a;
    outputs(3499) <= not (a xor b);
    outputs(3500) <= a;
    outputs(3501) <= not (a or b);
    outputs(3502) <= not (a and b);
    outputs(3503) <= a and b;
    outputs(3504) <= a and b;
    outputs(3505) <= a;
    outputs(3506) <= not (a or b);
    outputs(3507) <= not b;
    outputs(3508) <= not (a xor b);
    outputs(3509) <= not b;
    outputs(3510) <= a xor b;
    outputs(3511) <= not (a and b);
    outputs(3512) <= b and not a;
    outputs(3513) <= not a;
    outputs(3514) <= not b;
    outputs(3515) <= a xor b;
    outputs(3516) <= b;
    outputs(3517) <= a xor b;
    outputs(3518) <= not a or b;
    outputs(3519) <= a;
    outputs(3520) <= not (a xor b);
    outputs(3521) <= not (a xor b);
    outputs(3522) <= a;
    outputs(3523) <= not (a or b);
    outputs(3524) <= not (a xor b);
    outputs(3525) <= not b;
    outputs(3526) <= b;
    outputs(3527) <= a;
    outputs(3528) <= not (a and b);
    outputs(3529) <= a and not b;
    outputs(3530) <= not (a xor b);
    outputs(3531) <= not b;
    outputs(3532) <= not a;
    outputs(3533) <= a;
    outputs(3534) <= not (a xor b);
    outputs(3535) <= a;
    outputs(3536) <= a;
    outputs(3537) <= b;
    outputs(3538) <= not (a and b);
    outputs(3539) <= not b;
    outputs(3540) <= a and b;
    outputs(3541) <= b;
    outputs(3542) <= b;
    outputs(3543) <= not (a or b);
    outputs(3544) <= not (a xor b);
    outputs(3545) <= a and not b;
    outputs(3546) <= not (a and b);
    outputs(3547) <= b;
    outputs(3548) <= not (a and b);
    outputs(3549) <= not b;
    outputs(3550) <= a xor b;
    outputs(3551) <= not (a xor b);
    outputs(3552) <= a;
    outputs(3553) <= a xor b;
    outputs(3554) <= not (a xor b);
    outputs(3555) <= not b or a;
    outputs(3556) <= a xor b;
    outputs(3557) <= not (a or b);
    outputs(3558) <= not b;
    outputs(3559) <= a or b;
    outputs(3560) <= a xor b;
    outputs(3561) <= a;
    outputs(3562) <= a and not b;
    outputs(3563) <= not (a xor b);
    outputs(3564) <= a and not b;
    outputs(3565) <= not (a or b);
    outputs(3566) <= a xor b;
    outputs(3567) <= not b;
    outputs(3568) <= not (a xor b);
    outputs(3569) <= not a;
    outputs(3570) <= not b or a;
    outputs(3571) <= a and not b;
    outputs(3572) <= not b;
    outputs(3573) <= a and not b;
    outputs(3574) <= not b;
    outputs(3575) <= a;
    outputs(3576) <= b;
    outputs(3577) <= b;
    outputs(3578) <= a xor b;
    outputs(3579) <= not a;
    outputs(3580) <= not (a xor b);
    outputs(3581) <= not a;
    outputs(3582) <= not a or b;
    outputs(3583) <= not (a xor b);
    outputs(3584) <= not a;
    outputs(3585) <= a and not b;
    outputs(3586) <= not (a or b);
    outputs(3587) <= not b;
    outputs(3588) <= not b or a;
    outputs(3589) <= not (a xor b);
    outputs(3590) <= a;
    outputs(3591) <= a xor b;
    outputs(3592) <= a xor b;
    outputs(3593) <= a and not b;
    outputs(3594) <= a and not b;
    outputs(3595) <= a;
    outputs(3596) <= not a;
    outputs(3597) <= b;
    outputs(3598) <= a and b;
    outputs(3599) <= a and b;
    outputs(3600) <= not a or b;
    outputs(3601) <= not b;
    outputs(3602) <= a and b;
    outputs(3603) <= a or b;
    outputs(3604) <= not a;
    outputs(3605) <= not b;
    outputs(3606) <= a and not b;
    outputs(3607) <= not a;
    outputs(3608) <= b and not a;
    outputs(3609) <= not (a xor b);
    outputs(3610) <= b and not a;
    outputs(3611) <= a and not b;
    outputs(3612) <= a xor b;
    outputs(3613) <= not b;
    outputs(3614) <= a and not b;
    outputs(3615) <= not a;
    outputs(3616) <= not (a and b);
    outputs(3617) <= not (a xor b);
    outputs(3618) <= not (a or b);
    outputs(3619) <= a and not b;
    outputs(3620) <= a and b;
    outputs(3621) <= a;
    outputs(3622) <= not (a xor b);
    outputs(3623) <= a;
    outputs(3624) <= not (a xor b);
    outputs(3625) <= a and not b;
    outputs(3626) <= a xor b;
    outputs(3627) <= not a;
    outputs(3628) <= not (a xor b);
    outputs(3629) <= a xor b;
    outputs(3630) <= a or b;
    outputs(3631) <= a xor b;
    outputs(3632) <= a and b;
    outputs(3633) <= a xor b;
    outputs(3634) <= not b;
    outputs(3635) <= a xor b;
    outputs(3636) <= b;
    outputs(3637) <= not (a xor b);
    outputs(3638) <= b and not a;
    outputs(3639) <= not b;
    outputs(3640) <= not (a xor b);
    outputs(3641) <= a and b;
    outputs(3642) <= not b or a;
    outputs(3643) <= a;
    outputs(3644) <= a xor b;
    outputs(3645) <= b;
    outputs(3646) <= b;
    outputs(3647) <= not b;
    outputs(3648) <= not b;
    outputs(3649) <= not (a xor b);
    outputs(3650) <= a and not b;
    outputs(3651) <= a;
    outputs(3652) <= not b;
    outputs(3653) <= not b;
    outputs(3654) <= a;
    outputs(3655) <= b;
    outputs(3656) <= not b;
    outputs(3657) <= not b;
    outputs(3658) <= not a;
    outputs(3659) <= a and not b;
    outputs(3660) <= a xor b;
    outputs(3661) <= a and not b;
    outputs(3662) <= a xor b;
    outputs(3663) <= b;
    outputs(3664) <= b;
    outputs(3665) <= not (a or b);
    outputs(3666) <= not b;
    outputs(3667) <= not a;
    outputs(3668) <= a;
    outputs(3669) <= not a;
    outputs(3670) <= a and not b;
    outputs(3671) <= not b;
    outputs(3672) <= a;
    outputs(3673) <= b;
    outputs(3674) <= a and not b;
    outputs(3675) <= not b or a;
    outputs(3676) <= a xor b;
    outputs(3677) <= not (a xor b);
    outputs(3678) <= a xor b;
    outputs(3679) <= not a;
    outputs(3680) <= not b;
    outputs(3681) <= a;
    outputs(3682) <= a and not b;
    outputs(3683) <= a and not b;
    outputs(3684) <= not a or b;
    outputs(3685) <= not b;
    outputs(3686) <= not (a xor b);
    outputs(3687) <= not (a xor b);
    outputs(3688) <= b;
    outputs(3689) <= a;
    outputs(3690) <= not a or b;
    outputs(3691) <= a xor b;
    outputs(3692) <= not b;
    outputs(3693) <= b and not a;
    outputs(3694) <= not a;
    outputs(3695) <= not b;
    outputs(3696) <= not a;
    outputs(3697) <= not (a xor b);
    outputs(3698) <= b;
    outputs(3699) <= not a;
    outputs(3700) <= not a;
    outputs(3701) <= b and not a;
    outputs(3702) <= a xor b;
    outputs(3703) <= not b;
    outputs(3704) <= not a;
    outputs(3705) <= b;
    outputs(3706) <= not (a and b);
    outputs(3707) <= not b;
    outputs(3708) <= not (a or b);
    outputs(3709) <= a;
    outputs(3710) <= a or b;
    outputs(3711) <= a xor b;
    outputs(3712) <= not b;
    outputs(3713) <= not (a xor b);
    outputs(3714) <= a xor b;
    outputs(3715) <= a xor b;
    outputs(3716) <= not b;
    outputs(3717) <= a xor b;
    outputs(3718) <= not b;
    outputs(3719) <= not (a xor b);
    outputs(3720) <= a and b;
    outputs(3721) <= a xor b;
    outputs(3722) <= not a;
    outputs(3723) <= b;
    outputs(3724) <= a;
    outputs(3725) <= b;
    outputs(3726) <= b and not a;
    outputs(3727) <= not a;
    outputs(3728) <= b;
    outputs(3729) <= a and not b;
    outputs(3730) <= not (a xor b);
    outputs(3731) <= not a or b;
    outputs(3732) <= not a;
    outputs(3733) <= not a;
    outputs(3734) <= a;
    outputs(3735) <= a xor b;
    outputs(3736) <= not b;
    outputs(3737) <= not (a xor b);
    outputs(3738) <= b;
    outputs(3739) <= a;
    outputs(3740) <= not b;
    outputs(3741) <= b;
    outputs(3742) <= a xor b;
    outputs(3743) <= a xor b;
    outputs(3744) <= not (a and b);
    outputs(3745) <= b and not a;
    outputs(3746) <= a;
    outputs(3747) <= b;
    outputs(3748) <= not (a xor b);
    outputs(3749) <= a and b;
    outputs(3750) <= not (a or b);
    outputs(3751) <= b;
    outputs(3752) <= a or b;
    outputs(3753) <= not (a xor b);
    outputs(3754) <= not b or a;
    outputs(3755) <= a and b;
    outputs(3756) <= a;
    outputs(3757) <= not b or a;
    outputs(3758) <= not (a xor b);
    outputs(3759) <= a and not b;
    outputs(3760) <= b and not a;
    outputs(3761) <= a xor b;
    outputs(3762) <= b;
    outputs(3763) <= a;
    outputs(3764) <= a xor b;
    outputs(3765) <= not a;
    outputs(3766) <= not (a xor b);
    outputs(3767) <= a or b;
    outputs(3768) <= a xor b;
    outputs(3769) <= not a;
    outputs(3770) <= not (a or b);
    outputs(3771) <= not a;
    outputs(3772) <= b and not a;
    outputs(3773) <= b and not a;
    outputs(3774) <= not (a xor b);
    outputs(3775) <= not a;
    outputs(3776) <= not b;
    outputs(3777) <= b;
    outputs(3778) <= a xor b;
    outputs(3779) <= not (a xor b);
    outputs(3780) <= not b;
    outputs(3781) <= not b;
    outputs(3782) <= a xor b;
    outputs(3783) <= b;
    outputs(3784) <= a and b;
    outputs(3785) <= a xor b;
    outputs(3786) <= not a;
    outputs(3787) <= not a;
    outputs(3788) <= not (a and b);
    outputs(3789) <= a;
    outputs(3790) <= a;
    outputs(3791) <= a;
    outputs(3792) <= not a;
    outputs(3793) <= a xor b;
    outputs(3794) <= not b;
    outputs(3795) <= not (a and b);
    outputs(3796) <= not (a or b);
    outputs(3797) <= not (a xor b);
    outputs(3798) <= b;
    outputs(3799) <= not b;
    outputs(3800) <= a or b;
    outputs(3801) <= a and b;
    outputs(3802) <= not (a or b);
    outputs(3803) <= not a;
    outputs(3804) <= not a;
    outputs(3805) <= not (a xor b);
    outputs(3806) <= not b;
    outputs(3807) <= b;
    outputs(3808) <= a;
    outputs(3809) <= not (a or b);
    outputs(3810) <= a and not b;
    outputs(3811) <= not a;
    outputs(3812) <= a;
    outputs(3813) <= not b;
    outputs(3814) <= b and not a;
    outputs(3815) <= not (a or b);
    outputs(3816) <= a;
    outputs(3817) <= b;
    outputs(3818) <= b;
    outputs(3819) <= not b;
    outputs(3820) <= a and b;
    outputs(3821) <= a xor b;
    outputs(3822) <= not b or a;
    outputs(3823) <= a xor b;
    outputs(3824) <= not b;
    outputs(3825) <= a and b;
    outputs(3826) <= b;
    outputs(3827) <= not a;
    outputs(3828) <= a xor b;
    outputs(3829) <= not (a xor b);
    outputs(3830) <= not (a or b);
    outputs(3831) <= not b;
    outputs(3832) <= not (a xor b);
    outputs(3833) <= a xor b;
    outputs(3834) <= a xor b;
    outputs(3835) <= not b;
    outputs(3836) <= a;
    outputs(3837) <= not (a or b);
    outputs(3838) <= not a;
    outputs(3839) <= a;
    outputs(3840) <= not a;
    outputs(3841) <= not (a xor b);
    outputs(3842) <= a;
    outputs(3843) <= b;
    outputs(3844) <= a and b;
    outputs(3845) <= a and b;
    outputs(3846) <= not a;
    outputs(3847) <= a or b;
    outputs(3848) <= a and b;
    outputs(3849) <= a and b;
    outputs(3850) <= b;
    outputs(3851) <= not b;
    outputs(3852) <= a;
    outputs(3853) <= a and not b;
    outputs(3854) <= not b;
    outputs(3855) <= a and not b;
    outputs(3856) <= a;
    outputs(3857) <= not (a xor b);
    outputs(3858) <= b and not a;
    outputs(3859) <= a xor b;
    outputs(3860) <= a and not b;
    outputs(3861) <= not (a xor b);
    outputs(3862) <= not b or a;
    outputs(3863) <= a xor b;
    outputs(3864) <= not a;
    outputs(3865) <= not a;
    outputs(3866) <= b and not a;
    outputs(3867) <= b and not a;
    outputs(3868) <= a xor b;
    outputs(3869) <= not (a xor b);
    outputs(3870) <= b;
    outputs(3871) <= b and not a;
    outputs(3872) <= a and b;
    outputs(3873) <= a;
    outputs(3874) <= not b;
    outputs(3875) <= not a;
    outputs(3876) <= not (a xor b);
    outputs(3877) <= not (a or b);
    outputs(3878) <= not (a xor b);
    outputs(3879) <= a and not b;
    outputs(3880) <= not (a or b);
    outputs(3881) <= b;
    outputs(3882) <= a;
    outputs(3883) <= not a;
    outputs(3884) <= not (a xor b);
    outputs(3885) <= a or b;
    outputs(3886) <= a xor b;
    outputs(3887) <= a or b;
    outputs(3888) <= b;
    outputs(3889) <= not a;
    outputs(3890) <= a;
    outputs(3891) <= a;
    outputs(3892) <= not (a xor b);
    outputs(3893) <= b;
    outputs(3894) <= a;
    outputs(3895) <= b;
    outputs(3896) <= not (a xor b);
    outputs(3897) <= a and b;
    outputs(3898) <= a and not b;
    outputs(3899) <= not b;
    outputs(3900) <= b;
    outputs(3901) <= not (a and b);
    outputs(3902) <= not (a xor b);
    outputs(3903) <= not a or b;
    outputs(3904) <= not (a or b);
    outputs(3905) <= not b;
    outputs(3906) <= not a;
    outputs(3907) <= a xor b;
    outputs(3908) <= b;
    outputs(3909) <= not (a xor b);
    outputs(3910) <= b;
    outputs(3911) <= b;
    outputs(3912) <= not b;
    outputs(3913) <= not a;
    outputs(3914) <= not a;
    outputs(3915) <= a and not b;
    outputs(3916) <= a and not b;
    outputs(3917) <= a or b;
    outputs(3918) <= not a or b;
    outputs(3919) <= not b;
    outputs(3920) <= not (a xor b);
    outputs(3921) <= a;
    outputs(3922) <= a;
    outputs(3923) <= a or b;
    outputs(3924) <= a xor b;
    outputs(3925) <= a and not b;
    outputs(3926) <= a and b;
    outputs(3927) <= a;
    outputs(3928) <= b;
    outputs(3929) <= not a;
    outputs(3930) <= a and b;
    outputs(3931) <= a and not b;
    outputs(3932) <= not a;
    outputs(3933) <= not a;
    outputs(3934) <= not a;
    outputs(3935) <= b;
    outputs(3936) <= b;
    outputs(3937) <= b;
    outputs(3938) <= a xor b;
    outputs(3939) <= b and not a;
    outputs(3940) <= not a;
    outputs(3941) <= b;
    outputs(3942) <= not (a or b);
    outputs(3943) <= a or b;
    outputs(3944) <= b and not a;
    outputs(3945) <= not a;
    outputs(3946) <= a;
    outputs(3947) <= not b;
    outputs(3948) <= not a;
    outputs(3949) <= not (a or b);
    outputs(3950) <= b;
    outputs(3951) <= not (a or b);
    outputs(3952) <= not (a or b);
    outputs(3953) <= a and b;
    outputs(3954) <= a and b;
    outputs(3955) <= not (a xor b);
    outputs(3956) <= not b;
    outputs(3957) <= b;
    outputs(3958) <= a xor b;
    outputs(3959) <= b;
    outputs(3960) <= not b or a;
    outputs(3961) <= a;
    outputs(3962) <= a xor b;
    outputs(3963) <= a and b;
    outputs(3964) <= a;
    outputs(3965) <= not a or b;
    outputs(3966) <= not (a or b);
    outputs(3967) <= not (a or b);
    outputs(3968) <= not a;
    outputs(3969) <= not (a xor b);
    outputs(3970) <= not (a xor b);
    outputs(3971) <= not (a or b);
    outputs(3972) <= not (a or b);
    outputs(3973) <= a and b;
    outputs(3974) <= a and not b;
    outputs(3975) <= not (a or b);
    outputs(3976) <= not (a and b);
    outputs(3977) <= a;
    outputs(3978) <= not (a xor b);
    outputs(3979) <= a xor b;
    outputs(3980) <= not (a xor b);
    outputs(3981) <= not a;
    outputs(3982) <= a and not b;
    outputs(3983) <= not a;
    outputs(3984) <= not b;
    outputs(3985) <= not b;
    outputs(3986) <= a xor b;
    outputs(3987) <= not (a xor b);
    outputs(3988) <= not b;
    outputs(3989) <= b;
    outputs(3990) <= a and not b;
    outputs(3991) <= not b or a;
    outputs(3992) <= a and not b;
    outputs(3993) <= not b;
    outputs(3994) <= a xor b;
    outputs(3995) <= not b;
    outputs(3996) <= a xor b;
    outputs(3997) <= b and not a;
    outputs(3998) <= not (a xor b);
    outputs(3999) <= not (a xor b);
    outputs(4000) <= a xor b;
    outputs(4001) <= a;
    outputs(4002) <= a or b;
    outputs(4003) <= b;
    outputs(4004) <= a;
    outputs(4005) <= not (a or b);
    outputs(4006) <= a;
    outputs(4007) <= not (a xor b);
    outputs(4008) <= not b;
    outputs(4009) <= a and not b;
    outputs(4010) <= not (a or b);
    outputs(4011) <= b;
    outputs(4012) <= b;
    outputs(4013) <= not b;
    outputs(4014) <= a and b;
    outputs(4015) <= a and not b;
    outputs(4016) <= not a;
    outputs(4017) <= b;
    outputs(4018) <= not a;
    outputs(4019) <= not b;
    outputs(4020) <= a and not b;
    outputs(4021) <= not b;
    outputs(4022) <= a;
    outputs(4023) <= not a;
    outputs(4024) <= b;
    outputs(4025) <= not (a xor b);
    outputs(4026) <= a and not b;
    outputs(4027) <= not b;
    outputs(4028) <= a;
    outputs(4029) <= not (a and b);
    outputs(4030) <= a and not b;
    outputs(4031) <= a and b;
    outputs(4032) <= not a;
    outputs(4033) <= a and b;
    outputs(4034) <= b and not a;
    outputs(4035) <= b and not a;
    outputs(4036) <= a and b;
    outputs(4037) <= a;
    outputs(4038) <= not (a xor b);
    outputs(4039) <= a and not b;
    outputs(4040) <= not a;
    outputs(4041) <= a;
    outputs(4042) <= b;
    outputs(4043) <= a xor b;
    outputs(4044) <= a xor b;
    outputs(4045) <= not (a xor b);
    outputs(4046) <= not (a xor b);
    outputs(4047) <= b;
    outputs(4048) <= not (a xor b);
    outputs(4049) <= b;
    outputs(4050) <= b;
    outputs(4051) <= not b;
    outputs(4052) <= a xor b;
    outputs(4053) <= not (a or b);
    outputs(4054) <= a and b;
    outputs(4055) <= b;
    outputs(4056) <= a and not b;
    outputs(4057) <= not b or a;
    outputs(4058) <= not b;
    outputs(4059) <= not a or b;
    outputs(4060) <= a and b;
    outputs(4061) <= not a or b;
    outputs(4062) <= b and not a;
    outputs(4063) <= b;
    outputs(4064) <= not b;
    outputs(4065) <= a and not b;
    outputs(4066) <= not b;
    outputs(4067) <= a and not b;
    outputs(4068) <= not b;
    outputs(4069) <= not b or a;
    outputs(4070) <= not (a xor b);
    outputs(4071) <= not a;
    outputs(4072) <= a xor b;
    outputs(4073) <= a or b;
    outputs(4074) <= b;
    outputs(4075) <= not (a or b);
    outputs(4076) <= not b;
    outputs(4077) <= b;
    outputs(4078) <= b and not a;
    outputs(4079) <= a or b;
    outputs(4080) <= a;
    outputs(4081) <= b and not a;
    outputs(4082) <= b;
    outputs(4083) <= a;
    outputs(4084) <= a;
    outputs(4085) <= b;
    outputs(4086) <= not a;
    outputs(4087) <= a or b;
    outputs(4088) <= not a;
    outputs(4089) <= a;
    outputs(4090) <= b and not a;
    outputs(4091) <= not a;
    outputs(4092) <= b;
    outputs(4093) <= not b;
    outputs(4094) <= a;
    outputs(4095) <= a or b;
    outputs(4096) <= not (a xor b);
    outputs(4097) <= a;
    outputs(4098) <= not b;
    outputs(4099) <= a;
    outputs(4100) <= not b or a;
    outputs(4101) <= b;
    outputs(4102) <= not (a xor b);
    outputs(4103) <= not b;
    outputs(4104) <= b;
    outputs(4105) <= not b or a;
    outputs(4106) <= not (a or b);
    outputs(4107) <= a and b;
    outputs(4108) <= not (a xor b);
    outputs(4109) <= a xor b;
    outputs(4110) <= not (a xor b);
    outputs(4111) <= not a;
    outputs(4112) <= not b or a;
    outputs(4113) <= a xor b;
    outputs(4114) <= a xor b;
    outputs(4115) <= not (a xor b);
    outputs(4116) <= a and b;
    outputs(4117) <= a;
    outputs(4118) <= not a;
    outputs(4119) <= not a;
    outputs(4120) <= not b;
    outputs(4121) <= a and b;
    outputs(4122) <= a or b;
    outputs(4123) <= not (a xor b);
    outputs(4124) <= a xor b;
    outputs(4125) <= a xor b;
    outputs(4126) <= b;
    outputs(4127) <= not (a xor b);
    outputs(4128) <= not (a xor b);
    outputs(4129) <= a xor b;
    outputs(4130) <= a xor b;
    outputs(4131) <= a;
    outputs(4132) <= not (a xor b);
    outputs(4133) <= a;
    outputs(4134) <= b;
    outputs(4135) <= not (a and b);
    outputs(4136) <= a and b;
    outputs(4137) <= not a or b;
    outputs(4138) <= not (a xor b);
    outputs(4139) <= not b;
    outputs(4140) <= a;
    outputs(4141) <= not (a xor b);
    outputs(4142) <= not (a and b);
    outputs(4143) <= a;
    outputs(4144) <= b;
    outputs(4145) <= not b;
    outputs(4146) <= not b;
    outputs(4147) <= a or b;
    outputs(4148) <= a or b;
    outputs(4149) <= b;
    outputs(4150) <= a and b;
    outputs(4151) <= not b;
    outputs(4152) <= not (a xor b);
    outputs(4153) <= not (a xor b);
    outputs(4154) <= a and b;
    outputs(4155) <= a xor b;
    outputs(4156) <= a xor b;
    outputs(4157) <= not b;
    outputs(4158) <= not b;
    outputs(4159) <= not a;
    outputs(4160) <= not a;
    outputs(4161) <= b and not a;
    outputs(4162) <= a and b;
    outputs(4163) <= not (a xor b);
    outputs(4164) <= not b;
    outputs(4165) <= a or b;
    outputs(4166) <= not b;
    outputs(4167) <= b;
    outputs(4168) <= b;
    outputs(4169) <= not (a or b);
    outputs(4170) <= b;
    outputs(4171) <= a;
    outputs(4172) <= a xor b;
    outputs(4173) <= b;
    outputs(4174) <= a;
    outputs(4175) <= a;
    outputs(4176) <= not (a xor b);
    outputs(4177) <= b;
    outputs(4178) <= not b;
    outputs(4179) <= not b;
    outputs(4180) <= not (a xor b);
    outputs(4181) <= a or b;
    outputs(4182) <= not a;
    outputs(4183) <= a and not b;
    outputs(4184) <= not a or b;
    outputs(4185) <= a;
    outputs(4186) <= not b;
    outputs(4187) <= a and b;
    outputs(4188) <= a xor b;
    outputs(4189) <= not a;
    outputs(4190) <= not b;
    outputs(4191) <= not (a and b);
    outputs(4192) <= a xor b;
    outputs(4193) <= a xor b;
    outputs(4194) <= not (a or b);
    outputs(4195) <= not (a xor b);
    outputs(4196) <= not a or b;
    outputs(4197) <= a xor b;
    outputs(4198) <= a xor b;
    outputs(4199) <= not (a or b);
    outputs(4200) <= a xor b;
    outputs(4201) <= a and not b;
    outputs(4202) <= b;
    outputs(4203) <= a and b;
    outputs(4204) <= not b or a;
    outputs(4205) <= not (a xor b);
    outputs(4206) <= a;
    outputs(4207) <= a;
    outputs(4208) <= a;
    outputs(4209) <= a;
    outputs(4210) <= not b;
    outputs(4211) <= a or b;
    outputs(4212) <= a;
    outputs(4213) <= a xor b;
    outputs(4214) <= a;
    outputs(4215) <= a;
    outputs(4216) <= a and b;
    outputs(4217) <= not (a or b);
    outputs(4218) <= not b;
    outputs(4219) <= b;
    outputs(4220) <= not a;
    outputs(4221) <= b;
    outputs(4222) <= a and b;
    outputs(4223) <= a and b;
    outputs(4224) <= a and not b;
    outputs(4225) <= not a;
    outputs(4226) <= a and not b;
    outputs(4227) <= a and b;
    outputs(4228) <= a xor b;
    outputs(4229) <= b;
    outputs(4230) <= not a;
    outputs(4231) <= a or b;
    outputs(4232) <= a;
    outputs(4233) <= not (a and b);
    outputs(4234) <= a xor b;
    outputs(4235) <= a xor b;
    outputs(4236) <= b and not a;
    outputs(4237) <= not b or a;
    outputs(4238) <= a;
    outputs(4239) <= a xor b;
    outputs(4240) <= a xor b;
    outputs(4241) <= not b;
    outputs(4242) <= not (a xor b);
    outputs(4243) <= a xor b;
    outputs(4244) <= not a;
    outputs(4245) <= b and not a;
    outputs(4246) <= not (a xor b);
    outputs(4247) <= not (a xor b);
    outputs(4248) <= b;
    outputs(4249) <= not b;
    outputs(4250) <= not a;
    outputs(4251) <= not a or b;
    outputs(4252) <= b;
    outputs(4253) <= not (a xor b);
    outputs(4254) <= not (a xor b);
    outputs(4255) <= a xor b;
    outputs(4256) <= not a or b;
    outputs(4257) <= a;
    outputs(4258) <= not b;
    outputs(4259) <= a xor b;
    outputs(4260) <= b and not a;
    outputs(4261) <= not (a xor b);
    outputs(4262) <= not (a xor b);
    outputs(4263) <= b;
    outputs(4264) <= a and not b;
    outputs(4265) <= a xor b;
    outputs(4266) <= a and b;
    outputs(4267) <= b;
    outputs(4268) <= not a;
    outputs(4269) <= a xor b;
    outputs(4270) <= a;
    outputs(4271) <= not b;
    outputs(4272) <= b and not a;
    outputs(4273) <= a xor b;
    outputs(4274) <= a xor b;
    outputs(4275) <= b;
    outputs(4276) <= not (a xor b);
    outputs(4277) <= a;
    outputs(4278) <= not (a xor b);
    outputs(4279) <= not (a xor b);
    outputs(4280) <= not (a and b);
    outputs(4281) <= not (a xor b);
    outputs(4282) <= b and not a;
    outputs(4283) <= not (a or b);
    outputs(4284) <= a;
    outputs(4285) <= b;
    outputs(4286) <= not a or b;
    outputs(4287) <= a xor b;
    outputs(4288) <= not a;
    outputs(4289) <= not (a xor b);
    outputs(4290) <= not (a or b);
    outputs(4291) <= b;
    outputs(4292) <= a xor b;
    outputs(4293) <= not a;
    outputs(4294) <= not (a xor b);
    outputs(4295) <= not (a or b);
    outputs(4296) <= not a or b;
    outputs(4297) <= a xor b;
    outputs(4298) <= not (a xor b);
    outputs(4299) <= not (a and b);
    outputs(4300) <= a and b;
    outputs(4301) <= a or b;
    outputs(4302) <= not a;
    outputs(4303) <= a or b;
    outputs(4304) <= a xor b;
    outputs(4305) <= not b;
    outputs(4306) <= b;
    outputs(4307) <= b;
    outputs(4308) <= b;
    outputs(4309) <= a;
    outputs(4310) <= not b or a;
    outputs(4311) <= not a;
    outputs(4312) <= not (a xor b);
    outputs(4313) <= not (a xor b);
    outputs(4314) <= a;
    outputs(4315) <= a and not b;
    outputs(4316) <= not (a and b);
    outputs(4317) <= not a;
    outputs(4318) <= b and not a;
    outputs(4319) <= a and b;
    outputs(4320) <= not (a xor b);
    outputs(4321) <= a and b;
    outputs(4322) <= not (a and b);
    outputs(4323) <= not (a xor b);
    outputs(4324) <= a;
    outputs(4325) <= not a;
    outputs(4326) <= not b;
    outputs(4327) <= not (a and b);
    outputs(4328) <= not a;
    outputs(4329) <= not (a xor b);
    outputs(4330) <= a;
    outputs(4331) <= not b;
    outputs(4332) <= not (a xor b);
    outputs(4333) <= not (a xor b);
    outputs(4334) <= a and b;
    outputs(4335) <= a xor b;
    outputs(4336) <= not (a xor b);
    outputs(4337) <= b;
    outputs(4338) <= not b;
    outputs(4339) <= a xor b;
    outputs(4340) <= not (a xor b);
    outputs(4341) <= b;
    outputs(4342) <= not a;
    outputs(4343) <= a xor b;
    outputs(4344) <= a xor b;
    outputs(4345) <= not b or a;
    outputs(4346) <= not b or a;
    outputs(4347) <= a;
    outputs(4348) <= not (a xor b);
    outputs(4349) <= a;
    outputs(4350) <= not (a xor b);
    outputs(4351) <= a;
    outputs(4352) <= a;
    outputs(4353) <= not a;
    outputs(4354) <= a;
    outputs(4355) <= a and not b;
    outputs(4356) <= not (a or b);
    outputs(4357) <= a;
    outputs(4358) <= a xor b;
    outputs(4359) <= not (a xor b);
    outputs(4360) <= b;
    outputs(4361) <= not (a xor b);
    outputs(4362) <= not (a xor b);
    outputs(4363) <= a xor b;
    outputs(4364) <= not (a or b);
    outputs(4365) <= not b;
    outputs(4366) <= not (a and b);
    outputs(4367) <= not (a xor b);
    outputs(4368) <= not b;
    outputs(4369) <= a xor b;
    outputs(4370) <= not (a and b);
    outputs(4371) <= not b;
    outputs(4372) <= not (a xor b);
    outputs(4373) <= not (a xor b);
    outputs(4374) <= not (a or b);
    outputs(4375) <= not (a xor b);
    outputs(4376) <= not (a xor b);
    outputs(4377) <= not a;
    outputs(4378) <= a;
    outputs(4379) <= not (a xor b);
    outputs(4380) <= not (a and b);
    outputs(4381) <= b and not a;
    outputs(4382) <= a xor b;
    outputs(4383) <= not a;
    outputs(4384) <= not b;
    outputs(4385) <= a xor b;
    outputs(4386) <= a or b;
    outputs(4387) <= b;
    outputs(4388) <= not a;
    outputs(4389) <= not a;
    outputs(4390) <= not b;
    outputs(4391) <= a xor b;
    outputs(4392) <= a;
    outputs(4393) <= not b;
    outputs(4394) <= not b or a;
    outputs(4395) <= not a;
    outputs(4396) <= not a;
    outputs(4397) <= b;
    outputs(4398) <= a;
    outputs(4399) <= not (a xor b);
    outputs(4400) <= a xor b;
    outputs(4401) <= a xor b;
    outputs(4402) <= not b;
    outputs(4403) <= a xor b;
    outputs(4404) <= not (a xor b);
    outputs(4405) <= not (a xor b);
    outputs(4406) <= a and b;
    outputs(4407) <= not a;
    outputs(4408) <= a;
    outputs(4409) <= a xor b;
    outputs(4410) <= a xor b;
    outputs(4411) <= a xor b;
    outputs(4412) <= b;
    outputs(4413) <= a and not b;
    outputs(4414) <= a and not b;
    outputs(4415) <= a xor b;
    outputs(4416) <= not (a xor b);
    outputs(4417) <= a xor b;
    outputs(4418) <= a or b;
    outputs(4419) <= a;
    outputs(4420) <= not a;
    outputs(4421) <= a and not b;
    outputs(4422) <= not (a xor b);
    outputs(4423) <= not b;
    outputs(4424) <= b and not a;
    outputs(4425) <= a and not b;
    outputs(4426) <= a xor b;
    outputs(4427) <= not (a xor b);
    outputs(4428) <= a and not b;
    outputs(4429) <= b and not a;
    outputs(4430) <= not b;
    outputs(4431) <= b and not a;
    outputs(4432) <= a xor b;
    outputs(4433) <= not (a xor b);
    outputs(4434) <= a;
    outputs(4435) <= a xor b;
    outputs(4436) <= a;
    outputs(4437) <= not (a xor b);
    outputs(4438) <= not b or a;
    outputs(4439) <= not a;
    outputs(4440) <= b;
    outputs(4441) <= a;
    outputs(4442) <= a xor b;
    outputs(4443) <= not (a xor b);
    outputs(4444) <= not a;
    outputs(4445) <= a xor b;
    outputs(4446) <= not b;
    outputs(4447) <= not b;
    outputs(4448) <= not b;
    outputs(4449) <= a xor b;
    outputs(4450) <= not (a xor b);
    outputs(4451) <= a or b;
    outputs(4452) <= not (a xor b);
    outputs(4453) <= not a;
    outputs(4454) <= not (a xor b);
    outputs(4455) <= not (a xor b);
    outputs(4456) <= b;
    outputs(4457) <= not b;
    outputs(4458) <= not a;
    outputs(4459) <= b and not a;
    outputs(4460) <= b;
    outputs(4461) <= b;
    outputs(4462) <= a xor b;
    outputs(4463) <= not b;
    outputs(4464) <= not a;
    outputs(4465) <= not (a xor b);
    outputs(4466) <= not (a xor b);
    outputs(4467) <= a xor b;
    outputs(4468) <= not (a or b);
    outputs(4469) <= not a or b;
    outputs(4470) <= b;
    outputs(4471) <= b;
    outputs(4472) <= b;
    outputs(4473) <= b;
    outputs(4474) <= a xor b;
    outputs(4475) <= a;
    outputs(4476) <= not b;
    outputs(4477) <= not (a or b);
    outputs(4478) <= a xor b;
    outputs(4479) <= not b;
    outputs(4480) <= a;
    outputs(4481) <= b;
    outputs(4482) <= not (a xor b);
    outputs(4483) <= a and b;
    outputs(4484) <= b;
    outputs(4485) <= not (a xor b);
    outputs(4486) <= a xor b;
    outputs(4487) <= a;
    outputs(4488) <= a xor b;
    outputs(4489) <= not b;
    outputs(4490) <= a xor b;
    outputs(4491) <= a xor b;
    outputs(4492) <= not b;
    outputs(4493) <= a or b;
    outputs(4494) <= b and not a;
    outputs(4495) <= not a;
    outputs(4496) <= not (a xor b);
    outputs(4497) <= not b;
    outputs(4498) <= not a;
    outputs(4499) <= not (a xor b);
    outputs(4500) <= b;
    outputs(4501) <= a xor b;
    outputs(4502) <= a or b;
    outputs(4503) <= not b;
    outputs(4504) <= b;
    outputs(4505) <= not (a xor b);
    outputs(4506) <= a xor b;
    outputs(4507) <= a and b;
    outputs(4508) <= not b;
    outputs(4509) <= not (a xor b);
    outputs(4510) <= a xor b;
    outputs(4511) <= not a;
    outputs(4512) <= not (a xor b);
    outputs(4513) <= a xor b;
    outputs(4514) <= a xor b;
    outputs(4515) <= not b;
    outputs(4516) <= not b;
    outputs(4517) <= a xor b;
    outputs(4518) <= a xor b;
    outputs(4519) <= not a or b;
    outputs(4520) <= b and not a;
    outputs(4521) <= not (a and b);
    outputs(4522) <= a;
    outputs(4523) <= b;
    outputs(4524) <= b and not a;
    outputs(4525) <= b and not a;
    outputs(4526) <= a and not b;
    outputs(4527) <= not (a xor b);
    outputs(4528) <= a and not b;
    outputs(4529) <= not a;
    outputs(4530) <= a xor b;
    outputs(4531) <= a and b;
    outputs(4532) <= a and not b;
    outputs(4533) <= b and not a;
    outputs(4534) <= not a;
    outputs(4535) <= b;
    outputs(4536) <= not b or a;
    outputs(4537) <= a xor b;
    outputs(4538) <= not (a xor b);
    outputs(4539) <= not b or a;
    outputs(4540) <= a;
    outputs(4541) <= b;
    outputs(4542) <= not a;
    outputs(4543) <= not b;
    outputs(4544) <= not b;
    outputs(4545) <= b;
    outputs(4546) <= not b;
    outputs(4547) <= a;
    outputs(4548) <= not (a xor b);
    outputs(4549) <= b and not a;
    outputs(4550) <= a xor b;
    outputs(4551) <= not b;
    outputs(4552) <= not (a xor b);
    outputs(4553) <= not b;
    outputs(4554) <= a or b;
    outputs(4555) <= not (a xor b);
    outputs(4556) <= b;
    outputs(4557) <= not a;
    outputs(4558) <= not (a xor b);
    outputs(4559) <= not (a xor b);
    outputs(4560) <= a xor b;
    outputs(4561) <= not b;
    outputs(4562) <= a;
    outputs(4563) <= not a;
    outputs(4564) <= not a or b;
    outputs(4565) <= not (a and b);
    outputs(4566) <= a and not b;
    outputs(4567) <= a xor b;
    outputs(4568) <= not a;
    outputs(4569) <= not (a xor b);
    outputs(4570) <= a;
    outputs(4571) <= not (a or b);
    outputs(4572) <= a xor b;
    outputs(4573) <= a or b;
    outputs(4574) <= not a;
    outputs(4575) <= a xor b;
    outputs(4576) <= a;
    outputs(4577) <= not b;
    outputs(4578) <= a xor b;
    outputs(4579) <= not b;
    outputs(4580) <= not b;
    outputs(4581) <= not b;
    outputs(4582) <= not b;
    outputs(4583) <= not (a xor b);
    outputs(4584) <= not (a or b);
    outputs(4585) <= not a;
    outputs(4586) <= b;
    outputs(4587) <= b;
    outputs(4588) <= not a;
    outputs(4589) <= not a;
    outputs(4590) <= not a or b;
    outputs(4591) <= not (a xor b);
    outputs(4592) <= not a;
    outputs(4593) <= not a;
    outputs(4594) <= not (a xor b);
    outputs(4595) <= a;
    outputs(4596) <= b;
    outputs(4597) <= not (a xor b);
    outputs(4598) <= b;
    outputs(4599) <= a;
    outputs(4600) <= b;
    outputs(4601) <= not (a xor b);
    outputs(4602) <= b;
    outputs(4603) <= a;
    outputs(4604) <= a xor b;
    outputs(4605) <= a xor b;
    outputs(4606) <= a;
    outputs(4607) <= a xor b;
    outputs(4608) <= not (a or b);
    outputs(4609) <= a and not b;
    outputs(4610) <= b;
    outputs(4611) <= b and not a;
    outputs(4612) <= a and b;
    outputs(4613) <= a xor b;
    outputs(4614) <= a and b;
    outputs(4615) <= not a;
    outputs(4616) <= a or b;
    outputs(4617) <= a xor b;
    outputs(4618) <= a xor b;
    outputs(4619) <= b;
    outputs(4620) <= not (a or b);
    outputs(4621) <= a xor b;
    outputs(4622) <= b;
    outputs(4623) <= not a;
    outputs(4624) <= a and b;
    outputs(4625) <= a;
    outputs(4626) <= b and not a;
    outputs(4627) <= not a;
    outputs(4628) <= not (a and b);
    outputs(4629) <= not b;
    outputs(4630) <= b and not a;
    outputs(4631) <= not a;
    outputs(4632) <= b and not a;
    outputs(4633) <= a;
    outputs(4634) <= a xor b;
    outputs(4635) <= a xor b;
    outputs(4636) <= not (a xor b);
    outputs(4637) <= a;
    outputs(4638) <= a xor b;
    outputs(4639) <= not (a xor b);
    outputs(4640) <= a xor b;
    outputs(4641) <= a;
    outputs(4642) <= not (a xor b);
    outputs(4643) <= not a or b;
    outputs(4644) <= a and b;
    outputs(4645) <= not b;
    outputs(4646) <= b;
    outputs(4647) <= not a;
    outputs(4648) <= a and not b;
    outputs(4649) <= not (a or b);
    outputs(4650) <= not b;
    outputs(4651) <= b;
    outputs(4652) <= not a;
    outputs(4653) <= not a;
    outputs(4654) <= not a;
    outputs(4655) <= a;
    outputs(4656) <= not (a or b);
    outputs(4657) <= a xor b;
    outputs(4658) <= not b;
    outputs(4659) <= a and not b;
    outputs(4660) <= a and not b;
    outputs(4661) <= a and b;
    outputs(4662) <= b and not a;
    outputs(4663) <= b;
    outputs(4664) <= a;
    outputs(4665) <= b;
    outputs(4666) <= a xor b;
    outputs(4667) <= a xor b;
    outputs(4668) <= a;
    outputs(4669) <= a xor b;
    outputs(4670) <= a and not b;
    outputs(4671) <= b;
    outputs(4672) <= not (a xor b);
    outputs(4673) <= a xor b;
    outputs(4674) <= a and b;
    outputs(4675) <= not a or b;
    outputs(4676) <= b and not a;
    outputs(4677) <= not (a or b);
    outputs(4678) <= a xor b;
    outputs(4679) <= b;
    outputs(4680) <= not (a and b);
    outputs(4681) <= b;
    outputs(4682) <= not (a xor b);
    outputs(4683) <= a or b;
    outputs(4684) <= not b;
    outputs(4685) <= a and b;
    outputs(4686) <= not (a xor b);
    outputs(4687) <= a xor b;
    outputs(4688) <= not b;
    outputs(4689) <= not (a and b);
    outputs(4690) <= b and not a;
    outputs(4691) <= a xor b;
    outputs(4692) <= a and b;
    outputs(4693) <= a xor b;
    outputs(4694) <= b;
    outputs(4695) <= a;
    outputs(4696) <= a xor b;
    outputs(4697) <= not (a xor b);
    outputs(4698) <= b;
    outputs(4699) <= b and not a;
    outputs(4700) <= not a;
    outputs(4701) <= a;
    outputs(4702) <= a and not b;
    outputs(4703) <= b;
    outputs(4704) <= not a or b;
    outputs(4705) <= not (a xor b);
    outputs(4706) <= not (a xor b);
    outputs(4707) <= b and not a;
    outputs(4708) <= not (a and b);
    outputs(4709) <= a xor b;
    outputs(4710) <= a;
    outputs(4711) <= b;
    outputs(4712) <= b;
    outputs(4713) <= not (a or b);
    outputs(4714) <= b;
    outputs(4715) <= b;
    outputs(4716) <= not b;
    outputs(4717) <= not (a xor b);
    outputs(4718) <= a;
    outputs(4719) <= a xor b;
    outputs(4720) <= not (a or b);
    outputs(4721) <= a;
    outputs(4722) <= not b;
    outputs(4723) <= not a;
    outputs(4724) <= not (a xor b);
    outputs(4725) <= b;
    outputs(4726) <= not (a or b);
    outputs(4727) <= b and not a;
    outputs(4728) <= not a;
    outputs(4729) <= not b;
    outputs(4730) <= a;
    outputs(4731) <= a and b;
    outputs(4732) <= a xor b;
    outputs(4733) <= not a;
    outputs(4734) <= not (a xor b);
    outputs(4735) <= a xor b;
    outputs(4736) <= not (a xor b);
    outputs(4737) <= b;
    outputs(4738) <= not b;
    outputs(4739) <= not b;
    outputs(4740) <= not (a xor b);
    outputs(4741) <= not (a xor b);
    outputs(4742) <= b;
    outputs(4743) <= b;
    outputs(4744) <= not a;
    outputs(4745) <= b;
    outputs(4746) <= b;
    outputs(4747) <= a or b;
    outputs(4748) <= not b;
    outputs(4749) <= not (a or b);
    outputs(4750) <= not (a xor b);
    outputs(4751) <= a;
    outputs(4752) <= not a or b;
    outputs(4753) <= not (a xor b);
    outputs(4754) <= not b;
    outputs(4755) <= not a;
    outputs(4756) <= b;
    outputs(4757) <= not (a xor b);
    outputs(4758) <= a and not b;
    outputs(4759) <= b;
    outputs(4760) <= not a;
    outputs(4761) <= a;
    outputs(4762) <= b;
    outputs(4763) <= not a;
    outputs(4764) <= not a;
    outputs(4765) <= b;
    outputs(4766) <= not (a xor b);
    outputs(4767) <= not (a xor b);
    outputs(4768) <= not (a and b);
    outputs(4769) <= not a;
    outputs(4770) <= not (a xor b);
    outputs(4771) <= a;
    outputs(4772) <= b;
    outputs(4773) <= not b;
    outputs(4774) <= not (a xor b);
    outputs(4775) <= not b;
    outputs(4776) <= a and b;
    outputs(4777) <= a and b;
    outputs(4778) <= a or b;
    outputs(4779) <= not a;
    outputs(4780) <= a;
    outputs(4781) <= not (a or b);
    outputs(4782) <= not b;
    outputs(4783) <= a and not b;
    outputs(4784) <= not a;
    outputs(4785) <= a xor b;
    outputs(4786) <= b;
    outputs(4787) <= not (a or b);
    outputs(4788) <= not (a or b);
    outputs(4789) <= not a;
    outputs(4790) <= a and b;
    outputs(4791) <= a xor b;
    outputs(4792) <= a and not b;
    outputs(4793) <= a xor b;
    outputs(4794) <= not (a xor b);
    outputs(4795) <= a and not b;
    outputs(4796) <= a xor b;
    outputs(4797) <= b;
    outputs(4798) <= a xor b;
    outputs(4799) <= not b;
    outputs(4800) <= b and not a;
    outputs(4801) <= not (a xor b);
    outputs(4802) <= a xor b;
    outputs(4803) <= b;
    outputs(4804) <= b;
    outputs(4805) <= a;
    outputs(4806) <= a xor b;
    outputs(4807) <= a xor b;
    outputs(4808) <= a xor b;
    outputs(4809) <= a xor b;
    outputs(4810) <= b and not a;
    outputs(4811) <= not b;
    outputs(4812) <= a xor b;
    outputs(4813) <= not (a and b);
    outputs(4814) <= b;
    outputs(4815) <= a;
    outputs(4816) <= not (a xor b);
    outputs(4817) <= not b;
    outputs(4818) <= not a;
    outputs(4819) <= not a or b;
    outputs(4820) <= not a;
    outputs(4821) <= not (a xor b);
    outputs(4822) <= not a;
    outputs(4823) <= b and not a;
    outputs(4824) <= b;
    outputs(4825) <= b and not a;
    outputs(4826) <= a xor b;
    outputs(4827) <= a;
    outputs(4828) <= a or b;
    outputs(4829) <= not (a xor b);
    outputs(4830) <= a xor b;
    outputs(4831) <= a or b;
    outputs(4832) <= not a;
    outputs(4833) <= a xor b;
    outputs(4834) <= not a;
    outputs(4835) <= a xor b;
    outputs(4836) <= a xor b;
    outputs(4837) <= not b;
    outputs(4838) <= not b;
    outputs(4839) <= b;
    outputs(4840) <= not a;
    outputs(4841) <= not (a or b);
    outputs(4842) <= not b;
    outputs(4843) <= not b;
    outputs(4844) <= not b;
    outputs(4845) <= a xor b;
    outputs(4846) <= not (a xor b);
    outputs(4847) <= b and not a;
    outputs(4848) <= not a;
    outputs(4849) <= a;
    outputs(4850) <= not b;
    outputs(4851) <= not (a xor b);
    outputs(4852) <= a xor b;
    outputs(4853) <= not (a or b);
    outputs(4854) <= b;
    outputs(4855) <= not a;
    outputs(4856) <= a or b;
    outputs(4857) <= a and not b;
    outputs(4858) <= not (a xor b);
    outputs(4859) <= not b;
    outputs(4860) <= not (a xor b);
    outputs(4861) <= a xor b;
    outputs(4862) <= not b;
    outputs(4863) <= b;
    outputs(4864) <= not b or a;
    outputs(4865) <= b;
    outputs(4866) <= not b;
    outputs(4867) <= not b;
    outputs(4868) <= not a;
    outputs(4869) <= a and not b;
    outputs(4870) <= a;
    outputs(4871) <= not (a and b);
    outputs(4872) <= a xor b;
    outputs(4873) <= not (a and b);
    outputs(4874) <= a and b;
    outputs(4875) <= not (a xor b);
    outputs(4876) <= a and not b;
    outputs(4877) <= b;
    outputs(4878) <= a and b;
    outputs(4879) <= '1';
    outputs(4880) <= a xor b;
    outputs(4881) <= not a;
    outputs(4882) <= not b;
    outputs(4883) <= a or b;
    outputs(4884) <= not (a or b);
    outputs(4885) <= a and not b;
    outputs(4886) <= b;
    outputs(4887) <= not a;
    outputs(4888) <= not (a or b);
    outputs(4889) <= not (a or b);
    outputs(4890) <= a;
    outputs(4891) <= not b;
    outputs(4892) <= a xor b;
    outputs(4893) <= not (a and b);
    outputs(4894) <= a and not b;
    outputs(4895) <= b;
    outputs(4896) <= b and not a;
    outputs(4897) <= a xor b;
    outputs(4898) <= not b or a;
    outputs(4899) <= a or b;
    outputs(4900) <= a and not b;
    outputs(4901) <= a and b;
    outputs(4902) <= a or b;
    outputs(4903) <= b;
    outputs(4904) <= not (a xor b);
    outputs(4905) <= not (a and b);
    outputs(4906) <= b;
    outputs(4907) <= not (a xor b);
    outputs(4908) <= not a;
    outputs(4909) <= not a;
    outputs(4910) <= not a;
    outputs(4911) <= not b;
    outputs(4912) <= not a or b;
    outputs(4913) <= a xor b;
    outputs(4914) <= b;
    outputs(4915) <= not a;
    outputs(4916) <= not a;
    outputs(4917) <= a;
    outputs(4918) <= a xor b;
    outputs(4919) <= a and b;
    outputs(4920) <= not (a or b);
    outputs(4921) <= a and not b;
    outputs(4922) <= a;
    outputs(4923) <= not (a xor b);
    outputs(4924) <= not a;
    outputs(4925) <= b;
    outputs(4926) <= not b or a;
    outputs(4927) <= b;
    outputs(4928) <= not (a xor b);
    outputs(4929) <= a and b;
    outputs(4930) <= b and not a;
    outputs(4931) <= not a;
    outputs(4932) <= not (a xor b);
    outputs(4933) <= a and b;
    outputs(4934) <= not (a xor b);
    outputs(4935) <= not (a xor b);
    outputs(4936) <= b;
    outputs(4937) <= not (a xor b);
    outputs(4938) <= not b;
    outputs(4939) <= not a;
    outputs(4940) <= b;
    outputs(4941) <= not b;
    outputs(4942) <= not (a or b);
    outputs(4943) <= not (a xor b);
    outputs(4944) <= not a;
    outputs(4945) <= not b;
    outputs(4946) <= b;
    outputs(4947) <= not (a or b);
    outputs(4948) <= a;
    outputs(4949) <= not a;
    outputs(4950) <= not (a or b);
    outputs(4951) <= a;
    outputs(4952) <= a;
    outputs(4953) <= not (a xor b);
    outputs(4954) <= not a;
    outputs(4955) <= not (a xor b);
    outputs(4956) <= a xor b;
    outputs(4957) <= not b;
    outputs(4958) <= not b;
    outputs(4959) <= a and not b;
    outputs(4960) <= b;
    outputs(4961) <= a or b;
    outputs(4962) <= not (a xor b);
    outputs(4963) <= a and not b;
    outputs(4964) <= b and not a;
    outputs(4965) <= not a;
    outputs(4966) <= a xor b;
    outputs(4967) <= not a;
    outputs(4968) <= a xor b;
    outputs(4969) <= a xor b;
    outputs(4970) <= a xor b;
    outputs(4971) <= a and not b;
    outputs(4972) <= not b;
    outputs(4973) <= a;
    outputs(4974) <= b and not a;
    outputs(4975) <= b;
    outputs(4976) <= not (a xor b);
    outputs(4977) <= not b;
    outputs(4978) <= a and b;
    outputs(4979) <= a;
    outputs(4980) <= not (a and b);
    outputs(4981) <= not b;
    outputs(4982) <= a;
    outputs(4983) <= a and b;
    outputs(4984) <= not (a xor b);
    outputs(4985) <= not (a and b);
    outputs(4986) <= not (a and b);
    outputs(4987) <= not (a or b);
    outputs(4988) <= a xor b;
    outputs(4989) <= b and not a;
    outputs(4990) <= b;
    outputs(4991) <= a or b;
    outputs(4992) <= not a;
    outputs(4993) <= a xor b;
    outputs(4994) <= a xor b;
    outputs(4995) <= not (a and b);
    outputs(4996) <= b and not a;
    outputs(4997) <= b;
    outputs(4998) <= not a;
    outputs(4999) <= a xor b;
    outputs(5000) <= a xor b;
    outputs(5001) <= not (a or b);
    outputs(5002) <= a;
    outputs(5003) <= not a;
    outputs(5004) <= not (a or b);
    outputs(5005) <= not (a xor b);
    outputs(5006) <= a xor b;
    outputs(5007) <= not b;
    outputs(5008) <= a;
    outputs(5009) <= b;
    outputs(5010) <= not b;
    outputs(5011) <= a or b;
    outputs(5012) <= a;
    outputs(5013) <= not b or a;
    outputs(5014) <= not b or a;
    outputs(5015) <= a and not b;
    outputs(5016) <= not a;
    outputs(5017) <= b;
    outputs(5018) <= not (a xor b);
    outputs(5019) <= not b;
    outputs(5020) <= a and not b;
    outputs(5021) <= b and not a;
    outputs(5022) <= a and b;
    outputs(5023) <= a xor b;
    outputs(5024) <= not (a xor b);
    outputs(5025) <= a and b;
    outputs(5026) <= a xor b;
    outputs(5027) <= not (a or b);
    outputs(5028) <= b;
    outputs(5029) <= not b;
    outputs(5030) <= not b;
    outputs(5031) <= a xor b;
    outputs(5032) <= a and not b;
    outputs(5033) <= not (a xor b);
    outputs(5034) <= b;
    outputs(5035) <= not b;
    outputs(5036) <= a and b;
    outputs(5037) <= not (a or b);
    outputs(5038) <= a xor b;
    outputs(5039) <= a and b;
    outputs(5040) <= not (a xor b);
    outputs(5041) <= not (a xor b);
    outputs(5042) <= b and not a;
    outputs(5043) <= not (a xor b);
    outputs(5044) <= not (a or b);
    outputs(5045) <= a;
    outputs(5046) <= not (a xor b);
    outputs(5047) <= not (a or b);
    outputs(5048) <= not a;
    outputs(5049) <= b;
    outputs(5050) <= b;
    outputs(5051) <= a and b;
    outputs(5052) <= not b;
    outputs(5053) <= not b;
    outputs(5054) <= a or b;
    outputs(5055) <= b;
    outputs(5056) <= not (a or b);
    outputs(5057) <= not b;
    outputs(5058) <= a and not b;
    outputs(5059) <= not (a xor b);
    outputs(5060) <= not (a or b);
    outputs(5061) <= b and not a;
    outputs(5062) <= a and not b;
    outputs(5063) <= b;
    outputs(5064) <= not a;
    outputs(5065) <= not (a xor b);
    outputs(5066) <= a and not b;
    outputs(5067) <= a xor b;
    outputs(5068) <= not (a xor b);
    outputs(5069) <= a;
    outputs(5070) <= a or b;
    outputs(5071) <= a;
    outputs(5072) <= b;
    outputs(5073) <= b;
    outputs(5074) <= not (a or b);
    outputs(5075) <= not (a or b);
    outputs(5076) <= a;
    outputs(5077) <= not a;
    outputs(5078) <= not (a xor b);
    outputs(5079) <= not a;
    outputs(5080) <= b and not a;
    outputs(5081) <= not a or b;
    outputs(5082) <= not (a xor b);
    outputs(5083) <= a and not b;
    outputs(5084) <= a;
    outputs(5085) <= b and not a;
    outputs(5086) <= a and b;
    outputs(5087) <= a;
    outputs(5088) <= not (a or b);
    outputs(5089) <= b and not a;
    outputs(5090) <= not a;
    outputs(5091) <= not (a xor b);
    outputs(5092) <= a xor b;
    outputs(5093) <= not a;
    outputs(5094) <= not b;
    outputs(5095) <= not (a xor b);
    outputs(5096) <= b;
    outputs(5097) <= not b;
    outputs(5098) <= not b;
    outputs(5099) <= b and not a;
    outputs(5100) <= not b;
    outputs(5101) <= b and not a;
    outputs(5102) <= not (a xor b);
    outputs(5103) <= not b;
    outputs(5104) <= not a;
    outputs(5105) <= a;
    outputs(5106) <= not a;
    outputs(5107) <= a and not b;
    outputs(5108) <= b;
    outputs(5109) <= not b;
    outputs(5110) <= a;
    outputs(5111) <= not a or b;
    outputs(5112) <= not a or b;
    outputs(5113) <= b;
    outputs(5114) <= a;
    outputs(5115) <= a xor b;
    outputs(5116) <= a and b;
    outputs(5117) <= a;
    outputs(5118) <= not (a xor b);
    outputs(5119) <= not (a xor b);
end Behavioral;
