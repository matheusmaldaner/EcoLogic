library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs: in std_logic_vector(1023 downto 0);
        outputs: out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs: std_logic_vector(5119 downto 0);

begin
    layer0_outputs(0) <= not (a or b);
    layer0_outputs(1) <= b;
    layer0_outputs(2) <= a xor b;
    layer0_outputs(3) <= a or b;
    layer0_outputs(4) <= not a or b;
    layer0_outputs(5) <= not (a or b);
    layer0_outputs(6) <= a xor b;
    layer0_outputs(7) <= not a or b;
    layer0_outputs(8) <= not b or a;
    layer0_outputs(9) <= a and b;
    layer0_outputs(10) <= not (a or b);
    layer0_outputs(11) <= a xor b;
    layer0_outputs(12) <= a and not b;
    layer0_outputs(13) <= not b or a;
    layer0_outputs(14) <= b;
    layer0_outputs(15) <= a or b;
    layer0_outputs(16) <= not (a or b);
    layer0_outputs(17) <= a;
    layer0_outputs(18) <= a xor b;
    layer0_outputs(19) <= a or b;
    layer0_outputs(20) <= a and b;
    layer0_outputs(21) <= b;
    layer0_outputs(22) <= not (a xor b);
    layer0_outputs(23) <= not a or b;
    layer0_outputs(24) <= not b or a;
    layer0_outputs(25) <= a or b;
    layer0_outputs(26) <= not b or a;
    layer0_outputs(27) <= a or b;
    layer0_outputs(28) <= a xor b;
    layer0_outputs(29) <= '1';
    layer0_outputs(30) <= not a or b;
    layer0_outputs(31) <= not (a or b);
    layer0_outputs(32) <= not (a or b);
    layer0_outputs(33) <= '0';
    layer0_outputs(34) <= b and not a;
    layer0_outputs(35) <= not b;
    layer0_outputs(36) <= not (a or b);
    layer0_outputs(37) <= not b or a;
    layer0_outputs(38) <= a;
    layer0_outputs(39) <= a;
    layer0_outputs(40) <= not (a xor b);
    layer0_outputs(41) <= b and not a;
    layer0_outputs(42) <= a xor b;
    layer0_outputs(43) <= b;
    layer0_outputs(44) <= a;
    layer0_outputs(45) <= not b or a;
    layer0_outputs(46) <= a and not b;
    layer0_outputs(47) <= not a;
    layer0_outputs(48) <= not (a xor b);
    layer0_outputs(49) <= a;
    layer0_outputs(50) <= not b;
    layer0_outputs(51) <= not (a or b);
    layer0_outputs(52) <= not a;
    layer0_outputs(53) <= b and not a;
    layer0_outputs(54) <= not (a xor b);
    layer0_outputs(55) <= b and not a;
    layer0_outputs(56) <= a and not b;
    layer0_outputs(57) <= a or b;
    layer0_outputs(58) <= not a;
    layer0_outputs(59) <= b;
    layer0_outputs(60) <= a xor b;
    layer0_outputs(61) <= not b or a;
    layer0_outputs(62) <= not (a xor b);
    layer0_outputs(63) <= a;
    layer0_outputs(64) <= a;
    layer0_outputs(65) <= not (a or b);
    layer0_outputs(66) <= not a or b;
    layer0_outputs(67) <= b and not a;
    layer0_outputs(68) <= a xor b;
    layer0_outputs(69) <= a or b;
    layer0_outputs(70) <= not b;
    layer0_outputs(71) <= not (a and b);
    layer0_outputs(72) <= a or b;
    layer0_outputs(73) <= a or b;
    layer0_outputs(74) <= a;
    layer0_outputs(75) <= b and not a;
    layer0_outputs(76) <= not (a or b);
    layer0_outputs(77) <= b;
    layer0_outputs(78) <= not b;
    layer0_outputs(79) <= not b;
    layer0_outputs(80) <= not (a or b);
    layer0_outputs(81) <= a or b;
    layer0_outputs(82) <= a or b;
    layer0_outputs(83) <= not b;
    layer0_outputs(84) <= b;
    layer0_outputs(85) <= not a;
    layer0_outputs(86) <= not (a or b);
    layer0_outputs(87) <= a or b;
    layer0_outputs(88) <= not b;
    layer0_outputs(89) <= not b;
    layer0_outputs(90) <= not (a xor b);
    layer0_outputs(91) <= not (a or b);
    layer0_outputs(92) <= b;
    layer0_outputs(93) <= not (a xor b);
    layer0_outputs(94) <= not b;
    layer0_outputs(95) <= not (a or b);
    layer0_outputs(96) <= not a;
    layer0_outputs(97) <= a xor b;
    layer0_outputs(98) <= not (a or b);
    layer0_outputs(99) <= a and not b;
    layer0_outputs(100) <= b;
    layer0_outputs(101) <= '0';
    layer0_outputs(102) <= not b;
    layer0_outputs(103) <= a xor b;
    layer0_outputs(104) <= b and not a;
    layer0_outputs(105) <= b;
    layer0_outputs(106) <= b;
    layer0_outputs(107) <= a xor b;
    layer0_outputs(108) <= a and not b;
    layer0_outputs(109) <= b;
    layer0_outputs(110) <= a xor b;
    layer0_outputs(111) <= a and not b;
    layer0_outputs(112) <= not a;
    layer0_outputs(113) <= b;
    layer0_outputs(114) <= b;
    layer0_outputs(115) <= not (a xor b);
    layer0_outputs(116) <= a or b;
    layer0_outputs(117) <= a and not b;
    layer0_outputs(118) <= b and not a;
    layer0_outputs(119) <= a and not b;
    layer0_outputs(120) <= not a or b;
    layer0_outputs(121) <= a or b;
    layer0_outputs(122) <= not b or a;
    layer0_outputs(123) <= a or b;
    layer0_outputs(124) <= a or b;
    layer0_outputs(125) <= a;
    layer0_outputs(126) <= a or b;
    layer0_outputs(127) <= not (a xor b);
    layer0_outputs(128) <= not b;
    layer0_outputs(129) <= b and not a;
    layer0_outputs(130) <= not b;
    layer0_outputs(131) <= a and not b;
    layer0_outputs(132) <= not (a xor b);
    layer0_outputs(133) <= not (a xor b);
    layer0_outputs(134) <= b;
    layer0_outputs(135) <= b;
    layer0_outputs(136) <= not a or b;
    layer0_outputs(137) <= a xor b;
    layer0_outputs(138) <= not b;
    layer0_outputs(139) <= not (a xor b);
    layer0_outputs(140) <= not (a or b);
    layer0_outputs(141) <= not a;
    layer0_outputs(142) <= a xor b;
    layer0_outputs(143) <= not b or a;
    layer0_outputs(144) <= not b;
    layer0_outputs(145) <= b and not a;
    layer0_outputs(146) <= a;
    layer0_outputs(147) <= not (a xor b);
    layer0_outputs(148) <= a and not b;
    layer0_outputs(149) <= a or b;
    layer0_outputs(150) <= b;
    layer0_outputs(151) <= a and not b;
    layer0_outputs(152) <= a and not b;
    layer0_outputs(153) <= not (a and b);
    layer0_outputs(154) <= b;
    layer0_outputs(155) <= b and not a;
    layer0_outputs(156) <= not b;
    layer0_outputs(157) <= '0';
    layer0_outputs(158) <= '1';
    layer0_outputs(159) <= a xor b;
    layer0_outputs(160) <= a and not b;
    layer0_outputs(161) <= not (a or b);
    layer0_outputs(162) <= a or b;
    layer0_outputs(163) <= a and not b;
    layer0_outputs(164) <= a;
    layer0_outputs(165) <= '1';
    layer0_outputs(166) <= not b or a;
    layer0_outputs(167) <= not b or a;
    layer0_outputs(168) <= a;
    layer0_outputs(169) <= not a or b;
    layer0_outputs(170) <= '1';
    layer0_outputs(171) <= not (a or b);
    layer0_outputs(172) <= not (a or b);
    layer0_outputs(173) <= not (a or b);
    layer0_outputs(174) <= a and not b;
    layer0_outputs(175) <= b;
    layer0_outputs(176) <= not (a and b);
    layer0_outputs(177) <= not (a and b);
    layer0_outputs(178) <= b;
    layer0_outputs(179) <= not (a xor b);
    layer0_outputs(180) <= a or b;
    layer0_outputs(181) <= a;
    layer0_outputs(182) <= not (a or b);
    layer0_outputs(183) <= not (a or b);
    layer0_outputs(184) <= a xor b;
    layer0_outputs(185) <= not (a or b);
    layer0_outputs(186) <= b;
    layer0_outputs(187) <= a;
    layer0_outputs(188) <= a or b;
    layer0_outputs(189) <= not (a and b);
    layer0_outputs(190) <= not (a xor b);
    layer0_outputs(191) <= not (a or b);
    layer0_outputs(192) <= not (a xor b);
    layer0_outputs(193) <= not b;
    layer0_outputs(194) <= not b or a;
    layer0_outputs(195) <= '1';
    layer0_outputs(196) <= not b;
    layer0_outputs(197) <= not (a or b);
    layer0_outputs(198) <= a or b;
    layer0_outputs(199) <= a or b;
    layer0_outputs(200) <= not a or b;
    layer0_outputs(201) <= not (a or b);
    layer0_outputs(202) <= a;
    layer0_outputs(203) <= not (a or b);
    layer0_outputs(204) <= a or b;
    layer0_outputs(205) <= not a or b;
    layer0_outputs(206) <= not b or a;
    layer0_outputs(207) <= b;
    layer0_outputs(208) <= a;
    layer0_outputs(209) <= '1';
    layer0_outputs(210) <= a or b;
    layer0_outputs(211) <= a and not b;
    layer0_outputs(212) <= a and not b;
    layer0_outputs(213) <= not (a xor b);
    layer0_outputs(214) <= not b;
    layer0_outputs(215) <= a xor b;
    layer0_outputs(216) <= not (a or b);
    layer0_outputs(217) <= a;
    layer0_outputs(218) <= not (a or b);
    layer0_outputs(219) <= not a;
    layer0_outputs(220) <= a or b;
    layer0_outputs(221) <= not (a xor b);
    layer0_outputs(222) <= not (a or b);
    layer0_outputs(223) <= not a;
    layer0_outputs(224) <= not a;
    layer0_outputs(225) <= a or b;
    layer0_outputs(226) <= a or b;
    layer0_outputs(227) <= not b;
    layer0_outputs(228) <= b;
    layer0_outputs(229) <= not a;
    layer0_outputs(230) <= b;
    layer0_outputs(231) <= a;
    layer0_outputs(232) <= not (a or b);
    layer0_outputs(233) <= not (a or b);
    layer0_outputs(234) <= a and not b;
    layer0_outputs(235) <= a or b;
    layer0_outputs(236) <= not (a or b);
    layer0_outputs(237) <= a;
    layer0_outputs(238) <= b;
    layer0_outputs(239) <= a and not b;
    layer0_outputs(240) <= a and not b;
    layer0_outputs(241) <= not a;
    layer0_outputs(242) <= a or b;
    layer0_outputs(243) <= b;
    layer0_outputs(244) <= a or b;
    layer0_outputs(245) <= not (a or b);
    layer0_outputs(246) <= b;
    layer0_outputs(247) <= a and not b;
    layer0_outputs(248) <= not (a or b);
    layer0_outputs(249) <= not (a xor b);
    layer0_outputs(250) <= not a;
    layer0_outputs(251) <= a xor b;
    layer0_outputs(252) <= not a or b;
    layer0_outputs(253) <= not b;
    layer0_outputs(254) <= a;
    layer0_outputs(255) <= not b;
    layer0_outputs(256) <= a xor b;
    layer0_outputs(257) <= not (a xor b);
    layer0_outputs(258) <= not b;
    layer0_outputs(259) <= not b;
    layer0_outputs(260) <= not b;
    layer0_outputs(261) <= not b or a;
    layer0_outputs(262) <= a;
    layer0_outputs(263) <= a;
    layer0_outputs(264) <= not (a and b);
    layer0_outputs(265) <= a or b;
    layer0_outputs(266) <= not (a and b);
    layer0_outputs(267) <= a and not b;
    layer0_outputs(268) <= not a or b;
    layer0_outputs(269) <= not a or b;
    layer0_outputs(270) <= not (a or b);
    layer0_outputs(271) <= not a;
    layer0_outputs(272) <= not b;
    layer0_outputs(273) <= a and not b;
    layer0_outputs(274) <= not (a xor b);
    layer0_outputs(275) <= not b or a;
    layer0_outputs(276) <= a;
    layer0_outputs(277) <= a and not b;
    layer0_outputs(278) <= not b;
    layer0_outputs(279) <= a or b;
    layer0_outputs(280) <= b and not a;
    layer0_outputs(281) <= a and not b;
    layer0_outputs(282) <= b and not a;
    layer0_outputs(283) <= a;
    layer0_outputs(284) <= a;
    layer0_outputs(285) <= a and not b;
    layer0_outputs(286) <= a xor b;
    layer0_outputs(287) <= a or b;
    layer0_outputs(288) <= not a or b;
    layer0_outputs(289) <= not b or a;
    layer0_outputs(290) <= a and not b;
    layer0_outputs(291) <= b and not a;
    layer0_outputs(292) <= a;
    layer0_outputs(293) <= a or b;
    layer0_outputs(294) <= not (a or b);
    layer0_outputs(295) <= not (a and b);
    layer0_outputs(296) <= not b;
    layer0_outputs(297) <= b and not a;
    layer0_outputs(298) <= not (a xor b);
    layer0_outputs(299) <= not b;
    layer0_outputs(300) <= a xor b;
    layer0_outputs(301) <= not (a or b);
    layer0_outputs(302) <= not b or a;
    layer0_outputs(303) <= a and not b;
    layer0_outputs(304) <= not (a or b);
    layer0_outputs(305) <= not a;
    layer0_outputs(306) <= not (a and b);
    layer0_outputs(307) <= a or b;
    layer0_outputs(308) <= not (a or b);
    layer0_outputs(309) <= '1';
    layer0_outputs(310) <= a or b;
    layer0_outputs(311) <= not (a or b);
    layer0_outputs(312) <= not b or a;
    layer0_outputs(313) <= a;
    layer0_outputs(314) <= not a or b;
    layer0_outputs(315) <= a or b;
    layer0_outputs(316) <= a or b;
    layer0_outputs(317) <= a or b;
    layer0_outputs(318) <= a;
    layer0_outputs(319) <= b;
    layer0_outputs(320) <= not (a xor b);
    layer0_outputs(321) <= '0';
    layer0_outputs(322) <= b and not a;
    layer0_outputs(323) <= a and b;
    layer0_outputs(324) <= not b or a;
    layer0_outputs(325) <= not (a or b);
    layer0_outputs(326) <= not a or b;
    layer0_outputs(327) <= a;
    layer0_outputs(328) <= a xor b;
    layer0_outputs(329) <= not a;
    layer0_outputs(330) <= a or b;
    layer0_outputs(331) <= not b or a;
    layer0_outputs(332) <= not a or b;
    layer0_outputs(333) <= not (a or b);
    layer0_outputs(334) <= a;
    layer0_outputs(335) <= not (a or b);
    layer0_outputs(336) <= not (a or b);
    layer0_outputs(337) <= not b;
    layer0_outputs(338) <= a xor b;
    layer0_outputs(339) <= a xor b;
    layer0_outputs(340) <= a or b;
    layer0_outputs(341) <= not (a or b);
    layer0_outputs(342) <= not (a or b);
    layer0_outputs(343) <= a xor b;
    layer0_outputs(344) <= b and not a;
    layer0_outputs(345) <= not (a or b);
    layer0_outputs(346) <= not (a or b);
    layer0_outputs(347) <= not (a or b);
    layer0_outputs(348) <= a;
    layer0_outputs(349) <= a and not b;
    layer0_outputs(350) <= not b;
    layer0_outputs(351) <= not (a or b);
    layer0_outputs(352) <= a or b;
    layer0_outputs(353) <= a or b;
    layer0_outputs(354) <= '0';
    layer0_outputs(355) <= not a or b;
    layer0_outputs(356) <= a or b;
    layer0_outputs(357) <= not a;
    layer0_outputs(358) <= b;
    layer0_outputs(359) <= not a;
    layer0_outputs(360) <= a xor b;
    layer0_outputs(361) <= not a or b;
    layer0_outputs(362) <= a or b;
    layer0_outputs(363) <= b and not a;
    layer0_outputs(364) <= a or b;
    layer0_outputs(365) <= '0';
    layer0_outputs(366) <= a or b;
    layer0_outputs(367) <= not (a xor b);
    layer0_outputs(368) <= a or b;
    layer0_outputs(369) <= a and b;
    layer0_outputs(370) <= a;
    layer0_outputs(371) <= a xor b;
    layer0_outputs(372) <= a or b;
    layer0_outputs(373) <= not (a xor b);
    layer0_outputs(374) <= a or b;
    layer0_outputs(375) <= not (a or b);
    layer0_outputs(376) <= not a;
    layer0_outputs(377) <= not (a or b);
    layer0_outputs(378) <= a xor b;
    layer0_outputs(379) <= not a;
    layer0_outputs(380) <= not b or a;
    layer0_outputs(381) <= not (a or b);
    layer0_outputs(382) <= not (a or b);
    layer0_outputs(383) <= not (a or b);
    layer0_outputs(384) <= not b or a;
    layer0_outputs(385) <= not b or a;
    layer0_outputs(386) <= a;
    layer0_outputs(387) <= a;
    layer0_outputs(388) <= a and not b;
    layer0_outputs(389) <= b;
    layer0_outputs(390) <= not (a xor b);
    layer0_outputs(391) <= not b or a;
    layer0_outputs(392) <= a xor b;
    layer0_outputs(393) <= b and not a;
    layer0_outputs(394) <= a or b;
    layer0_outputs(395) <= b and not a;
    layer0_outputs(396) <= not (a or b);
    layer0_outputs(397) <= a and b;
    layer0_outputs(398) <= not (a and b);
    layer0_outputs(399) <= b;
    layer0_outputs(400) <= not (a or b);
    layer0_outputs(401) <= a and not b;
    layer0_outputs(402) <= not b or a;
    layer0_outputs(403) <= not b;
    layer0_outputs(404) <= a xor b;
    layer0_outputs(405) <= not (a or b);
    layer0_outputs(406) <= b and not a;
    layer0_outputs(407) <= not a;
    layer0_outputs(408) <= not (a xor b);
    layer0_outputs(409) <= not a or b;
    layer0_outputs(410) <= a;
    layer0_outputs(411) <= not a or b;
    layer0_outputs(412) <= not a;
    layer0_outputs(413) <= a or b;
    layer0_outputs(414) <= a or b;
    layer0_outputs(415) <= not b or a;
    layer0_outputs(416) <= not b;
    layer0_outputs(417) <= not (a or b);
    layer0_outputs(418) <= not (a xor b);
    layer0_outputs(419) <= a or b;
    layer0_outputs(420) <= a and not b;
    layer0_outputs(421) <= a or b;
    layer0_outputs(422) <= not (a or b);
    layer0_outputs(423) <= not (a or b);
    layer0_outputs(424) <= not b;
    layer0_outputs(425) <= not (a and b);
    layer0_outputs(426) <= not b;
    layer0_outputs(427) <= a;
    layer0_outputs(428) <= not b;
    layer0_outputs(429) <= a and not b;
    layer0_outputs(430) <= not b or a;
    layer0_outputs(431) <= '0';
    layer0_outputs(432) <= a or b;
    layer0_outputs(433) <= b and not a;
    layer0_outputs(434) <= '1';
    layer0_outputs(435) <= not b;
    layer0_outputs(436) <= a xor b;
    layer0_outputs(437) <= a xor b;
    layer0_outputs(438) <= a;
    layer0_outputs(439) <= a xor b;
    layer0_outputs(440) <= a xor b;
    layer0_outputs(441) <= not (a or b);
    layer0_outputs(442) <= a or b;
    layer0_outputs(443) <= a or b;
    layer0_outputs(444) <= not (a xor b);
    layer0_outputs(445) <= not b or a;
    layer0_outputs(446) <= a;
    layer0_outputs(447) <= not (a and b);
    layer0_outputs(448) <= not (a and b);
    layer0_outputs(449) <= not b or a;
    layer0_outputs(450) <= not (a or b);
    layer0_outputs(451) <= b;
    layer0_outputs(452) <= b and not a;
    layer0_outputs(453) <= not (a and b);
    layer0_outputs(454) <= b and not a;
    layer0_outputs(455) <= not (a xor b);
    layer0_outputs(456) <= not a or b;
    layer0_outputs(457) <= a xor b;
    layer0_outputs(458) <= not a;
    layer0_outputs(459) <= not b or a;
    layer0_outputs(460) <= a or b;
    layer0_outputs(461) <= a and not b;
    layer0_outputs(462) <= not (a or b);
    layer0_outputs(463) <= not (a or b);
    layer0_outputs(464) <= not (a or b);
    layer0_outputs(465) <= not a or b;
    layer0_outputs(466) <= b and not a;
    layer0_outputs(467) <= a xor b;
    layer0_outputs(468) <= not a;
    layer0_outputs(469) <= not a or b;
    layer0_outputs(470) <= a or b;
    layer0_outputs(471) <= not b or a;
    layer0_outputs(472) <= a or b;
    layer0_outputs(473) <= not a or b;
    layer0_outputs(474) <= a or b;
    layer0_outputs(475) <= a or b;
    layer0_outputs(476) <= a and b;
    layer0_outputs(477) <= not (a or b);
    layer0_outputs(478) <= not a or b;
    layer0_outputs(479) <= not b or a;
    layer0_outputs(480) <= not (a xor b);
    layer0_outputs(481) <= a xor b;
    layer0_outputs(482) <= not a or b;
    layer0_outputs(483) <= not (a or b);
    layer0_outputs(484) <= not b;
    layer0_outputs(485) <= not (a xor b);
    layer0_outputs(486) <= a and not b;
    layer0_outputs(487) <= not (a xor b);
    layer0_outputs(488) <= '1';
    layer0_outputs(489) <= b;
    layer0_outputs(490) <= a;
    layer0_outputs(491) <= b and not a;
    layer0_outputs(492) <= a xor b;
    layer0_outputs(493) <= not (a or b);
    layer0_outputs(494) <= b;
    layer0_outputs(495) <= a and not b;
    layer0_outputs(496) <= b;
    layer0_outputs(497) <= '0';
    layer0_outputs(498) <= a and not b;
    layer0_outputs(499) <= b;
    layer0_outputs(500) <= a or b;
    layer0_outputs(501) <= not b;
    layer0_outputs(502) <= not (a or b);
    layer0_outputs(503) <= a xor b;
    layer0_outputs(504) <= not a;
    layer0_outputs(505) <= a xor b;
    layer0_outputs(506) <= a xor b;
    layer0_outputs(507) <= not b;
    layer0_outputs(508) <= b and not a;
    layer0_outputs(509) <= '1';
    layer0_outputs(510) <= not (a or b);
    layer0_outputs(511) <= not (a or b);
    layer0_outputs(512) <= b;
    layer0_outputs(513) <= not (a or b);
    layer0_outputs(514) <= a or b;
    layer0_outputs(515) <= not b;
    layer0_outputs(516) <= not (a or b);
    layer0_outputs(517) <= a or b;
    layer0_outputs(518) <= not b;
    layer0_outputs(519) <= a or b;
    layer0_outputs(520) <= a;
    layer0_outputs(521) <= not a or b;
    layer0_outputs(522) <= not b or a;
    layer0_outputs(523) <= a xor b;
    layer0_outputs(524) <= not a;
    layer0_outputs(525) <= b;
    layer0_outputs(526) <= a and not b;
    layer0_outputs(527) <= a xor b;
    layer0_outputs(528) <= not (a and b);
    layer0_outputs(529) <= a;
    layer0_outputs(530) <= '1';
    layer0_outputs(531) <= not (a xor b);
    layer0_outputs(532) <= a;
    layer0_outputs(533) <= b;
    layer0_outputs(534) <= not b or a;
    layer0_outputs(535) <= a;
    layer0_outputs(536) <= a and b;
    layer0_outputs(537) <= b and not a;
    layer0_outputs(538) <= not a;
    layer0_outputs(539) <= not a or b;
    layer0_outputs(540) <= not b or a;
    layer0_outputs(541) <= a;
    layer0_outputs(542) <= not (a or b);
    layer0_outputs(543) <= a or b;
    layer0_outputs(544) <= a;
    layer0_outputs(545) <= a xor b;
    layer0_outputs(546) <= a or b;
    layer0_outputs(547) <= not b;
    layer0_outputs(548) <= a xor b;
    layer0_outputs(549) <= b and not a;
    layer0_outputs(550) <= not (a or b);
    layer0_outputs(551) <= not (a or b);
    layer0_outputs(552) <= a or b;
    layer0_outputs(553) <= not a;
    layer0_outputs(554) <= a;
    layer0_outputs(555) <= not a;
    layer0_outputs(556) <= a or b;
    layer0_outputs(557) <= not a or b;
    layer0_outputs(558) <= a;
    layer0_outputs(559) <= b and not a;
    layer0_outputs(560) <= not (a or b);
    layer0_outputs(561) <= not (a or b);
    layer0_outputs(562) <= b;
    layer0_outputs(563) <= b;
    layer0_outputs(564) <= not b;
    layer0_outputs(565) <= a;
    layer0_outputs(566) <= not (a and b);
    layer0_outputs(567) <= a or b;
    layer0_outputs(568) <= not (a or b);
    layer0_outputs(569) <= not (a or b);
    layer0_outputs(570) <= b;
    layer0_outputs(571) <= not b;
    layer0_outputs(572) <= not (a or b);
    layer0_outputs(573) <= not (a xor b);
    layer0_outputs(574) <= not b;
    layer0_outputs(575) <= not (a or b);
    layer0_outputs(576) <= b and not a;
    layer0_outputs(577) <= b;
    layer0_outputs(578) <= b and not a;
    layer0_outputs(579) <= a and not b;
    layer0_outputs(580) <= a or b;
    layer0_outputs(581) <= b;
    layer0_outputs(582) <= not b;
    layer0_outputs(583) <= b and not a;
    layer0_outputs(584) <= not b or a;
    layer0_outputs(585) <= not b;
    layer0_outputs(586) <= b;
    layer0_outputs(587) <= b;
    layer0_outputs(588) <= not b;
    layer0_outputs(589) <= not (a or b);
    layer0_outputs(590) <= not (a or b);
    layer0_outputs(591) <= not b;
    layer0_outputs(592) <= a xor b;
    layer0_outputs(593) <= b;
    layer0_outputs(594) <= not a;
    layer0_outputs(595) <= not b or a;
    layer0_outputs(596) <= b;
    layer0_outputs(597) <= a or b;
    layer0_outputs(598) <= not (a or b);
    layer0_outputs(599) <= '0';
    layer0_outputs(600) <= a and not b;
    layer0_outputs(601) <= not (a and b);
    layer0_outputs(602) <= not (a and b);
    layer0_outputs(603) <= not (a xor b);
    layer0_outputs(604) <= a xor b;
    layer0_outputs(605) <= not b;
    layer0_outputs(606) <= not a;
    layer0_outputs(607) <= not b or a;
    layer0_outputs(608) <= not (a or b);
    layer0_outputs(609) <= a and b;
    layer0_outputs(610) <= not b or a;
    layer0_outputs(611) <= not b;
    layer0_outputs(612) <= a or b;
    layer0_outputs(613) <= '0';
    layer0_outputs(614) <= not (a or b);
    layer0_outputs(615) <= a;
    layer0_outputs(616) <= not b;
    layer0_outputs(617) <= a or b;
    layer0_outputs(618) <= a or b;
    layer0_outputs(619) <= not (a or b);
    layer0_outputs(620) <= a;
    layer0_outputs(621) <= not a or b;
    layer0_outputs(622) <= '1';
    layer0_outputs(623) <= not a or b;
    layer0_outputs(624) <= not a;
    layer0_outputs(625) <= not (a or b);
    layer0_outputs(626) <= not (a or b);
    layer0_outputs(627) <= not (a or b);
    layer0_outputs(628) <= not (a xor b);
    layer0_outputs(629) <= a;
    layer0_outputs(630) <= not b;
    layer0_outputs(631) <= not (a or b);
    layer0_outputs(632) <= '1';
    layer0_outputs(633) <= a or b;
    layer0_outputs(634) <= a xor b;
    layer0_outputs(635) <= a and not b;
    layer0_outputs(636) <= not (a or b);
    layer0_outputs(637) <= b;
    layer0_outputs(638) <= not b or a;
    layer0_outputs(639) <= not (a or b);
    layer0_outputs(640) <= a or b;
    layer0_outputs(641) <= a xor b;
    layer0_outputs(642) <= a or b;
    layer0_outputs(643) <= b and not a;
    layer0_outputs(644) <= b;
    layer0_outputs(645) <= not (a xor b);
    layer0_outputs(646) <= not b;
    layer0_outputs(647) <= a or b;
    layer0_outputs(648) <= a and b;
    layer0_outputs(649) <= b;
    layer0_outputs(650) <= not b;
    layer0_outputs(651) <= not a;
    layer0_outputs(652) <= not (a or b);
    layer0_outputs(653) <= b;
    layer0_outputs(654) <= a or b;
    layer0_outputs(655) <= b and not a;
    layer0_outputs(656) <= b;
    layer0_outputs(657) <= not a;
    layer0_outputs(658) <= not (a or b);
    layer0_outputs(659) <= not (a xor b);
    layer0_outputs(660) <= not b or a;
    layer0_outputs(661) <= a and not b;
    layer0_outputs(662) <= not (a xor b);
    layer0_outputs(663) <= b;
    layer0_outputs(664) <= a xor b;
    layer0_outputs(665) <= not b or a;
    layer0_outputs(666) <= b;
    layer0_outputs(667) <= not b or a;
    layer0_outputs(668) <= b;
    layer0_outputs(669) <= not (a or b);
    layer0_outputs(670) <= not (a or b);
    layer0_outputs(671) <= a or b;
    layer0_outputs(672) <= a;
    layer0_outputs(673) <= b;
    layer0_outputs(674) <= a or b;
    layer0_outputs(675) <= b;
    layer0_outputs(676) <= a xor b;
    layer0_outputs(677) <= not (a or b);
    layer0_outputs(678) <= not (a or b);
    layer0_outputs(679) <= not (a or b);
    layer0_outputs(680) <= not (a or b);
    layer0_outputs(681) <= b and not a;
    layer0_outputs(682) <= a and not b;
    layer0_outputs(683) <= a or b;
    layer0_outputs(684) <= not (a or b);
    layer0_outputs(685) <= a xor b;
    layer0_outputs(686) <= not a or b;
    layer0_outputs(687) <= a and not b;
    layer0_outputs(688) <= '1';
    layer0_outputs(689) <= not a or b;
    layer0_outputs(690) <= not (a xor b);
    layer0_outputs(691) <= not a or b;
    layer0_outputs(692) <= a and b;
    layer0_outputs(693) <= a;
    layer0_outputs(694) <= a;
    layer0_outputs(695) <= not (a or b);
    layer0_outputs(696) <= not a or b;
    layer0_outputs(697) <= a or b;
    layer0_outputs(698) <= a or b;
    layer0_outputs(699) <= a or b;
    layer0_outputs(700) <= not a;
    layer0_outputs(701) <= b;
    layer0_outputs(702) <= not (a xor b);
    layer0_outputs(703) <= a and b;
    layer0_outputs(704) <= a or b;
    layer0_outputs(705) <= not (a or b);
    layer0_outputs(706) <= a or b;
    layer0_outputs(707) <= b;
    layer0_outputs(708) <= not b or a;
    layer0_outputs(709) <= b and not a;
    layer0_outputs(710) <= not b;
    layer0_outputs(711) <= not a;
    layer0_outputs(712) <= a or b;
    layer0_outputs(713) <= not (a or b);
    layer0_outputs(714) <= b;
    layer0_outputs(715) <= not b;
    layer0_outputs(716) <= not (a xor b);
    layer0_outputs(717) <= a xor b;
    layer0_outputs(718) <= not (a or b);
    layer0_outputs(719) <= a and not b;
    layer0_outputs(720) <= a xor b;
    layer0_outputs(721) <= not (a or b);
    layer0_outputs(722) <= a;
    layer0_outputs(723) <= a;
    layer0_outputs(724) <= b and not a;
    layer0_outputs(725) <= not a;
    layer0_outputs(726) <= not (a and b);
    layer0_outputs(727) <= a or b;
    layer0_outputs(728) <= a and not b;
    layer0_outputs(729) <= not a or b;
    layer0_outputs(730) <= not (a xor b);
    layer0_outputs(731) <= a and not b;
    layer0_outputs(732) <= a and not b;
    layer0_outputs(733) <= a and not b;
    layer0_outputs(734) <= not (a or b);
    layer0_outputs(735) <= a or b;
    layer0_outputs(736) <= not (a or b);
    layer0_outputs(737) <= not (a or b);
    layer0_outputs(738) <= not (a and b);
    layer0_outputs(739) <= a;
    layer0_outputs(740) <= b and not a;
    layer0_outputs(741) <= a or b;
    layer0_outputs(742) <= a or b;
    layer0_outputs(743) <= a and not b;
    layer0_outputs(744) <= not b;
    layer0_outputs(745) <= a;
    layer0_outputs(746) <= not a;
    layer0_outputs(747) <= a and not b;
    layer0_outputs(748) <= not a or b;
    layer0_outputs(749) <= b and not a;
    layer0_outputs(750) <= '1';
    layer0_outputs(751) <= a and not b;
    layer0_outputs(752) <= a;
    layer0_outputs(753) <= not a or b;
    layer0_outputs(754) <= not (a or b);
    layer0_outputs(755) <= not (a xor b);
    layer0_outputs(756) <= not (a or b);
    layer0_outputs(757) <= a;
    layer0_outputs(758) <= a or b;
    layer0_outputs(759) <= not a or b;
    layer0_outputs(760) <= a or b;
    layer0_outputs(761) <= b and not a;
    layer0_outputs(762) <= '0';
    layer0_outputs(763) <= not (a or b);
    layer0_outputs(764) <= a xor b;
    layer0_outputs(765) <= a xor b;
    layer0_outputs(766) <= b and not a;
    layer0_outputs(767) <= not a or b;
    layer0_outputs(768) <= not (a xor b);
    layer0_outputs(769) <= a or b;
    layer0_outputs(770) <= a and not b;
    layer0_outputs(771) <= not b or a;
    layer0_outputs(772) <= '0';
    layer0_outputs(773) <= not (a xor b);
    layer0_outputs(774) <= not (a or b);
    layer0_outputs(775) <= not (a or b);
    layer0_outputs(776) <= not (a or b);
    layer0_outputs(777) <= not a;
    layer0_outputs(778) <= a or b;
    layer0_outputs(779) <= a;
    layer0_outputs(780) <= b;
    layer0_outputs(781) <= not (a xor b);
    layer0_outputs(782) <= not b;
    layer0_outputs(783) <= a;
    layer0_outputs(784) <= b and not a;
    layer0_outputs(785) <= not b or a;
    layer0_outputs(786) <= not a or b;
    layer0_outputs(787) <= not b or a;
    layer0_outputs(788) <= a;
    layer0_outputs(789) <= a and not b;
    layer0_outputs(790) <= b;
    layer0_outputs(791) <= not (a or b);
    layer0_outputs(792) <= not b or a;
    layer0_outputs(793) <= a and b;
    layer0_outputs(794) <= b and not a;
    layer0_outputs(795) <= not (a xor b);
    layer0_outputs(796) <= not b;
    layer0_outputs(797) <= a;
    layer0_outputs(798) <= not b;
    layer0_outputs(799) <= not a;
    layer0_outputs(800) <= not (a xor b);
    layer0_outputs(801) <= not (a or b);
    layer0_outputs(802) <= not b or a;
    layer0_outputs(803) <= not (a or b);
    layer0_outputs(804) <= a or b;
    layer0_outputs(805) <= not b or a;
    layer0_outputs(806) <= not b;
    layer0_outputs(807) <= not (a or b);
    layer0_outputs(808) <= a;
    layer0_outputs(809) <= b and not a;
    layer0_outputs(810) <= b;
    layer0_outputs(811) <= not b or a;
    layer0_outputs(812) <= b;
    layer0_outputs(813) <= a;
    layer0_outputs(814) <= a or b;
    layer0_outputs(815) <= not (a xor b);
    layer0_outputs(816) <= a and not b;
    layer0_outputs(817) <= a and b;
    layer0_outputs(818) <= a and not b;
    layer0_outputs(819) <= b;
    layer0_outputs(820) <= b;
    layer0_outputs(821) <= a or b;
    layer0_outputs(822) <= a and not b;
    layer0_outputs(823) <= not a or b;
    layer0_outputs(824) <= not b or a;
    layer0_outputs(825) <= a or b;
    layer0_outputs(826) <= a or b;
    layer0_outputs(827) <= not (a or b);
    layer0_outputs(828) <= a or b;
    layer0_outputs(829) <= not (a or b);
    layer0_outputs(830) <= a xor b;
    layer0_outputs(831) <= a or b;
    layer0_outputs(832) <= a;
    layer0_outputs(833) <= not (a or b);
    layer0_outputs(834) <= a or b;
    layer0_outputs(835) <= a and not b;
    layer0_outputs(836) <= not (a or b);
    layer0_outputs(837) <= not b or a;
    layer0_outputs(838) <= a and not b;
    layer0_outputs(839) <= not (a or b);
    layer0_outputs(840) <= not b or a;
    layer0_outputs(841) <= b;
    layer0_outputs(842) <= a xor b;
    layer0_outputs(843) <= not b or a;
    layer0_outputs(844) <= a or b;
    layer0_outputs(845) <= b;
    layer0_outputs(846) <= not b;
    layer0_outputs(847) <= b;
    layer0_outputs(848) <= not b;
    layer0_outputs(849) <= not (a xor b);
    layer0_outputs(850) <= not (a xor b);
    layer0_outputs(851) <= not (a xor b);
    layer0_outputs(852) <= a and not b;
    layer0_outputs(853) <= a;
    layer0_outputs(854) <= not a;
    layer0_outputs(855) <= b and not a;
    layer0_outputs(856) <= a or b;
    layer0_outputs(857) <= not a;
    layer0_outputs(858) <= a;
    layer0_outputs(859) <= not a;
    layer0_outputs(860) <= b;
    layer0_outputs(861) <= not a or b;
    layer0_outputs(862) <= b and not a;
    layer0_outputs(863) <= a or b;
    layer0_outputs(864) <= a xor b;
    layer0_outputs(865) <= a or b;
    layer0_outputs(866) <= not a;
    layer0_outputs(867) <= b;
    layer0_outputs(868) <= a;
    layer0_outputs(869) <= a or b;
    layer0_outputs(870) <= a xor b;
    layer0_outputs(871) <= not (a or b);
    layer0_outputs(872) <= not a;
    layer0_outputs(873) <= a or b;
    layer0_outputs(874) <= a and not b;
    layer0_outputs(875) <= not b;
    layer0_outputs(876) <= a or b;
    layer0_outputs(877) <= a or b;
    layer0_outputs(878) <= a;
    layer0_outputs(879) <= not (a or b);
    layer0_outputs(880) <= a;
    layer0_outputs(881) <= not a;
    layer0_outputs(882) <= '0';
    layer0_outputs(883) <= a or b;
    layer0_outputs(884) <= not (a xor b);
    layer0_outputs(885) <= a and not b;
    layer0_outputs(886) <= a and not b;
    layer0_outputs(887) <= a or b;
    layer0_outputs(888) <= not (a or b);
    layer0_outputs(889) <= a and not b;
    layer0_outputs(890) <= not a;
    layer0_outputs(891) <= a or b;
    layer0_outputs(892) <= not (a xor b);
    layer0_outputs(893) <= not (a xor b);
    layer0_outputs(894) <= a;
    layer0_outputs(895) <= not (a or b);
    layer0_outputs(896) <= a or b;
    layer0_outputs(897) <= a;
    layer0_outputs(898) <= b and not a;
    layer0_outputs(899) <= not b or a;
    layer0_outputs(900) <= a xor b;
    layer0_outputs(901) <= a xor b;
    layer0_outputs(902) <= not (a or b);
    layer0_outputs(903) <= a or b;
    layer0_outputs(904) <= not a;
    layer0_outputs(905) <= a or b;
    layer0_outputs(906) <= a and b;
    layer0_outputs(907) <= a or b;
    layer0_outputs(908) <= not b or a;
    layer0_outputs(909) <= a xor b;
    layer0_outputs(910) <= not b or a;
    layer0_outputs(911) <= not a or b;
    layer0_outputs(912) <= not b;
    layer0_outputs(913) <= not (a or b);
    layer0_outputs(914) <= a;
    layer0_outputs(915) <= not a or b;
    layer0_outputs(916) <= not a or b;
    layer0_outputs(917) <= a;
    layer0_outputs(918) <= a;
    layer0_outputs(919) <= b and not a;
    layer0_outputs(920) <= not b;
    layer0_outputs(921) <= a and not b;
    layer0_outputs(922) <= b;
    layer0_outputs(923) <= b;
    layer0_outputs(924) <= a xor b;
    layer0_outputs(925) <= not (a xor b);
    layer0_outputs(926) <= not (a or b);
    layer0_outputs(927) <= not (a or b);
    layer0_outputs(928) <= b;
    layer0_outputs(929) <= not (a xor b);
    layer0_outputs(930) <= b and not a;
    layer0_outputs(931) <= a or b;
    layer0_outputs(932) <= b and not a;
    layer0_outputs(933) <= not (a or b);
    layer0_outputs(934) <= not (a xor b);
    layer0_outputs(935) <= not b;
    layer0_outputs(936) <= not a;
    layer0_outputs(937) <= not a;
    layer0_outputs(938) <= b and not a;
    layer0_outputs(939) <= b and not a;
    layer0_outputs(940) <= not (a or b);
    layer0_outputs(941) <= not (a or b);
    layer0_outputs(942) <= a;
    layer0_outputs(943) <= not a;
    layer0_outputs(944) <= not b or a;
    layer0_outputs(945) <= not a or b;
    layer0_outputs(946) <= a or b;
    layer0_outputs(947) <= b and not a;
    layer0_outputs(948) <= not a or b;
    layer0_outputs(949) <= a and b;
    layer0_outputs(950) <= not (a or b);
    layer0_outputs(951) <= a xor b;
    layer0_outputs(952) <= not a or b;
    layer0_outputs(953) <= a and b;
    layer0_outputs(954) <= not (a or b);
    layer0_outputs(955) <= a;
    layer0_outputs(956) <= '1';
    layer0_outputs(957) <= not (a or b);
    layer0_outputs(958) <= a;
    layer0_outputs(959) <= b and not a;
    layer0_outputs(960) <= b and not a;
    layer0_outputs(961) <= b and not a;
    layer0_outputs(962) <= '1';
    layer0_outputs(963) <= not a;
    layer0_outputs(964) <= not (a or b);
    layer0_outputs(965) <= a or b;
    layer0_outputs(966) <= b and not a;
    layer0_outputs(967) <= a or b;
    layer0_outputs(968) <= a and not b;
    layer0_outputs(969) <= not (a and b);
    layer0_outputs(970) <= not a or b;
    layer0_outputs(971) <= not a;
    layer0_outputs(972) <= a xor b;
    layer0_outputs(973) <= not (a or b);
    layer0_outputs(974) <= not b or a;
    layer0_outputs(975) <= not (a or b);
    layer0_outputs(976) <= not b or a;
    layer0_outputs(977) <= not (a xor b);
    layer0_outputs(978) <= not a or b;
    layer0_outputs(979) <= not b;
    layer0_outputs(980) <= b and not a;
    layer0_outputs(981) <= not a;
    layer0_outputs(982) <= a or b;
    layer0_outputs(983) <= not (a or b);
    layer0_outputs(984) <= not (a or b);
    layer0_outputs(985) <= not (a or b);
    layer0_outputs(986) <= b;
    layer0_outputs(987) <= not a or b;
    layer0_outputs(988) <= a or b;
    layer0_outputs(989) <= not (a xor b);
    layer0_outputs(990) <= not a;
    layer0_outputs(991) <= not (a xor b);
    layer0_outputs(992) <= b and not a;
    layer0_outputs(993) <= not b or a;
    layer0_outputs(994) <= not (a or b);
    layer0_outputs(995) <= b and not a;
    layer0_outputs(996) <= not (a xor b);
    layer0_outputs(997) <= a or b;
    layer0_outputs(998) <= not b;
    layer0_outputs(999) <= not b or a;
    layer0_outputs(1000) <= not a;
    layer0_outputs(1001) <= not (a or b);
    layer0_outputs(1002) <= not a;
    layer0_outputs(1003) <= b and not a;
    layer0_outputs(1004) <= a or b;
    layer0_outputs(1005) <= b;
    layer0_outputs(1006) <= a or b;
    layer0_outputs(1007) <= not b;
    layer0_outputs(1008) <= b;
    layer0_outputs(1009) <= not (a xor b);
    layer0_outputs(1010) <= b and not a;
    layer0_outputs(1011) <= b;
    layer0_outputs(1012) <= not a or b;
    layer0_outputs(1013) <= a;
    layer0_outputs(1014) <= not (a or b);
    layer0_outputs(1015) <= not a;
    layer0_outputs(1016) <= a or b;
    layer0_outputs(1017) <= not a or b;
    layer0_outputs(1018) <= a and not b;
    layer0_outputs(1019) <= '0';
    layer0_outputs(1020) <= b and not a;
    layer0_outputs(1021) <= not (a or b);
    layer0_outputs(1022) <= not (a or b);
    layer0_outputs(1023) <= a xor b;
    layer0_outputs(1024) <= a xor b;
    layer0_outputs(1025) <= not b;
    layer0_outputs(1026) <= a and b;
    layer0_outputs(1027) <= a or b;
    layer0_outputs(1028) <= a xor b;
    layer0_outputs(1029) <= not (a xor b);
    layer0_outputs(1030) <= a or b;
    layer0_outputs(1031) <= not a;
    layer0_outputs(1032) <= a and not b;
    layer0_outputs(1033) <= a or b;
    layer0_outputs(1034) <= a and not b;
    layer0_outputs(1035) <= not (a or b);
    layer0_outputs(1036) <= a xor b;
    layer0_outputs(1037) <= a xor b;
    layer0_outputs(1038) <= '0';
    layer0_outputs(1039) <= a and b;
    layer0_outputs(1040) <= a or b;
    layer0_outputs(1041) <= not (a or b);
    layer0_outputs(1042) <= a xor b;
    layer0_outputs(1043) <= a or b;
    layer0_outputs(1044) <= a and not b;
    layer0_outputs(1045) <= a and not b;
    layer0_outputs(1046) <= not a;
    layer0_outputs(1047) <= not a or b;
    layer0_outputs(1048) <= not a or b;
    layer0_outputs(1049) <= not (a xor b);
    layer0_outputs(1050) <= not (a or b);
    layer0_outputs(1051) <= not (a xor b);
    layer0_outputs(1052) <= not (a or b);
    layer0_outputs(1053) <= a or b;
    layer0_outputs(1054) <= not (a or b);
    layer0_outputs(1055) <= not a;
    layer0_outputs(1056) <= not (a or b);
    layer0_outputs(1057) <= b;
    layer0_outputs(1058) <= a or b;
    layer0_outputs(1059) <= not b;
    layer0_outputs(1060) <= a or b;
    layer0_outputs(1061) <= not (a or b);
    layer0_outputs(1062) <= not a or b;
    layer0_outputs(1063) <= a or b;
    layer0_outputs(1064) <= '0';
    layer0_outputs(1065) <= not b or a;
    layer0_outputs(1066) <= not b;
    layer0_outputs(1067) <= not b or a;
    layer0_outputs(1068) <= a or b;
    layer0_outputs(1069) <= not a;
    layer0_outputs(1070) <= a and b;
    layer0_outputs(1071) <= not b or a;
    layer0_outputs(1072) <= not (a or b);
    layer0_outputs(1073) <= a;
    layer0_outputs(1074) <= a or b;
    layer0_outputs(1075) <= not b;
    layer0_outputs(1076) <= not (a or b);
    layer0_outputs(1077) <= b;
    layer0_outputs(1078) <= b;
    layer0_outputs(1079) <= a xor b;
    layer0_outputs(1080) <= not a;
    layer0_outputs(1081) <= a xor b;
    layer0_outputs(1082) <= a or b;
    layer0_outputs(1083) <= a and not b;
    layer0_outputs(1084) <= a;
    layer0_outputs(1085) <= a or b;
    layer0_outputs(1086) <= not a;
    layer0_outputs(1087) <= b;
    layer0_outputs(1088) <= b;
    layer0_outputs(1089) <= a or b;
    layer0_outputs(1090) <= a or b;
    layer0_outputs(1091) <= not (a and b);
    layer0_outputs(1092) <= not a or b;
    layer0_outputs(1093) <= a xor b;
    layer0_outputs(1094) <= a or b;
    layer0_outputs(1095) <= '1';
    layer0_outputs(1096) <= b;
    layer0_outputs(1097) <= a or b;
    layer0_outputs(1098) <= not a;
    layer0_outputs(1099) <= not (a xor b);
    layer0_outputs(1100) <= b;
    layer0_outputs(1101) <= not a;
    layer0_outputs(1102) <= a and b;
    layer0_outputs(1103) <= b;
    layer0_outputs(1104) <= b and not a;
    layer0_outputs(1105) <= b and not a;
    layer0_outputs(1106) <= a;
    layer0_outputs(1107) <= '1';
    layer0_outputs(1108) <= not a;
    layer0_outputs(1109) <= not b;
    layer0_outputs(1110) <= a and not b;
    layer0_outputs(1111) <= not (a and b);
    layer0_outputs(1112) <= a or b;
    layer0_outputs(1113) <= not b or a;
    layer0_outputs(1114) <= a or b;
    layer0_outputs(1115) <= a;
    layer0_outputs(1116) <= not a or b;
    layer0_outputs(1117) <= not a or b;
    layer0_outputs(1118) <= a and not b;
    layer0_outputs(1119) <= b;
    layer0_outputs(1120) <= not b;
    layer0_outputs(1121) <= not (a or b);
    layer0_outputs(1122) <= a or b;
    layer0_outputs(1123) <= a xor b;
    layer0_outputs(1124) <= not (a or b);
    layer0_outputs(1125) <= b and not a;
    layer0_outputs(1126) <= a;
    layer0_outputs(1127) <= not (a xor b);
    layer0_outputs(1128) <= b;
    layer0_outputs(1129) <= not (a xor b);
    layer0_outputs(1130) <= a xor b;
    layer0_outputs(1131) <= b;
    layer0_outputs(1132) <= a xor b;
    layer0_outputs(1133) <= a or b;
    layer0_outputs(1134) <= not b or a;
    layer0_outputs(1135) <= not b;
    layer0_outputs(1136) <= a xor b;
    layer0_outputs(1137) <= not (a xor b);
    layer0_outputs(1138) <= not (a xor b);
    layer0_outputs(1139) <= a and not b;
    layer0_outputs(1140) <= not (a or b);
    layer0_outputs(1141) <= a;
    layer0_outputs(1142) <= b and not a;
    layer0_outputs(1143) <= not b;
    layer0_outputs(1144) <= not (a or b);
    layer0_outputs(1145) <= a xor b;
    layer0_outputs(1146) <= '0';
    layer0_outputs(1147) <= not b or a;
    layer0_outputs(1148) <= a or b;
    layer0_outputs(1149) <= not a or b;
    layer0_outputs(1150) <= b and not a;
    layer0_outputs(1151) <= a xor b;
    layer0_outputs(1152) <= not b;
    layer0_outputs(1153) <= a xor b;
    layer0_outputs(1154) <= b;
    layer0_outputs(1155) <= a;
    layer0_outputs(1156) <= a;
    layer0_outputs(1157) <= not (a or b);
    layer0_outputs(1158) <= not (a or b);
    layer0_outputs(1159) <= not (a or b);
    layer0_outputs(1160) <= a or b;
    layer0_outputs(1161) <= not (a xor b);
    layer0_outputs(1162) <= b and not a;
    layer0_outputs(1163) <= a or b;
    layer0_outputs(1164) <= not a;
    layer0_outputs(1165) <= a;
    layer0_outputs(1166) <= not (a and b);
    layer0_outputs(1167) <= a or b;
    layer0_outputs(1168) <= not (a and b);
    layer0_outputs(1169) <= not (a or b);
    layer0_outputs(1170) <= not b;
    layer0_outputs(1171) <= a or b;
    layer0_outputs(1172) <= b and not a;
    layer0_outputs(1173) <= b;
    layer0_outputs(1174) <= not b or a;
    layer0_outputs(1175) <= a and not b;
    layer0_outputs(1176) <= a or b;
    layer0_outputs(1177) <= a and not b;
    layer0_outputs(1178) <= b and not a;
    layer0_outputs(1179) <= not (a xor b);
    layer0_outputs(1180) <= not (a xor b);
    layer0_outputs(1181) <= not a or b;
    layer0_outputs(1182) <= a xor b;
    layer0_outputs(1183) <= a xor b;
    layer0_outputs(1184) <= a or b;
    layer0_outputs(1185) <= not b or a;
    layer0_outputs(1186) <= a or b;
    layer0_outputs(1187) <= not (a or b);
    layer0_outputs(1188) <= not (a or b);
    layer0_outputs(1189) <= b and not a;
    layer0_outputs(1190) <= a;
    layer0_outputs(1191) <= a xor b;
    layer0_outputs(1192) <= a xor b;
    layer0_outputs(1193) <= a and not b;
    layer0_outputs(1194) <= not (a or b);
    layer0_outputs(1195) <= a and b;
    layer0_outputs(1196) <= not (a xor b);
    layer0_outputs(1197) <= b;
    layer0_outputs(1198) <= not (a xor b);
    layer0_outputs(1199) <= not (a or b);
    layer0_outputs(1200) <= not b;
    layer0_outputs(1201) <= '1';
    layer0_outputs(1202) <= a or b;
    layer0_outputs(1203) <= a or b;
    layer0_outputs(1204) <= not a;
    layer0_outputs(1205) <= a;
    layer0_outputs(1206) <= a;
    layer0_outputs(1207) <= a or b;
    layer0_outputs(1208) <= b and not a;
    layer0_outputs(1209) <= not (a and b);
    layer0_outputs(1210) <= not (a or b);
    layer0_outputs(1211) <= b;
    layer0_outputs(1212) <= not a;
    layer0_outputs(1213) <= a and not b;
    layer0_outputs(1214) <= '1';
    layer0_outputs(1215) <= not (a xor b);
    layer0_outputs(1216) <= b;
    layer0_outputs(1217) <= not b;
    layer0_outputs(1218) <= '0';
    layer0_outputs(1219) <= a or b;
    layer0_outputs(1220) <= a and not b;
    layer0_outputs(1221) <= a or b;
    layer0_outputs(1222) <= not (a or b);
    layer0_outputs(1223) <= not (a or b);
    layer0_outputs(1224) <= not (a and b);
    layer0_outputs(1225) <= not (a xor b);
    layer0_outputs(1226) <= not (a and b);
    layer0_outputs(1227) <= a or b;
    layer0_outputs(1228) <= not a or b;
    layer0_outputs(1229) <= not a;
    layer0_outputs(1230) <= not (a or b);
    layer0_outputs(1231) <= not (a or b);
    layer0_outputs(1232) <= not b or a;
    layer0_outputs(1233) <= not (a or b);
    layer0_outputs(1234) <= a or b;
    layer0_outputs(1235) <= not (a or b);
    layer0_outputs(1236) <= b;
    layer0_outputs(1237) <= b and not a;
    layer0_outputs(1238) <= not a;
    layer0_outputs(1239) <= not (a or b);
    layer0_outputs(1240) <= not b;
    layer0_outputs(1241) <= a;
    layer0_outputs(1242) <= a or b;
    layer0_outputs(1243) <= not a or b;
    layer0_outputs(1244) <= a or b;
    layer0_outputs(1245) <= a or b;
    layer0_outputs(1246) <= '1';
    layer0_outputs(1247) <= '1';
    layer0_outputs(1248) <= not (a or b);
    layer0_outputs(1249) <= a and not b;
    layer0_outputs(1250) <= b;
    layer0_outputs(1251) <= b and not a;
    layer0_outputs(1252) <= not (a or b);
    layer0_outputs(1253) <= not a or b;
    layer0_outputs(1254) <= not (a and b);
    layer0_outputs(1255) <= a or b;
    layer0_outputs(1256) <= b;
    layer0_outputs(1257) <= a xor b;
    layer0_outputs(1258) <= a or b;
    layer0_outputs(1259) <= not (a xor b);
    layer0_outputs(1260) <= b;
    layer0_outputs(1261) <= not (a or b);
    layer0_outputs(1262) <= not a;
    layer0_outputs(1263) <= not (a or b);
    layer0_outputs(1264) <= a and not b;
    layer0_outputs(1265) <= a or b;
    layer0_outputs(1266) <= not a;
    layer0_outputs(1267) <= not (a or b);
    layer0_outputs(1268) <= not (a xor b);
    layer0_outputs(1269) <= a xor b;
    layer0_outputs(1270) <= not b or a;
    layer0_outputs(1271) <= a and not b;
    layer0_outputs(1272) <= b and not a;
    layer0_outputs(1273) <= '0';
    layer0_outputs(1274) <= a and b;
    layer0_outputs(1275) <= a;
    layer0_outputs(1276) <= a or b;
    layer0_outputs(1277) <= a or b;
    layer0_outputs(1278) <= a xor b;
    layer0_outputs(1279) <= '0';
    layer0_outputs(1280) <= not (a or b);
    layer0_outputs(1281) <= not b;
    layer0_outputs(1282) <= not a or b;
    layer0_outputs(1283) <= not b;
    layer0_outputs(1284) <= not b;
    layer0_outputs(1285) <= not a or b;
    layer0_outputs(1286) <= not (a or b);
    layer0_outputs(1287) <= a or b;
    layer0_outputs(1288) <= not (a xor b);
    layer0_outputs(1289) <= b and not a;
    layer0_outputs(1290) <= not (a or b);
    layer0_outputs(1291) <= not b or a;
    layer0_outputs(1292) <= a;
    layer0_outputs(1293) <= a or b;
    layer0_outputs(1294) <= not a or b;
    layer0_outputs(1295) <= not a or b;
    layer0_outputs(1296) <= not b or a;
    layer0_outputs(1297) <= a xor b;
    layer0_outputs(1298) <= not (a and b);
    layer0_outputs(1299) <= a and not b;
    layer0_outputs(1300) <= not (a or b);
    layer0_outputs(1301) <= not (a xor b);
    layer0_outputs(1302) <= not (a xor b);
    layer0_outputs(1303) <= not (a or b);
    layer0_outputs(1304) <= not (a xor b);
    layer0_outputs(1305) <= not a;
    layer0_outputs(1306) <= a or b;
    layer0_outputs(1307) <= a or b;
    layer0_outputs(1308) <= a;
    layer0_outputs(1309) <= a or b;
    layer0_outputs(1310) <= a xor b;
    layer0_outputs(1311) <= not b;
    layer0_outputs(1312) <= not (a or b);
    layer0_outputs(1313) <= b and not a;
    layer0_outputs(1314) <= not b;
    layer0_outputs(1315) <= not (a xor b);
    layer0_outputs(1316) <= a or b;
    layer0_outputs(1317) <= a xor b;
    layer0_outputs(1318) <= a and b;
    layer0_outputs(1319) <= not a;
    layer0_outputs(1320) <= b;
    layer0_outputs(1321) <= a and not b;
    layer0_outputs(1322) <= not (a xor b);
    layer0_outputs(1323) <= a xor b;
    layer0_outputs(1324) <= not a;
    layer0_outputs(1325) <= '1';
    layer0_outputs(1326) <= b and not a;
    layer0_outputs(1327) <= a or b;
    layer0_outputs(1328) <= not a or b;
    layer0_outputs(1329) <= not b or a;
    layer0_outputs(1330) <= b;
    layer0_outputs(1331) <= not b or a;
    layer0_outputs(1332) <= a xor b;
    layer0_outputs(1333) <= a and b;
    layer0_outputs(1334) <= not (a or b);
    layer0_outputs(1335) <= not a or b;
    layer0_outputs(1336) <= a xor b;
    layer0_outputs(1337) <= not b or a;
    layer0_outputs(1338) <= not b or a;
    layer0_outputs(1339) <= not (a or b);
    layer0_outputs(1340) <= not (a or b);
    layer0_outputs(1341) <= not (a or b);
    layer0_outputs(1342) <= a or b;
    layer0_outputs(1343) <= a and not b;
    layer0_outputs(1344) <= not b or a;
    layer0_outputs(1345) <= not (a or b);
    layer0_outputs(1346) <= not (a xor b);
    layer0_outputs(1347) <= b;
    layer0_outputs(1348) <= not (a or b);
    layer0_outputs(1349) <= not (a or b);
    layer0_outputs(1350) <= b;
    layer0_outputs(1351) <= a;
    layer0_outputs(1352) <= a or b;
    layer0_outputs(1353) <= a or b;
    layer0_outputs(1354) <= a or b;
    layer0_outputs(1355) <= a;
    layer0_outputs(1356) <= a or b;
    layer0_outputs(1357) <= b;
    layer0_outputs(1358) <= not b;
    layer0_outputs(1359) <= a and b;
    layer0_outputs(1360) <= a or b;
    layer0_outputs(1361) <= not a or b;
    layer0_outputs(1362) <= not (a xor b);
    layer0_outputs(1363) <= a;
    layer0_outputs(1364) <= not b or a;
    layer0_outputs(1365) <= not (a or b);
    layer0_outputs(1366) <= a and not b;
    layer0_outputs(1367) <= not (a xor b);
    layer0_outputs(1368) <= '0';
    layer0_outputs(1369) <= b and not a;
    layer0_outputs(1370) <= not a or b;
    layer0_outputs(1371) <= not (a or b);
    layer0_outputs(1372) <= not a;
    layer0_outputs(1373) <= not a;
    layer0_outputs(1374) <= a or b;
    layer0_outputs(1375) <= a or b;
    layer0_outputs(1376) <= not b or a;
    layer0_outputs(1377) <= not (a or b);
    layer0_outputs(1378) <= a xor b;
    layer0_outputs(1379) <= '1';
    layer0_outputs(1380) <= not b or a;
    layer0_outputs(1381) <= '0';
    layer0_outputs(1382) <= b;
    layer0_outputs(1383) <= b and not a;
    layer0_outputs(1384) <= not a or b;
    layer0_outputs(1385) <= a or b;
    layer0_outputs(1386) <= '0';
    layer0_outputs(1387) <= a;
    layer0_outputs(1388) <= not a or b;
    layer0_outputs(1389) <= b and not a;
    layer0_outputs(1390) <= a or b;
    layer0_outputs(1391) <= not (a xor b);
    layer0_outputs(1392) <= not a or b;
    layer0_outputs(1393) <= not b;
    layer0_outputs(1394) <= not (a or b);
    layer0_outputs(1395) <= b and not a;
    layer0_outputs(1396) <= not (a xor b);
    layer0_outputs(1397) <= a xor b;
    layer0_outputs(1398) <= not (a or b);
    layer0_outputs(1399) <= not (a or b);
    layer0_outputs(1400) <= not (a xor b);
    layer0_outputs(1401) <= not b;
    layer0_outputs(1402) <= not (a xor b);
    layer0_outputs(1403) <= not (a or b);
    layer0_outputs(1404) <= a or b;
    layer0_outputs(1405) <= not (a xor b);
    layer0_outputs(1406) <= not b;
    layer0_outputs(1407) <= not (a xor b);
    layer0_outputs(1408) <= not (a or b);
    layer0_outputs(1409) <= a xor b;
    layer0_outputs(1410) <= a;
    layer0_outputs(1411) <= b;
    layer0_outputs(1412) <= b and not a;
    layer0_outputs(1413) <= b;
    layer0_outputs(1414) <= not a or b;
    layer0_outputs(1415) <= not (a and b);
    layer0_outputs(1416) <= not (a or b);
    layer0_outputs(1417) <= not a;
    layer0_outputs(1418) <= not a or b;
    layer0_outputs(1419) <= not (a or b);
    layer0_outputs(1420) <= b;
    layer0_outputs(1421) <= a xor b;
    layer0_outputs(1422) <= not (a xor b);
    layer0_outputs(1423) <= not (a and b);
    layer0_outputs(1424) <= a xor b;
    layer0_outputs(1425) <= a or b;
    layer0_outputs(1426) <= not (a or b);
    layer0_outputs(1427) <= a or b;
    layer0_outputs(1428) <= not b or a;
    layer0_outputs(1429) <= not (a xor b);
    layer0_outputs(1430) <= not (a or b);
    layer0_outputs(1431) <= a and not b;
    layer0_outputs(1432) <= a;
    layer0_outputs(1433) <= a and not b;
    layer0_outputs(1434) <= not b;
    layer0_outputs(1435) <= not a or b;
    layer0_outputs(1436) <= not b or a;
    layer0_outputs(1437) <= b;
    layer0_outputs(1438) <= not b;
    layer0_outputs(1439) <= not (a or b);
    layer0_outputs(1440) <= a or b;
    layer0_outputs(1441) <= not (a or b);
    layer0_outputs(1442) <= a and b;
    layer0_outputs(1443) <= not b;
    layer0_outputs(1444) <= not (a or b);
    layer0_outputs(1445) <= a and b;
    layer0_outputs(1446) <= a xor b;
    layer0_outputs(1447) <= a;
    layer0_outputs(1448) <= not (a or b);
    layer0_outputs(1449) <= a and b;
    layer0_outputs(1450) <= not (a xor b);
    layer0_outputs(1451) <= not (a xor b);
    layer0_outputs(1452) <= not b;
    layer0_outputs(1453) <= not (a or b);
    layer0_outputs(1454) <= '0';
    layer0_outputs(1455) <= a or b;
    layer0_outputs(1456) <= not b or a;
    layer0_outputs(1457) <= not b;
    layer0_outputs(1458) <= b;
    layer0_outputs(1459) <= not (a or b);
    layer0_outputs(1460) <= a or b;
    layer0_outputs(1461) <= a;
    layer0_outputs(1462) <= b and not a;
    layer0_outputs(1463) <= a or b;
    layer0_outputs(1464) <= a or b;
    layer0_outputs(1465) <= a;
    layer0_outputs(1466) <= a xor b;
    layer0_outputs(1467) <= a or b;
    layer0_outputs(1468) <= not (a or b);
    layer0_outputs(1469) <= a or b;
    layer0_outputs(1470) <= a or b;
    layer0_outputs(1471) <= a and not b;
    layer0_outputs(1472) <= a or b;
    layer0_outputs(1473) <= not (a or b);
    layer0_outputs(1474) <= not b or a;
    layer0_outputs(1475) <= a or b;
    layer0_outputs(1476) <= not (a xor b);
    layer0_outputs(1477) <= not (a xor b);
    layer0_outputs(1478) <= b;
    layer0_outputs(1479) <= a and not b;
    layer0_outputs(1480) <= not a or b;
    layer0_outputs(1481) <= '0';
    layer0_outputs(1482) <= '1';
    layer0_outputs(1483) <= '1';
    layer0_outputs(1484) <= b and not a;
    layer0_outputs(1485) <= not (a or b);
    layer0_outputs(1486) <= not (a or b);
    layer0_outputs(1487) <= a xor b;
    layer0_outputs(1488) <= b;
    layer0_outputs(1489) <= a or b;
    layer0_outputs(1490) <= a or b;
    layer0_outputs(1491) <= not (a or b);
    layer0_outputs(1492) <= a or b;
    layer0_outputs(1493) <= '1';
    layer0_outputs(1494) <= b and not a;
    layer0_outputs(1495) <= not (a xor b);
    layer0_outputs(1496) <= not a or b;
    layer0_outputs(1497) <= a or b;
    layer0_outputs(1498) <= not (a or b);
    layer0_outputs(1499) <= a and not b;
    layer0_outputs(1500) <= a xor b;
    layer0_outputs(1501) <= b and not a;
    layer0_outputs(1502) <= a xor b;
    layer0_outputs(1503) <= a or b;
    layer0_outputs(1504) <= a or b;
    layer0_outputs(1505) <= not (a or b);
    layer0_outputs(1506) <= a and not b;
    layer0_outputs(1507) <= not a or b;
    layer0_outputs(1508) <= not a or b;
    layer0_outputs(1509) <= a;
    layer0_outputs(1510) <= not (a or b);
    layer0_outputs(1511) <= a or b;
    layer0_outputs(1512) <= not (a or b);
    layer0_outputs(1513) <= a and not b;
    layer0_outputs(1514) <= not a or b;
    layer0_outputs(1515) <= not (a and b);
    layer0_outputs(1516) <= not a;
    layer0_outputs(1517) <= not a;
    layer0_outputs(1518) <= a or b;
    layer0_outputs(1519) <= not b;
    layer0_outputs(1520) <= b and not a;
    layer0_outputs(1521) <= not b or a;
    layer0_outputs(1522) <= a;
    layer0_outputs(1523) <= not (a or b);
    layer0_outputs(1524) <= b and not a;
    layer0_outputs(1525) <= a and b;
    layer0_outputs(1526) <= b and not a;
    layer0_outputs(1527) <= a and not b;
    layer0_outputs(1528) <= a;
    layer0_outputs(1529) <= a or b;
    layer0_outputs(1530) <= a xor b;
    layer0_outputs(1531) <= not a or b;
    layer0_outputs(1532) <= not a;
    layer0_outputs(1533) <= not a or b;
    layer0_outputs(1534) <= a or b;
    layer0_outputs(1535) <= not b;
    layer0_outputs(1536) <= not a or b;
    layer0_outputs(1537) <= not (a or b);
    layer0_outputs(1538) <= not (a or b);
    layer0_outputs(1539) <= not b or a;
    layer0_outputs(1540) <= not b;
    layer0_outputs(1541) <= a or b;
    layer0_outputs(1542) <= a or b;
    layer0_outputs(1543) <= a xor b;
    layer0_outputs(1544) <= a or b;
    layer0_outputs(1545) <= not a or b;
    layer0_outputs(1546) <= a or b;
    layer0_outputs(1547) <= a xor b;
    layer0_outputs(1548) <= a and not b;
    layer0_outputs(1549) <= b;
    layer0_outputs(1550) <= a or b;
    layer0_outputs(1551) <= a or b;
    layer0_outputs(1552) <= '0';
    layer0_outputs(1553) <= not (a xor b);
    layer0_outputs(1554) <= not (a xor b);
    layer0_outputs(1555) <= not b;
    layer0_outputs(1556) <= not b or a;
    layer0_outputs(1557) <= not (a or b);
    layer0_outputs(1558) <= not (a or b);
    layer0_outputs(1559) <= not a;
    layer0_outputs(1560) <= b and not a;
    layer0_outputs(1561) <= not (a or b);
    layer0_outputs(1562) <= a and not b;
    layer0_outputs(1563) <= a;
    layer0_outputs(1564) <= a or b;
    layer0_outputs(1565) <= not (a or b);
    layer0_outputs(1566) <= '1';
    layer0_outputs(1567) <= '1';
    layer0_outputs(1568) <= a;
    layer0_outputs(1569) <= a and not b;
    layer0_outputs(1570) <= a and not b;
    layer0_outputs(1571) <= not (a and b);
    layer0_outputs(1572) <= not b;
    layer0_outputs(1573) <= '1';
    layer0_outputs(1574) <= not a or b;
    layer0_outputs(1575) <= not (a or b);
    layer0_outputs(1576) <= a xor b;
    layer0_outputs(1577) <= a;
    layer0_outputs(1578) <= b;
    layer0_outputs(1579) <= not a or b;
    layer0_outputs(1580) <= a or b;
    layer0_outputs(1581) <= not (a xor b);
    layer0_outputs(1582) <= a xor b;
    layer0_outputs(1583) <= not b;
    layer0_outputs(1584) <= not a;
    layer0_outputs(1585) <= a or b;
    layer0_outputs(1586) <= not (a or b);
    layer0_outputs(1587) <= a;
    layer0_outputs(1588) <= not (a or b);
    layer0_outputs(1589) <= not b or a;
    layer0_outputs(1590) <= a or b;
    layer0_outputs(1591) <= a;
    layer0_outputs(1592) <= not a or b;
    layer0_outputs(1593) <= a and not b;
    layer0_outputs(1594) <= a or b;
    layer0_outputs(1595) <= a or b;
    layer0_outputs(1596) <= a;
    layer0_outputs(1597) <= a or b;
    layer0_outputs(1598) <= not (a xor b);
    layer0_outputs(1599) <= a and not b;
    layer0_outputs(1600) <= b and not a;
    layer0_outputs(1601) <= a and b;
    layer0_outputs(1602) <= not (a xor b);
    layer0_outputs(1603) <= not (a xor b);
    layer0_outputs(1604) <= a;
    layer0_outputs(1605) <= b;
    layer0_outputs(1606) <= a and not b;
    layer0_outputs(1607) <= b;
    layer0_outputs(1608) <= not (a or b);
    layer0_outputs(1609) <= b and not a;
    layer0_outputs(1610) <= a xor b;
    layer0_outputs(1611) <= not (a or b);
    layer0_outputs(1612) <= a xor b;
    layer0_outputs(1613) <= a xor b;
    layer0_outputs(1614) <= a and not b;
    layer0_outputs(1615) <= b and not a;
    layer0_outputs(1616) <= not (a or b);
    layer0_outputs(1617) <= not b;
    layer0_outputs(1618) <= not (a or b);
    layer0_outputs(1619) <= not (a or b);
    layer0_outputs(1620) <= not (a xor b);
    layer0_outputs(1621) <= not (a or b);
    layer0_outputs(1622) <= a xor b;
    layer0_outputs(1623) <= not (a or b);
    layer0_outputs(1624) <= '0';
    layer0_outputs(1625) <= not b or a;
    layer0_outputs(1626) <= a or b;
    layer0_outputs(1627) <= not (a xor b);
    layer0_outputs(1628) <= b;
    layer0_outputs(1629) <= a;
    layer0_outputs(1630) <= not (a or b);
    layer0_outputs(1631) <= a and not b;
    layer0_outputs(1632) <= a xor b;
    layer0_outputs(1633) <= not a or b;
    layer0_outputs(1634) <= not b or a;
    layer0_outputs(1635) <= not (a and b);
    layer0_outputs(1636) <= a or b;
    layer0_outputs(1637) <= a xor b;
    layer0_outputs(1638) <= a xor b;
    layer0_outputs(1639) <= not a or b;
    layer0_outputs(1640) <= a;
    layer0_outputs(1641) <= not (a or b);
    layer0_outputs(1642) <= not a or b;
    layer0_outputs(1643) <= not (a xor b);
    layer0_outputs(1644) <= not a or b;
    layer0_outputs(1645) <= not b or a;
    layer0_outputs(1646) <= not a or b;
    layer0_outputs(1647) <= a;
    layer0_outputs(1648) <= b and not a;
    layer0_outputs(1649) <= not (a xor b);
    layer0_outputs(1650) <= not b;
    layer0_outputs(1651) <= not a or b;
    layer0_outputs(1652) <= not a;
    layer0_outputs(1653) <= a and not b;
    layer0_outputs(1654) <= not (a or b);
    layer0_outputs(1655) <= not b;
    layer0_outputs(1656) <= not a or b;
    layer0_outputs(1657) <= a xor b;
    layer0_outputs(1658) <= a xor b;
    layer0_outputs(1659) <= b;
    layer0_outputs(1660) <= b and not a;
    layer0_outputs(1661) <= a xor b;
    layer0_outputs(1662) <= not (a or b);
    layer0_outputs(1663) <= a;
    layer0_outputs(1664) <= not (a or b);
    layer0_outputs(1665) <= not (a or b);
    layer0_outputs(1666) <= a or b;
    layer0_outputs(1667) <= not a or b;
    layer0_outputs(1668) <= a or b;
    layer0_outputs(1669) <= not a or b;
    layer0_outputs(1670) <= a and not b;
    layer0_outputs(1671) <= not (a or b);
    layer0_outputs(1672) <= b;
    layer0_outputs(1673) <= b;
    layer0_outputs(1674) <= not b or a;
    layer0_outputs(1675) <= not a or b;
    layer0_outputs(1676) <= a and b;
    layer0_outputs(1677) <= a xor b;
    layer0_outputs(1678) <= not a;
    layer0_outputs(1679) <= a or b;
    layer0_outputs(1680) <= a or b;
    layer0_outputs(1681) <= '1';
    layer0_outputs(1682) <= not (a or b);
    layer0_outputs(1683) <= a xor b;
    layer0_outputs(1684) <= a or b;
    layer0_outputs(1685) <= b;
    layer0_outputs(1686) <= not (a xor b);
    layer0_outputs(1687) <= b;
    layer0_outputs(1688) <= not b;
    layer0_outputs(1689) <= b and not a;
    layer0_outputs(1690) <= not (a or b);
    layer0_outputs(1691) <= not (a or b);
    layer0_outputs(1692) <= a xor b;
    layer0_outputs(1693) <= b;
    layer0_outputs(1694) <= not (a xor b);
    layer0_outputs(1695) <= not (a xor b);
    layer0_outputs(1696) <= not (a or b);
    layer0_outputs(1697) <= b and not a;
    layer0_outputs(1698) <= a;
    layer0_outputs(1699) <= not (a or b);
    layer0_outputs(1700) <= not (a or b);
    layer0_outputs(1701) <= b;
    layer0_outputs(1702) <= not a;
    layer0_outputs(1703) <= not (a or b);
    layer0_outputs(1704) <= not b;
    layer0_outputs(1705) <= a or b;
    layer0_outputs(1706) <= not (a or b);
    layer0_outputs(1707) <= not a;
    layer0_outputs(1708) <= a xor b;
    layer0_outputs(1709) <= a and not b;
    layer0_outputs(1710) <= not a or b;
    layer0_outputs(1711) <= a and not b;
    layer0_outputs(1712) <= not a or b;
    layer0_outputs(1713) <= not (a or b);
    layer0_outputs(1714) <= not b;
    layer0_outputs(1715) <= not (a or b);
    layer0_outputs(1716) <= a xor b;
    layer0_outputs(1717) <= not (a or b);
    layer0_outputs(1718) <= not a or b;
    layer0_outputs(1719) <= a;
    layer0_outputs(1720) <= b and not a;
    layer0_outputs(1721) <= a and b;
    layer0_outputs(1722) <= a or b;
    layer0_outputs(1723) <= not b or a;
    layer0_outputs(1724) <= a;
    layer0_outputs(1725) <= a;
    layer0_outputs(1726) <= a xor b;
    layer0_outputs(1727) <= a or b;
    layer0_outputs(1728) <= a or b;
    layer0_outputs(1729) <= a xor b;
    layer0_outputs(1730) <= not b;
    layer0_outputs(1731) <= not b;
    layer0_outputs(1732) <= not (a or b);
    layer0_outputs(1733) <= b and not a;
    layer0_outputs(1734) <= a xor b;
    layer0_outputs(1735) <= not b;
    layer0_outputs(1736) <= not a or b;
    layer0_outputs(1737) <= not a or b;
    layer0_outputs(1738) <= a xor b;
    layer0_outputs(1739) <= not b;
    layer0_outputs(1740) <= not (a or b);
    layer0_outputs(1741) <= '0';
    layer0_outputs(1742) <= not (a xor b);
    layer0_outputs(1743) <= b;
    layer0_outputs(1744) <= a or b;
    layer0_outputs(1745) <= a and not b;
    layer0_outputs(1746) <= '0';
    layer0_outputs(1747) <= a and b;
    layer0_outputs(1748) <= a or b;
    layer0_outputs(1749) <= '0';
    layer0_outputs(1750) <= b and not a;
    layer0_outputs(1751) <= a and not b;
    layer0_outputs(1752) <= a xor b;
    layer0_outputs(1753) <= not (a or b);
    layer0_outputs(1754) <= a or b;
    layer0_outputs(1755) <= a xor b;
    layer0_outputs(1756) <= not b;
    layer0_outputs(1757) <= not a or b;
    layer0_outputs(1758) <= not (a or b);
    layer0_outputs(1759) <= b;
    layer0_outputs(1760) <= not a or b;
    layer0_outputs(1761) <= a or b;
    layer0_outputs(1762) <= a;
    layer0_outputs(1763) <= b and not a;
    layer0_outputs(1764) <= not (a and b);
    layer0_outputs(1765) <= not (a or b);
    layer0_outputs(1766) <= not a or b;
    layer0_outputs(1767) <= a or b;
    layer0_outputs(1768) <= a xor b;
    layer0_outputs(1769) <= b and not a;
    layer0_outputs(1770) <= '0';
    layer0_outputs(1771) <= a xor b;
    layer0_outputs(1772) <= a xor b;
    layer0_outputs(1773) <= not (a xor b);
    layer0_outputs(1774) <= not (a or b);
    layer0_outputs(1775) <= a or b;
    layer0_outputs(1776) <= not (a or b);
    layer0_outputs(1777) <= a xor b;
    layer0_outputs(1778) <= b and not a;
    layer0_outputs(1779) <= not (a or b);
    layer0_outputs(1780) <= not a or b;
    layer0_outputs(1781) <= a xor b;
    layer0_outputs(1782) <= not (a xor b);
    layer0_outputs(1783) <= a or b;
    layer0_outputs(1784) <= b and not a;
    layer0_outputs(1785) <= not b or a;
    layer0_outputs(1786) <= not (a xor b);
    layer0_outputs(1787) <= a and not b;
    layer0_outputs(1788) <= not (a and b);
    layer0_outputs(1789) <= not (a xor b);
    layer0_outputs(1790) <= not a or b;
    layer0_outputs(1791) <= b;
    layer0_outputs(1792) <= b and not a;
    layer0_outputs(1793) <= '0';
    layer0_outputs(1794) <= not (a or b);
    layer0_outputs(1795) <= not (a or b);
    layer0_outputs(1796) <= not (a xor b);
    layer0_outputs(1797) <= a or b;
    layer0_outputs(1798) <= not b or a;
    layer0_outputs(1799) <= not a or b;
    layer0_outputs(1800) <= '0';
    layer0_outputs(1801) <= a xor b;
    layer0_outputs(1802) <= not a;
    layer0_outputs(1803) <= not (a or b);
    layer0_outputs(1804) <= not (a xor b);
    layer0_outputs(1805) <= b;
    layer0_outputs(1806) <= not b;
    layer0_outputs(1807) <= not (a or b);
    layer0_outputs(1808) <= not (a xor b);
    layer0_outputs(1809) <= not b;
    layer0_outputs(1810) <= b;
    layer0_outputs(1811) <= not (a or b);
    layer0_outputs(1812) <= a or b;
    layer0_outputs(1813) <= not b;
    layer0_outputs(1814) <= not b or a;
    layer0_outputs(1815) <= not b;
    layer0_outputs(1816) <= not b or a;
    layer0_outputs(1817) <= '0';
    layer0_outputs(1818) <= not (a xor b);
    layer0_outputs(1819) <= b and not a;
    layer0_outputs(1820) <= b and not a;
    layer0_outputs(1821) <= not (a or b);
    layer0_outputs(1822) <= not a;
    layer0_outputs(1823) <= not (a or b);
    layer0_outputs(1824) <= not (a or b);
    layer0_outputs(1825) <= a and not b;
    layer0_outputs(1826) <= not a;
    layer0_outputs(1827) <= a;
    layer0_outputs(1828) <= not (a or b);
    layer0_outputs(1829) <= not (a or b);
    layer0_outputs(1830) <= b;
    layer0_outputs(1831) <= not b;
    layer0_outputs(1832) <= a;
    layer0_outputs(1833) <= not a or b;
    layer0_outputs(1834) <= b;
    layer0_outputs(1835) <= not b or a;
    layer0_outputs(1836) <= not (a or b);
    layer0_outputs(1837) <= not b or a;
    layer0_outputs(1838) <= a and not b;
    layer0_outputs(1839) <= not b or a;
    layer0_outputs(1840) <= a or b;
    layer0_outputs(1841) <= not a or b;
    layer0_outputs(1842) <= a and not b;
    layer0_outputs(1843) <= a xor b;
    layer0_outputs(1844) <= a or b;
    layer0_outputs(1845) <= not (a or b);
    layer0_outputs(1846) <= a or b;
    layer0_outputs(1847) <= a;
    layer0_outputs(1848) <= a or b;
    layer0_outputs(1849) <= b;
    layer0_outputs(1850) <= not (a or b);
    layer0_outputs(1851) <= a and b;
    layer0_outputs(1852) <= a xor b;
    layer0_outputs(1853) <= not (a xor b);
    layer0_outputs(1854) <= not (a or b);
    layer0_outputs(1855) <= b;
    layer0_outputs(1856) <= b and not a;
    layer0_outputs(1857) <= not a;
    layer0_outputs(1858) <= '0';
    layer0_outputs(1859) <= a or b;
    layer0_outputs(1860) <= a xor b;
    layer0_outputs(1861) <= not b;
    layer0_outputs(1862) <= '1';
    layer0_outputs(1863) <= not b;
    layer0_outputs(1864) <= a xor b;
    layer0_outputs(1865) <= a or b;
    layer0_outputs(1866) <= not (a or b);
    layer0_outputs(1867) <= b;
    layer0_outputs(1868) <= not a;
    layer0_outputs(1869) <= not (a or b);
    layer0_outputs(1870) <= a or b;
    layer0_outputs(1871) <= not a or b;
    layer0_outputs(1872) <= a xor b;
    layer0_outputs(1873) <= not b;
    layer0_outputs(1874) <= not (a xor b);
    layer0_outputs(1875) <= '0';
    layer0_outputs(1876) <= b and not a;
    layer0_outputs(1877) <= a or b;
    layer0_outputs(1878) <= a;
    layer0_outputs(1879) <= not (a or b);
    layer0_outputs(1880) <= a;
    layer0_outputs(1881) <= b;
    layer0_outputs(1882) <= b;
    layer0_outputs(1883) <= not a;
    layer0_outputs(1884) <= a or b;
    layer0_outputs(1885) <= a and b;
    layer0_outputs(1886) <= not (a or b);
    layer0_outputs(1887) <= not (a xor b);
    layer0_outputs(1888) <= a xor b;
    layer0_outputs(1889) <= not (a or b);
    layer0_outputs(1890) <= b;
    layer0_outputs(1891) <= b and not a;
    layer0_outputs(1892) <= not b;
    layer0_outputs(1893) <= b;
    layer0_outputs(1894) <= not b or a;
    layer0_outputs(1895) <= a and not b;
    layer0_outputs(1896) <= '0';
    layer0_outputs(1897) <= a or b;
    layer0_outputs(1898) <= a and not b;
    layer0_outputs(1899) <= a xor b;
    layer0_outputs(1900) <= a and not b;
    layer0_outputs(1901) <= a;
    layer0_outputs(1902) <= not (a or b);
    layer0_outputs(1903) <= not (a xor b);
    layer0_outputs(1904) <= a and not b;
    layer0_outputs(1905) <= not a or b;
    layer0_outputs(1906) <= a and not b;
    layer0_outputs(1907) <= a and not b;
    layer0_outputs(1908) <= a or b;
    layer0_outputs(1909) <= not a or b;
    layer0_outputs(1910) <= not b;
    layer0_outputs(1911) <= not (a or b);
    layer0_outputs(1912) <= not (a or b);
    layer0_outputs(1913) <= not b or a;
    layer0_outputs(1914) <= not a or b;
    layer0_outputs(1915) <= not a or b;
    layer0_outputs(1916) <= not (a xor b);
    layer0_outputs(1917) <= a or b;
    layer0_outputs(1918) <= a;
    layer0_outputs(1919) <= b and not a;
    layer0_outputs(1920) <= not a or b;
    layer0_outputs(1921) <= b;
    layer0_outputs(1922) <= b;
    layer0_outputs(1923) <= a;
    layer0_outputs(1924) <= not (a xor b);
    layer0_outputs(1925) <= not (a or b);
    layer0_outputs(1926) <= not b;
    layer0_outputs(1927) <= a xor b;
    layer0_outputs(1928) <= not (a or b);
    layer0_outputs(1929) <= a xor b;
    layer0_outputs(1930) <= not a or b;
    layer0_outputs(1931) <= a or b;
    layer0_outputs(1932) <= a xor b;
    layer0_outputs(1933) <= not b;
    layer0_outputs(1934) <= a and not b;
    layer0_outputs(1935) <= not a or b;
    layer0_outputs(1936) <= '0';
    layer0_outputs(1937) <= not (a or b);
    layer0_outputs(1938) <= not b or a;
    layer0_outputs(1939) <= not b or a;
    layer0_outputs(1940) <= not b;
    layer0_outputs(1941) <= not (a or b);
    layer0_outputs(1942) <= a xor b;
    layer0_outputs(1943) <= not b;
    layer0_outputs(1944) <= not (a or b);
    layer0_outputs(1945) <= a and not b;
    layer0_outputs(1946) <= a;
    layer0_outputs(1947) <= a and not b;
    layer0_outputs(1948) <= a or b;
    layer0_outputs(1949) <= a xor b;
    layer0_outputs(1950) <= not (a xor b);
    layer0_outputs(1951) <= not a;
    layer0_outputs(1952) <= a;
    layer0_outputs(1953) <= a or b;
    layer0_outputs(1954) <= a or b;
    layer0_outputs(1955) <= a or b;
    layer0_outputs(1956) <= a or b;
    layer0_outputs(1957) <= not (a xor b);
    layer0_outputs(1958) <= a xor b;
    layer0_outputs(1959) <= not (a or b);
    layer0_outputs(1960) <= b and not a;
    layer0_outputs(1961) <= not a or b;
    layer0_outputs(1962) <= not (a xor b);
    layer0_outputs(1963) <= not (a or b);
    layer0_outputs(1964) <= a or b;
    layer0_outputs(1965) <= not (a xor b);
    layer0_outputs(1966) <= not (a and b);
    layer0_outputs(1967) <= a and not b;
    layer0_outputs(1968) <= not a or b;
    layer0_outputs(1969) <= b and not a;
    layer0_outputs(1970) <= b;
    layer0_outputs(1971) <= a and b;
    layer0_outputs(1972) <= a or b;
    layer0_outputs(1973) <= not a or b;
    layer0_outputs(1974) <= not (a or b);
    layer0_outputs(1975) <= a or b;
    layer0_outputs(1976) <= not b;
    layer0_outputs(1977) <= not a;
    layer0_outputs(1978) <= not b;
    layer0_outputs(1979) <= not (a or b);
    layer0_outputs(1980) <= a and b;
    layer0_outputs(1981) <= not (a or b);
    layer0_outputs(1982) <= a xor b;
    layer0_outputs(1983) <= not (a or b);
    layer0_outputs(1984) <= not b or a;
    layer0_outputs(1985) <= a xor b;
    layer0_outputs(1986) <= b and not a;
    layer0_outputs(1987) <= not a or b;
    layer0_outputs(1988) <= not (a or b);
    layer0_outputs(1989) <= a;
    layer0_outputs(1990) <= b and not a;
    layer0_outputs(1991) <= a or b;
    layer0_outputs(1992) <= not a;
    layer0_outputs(1993) <= a;
    layer0_outputs(1994) <= not (a and b);
    layer0_outputs(1995) <= a or b;
    layer0_outputs(1996) <= not a or b;
    layer0_outputs(1997) <= not (a or b);
    layer0_outputs(1998) <= not b or a;
    layer0_outputs(1999) <= a or b;
    layer0_outputs(2000) <= a or b;
    layer0_outputs(2001) <= not a or b;
    layer0_outputs(2002) <= not (a or b);
    layer0_outputs(2003) <= not (a or b);
    layer0_outputs(2004) <= b and not a;
    layer0_outputs(2005) <= a;
    layer0_outputs(2006) <= not a or b;
    layer0_outputs(2007) <= a or b;
    layer0_outputs(2008) <= b and not a;
    layer0_outputs(2009) <= not b;
    layer0_outputs(2010) <= not a or b;
    layer0_outputs(2011) <= b and not a;
    layer0_outputs(2012) <= not b or a;
    layer0_outputs(2013) <= a;
    layer0_outputs(2014) <= a or b;
    layer0_outputs(2015) <= not a;
    layer0_outputs(2016) <= a or b;
    layer0_outputs(2017) <= not (a or b);
    layer0_outputs(2018) <= b and not a;
    layer0_outputs(2019) <= not b or a;
    layer0_outputs(2020) <= a or b;
    layer0_outputs(2021) <= b and not a;
    layer0_outputs(2022) <= a xor b;
    layer0_outputs(2023) <= b and not a;
    layer0_outputs(2024) <= b;
    layer0_outputs(2025) <= a or b;
    layer0_outputs(2026) <= a and b;
    layer0_outputs(2027) <= a xor b;
    layer0_outputs(2028) <= a;
    layer0_outputs(2029) <= not b;
    layer0_outputs(2030) <= not b;
    layer0_outputs(2031) <= a or b;
    layer0_outputs(2032) <= not (a or b);
    layer0_outputs(2033) <= not a or b;
    layer0_outputs(2034) <= not (a xor b);
    layer0_outputs(2035) <= a or b;
    layer0_outputs(2036) <= not b or a;
    layer0_outputs(2037) <= not b;
    layer0_outputs(2038) <= not b;
    layer0_outputs(2039) <= not a;
    layer0_outputs(2040) <= a;
    layer0_outputs(2041) <= a or b;
    layer0_outputs(2042) <= not (a or b);
    layer0_outputs(2043) <= a or b;
    layer0_outputs(2044) <= a;
    layer0_outputs(2045) <= not (a xor b);
    layer0_outputs(2046) <= a;
    layer0_outputs(2047) <= not (a or b);
    layer0_outputs(2048) <= b and not a;
    layer0_outputs(2049) <= b and not a;
    layer0_outputs(2050) <= not a or b;
    layer0_outputs(2051) <= not a or b;
    layer0_outputs(2052) <= a or b;
    layer0_outputs(2053) <= '0';
    layer0_outputs(2054) <= not a;
    layer0_outputs(2055) <= not (a or b);
    layer0_outputs(2056) <= not a;
    layer0_outputs(2057) <= not b or a;
    layer0_outputs(2058) <= a;
    layer0_outputs(2059) <= not a;
    layer0_outputs(2060) <= b and not a;
    layer0_outputs(2061) <= a xor b;
    layer0_outputs(2062) <= a and b;
    layer0_outputs(2063) <= '0';
    layer0_outputs(2064) <= a or b;
    layer0_outputs(2065) <= not (a or b);
    layer0_outputs(2066) <= not b or a;
    layer0_outputs(2067) <= a;
    layer0_outputs(2068) <= a xor b;
    layer0_outputs(2069) <= not b or a;
    layer0_outputs(2070) <= a and b;
    layer0_outputs(2071) <= not (a and b);
    layer0_outputs(2072) <= not (a or b);
    layer0_outputs(2073) <= not (a or b);
    layer0_outputs(2074) <= b;
    layer0_outputs(2075) <= b and not a;
    layer0_outputs(2076) <= a and not b;
    layer0_outputs(2077) <= a xor b;
    layer0_outputs(2078) <= a or b;
    layer0_outputs(2079) <= not (a xor b);
    layer0_outputs(2080) <= a;
    layer0_outputs(2081) <= not a;
    layer0_outputs(2082) <= not b;
    layer0_outputs(2083) <= a or b;
    layer0_outputs(2084) <= not a or b;
    layer0_outputs(2085) <= a or b;
    layer0_outputs(2086) <= b and not a;
    layer0_outputs(2087) <= a or b;
    layer0_outputs(2088) <= a or b;
    layer0_outputs(2089) <= a;
    layer0_outputs(2090) <= not (a or b);
    layer0_outputs(2091) <= a or b;
    layer0_outputs(2092) <= '0';
    layer0_outputs(2093) <= not (a or b);
    layer0_outputs(2094) <= a;
    layer0_outputs(2095) <= '0';
    layer0_outputs(2096) <= a xor b;
    layer0_outputs(2097) <= not a;
    layer0_outputs(2098) <= '1';
    layer0_outputs(2099) <= not a or b;
    layer0_outputs(2100) <= not b;
    layer0_outputs(2101) <= not (a or b);
    layer0_outputs(2102) <= not (a or b);
    layer0_outputs(2103) <= '1';
    layer0_outputs(2104) <= not b or a;
    layer0_outputs(2105) <= not (a or b);
    layer0_outputs(2106) <= b;
    layer0_outputs(2107) <= '1';
    layer0_outputs(2108) <= a xor b;
    layer0_outputs(2109) <= not b;
    layer0_outputs(2110) <= not (a or b);
    layer0_outputs(2111) <= not (a or b);
    layer0_outputs(2112) <= not b;
    layer0_outputs(2113) <= a and not b;
    layer0_outputs(2114) <= a or b;
    layer0_outputs(2115) <= not a or b;
    layer0_outputs(2116) <= a and not b;
    layer0_outputs(2117) <= a or b;
    layer0_outputs(2118) <= not (a or b);
    layer0_outputs(2119) <= not (a or b);
    layer0_outputs(2120) <= not (a or b);
    layer0_outputs(2121) <= b and not a;
    layer0_outputs(2122) <= not b or a;
    layer0_outputs(2123) <= b;
    layer0_outputs(2124) <= not b;
    layer0_outputs(2125) <= not b;
    layer0_outputs(2126) <= not b or a;
    layer0_outputs(2127) <= not (a and b);
    layer0_outputs(2128) <= not b or a;
    layer0_outputs(2129) <= a or b;
    layer0_outputs(2130) <= a and not b;
    layer0_outputs(2131) <= not a or b;
    layer0_outputs(2132) <= not a or b;
    layer0_outputs(2133) <= b;
    layer0_outputs(2134) <= a;
    layer0_outputs(2135) <= not a;
    layer0_outputs(2136) <= not a;
    layer0_outputs(2137) <= a xor b;
    layer0_outputs(2138) <= a or b;
    layer0_outputs(2139) <= not b;
    layer0_outputs(2140) <= not b;
    layer0_outputs(2141) <= not (a or b);
    layer0_outputs(2142) <= a and not b;
    layer0_outputs(2143) <= not b or a;
    layer0_outputs(2144) <= not a;
    layer0_outputs(2145) <= a or b;
    layer0_outputs(2146) <= not a or b;
    layer0_outputs(2147) <= not (a xor b);
    layer0_outputs(2148) <= a or b;
    layer0_outputs(2149) <= not b or a;
    layer0_outputs(2150) <= not a;
    layer0_outputs(2151) <= a and not b;
    layer0_outputs(2152) <= a or b;
    layer0_outputs(2153) <= a xor b;
    layer0_outputs(2154) <= a and not b;
    layer0_outputs(2155) <= not b;
    layer0_outputs(2156) <= '0';
    layer0_outputs(2157) <= not (a or b);
    layer0_outputs(2158) <= not (a or b);
    layer0_outputs(2159) <= a or b;
    layer0_outputs(2160) <= a xor b;
    layer0_outputs(2161) <= b;
    layer0_outputs(2162) <= a or b;
    layer0_outputs(2163) <= '1';
    layer0_outputs(2164) <= not b;
    layer0_outputs(2165) <= not (a or b);
    layer0_outputs(2166) <= a and not b;
    layer0_outputs(2167) <= a;
    layer0_outputs(2168) <= '0';
    layer0_outputs(2169) <= b;
    layer0_outputs(2170) <= a xor b;
    layer0_outputs(2171) <= b and not a;
    layer0_outputs(2172) <= not (a xor b);
    layer0_outputs(2173) <= not b;
    layer0_outputs(2174) <= a and b;
    layer0_outputs(2175) <= a xor b;
    layer0_outputs(2176) <= not b;
    layer0_outputs(2177) <= not (a xor b);
    layer0_outputs(2178) <= not a;
    layer0_outputs(2179) <= not b or a;
    layer0_outputs(2180) <= a or b;
    layer0_outputs(2181) <= a and not b;
    layer0_outputs(2182) <= b;
    layer0_outputs(2183) <= not (a or b);
    layer0_outputs(2184) <= not b;
    layer0_outputs(2185) <= a xor b;
    layer0_outputs(2186) <= a xor b;
    layer0_outputs(2187) <= not (a or b);
    layer0_outputs(2188) <= not (a and b);
    layer0_outputs(2189) <= a xor b;
    layer0_outputs(2190) <= a;
    layer0_outputs(2191) <= a or b;
    layer0_outputs(2192) <= not (a or b);
    layer0_outputs(2193) <= not b or a;
    layer0_outputs(2194) <= a or b;
    layer0_outputs(2195) <= '0';
    layer0_outputs(2196) <= a and not b;
    layer0_outputs(2197) <= '1';
    layer0_outputs(2198) <= not b;
    layer0_outputs(2199) <= not a or b;
    layer0_outputs(2200) <= a or b;
    layer0_outputs(2201) <= not a or b;
    layer0_outputs(2202) <= not (a or b);
    layer0_outputs(2203) <= a or b;
    layer0_outputs(2204) <= not b or a;
    layer0_outputs(2205) <= not b or a;
    layer0_outputs(2206) <= not a;
    layer0_outputs(2207) <= a and not b;
    layer0_outputs(2208) <= a;
    layer0_outputs(2209) <= not (a xor b);
    layer0_outputs(2210) <= not b;
    layer0_outputs(2211) <= a and not b;
    layer0_outputs(2212) <= not (a or b);
    layer0_outputs(2213) <= a xor b;
    layer0_outputs(2214) <= not (a or b);
    layer0_outputs(2215) <= '1';
    layer0_outputs(2216) <= not b;
    layer0_outputs(2217) <= not (a xor b);
    layer0_outputs(2218) <= b;
    layer0_outputs(2219) <= a;
    layer0_outputs(2220) <= not (a or b);
    layer0_outputs(2221) <= not a or b;
    layer0_outputs(2222) <= not (a and b);
    layer0_outputs(2223) <= not b;
    layer0_outputs(2224) <= '1';
    layer0_outputs(2225) <= not (a xor b);
    layer0_outputs(2226) <= a xor b;
    layer0_outputs(2227) <= b;
    layer0_outputs(2228) <= not a;
    layer0_outputs(2229) <= b and not a;
    layer0_outputs(2230) <= not a;
    layer0_outputs(2231) <= not (a and b);
    layer0_outputs(2232) <= not a;
    layer0_outputs(2233) <= not a or b;
    layer0_outputs(2234) <= b;
    layer0_outputs(2235) <= not (a or b);
    layer0_outputs(2236) <= not (a or b);
    layer0_outputs(2237) <= not b;
    layer0_outputs(2238) <= a or b;
    layer0_outputs(2239) <= a and not b;
    layer0_outputs(2240) <= a or b;
    layer0_outputs(2241) <= b;
    layer0_outputs(2242) <= not (a or b);
    layer0_outputs(2243) <= not (a or b);
    layer0_outputs(2244) <= a and not b;
    layer0_outputs(2245) <= b;
    layer0_outputs(2246) <= not (a xor b);
    layer0_outputs(2247) <= a and b;
    layer0_outputs(2248) <= b;
    layer0_outputs(2249) <= not (a or b);
    layer0_outputs(2250) <= a or b;
    layer0_outputs(2251) <= '1';
    layer0_outputs(2252) <= a or b;
    layer0_outputs(2253) <= not b;
    layer0_outputs(2254) <= not a or b;
    layer0_outputs(2255) <= a xor b;
    layer0_outputs(2256) <= a and not b;
    layer0_outputs(2257) <= b and not a;
    layer0_outputs(2258) <= not a or b;
    layer0_outputs(2259) <= '1';
    layer0_outputs(2260) <= a or b;
    layer0_outputs(2261) <= not a;
    layer0_outputs(2262) <= not (a or b);
    layer0_outputs(2263) <= not (a or b);
    layer0_outputs(2264) <= b;
    layer0_outputs(2265) <= not (a or b);
    layer0_outputs(2266) <= not (a or b);
    layer0_outputs(2267) <= not a or b;
    layer0_outputs(2268) <= not (a or b);
    layer0_outputs(2269) <= a or b;
    layer0_outputs(2270) <= not b;
    layer0_outputs(2271) <= a;
    layer0_outputs(2272) <= '0';
    layer0_outputs(2273) <= a or b;
    layer0_outputs(2274) <= a or b;
    layer0_outputs(2275) <= a and b;
    layer0_outputs(2276) <= a;
    layer0_outputs(2277) <= not a;
    layer0_outputs(2278) <= b and not a;
    layer0_outputs(2279) <= a xor b;
    layer0_outputs(2280) <= '1';
    layer0_outputs(2281) <= b and not a;
    layer0_outputs(2282) <= not a;
    layer0_outputs(2283) <= not (a or b);
    layer0_outputs(2284) <= not b;
    layer0_outputs(2285) <= a and not b;
    layer0_outputs(2286) <= not (a xor b);
    layer0_outputs(2287) <= a or b;
    layer0_outputs(2288) <= not (a xor b);
    layer0_outputs(2289) <= a and not b;
    layer0_outputs(2290) <= not (a xor b);
    layer0_outputs(2291) <= b and not a;
    layer0_outputs(2292) <= not a;
    layer0_outputs(2293) <= not (a or b);
    layer0_outputs(2294) <= a or b;
    layer0_outputs(2295) <= not b;
    layer0_outputs(2296) <= a and not b;
    layer0_outputs(2297) <= a or b;
    layer0_outputs(2298) <= not a;
    layer0_outputs(2299) <= not (a and b);
    layer0_outputs(2300) <= a and b;
    layer0_outputs(2301) <= a xor b;
    layer0_outputs(2302) <= not (a xor b);
    layer0_outputs(2303) <= not (a and b);
    layer0_outputs(2304) <= not b;
    layer0_outputs(2305) <= b;
    layer0_outputs(2306) <= not (a or b);
    layer0_outputs(2307) <= a or b;
    layer0_outputs(2308) <= b;
    layer0_outputs(2309) <= not a;
    layer0_outputs(2310) <= not (a and b);
    layer0_outputs(2311) <= not b or a;
    layer0_outputs(2312) <= a or b;
    layer0_outputs(2313) <= not (a or b);
    layer0_outputs(2314) <= not a or b;
    layer0_outputs(2315) <= a or b;
    layer0_outputs(2316) <= a xor b;
    layer0_outputs(2317) <= not (a or b);
    layer0_outputs(2318) <= '0';
    layer0_outputs(2319) <= a xor b;
    layer0_outputs(2320) <= a or b;
    layer0_outputs(2321) <= a or b;
    layer0_outputs(2322) <= a;
    layer0_outputs(2323) <= a or b;
    layer0_outputs(2324) <= a and not b;
    layer0_outputs(2325) <= b and not a;
    layer0_outputs(2326) <= not (a xor b);
    layer0_outputs(2327) <= a xor b;
    layer0_outputs(2328) <= b;
    layer0_outputs(2329) <= a or b;
    layer0_outputs(2330) <= a or b;
    layer0_outputs(2331) <= b and not a;
    layer0_outputs(2332) <= not (a or b);
    layer0_outputs(2333) <= not b;
    layer0_outputs(2334) <= a or b;
    layer0_outputs(2335) <= b and not a;
    layer0_outputs(2336) <= a xor b;
    layer0_outputs(2337) <= a xor b;
    layer0_outputs(2338) <= a;
    layer0_outputs(2339) <= not b;
    layer0_outputs(2340) <= not b or a;
    layer0_outputs(2341) <= a xor b;
    layer0_outputs(2342) <= not (a xor b);
    layer0_outputs(2343) <= not (a or b);
    layer0_outputs(2344) <= not a or b;
    layer0_outputs(2345) <= a and not b;
    layer0_outputs(2346) <= a or b;
    layer0_outputs(2347) <= not (a xor b);
    layer0_outputs(2348) <= '1';
    layer0_outputs(2349) <= a xor b;
    layer0_outputs(2350) <= not (a or b);
    layer0_outputs(2351) <= a;
    layer0_outputs(2352) <= not a;
    layer0_outputs(2353) <= a xor b;
    layer0_outputs(2354) <= a or b;
    layer0_outputs(2355) <= not a;
    layer0_outputs(2356) <= a or b;
    layer0_outputs(2357) <= not b;
    layer0_outputs(2358) <= b;
    layer0_outputs(2359) <= a xor b;
    layer0_outputs(2360) <= a xor b;
    layer0_outputs(2361) <= a;
    layer0_outputs(2362) <= not (a or b);
    layer0_outputs(2363) <= not (a xor b);
    layer0_outputs(2364) <= '1';
    layer0_outputs(2365) <= not (a or b);
    layer0_outputs(2366) <= b and not a;
    layer0_outputs(2367) <= '1';
    layer0_outputs(2368) <= a;
    layer0_outputs(2369) <= a and not b;
    layer0_outputs(2370) <= a;
    layer0_outputs(2371) <= not a or b;
    layer0_outputs(2372) <= a or b;
    layer0_outputs(2373) <= not (a or b);
    layer0_outputs(2374) <= a or b;
    layer0_outputs(2375) <= not a or b;
    layer0_outputs(2376) <= '1';
    layer0_outputs(2377) <= b and not a;
    layer0_outputs(2378) <= not (a and b);
    layer0_outputs(2379) <= not b;
    layer0_outputs(2380) <= a or b;
    layer0_outputs(2381) <= a or b;
    layer0_outputs(2382) <= a and b;
    layer0_outputs(2383) <= a and b;
    layer0_outputs(2384) <= not a;
    layer0_outputs(2385) <= a xor b;
    layer0_outputs(2386) <= b;
    layer0_outputs(2387) <= a or b;
    layer0_outputs(2388) <= a and b;
    layer0_outputs(2389) <= not a or b;
    layer0_outputs(2390) <= not (a or b);
    layer0_outputs(2391) <= not b or a;
    layer0_outputs(2392) <= a;
    layer0_outputs(2393) <= not a;
    layer0_outputs(2394) <= a xor b;
    layer0_outputs(2395) <= not (a or b);
    layer0_outputs(2396) <= '1';
    layer0_outputs(2397) <= '1';
    layer0_outputs(2398) <= a xor b;
    layer0_outputs(2399) <= a;
    layer0_outputs(2400) <= not b or a;
    layer0_outputs(2401) <= not b;
    layer0_outputs(2402) <= not (a or b);
    layer0_outputs(2403) <= not (a xor b);
    layer0_outputs(2404) <= not b;
    layer0_outputs(2405) <= a;
    layer0_outputs(2406) <= not a;
    layer0_outputs(2407) <= not a;
    layer0_outputs(2408) <= not (a and b);
    layer0_outputs(2409) <= b;
    layer0_outputs(2410) <= not (a xor b);
    layer0_outputs(2411) <= a;
    layer0_outputs(2412) <= b;
    layer0_outputs(2413) <= a or b;
    layer0_outputs(2414) <= not a;
    layer0_outputs(2415) <= a and not b;
    layer0_outputs(2416) <= not (a or b);
    layer0_outputs(2417) <= a xor b;
    layer0_outputs(2418) <= not (a xor b);
    layer0_outputs(2419) <= a and not b;
    layer0_outputs(2420) <= a or b;
    layer0_outputs(2421) <= a and b;
    layer0_outputs(2422) <= a or b;
    layer0_outputs(2423) <= a and not b;
    layer0_outputs(2424) <= not (a xor b);
    layer0_outputs(2425) <= not a;
    layer0_outputs(2426) <= a xor b;
    layer0_outputs(2427) <= a or b;
    layer0_outputs(2428) <= not b;
    layer0_outputs(2429) <= a and b;
    layer0_outputs(2430) <= not b;
    layer0_outputs(2431) <= a and b;
    layer0_outputs(2432) <= a or b;
    layer0_outputs(2433) <= not (a or b);
    layer0_outputs(2434) <= a or b;
    layer0_outputs(2435) <= a or b;
    layer0_outputs(2436) <= not (a or b);
    layer0_outputs(2437) <= a;
    layer0_outputs(2438) <= not (a xor b);
    layer0_outputs(2439) <= a and b;
    layer0_outputs(2440) <= not b or a;
    layer0_outputs(2441) <= not (a xor b);
    layer0_outputs(2442) <= not b or a;
    layer0_outputs(2443) <= not (a xor b);
    layer0_outputs(2444) <= not (a or b);
    layer0_outputs(2445) <= not b;
    layer0_outputs(2446) <= not (a and b);
    layer0_outputs(2447) <= not (a xor b);
    layer0_outputs(2448) <= b and not a;
    layer0_outputs(2449) <= not (a xor b);
    layer0_outputs(2450) <= not a or b;
    layer0_outputs(2451) <= a and not b;
    layer0_outputs(2452) <= not (a or b);
    layer0_outputs(2453) <= '1';
    layer0_outputs(2454) <= '1';
    layer0_outputs(2455) <= not (a xor b);
    layer0_outputs(2456) <= not b or a;
    layer0_outputs(2457) <= a xor b;
    layer0_outputs(2458) <= '0';
    layer0_outputs(2459) <= not (a and b);
    layer0_outputs(2460) <= a xor b;
    layer0_outputs(2461) <= a xor b;
    layer0_outputs(2462) <= not b;
    layer0_outputs(2463) <= not (a or b);
    layer0_outputs(2464) <= b;
    layer0_outputs(2465) <= not (a or b);
    layer0_outputs(2466) <= not a or b;
    layer0_outputs(2467) <= a or b;
    layer0_outputs(2468) <= a;
    layer0_outputs(2469) <= b;
    layer0_outputs(2470) <= '0';
    layer0_outputs(2471) <= not (a or b);
    layer0_outputs(2472) <= a;
    layer0_outputs(2473) <= a or b;
    layer0_outputs(2474) <= b;
    layer0_outputs(2475) <= a or b;
    layer0_outputs(2476) <= '0';
    layer0_outputs(2477) <= not (a xor b);
    layer0_outputs(2478) <= '1';
    layer0_outputs(2479) <= not b;
    layer0_outputs(2480) <= b;
    layer0_outputs(2481) <= a or b;
    layer0_outputs(2482) <= a xor b;
    layer0_outputs(2483) <= not (a xor b);
    layer0_outputs(2484) <= not (a or b);
    layer0_outputs(2485) <= b;
    layer0_outputs(2486) <= a;
    layer0_outputs(2487) <= not a;
    layer0_outputs(2488) <= not (a or b);
    layer0_outputs(2489) <= not a or b;
    layer0_outputs(2490) <= not a or b;
    layer0_outputs(2491) <= a xor b;
    layer0_outputs(2492) <= b and not a;
    layer0_outputs(2493) <= not (a or b);
    layer0_outputs(2494) <= a;
    layer0_outputs(2495) <= a xor b;
    layer0_outputs(2496) <= b and not a;
    layer0_outputs(2497) <= not (a or b);
    layer0_outputs(2498) <= not (a and b);
    layer0_outputs(2499) <= not (a or b);
    layer0_outputs(2500) <= not (a or b);
    layer0_outputs(2501) <= not b;
    layer0_outputs(2502) <= a and not b;
    layer0_outputs(2503) <= not a or b;
    layer0_outputs(2504) <= not a or b;
    layer0_outputs(2505) <= a and not b;
    layer0_outputs(2506) <= not a;
    layer0_outputs(2507) <= not (a or b);
    layer0_outputs(2508) <= a;
    layer0_outputs(2509) <= not (a or b);
    layer0_outputs(2510) <= b and not a;
    layer0_outputs(2511) <= not (a or b);
    layer0_outputs(2512) <= '1';
    layer0_outputs(2513) <= not (a or b);
    layer0_outputs(2514) <= b;
    layer0_outputs(2515) <= a or b;
    layer0_outputs(2516) <= b and not a;
    layer0_outputs(2517) <= a or b;
    layer0_outputs(2518) <= not (a or b);
    layer0_outputs(2519) <= not b;
    layer0_outputs(2520) <= a or b;
    layer0_outputs(2521) <= b;
    layer0_outputs(2522) <= not (a or b);
    layer0_outputs(2523) <= b and not a;
    layer0_outputs(2524) <= not a;
    layer0_outputs(2525) <= not (a or b);
    layer0_outputs(2526) <= not a or b;
    layer0_outputs(2527) <= a or b;
    layer0_outputs(2528) <= not (a or b);
    layer0_outputs(2529) <= a and not b;
    layer0_outputs(2530) <= not (a xor b);
    layer0_outputs(2531) <= not a or b;
    layer0_outputs(2532) <= not (a or b);
    layer0_outputs(2533) <= a or b;
    layer0_outputs(2534) <= not (a or b);
    layer0_outputs(2535) <= not b or a;
    layer0_outputs(2536) <= a xor b;
    layer0_outputs(2537) <= not (a or b);
    layer0_outputs(2538) <= a xor b;
    layer0_outputs(2539) <= a xor b;
    layer0_outputs(2540) <= not a;
    layer0_outputs(2541) <= not b or a;
    layer0_outputs(2542) <= not (a or b);
    layer0_outputs(2543) <= a or b;
    layer0_outputs(2544) <= not (a or b);
    layer0_outputs(2545) <= a and not b;
    layer0_outputs(2546) <= a xor b;
    layer0_outputs(2547) <= a and not b;
    layer0_outputs(2548) <= not (a xor b);
    layer0_outputs(2549) <= not (a or b);
    layer0_outputs(2550) <= not (a or b);
    layer0_outputs(2551) <= a or b;
    layer0_outputs(2552) <= b;
    layer0_outputs(2553) <= a or b;
    layer0_outputs(2554) <= a or b;
    layer0_outputs(2555) <= a or b;
    layer0_outputs(2556) <= not b;
    layer0_outputs(2557) <= not (a and b);
    layer0_outputs(2558) <= a and not b;
    layer0_outputs(2559) <= a or b;
    layer0_outputs(2560) <= a xor b;
    layer0_outputs(2561) <= not (a and b);
    layer0_outputs(2562) <= a and not b;
    layer0_outputs(2563) <= a or b;
    layer0_outputs(2564) <= not a;
    layer0_outputs(2565) <= not (a xor b);
    layer0_outputs(2566) <= not b;
    layer0_outputs(2567) <= a and not b;
    layer0_outputs(2568) <= not a;
    layer0_outputs(2569) <= a or b;
    layer0_outputs(2570) <= b and not a;
    layer0_outputs(2571) <= a xor b;
    layer0_outputs(2572) <= a or b;
    layer0_outputs(2573) <= not b or a;
    layer0_outputs(2574) <= not b or a;
    layer0_outputs(2575) <= a or b;
    layer0_outputs(2576) <= a or b;
    layer0_outputs(2577) <= not (a xor b);
    layer0_outputs(2578) <= not (a xor b);
    layer0_outputs(2579) <= a;
    layer0_outputs(2580) <= a or b;
    layer0_outputs(2581) <= b;
    layer0_outputs(2582) <= not a or b;
    layer0_outputs(2583) <= not b;
    layer0_outputs(2584) <= not b;
    layer0_outputs(2585) <= a;
    layer0_outputs(2586) <= a and not b;
    layer0_outputs(2587) <= not (a xor b);
    layer0_outputs(2588) <= b and not a;
    layer0_outputs(2589) <= '1';
    layer0_outputs(2590) <= not b;
    layer0_outputs(2591) <= not (a or b);
    layer0_outputs(2592) <= a or b;
    layer0_outputs(2593) <= a or b;
    layer0_outputs(2594) <= a xor b;
    layer0_outputs(2595) <= b;
    layer0_outputs(2596) <= not b;
    layer0_outputs(2597) <= not a or b;
    layer0_outputs(2598) <= b and not a;
    layer0_outputs(2599) <= b;
    layer0_outputs(2600) <= not (a or b);
    layer0_outputs(2601) <= a or b;
    layer0_outputs(2602) <= not a or b;
    layer0_outputs(2603) <= not (a xor b);
    layer0_outputs(2604) <= not b or a;
    layer0_outputs(2605) <= not (a or b);
    layer0_outputs(2606) <= not (a or b);
    layer0_outputs(2607) <= a and not b;
    layer0_outputs(2608) <= not a or b;
    layer0_outputs(2609) <= not (a or b);
    layer0_outputs(2610) <= not a or b;
    layer0_outputs(2611) <= b;
    layer0_outputs(2612) <= a xor b;
    layer0_outputs(2613) <= a;
    layer0_outputs(2614) <= not (a or b);
    layer0_outputs(2615) <= not b;
    layer0_outputs(2616) <= not a or b;
    layer0_outputs(2617) <= a or b;
    layer0_outputs(2618) <= not (a or b);
    layer0_outputs(2619) <= not b;
    layer0_outputs(2620) <= a and not b;
    layer0_outputs(2621) <= not (a or b);
    layer0_outputs(2622) <= not (a or b);
    layer0_outputs(2623) <= a xor b;
    layer0_outputs(2624) <= not a;
    layer0_outputs(2625) <= not b;
    layer0_outputs(2626) <= not (a xor b);
    layer0_outputs(2627) <= not b or a;
    layer0_outputs(2628) <= b;
    layer0_outputs(2629) <= not (a xor b);
    layer0_outputs(2630) <= not b or a;
    layer0_outputs(2631) <= not a;
    layer0_outputs(2632) <= not a or b;
    layer0_outputs(2633) <= b;
    layer0_outputs(2634) <= not (a or b);
    layer0_outputs(2635) <= '0';
    layer0_outputs(2636) <= not a or b;
    layer0_outputs(2637) <= not b or a;
    layer0_outputs(2638) <= not a;
    layer0_outputs(2639) <= '0';
    layer0_outputs(2640) <= a or b;
    layer0_outputs(2641) <= a or b;
    layer0_outputs(2642) <= not (a and b);
    layer0_outputs(2643) <= not (a or b);
    layer0_outputs(2644) <= not (a or b);
    layer0_outputs(2645) <= not a or b;
    layer0_outputs(2646) <= a or b;
    layer0_outputs(2647) <= not (a or b);
    layer0_outputs(2648) <= a and b;
    layer0_outputs(2649) <= not (a xor b);
    layer0_outputs(2650) <= b and not a;
    layer0_outputs(2651) <= not (a xor b);
    layer0_outputs(2652) <= not b or a;
    layer0_outputs(2653) <= a and not b;
    layer0_outputs(2654) <= not (a or b);
    layer0_outputs(2655) <= not (a xor b);
    layer0_outputs(2656) <= b;
    layer0_outputs(2657) <= a or b;
    layer0_outputs(2658) <= a;
    layer0_outputs(2659) <= b;
    layer0_outputs(2660) <= a and not b;
    layer0_outputs(2661) <= not (a or b);
    layer0_outputs(2662) <= not a or b;
    layer0_outputs(2663) <= not (a xor b);
    layer0_outputs(2664) <= not a;
    layer0_outputs(2665) <= a;
    layer0_outputs(2666) <= not (a or b);
    layer0_outputs(2667) <= not (a or b);
    layer0_outputs(2668) <= a and not b;
    layer0_outputs(2669) <= a;
    layer0_outputs(2670) <= not a;
    layer0_outputs(2671) <= a or b;
    layer0_outputs(2672) <= a xor b;
    layer0_outputs(2673) <= a;
    layer0_outputs(2674) <= a;
    layer0_outputs(2675) <= a or b;
    layer0_outputs(2676) <= a;
    layer0_outputs(2677) <= not (a or b);
    layer0_outputs(2678) <= b;
    layer0_outputs(2679) <= a;
    layer0_outputs(2680) <= a or b;
    layer0_outputs(2681) <= not a or b;
    layer0_outputs(2682) <= not (a or b);
    layer0_outputs(2683) <= a and b;
    layer0_outputs(2684) <= a xor b;
    layer0_outputs(2685) <= a or b;
    layer0_outputs(2686) <= a xor b;
    layer0_outputs(2687) <= not b;
    layer0_outputs(2688) <= a or b;
    layer0_outputs(2689) <= not (a or b);
    layer0_outputs(2690) <= a or b;
    layer0_outputs(2691) <= not b;
    layer0_outputs(2692) <= not b;
    layer0_outputs(2693) <= not (a or b);
    layer0_outputs(2694) <= not (a xor b);
    layer0_outputs(2695) <= a xor b;
    layer0_outputs(2696) <= not b;
    layer0_outputs(2697) <= b;
    layer0_outputs(2698) <= not (a or b);
    layer0_outputs(2699) <= '1';
    layer0_outputs(2700) <= not (a or b);
    layer0_outputs(2701) <= b;
    layer0_outputs(2702) <= a xor b;
    layer0_outputs(2703) <= not a;
    layer0_outputs(2704) <= a or b;
    layer0_outputs(2705) <= b;
    layer0_outputs(2706) <= not (a or b);
    layer0_outputs(2707) <= a or b;
    layer0_outputs(2708) <= b;
    layer0_outputs(2709) <= not b;
    layer0_outputs(2710) <= not b or a;
    layer0_outputs(2711) <= not a or b;
    layer0_outputs(2712) <= a or b;
    layer0_outputs(2713) <= a;
    layer0_outputs(2714) <= '1';
    layer0_outputs(2715) <= not b or a;
    layer0_outputs(2716) <= a xor b;
    layer0_outputs(2717) <= a or b;
    layer0_outputs(2718) <= not (a or b);
    layer0_outputs(2719) <= a or b;
    layer0_outputs(2720) <= a and not b;
    layer0_outputs(2721) <= not a or b;
    layer0_outputs(2722) <= a or b;
    layer0_outputs(2723) <= b and not a;
    layer0_outputs(2724) <= a xor b;
    layer0_outputs(2725) <= b and not a;
    layer0_outputs(2726) <= b and not a;
    layer0_outputs(2727) <= a;
    layer0_outputs(2728) <= b;
    layer0_outputs(2729) <= b;
    layer0_outputs(2730) <= not a or b;
    layer0_outputs(2731) <= not (a or b);
    layer0_outputs(2732) <= b and not a;
    layer0_outputs(2733) <= not (a or b);
    layer0_outputs(2734) <= b and not a;
    layer0_outputs(2735) <= not a or b;
    layer0_outputs(2736) <= a and not b;
    layer0_outputs(2737) <= not b;
    layer0_outputs(2738) <= a;
    layer0_outputs(2739) <= a or b;
    layer0_outputs(2740) <= a;
    layer0_outputs(2741) <= a or b;
    layer0_outputs(2742) <= not (a or b);
    layer0_outputs(2743) <= '1';
    layer0_outputs(2744) <= a;
    layer0_outputs(2745) <= a or b;
    layer0_outputs(2746) <= a or b;
    layer0_outputs(2747) <= a xor b;
    layer0_outputs(2748) <= a xor b;
    layer0_outputs(2749) <= not b or a;
    layer0_outputs(2750) <= a and not b;
    layer0_outputs(2751) <= not b or a;
    layer0_outputs(2752) <= not (a xor b);
    layer0_outputs(2753) <= b;
    layer0_outputs(2754) <= not a or b;
    layer0_outputs(2755) <= a xor b;
    layer0_outputs(2756) <= not a;
    layer0_outputs(2757) <= a;
    layer0_outputs(2758) <= b and not a;
    layer0_outputs(2759) <= not b or a;
    layer0_outputs(2760) <= '1';
    layer0_outputs(2761) <= a;
    layer0_outputs(2762) <= '1';
    layer0_outputs(2763) <= not a or b;
    layer0_outputs(2764) <= not b;
    layer0_outputs(2765) <= not a or b;
    layer0_outputs(2766) <= a and not b;
    layer0_outputs(2767) <= not a;
    layer0_outputs(2768) <= not a or b;
    layer0_outputs(2769) <= not b or a;
    layer0_outputs(2770) <= b;
    layer0_outputs(2771) <= a or b;
    layer0_outputs(2772) <= a and not b;
    layer0_outputs(2773) <= a or b;
    layer0_outputs(2774) <= not (a xor b);
    layer0_outputs(2775) <= a and b;
    layer0_outputs(2776) <= a and not b;
    layer0_outputs(2777) <= not b;
    layer0_outputs(2778) <= not b or a;
    layer0_outputs(2779) <= a xor b;
    layer0_outputs(2780) <= a and not b;
    layer0_outputs(2781) <= b and not a;
    layer0_outputs(2782) <= b;
    layer0_outputs(2783) <= not (a xor b);
    layer0_outputs(2784) <= a or b;
    layer0_outputs(2785) <= a;
    layer0_outputs(2786) <= not (a xor b);
    layer0_outputs(2787) <= not a;
    layer0_outputs(2788) <= not (a xor b);
    layer0_outputs(2789) <= not (a or b);
    layer0_outputs(2790) <= not (a or b);
    layer0_outputs(2791) <= b;
    layer0_outputs(2792) <= not a or b;
    layer0_outputs(2793) <= '0';
    layer0_outputs(2794) <= a or b;
    layer0_outputs(2795) <= a or b;
    layer0_outputs(2796) <= not b or a;
    layer0_outputs(2797) <= not (a or b);
    layer0_outputs(2798) <= not (a or b);
    layer0_outputs(2799) <= a;
    layer0_outputs(2800) <= not a or b;
    layer0_outputs(2801) <= not (a or b);
    layer0_outputs(2802) <= not b;
    layer0_outputs(2803) <= not (a or b);
    layer0_outputs(2804) <= not b or a;
    layer0_outputs(2805) <= a xor b;
    layer0_outputs(2806) <= not (a xor b);
    layer0_outputs(2807) <= a and not b;
    layer0_outputs(2808) <= a or b;
    layer0_outputs(2809) <= not (a or b);
    layer0_outputs(2810) <= '0';
    layer0_outputs(2811) <= not a;
    layer0_outputs(2812) <= a or b;
    layer0_outputs(2813) <= a and not b;
    layer0_outputs(2814) <= b and not a;
    layer0_outputs(2815) <= not b or a;
    layer0_outputs(2816) <= not b or a;
    layer0_outputs(2817) <= a and b;
    layer0_outputs(2818) <= a xor b;
    layer0_outputs(2819) <= not (a or b);
    layer0_outputs(2820) <= a;
    layer0_outputs(2821) <= a xor b;
    layer0_outputs(2822) <= not (a or b);
    layer0_outputs(2823) <= b;
    layer0_outputs(2824) <= not (a xor b);
    layer0_outputs(2825) <= not b or a;
    layer0_outputs(2826) <= a xor b;
    layer0_outputs(2827) <= not b or a;
    layer0_outputs(2828) <= not b or a;
    layer0_outputs(2829) <= a xor b;
    layer0_outputs(2830) <= a and not b;
    layer0_outputs(2831) <= not a;
    layer0_outputs(2832) <= b;
    layer0_outputs(2833) <= b;
    layer0_outputs(2834) <= a or b;
    layer0_outputs(2835) <= b;
    layer0_outputs(2836) <= not (a xor b);
    layer0_outputs(2837) <= not b;
    layer0_outputs(2838) <= not (a or b);
    layer0_outputs(2839) <= a and not b;
    layer0_outputs(2840) <= a or b;
    layer0_outputs(2841) <= not (a or b);
    layer0_outputs(2842) <= not a or b;
    layer0_outputs(2843) <= not b;
    layer0_outputs(2844) <= not a;
    layer0_outputs(2845) <= not (a xor b);
    layer0_outputs(2846) <= not (a xor b);
    layer0_outputs(2847) <= not (a or b);
    layer0_outputs(2848) <= not (a or b);
    layer0_outputs(2849) <= a xor b;
    layer0_outputs(2850) <= not b;
    layer0_outputs(2851) <= not b or a;
    layer0_outputs(2852) <= not (a or b);
    layer0_outputs(2853) <= a or b;
    layer0_outputs(2854) <= a or b;
    layer0_outputs(2855) <= '0';
    layer0_outputs(2856) <= not (a and b);
    layer0_outputs(2857) <= not (a or b);
    layer0_outputs(2858) <= not a;
    layer0_outputs(2859) <= not (a or b);
    layer0_outputs(2860) <= a xor b;
    layer0_outputs(2861) <= a or b;
    layer0_outputs(2862) <= not b or a;
    layer0_outputs(2863) <= not b or a;
    layer0_outputs(2864) <= not a;
    layer0_outputs(2865) <= a;
    layer0_outputs(2866) <= b;
    layer0_outputs(2867) <= not a or b;
    layer0_outputs(2868) <= b;
    layer0_outputs(2869) <= a;
    layer0_outputs(2870) <= a and not b;
    layer0_outputs(2871) <= b;
    layer0_outputs(2872) <= '1';
    layer0_outputs(2873) <= a and not b;
    layer0_outputs(2874) <= not (a or b);
    layer0_outputs(2875) <= not (a or b);
    layer0_outputs(2876) <= a;
    layer0_outputs(2877) <= a and b;
    layer0_outputs(2878) <= not (a or b);
    layer0_outputs(2879) <= not (a and b);
    layer0_outputs(2880) <= not a or b;
    layer0_outputs(2881) <= not (a or b);
    layer0_outputs(2882) <= not (a and b);
    layer0_outputs(2883) <= a;
    layer0_outputs(2884) <= a or b;
    layer0_outputs(2885) <= a xor b;
    layer0_outputs(2886) <= not (a xor b);
    layer0_outputs(2887) <= a or b;
    layer0_outputs(2888) <= a xor b;
    layer0_outputs(2889) <= a or b;
    layer0_outputs(2890) <= not a or b;
    layer0_outputs(2891) <= not a;
    layer0_outputs(2892) <= not a;
    layer0_outputs(2893) <= a and b;
    layer0_outputs(2894) <= not (a or b);
    layer0_outputs(2895) <= not b or a;
    layer0_outputs(2896) <= a xor b;
    layer0_outputs(2897) <= '1';
    layer0_outputs(2898) <= not (a xor b);
    layer0_outputs(2899) <= b;
    layer0_outputs(2900) <= not (a or b);
    layer0_outputs(2901) <= a xor b;
    layer0_outputs(2902) <= not a;
    layer0_outputs(2903) <= a;
    layer0_outputs(2904) <= a xor b;
    layer0_outputs(2905) <= a;
    layer0_outputs(2906) <= not b;
    layer0_outputs(2907) <= a or b;
    layer0_outputs(2908) <= not (a or b);
    layer0_outputs(2909) <= a xor b;
    layer0_outputs(2910) <= not (a xor b);
    layer0_outputs(2911) <= not a or b;
    layer0_outputs(2912) <= not a;
    layer0_outputs(2913) <= not (a or b);
    layer0_outputs(2914) <= not (a or b);
    layer0_outputs(2915) <= not b or a;
    layer0_outputs(2916) <= a or b;
    layer0_outputs(2917) <= a or b;
    layer0_outputs(2918) <= a or b;
    layer0_outputs(2919) <= not a;
    layer0_outputs(2920) <= not (a xor b);
    layer0_outputs(2921) <= not (a xor b);
    layer0_outputs(2922) <= not (a or b);
    layer0_outputs(2923) <= a and not b;
    layer0_outputs(2924) <= b;
    layer0_outputs(2925) <= '0';
    layer0_outputs(2926) <= not a or b;
    layer0_outputs(2927) <= not b or a;
    layer0_outputs(2928) <= not b;
    layer0_outputs(2929) <= not (a or b);
    layer0_outputs(2930) <= not (a or b);
    layer0_outputs(2931) <= a xor b;
    layer0_outputs(2932) <= a or b;
    layer0_outputs(2933) <= not b;
    layer0_outputs(2934) <= a or b;
    layer0_outputs(2935) <= not (a xor b);
    layer0_outputs(2936) <= not (a or b);
    layer0_outputs(2937) <= a or b;
    layer0_outputs(2938) <= not b or a;
    layer0_outputs(2939) <= not (a or b);
    layer0_outputs(2940) <= not a or b;
    layer0_outputs(2941) <= not b;
    layer0_outputs(2942) <= a or b;
    layer0_outputs(2943) <= a or b;
    layer0_outputs(2944) <= not (a or b);
    layer0_outputs(2945) <= not (a or b);
    layer0_outputs(2946) <= a xor b;
    layer0_outputs(2947) <= a and not b;
    layer0_outputs(2948) <= a or b;
    layer0_outputs(2949) <= a or b;
    layer0_outputs(2950) <= a and not b;
    layer0_outputs(2951) <= a and not b;
    layer0_outputs(2952) <= '0';
    layer0_outputs(2953) <= not b;
    layer0_outputs(2954) <= not (a xor b);
    layer0_outputs(2955) <= not (a or b);
    layer0_outputs(2956) <= not (a or b);
    layer0_outputs(2957) <= not (a or b);
    layer0_outputs(2958) <= b and not a;
    layer0_outputs(2959) <= a or b;
    layer0_outputs(2960) <= not a or b;
    layer0_outputs(2961) <= not (a or b);
    layer0_outputs(2962) <= '1';
    layer0_outputs(2963) <= not a;
    layer0_outputs(2964) <= a xor b;
    layer0_outputs(2965) <= not b;
    layer0_outputs(2966) <= not (a or b);
    layer0_outputs(2967) <= a and not b;
    layer0_outputs(2968) <= not (a or b);
    layer0_outputs(2969) <= a or b;
    layer0_outputs(2970) <= b and not a;
    layer0_outputs(2971) <= a and not b;
    layer0_outputs(2972) <= b and not a;
    layer0_outputs(2973) <= not (a or b);
    layer0_outputs(2974) <= not a;
    layer0_outputs(2975) <= a;
    layer0_outputs(2976) <= not b;
    layer0_outputs(2977) <= a and not b;
    layer0_outputs(2978) <= a or b;
    layer0_outputs(2979) <= not (a or b);
    layer0_outputs(2980) <= not b;
    layer0_outputs(2981) <= a or b;
    layer0_outputs(2982) <= not b;
    layer0_outputs(2983) <= a xor b;
    layer0_outputs(2984) <= not a or b;
    layer0_outputs(2985) <= not (a and b);
    layer0_outputs(2986) <= a or b;
    layer0_outputs(2987) <= a;
    layer0_outputs(2988) <= not (a or b);
    layer0_outputs(2989) <= b;
    layer0_outputs(2990) <= not (a or b);
    layer0_outputs(2991) <= not (a or b);
    layer0_outputs(2992) <= not (a xor b);
    layer0_outputs(2993) <= not b or a;
    layer0_outputs(2994) <= not a or b;
    layer0_outputs(2995) <= a or b;
    layer0_outputs(2996) <= not a;
    layer0_outputs(2997) <= not (a xor b);
    layer0_outputs(2998) <= a or b;
    layer0_outputs(2999) <= a or b;
    layer0_outputs(3000) <= a and not b;
    layer0_outputs(3001) <= a or b;
    layer0_outputs(3002) <= not b or a;
    layer0_outputs(3003) <= not a or b;
    layer0_outputs(3004) <= not b;
    layer0_outputs(3005) <= not b or a;
    layer0_outputs(3006) <= not a or b;
    layer0_outputs(3007) <= a;
    layer0_outputs(3008) <= a or b;
    layer0_outputs(3009) <= '0';
    layer0_outputs(3010) <= not (a xor b);
    layer0_outputs(3011) <= not (a or b);
    layer0_outputs(3012) <= a xor b;
    layer0_outputs(3013) <= not (a xor b);
    layer0_outputs(3014) <= b and not a;
    layer0_outputs(3015) <= a and not b;
    layer0_outputs(3016) <= a or b;
    layer0_outputs(3017) <= not b;
    layer0_outputs(3018) <= b and not a;
    layer0_outputs(3019) <= a xor b;
    layer0_outputs(3020) <= not b or a;
    layer0_outputs(3021) <= not (a and b);
    layer0_outputs(3022) <= a xor b;
    layer0_outputs(3023) <= not a;
    layer0_outputs(3024) <= not a or b;
    layer0_outputs(3025) <= a xor b;
    layer0_outputs(3026) <= a and not b;
    layer0_outputs(3027) <= b;
    layer0_outputs(3028) <= not (a or b);
    layer0_outputs(3029) <= a and not b;
    layer0_outputs(3030) <= b and not a;
    layer0_outputs(3031) <= a or b;
    layer0_outputs(3032) <= a;
    layer0_outputs(3033) <= not (a xor b);
    layer0_outputs(3034) <= '1';
    layer0_outputs(3035) <= a;
    layer0_outputs(3036) <= not b or a;
    layer0_outputs(3037) <= a or b;
    layer0_outputs(3038) <= '1';
    layer0_outputs(3039) <= a and not b;
    layer0_outputs(3040) <= a;
    layer0_outputs(3041) <= not (a or b);
    layer0_outputs(3042) <= a or b;
    layer0_outputs(3043) <= not a;
    layer0_outputs(3044) <= a or b;
    layer0_outputs(3045) <= a and not b;
    layer0_outputs(3046) <= not (a or b);
    layer0_outputs(3047) <= a or b;
    layer0_outputs(3048) <= a xor b;
    layer0_outputs(3049) <= not b;
    layer0_outputs(3050) <= a or b;
    layer0_outputs(3051) <= not (a or b);
    layer0_outputs(3052) <= not (a or b);
    layer0_outputs(3053) <= not (a or b);
    layer0_outputs(3054) <= not (a and b);
    layer0_outputs(3055) <= not (a or b);
    layer0_outputs(3056) <= b;
    layer0_outputs(3057) <= a;
    layer0_outputs(3058) <= a;
    layer0_outputs(3059) <= not a or b;
    layer0_outputs(3060) <= not (a or b);
    layer0_outputs(3061) <= not a or b;
    layer0_outputs(3062) <= a and not b;
    layer0_outputs(3063) <= not b or a;
    layer0_outputs(3064) <= not b;
    layer0_outputs(3065) <= a and not b;
    layer0_outputs(3066) <= not (a or b);
    layer0_outputs(3067) <= a;
    layer0_outputs(3068) <= a or b;
    layer0_outputs(3069) <= not b;
    layer0_outputs(3070) <= b and not a;
    layer0_outputs(3071) <= not a;
    layer0_outputs(3072) <= not (a xor b);
    layer0_outputs(3073) <= a or b;
    layer0_outputs(3074) <= a and b;
    layer0_outputs(3075) <= not (a and b);
    layer0_outputs(3076) <= not b;
    layer0_outputs(3077) <= b;
    layer0_outputs(3078) <= a xor b;
    layer0_outputs(3079) <= a and not b;
    layer0_outputs(3080) <= a or b;
    layer0_outputs(3081) <= not b or a;
    layer0_outputs(3082) <= a;
    layer0_outputs(3083) <= b;
    layer0_outputs(3084) <= not b;
    layer0_outputs(3085) <= not (a or b);
    layer0_outputs(3086) <= not (a or b);
    layer0_outputs(3087) <= not a;
    layer0_outputs(3088) <= not (a xor b);
    layer0_outputs(3089) <= not b or a;
    layer0_outputs(3090) <= a xor b;
    layer0_outputs(3091) <= b;
    layer0_outputs(3092) <= '1';
    layer0_outputs(3093) <= a or b;
    layer0_outputs(3094) <= not (a or b);
    layer0_outputs(3095) <= b;
    layer0_outputs(3096) <= b;
    layer0_outputs(3097) <= not a or b;
    layer0_outputs(3098) <= not (a or b);
    layer0_outputs(3099) <= not (a or b);
    layer0_outputs(3100) <= not b or a;
    layer0_outputs(3101) <= '0';
    layer0_outputs(3102) <= not b;
    layer0_outputs(3103) <= not (a and b);
    layer0_outputs(3104) <= a;
    layer0_outputs(3105) <= b;
    layer0_outputs(3106) <= a and b;
    layer0_outputs(3107) <= not (a or b);
    layer0_outputs(3108) <= not b or a;
    layer0_outputs(3109) <= not b or a;
    layer0_outputs(3110) <= a and not b;
    layer0_outputs(3111) <= not a;
    layer0_outputs(3112) <= a or b;
    layer0_outputs(3113) <= a or b;
    layer0_outputs(3114) <= b and not a;
    layer0_outputs(3115) <= not a or b;
    layer0_outputs(3116) <= '1';
    layer0_outputs(3117) <= a and not b;
    layer0_outputs(3118) <= not (a or b);
    layer0_outputs(3119) <= not a;
    layer0_outputs(3120) <= not (a or b);
    layer0_outputs(3121) <= a;
    layer0_outputs(3122) <= not a;
    layer0_outputs(3123) <= not (a xor b);
    layer0_outputs(3124) <= not (a or b);
    layer0_outputs(3125) <= a or b;
    layer0_outputs(3126) <= not (a or b);
    layer0_outputs(3127) <= a or b;
    layer0_outputs(3128) <= not a or b;
    layer0_outputs(3129) <= not (a or b);
    layer0_outputs(3130) <= not (a or b);
    layer0_outputs(3131) <= b and not a;
    layer0_outputs(3132) <= a;
    layer0_outputs(3133) <= a;
    layer0_outputs(3134) <= not b;
    layer0_outputs(3135) <= a;
    layer0_outputs(3136) <= b;
    layer0_outputs(3137) <= not (a xor b);
    layer0_outputs(3138) <= '0';
    layer0_outputs(3139) <= not (a or b);
    layer0_outputs(3140) <= a xor b;
    layer0_outputs(3141) <= a or b;
    layer0_outputs(3142) <= not (a and b);
    layer0_outputs(3143) <= b;
    layer0_outputs(3144) <= a xor b;
    layer0_outputs(3145) <= not (a or b);
    layer0_outputs(3146) <= a or b;
    layer0_outputs(3147) <= not b;
    layer0_outputs(3148) <= not b;
    layer0_outputs(3149) <= a or b;
    layer0_outputs(3150) <= b;
    layer0_outputs(3151) <= a or b;
    layer0_outputs(3152) <= not a;
    layer0_outputs(3153) <= a xor b;
    layer0_outputs(3154) <= b and not a;
    layer0_outputs(3155) <= a or b;
    layer0_outputs(3156) <= not (a or b);
    layer0_outputs(3157) <= a or b;
    layer0_outputs(3158) <= a xor b;
    layer0_outputs(3159) <= a xor b;
    layer0_outputs(3160) <= not (a or b);
    layer0_outputs(3161) <= not (a or b);
    layer0_outputs(3162) <= not a or b;
    layer0_outputs(3163) <= not (a or b);
    layer0_outputs(3164) <= a or b;
    layer0_outputs(3165) <= not b;
    layer0_outputs(3166) <= not a;
    layer0_outputs(3167) <= '1';
    layer0_outputs(3168) <= a;
    layer0_outputs(3169) <= b and not a;
    layer0_outputs(3170) <= a or b;
    layer0_outputs(3171) <= not (a or b);
    layer0_outputs(3172) <= a xor b;
    layer0_outputs(3173) <= a or b;
    layer0_outputs(3174) <= not (a or b);
    layer0_outputs(3175) <= a and not b;
    layer0_outputs(3176) <= a xor b;
    layer0_outputs(3177) <= not b;
    layer0_outputs(3178) <= not a;
    layer0_outputs(3179) <= a or b;
    layer0_outputs(3180) <= not a;
    layer0_outputs(3181) <= a xor b;
    layer0_outputs(3182) <= not (a or b);
    layer0_outputs(3183) <= not (a or b);
    layer0_outputs(3184) <= not (a or b);
    layer0_outputs(3185) <= a;
    layer0_outputs(3186) <= not (a or b);
    layer0_outputs(3187) <= a or b;
    layer0_outputs(3188) <= not b or a;
    layer0_outputs(3189) <= not (a or b);
    layer0_outputs(3190) <= not (a or b);
    layer0_outputs(3191) <= a or b;
    layer0_outputs(3192) <= not (a xor b);
    layer0_outputs(3193) <= not (a xor b);
    layer0_outputs(3194) <= '0';
    layer0_outputs(3195) <= not (a or b);
    layer0_outputs(3196) <= b and not a;
    layer0_outputs(3197) <= not (a or b);
    layer0_outputs(3198) <= not a;
    layer0_outputs(3199) <= not b or a;
    layer0_outputs(3200) <= not (a or b);
    layer0_outputs(3201) <= a;
    layer0_outputs(3202) <= not (a xor b);
    layer0_outputs(3203) <= not b;
    layer0_outputs(3204) <= a xor b;
    layer0_outputs(3205) <= a or b;
    layer0_outputs(3206) <= a or b;
    layer0_outputs(3207) <= not (a xor b);
    layer0_outputs(3208) <= a;
    layer0_outputs(3209) <= b;
    layer0_outputs(3210) <= not b or a;
    layer0_outputs(3211) <= b and not a;
    layer0_outputs(3212) <= not (a or b);
    layer0_outputs(3213) <= b;
    layer0_outputs(3214) <= not b or a;
    layer0_outputs(3215) <= b and not a;
    layer0_outputs(3216) <= a or b;
    layer0_outputs(3217) <= not (a or b);
    layer0_outputs(3218) <= not (a xor b);
    layer0_outputs(3219) <= a;
    layer0_outputs(3220) <= not (a or b);
    layer0_outputs(3221) <= not (a or b);
    layer0_outputs(3222) <= not b;
    layer0_outputs(3223) <= b;
    layer0_outputs(3224) <= a and not b;
    layer0_outputs(3225) <= a;
    layer0_outputs(3226) <= not a;
    layer0_outputs(3227) <= b;
    layer0_outputs(3228) <= b and not a;
    layer0_outputs(3229) <= not b;
    layer0_outputs(3230) <= a or b;
    layer0_outputs(3231) <= not b or a;
    layer0_outputs(3232) <= not a or b;
    layer0_outputs(3233) <= a or b;
    layer0_outputs(3234) <= not (a or b);
    layer0_outputs(3235) <= a and not b;
    layer0_outputs(3236) <= a or b;
    layer0_outputs(3237) <= not b or a;
    layer0_outputs(3238) <= not (a or b);
    layer0_outputs(3239) <= a and not b;
    layer0_outputs(3240) <= a or b;
    layer0_outputs(3241) <= not (a or b);
    layer0_outputs(3242) <= b and not a;
    layer0_outputs(3243) <= not (a or b);
    layer0_outputs(3244) <= not b or a;
    layer0_outputs(3245) <= not (a or b);
    layer0_outputs(3246) <= a xor b;
    layer0_outputs(3247) <= not (a or b);
    layer0_outputs(3248) <= a or b;
    layer0_outputs(3249) <= a;
    layer0_outputs(3250) <= '1';
    layer0_outputs(3251) <= b and not a;
    layer0_outputs(3252) <= not b or a;
    layer0_outputs(3253) <= a or b;
    layer0_outputs(3254) <= not a;
    layer0_outputs(3255) <= not (a or b);
    layer0_outputs(3256) <= not (a xor b);
    layer0_outputs(3257) <= not (a or b);
    layer0_outputs(3258) <= not b or a;
    layer0_outputs(3259) <= not b;
    layer0_outputs(3260) <= not (a xor b);
    layer0_outputs(3261) <= a xor b;
    layer0_outputs(3262) <= a xor b;
    layer0_outputs(3263) <= a xor b;
    layer0_outputs(3264) <= a;
    layer0_outputs(3265) <= not b;
    layer0_outputs(3266) <= a or b;
    layer0_outputs(3267) <= a;
    layer0_outputs(3268) <= not (a or b);
    layer0_outputs(3269) <= a;
    layer0_outputs(3270) <= not b;
    layer0_outputs(3271) <= b and not a;
    layer0_outputs(3272) <= not a;
    layer0_outputs(3273) <= a or b;
    layer0_outputs(3274) <= a and b;
    layer0_outputs(3275) <= a xor b;
    layer0_outputs(3276) <= not (a xor b);
    layer0_outputs(3277) <= not (a xor b);
    layer0_outputs(3278) <= not b or a;
    layer0_outputs(3279) <= not (a or b);
    layer0_outputs(3280) <= a xor b;
    layer0_outputs(3281) <= not (a or b);
    layer0_outputs(3282) <= a;
    layer0_outputs(3283) <= a or b;
    layer0_outputs(3284) <= a xor b;
    layer0_outputs(3285) <= a xor b;
    layer0_outputs(3286) <= a;
    layer0_outputs(3287) <= a xor b;
    layer0_outputs(3288) <= not (a or b);
    layer0_outputs(3289) <= a or b;
    layer0_outputs(3290) <= not (a xor b);
    layer0_outputs(3291) <= a xor b;
    layer0_outputs(3292) <= not (a or b);
    layer0_outputs(3293) <= not b;
    layer0_outputs(3294) <= not (a or b);
    layer0_outputs(3295) <= a xor b;
    layer0_outputs(3296) <= a xor b;
    layer0_outputs(3297) <= a or b;
    layer0_outputs(3298) <= a;
    layer0_outputs(3299) <= not a;
    layer0_outputs(3300) <= not b;
    layer0_outputs(3301) <= not (a or b);
    layer0_outputs(3302) <= not a;
    layer0_outputs(3303) <= b and not a;
    layer0_outputs(3304) <= not (a xor b);
    layer0_outputs(3305) <= a xor b;
    layer0_outputs(3306) <= not a;
    layer0_outputs(3307) <= not (a or b);
    layer0_outputs(3308) <= not (a xor b);
    layer0_outputs(3309) <= not b;
    layer0_outputs(3310) <= not (a xor b);
    layer0_outputs(3311) <= not (a xor b);
    layer0_outputs(3312) <= '0';
    layer0_outputs(3313) <= not (a or b);
    layer0_outputs(3314) <= not a or b;
    layer0_outputs(3315) <= not (a or b);
    layer0_outputs(3316) <= '0';
    layer0_outputs(3317) <= b and not a;
    layer0_outputs(3318) <= a and not b;
    layer0_outputs(3319) <= a or b;
    layer0_outputs(3320) <= not a;
    layer0_outputs(3321) <= '1';
    layer0_outputs(3322) <= b and not a;
    layer0_outputs(3323) <= '1';
    layer0_outputs(3324) <= not b;
    layer0_outputs(3325) <= b;
    layer0_outputs(3326) <= b and not a;
    layer0_outputs(3327) <= not b;
    layer0_outputs(3328) <= not (a or b);
    layer0_outputs(3329) <= not a;
    layer0_outputs(3330) <= b;
    layer0_outputs(3331) <= not (a or b);
    layer0_outputs(3332) <= a or b;
    layer0_outputs(3333) <= not (a xor b);
    layer0_outputs(3334) <= not (a xor b);
    layer0_outputs(3335) <= b;
    layer0_outputs(3336) <= not (a xor b);
    layer0_outputs(3337) <= b;
    layer0_outputs(3338) <= not b;
    layer0_outputs(3339) <= not (a or b);
    layer0_outputs(3340) <= a;
    layer0_outputs(3341) <= a;
    layer0_outputs(3342) <= not (a xor b);
    layer0_outputs(3343) <= a or b;
    layer0_outputs(3344) <= not b;
    layer0_outputs(3345) <= a xor b;
    layer0_outputs(3346) <= b and not a;
    layer0_outputs(3347) <= not (a or b);
    layer0_outputs(3348) <= not a;
    layer0_outputs(3349) <= b and not a;
    layer0_outputs(3350) <= not a;
    layer0_outputs(3351) <= a;
    layer0_outputs(3352) <= b;
    layer0_outputs(3353) <= a;
    layer0_outputs(3354) <= a or b;
    layer0_outputs(3355) <= b;
    layer0_outputs(3356) <= a xor b;
    layer0_outputs(3357) <= not (a xor b);
    layer0_outputs(3358) <= a or b;
    layer0_outputs(3359) <= a xor b;
    layer0_outputs(3360) <= not b or a;
    layer0_outputs(3361) <= not b;
    layer0_outputs(3362) <= a or b;
    layer0_outputs(3363) <= a and not b;
    layer0_outputs(3364) <= not (a or b);
    layer0_outputs(3365) <= not b or a;
    layer0_outputs(3366) <= not (a or b);
    layer0_outputs(3367) <= a or b;
    layer0_outputs(3368) <= a and b;
    layer0_outputs(3369) <= not (a and b);
    layer0_outputs(3370) <= not (a xor b);
    layer0_outputs(3371) <= not b or a;
    layer0_outputs(3372) <= not (a or b);
    layer0_outputs(3373) <= a or b;
    layer0_outputs(3374) <= not b or a;
    layer0_outputs(3375) <= a or b;
    layer0_outputs(3376) <= not a;
    layer0_outputs(3377) <= a or b;
    layer0_outputs(3378) <= a and not b;
    layer0_outputs(3379) <= not (a or b);
    layer0_outputs(3380) <= b;
    layer0_outputs(3381) <= a;
    layer0_outputs(3382) <= a;
    layer0_outputs(3383) <= not (a xor b);
    layer0_outputs(3384) <= not (a or b);
    layer0_outputs(3385) <= not (a xor b);
    layer0_outputs(3386) <= not b;
    layer0_outputs(3387) <= b and not a;
    layer0_outputs(3388) <= b and not a;
    layer0_outputs(3389) <= not b or a;
    layer0_outputs(3390) <= not (a or b);
    layer0_outputs(3391) <= a;
    layer0_outputs(3392) <= a xor b;
    layer0_outputs(3393) <= a or b;
    layer0_outputs(3394) <= not (a or b);
    layer0_outputs(3395) <= '1';
    layer0_outputs(3396) <= not b or a;
    layer0_outputs(3397) <= not b or a;
    layer0_outputs(3398) <= not b or a;
    layer0_outputs(3399) <= a or b;
    layer0_outputs(3400) <= not (a xor b);
    layer0_outputs(3401) <= a;
    layer0_outputs(3402) <= not a;
    layer0_outputs(3403) <= a or b;
    layer0_outputs(3404) <= b;
    layer0_outputs(3405) <= a;
    layer0_outputs(3406) <= a;
    layer0_outputs(3407) <= not (a or b);
    layer0_outputs(3408) <= b and not a;
    layer0_outputs(3409) <= a or b;
    layer0_outputs(3410) <= b and not a;
    layer0_outputs(3411) <= a and not b;
    layer0_outputs(3412) <= not (a or b);
    layer0_outputs(3413) <= a xor b;
    layer0_outputs(3414) <= '1';
    layer0_outputs(3415) <= a and not b;
    layer0_outputs(3416) <= a or b;
    layer0_outputs(3417) <= not b;
    layer0_outputs(3418) <= not a;
    layer0_outputs(3419) <= a or b;
    layer0_outputs(3420) <= a and not b;
    layer0_outputs(3421) <= b and not a;
    layer0_outputs(3422) <= a and b;
    layer0_outputs(3423) <= not a;
    layer0_outputs(3424) <= not a;
    layer0_outputs(3425) <= not b;
    layer0_outputs(3426) <= a or b;
    layer0_outputs(3427) <= a;
    layer0_outputs(3428) <= a or b;
    layer0_outputs(3429) <= not (a or b);
    layer0_outputs(3430) <= a xor b;
    layer0_outputs(3431) <= not b or a;
    layer0_outputs(3432) <= b;
    layer0_outputs(3433) <= b;
    layer0_outputs(3434) <= not b;
    layer0_outputs(3435) <= not (a or b);
    layer0_outputs(3436) <= b;
    layer0_outputs(3437) <= not b or a;
    layer0_outputs(3438) <= a or b;
    layer0_outputs(3439) <= a and b;
    layer0_outputs(3440) <= a or b;
    layer0_outputs(3441) <= b and not a;
    layer0_outputs(3442) <= not (a xor b);
    layer0_outputs(3443) <= b and not a;
    layer0_outputs(3444) <= b;
    layer0_outputs(3445) <= not a or b;
    layer0_outputs(3446) <= not a or b;
    layer0_outputs(3447) <= not (a or b);
    layer0_outputs(3448) <= not a;
    layer0_outputs(3449) <= not (a xor b);
    layer0_outputs(3450) <= not (a or b);
    layer0_outputs(3451) <= a and not b;
    layer0_outputs(3452) <= not (a or b);
    layer0_outputs(3453) <= a xor b;
    layer0_outputs(3454) <= not a;
    layer0_outputs(3455) <= a xor b;
    layer0_outputs(3456) <= a xor b;
    layer0_outputs(3457) <= not b or a;
    layer0_outputs(3458) <= b and not a;
    layer0_outputs(3459) <= a and not b;
    layer0_outputs(3460) <= not a or b;
    layer0_outputs(3461) <= a or b;
    layer0_outputs(3462) <= not a;
    layer0_outputs(3463) <= not (a or b);
    layer0_outputs(3464) <= a or b;
    layer0_outputs(3465) <= not a or b;
    layer0_outputs(3466) <= not (a xor b);
    layer0_outputs(3467) <= not a;
    layer0_outputs(3468) <= not b;
    layer0_outputs(3469) <= not (a and b);
    layer0_outputs(3470) <= not (a or b);
    layer0_outputs(3471) <= not b or a;
    layer0_outputs(3472) <= not a or b;
    layer0_outputs(3473) <= not (a and b);
    layer0_outputs(3474) <= not (a and b);
    layer0_outputs(3475) <= not (a or b);
    layer0_outputs(3476) <= not (a or b);
    layer0_outputs(3477) <= a or b;
    layer0_outputs(3478) <= a and not b;
    layer0_outputs(3479) <= a or b;
    layer0_outputs(3480) <= not (a and b);
    layer0_outputs(3481) <= a or b;
    layer0_outputs(3482) <= not (a xor b);
    layer0_outputs(3483) <= a xor b;
    layer0_outputs(3484) <= '1';
    layer0_outputs(3485) <= a or b;
    layer0_outputs(3486) <= a xor b;
    layer0_outputs(3487) <= b;
    layer0_outputs(3488) <= not a;
    layer0_outputs(3489) <= b and not a;
    layer0_outputs(3490) <= b;
    layer0_outputs(3491) <= not b or a;
    layer0_outputs(3492) <= a or b;
    layer0_outputs(3493) <= a or b;
    layer0_outputs(3494) <= not a;
    layer0_outputs(3495) <= not a;
    layer0_outputs(3496) <= a xor b;
    layer0_outputs(3497) <= a or b;
    layer0_outputs(3498) <= not b or a;
    layer0_outputs(3499) <= b and not a;
    layer0_outputs(3500) <= a and b;
    layer0_outputs(3501) <= a xor b;
    layer0_outputs(3502) <= a and not b;
    layer0_outputs(3503) <= a or b;
    layer0_outputs(3504) <= a and not b;
    layer0_outputs(3505) <= not (a or b);
    layer0_outputs(3506) <= not b;
    layer0_outputs(3507) <= not a or b;
    layer0_outputs(3508) <= not a;
    layer0_outputs(3509) <= a;
    layer0_outputs(3510) <= not a;
    layer0_outputs(3511) <= a or b;
    layer0_outputs(3512) <= not (a or b);
    layer0_outputs(3513) <= b;
    layer0_outputs(3514) <= a xor b;
    layer0_outputs(3515) <= not (a xor b);
    layer0_outputs(3516) <= not (a xor b);
    layer0_outputs(3517) <= a or b;
    layer0_outputs(3518) <= not a;
    layer0_outputs(3519) <= b and not a;
    layer0_outputs(3520) <= not b or a;
    layer0_outputs(3521) <= a;
    layer0_outputs(3522) <= b;
    layer0_outputs(3523) <= a xor b;
    layer0_outputs(3524) <= b and not a;
    layer0_outputs(3525) <= not a or b;
    layer0_outputs(3526) <= not (a or b);
    layer0_outputs(3527) <= not a or b;
    layer0_outputs(3528) <= not (a xor b);
    layer0_outputs(3529) <= not (a or b);
    layer0_outputs(3530) <= b and not a;
    layer0_outputs(3531) <= a xor b;
    layer0_outputs(3532) <= b and not a;
    layer0_outputs(3533) <= not a;
    layer0_outputs(3534) <= b;
    layer0_outputs(3535) <= not a or b;
    layer0_outputs(3536) <= not (a or b);
    layer0_outputs(3537) <= not (a or b);
    layer0_outputs(3538) <= not b;
    layer0_outputs(3539) <= a and not b;
    layer0_outputs(3540) <= not (a xor b);
    layer0_outputs(3541) <= not (a or b);
    layer0_outputs(3542) <= a or b;
    layer0_outputs(3543) <= not b;
    layer0_outputs(3544) <= a xor b;
    layer0_outputs(3545) <= not b;
    layer0_outputs(3546) <= a;
    layer0_outputs(3547) <= not b;
    layer0_outputs(3548) <= not b or a;
    layer0_outputs(3549) <= not a;
    layer0_outputs(3550) <= b and not a;
    layer0_outputs(3551) <= not a or b;
    layer0_outputs(3552) <= a or b;
    layer0_outputs(3553) <= a or b;
    layer0_outputs(3554) <= not (a xor b);
    layer0_outputs(3555) <= a;
    layer0_outputs(3556) <= not a;
    layer0_outputs(3557) <= a;
    layer0_outputs(3558) <= not (a or b);
    layer0_outputs(3559) <= a or b;
    layer0_outputs(3560) <= a;
    layer0_outputs(3561) <= a and not b;
    layer0_outputs(3562) <= not (a or b);
    layer0_outputs(3563) <= a xor b;
    layer0_outputs(3564) <= b;
    layer0_outputs(3565) <= a;
    layer0_outputs(3566) <= not (a or b);
    layer0_outputs(3567) <= not a;
    layer0_outputs(3568) <= a or b;
    layer0_outputs(3569) <= '1';
    layer0_outputs(3570) <= not (a or b);
    layer0_outputs(3571) <= a xor b;
    layer0_outputs(3572) <= a or b;
    layer0_outputs(3573) <= b;
    layer0_outputs(3574) <= not (a xor b);
    layer0_outputs(3575) <= not a;
    layer0_outputs(3576) <= a or b;
    layer0_outputs(3577) <= b and not a;
    layer0_outputs(3578) <= a or b;
    layer0_outputs(3579) <= a xor b;
    layer0_outputs(3580) <= a or b;
    layer0_outputs(3581) <= b;
    layer0_outputs(3582) <= a and not b;
    layer0_outputs(3583) <= not b or a;
    layer0_outputs(3584) <= not a;
    layer0_outputs(3585) <= a and not b;
    layer0_outputs(3586) <= not b;
    layer0_outputs(3587) <= a or b;
    layer0_outputs(3588) <= '1';
    layer0_outputs(3589) <= not a;
    layer0_outputs(3590) <= not (a xor b);
    layer0_outputs(3591) <= a and not b;
    layer0_outputs(3592) <= not (a xor b);
    layer0_outputs(3593) <= not a or b;
    layer0_outputs(3594) <= not a;
    layer0_outputs(3595) <= not a;
    layer0_outputs(3596) <= a and not b;
    layer0_outputs(3597) <= a and b;
    layer0_outputs(3598) <= not a or b;
    layer0_outputs(3599) <= not a;
    layer0_outputs(3600) <= not b or a;
    layer0_outputs(3601) <= not (a or b);
    layer0_outputs(3602) <= a or b;
    layer0_outputs(3603) <= b and not a;
    layer0_outputs(3604) <= not a;
    layer0_outputs(3605) <= a;
    layer0_outputs(3606) <= a or b;
    layer0_outputs(3607) <= not a;
    layer0_outputs(3608) <= a;
    layer0_outputs(3609) <= '1';
    layer0_outputs(3610) <= not a;
    layer0_outputs(3611) <= a xor b;
    layer0_outputs(3612) <= a;
    layer0_outputs(3613) <= '1';
    layer0_outputs(3614) <= a and not b;
    layer0_outputs(3615) <= b;
    layer0_outputs(3616) <= b and not a;
    layer0_outputs(3617) <= not (a and b);
    layer0_outputs(3618) <= a xor b;
    layer0_outputs(3619) <= a and not b;
    layer0_outputs(3620) <= not b;
    layer0_outputs(3621) <= a xor b;
    layer0_outputs(3622) <= a xor b;
    layer0_outputs(3623) <= not b;
    layer0_outputs(3624) <= a xor b;
    layer0_outputs(3625) <= a xor b;
    layer0_outputs(3626) <= not (a or b);
    layer0_outputs(3627) <= not a;
    layer0_outputs(3628) <= not b;
    layer0_outputs(3629) <= not b;
    layer0_outputs(3630) <= not (a or b);
    layer0_outputs(3631) <= '1';
    layer0_outputs(3632) <= a or b;
    layer0_outputs(3633) <= a or b;
    layer0_outputs(3634) <= a xor b;
    layer0_outputs(3635) <= a or b;
    layer0_outputs(3636) <= a;
    layer0_outputs(3637) <= b;
    layer0_outputs(3638) <= not b or a;
    layer0_outputs(3639) <= not b or a;
    layer0_outputs(3640) <= not (a and b);
    layer0_outputs(3641) <= not (a and b);
    layer0_outputs(3642) <= not (a or b);
    layer0_outputs(3643) <= not b or a;
    layer0_outputs(3644) <= not (a or b);
    layer0_outputs(3645) <= not (a or b);
    layer0_outputs(3646) <= a or b;
    layer0_outputs(3647) <= a or b;
    layer0_outputs(3648) <= a and not b;
    layer0_outputs(3649) <= not (a or b);
    layer0_outputs(3650) <= not (a xor b);
    layer0_outputs(3651) <= '1';
    layer0_outputs(3652) <= a and b;
    layer0_outputs(3653) <= b;
    layer0_outputs(3654) <= not (a or b);
    layer0_outputs(3655) <= not (a or b);
    layer0_outputs(3656) <= not b;
    layer0_outputs(3657) <= a;
    layer0_outputs(3658) <= a and b;
    layer0_outputs(3659) <= not (a or b);
    layer0_outputs(3660) <= a or b;
    layer0_outputs(3661) <= a;
    layer0_outputs(3662) <= a xor b;
    layer0_outputs(3663) <= not b;
    layer0_outputs(3664) <= not (a or b);
    layer0_outputs(3665) <= not a or b;
    layer0_outputs(3666) <= not b or a;
    layer0_outputs(3667) <= a;
    layer0_outputs(3668) <= not a or b;
    layer0_outputs(3669) <= not (a and b);
    layer0_outputs(3670) <= a xor b;
    layer0_outputs(3671) <= not (a and b);
    layer0_outputs(3672) <= not a;
    layer0_outputs(3673) <= a or b;
    layer0_outputs(3674) <= a xor b;
    layer0_outputs(3675) <= a or b;
    layer0_outputs(3676) <= a;
    layer0_outputs(3677) <= a;
    layer0_outputs(3678) <= a xor b;
    layer0_outputs(3679) <= not (a or b);
    layer0_outputs(3680) <= not (a and b);
    layer0_outputs(3681) <= not a or b;
    layer0_outputs(3682) <= a xor b;
    layer0_outputs(3683) <= '1';
    layer0_outputs(3684) <= not (a xor b);
    layer0_outputs(3685) <= not (a and b);
    layer0_outputs(3686) <= not b or a;
    layer0_outputs(3687) <= not b or a;
    layer0_outputs(3688) <= not (a xor b);
    layer0_outputs(3689) <= not b;
    layer0_outputs(3690) <= a or b;
    layer0_outputs(3691) <= not a or b;
    layer0_outputs(3692) <= b and not a;
    layer0_outputs(3693) <= a or b;
    layer0_outputs(3694) <= a or b;
    layer0_outputs(3695) <= b;
    layer0_outputs(3696) <= a or b;
    layer0_outputs(3697) <= not b or a;
    layer0_outputs(3698) <= b and not a;
    layer0_outputs(3699) <= not (a xor b);
    layer0_outputs(3700) <= not (a or b);
    layer0_outputs(3701) <= a or b;
    layer0_outputs(3702) <= a;
    layer0_outputs(3703) <= a xor b;
    layer0_outputs(3704) <= a or b;
    layer0_outputs(3705) <= not (a or b);
    layer0_outputs(3706) <= not a;
    layer0_outputs(3707) <= not a;
    layer0_outputs(3708) <= a or b;
    layer0_outputs(3709) <= a xor b;
    layer0_outputs(3710) <= not a or b;
    layer0_outputs(3711) <= not a or b;
    layer0_outputs(3712) <= a and b;
    layer0_outputs(3713) <= not (a or b);
    layer0_outputs(3714) <= a and not b;
    layer0_outputs(3715) <= a;
    layer0_outputs(3716) <= a xor b;
    layer0_outputs(3717) <= a or b;
    layer0_outputs(3718) <= not (a or b);
    layer0_outputs(3719) <= b and not a;
    layer0_outputs(3720) <= not a or b;
    layer0_outputs(3721) <= not (a or b);
    layer0_outputs(3722) <= not b;
    layer0_outputs(3723) <= a or b;
    layer0_outputs(3724) <= not (a or b);
    layer0_outputs(3725) <= not b;
    layer0_outputs(3726) <= not (a xor b);
    layer0_outputs(3727) <= b and not a;
    layer0_outputs(3728) <= a or b;
    layer0_outputs(3729) <= not (a or b);
    layer0_outputs(3730) <= not a;
    layer0_outputs(3731) <= not b or a;
    layer0_outputs(3732) <= b;
    layer0_outputs(3733) <= a and not b;
    layer0_outputs(3734) <= not a or b;
    layer0_outputs(3735) <= b;
    layer0_outputs(3736) <= a and not b;
    layer0_outputs(3737) <= not (a xor b);
    layer0_outputs(3738) <= not a or b;
    layer0_outputs(3739) <= a xor b;
    layer0_outputs(3740) <= not (a or b);
    layer0_outputs(3741) <= not (a or b);
    layer0_outputs(3742) <= not a or b;
    layer0_outputs(3743) <= not b;
    layer0_outputs(3744) <= b and not a;
    layer0_outputs(3745) <= not (a or b);
    layer0_outputs(3746) <= not (a or b);
    layer0_outputs(3747) <= a and not b;
    layer0_outputs(3748) <= a or b;
    layer0_outputs(3749) <= a xor b;
    layer0_outputs(3750) <= not b or a;
    layer0_outputs(3751) <= not b or a;
    layer0_outputs(3752) <= not b or a;
    layer0_outputs(3753) <= a xor b;
    layer0_outputs(3754) <= not a or b;
    layer0_outputs(3755) <= not b or a;
    layer0_outputs(3756) <= a;
    layer0_outputs(3757) <= '1';
    layer0_outputs(3758) <= b;
    layer0_outputs(3759) <= not b or a;
    layer0_outputs(3760) <= not (a or b);
    layer0_outputs(3761) <= a and not b;
    layer0_outputs(3762) <= not b;
    layer0_outputs(3763) <= b;
    layer0_outputs(3764) <= a and not b;
    layer0_outputs(3765) <= a or b;
    layer0_outputs(3766) <= not (a xor b);
    layer0_outputs(3767) <= '1';
    layer0_outputs(3768) <= a or b;
    layer0_outputs(3769) <= a or b;
    layer0_outputs(3770) <= not b;
    layer0_outputs(3771) <= b;
    layer0_outputs(3772) <= a and not b;
    layer0_outputs(3773) <= not (a xor b);
    layer0_outputs(3774) <= a or b;
    layer0_outputs(3775) <= a xor b;
    layer0_outputs(3776) <= not a or b;
    layer0_outputs(3777) <= a or b;
    layer0_outputs(3778) <= not a or b;
    layer0_outputs(3779) <= not (a xor b);
    layer0_outputs(3780) <= a and not b;
    layer0_outputs(3781) <= not a;
    layer0_outputs(3782) <= a or b;
    layer0_outputs(3783) <= not (a or b);
    layer0_outputs(3784) <= not a or b;
    layer0_outputs(3785) <= a or b;
    layer0_outputs(3786) <= '1';
    layer0_outputs(3787) <= a xor b;
    layer0_outputs(3788) <= a or b;
    layer0_outputs(3789) <= a and b;
    layer0_outputs(3790) <= a;
    layer0_outputs(3791) <= not (a xor b);
    layer0_outputs(3792) <= b and not a;
    layer0_outputs(3793) <= a and not b;
    layer0_outputs(3794) <= b;
    layer0_outputs(3795) <= not b;
    layer0_outputs(3796) <= a and not b;
    layer0_outputs(3797) <= not b or a;
    layer0_outputs(3798) <= not a or b;
    layer0_outputs(3799) <= a and not b;
    layer0_outputs(3800) <= a or b;
    layer0_outputs(3801) <= not b;
    layer0_outputs(3802) <= not a;
    layer0_outputs(3803) <= a or b;
    layer0_outputs(3804) <= a;
    layer0_outputs(3805) <= a or b;
    layer0_outputs(3806) <= a xor b;
    layer0_outputs(3807) <= a;
    layer0_outputs(3808) <= not (a and b);
    layer0_outputs(3809) <= not b;
    layer0_outputs(3810) <= a or b;
    layer0_outputs(3811) <= a;
    layer0_outputs(3812) <= not (a xor b);
    layer0_outputs(3813) <= b;
    layer0_outputs(3814) <= not b;
    layer0_outputs(3815) <= a and b;
    layer0_outputs(3816) <= a or b;
    layer0_outputs(3817) <= not (a xor b);
    layer0_outputs(3818) <= b;
    layer0_outputs(3819) <= not a;
    layer0_outputs(3820) <= b;
    layer0_outputs(3821) <= not (a or b);
    layer0_outputs(3822) <= a and not b;
    layer0_outputs(3823) <= not b;
    layer0_outputs(3824) <= a and not b;
    layer0_outputs(3825) <= a xor b;
    layer0_outputs(3826) <= a or b;
    layer0_outputs(3827) <= not a or b;
    layer0_outputs(3828) <= a and not b;
    layer0_outputs(3829) <= not (a or b);
    layer0_outputs(3830) <= a;
    layer0_outputs(3831) <= a or b;
    layer0_outputs(3832) <= not a or b;
    layer0_outputs(3833) <= a or b;
    layer0_outputs(3834) <= not (a or b);
    layer0_outputs(3835) <= b and not a;
    layer0_outputs(3836) <= not a;
    layer0_outputs(3837) <= not b;
    layer0_outputs(3838) <= not b;
    layer0_outputs(3839) <= not (a xor b);
    layer0_outputs(3840) <= not (a or b);
    layer0_outputs(3841) <= a or b;
    layer0_outputs(3842) <= a xor b;
    layer0_outputs(3843) <= a or b;
    layer0_outputs(3844) <= b and not a;
    layer0_outputs(3845) <= b;
    layer0_outputs(3846) <= a or b;
    layer0_outputs(3847) <= a xor b;
    layer0_outputs(3848) <= a and not b;
    layer0_outputs(3849) <= a and not b;
    layer0_outputs(3850) <= a or b;
    layer0_outputs(3851) <= a;
    layer0_outputs(3852) <= not a;
    layer0_outputs(3853) <= b;
    layer0_outputs(3854) <= a or b;
    layer0_outputs(3855) <= a or b;
    layer0_outputs(3856) <= a or b;
    layer0_outputs(3857) <= not b;
    layer0_outputs(3858) <= not (a or b);
    layer0_outputs(3859) <= not (a or b);
    layer0_outputs(3860) <= not a or b;
    layer0_outputs(3861) <= a;
    layer0_outputs(3862) <= a;
    layer0_outputs(3863) <= not a;
    layer0_outputs(3864) <= not a;
    layer0_outputs(3865) <= not (a or b);
    layer0_outputs(3866) <= a xor b;
    layer0_outputs(3867) <= b and not a;
    layer0_outputs(3868) <= a or b;
    layer0_outputs(3869) <= a xor b;
    layer0_outputs(3870) <= a xor b;
    layer0_outputs(3871) <= a or b;
    layer0_outputs(3872) <= not a or b;
    layer0_outputs(3873) <= not a or b;
    layer0_outputs(3874) <= a or b;
    layer0_outputs(3875) <= b and not a;
    layer0_outputs(3876) <= a or b;
    layer0_outputs(3877) <= not (a xor b);
    layer0_outputs(3878) <= not b;
    layer0_outputs(3879) <= a or b;
    layer0_outputs(3880) <= a xor b;
    layer0_outputs(3881) <= a xor b;
    layer0_outputs(3882) <= a;
    layer0_outputs(3883) <= '0';
    layer0_outputs(3884) <= a;
    layer0_outputs(3885) <= a and b;
    layer0_outputs(3886) <= not b or a;
    layer0_outputs(3887) <= not (a and b);
    layer0_outputs(3888) <= not (a or b);
    layer0_outputs(3889) <= not a;
    layer0_outputs(3890) <= not a;
    layer0_outputs(3891) <= not (a or b);
    layer0_outputs(3892) <= not (a or b);
    layer0_outputs(3893) <= not (a and b);
    layer0_outputs(3894) <= not (a or b);
    layer0_outputs(3895) <= a or b;
    layer0_outputs(3896) <= not (a xor b);
    layer0_outputs(3897) <= not (a or b);
    layer0_outputs(3898) <= b and not a;
    layer0_outputs(3899) <= not (a xor b);
    layer0_outputs(3900) <= not (a or b);
    layer0_outputs(3901) <= b;
    layer0_outputs(3902) <= not (a or b);
    layer0_outputs(3903) <= not (a xor b);
    layer0_outputs(3904) <= '0';
    layer0_outputs(3905) <= a;
    layer0_outputs(3906) <= a xor b;
    layer0_outputs(3907) <= not a;
    layer0_outputs(3908) <= not (a or b);
    layer0_outputs(3909) <= a or b;
    layer0_outputs(3910) <= b;
    layer0_outputs(3911) <= a or b;
    layer0_outputs(3912) <= a;
    layer0_outputs(3913) <= not a;
    layer0_outputs(3914) <= a or b;
    layer0_outputs(3915) <= a xor b;
    layer0_outputs(3916) <= not (a or b);
    layer0_outputs(3917) <= b;
    layer0_outputs(3918) <= b;
    layer0_outputs(3919) <= not (a or b);
    layer0_outputs(3920) <= not a or b;
    layer0_outputs(3921) <= a or b;
    layer0_outputs(3922) <= not (a or b);
    layer0_outputs(3923) <= not (a or b);
    layer0_outputs(3924) <= b;
    layer0_outputs(3925) <= a and not b;
    layer0_outputs(3926) <= a xor b;
    layer0_outputs(3927) <= b and not a;
    layer0_outputs(3928) <= not a;
    layer0_outputs(3929) <= not b or a;
    layer0_outputs(3930) <= a and not b;
    layer0_outputs(3931) <= not (a or b);
    layer0_outputs(3932) <= a xor b;
    layer0_outputs(3933) <= a and not b;
    layer0_outputs(3934) <= not b or a;
    layer0_outputs(3935) <= not (a or b);
    layer0_outputs(3936) <= not (a or b);
    layer0_outputs(3937) <= b;
    layer0_outputs(3938) <= not (a or b);
    layer0_outputs(3939) <= a or b;
    layer0_outputs(3940) <= not (a and b);
    layer0_outputs(3941) <= a xor b;
    layer0_outputs(3942) <= '0';
    layer0_outputs(3943) <= not (a or b);
    layer0_outputs(3944) <= not (a or b);
    layer0_outputs(3945) <= not b;
    layer0_outputs(3946) <= not b or a;
    layer0_outputs(3947) <= a and not b;
    layer0_outputs(3948) <= a and b;
    layer0_outputs(3949) <= b and not a;
    layer0_outputs(3950) <= b and not a;
    layer0_outputs(3951) <= a xor b;
    layer0_outputs(3952) <= not b;
    layer0_outputs(3953) <= not (a or b);
    layer0_outputs(3954) <= not b;
    layer0_outputs(3955) <= not (a and b);
    layer0_outputs(3956) <= a or b;
    layer0_outputs(3957) <= a and b;
    layer0_outputs(3958) <= a and not b;
    layer0_outputs(3959) <= not (a or b);
    layer0_outputs(3960) <= a;
    layer0_outputs(3961) <= a or b;
    layer0_outputs(3962) <= b and not a;
    layer0_outputs(3963) <= not (a xor b);
    layer0_outputs(3964) <= not b;
    layer0_outputs(3965) <= a xor b;
    layer0_outputs(3966) <= not a or b;
    layer0_outputs(3967) <= a or b;
    layer0_outputs(3968) <= a and not b;
    layer0_outputs(3969) <= a or b;
    layer0_outputs(3970) <= a;
    layer0_outputs(3971) <= a or b;
    layer0_outputs(3972) <= a or b;
    layer0_outputs(3973) <= not (a or b);
    layer0_outputs(3974) <= a or b;
    layer0_outputs(3975) <= a and not b;
    layer0_outputs(3976) <= not (a xor b);
    layer0_outputs(3977) <= a or b;
    layer0_outputs(3978) <= not b;
    layer0_outputs(3979) <= '1';
    layer0_outputs(3980) <= b;
    layer0_outputs(3981) <= not (a and b);
    layer0_outputs(3982) <= '0';
    layer0_outputs(3983) <= b;
    layer0_outputs(3984) <= a or b;
    layer0_outputs(3985) <= not (a or b);
    layer0_outputs(3986) <= not (a or b);
    layer0_outputs(3987) <= not (a xor b);
    layer0_outputs(3988) <= not (a or b);
    layer0_outputs(3989) <= not a;
    layer0_outputs(3990) <= a or b;
    layer0_outputs(3991) <= not b;
    layer0_outputs(3992) <= a and not b;
    layer0_outputs(3993) <= not a or b;
    layer0_outputs(3994) <= a or b;
    layer0_outputs(3995) <= not (a or b);
    layer0_outputs(3996) <= b and not a;
    layer0_outputs(3997) <= a or b;
    layer0_outputs(3998) <= not b or a;
    layer0_outputs(3999) <= not b;
    layer0_outputs(4000) <= a and not b;
    layer0_outputs(4001) <= b and not a;
    layer0_outputs(4002) <= b and not a;
    layer0_outputs(4003) <= not b;
    layer0_outputs(4004) <= not a or b;
    layer0_outputs(4005) <= not (a or b);
    layer0_outputs(4006) <= not b;
    layer0_outputs(4007) <= b;
    layer0_outputs(4008) <= a;
    layer0_outputs(4009) <= not a or b;
    layer0_outputs(4010) <= a;
    layer0_outputs(4011) <= a;
    layer0_outputs(4012) <= not (a xor b);
    layer0_outputs(4013) <= a;
    layer0_outputs(4014) <= not (a or b);
    layer0_outputs(4015) <= not (a or b);
    layer0_outputs(4016) <= not (a and b);
    layer0_outputs(4017) <= not b;
    layer0_outputs(4018) <= not (a or b);
    layer0_outputs(4019) <= a or b;
    layer0_outputs(4020) <= a;
    layer0_outputs(4021) <= a and not b;
    layer0_outputs(4022) <= not a or b;
    layer0_outputs(4023) <= a;
    layer0_outputs(4024) <= a or b;
    layer0_outputs(4025) <= a or b;
    layer0_outputs(4026) <= a and not b;
    layer0_outputs(4027) <= a;
    layer0_outputs(4028) <= a and not b;
    layer0_outputs(4029) <= a or b;
    layer0_outputs(4030) <= not b;
    layer0_outputs(4031) <= not (a xor b);
    layer0_outputs(4032) <= not (a or b);
    layer0_outputs(4033) <= a and not b;
    layer0_outputs(4034) <= b;
    layer0_outputs(4035) <= not a;
    layer0_outputs(4036) <= not (a xor b);
    layer0_outputs(4037) <= a;
    layer0_outputs(4038) <= not (a or b);
    layer0_outputs(4039) <= not (a and b);
    layer0_outputs(4040) <= not (a or b);
    layer0_outputs(4041) <= not (a xor b);
    layer0_outputs(4042) <= b and not a;
    layer0_outputs(4043) <= not b;
    layer0_outputs(4044) <= not a or b;
    layer0_outputs(4045) <= b and not a;
    layer0_outputs(4046) <= a;
    layer0_outputs(4047) <= a and not b;
    layer0_outputs(4048) <= '1';
    layer0_outputs(4049) <= a;
    layer0_outputs(4050) <= a or b;
    layer0_outputs(4051) <= not a;
    layer0_outputs(4052) <= not (a or b);
    layer0_outputs(4053) <= not (a or b);
    layer0_outputs(4054) <= not (a xor b);
    layer0_outputs(4055) <= a and b;
    layer0_outputs(4056) <= not (a or b);
    layer0_outputs(4057) <= not (a xor b);
    layer0_outputs(4058) <= not (a or b);
    layer0_outputs(4059) <= a or b;
    layer0_outputs(4060) <= not (a xor b);
    layer0_outputs(4061) <= not (a or b);
    layer0_outputs(4062) <= '1';
    layer0_outputs(4063) <= not (a or b);
    layer0_outputs(4064) <= not (a or b);
    layer0_outputs(4065) <= not b or a;
    layer0_outputs(4066) <= not b;
    layer0_outputs(4067) <= not a or b;
    layer0_outputs(4068) <= b and not a;
    layer0_outputs(4069) <= '0';
    layer0_outputs(4070) <= not (a xor b);
    layer0_outputs(4071) <= a or b;
    layer0_outputs(4072) <= a xor b;
    layer0_outputs(4073) <= not (a or b);
    layer0_outputs(4074) <= '1';
    layer0_outputs(4075) <= not (a or b);
    layer0_outputs(4076) <= a xor b;
    layer0_outputs(4077) <= not (a or b);
    layer0_outputs(4078) <= b;
    layer0_outputs(4079) <= not a or b;
    layer0_outputs(4080) <= a or b;
    layer0_outputs(4081) <= b;
    layer0_outputs(4082) <= not (a or b);
    layer0_outputs(4083) <= not b or a;
    layer0_outputs(4084) <= not b;
    layer0_outputs(4085) <= not b;
    layer0_outputs(4086) <= not (a or b);
    layer0_outputs(4087) <= not (a or b);
    layer0_outputs(4088) <= not a or b;
    layer0_outputs(4089) <= b;
    layer0_outputs(4090) <= a xor b;
    layer0_outputs(4091) <= not a or b;
    layer0_outputs(4092) <= b;
    layer0_outputs(4093) <= not (a or b);
    layer0_outputs(4094) <= not (a xor b);
    layer0_outputs(4095) <= not (a or b);
    layer0_outputs(4096) <= a and not b;
    layer0_outputs(4097) <= b and not a;
    layer0_outputs(4098) <= not b;
    layer0_outputs(4099) <= not a;
    layer0_outputs(4100) <= a;
    layer0_outputs(4101) <= not (a or b);
    layer0_outputs(4102) <= a or b;
    layer0_outputs(4103) <= not b or a;
    layer0_outputs(4104) <= not (a or b);
    layer0_outputs(4105) <= not (a or b);
    layer0_outputs(4106) <= b and not a;
    layer0_outputs(4107) <= not (a xor b);
    layer0_outputs(4108) <= not (a or b);
    layer0_outputs(4109) <= not a;
    layer0_outputs(4110) <= a;
    layer0_outputs(4111) <= '1';
    layer0_outputs(4112) <= not a;
    layer0_outputs(4113) <= b;
    layer0_outputs(4114) <= not (a xor b);
    layer0_outputs(4115) <= not a or b;
    layer0_outputs(4116) <= a;
    layer0_outputs(4117) <= b;
    layer0_outputs(4118) <= not b or a;
    layer0_outputs(4119) <= a or b;
    layer0_outputs(4120) <= not (a xor b);
    layer0_outputs(4121) <= not (a or b);
    layer0_outputs(4122) <= a and not b;
    layer0_outputs(4123) <= b and not a;
    layer0_outputs(4124) <= '1';
    layer0_outputs(4125) <= not b or a;
    layer0_outputs(4126) <= a and b;
    layer0_outputs(4127) <= not b;
    layer0_outputs(4128) <= b and not a;
    layer0_outputs(4129) <= not a or b;
    layer0_outputs(4130) <= not b or a;
    layer0_outputs(4131) <= not b;
    layer0_outputs(4132) <= b and not a;
    layer0_outputs(4133) <= a or b;
    layer0_outputs(4134) <= not (a xor b);
    layer0_outputs(4135) <= b and not a;
    layer0_outputs(4136) <= not (a xor b);
    layer0_outputs(4137) <= not b;
    layer0_outputs(4138) <= b and not a;
    layer0_outputs(4139) <= b;
    layer0_outputs(4140) <= a and b;
    layer0_outputs(4141) <= not (a or b);
    layer0_outputs(4142) <= not a;
    layer0_outputs(4143) <= not (a and b);
    layer0_outputs(4144) <= b;
    layer0_outputs(4145) <= b and not a;
    layer0_outputs(4146) <= a xor b;
    layer0_outputs(4147) <= not (a and b);
    layer0_outputs(4148) <= a and not b;
    layer0_outputs(4149) <= a and b;
    layer0_outputs(4150) <= not (a or b);
    layer0_outputs(4151) <= not b or a;
    layer0_outputs(4152) <= not a or b;
    layer0_outputs(4153) <= a or b;
    layer0_outputs(4154) <= not b;
    layer0_outputs(4155) <= not (a or b);
    layer0_outputs(4156) <= b and not a;
    layer0_outputs(4157) <= not b or a;
    layer0_outputs(4158) <= b;
    layer0_outputs(4159) <= not b;
    layer0_outputs(4160) <= not (a xor b);
    layer0_outputs(4161) <= not (a or b);
    layer0_outputs(4162) <= not a;
    layer0_outputs(4163) <= a or b;
    layer0_outputs(4164) <= a;
    layer0_outputs(4165) <= not a;
    layer0_outputs(4166) <= not (a or b);
    layer0_outputs(4167) <= not a;
    layer0_outputs(4168) <= a xor b;
    layer0_outputs(4169) <= a or b;
    layer0_outputs(4170) <= a and not b;
    layer0_outputs(4171) <= not a or b;
    layer0_outputs(4172) <= a or b;
    layer0_outputs(4173) <= a;
    layer0_outputs(4174) <= a or b;
    layer0_outputs(4175) <= not a;
    layer0_outputs(4176) <= not (a or b);
    layer0_outputs(4177) <= not b or a;
    layer0_outputs(4178) <= not a;
    layer0_outputs(4179) <= a;
    layer0_outputs(4180) <= a and not b;
    layer0_outputs(4181) <= not b or a;
    layer0_outputs(4182) <= not b;
    layer0_outputs(4183) <= b;
    layer0_outputs(4184) <= a or b;
    layer0_outputs(4185) <= not b;
    layer0_outputs(4186) <= not (a or b);
    layer0_outputs(4187) <= '1';
    layer0_outputs(4188) <= not a or b;
    layer0_outputs(4189) <= not (a or b);
    layer0_outputs(4190) <= not a or b;
    layer0_outputs(4191) <= not (a xor b);
    layer0_outputs(4192) <= b;
    layer0_outputs(4193) <= a and b;
    layer0_outputs(4194) <= not a or b;
    layer0_outputs(4195) <= b;
    layer0_outputs(4196) <= not a or b;
    layer0_outputs(4197) <= a or b;
    layer0_outputs(4198) <= not b;
    layer0_outputs(4199) <= not (a xor b);
    layer0_outputs(4200) <= not a or b;
    layer0_outputs(4201) <= a or b;
    layer0_outputs(4202) <= a or b;
    layer0_outputs(4203) <= not (a xor b);
    layer0_outputs(4204) <= a;
    layer0_outputs(4205) <= not b;
    layer0_outputs(4206) <= not (a or b);
    layer0_outputs(4207) <= a;
    layer0_outputs(4208) <= b and not a;
    layer0_outputs(4209) <= not b;
    layer0_outputs(4210) <= not (a xor b);
    layer0_outputs(4211) <= a xor b;
    layer0_outputs(4212) <= a xor b;
    layer0_outputs(4213) <= not b;
    layer0_outputs(4214) <= a or b;
    layer0_outputs(4215) <= not (a or b);
    layer0_outputs(4216) <= not a;
    layer0_outputs(4217) <= a or b;
    layer0_outputs(4218) <= not (a xor b);
    layer0_outputs(4219) <= not b or a;
    layer0_outputs(4220) <= not b;
    layer0_outputs(4221) <= a and b;
    layer0_outputs(4222) <= a;
    layer0_outputs(4223) <= not b or a;
    layer0_outputs(4224) <= not b or a;
    layer0_outputs(4225) <= b;
    layer0_outputs(4226) <= a xor b;
    layer0_outputs(4227) <= a xor b;
    layer0_outputs(4228) <= not b;
    layer0_outputs(4229) <= not a;
    layer0_outputs(4230) <= a and not b;
    layer0_outputs(4231) <= not b;
    layer0_outputs(4232) <= not a;
    layer0_outputs(4233) <= not (a and b);
    layer0_outputs(4234) <= a xor b;
    layer0_outputs(4235) <= not (a or b);
    layer0_outputs(4236) <= a and not b;
    layer0_outputs(4237) <= b;
    layer0_outputs(4238) <= a or b;
    layer0_outputs(4239) <= a xor b;
    layer0_outputs(4240) <= not (a or b);
    layer0_outputs(4241) <= a and not b;
    layer0_outputs(4242) <= a or b;
    layer0_outputs(4243) <= a and not b;
    layer0_outputs(4244) <= not (a xor b);
    layer0_outputs(4245) <= not b or a;
    layer0_outputs(4246) <= b and not a;
    layer0_outputs(4247) <= a or b;
    layer0_outputs(4248) <= a xor b;
    layer0_outputs(4249) <= b;
    layer0_outputs(4250) <= not (a xor b);
    layer0_outputs(4251) <= not (a or b);
    layer0_outputs(4252) <= not a or b;
    layer0_outputs(4253) <= '1';
    layer0_outputs(4254) <= a or b;
    layer0_outputs(4255) <= not (a xor b);
    layer0_outputs(4256) <= not a or b;
    layer0_outputs(4257) <= not (a or b);
    layer0_outputs(4258) <= b and not a;
    layer0_outputs(4259) <= a and not b;
    layer0_outputs(4260) <= '0';
    layer0_outputs(4261) <= a and not b;
    layer0_outputs(4262) <= b;
    layer0_outputs(4263) <= b and not a;
    layer0_outputs(4264) <= not (a or b);
    layer0_outputs(4265) <= not a or b;
    layer0_outputs(4266) <= not a;
    layer0_outputs(4267) <= b and not a;
    layer0_outputs(4268) <= b;
    layer0_outputs(4269) <= b and not a;
    layer0_outputs(4270) <= not a or b;
    layer0_outputs(4271) <= not a or b;
    layer0_outputs(4272) <= not (a xor b);
    layer0_outputs(4273) <= a or b;
    layer0_outputs(4274) <= a or b;
    layer0_outputs(4275) <= '1';
    layer0_outputs(4276) <= a or b;
    layer0_outputs(4277) <= not b or a;
    layer0_outputs(4278) <= a and not b;
    layer0_outputs(4279) <= not a or b;
    layer0_outputs(4280) <= not a;
    layer0_outputs(4281) <= not a;
    layer0_outputs(4282) <= not (a or b);
    layer0_outputs(4283) <= '0';
    layer0_outputs(4284) <= b and not a;
    layer0_outputs(4285) <= not (a xor b);
    layer0_outputs(4286) <= b;
    layer0_outputs(4287) <= a or b;
    layer0_outputs(4288) <= a or b;
    layer0_outputs(4289) <= b and not a;
    layer0_outputs(4290) <= not b;
    layer0_outputs(4291) <= not a;
    layer0_outputs(4292) <= a or b;
    layer0_outputs(4293) <= b;
    layer0_outputs(4294) <= not b;
    layer0_outputs(4295) <= a or b;
    layer0_outputs(4296) <= b;
    layer0_outputs(4297) <= b;
    layer0_outputs(4298) <= b;
    layer0_outputs(4299) <= not (a xor b);
    layer0_outputs(4300) <= not a;
    layer0_outputs(4301) <= b;
    layer0_outputs(4302) <= not (a or b);
    layer0_outputs(4303) <= b;
    layer0_outputs(4304) <= a xor b;
    layer0_outputs(4305) <= not (a and b);
    layer0_outputs(4306) <= not b or a;
    layer0_outputs(4307) <= a and b;
    layer0_outputs(4308) <= not (a or b);
    layer0_outputs(4309) <= not b or a;
    layer0_outputs(4310) <= not b;
    layer0_outputs(4311) <= not (a and b);
    layer0_outputs(4312) <= a and not b;
    layer0_outputs(4313) <= not (a xor b);
    layer0_outputs(4314) <= a;
    layer0_outputs(4315) <= not b;
    layer0_outputs(4316) <= not (a xor b);
    layer0_outputs(4317) <= not b or a;
    layer0_outputs(4318) <= not a or b;
    layer0_outputs(4319) <= not a or b;
    layer0_outputs(4320) <= a xor b;
    layer0_outputs(4321) <= b;
    layer0_outputs(4322) <= a or b;
    layer0_outputs(4323) <= b and not a;
    layer0_outputs(4324) <= not (a and b);
    layer0_outputs(4325) <= a;
    layer0_outputs(4326) <= a and not b;
    layer0_outputs(4327) <= not a or b;
    layer0_outputs(4328) <= not b;
    layer0_outputs(4329) <= a xor b;
    layer0_outputs(4330) <= a and not b;
    layer0_outputs(4331) <= not (a xor b);
    layer0_outputs(4332) <= a and not b;
    layer0_outputs(4333) <= b;
    layer0_outputs(4334) <= a or b;
    layer0_outputs(4335) <= not a or b;
    layer0_outputs(4336) <= not (a or b);
    layer0_outputs(4337) <= b and not a;
    layer0_outputs(4338) <= not a or b;
    layer0_outputs(4339) <= a xor b;
    layer0_outputs(4340) <= a or b;
    layer0_outputs(4341) <= not (a xor b);
    layer0_outputs(4342) <= '1';
    layer0_outputs(4343) <= not (a or b);
    layer0_outputs(4344) <= not a or b;
    layer0_outputs(4345) <= not (a or b);
    layer0_outputs(4346) <= a and b;
    layer0_outputs(4347) <= a and not b;
    layer0_outputs(4348) <= not a or b;
    layer0_outputs(4349) <= a and b;
    layer0_outputs(4350) <= not (a or b);
    layer0_outputs(4351) <= a xor b;
    layer0_outputs(4352) <= not a;
    layer0_outputs(4353) <= not (a and b);
    layer0_outputs(4354) <= not (a or b);
    layer0_outputs(4355) <= a or b;
    layer0_outputs(4356) <= a or b;
    layer0_outputs(4357) <= not (a or b);
    layer0_outputs(4358) <= a or b;
    layer0_outputs(4359) <= a and not b;
    layer0_outputs(4360) <= not (a or b);
    layer0_outputs(4361) <= a or b;
    layer0_outputs(4362) <= not b;
    layer0_outputs(4363) <= b;
    layer0_outputs(4364) <= not (a or b);
    layer0_outputs(4365) <= b and not a;
    layer0_outputs(4366) <= a and not b;
    layer0_outputs(4367) <= not (a or b);
    layer0_outputs(4368) <= not a or b;
    layer0_outputs(4369) <= a and not b;
    layer0_outputs(4370) <= b;
    layer0_outputs(4371) <= not a or b;
    layer0_outputs(4372) <= a or b;
    layer0_outputs(4373) <= a;
    layer0_outputs(4374) <= not (a xor b);
    layer0_outputs(4375) <= a xor b;
    layer0_outputs(4376) <= not (a xor b);
    layer0_outputs(4377) <= not a;
    layer0_outputs(4378) <= not (a xor b);
    layer0_outputs(4379) <= b and not a;
    layer0_outputs(4380) <= a or b;
    layer0_outputs(4381) <= a or b;
    layer0_outputs(4382) <= a xor b;
    layer0_outputs(4383) <= not a;
    layer0_outputs(4384) <= not (a or b);
    layer0_outputs(4385) <= a or b;
    layer0_outputs(4386) <= not (a or b);
    layer0_outputs(4387) <= not b;
    layer0_outputs(4388) <= b and not a;
    layer0_outputs(4389) <= not (a or b);
    layer0_outputs(4390) <= not a;
    layer0_outputs(4391) <= b;
    layer0_outputs(4392) <= a and not b;
    layer0_outputs(4393) <= a or b;
    layer0_outputs(4394) <= a or b;
    layer0_outputs(4395) <= not (a or b);
    layer0_outputs(4396) <= b and not a;
    layer0_outputs(4397) <= b and not a;
    layer0_outputs(4398) <= a or b;
    layer0_outputs(4399) <= not a or b;
    layer0_outputs(4400) <= not (a and b);
    layer0_outputs(4401) <= a or b;
    layer0_outputs(4402) <= a and not b;
    layer0_outputs(4403) <= a xor b;
    layer0_outputs(4404) <= a or b;
    layer0_outputs(4405) <= not b;
    layer0_outputs(4406) <= not (a or b);
    layer0_outputs(4407) <= not b;
    layer0_outputs(4408) <= a xor b;
    layer0_outputs(4409) <= a;
    layer0_outputs(4410) <= not b;
    layer0_outputs(4411) <= b and not a;
    layer0_outputs(4412) <= not (a or b);
    layer0_outputs(4413) <= a and b;
    layer0_outputs(4414) <= not (a or b);
    layer0_outputs(4415) <= not a;
    layer0_outputs(4416) <= a;
    layer0_outputs(4417) <= b and not a;
    layer0_outputs(4418) <= a;
    layer0_outputs(4419) <= a or b;
    layer0_outputs(4420) <= b;
    layer0_outputs(4421) <= not a;
    layer0_outputs(4422) <= not b;
    layer0_outputs(4423) <= a or b;
    layer0_outputs(4424) <= not b;
    layer0_outputs(4425) <= '1';
    layer0_outputs(4426) <= a and b;
    layer0_outputs(4427) <= a or b;
    layer0_outputs(4428) <= not (a and b);
    layer0_outputs(4429) <= a or b;
    layer0_outputs(4430) <= a or b;
    layer0_outputs(4431) <= not a;
    layer0_outputs(4432) <= b;
    layer0_outputs(4433) <= not b or a;
    layer0_outputs(4434) <= a;
    layer0_outputs(4435) <= '1';
    layer0_outputs(4436) <= not (a and b);
    layer0_outputs(4437) <= b;
    layer0_outputs(4438) <= not a or b;
    layer0_outputs(4439) <= not b;
    layer0_outputs(4440) <= not b;
    layer0_outputs(4441) <= not (a or b);
    layer0_outputs(4442) <= not b or a;
    layer0_outputs(4443) <= not b;
    layer0_outputs(4444) <= a xor b;
    layer0_outputs(4445) <= a or b;
    layer0_outputs(4446) <= not (a xor b);
    layer0_outputs(4447) <= not (a or b);
    layer0_outputs(4448) <= not b or a;
    layer0_outputs(4449) <= a and not b;
    layer0_outputs(4450) <= b and not a;
    layer0_outputs(4451) <= not b;
    layer0_outputs(4452) <= not a;
    layer0_outputs(4453) <= b and not a;
    layer0_outputs(4454) <= a and not b;
    layer0_outputs(4455) <= a or b;
    layer0_outputs(4456) <= a xor b;
    layer0_outputs(4457) <= a or b;
    layer0_outputs(4458) <= a xor b;
    layer0_outputs(4459) <= a xor b;
    layer0_outputs(4460) <= not (a or b);
    layer0_outputs(4461) <= not (a or b);
    layer0_outputs(4462) <= not (a xor b);
    layer0_outputs(4463) <= not (a or b);
    layer0_outputs(4464) <= b and not a;
    layer0_outputs(4465) <= not (a or b);
    layer0_outputs(4466) <= not a;
    layer0_outputs(4467) <= a or b;
    layer0_outputs(4468) <= not (a or b);
    layer0_outputs(4469) <= b;
    layer0_outputs(4470) <= not b;
    layer0_outputs(4471) <= not b or a;
    layer0_outputs(4472) <= a or b;
    layer0_outputs(4473) <= not (a or b);
    layer0_outputs(4474) <= not (a and b);
    layer0_outputs(4475) <= b;
    layer0_outputs(4476) <= not (a or b);
    layer0_outputs(4477) <= not b or a;
    layer0_outputs(4478) <= not (a xor b);
    layer0_outputs(4479) <= not (a or b);
    layer0_outputs(4480) <= not b or a;
    layer0_outputs(4481) <= a and not b;
    layer0_outputs(4482) <= a or b;
    layer0_outputs(4483) <= not a;
    layer0_outputs(4484) <= a;
    layer0_outputs(4485) <= not (a or b);
    layer0_outputs(4486) <= not (a or b);
    layer0_outputs(4487) <= b and not a;
    layer0_outputs(4488) <= not (a or b);
    layer0_outputs(4489) <= a or b;
    layer0_outputs(4490) <= a xor b;
    layer0_outputs(4491) <= b;
    layer0_outputs(4492) <= a;
    layer0_outputs(4493) <= a or b;
    layer0_outputs(4494) <= not (a or b);
    layer0_outputs(4495) <= '1';
    layer0_outputs(4496) <= not (a xor b);
    layer0_outputs(4497) <= not a;
    layer0_outputs(4498) <= a xor b;
    layer0_outputs(4499) <= a or b;
    layer0_outputs(4500) <= a;
    layer0_outputs(4501) <= a xor b;
    layer0_outputs(4502) <= b and not a;
    layer0_outputs(4503) <= not (a xor b);
    layer0_outputs(4504) <= a xor b;
    layer0_outputs(4505) <= not a or b;
    layer0_outputs(4506) <= not a;
    layer0_outputs(4507) <= not (a xor b);
    layer0_outputs(4508) <= b;
    layer0_outputs(4509) <= a or b;
    layer0_outputs(4510) <= a and not b;
    layer0_outputs(4511) <= a xor b;
    layer0_outputs(4512) <= b;
    layer0_outputs(4513) <= not b or a;
    layer0_outputs(4514) <= '0';
    layer0_outputs(4515) <= '1';
    layer0_outputs(4516) <= a xor b;
    layer0_outputs(4517) <= b and not a;
    layer0_outputs(4518) <= not (a xor b);
    layer0_outputs(4519) <= a;
    layer0_outputs(4520) <= not (a xor b);
    layer0_outputs(4521) <= a or b;
    layer0_outputs(4522) <= not (a or b);
    layer0_outputs(4523) <= not (a xor b);
    layer0_outputs(4524) <= a;
    layer0_outputs(4525) <= not (a or b);
    layer0_outputs(4526) <= '0';
    layer0_outputs(4527) <= not (a or b);
    layer0_outputs(4528) <= a;
    layer0_outputs(4529) <= not (a or b);
    layer0_outputs(4530) <= b and not a;
    layer0_outputs(4531) <= a or b;
    layer0_outputs(4532) <= not (a xor b);
    layer0_outputs(4533) <= a and not b;
    layer0_outputs(4534) <= not (a or b);
    layer0_outputs(4535) <= not b;
    layer0_outputs(4536) <= a or b;
    layer0_outputs(4537) <= a xor b;
    layer0_outputs(4538) <= not a;
    layer0_outputs(4539) <= not (a or b);
    layer0_outputs(4540) <= a;
    layer0_outputs(4541) <= a xor b;
    layer0_outputs(4542) <= not a;
    layer0_outputs(4543) <= a or b;
    layer0_outputs(4544) <= not (a xor b);
    layer0_outputs(4545) <= b and not a;
    layer0_outputs(4546) <= b and not a;
    layer0_outputs(4547) <= not b or a;
    layer0_outputs(4548) <= not (a or b);
    layer0_outputs(4549) <= a or b;
    layer0_outputs(4550) <= not (a or b);
    layer0_outputs(4551) <= b and not a;
    layer0_outputs(4552) <= not (a or b);
    layer0_outputs(4553) <= not (a xor b);
    layer0_outputs(4554) <= not (a and b);
    layer0_outputs(4555) <= not b;
    layer0_outputs(4556) <= a or b;
    layer0_outputs(4557) <= a;
    layer0_outputs(4558) <= not b;
    layer0_outputs(4559) <= not (a xor b);
    layer0_outputs(4560) <= b;
    layer0_outputs(4561) <= a or b;
    layer0_outputs(4562) <= a or b;
    layer0_outputs(4563) <= a and not b;
    layer0_outputs(4564) <= not b or a;
    layer0_outputs(4565) <= not b;
    layer0_outputs(4566) <= a;
    layer0_outputs(4567) <= not (a xor b);
    layer0_outputs(4568) <= a or b;
    layer0_outputs(4569) <= b;
    layer0_outputs(4570) <= a or b;
    layer0_outputs(4571) <= not (a or b);
    layer0_outputs(4572) <= a and not b;
    layer0_outputs(4573) <= not a;
    layer0_outputs(4574) <= not b;
    layer0_outputs(4575) <= a and b;
    layer0_outputs(4576) <= a;
    layer0_outputs(4577) <= b;
    layer0_outputs(4578) <= not b or a;
    layer0_outputs(4579) <= b and not a;
    layer0_outputs(4580) <= not (a or b);
    layer0_outputs(4581) <= not (a or b);
    layer0_outputs(4582) <= not (a or b);
    layer0_outputs(4583) <= a or b;
    layer0_outputs(4584) <= b and not a;
    layer0_outputs(4585) <= a;
    layer0_outputs(4586) <= not (a xor b);
    layer0_outputs(4587) <= not b or a;
    layer0_outputs(4588) <= a or b;
    layer0_outputs(4589) <= not a or b;
    layer0_outputs(4590) <= a;
    layer0_outputs(4591) <= not b or a;
    layer0_outputs(4592) <= not (a and b);
    layer0_outputs(4593) <= a xor b;
    layer0_outputs(4594) <= a xor b;
    layer0_outputs(4595) <= not (a or b);
    layer0_outputs(4596) <= not a or b;
    layer0_outputs(4597) <= not a or b;
    layer0_outputs(4598) <= not (a xor b);
    layer0_outputs(4599) <= not (a or b);
    layer0_outputs(4600) <= not a or b;
    layer0_outputs(4601) <= a and not b;
    layer0_outputs(4602) <= not b or a;
    layer0_outputs(4603) <= not a or b;
    layer0_outputs(4604) <= a xor b;
    layer0_outputs(4605) <= b;
    layer0_outputs(4606) <= not b;
    layer0_outputs(4607) <= not (a xor b);
    layer0_outputs(4608) <= not b;
    layer0_outputs(4609) <= not a;
    layer0_outputs(4610) <= '0';
    layer0_outputs(4611) <= a xor b;
    layer0_outputs(4612) <= b and not a;
    layer0_outputs(4613) <= not a;
    layer0_outputs(4614) <= a or b;
    layer0_outputs(4615) <= not a;
    layer0_outputs(4616) <= '0';
    layer0_outputs(4617) <= not b;
    layer0_outputs(4618) <= b and not a;
    layer0_outputs(4619) <= a or b;
    layer0_outputs(4620) <= a xor b;
    layer0_outputs(4621) <= not (a or b);
    layer0_outputs(4622) <= a or b;
    layer0_outputs(4623) <= not a;
    layer0_outputs(4624) <= a;
    layer0_outputs(4625) <= a and not b;
    layer0_outputs(4626) <= not (a or b);
    layer0_outputs(4627) <= not a or b;
    layer0_outputs(4628) <= not (a and b);
    layer0_outputs(4629) <= a and b;
    layer0_outputs(4630) <= b and not a;
    layer0_outputs(4631) <= not a or b;
    layer0_outputs(4632) <= b and not a;
    layer0_outputs(4633) <= not b or a;
    layer0_outputs(4634) <= a or b;
    layer0_outputs(4635) <= not b;
    layer0_outputs(4636) <= a and not b;
    layer0_outputs(4637) <= b;
    layer0_outputs(4638) <= '0';
    layer0_outputs(4639) <= '1';
    layer0_outputs(4640) <= not (a and b);
    layer0_outputs(4641) <= not b;
    layer0_outputs(4642) <= a xor b;
    layer0_outputs(4643) <= a and b;
    layer0_outputs(4644) <= not (a xor b);
    layer0_outputs(4645) <= not b;
    layer0_outputs(4646) <= not a or b;
    layer0_outputs(4647) <= not b or a;
    layer0_outputs(4648) <= not (a or b);
    layer0_outputs(4649) <= a and b;
    layer0_outputs(4650) <= not a or b;
    layer0_outputs(4651) <= not a or b;
    layer0_outputs(4652) <= not (a or b);
    layer0_outputs(4653) <= a and not b;
    layer0_outputs(4654) <= not (a or b);
    layer0_outputs(4655) <= a;
    layer0_outputs(4656) <= a and not b;
    layer0_outputs(4657) <= b and not a;
    layer0_outputs(4658) <= a or b;
    layer0_outputs(4659) <= b;
    layer0_outputs(4660) <= a or b;
    layer0_outputs(4661) <= not a;
    layer0_outputs(4662) <= b and not a;
    layer0_outputs(4663) <= a xor b;
    layer0_outputs(4664) <= '1';
    layer0_outputs(4665) <= a or b;
    layer0_outputs(4666) <= a or b;
    layer0_outputs(4667) <= not a or b;
    layer0_outputs(4668) <= not b or a;
    layer0_outputs(4669) <= not (a or b);
    layer0_outputs(4670) <= a;
    layer0_outputs(4671) <= not (a xor b);
    layer0_outputs(4672) <= a xor b;
    layer0_outputs(4673) <= not a or b;
    layer0_outputs(4674) <= not (a or b);
    layer0_outputs(4675) <= b and not a;
    layer0_outputs(4676) <= not b or a;
    layer0_outputs(4677) <= a;
    layer0_outputs(4678) <= not (a xor b);
    layer0_outputs(4679) <= not b;
    layer0_outputs(4680) <= a xor b;
    layer0_outputs(4681) <= not a or b;
    layer0_outputs(4682) <= a or b;
    layer0_outputs(4683) <= not a;
    layer0_outputs(4684) <= not (a or b);
    layer0_outputs(4685) <= a xor b;
    layer0_outputs(4686) <= not a or b;
    layer0_outputs(4687) <= a xor b;
    layer0_outputs(4688) <= '0';
    layer0_outputs(4689) <= not (a or b);
    layer0_outputs(4690) <= a xor b;
    layer0_outputs(4691) <= a or b;
    layer0_outputs(4692) <= not (a or b);
    layer0_outputs(4693) <= not (a xor b);
    layer0_outputs(4694) <= not (a or b);
    layer0_outputs(4695) <= not b or a;
    layer0_outputs(4696) <= a xor b;
    layer0_outputs(4697) <= not b or a;
    layer0_outputs(4698) <= a or b;
    layer0_outputs(4699) <= b;
    layer0_outputs(4700) <= not b;
    layer0_outputs(4701) <= not a;
    layer0_outputs(4702) <= '1';
    layer0_outputs(4703) <= not (a xor b);
    layer0_outputs(4704) <= not a;
    layer0_outputs(4705) <= a or b;
    layer0_outputs(4706) <= not (a xor b);
    layer0_outputs(4707) <= '0';
    layer0_outputs(4708) <= not (a or b);
    layer0_outputs(4709) <= not (a or b);
    layer0_outputs(4710) <= a xor b;
    layer0_outputs(4711) <= a xor b;
    layer0_outputs(4712) <= not b;
    layer0_outputs(4713) <= b and not a;
    layer0_outputs(4714) <= not b;
    layer0_outputs(4715) <= a xor b;
    layer0_outputs(4716) <= a xor b;
    layer0_outputs(4717) <= a or b;
    layer0_outputs(4718) <= not a;
    layer0_outputs(4719) <= not (a or b);
    layer0_outputs(4720) <= b;
    layer0_outputs(4721) <= not b;
    layer0_outputs(4722) <= b and not a;
    layer0_outputs(4723) <= a or b;
    layer0_outputs(4724) <= not (a or b);
    layer0_outputs(4725) <= a;
    layer0_outputs(4726) <= a and not b;
    layer0_outputs(4727) <= not b;
    layer0_outputs(4728) <= not b or a;
    layer0_outputs(4729) <= a or b;
    layer0_outputs(4730) <= a xor b;
    layer0_outputs(4731) <= not (a or b);
    layer0_outputs(4732) <= a or b;
    layer0_outputs(4733) <= b and not a;
    layer0_outputs(4734) <= not a;
    layer0_outputs(4735) <= not a;
    layer0_outputs(4736) <= not (a or b);
    layer0_outputs(4737) <= '1';
    layer0_outputs(4738) <= not (a xor b);
    layer0_outputs(4739) <= a and not b;
    layer0_outputs(4740) <= a or b;
    layer0_outputs(4741) <= a and not b;
    layer0_outputs(4742) <= not (a and b);
    layer0_outputs(4743) <= a or b;
    layer0_outputs(4744) <= not (a and b);
    layer0_outputs(4745) <= a and b;
    layer0_outputs(4746) <= not b;
    layer0_outputs(4747) <= a and not b;
    layer0_outputs(4748) <= not (a or b);
    layer0_outputs(4749) <= not (a or b);
    layer0_outputs(4750) <= a or b;
    layer0_outputs(4751) <= a or b;
    layer0_outputs(4752) <= not b or a;
    layer0_outputs(4753) <= not b;
    layer0_outputs(4754) <= a;
    layer0_outputs(4755) <= not b or a;
    layer0_outputs(4756) <= not (a and b);
    layer0_outputs(4757) <= a or b;
    layer0_outputs(4758) <= not a or b;
    layer0_outputs(4759) <= not (a or b);
    layer0_outputs(4760) <= a or b;
    layer0_outputs(4761) <= not a or b;
    layer0_outputs(4762) <= b;
    layer0_outputs(4763) <= a xor b;
    layer0_outputs(4764) <= not b or a;
    layer0_outputs(4765) <= a or b;
    layer0_outputs(4766) <= '1';
    layer0_outputs(4767) <= a or b;
    layer0_outputs(4768) <= not a or b;
    layer0_outputs(4769) <= '1';
    layer0_outputs(4770) <= not a;
    layer0_outputs(4771) <= a;
    layer0_outputs(4772) <= a or b;
    layer0_outputs(4773) <= a xor b;
    layer0_outputs(4774) <= not (a or b);
    layer0_outputs(4775) <= not (a xor b);
    layer0_outputs(4776) <= a;
    layer0_outputs(4777) <= a or b;
    layer0_outputs(4778) <= not b or a;
    layer0_outputs(4779) <= b and not a;
    layer0_outputs(4780) <= not a or b;
    layer0_outputs(4781) <= not a or b;
    layer0_outputs(4782) <= not (a or b);
    layer0_outputs(4783) <= a;
    layer0_outputs(4784) <= a and not b;
    layer0_outputs(4785) <= a xor b;
    layer0_outputs(4786) <= b;
    layer0_outputs(4787) <= a and not b;
    layer0_outputs(4788) <= a xor b;
    layer0_outputs(4789) <= b and not a;
    layer0_outputs(4790) <= not a;
    layer0_outputs(4791) <= a and not b;
    layer0_outputs(4792) <= not a;
    layer0_outputs(4793) <= a and not b;
    layer0_outputs(4794) <= not (a or b);
    layer0_outputs(4795) <= a or b;
    layer0_outputs(4796) <= not a or b;
    layer0_outputs(4797) <= not (a or b);
    layer0_outputs(4798) <= a;
    layer0_outputs(4799) <= a or b;
    layer0_outputs(4800) <= not (a or b);
    layer0_outputs(4801) <= not a;
    layer0_outputs(4802) <= not a;
    layer0_outputs(4803) <= not b or a;
    layer0_outputs(4804) <= not (a or b);
    layer0_outputs(4805) <= b and not a;
    layer0_outputs(4806) <= b;
    layer0_outputs(4807) <= b and not a;
    layer0_outputs(4808) <= not b;
    layer0_outputs(4809) <= not (a or b);
    layer0_outputs(4810) <= b and not a;
    layer0_outputs(4811) <= a or b;
    layer0_outputs(4812) <= not (a or b);
    layer0_outputs(4813) <= a and b;
    layer0_outputs(4814) <= b and not a;
    layer0_outputs(4815) <= not (a or b);
    layer0_outputs(4816) <= not a or b;
    layer0_outputs(4817) <= a xor b;
    layer0_outputs(4818) <= '0';
    layer0_outputs(4819) <= a or b;
    layer0_outputs(4820) <= not (a xor b);
    layer0_outputs(4821) <= not (a xor b);
    layer0_outputs(4822) <= b and not a;
    layer0_outputs(4823) <= not (a xor b);
    layer0_outputs(4824) <= a or b;
    layer0_outputs(4825) <= a xor b;
    layer0_outputs(4826) <= a and not b;
    layer0_outputs(4827) <= not a;
    layer0_outputs(4828) <= not (a or b);
    layer0_outputs(4829) <= a or b;
    layer0_outputs(4830) <= a and not b;
    layer0_outputs(4831) <= '0';
    layer0_outputs(4832) <= not a or b;
    layer0_outputs(4833) <= not b or a;
    layer0_outputs(4834) <= a or b;
    layer0_outputs(4835) <= not a;
    layer0_outputs(4836) <= not (a xor b);
    layer0_outputs(4837) <= not b or a;
    layer0_outputs(4838) <= b;
    layer0_outputs(4839) <= not a or b;
    layer0_outputs(4840) <= a and not b;
    layer0_outputs(4841) <= b;
    layer0_outputs(4842) <= a and not b;
    layer0_outputs(4843) <= '1';
    layer0_outputs(4844) <= a or b;
    layer0_outputs(4845) <= not a;
    layer0_outputs(4846) <= not (a xor b);
    layer0_outputs(4847) <= b;
    layer0_outputs(4848) <= b;
    layer0_outputs(4849) <= not b or a;
    layer0_outputs(4850) <= not b;
    layer0_outputs(4851) <= not (a or b);
    layer0_outputs(4852) <= a;
    layer0_outputs(4853) <= not (a or b);
    layer0_outputs(4854) <= '0';
    layer0_outputs(4855) <= not (a or b);
    layer0_outputs(4856) <= not b or a;
    layer0_outputs(4857) <= b and not a;
    layer0_outputs(4858) <= b;
    layer0_outputs(4859) <= a and not b;
    layer0_outputs(4860) <= not (a xor b);
    layer0_outputs(4861) <= a;
    layer0_outputs(4862) <= a or b;
    layer0_outputs(4863) <= not b;
    layer0_outputs(4864) <= a;
    layer0_outputs(4865) <= '1';
    layer0_outputs(4866) <= not (a or b);
    layer0_outputs(4867) <= a or b;
    layer0_outputs(4868) <= not (a or b);
    layer0_outputs(4869) <= not (a xor b);
    layer0_outputs(4870) <= b;
    layer0_outputs(4871) <= not (a or b);
    layer0_outputs(4872) <= b and not a;
    layer0_outputs(4873) <= not (a xor b);
    layer0_outputs(4874) <= b and not a;
    layer0_outputs(4875) <= not b or a;
    layer0_outputs(4876) <= a or b;
    layer0_outputs(4877) <= not (a or b);
    layer0_outputs(4878) <= a and not b;
    layer0_outputs(4879) <= a or b;
    layer0_outputs(4880) <= not b;
    layer0_outputs(4881) <= a or b;
    layer0_outputs(4882) <= not (a or b);
    layer0_outputs(4883) <= a or b;
    layer0_outputs(4884) <= not (a or b);
    layer0_outputs(4885) <= not a or b;
    layer0_outputs(4886) <= not (a xor b);
    layer0_outputs(4887) <= not (a or b);
    layer0_outputs(4888) <= not (a and b);
    layer0_outputs(4889) <= not (a xor b);
    layer0_outputs(4890) <= a xor b;
    layer0_outputs(4891) <= b;
    layer0_outputs(4892) <= b and not a;
    layer0_outputs(4893) <= b and not a;
    layer0_outputs(4894) <= b and not a;
    layer0_outputs(4895) <= not b or a;
    layer0_outputs(4896) <= not a or b;
    layer0_outputs(4897) <= not (a or b);
    layer0_outputs(4898) <= not (a or b);
    layer0_outputs(4899) <= not (a xor b);
    layer0_outputs(4900) <= a or b;
    layer0_outputs(4901) <= a;
    layer0_outputs(4902) <= '0';
    layer0_outputs(4903) <= b;
    layer0_outputs(4904) <= a xor b;
    layer0_outputs(4905) <= a and not b;
    layer0_outputs(4906) <= a xor b;
    layer0_outputs(4907) <= not a or b;
    layer0_outputs(4908) <= a xor b;
    layer0_outputs(4909) <= not a or b;
    layer0_outputs(4910) <= not a or b;
    layer0_outputs(4911) <= not (a or b);
    layer0_outputs(4912) <= a or b;
    layer0_outputs(4913) <= a or b;
    layer0_outputs(4914) <= a or b;
    layer0_outputs(4915) <= not b;
    layer0_outputs(4916) <= a xor b;
    layer0_outputs(4917) <= not a;
    layer0_outputs(4918) <= a xor b;
    layer0_outputs(4919) <= a and not b;
    layer0_outputs(4920) <= a or b;
    layer0_outputs(4921) <= not (a or b);
    layer0_outputs(4922) <= not b or a;
    layer0_outputs(4923) <= a;
    layer0_outputs(4924) <= not b;
    layer0_outputs(4925) <= b and not a;
    layer0_outputs(4926) <= b;
    layer0_outputs(4927) <= a and b;
    layer0_outputs(4928) <= a or b;
    layer0_outputs(4929) <= not (a xor b);
    layer0_outputs(4930) <= a or b;
    layer0_outputs(4931) <= a or b;
    layer0_outputs(4932) <= a or b;
    layer0_outputs(4933) <= a;
    layer0_outputs(4934) <= not a;
    layer0_outputs(4935) <= not a or b;
    layer0_outputs(4936) <= a or b;
    layer0_outputs(4937) <= not a;
    layer0_outputs(4938) <= not (a or b);
    layer0_outputs(4939) <= a xor b;
    layer0_outputs(4940) <= not a or b;
    layer0_outputs(4941) <= a;
    layer0_outputs(4942) <= not a or b;
    layer0_outputs(4943) <= a or b;
    layer0_outputs(4944) <= a;
    layer0_outputs(4945) <= a xor b;
    layer0_outputs(4946) <= a xor b;
    layer0_outputs(4947) <= a or b;
    layer0_outputs(4948) <= a or b;
    layer0_outputs(4949) <= a and not b;
    layer0_outputs(4950) <= a or b;
    layer0_outputs(4951) <= '0';
    layer0_outputs(4952) <= a or b;
    layer0_outputs(4953) <= a or b;
    layer0_outputs(4954) <= not (a or b);
    layer0_outputs(4955) <= b and not a;
    layer0_outputs(4956) <= not (a or b);
    layer0_outputs(4957) <= not a or b;
    layer0_outputs(4958) <= not (a xor b);
    layer0_outputs(4959) <= '1';
    layer0_outputs(4960) <= a or b;
    layer0_outputs(4961) <= a or b;
    layer0_outputs(4962) <= not (a or b);
    layer0_outputs(4963) <= not (a or b);
    layer0_outputs(4964) <= not a;
    layer0_outputs(4965) <= not a or b;
    layer0_outputs(4966) <= not b or a;
    layer0_outputs(4967) <= b;
    layer0_outputs(4968) <= a or b;
    layer0_outputs(4969) <= not a or b;
    layer0_outputs(4970) <= b and not a;
    layer0_outputs(4971) <= not b;
    layer0_outputs(4972) <= not (a or b);
    layer0_outputs(4973) <= a or b;
    layer0_outputs(4974) <= not (a and b);
    layer0_outputs(4975) <= not (a or b);
    layer0_outputs(4976) <= a and not b;
    layer0_outputs(4977) <= b;
    layer0_outputs(4978) <= not (a xor b);
    layer0_outputs(4979) <= a and not b;
    layer0_outputs(4980) <= a xor b;
    layer0_outputs(4981) <= not b;
    layer0_outputs(4982) <= not (a or b);
    layer0_outputs(4983) <= '0';
    layer0_outputs(4984) <= not (a and b);
    layer0_outputs(4985) <= b;
    layer0_outputs(4986) <= a or b;
    layer0_outputs(4987) <= not (a and b);
    layer0_outputs(4988) <= b and not a;
    layer0_outputs(4989) <= a xor b;
    layer0_outputs(4990) <= a;
    layer0_outputs(4991) <= not (a or b);
    layer0_outputs(4992) <= not a or b;
    layer0_outputs(4993) <= not b;
    layer0_outputs(4994) <= not (a or b);
    layer0_outputs(4995) <= not (a or b);
    layer0_outputs(4996) <= not (a or b);
    layer0_outputs(4997) <= a or b;
    layer0_outputs(4998) <= not (a xor b);
    layer0_outputs(4999) <= a or b;
    layer0_outputs(5000) <= not b;
    layer0_outputs(5001) <= a or b;
    layer0_outputs(5002) <= a and not b;
    layer0_outputs(5003) <= not a or b;
    layer0_outputs(5004) <= not (a or b);
    layer0_outputs(5005) <= b and not a;
    layer0_outputs(5006) <= not (a and b);
    layer0_outputs(5007) <= not (a xor b);
    layer0_outputs(5008) <= not (a or b);
    layer0_outputs(5009) <= not a or b;
    layer0_outputs(5010) <= not a or b;
    layer0_outputs(5011) <= not a;
    layer0_outputs(5012) <= a;
    layer0_outputs(5013) <= a or b;
    layer0_outputs(5014) <= a and not b;
    layer0_outputs(5015) <= not b;
    layer0_outputs(5016) <= not a;
    layer0_outputs(5017) <= not (a or b);
    layer0_outputs(5018) <= not b or a;
    layer0_outputs(5019) <= not b;
    layer0_outputs(5020) <= a xor b;
    layer0_outputs(5021) <= not (a or b);
    layer0_outputs(5022) <= b and not a;
    layer0_outputs(5023) <= not (a or b);
    layer0_outputs(5024) <= not a;
    layer0_outputs(5025) <= not b or a;
    layer0_outputs(5026) <= not (a or b);
    layer0_outputs(5027) <= not (a or b);
    layer0_outputs(5028) <= a xor b;
    layer0_outputs(5029) <= a or b;
    layer0_outputs(5030) <= a or b;
    layer0_outputs(5031) <= not (a or b);
    layer0_outputs(5032) <= not a or b;
    layer0_outputs(5033) <= not (a or b);
    layer0_outputs(5034) <= not (a and b);
    layer0_outputs(5035) <= not b;
    layer0_outputs(5036) <= a or b;
    layer0_outputs(5037) <= not (a or b);
    layer0_outputs(5038) <= a xor b;
    layer0_outputs(5039) <= not b or a;
    layer0_outputs(5040) <= b;
    layer0_outputs(5041) <= not (a and b);
    layer0_outputs(5042) <= not b;
    layer0_outputs(5043) <= b and not a;
    layer0_outputs(5044) <= a and not b;
    layer0_outputs(5045) <= a;
    layer0_outputs(5046) <= a;
    layer0_outputs(5047) <= not b;
    layer0_outputs(5048) <= not (a xor b);
    layer0_outputs(5049) <= not (a and b);
    layer0_outputs(5050) <= b;
    layer0_outputs(5051) <= a xor b;
    layer0_outputs(5052) <= not b or a;
    layer0_outputs(5053) <= not (a xor b);
    layer0_outputs(5054) <= not (a or b);
    layer0_outputs(5055) <= not (a and b);
    layer0_outputs(5056) <= not b;
    layer0_outputs(5057) <= not (a or b);
    layer0_outputs(5058) <= a or b;
    layer0_outputs(5059) <= not (a or b);
    layer0_outputs(5060) <= not a or b;
    layer0_outputs(5061) <= not (a xor b);
    layer0_outputs(5062) <= not (a or b);
    layer0_outputs(5063) <= not (a or b);
    layer0_outputs(5064) <= a or b;
    layer0_outputs(5065) <= not b;
    layer0_outputs(5066) <= '0';
    layer0_outputs(5067) <= not (a xor b);
    layer0_outputs(5068) <= not a or b;
    layer0_outputs(5069) <= not (a or b);
    layer0_outputs(5070) <= a xor b;
    layer0_outputs(5071) <= not (a or b);
    layer0_outputs(5072) <= not (a or b);
    layer0_outputs(5073) <= a or b;
    layer0_outputs(5074) <= '1';
    layer0_outputs(5075) <= not a;
    layer0_outputs(5076) <= not (a and b);
    layer0_outputs(5077) <= a xor b;
    layer0_outputs(5078) <= '1';
    layer0_outputs(5079) <= b;
    layer0_outputs(5080) <= not a;
    layer0_outputs(5081) <= not a or b;
    layer0_outputs(5082) <= not (a xor b);
    layer0_outputs(5083) <= not a;
    layer0_outputs(5084) <= b and not a;
    layer0_outputs(5085) <= b;
    layer0_outputs(5086) <= not (a or b);
    layer0_outputs(5087) <= b and not a;
    layer0_outputs(5088) <= a xor b;
    layer0_outputs(5089) <= '0';
    layer0_outputs(5090) <= a or b;
    layer0_outputs(5091) <= b and not a;
    layer0_outputs(5092) <= b and not a;
    layer0_outputs(5093) <= b and not a;
    layer0_outputs(5094) <= a and not b;
    layer0_outputs(5095) <= b and not a;
    layer0_outputs(5096) <= not b;
    layer0_outputs(5097) <= not (a or b);
    layer0_outputs(5098) <= not (a or b);
    layer0_outputs(5099) <= not a;
    layer0_outputs(5100) <= a and b;
    layer0_outputs(5101) <= not b;
    layer0_outputs(5102) <= not b;
    layer0_outputs(5103) <= a and not b;
    layer0_outputs(5104) <= b and not a;
    layer0_outputs(5105) <= not (a or b);
    layer0_outputs(5106) <= a and not b;
    layer0_outputs(5107) <= a or b;
    layer0_outputs(5108) <= a xor b;
    layer0_outputs(5109) <= not (a or b);
    layer0_outputs(5110) <= a or b;
    layer0_outputs(5111) <= not a;
    layer0_outputs(5112) <= not (a or b);
    layer0_outputs(5113) <= not (a xor b);
    layer0_outputs(5114) <= a or b;
    layer0_outputs(5115) <= not (a xor b);
    layer0_outputs(5116) <= not a;
    layer0_outputs(5117) <= not (a xor b);
    layer0_outputs(5118) <= not b or a;
    layer0_outputs(5119) <= b;
    outputs(0) <= not a;
    outputs(1) <= not (a or b);
    outputs(2) <= b;
    outputs(3) <= not (a xor b);
    outputs(4) <= not b;
    outputs(5) <= not a;
    outputs(6) <= not (a and b);
    outputs(7) <= not (a or b);
    outputs(8) <= not (a and b);
    outputs(9) <= a;
    outputs(10) <= not (a or b);
    outputs(11) <= b;
    outputs(12) <= not (a and b);
    outputs(13) <= not (a and b);
    outputs(14) <= a and not b;
    outputs(15) <= not b or a;
    outputs(16) <= not (a xor b);
    outputs(17) <= not (a or b);
    outputs(18) <= b;
    outputs(19) <= a;
    outputs(20) <= not (a xor b);
    outputs(21) <= b;
    outputs(22) <= not a;
    outputs(23) <= a;
    outputs(24) <= not a;
    outputs(25) <= a xor b;
    outputs(26) <= not a;
    outputs(27) <= a or b;
    outputs(28) <= b;
    outputs(29) <= not (a and b);
    outputs(30) <= not (a or b);
    outputs(31) <= a and b;
    outputs(32) <= not (a xor b);
    outputs(33) <= not (a or b);
    outputs(34) <= not (a xor b);
    outputs(35) <= not b;
    outputs(36) <= b and not a;
    outputs(37) <= a;
    outputs(38) <= b;
    outputs(39) <= b and not a;
    outputs(40) <= not (a xor b);
    outputs(41) <= a;
    outputs(42) <= a xor b;
    outputs(43) <= a xor b;
    outputs(44) <= not (a xor b);
    outputs(45) <= b;
    outputs(46) <= not a;
    outputs(47) <= a xor b;
    outputs(48) <= a xor b;
    outputs(49) <= not (a and b);
    outputs(50) <= not (a or b);
    outputs(51) <= not b or a;
    outputs(52) <= not (a or b);
    outputs(53) <= a and not b;
    outputs(54) <= not (a or b);
    outputs(55) <= not (a and b);
    outputs(56) <= not b or a;
    outputs(57) <= a xor b;
    outputs(58) <= a and b;
    outputs(59) <= not b or a;
    outputs(60) <= a;
    outputs(61) <= b and not a;
    outputs(62) <= b;
    outputs(63) <= a;
    outputs(64) <= b;
    outputs(65) <= not b;
    outputs(66) <= a xor b;
    outputs(67) <= a and not b;
    outputs(68) <= b;
    outputs(69) <= a;
    outputs(70) <= a;
    outputs(71) <= not (a xor b);
    outputs(72) <= a and b;
    outputs(73) <= a and b;
    outputs(74) <= a and b;
    outputs(75) <= a or b;
    outputs(76) <= a and b;
    outputs(77) <= not (a and b);
    outputs(78) <= not (a xor b);
    outputs(79) <= b;
    outputs(80) <= a;
    outputs(81) <= b;
    outputs(82) <= a xor b;
    outputs(83) <= not b or a;
    outputs(84) <= a;
    outputs(85) <= a and not b;
    outputs(86) <= a xor b;
    outputs(87) <= a and not b;
    outputs(88) <= not (a or b);
    outputs(89) <= a;
    outputs(90) <= not b or a;
    outputs(91) <= a;
    outputs(92) <= a and b;
    outputs(93) <= b;
    outputs(94) <= a and not b;
    outputs(95) <= not a;
    outputs(96) <= not (a xor b);
    outputs(97) <= b and not a;
    outputs(98) <= not b or a;
    outputs(99) <= not a or b;
    outputs(100) <= b and not a;
    outputs(101) <= b;
    outputs(102) <= a;
    outputs(103) <= a and not b;
    outputs(104) <= a;
    outputs(105) <= not (a and b);
    outputs(106) <= a;
    outputs(107) <= a;
    outputs(108) <= a and b;
    outputs(109) <= b and not a;
    outputs(110) <= a xor b;
    outputs(111) <= b and not a;
    outputs(112) <= a;
    outputs(113) <= not a or b;
    outputs(114) <= not (a and b);
    outputs(115) <= not (a xor b);
    outputs(116) <= b;
    outputs(117) <= a or b;
    outputs(118) <= not (a xor b);
    outputs(119) <= not b;
    outputs(120) <= a and not b;
    outputs(121) <= a;
    outputs(122) <= b;
    outputs(123) <= not a;
    outputs(124) <= not a;
    outputs(125) <= not b or a;
    outputs(126) <= a;
    outputs(127) <= a and not b;
    outputs(128) <= not b;
    outputs(129) <= b;
    outputs(130) <= a;
    outputs(131) <= not b;
    outputs(132) <= a xor b;
    outputs(133) <= a and not b;
    outputs(134) <= not a or b;
    outputs(135) <= not (a xor b);
    outputs(136) <= b and not a;
    outputs(137) <= b and not a;
    outputs(138) <= b and not a;
    outputs(139) <= a and b;
    outputs(140) <= a and not b;
    outputs(141) <= a;
    outputs(142) <= not (a xor b);
    outputs(143) <= b;
    outputs(144) <= a;
    outputs(145) <= a or b;
    outputs(146) <= a xor b;
    outputs(147) <= not (a xor b);
    outputs(148) <= a;
    outputs(149) <= not b;
    outputs(150) <= a;
    outputs(151) <= not b or a;
    outputs(152) <= not (a or b);
    outputs(153) <= b;
    outputs(154) <= not (a and b);
    outputs(155) <= a;
    outputs(156) <= not (a xor b);
    outputs(157) <= a and b;
    outputs(158) <= not a;
    outputs(159) <= not (a and b);
    outputs(160) <= b;
    outputs(161) <= a and not b;
    outputs(162) <= not (a or b);
    outputs(163) <= b;
    outputs(164) <= a;
    outputs(165) <= not b;
    outputs(166) <= not (a or b);
    outputs(167) <= not (a xor b);
    outputs(168) <= not (a xor b);
    outputs(169) <= b;
    outputs(170) <= a;
    outputs(171) <= a and not b;
    outputs(172) <= a xor b;
    outputs(173) <= not (a and b);
    outputs(174) <= not a;
    outputs(175) <= a;
    outputs(176) <= a and not b;
    outputs(177) <= a;
    outputs(178) <= b;
    outputs(179) <= b;
    outputs(180) <= not b;
    outputs(181) <= b;
    outputs(182) <= a xor b;
    outputs(183) <= b;
    outputs(184) <= not a;
    outputs(185) <= not (a xor b);
    outputs(186) <= a xor b;
    outputs(187) <= b;
    outputs(188) <= b;
    outputs(189) <= a and not b;
    outputs(190) <= b;
    outputs(191) <= not (a and b);
    outputs(192) <= a xor b;
    outputs(193) <= a;
    outputs(194) <= not (a and b);
    outputs(195) <= not (a xor b);
    outputs(196) <= not (a or b);
    outputs(197) <= not b;
    outputs(198) <= b;
    outputs(199) <= not (a or b);
    outputs(200) <= not b;
    outputs(201) <= a xor b;
    outputs(202) <= not b or a;
    outputs(203) <= b;
    outputs(204) <= not a;
    outputs(205) <= not (a or b);
    outputs(206) <= not (a xor b);
    outputs(207) <= a xor b;
    outputs(208) <= a;
    outputs(209) <= b and not a;
    outputs(210) <= not a;
    outputs(211) <= b;
    outputs(212) <= not (a or b);
    outputs(213) <= not a;
    outputs(214) <= b;
    outputs(215) <= a and not b;
    outputs(216) <= a and b;
    outputs(217) <= not b;
    outputs(218) <= not (a xor b);
    outputs(219) <= not (a xor b);
    outputs(220) <= b;
    outputs(221) <= a and b;
    outputs(222) <= a and not b;
    outputs(223) <= b;
    outputs(224) <= a xor b;
    outputs(225) <= a and not b;
    outputs(226) <= a xor b;
    outputs(227) <= not a;
    outputs(228) <= a;
    outputs(229) <= a and b;
    outputs(230) <= a;
    outputs(231) <= not (a or b);
    outputs(232) <= a and b;
    outputs(233) <= not (a xor b);
    outputs(234) <= not (a or b);
    outputs(235) <= a;
    outputs(236) <= not (a xor b);
    outputs(237) <= not (a and b);
    outputs(238) <= a and b;
    outputs(239) <= not a;
    outputs(240) <= not (a xor b);
    outputs(241) <= not b;
    outputs(242) <= not b;
    outputs(243) <= not b;
    outputs(244) <= a xor b;
    outputs(245) <= not b;
    outputs(246) <= not b or a;
    outputs(247) <= not a;
    outputs(248) <= b;
    outputs(249) <= not (a and b);
    outputs(250) <= a or b;
    outputs(251) <= not a;
    outputs(252) <= a;
    outputs(253) <= not b or a;
    outputs(254) <= not (a xor b);
    outputs(255) <= a xor b;
    outputs(256) <= b;
    outputs(257) <= not b;
    outputs(258) <= a xor b;
    outputs(259) <= not (a xor b);
    outputs(260) <= a xor b;
    outputs(261) <= not a;
    outputs(262) <= a or b;
    outputs(263) <= not (a or b);
    outputs(264) <= not (a xor b);
    outputs(265) <= a xor b;
    outputs(266) <= not b;
    outputs(267) <= not a or b;
    outputs(268) <= not a;
    outputs(269) <= a;
    outputs(270) <= not a;
    outputs(271) <= not (a or b);
    outputs(272) <= not (a and b);
    outputs(273) <= a;
    outputs(274) <= a or b;
    outputs(275) <= b;
    outputs(276) <= a;
    outputs(277) <= not b;
    outputs(278) <= not (a or b);
    outputs(279) <= a or b;
    outputs(280) <= a xor b;
    outputs(281) <= not a;
    outputs(282) <= a or b;
    outputs(283) <= not b;
    outputs(284) <= b;
    outputs(285) <= a and b;
    outputs(286) <= b;
    outputs(287) <= not (a xor b);
    outputs(288) <= not (a xor b);
    outputs(289) <= b and not a;
    outputs(290) <= b and not a;
    outputs(291) <= not a;
    outputs(292) <= not b;
    outputs(293) <= a and b;
    outputs(294) <= not (a and b);
    outputs(295) <= not b or a;
    outputs(296) <= a xor b;
    outputs(297) <= a;
    outputs(298) <= a xor b;
    outputs(299) <= not a;
    outputs(300) <= a;
    outputs(301) <= a;
    outputs(302) <= b and not a;
    outputs(303) <= b;
    outputs(304) <= a xor b;
    outputs(305) <= a xor b;
    outputs(306) <= a;
    outputs(307) <= b;
    outputs(308) <= a;
    outputs(309) <= b;
    outputs(310) <= a xor b;
    outputs(311) <= b;
    outputs(312) <= not (a xor b);
    outputs(313) <= a and b;
    outputs(314) <= b;
    outputs(315) <= a xor b;
    outputs(316) <= not (a or b);
    outputs(317) <= not (a or b);
    outputs(318) <= not a;
    outputs(319) <= b;
    outputs(320) <= b;
    outputs(321) <= a xor b;
    outputs(322) <= not (a or b);
    outputs(323) <= b;
    outputs(324) <= a;
    outputs(325) <= a and not b;
    outputs(326) <= b;
    outputs(327) <= not b;
    outputs(328) <= a and b;
    outputs(329) <= a and not b;
    outputs(330) <= not (a xor b);
    outputs(331) <= a or b;
    outputs(332) <= not (a or b);
    outputs(333) <= not a;
    outputs(334) <= not (a xor b);
    outputs(335) <= a;
    outputs(336) <= a;
    outputs(337) <= not b;
    outputs(338) <= not (a or b);
    outputs(339) <= b and not a;
    outputs(340) <= b and not a;
    outputs(341) <= a xor b;
    outputs(342) <= a;
    outputs(343) <= not b;
    outputs(344) <= b and not a;
    outputs(345) <= a;
    outputs(346) <= a and b;
    outputs(347) <= not (a xor b);
    outputs(348) <= a and not b;
    outputs(349) <= b and not a;
    outputs(350) <= not (a xor b);
    outputs(351) <= a or b;
    outputs(352) <= not (a and b);
    outputs(353) <= b;
    outputs(354) <= a xor b;
    outputs(355) <= a xor b;
    outputs(356) <= a xor b;
    outputs(357) <= b;
    outputs(358) <= b;
    outputs(359) <= b and not a;
    outputs(360) <= not (a xor b);
    outputs(361) <= b;
    outputs(362) <= not a;
    outputs(363) <= a and b;
    outputs(364) <= not (a or b);
    outputs(365) <= a xor b;
    outputs(366) <= not (a xor b);
    outputs(367) <= a or b;
    outputs(368) <= a;
    outputs(369) <= not b;
    outputs(370) <= not b;
    outputs(371) <= not (a xor b);
    outputs(372) <= not b or a;
    outputs(373) <= b;
    outputs(374) <= a xor b;
    outputs(375) <= not (a or b);
    outputs(376) <= not b;
    outputs(377) <= b;
    outputs(378) <= not a;
    outputs(379) <= not b;
    outputs(380) <= not b;
    outputs(381) <= a and b;
    outputs(382) <= a and b;
    outputs(383) <= b;
    outputs(384) <= not a or b;
    outputs(385) <= not a;
    outputs(386) <= b;
    outputs(387) <= a xor b;
    outputs(388) <= not a;
    outputs(389) <= b and not a;
    outputs(390) <= not (a xor b);
    outputs(391) <= a and b;
    outputs(392) <= a xor b;
    outputs(393) <= a xor b;
    outputs(394) <= a and not b;
    outputs(395) <= b and not a;
    outputs(396) <= b;
    outputs(397) <= not b;
    outputs(398) <= not a;
    outputs(399) <= a and not b;
    outputs(400) <= not a;
    outputs(401) <= not (a xor b);
    outputs(402) <= not a or b;
    outputs(403) <= b;
    outputs(404) <= b;
    outputs(405) <= b;
    outputs(406) <= not (a or b);
    outputs(407) <= not b;
    outputs(408) <= not (a or b);
    outputs(409) <= a;
    outputs(410) <= b;
    outputs(411) <= not (a or b);
    outputs(412) <= b and not a;
    outputs(413) <= b and not a;
    outputs(414) <= a and b;
    outputs(415) <= not (a or b);
    outputs(416) <= '1';
    outputs(417) <= not a;
    outputs(418) <= not a;
    outputs(419) <= not b;
    outputs(420) <= not a or b;
    outputs(421) <= not (a xor b);
    outputs(422) <= a xor b;
    outputs(423) <= a xor b;
    outputs(424) <= not b;
    outputs(425) <= a xor b;
    outputs(426) <= not b;
    outputs(427) <= a;
    outputs(428) <= not (a xor b);
    outputs(429) <= not a or b;
    outputs(430) <= b;
    outputs(431) <= not (a and b);
    outputs(432) <= not b;
    outputs(433) <= a;
    outputs(434) <= a;
    outputs(435) <= not a or b;
    outputs(436) <= a;
    outputs(437) <= not b;
    outputs(438) <= a xor b;
    outputs(439) <= a xor b;
    outputs(440) <= a xor b;
    outputs(441) <= not b;
    outputs(442) <= b;
    outputs(443) <= not b or a;
    outputs(444) <= b;
    outputs(445) <= not b;
    outputs(446) <= b;
    outputs(447) <= not (a and b);
    outputs(448) <= b;
    outputs(449) <= a or b;
    outputs(450) <= a xor b;
    outputs(451) <= not b;
    outputs(452) <= not b or a;
    outputs(453) <= a and not b;
    outputs(454) <= not a;
    outputs(455) <= not (a xor b);
    outputs(456) <= not (a xor b);
    outputs(457) <= not (a xor b);
    outputs(458) <= b and not a;
    outputs(459) <= b and not a;
    outputs(460) <= a and not b;
    outputs(461) <= not a or b;
    outputs(462) <= a or b;
    outputs(463) <= a;
    outputs(464) <= not b;
    outputs(465) <= a and not b;
    outputs(466) <= not (a or b);
    outputs(467) <= a and not b;
    outputs(468) <= not (a or b);
    outputs(469) <= a or b;
    outputs(470) <= a or b;
    outputs(471) <= a and not b;
    outputs(472) <= a;
    outputs(473) <= a and b;
    outputs(474) <= a;
    outputs(475) <= a or b;
    outputs(476) <= not (a xor b);
    outputs(477) <= not (a or b);
    outputs(478) <= not (a or b);
    outputs(479) <= a and not b;
    outputs(480) <= b;
    outputs(481) <= not (a or b);
    outputs(482) <= not a or b;
    outputs(483) <= not (a and b);
    outputs(484) <= b and not a;
    outputs(485) <= a xor b;
    outputs(486) <= not (a or b);
    outputs(487) <= not a or b;
    outputs(488) <= b;
    outputs(489) <= b;
    outputs(490) <= a and not b;
    outputs(491) <= not (a or b);
    outputs(492) <= not (a and b);
    outputs(493) <= not (a xor b);
    outputs(494) <= b;
    outputs(495) <= not (a xor b);
    outputs(496) <= not (a or b);
    outputs(497) <= not (a xor b);
    outputs(498) <= not b;
    outputs(499) <= not (a and b);
    outputs(500) <= not a;
    outputs(501) <= not a;
    outputs(502) <= not (a xor b);
    outputs(503) <= not (a or b);
    outputs(504) <= b;
    outputs(505) <= not (a or b);
    outputs(506) <= a;
    outputs(507) <= a and not b;
    outputs(508) <= not b;
    outputs(509) <= b;
    outputs(510) <= a and not b;
    outputs(511) <= a;
    outputs(512) <= a and b;
    outputs(513) <= a;
    outputs(514) <= not a;
    outputs(515) <= not a;
    outputs(516) <= a and not b;
    outputs(517) <= b and not a;
    outputs(518) <= a and not b;
    outputs(519) <= a and b;
    outputs(520) <= b and not a;
    outputs(521) <= not (a or b);
    outputs(522) <= b and not a;
    outputs(523) <= b;
    outputs(524) <= a and not b;
    outputs(525) <= a and not b;
    outputs(526) <= a and not b;
    outputs(527) <= not (a or b);
    outputs(528) <= '0';
    outputs(529) <= a;
    outputs(530) <= not b;
    outputs(531) <= a and b;
    outputs(532) <= a and not b;
    outputs(533) <= a and b;
    outputs(534) <= not (a xor b);
    outputs(535) <= not (a or b);
    outputs(536) <= a and not b;
    outputs(537) <= not b;
    outputs(538) <= a xor b;
    outputs(539) <= b and not a;
    outputs(540) <= a and not b;
    outputs(541) <= a;
    outputs(542) <= not (a or b);
    outputs(543) <= a and not b;
    outputs(544) <= b and not a;
    outputs(545) <= a and b;
    outputs(546) <= b and not a;
    outputs(547) <= a xor b;
    outputs(548) <= not a;
    outputs(549) <= not (a or b);
    outputs(550) <= not (a xor b);
    outputs(551) <= not (a or b);
    outputs(552) <= not b;
    outputs(553) <= b;
    outputs(554) <= b;
    outputs(555) <= not a;
    outputs(556) <= not (a xor b);
    outputs(557) <= not a;
    outputs(558) <= b;
    outputs(559) <= a and not b;
    outputs(560) <= not (a xor b);
    outputs(561) <= a and b;
    outputs(562) <= a and not b;
    outputs(563) <= a;
    outputs(564) <= a and not b;
    outputs(565) <= not (a or b);
    outputs(566) <= b and not a;
    outputs(567) <= '0';
    outputs(568) <= not b;
    outputs(569) <= a and not b;
    outputs(570) <= a and b;
    outputs(571) <= a and b;
    outputs(572) <= a and b;
    outputs(573) <= b;
    outputs(574) <= a and not b;
    outputs(575) <= a and b;
    outputs(576) <= not (a or b);
    outputs(577) <= not (a or b);
    outputs(578) <= not (a or b);
    outputs(579) <= a xor b;
    outputs(580) <= a and b;
    outputs(581) <= not (a or b);
    outputs(582) <= '0';
    outputs(583) <= b and not a;
    outputs(584) <= a and b;
    outputs(585) <= b and not a;
    outputs(586) <= b and not a;
    outputs(587) <= not (a or b);
    outputs(588) <= not (a or b);
    outputs(589) <= b and not a;
    outputs(590) <= a and b;
    outputs(591) <= not b;
    outputs(592) <= not (a or b);
    outputs(593) <= a and not b;
    outputs(594) <= a;
    outputs(595) <= b and not a;
    outputs(596) <= b and not a;
    outputs(597) <= not b;
    outputs(598) <= '0';
    outputs(599) <= a xor b;
    outputs(600) <= not a;
    outputs(601) <= not (a or b);
    outputs(602) <= not a;
    outputs(603) <= '0';
    outputs(604) <= not a;
    outputs(605) <= a and b;
    outputs(606) <= a and b;
    outputs(607) <= b and not a;
    outputs(608) <= a and b;
    outputs(609) <= not (a xor b);
    outputs(610) <= b and not a;
    outputs(611) <= not (a or b);
    outputs(612) <= a xor b;
    outputs(613) <= a and b;
    outputs(614) <= a and b;
    outputs(615) <= a;
    outputs(616) <= a and not b;
    outputs(617) <= a;
    outputs(618) <= a and b;
    outputs(619) <= not (a or b);
    outputs(620) <= a and b;
    outputs(621) <= not (a or b);
    outputs(622) <= a and not b;
    outputs(623) <= a and b;
    outputs(624) <= not (a xor b);
    outputs(625) <= a xor b;
    outputs(626) <= not (a or b);
    outputs(627) <= not (a xor b);
    outputs(628) <= a;
    outputs(629) <= a and not b;
    outputs(630) <= a xor b;
    outputs(631) <= not (a or b);
    outputs(632) <= not (a xor b);
    outputs(633) <= not (a or b);
    outputs(634) <= not (a or b);
    outputs(635) <= b and not a;
    outputs(636) <= not (a xor b);
    outputs(637) <= a and not b;
    outputs(638) <= not (a or b);
    outputs(639) <= not (a or b);
    outputs(640) <= a and b;
    outputs(641) <= not (a or b);
    outputs(642) <= not (a or b);
    outputs(643) <= a xor b;
    outputs(644) <= a and b;
    outputs(645) <= a and not b;
    outputs(646) <= a and b;
    outputs(647) <= a and b;
    outputs(648) <= a and not b;
    outputs(649) <= b and not a;
    outputs(650) <= b and not a;
    outputs(651) <= a;
    outputs(652) <= not (a or b);
    outputs(653) <= a and b;
    outputs(654) <= not a;
    outputs(655) <= a;
    outputs(656) <= a and not b;
    outputs(657) <= not a;
    outputs(658) <= not (a or b);
    outputs(659) <= not (a or b);
    outputs(660) <= not b;
    outputs(661) <= b and not a;
    outputs(662) <= a and b;
    outputs(663) <= not b;
    outputs(664) <= a and b;
    outputs(665) <= a and not b;
    outputs(666) <= a and not b;
    outputs(667) <= '0';
    outputs(668) <= b and not a;
    outputs(669) <= a and b;
    outputs(670) <= a and not b;
    outputs(671) <= a and b;
    outputs(672) <= not a;
    outputs(673) <= not b;
    outputs(674) <= b and not a;
    outputs(675) <= not b;
    outputs(676) <= not (a or b);
    outputs(677) <= not (a or b);
    outputs(678) <= b and not a;
    outputs(679) <= a and not b;
    outputs(680) <= not (a or b);
    outputs(681) <= a xor b;
    outputs(682) <= not a or b;
    outputs(683) <= a and b;
    outputs(684) <= not (a or b);
    outputs(685) <= a and b;
    outputs(686) <= a and b;
    outputs(687) <= b;
    outputs(688) <= a and not b;
    outputs(689) <= not (a xor b);
    outputs(690) <= not (a or b);
    outputs(691) <= a;
    outputs(692) <= not (a or b);
    outputs(693) <= '0';
    outputs(694) <= a and not b;
    outputs(695) <= not (a or b);
    outputs(696) <= b and not a;
    outputs(697) <= not b;
    outputs(698) <= b and not a;
    outputs(699) <= not b;
    outputs(700) <= not (a or b);
    outputs(701) <= not (a or b);
    outputs(702) <= not a;
    outputs(703) <= not b;
    outputs(704) <= a and b;
    outputs(705) <= not (a xor b);
    outputs(706) <= a and b;
    outputs(707) <= not (a or b);
    outputs(708) <= not b;
    outputs(709) <= a xor b;
    outputs(710) <= not (a or b);
    outputs(711) <= '0';
    outputs(712) <= b and not a;
    outputs(713) <= not (a or b);
    outputs(714) <= b;
    outputs(715) <= a and b;
    outputs(716) <= not (a xor b);
    outputs(717) <= a and not b;
    outputs(718) <= a;
    outputs(719) <= not (a or b);
    outputs(720) <= b and not a;
    outputs(721) <= b and not a;
    outputs(722) <= b and not a;
    outputs(723) <= not b;
    outputs(724) <= a and not b;
    outputs(725) <= not (a or b);
    outputs(726) <= a and b;
    outputs(727) <= '0';
    outputs(728) <= not b;
    outputs(729) <= not a;
    outputs(730) <= a xor b;
    outputs(731) <= not (a or b);
    outputs(732) <= not a or b;
    outputs(733) <= not (a or b);
    outputs(734) <= not a;
    outputs(735) <= a and not b;
    outputs(736) <= not a;
    outputs(737) <= a xor b;
    outputs(738) <= not b;
    outputs(739) <= a and not b;
    outputs(740) <= a and b;
    outputs(741) <= b and not a;
    outputs(742) <= b and not a;
    outputs(743) <= a xor b;
    outputs(744) <= b and not a;
    outputs(745) <= not a;
    outputs(746) <= a and b;
    outputs(747) <= a and b;
    outputs(748) <= b and not a;
    outputs(749) <= not (a or b);
    outputs(750) <= b and not a;
    outputs(751) <= not b;
    outputs(752) <= a xor b;
    outputs(753) <= a and not b;
    outputs(754) <= a and b;
    outputs(755) <= a;
    outputs(756) <= a and not b;
    outputs(757) <= b and not a;
    outputs(758) <= a;
    outputs(759) <= a;
    outputs(760) <= '0';
    outputs(761) <= not (a or b);
    outputs(762) <= a xor b;
    outputs(763) <= not (a xor b);
    outputs(764) <= b and not a;
    outputs(765) <= not a;
    outputs(766) <= b and not a;
    outputs(767) <= a and b;
    outputs(768) <= not (a or b);
    outputs(769) <= a and not b;
    outputs(770) <= a and not b;
    outputs(771) <= a and b;
    outputs(772) <= b and not a;
    outputs(773) <= not (a xor b);
    outputs(774) <= not (a xor b);
    outputs(775) <= a and not b;
    outputs(776) <= not b;
    outputs(777) <= a xor b;
    outputs(778) <= a and b;
    outputs(779) <= b and not a;
    outputs(780) <= a and b;
    outputs(781) <= not a;
    outputs(782) <= b and not a;
    outputs(783) <= a;
    outputs(784) <= a and b;
    outputs(785) <= a and b;
    outputs(786) <= not b;
    outputs(787) <= not (a or b);
    outputs(788) <= a and b;
    outputs(789) <= not a;
    outputs(790) <= b;
    outputs(791) <= b and not a;
    outputs(792) <= a and b;
    outputs(793) <= not (a or b);
    outputs(794) <= not (a xor b);
    outputs(795) <= b;
    outputs(796) <= not (a or b);
    outputs(797) <= b and not a;
    outputs(798) <= not (a or b);
    outputs(799) <= not a;
    outputs(800) <= a and b;
    outputs(801) <= b and not a;
    outputs(802) <= not a;
    outputs(803) <= '0';
    outputs(804) <= not (a or b);
    outputs(805) <= not a;
    outputs(806) <= not (a or b);
    outputs(807) <= not (a or b);
    outputs(808) <= a and b;
    outputs(809) <= a and b;
    outputs(810) <= '0';
    outputs(811) <= b and not a;
    outputs(812) <= not a;
    outputs(813) <= not (a or b);
    outputs(814) <= b and not a;
    outputs(815) <= not a;
    outputs(816) <= not (a xor b);
    outputs(817) <= a and not b;
    outputs(818) <= not (a xor b);
    outputs(819) <= a and not b;
    outputs(820) <= not (a or b);
    outputs(821) <= not (a and b);
    outputs(822) <= a and b;
    outputs(823) <= a and not b;
    outputs(824) <= not (a or b);
    outputs(825) <= not a;
    outputs(826) <= b and not a;
    outputs(827) <= b;
    outputs(828) <= b and not a;
    outputs(829) <= a and b;
    outputs(830) <= not (a xor b);
    outputs(831) <= b and not a;
    outputs(832) <= a and b;
    outputs(833) <= not (a or b);
    outputs(834) <= a and not b;
    outputs(835) <= not (a xor b);
    outputs(836) <= b;
    outputs(837) <= not b;
    outputs(838) <= a and not b;
    outputs(839) <= not a;
    outputs(840) <= b;
    outputs(841) <= a and not b;
    outputs(842) <= not a;
    outputs(843) <= b and not a;
    outputs(844) <= a xor b;
    outputs(845) <= not a;
    outputs(846) <= a and b;
    outputs(847) <= a and b;
    outputs(848) <= not a or b;
    outputs(849) <= not (a or b);
    outputs(850) <= not (a or b);
    outputs(851) <= a xor b;
    outputs(852) <= b and not a;
    outputs(853) <= b and not a;
    outputs(854) <= not a;
    outputs(855) <= not a;
    outputs(856) <= a and not b;
    outputs(857) <= not a;
    outputs(858) <= b;
    outputs(859) <= not (a xor b);
    outputs(860) <= a and not b;
    outputs(861) <= not a;
    outputs(862) <= not b;
    outputs(863) <= a and not b;
    outputs(864) <= a and b;
    outputs(865) <= b and not a;
    outputs(866) <= not a or b;
    outputs(867) <= a and not b;
    outputs(868) <= b and not a;
    outputs(869) <= not (a or b);
    outputs(870) <= b and not a;
    outputs(871) <= a;
    outputs(872) <= b and not a;
    outputs(873) <= not (a or b);
    outputs(874) <= not (a and b);
    outputs(875) <= a and not b;
    outputs(876) <= a and b;
    outputs(877) <= a and b;
    outputs(878) <= not (a xor b);
    outputs(879) <= not (a xor b);
    outputs(880) <= b;
    outputs(881) <= b and not a;
    outputs(882) <= a and not b;
    outputs(883) <= not (a or b);
    outputs(884) <= a and b;
    outputs(885) <= a and b;
    outputs(886) <= not a;
    outputs(887) <= a and not b;
    outputs(888) <= not (a or b);
    outputs(889) <= b and not a;
    outputs(890) <= not (a xor b);
    outputs(891) <= not (a or b);
    outputs(892) <= a;
    outputs(893) <= a;
    outputs(894) <= not b;
    outputs(895) <= a and not b;
    outputs(896) <= a and not b;
    outputs(897) <= a and not b;
    outputs(898) <= not a;
    outputs(899) <= a and b;
    outputs(900) <= a xor b;
    outputs(901) <= b;
    outputs(902) <= a and not b;
    outputs(903) <= not (a or b);
    outputs(904) <= b and not a;
    outputs(905) <= a and not b;
    outputs(906) <= a and b;
    outputs(907) <= not (a or b);
    outputs(908) <= b and not a;
    outputs(909) <= a or b;
    outputs(910) <= a;
    outputs(911) <= not (a xor b);
    outputs(912) <= b and not a;
    outputs(913) <= a and not b;
    outputs(914) <= b and not a;
    outputs(915) <= a;
    outputs(916) <= b;
    outputs(917) <= b;
    outputs(918) <= a and not b;
    outputs(919) <= a xor b;
    outputs(920) <= b and not a;
    outputs(921) <= b and not a;
    outputs(922) <= b and not a;
    outputs(923) <= '0';
    outputs(924) <= b and not a;
    outputs(925) <= a xor b;
    outputs(926) <= a and not b;
    outputs(927) <= '0';
    outputs(928) <= not b;
    outputs(929) <= a and b;
    outputs(930) <= b;
    outputs(931) <= a and not b;
    outputs(932) <= a and not b;
    outputs(933) <= a and not b;
    outputs(934) <= not (a xor b);
    outputs(935) <= a and b;
    outputs(936) <= not a;
    outputs(937) <= not (a or b);
    outputs(938) <= not (a or b);
    outputs(939) <= not (a or b);
    outputs(940) <= b;
    outputs(941) <= b and not a;
    outputs(942) <= a and not b;
    outputs(943) <= b;
    outputs(944) <= a and b;
    outputs(945) <= not a;
    outputs(946) <= a xor b;
    outputs(947) <= not (a or b);
    outputs(948) <= b and not a;
    outputs(949) <= b and not a;
    outputs(950) <= not a;
    outputs(951) <= a and b;
    outputs(952) <= a and b;
    outputs(953) <= b and not a;
    outputs(954) <= not (a xor b);
    outputs(955) <= a and not b;
    outputs(956) <= b;
    outputs(957) <= a and not b;
    outputs(958) <= not a;
    outputs(959) <= a and b;
    outputs(960) <= b and not a;
    outputs(961) <= b and not a;
    outputs(962) <= b and not a;
    outputs(963) <= not (a xor b);
    outputs(964) <= not a;
    outputs(965) <= not (a xor b);
    outputs(966) <= not (a or b);
    outputs(967) <= a and b;
    outputs(968) <= not (a or b);
    outputs(969) <= b;
    outputs(970) <= not (a or b);
    outputs(971) <= a and not b;
    outputs(972) <= a and b;
    outputs(973) <= not a or b;
    outputs(974) <= not a;
    outputs(975) <= a and b;
    outputs(976) <= not (a or b);
    outputs(977) <= a and b;
    outputs(978) <= not (a or b);
    outputs(979) <= a and b;
    outputs(980) <= b;
    outputs(981) <= not b;
    outputs(982) <= not (a or b);
    outputs(983) <= a;
    outputs(984) <= b;
    outputs(985) <= not b;
    outputs(986) <= not b;
    outputs(987) <= b and not a;
    outputs(988) <= not (a or b);
    outputs(989) <= not b;
    outputs(990) <= a and not b;
    outputs(991) <= not b;
    outputs(992) <= a;
    outputs(993) <= a and not b;
    outputs(994) <= b and not a;
    outputs(995) <= a and not b;
    outputs(996) <= a and b;
    outputs(997) <= a xor b;
    outputs(998) <= not a;
    outputs(999) <= '0';
    outputs(1000) <= not a;
    outputs(1001) <= b and not a;
    outputs(1002) <= b and not a;
    outputs(1003) <= not (a or b);
    outputs(1004) <= not b;
    outputs(1005) <= a;
    outputs(1006) <= not (a xor b);
    outputs(1007) <= '0';
    outputs(1008) <= not (a or b);
    outputs(1009) <= a and not b;
    outputs(1010) <= b and not a;
    outputs(1011) <= a and b;
    outputs(1012) <= not (a or b);
    outputs(1013) <= a xor b;
    outputs(1014) <= a and not b;
    outputs(1015) <= a;
    outputs(1016) <= not (a or b);
    outputs(1017) <= b;
    outputs(1018) <= a and not b;
    outputs(1019) <= a and b;
    outputs(1020) <= a;
    outputs(1021) <= a;
    outputs(1022) <= b and not a;
    outputs(1023) <= a and b;
    outputs(1024) <= a;
    outputs(1025) <= not (a xor b);
    outputs(1026) <= not a;
    outputs(1027) <= a xor b;
    outputs(1028) <= a xor b;
    outputs(1029) <= not b or a;
    outputs(1030) <= not b or a;
    outputs(1031) <= not (a or b);
    outputs(1032) <= not a;
    outputs(1033) <= b and not a;
    outputs(1034) <= a;
    outputs(1035) <= b;
    outputs(1036) <= a or b;
    outputs(1037) <= not a;
    outputs(1038) <= b;
    outputs(1039) <= a or b;
    outputs(1040) <= b;
    outputs(1041) <= a;
    outputs(1042) <= not (a and b);
    outputs(1043) <= a xor b;
    outputs(1044) <= b;
    outputs(1045) <= not (a or b);
    outputs(1046) <= not (a xor b);
    outputs(1047) <= not (a xor b);
    outputs(1048) <= a or b;
    outputs(1049) <= a;
    outputs(1050) <= not b or a;
    outputs(1051) <= b;
    outputs(1052) <= a xor b;
    outputs(1053) <= not (a and b);
    outputs(1054) <= b;
    outputs(1055) <= a or b;
    outputs(1056) <= not (a xor b);
    outputs(1057) <= not (a or b);
    outputs(1058) <= b and not a;
    outputs(1059) <= not (a or b);
    outputs(1060) <= not b;
    outputs(1061) <= not a or b;
    outputs(1062) <= not (a xor b);
    outputs(1063) <= not b;
    outputs(1064) <= a;
    outputs(1065) <= not (a and b);
    outputs(1066) <= a or b;
    outputs(1067) <= b;
    outputs(1068) <= b;
    outputs(1069) <= not b or a;
    outputs(1070) <= b;
    outputs(1071) <= not (a xor b);
    outputs(1072) <= not a or b;
    outputs(1073) <= a or b;
    outputs(1074) <= not a or b;
    outputs(1075) <= not b;
    outputs(1076) <= not a;
    outputs(1077) <= a or b;
    outputs(1078) <= not (a or b);
    outputs(1079) <= not a;
    outputs(1080) <= not a;
    outputs(1081) <= not (a xor b);
    outputs(1082) <= a;
    outputs(1083) <= not a;
    outputs(1084) <= not b or a;
    outputs(1085) <= not (a xor b);
    outputs(1086) <= not b or a;
    outputs(1087) <= b and not a;
    outputs(1088) <= b;
    outputs(1089) <= not a;
    outputs(1090) <= a;
    outputs(1091) <= not b;
    outputs(1092) <= b;
    outputs(1093) <= not b or a;
    outputs(1094) <= not b;
    outputs(1095) <= not b or a;
    outputs(1096) <= b and not a;
    outputs(1097) <= not a or b;
    outputs(1098) <= not (a xor b);
    outputs(1099) <= not a or b;
    outputs(1100) <= b;
    outputs(1101) <= not (a xor b);
    outputs(1102) <= not (a and b);
    outputs(1103) <= a xor b;
    outputs(1104) <= not b;
    outputs(1105) <= b;
    outputs(1106) <= not (a or b);
    outputs(1107) <= not (a xor b);
    outputs(1108) <= not a or b;
    outputs(1109) <= not (a xor b);
    outputs(1110) <= b;
    outputs(1111) <= a and b;
    outputs(1112) <= not (a xor b);
    outputs(1113) <= a xor b;
    outputs(1114) <= not (a or b);
    outputs(1115) <= b;
    outputs(1116) <= not b or a;
    outputs(1117) <= b and not a;
    outputs(1118) <= not (a and b);
    outputs(1119) <= not a;
    outputs(1120) <= not (a or b);
    outputs(1121) <= not b;
    outputs(1122) <= a or b;
    outputs(1123) <= not (a and b);
    outputs(1124) <= not (a or b);
    outputs(1125) <= not (a or b);
    outputs(1126) <= a xor b;
    outputs(1127) <= a or b;
    outputs(1128) <= a or b;
    outputs(1129) <= not b;
    outputs(1130) <= a xor b;
    outputs(1131) <= not b;
    outputs(1132) <= a xor b;
    outputs(1133) <= not (a xor b);
    outputs(1134) <= a xor b;
    outputs(1135) <= not a;
    outputs(1136) <= not (a xor b);
    outputs(1137) <= not b;
    outputs(1138) <= b;
    outputs(1139) <= not (a xor b);
    outputs(1140) <= not b;
    outputs(1141) <= not (a xor b);
    outputs(1142) <= not b;
    outputs(1143) <= a and not b;
    outputs(1144) <= a xor b;
    outputs(1145) <= not (a xor b);
    outputs(1146) <= a;
    outputs(1147) <= a xor b;
    outputs(1148) <= not (a xor b);
    outputs(1149) <= not a;
    outputs(1150) <= not a or b;
    outputs(1151) <= a and b;
    outputs(1152) <= not (a xor b);
    outputs(1153) <= b and not a;
    outputs(1154) <= a xor b;
    outputs(1155) <= not (a and b);
    outputs(1156) <= a and not b;
    outputs(1157) <= a;
    outputs(1158) <= b;
    outputs(1159) <= not b or a;
    outputs(1160) <= a;
    outputs(1161) <= not (a or b);
    outputs(1162) <= a and b;
    outputs(1163) <= not (a and b);
    outputs(1164) <= a;
    outputs(1165) <= a;
    outputs(1166) <= not a;
    outputs(1167) <= not b or a;
    outputs(1168) <= not a;
    outputs(1169) <= a;
    outputs(1170) <= not a;
    outputs(1171) <= not (a and b);
    outputs(1172) <= a and not b;
    outputs(1173) <= not (a xor b);
    outputs(1174) <= not a;
    outputs(1175) <= a and b;
    outputs(1176) <= not b;
    outputs(1177) <= not (a or b);
    outputs(1178) <= not b or a;
    outputs(1179) <= '1';
    outputs(1180) <= not b;
    outputs(1181) <= not b;
    outputs(1182) <= a and not b;
    outputs(1183) <= b and not a;
    outputs(1184) <= not (a and b);
    outputs(1185) <= a xor b;
    outputs(1186) <= not a;
    outputs(1187) <= a and b;
    outputs(1188) <= not (a xor b);
    outputs(1189) <= not b;
    outputs(1190) <= not b;
    outputs(1191) <= not b or a;
    outputs(1192) <= not a;
    outputs(1193) <= b and not a;
    outputs(1194) <= not b or a;
    outputs(1195) <= not (a xor b);
    outputs(1196) <= not b;
    outputs(1197) <= not a or b;
    outputs(1198) <= a xor b;
    outputs(1199) <= not (a xor b);
    outputs(1200) <= not a;
    outputs(1201) <= not b;
    outputs(1202) <= not b;
    outputs(1203) <= not a or b;
    outputs(1204) <= a xor b;
    outputs(1205) <= not a or b;
    outputs(1206) <= b;
    outputs(1207) <= not b;
    outputs(1208) <= a;
    outputs(1209) <= b and not a;
    outputs(1210) <= not b;
    outputs(1211) <= a and b;
    outputs(1212) <= a xor b;
    outputs(1213) <= a xor b;
    outputs(1214) <= not (a and b);
    outputs(1215) <= not (a and b);
    outputs(1216) <= not b or a;
    outputs(1217) <= a;
    outputs(1218) <= not (a xor b);
    outputs(1219) <= not (a or b);
    outputs(1220) <= b;
    outputs(1221) <= a and b;
    outputs(1222) <= a and b;
    outputs(1223) <= not a or b;
    outputs(1224) <= a and not b;
    outputs(1225) <= a and not b;
    outputs(1226) <= not (a or b);
    outputs(1227) <= not a;
    outputs(1228) <= not a or b;
    outputs(1229) <= a and b;
    outputs(1230) <= a xor b;
    outputs(1231) <= not b or a;
    outputs(1232) <= a or b;
    outputs(1233) <= b;
    outputs(1234) <= a;
    outputs(1235) <= not a or b;
    outputs(1236) <= not b or a;
    outputs(1237) <= not a;
    outputs(1238) <= a xor b;
    outputs(1239) <= a xor b;
    outputs(1240) <= not (a xor b);
    outputs(1241) <= not a or b;
    outputs(1242) <= not a;
    outputs(1243) <= a;
    outputs(1244) <= a;
    outputs(1245) <= a xor b;
    outputs(1246) <= a;
    outputs(1247) <= a or b;
    outputs(1248) <= a or b;
    outputs(1249) <= a;
    outputs(1250) <= not b or a;
    outputs(1251) <= b;
    outputs(1252) <= a and b;
    outputs(1253) <= a and b;
    outputs(1254) <= a;
    outputs(1255) <= a;
    outputs(1256) <= not (a and b);
    outputs(1257) <= b and not a;
    outputs(1258) <= b;
    outputs(1259) <= not (a xor b);
    outputs(1260) <= not a;
    outputs(1261) <= not b or a;
    outputs(1262) <= not (a and b);
    outputs(1263) <= b and not a;
    outputs(1264) <= not b or a;
    outputs(1265) <= b and not a;
    outputs(1266) <= a xor b;
    outputs(1267) <= not a;
    outputs(1268) <= not a;
    outputs(1269) <= not a or b;
    outputs(1270) <= not b or a;
    outputs(1271) <= not b;
    outputs(1272) <= not (a or b);
    outputs(1273) <= b;
    outputs(1274) <= b and not a;
    outputs(1275) <= a;
    outputs(1276) <= not (a xor b);
    outputs(1277) <= not (a and b);
    outputs(1278) <= not a or b;
    outputs(1279) <= a;
    outputs(1280) <= b and not a;
    outputs(1281) <= not (a and b);
    outputs(1282) <= a and not b;
    outputs(1283) <= b and not a;
    outputs(1284) <= not a or b;
    outputs(1285) <= a;
    outputs(1286) <= not a;
    outputs(1287) <= not b or a;
    outputs(1288) <= a and not b;
    outputs(1289) <= not (a xor b);
    outputs(1290) <= not (a and b);
    outputs(1291) <= '1';
    outputs(1292) <= not a or b;
    outputs(1293) <= a xor b;
    outputs(1294) <= not (a xor b);
    outputs(1295) <= a and not b;
    outputs(1296) <= not (a xor b);
    outputs(1297) <= not a;
    outputs(1298) <= not b;
    outputs(1299) <= a and not b;
    outputs(1300) <= not (a or b);
    outputs(1301) <= a and b;
    outputs(1302) <= a xor b;
    outputs(1303) <= b;
    outputs(1304) <= not b;
    outputs(1305) <= not (a or b);
    outputs(1306) <= a or b;
    outputs(1307) <= b;
    outputs(1308) <= b and not a;
    outputs(1309) <= a;
    outputs(1310) <= a and not b;
    outputs(1311) <= a;
    outputs(1312) <= not (a and b);
    outputs(1313) <= a and not b;
    outputs(1314) <= not (a and b);
    outputs(1315) <= a and b;
    outputs(1316) <= not b or a;
    outputs(1317) <= not a or b;
    outputs(1318) <= a or b;
    outputs(1319) <= not a;
    outputs(1320) <= a;
    outputs(1321) <= a xor b;
    outputs(1322) <= a xor b;
    outputs(1323) <= not b or a;
    outputs(1324) <= not b or a;
    outputs(1325) <= not a or b;
    outputs(1326) <= a and not b;
    outputs(1327) <= not (a and b);
    outputs(1328) <= a;
    outputs(1329) <= not (a and b);
    outputs(1330) <= not b;
    outputs(1331) <= a or b;
    outputs(1332) <= not (a and b);
    outputs(1333) <= a and not b;
    outputs(1334) <= b;
    outputs(1335) <= b;
    outputs(1336) <= not (a or b);
    outputs(1337) <= not (a xor b);
    outputs(1338) <= b and not a;
    outputs(1339) <= not a;
    outputs(1340) <= a xor b;
    outputs(1341) <= a;
    outputs(1342) <= not a;
    outputs(1343) <= not b;
    outputs(1344) <= not (a or b);
    outputs(1345) <= not (a xor b);
    outputs(1346) <= a xor b;
    outputs(1347) <= not a or b;
    outputs(1348) <= not a or b;
    outputs(1349) <= not b or a;
    outputs(1350) <= a xor b;
    outputs(1351) <= not (a xor b);
    outputs(1352) <= a;
    outputs(1353) <= a xor b;
    outputs(1354) <= a or b;
    outputs(1355) <= not b or a;
    outputs(1356) <= not b;
    outputs(1357) <= b;
    outputs(1358) <= not (a or b);
    outputs(1359) <= b and not a;
    outputs(1360) <= not (a and b);
    outputs(1361) <= a or b;
    outputs(1362) <= a;
    outputs(1363) <= not a;
    outputs(1364) <= not b or a;
    outputs(1365) <= a or b;
    outputs(1366) <= not (a xor b);
    outputs(1367) <= b and not a;
    outputs(1368) <= not (a or b);
    outputs(1369) <= b and not a;
    outputs(1370) <= a or b;
    outputs(1371) <= not b or a;
    outputs(1372) <= a and b;
    outputs(1373) <= b;
    outputs(1374) <= not a;
    outputs(1375) <= b;
    outputs(1376) <= not (a xor b);
    outputs(1377) <= not (a and b);
    outputs(1378) <= a;
    outputs(1379) <= a and not b;
    outputs(1380) <= not (a xor b);
    outputs(1381) <= b and not a;
    outputs(1382) <= not b or a;
    outputs(1383) <= a xor b;
    outputs(1384) <= a;
    outputs(1385) <= b and not a;
    outputs(1386) <= not a;
    outputs(1387) <= not a;
    outputs(1388) <= a xor b;
    outputs(1389) <= a;
    outputs(1390) <= not (a xor b);
    outputs(1391) <= not a;
    outputs(1392) <= a;
    outputs(1393) <= b;
    outputs(1394) <= not b;
    outputs(1395) <= not (a or b);
    outputs(1396) <= not b or a;
    outputs(1397) <= a xor b;
    outputs(1398) <= a;
    outputs(1399) <= not b or a;
    outputs(1400) <= a and b;
    outputs(1401) <= not (a xor b);
    outputs(1402) <= b;
    outputs(1403) <= not (a or b);
    outputs(1404) <= not b;
    outputs(1405) <= not a or b;
    outputs(1406) <= not a;
    outputs(1407) <= b;
    outputs(1408) <= not (a xor b);
    outputs(1409) <= not a;
    outputs(1410) <= not (a xor b);
    outputs(1411) <= a and b;
    outputs(1412) <= a and not b;
    outputs(1413) <= not a;
    outputs(1414) <= b;
    outputs(1415) <= b;
    outputs(1416) <= a xor b;
    outputs(1417) <= a xor b;
    outputs(1418) <= not b or a;
    outputs(1419) <= a and not b;
    outputs(1420) <= not (a and b);
    outputs(1421) <= b;
    outputs(1422) <= not a or b;
    outputs(1423) <= a;
    outputs(1424) <= not (a xor b);
    outputs(1425) <= not b;
    outputs(1426) <= not (a and b);
    outputs(1427) <= a;
    outputs(1428) <= a;
    outputs(1429) <= not (a and b);
    outputs(1430) <= not b;
    outputs(1431) <= a;
    outputs(1432) <= a xor b;
    outputs(1433) <= not (a xor b);
    outputs(1434) <= not (a and b);
    outputs(1435) <= a xor b;
    outputs(1436) <= a xor b;
    outputs(1437) <= not a;
    outputs(1438) <= not a;
    outputs(1439) <= not (a xor b);
    outputs(1440) <= not (a and b);
    outputs(1441) <= a;
    outputs(1442) <= not (a and b);
    outputs(1443) <= a or b;
    outputs(1444) <= b;
    outputs(1445) <= not a;
    outputs(1446) <= not a or b;
    outputs(1447) <= not b;
    outputs(1448) <= not (a xor b);
    outputs(1449) <= not a;
    outputs(1450) <= a;
    outputs(1451) <= not b or a;
    outputs(1452) <= not (a or b);
    outputs(1453) <= not b;
    outputs(1454) <= a and not b;
    outputs(1455) <= not (a xor b);
    outputs(1456) <= not a;
    outputs(1457) <= not a or b;
    outputs(1458) <= a and b;
    outputs(1459) <= not b or a;
    outputs(1460) <= not (a or b);
    outputs(1461) <= not b;
    outputs(1462) <= not b or a;
    outputs(1463) <= a or b;
    outputs(1464) <= b;
    outputs(1465) <= a;
    outputs(1466) <= '1';
    outputs(1467) <= b;
    outputs(1468) <= a and not b;
    outputs(1469) <= a xor b;
    outputs(1470) <= b;
    outputs(1471) <= a;
    outputs(1472) <= b;
    outputs(1473) <= a and not b;
    outputs(1474) <= a and not b;
    outputs(1475) <= a and not b;
    outputs(1476) <= not b;
    outputs(1477) <= not a;
    outputs(1478) <= a and b;
    outputs(1479) <= not (a xor b);
    outputs(1480) <= not b;
    outputs(1481) <= not b;
    outputs(1482) <= not b or a;
    outputs(1483) <= a;
    outputs(1484) <= b;
    outputs(1485) <= a or b;
    outputs(1486) <= not a;
    outputs(1487) <= a and not b;
    outputs(1488) <= not (a and b);
    outputs(1489) <= not b;
    outputs(1490) <= a and b;
    outputs(1491) <= a and not b;
    outputs(1492) <= not b;
    outputs(1493) <= not (a or b);
    outputs(1494) <= a;
    outputs(1495) <= not (a or b);
    outputs(1496) <= a;
    outputs(1497) <= a and not b;
    outputs(1498) <= not (a or b);
    outputs(1499) <= a and not b;
    outputs(1500) <= a and b;
    outputs(1501) <= a xor b;
    outputs(1502) <= not (a or b);
    outputs(1503) <= not b;
    outputs(1504) <= b and not a;
    outputs(1505) <= b and not a;
    outputs(1506) <= a;
    outputs(1507) <= a and b;
    outputs(1508) <= not a or b;
    outputs(1509) <= not b;
    outputs(1510) <= a or b;
    outputs(1511) <= not b;
    outputs(1512) <= not (a or b);
    outputs(1513) <= a;
    outputs(1514) <= a xor b;
    outputs(1515) <= not (a xor b);
    outputs(1516) <= a and b;
    outputs(1517) <= not b;
    outputs(1518) <= not a;
    outputs(1519) <= not a;
    outputs(1520) <= a xor b;
    outputs(1521) <= not (a xor b);
    outputs(1522) <= a or b;
    outputs(1523) <= not b or a;
    outputs(1524) <= not a;
    outputs(1525) <= b and not a;
    outputs(1526) <= not a or b;
    outputs(1527) <= not b;
    outputs(1528) <= b and not a;
    outputs(1529) <= a xor b;
    outputs(1530) <= a and b;
    outputs(1531) <= a;
    outputs(1532) <= not b;
    outputs(1533) <= not a;
    outputs(1534) <= a;
    outputs(1535) <= not b;
    outputs(1536) <= a;
    outputs(1537) <= a;
    outputs(1538) <= not b;
    outputs(1539) <= not (a or b);
    outputs(1540) <= b and not a;
    outputs(1541) <= not (a or b);
    outputs(1542) <= not b;
    outputs(1543) <= a or b;
    outputs(1544) <= b;
    outputs(1545) <= a or b;
    outputs(1546) <= a;
    outputs(1547) <= not b;
    outputs(1548) <= not (a xor b);
    outputs(1549) <= not (a xor b);
    outputs(1550) <= b;
    outputs(1551) <= not b;
    outputs(1552) <= not b;
    outputs(1553) <= a and not b;
    outputs(1554) <= a and not b;
    outputs(1555) <= b and not a;
    outputs(1556) <= not (a or b);
    outputs(1557) <= a and not b;
    outputs(1558) <= a xor b;
    outputs(1559) <= a and b;
    outputs(1560) <= not a;
    outputs(1561) <= a xor b;
    outputs(1562) <= not a;
    outputs(1563) <= not a;
    outputs(1564) <= not b;
    outputs(1565) <= not b or a;
    outputs(1566) <= b and not a;
    outputs(1567) <= a;
    outputs(1568) <= not (a or b);
    outputs(1569) <= not a;
    outputs(1570) <= a and not b;
    outputs(1571) <= not (a or b);
    outputs(1572) <= not (a or b);
    outputs(1573) <= b;
    outputs(1574) <= not (a and b);
    outputs(1575) <= not b;
    outputs(1576) <= not a or b;
    outputs(1577) <= a and not b;
    outputs(1578) <= b and not a;
    outputs(1579) <= b and not a;
    outputs(1580) <= b and not a;
    outputs(1581) <= not b;
    outputs(1582) <= not (a xor b);
    outputs(1583) <= b and not a;
    outputs(1584) <= a and not b;
    outputs(1585) <= a and not b;
    outputs(1586) <= not a or b;
    outputs(1587) <= b;
    outputs(1588) <= b;
    outputs(1589) <= not (a xor b);
    outputs(1590) <= not a or b;
    outputs(1591) <= not a;
    outputs(1592) <= b;
    outputs(1593) <= a;
    outputs(1594) <= a and not b;
    outputs(1595) <= not a or b;
    outputs(1596) <= not a;
    outputs(1597) <= not (a or b);
    outputs(1598) <= b;
    outputs(1599) <= not b or a;
    outputs(1600) <= a xor b;
    outputs(1601) <= a and not b;
    outputs(1602) <= a;
    outputs(1603) <= a xor b;
    outputs(1604) <= not a or b;
    outputs(1605) <= not (a xor b);
    outputs(1606) <= not a;
    outputs(1607) <= b and not a;
    outputs(1608) <= a xor b;
    outputs(1609) <= b and not a;
    outputs(1610) <= not b;
    outputs(1611) <= b and not a;
    outputs(1612) <= not a;
    outputs(1613) <= a;
    outputs(1614) <= not a;
    outputs(1615) <= not b;
    outputs(1616) <= a xor b;
    outputs(1617) <= not b or a;
    outputs(1618) <= not (a xor b);
    outputs(1619) <= not (a or b);
    outputs(1620) <= not (a and b);
    outputs(1621) <= b;
    outputs(1622) <= not a or b;
    outputs(1623) <= b and not a;
    outputs(1624) <= not b;
    outputs(1625) <= a xor b;
    outputs(1626) <= not b;
    outputs(1627) <= not (a xor b);
    outputs(1628) <= a;
    outputs(1629) <= not a;
    outputs(1630) <= not (a xor b);
    outputs(1631) <= not (a and b);
    outputs(1632) <= not (a and b);
    outputs(1633) <= not a;
    outputs(1634) <= a xor b;
    outputs(1635) <= not a;
    outputs(1636) <= b and not a;
    outputs(1637) <= not b or a;
    outputs(1638) <= not b;
    outputs(1639) <= b and not a;
    outputs(1640) <= a xor b;
    outputs(1641) <= not (a or b);
    outputs(1642) <= a and not b;
    outputs(1643) <= not a or b;
    outputs(1644) <= b and not a;
    outputs(1645) <= a and not b;
    outputs(1646) <= a and b;
    outputs(1647) <= b and not a;
    outputs(1648) <= not (a xor b);
    outputs(1649) <= a;
    outputs(1650) <= a and not b;
    outputs(1651) <= not a;
    outputs(1652) <= a xor b;
    outputs(1653) <= not a;
    outputs(1654) <= a and b;
    outputs(1655) <= not a;
    outputs(1656) <= a and b;
    outputs(1657) <= a or b;
    outputs(1658) <= b and not a;
    outputs(1659) <= not (a or b);
    outputs(1660) <= b and not a;
    outputs(1661) <= not a;
    outputs(1662) <= a;
    outputs(1663) <= not (a xor b);
    outputs(1664) <= a;
    outputs(1665) <= not (a xor b);
    outputs(1666) <= a and b;
    outputs(1667) <= b;
    outputs(1668) <= a xor b;
    outputs(1669) <= not (a or b);
    outputs(1670) <= b;
    outputs(1671) <= not (a or b);
    outputs(1672) <= not a;
    outputs(1673) <= a or b;
    outputs(1674) <= not b;
    outputs(1675) <= not a or b;
    outputs(1676) <= b;
    outputs(1677) <= a and b;
    outputs(1678) <= b and not a;
    outputs(1679) <= not a;
    outputs(1680) <= a;
    outputs(1681) <= a xor b;
    outputs(1682) <= not (a or b);
    outputs(1683) <= not (a xor b);
    outputs(1684) <= a xor b;
    outputs(1685) <= a and not b;
    outputs(1686) <= a;
    outputs(1687) <= not (a xor b);
    outputs(1688) <= not (a or b);
    outputs(1689) <= b;
    outputs(1690) <= a and b;
    outputs(1691) <= b and not a;
    outputs(1692) <= not a;
    outputs(1693) <= not b or a;
    outputs(1694) <= a and not b;
    outputs(1695) <= not b;
    outputs(1696) <= a xor b;
    outputs(1697) <= not b;
    outputs(1698) <= not a;
    outputs(1699) <= a and b;
    outputs(1700) <= not b;
    outputs(1701) <= a xor b;
    outputs(1702) <= not b;
    outputs(1703) <= a and b;
    outputs(1704) <= not (a or b);
    outputs(1705) <= a and b;
    outputs(1706) <= not (a and b);
    outputs(1707) <= not (a xor b);
    outputs(1708) <= a xor b;
    outputs(1709) <= not (a xor b);
    outputs(1710) <= a or b;
    outputs(1711) <= a and not b;
    outputs(1712) <= b and not a;
    outputs(1713) <= a and not b;
    outputs(1714) <= not (a xor b);
    outputs(1715) <= not a or b;
    outputs(1716) <= not (a xor b);
    outputs(1717) <= b;
    outputs(1718) <= a;
    outputs(1719) <= a;
    outputs(1720) <= a xor b;
    outputs(1721) <= a and b;
    outputs(1722) <= a;
    outputs(1723) <= a;
    outputs(1724) <= not b;
    outputs(1725) <= not a or b;
    outputs(1726) <= b and not a;
    outputs(1727) <= not b;
    outputs(1728) <= not (a xor b);
    outputs(1729) <= a and b;
    outputs(1730) <= a and not b;
    outputs(1731) <= a and b;
    outputs(1732) <= not (a or b);
    outputs(1733) <= not a;
    outputs(1734) <= a xor b;
    outputs(1735) <= a xor b;
    outputs(1736) <= not b or a;
    outputs(1737) <= b and not a;
    outputs(1738) <= not (a and b);
    outputs(1739) <= a xor b;
    outputs(1740) <= not a or b;
    outputs(1741) <= a;
    outputs(1742) <= not (a and b);
    outputs(1743) <= a;
    outputs(1744) <= not b;
    outputs(1745) <= b;
    outputs(1746) <= a xor b;
    outputs(1747) <= a or b;
    outputs(1748) <= not (a xor b);
    outputs(1749) <= not a;
    outputs(1750) <= a xor b;
    outputs(1751) <= b;
    outputs(1752) <= b and not a;
    outputs(1753) <= b;
    outputs(1754) <= a xor b;
    outputs(1755) <= not a or b;
    outputs(1756) <= b;
    outputs(1757) <= a and not b;
    outputs(1758) <= not b;
    outputs(1759) <= not b;
    outputs(1760) <= not (a and b);
    outputs(1761) <= b and not a;
    outputs(1762) <= b;
    outputs(1763) <= a xor b;
    outputs(1764) <= not b or a;
    outputs(1765) <= not (a xor b);
    outputs(1766) <= not b;
    outputs(1767) <= a;
    outputs(1768) <= a and not b;
    outputs(1769) <= not b;
    outputs(1770) <= b;
    outputs(1771) <= not (a xor b);
    outputs(1772) <= a and not b;
    outputs(1773) <= a;
    outputs(1774) <= not (a or b);
    outputs(1775) <= not (a xor b);
    outputs(1776) <= b and not a;
    outputs(1777) <= a and b;
    outputs(1778) <= a and b;
    outputs(1779) <= not b or a;
    outputs(1780) <= not b;
    outputs(1781) <= a xor b;
    outputs(1782) <= a and not b;
    outputs(1783) <= not a or b;
    outputs(1784) <= not a;
    outputs(1785) <= b;
    outputs(1786) <= not b;
    outputs(1787) <= not b;
    outputs(1788) <= a and not b;
    outputs(1789) <= not b;
    outputs(1790) <= not a;
    outputs(1791) <= not b or a;
    outputs(1792) <= b and not a;
    outputs(1793) <= a xor b;
    outputs(1794) <= not a;
    outputs(1795) <= not (a or b);
    outputs(1796) <= a;
    outputs(1797) <= a and not b;
    outputs(1798) <= a and b;
    outputs(1799) <= b;
    outputs(1800) <= not (a and b);
    outputs(1801) <= not b;
    outputs(1802) <= not (a or b);
    outputs(1803) <= a xor b;
    outputs(1804) <= not (a or b);
    outputs(1805) <= b and not a;
    outputs(1806) <= a;
    outputs(1807) <= a and not b;
    outputs(1808) <= not b or a;
    outputs(1809) <= b and not a;
    outputs(1810) <= not (a and b);
    outputs(1811) <= a xor b;
    outputs(1812) <= a;
    outputs(1813) <= not a;
    outputs(1814) <= not a or b;
    outputs(1815) <= not a;
    outputs(1816) <= not b;
    outputs(1817) <= not (a or b);
    outputs(1818) <= not a;
    outputs(1819) <= b;
    outputs(1820) <= not a or b;
    outputs(1821) <= not b;
    outputs(1822) <= not a;
    outputs(1823) <= not b;
    outputs(1824) <= a xor b;
    outputs(1825) <= a;
    outputs(1826) <= not (a or b);
    outputs(1827) <= b;
    outputs(1828) <= b;
    outputs(1829) <= a;
    outputs(1830) <= not a;
    outputs(1831) <= not (a xor b);
    outputs(1832) <= a or b;
    outputs(1833) <= a;
    outputs(1834) <= a xor b;
    outputs(1835) <= not b or a;
    outputs(1836) <= not (a xor b);
    outputs(1837) <= not a;
    outputs(1838) <= not a;
    outputs(1839) <= not a;
    outputs(1840) <= not a;
    outputs(1841) <= not a;
    outputs(1842) <= a;
    outputs(1843) <= b;
    outputs(1844) <= not b;
    outputs(1845) <= a;
    outputs(1846) <= not a;
    outputs(1847) <= a and b;
    outputs(1848) <= not b;
    outputs(1849) <= a xor b;
    outputs(1850) <= a and not b;
    outputs(1851) <= not b;
    outputs(1852) <= not b;
    outputs(1853) <= a xor b;
    outputs(1854) <= not a or b;
    outputs(1855) <= not a or b;
    outputs(1856) <= a;
    outputs(1857) <= not a or b;
    outputs(1858) <= not a;
    outputs(1859) <= not a or b;
    outputs(1860) <= a xor b;
    outputs(1861) <= not (a or b);
    outputs(1862) <= not (a and b);
    outputs(1863) <= not a;
    outputs(1864) <= b and not a;
    outputs(1865) <= a or b;
    outputs(1866) <= b and not a;
    outputs(1867) <= not b;
    outputs(1868) <= a;
    outputs(1869) <= b and not a;
    outputs(1870) <= not (a xor b);
    outputs(1871) <= not (a or b);
    outputs(1872) <= a xor b;
    outputs(1873) <= a xor b;
    outputs(1874) <= b;
    outputs(1875) <= not (a or b);
    outputs(1876) <= b;
    outputs(1877) <= not b or a;
    outputs(1878) <= not (a and b);
    outputs(1879) <= not b;
    outputs(1880) <= not (a or b);
    outputs(1881) <= a and b;
    outputs(1882) <= not b;
    outputs(1883) <= not a or b;
    outputs(1884) <= not b or a;
    outputs(1885) <= not (a and b);
    outputs(1886) <= a xor b;
    outputs(1887) <= not (a xor b);
    outputs(1888) <= not (a xor b);
    outputs(1889) <= not b;
    outputs(1890) <= not b;
    outputs(1891) <= a and b;
    outputs(1892) <= not (a and b);
    outputs(1893) <= b;
    outputs(1894) <= b;
    outputs(1895) <= b;
    outputs(1896) <= b and not a;
    outputs(1897) <= b and not a;
    outputs(1898) <= not (a xor b);
    outputs(1899) <= not b or a;
    outputs(1900) <= b and not a;
    outputs(1901) <= not a;
    outputs(1902) <= a xor b;
    outputs(1903) <= a;
    outputs(1904) <= not a or b;
    outputs(1905) <= b and not a;
    outputs(1906) <= not a;
    outputs(1907) <= a;
    outputs(1908) <= b and not a;
    outputs(1909) <= b;
    outputs(1910) <= not (a or b);
    outputs(1911) <= b;
    outputs(1912) <= a and not b;
    outputs(1913) <= not (a xor b);
    outputs(1914) <= not a;
    outputs(1915) <= a and b;
    outputs(1916) <= b;
    outputs(1917) <= a and b;
    outputs(1918) <= not b or a;
    outputs(1919) <= not a;
    outputs(1920) <= a and not b;
    outputs(1921) <= not a;
    outputs(1922) <= not b or a;
    outputs(1923) <= b and not a;
    outputs(1924) <= a;
    outputs(1925) <= a and not b;
    outputs(1926) <= a and not b;
    outputs(1927) <= a or b;
    outputs(1928) <= not (a xor b);
    outputs(1929) <= b and not a;
    outputs(1930) <= not b;
    outputs(1931) <= not (a and b);
    outputs(1932) <= not b;
    outputs(1933) <= a and not b;
    outputs(1934) <= a xor b;
    outputs(1935) <= not a;
    outputs(1936) <= not b;
    outputs(1937) <= b and not a;
    outputs(1938) <= not (a and b);
    outputs(1939) <= a;
    outputs(1940) <= a;
    outputs(1941) <= a xor b;
    outputs(1942) <= not b;
    outputs(1943) <= not a;
    outputs(1944) <= a xor b;
    outputs(1945) <= not (a or b);
    outputs(1946) <= not a;
    outputs(1947) <= a xor b;
    outputs(1948) <= not b or a;
    outputs(1949) <= a and not b;
    outputs(1950) <= a and b;
    outputs(1951) <= a and not b;
    outputs(1952) <= b and not a;
    outputs(1953) <= not a;
    outputs(1954) <= a xor b;
    outputs(1955) <= a and b;
    outputs(1956) <= not b;
    outputs(1957) <= b and not a;
    outputs(1958) <= a xor b;
    outputs(1959) <= not b;
    outputs(1960) <= not (a or b);
    outputs(1961) <= a and b;
    outputs(1962) <= a and not b;
    outputs(1963) <= a or b;
    outputs(1964) <= a;
    outputs(1965) <= a;
    outputs(1966) <= a;
    outputs(1967) <= a and b;
    outputs(1968) <= not a or b;
    outputs(1969) <= a and b;
    outputs(1970) <= not (a and b);
    outputs(1971) <= a;
    outputs(1972) <= not b;
    outputs(1973) <= not (a or b);
    outputs(1974) <= b;
    outputs(1975) <= not (a or b);
    outputs(1976) <= not (a or b);
    outputs(1977) <= not b or a;
    outputs(1978) <= a xor b;
    outputs(1979) <= not b;
    outputs(1980) <= not (a or b);
    outputs(1981) <= not (a or b);
    outputs(1982) <= not (a or b);
    outputs(1983) <= b;
    outputs(1984) <= not b;
    outputs(1985) <= a;
    outputs(1986) <= b and not a;
    outputs(1987) <= not (a or b);
    outputs(1988) <= not a or b;
    outputs(1989) <= a and not b;
    outputs(1990) <= not b or a;
    outputs(1991) <= not b;
    outputs(1992) <= b and not a;
    outputs(1993) <= not a or b;
    outputs(1994) <= a and not b;
    outputs(1995) <= not (a xor b);
    outputs(1996) <= a xor b;
    outputs(1997) <= not (a xor b);
    outputs(1998) <= b and not a;
    outputs(1999) <= b and not a;
    outputs(2000) <= a;
    outputs(2001) <= not b;
    outputs(2002) <= not a or b;
    outputs(2003) <= a and b;
    outputs(2004) <= not (a and b);
    outputs(2005) <= a;
    outputs(2006) <= a and b;
    outputs(2007) <= a;
    outputs(2008) <= a xor b;
    outputs(2009) <= a and b;
    outputs(2010) <= not a;
    outputs(2011) <= a and b;
    outputs(2012) <= not a or b;
    outputs(2013) <= a xor b;
    outputs(2014) <= not a;
    outputs(2015) <= not (a xor b);
    outputs(2016) <= not a or b;
    outputs(2017) <= a and b;
    outputs(2018) <= b;
    outputs(2019) <= a and not b;
    outputs(2020) <= not a;
    outputs(2021) <= b;
    outputs(2022) <= a or b;
    outputs(2023) <= a;
    outputs(2024) <= b and not a;
    outputs(2025) <= not b;
    outputs(2026) <= not (a and b);
    outputs(2027) <= not b;
    outputs(2028) <= b and not a;
    outputs(2029) <= a and b;
    outputs(2030) <= a xor b;
    outputs(2031) <= not b or a;
    outputs(2032) <= not (a xor b);
    outputs(2033) <= a and b;
    outputs(2034) <= a xor b;
    outputs(2035) <= a xor b;
    outputs(2036) <= b;
    outputs(2037) <= a xor b;
    outputs(2038) <= not (a xor b);
    outputs(2039) <= a;
    outputs(2040) <= a;
    outputs(2041) <= not b or a;
    outputs(2042) <= not (a xor b);
    outputs(2043) <= not (a and b);
    outputs(2044) <= not (a or b);
    outputs(2045) <= a and b;
    outputs(2046) <= not (a or b);
    outputs(2047) <= not (a or b);
    outputs(2048) <= b;
    outputs(2049) <= not a;
    outputs(2050) <= a;
    outputs(2051) <= not (a xor b);
    outputs(2052) <= b and not a;
    outputs(2053) <= b;
    outputs(2054) <= not (a xor b);
    outputs(2055) <= not (a or b);
    outputs(2056) <= b and not a;
    outputs(2057) <= b;
    outputs(2058) <= a;
    outputs(2059) <= a and not b;
    outputs(2060) <= a;
    outputs(2061) <= not (a or b);
    outputs(2062) <= a and b;
    outputs(2063) <= not (a or b);
    outputs(2064) <= b and not a;
    outputs(2065) <= a and not b;
    outputs(2066) <= not (a or b);
    outputs(2067) <= a and b;
    outputs(2068) <= not b;
    outputs(2069) <= not a;
    outputs(2070) <= b and not a;
    outputs(2071) <= a xor b;
    outputs(2072) <= not (a or b);
    outputs(2073) <= b;
    outputs(2074) <= a and not b;
    outputs(2075) <= b and not a;
    outputs(2076) <= b and not a;
    outputs(2077) <= a and not b;
    outputs(2078) <= a;
    outputs(2079) <= not (a xor b);
    outputs(2080) <= a and not b;
    outputs(2081) <= a;
    outputs(2082) <= not a or b;
    outputs(2083) <= a and not b;
    outputs(2084) <= not (a xor b);
    outputs(2085) <= b and not a;
    outputs(2086) <= b;
    outputs(2087) <= not b or a;
    outputs(2088) <= not (a or b);
    outputs(2089) <= a;
    outputs(2090) <= not b;
    outputs(2091) <= not (a or b);
    outputs(2092) <= not a;
    outputs(2093) <= a;
    outputs(2094) <= not b;
    outputs(2095) <= a and b;
    outputs(2096) <= not b;
    outputs(2097) <= not b;
    outputs(2098) <= a xor b;
    outputs(2099) <= b;
    outputs(2100) <= a xor b;
    outputs(2101) <= b;
    outputs(2102) <= not b;
    outputs(2103) <= a and b;
    outputs(2104) <= a and not b;
    outputs(2105) <= b;
    outputs(2106) <= a;
    outputs(2107) <= not (a xor b);
    outputs(2108) <= not (a or b);
    outputs(2109) <= b;
    outputs(2110) <= not (a or b);
    outputs(2111) <= not a;
    outputs(2112) <= not (a or b);
    outputs(2113) <= a;
    outputs(2114) <= not a or b;
    outputs(2115) <= not b or a;
    outputs(2116) <= b and not a;
    outputs(2117) <= not b;
    outputs(2118) <= b;
    outputs(2119) <= a;
    outputs(2120) <= a;
    outputs(2121) <= a xor b;
    outputs(2122) <= not a or b;
    outputs(2123) <= not (a or b);
    outputs(2124) <= not (a xor b);
    outputs(2125) <= b and not a;
    outputs(2126) <= not (a or b);
    outputs(2127) <= a and not b;
    outputs(2128) <= a and b;
    outputs(2129) <= '0';
    outputs(2130) <= b and not a;
    outputs(2131) <= not a;
    outputs(2132) <= not a;
    outputs(2133) <= not a;
    outputs(2134) <= not (a or b);
    outputs(2135) <= b;
    outputs(2136) <= a and b;
    outputs(2137) <= a and b;
    outputs(2138) <= not a or b;
    outputs(2139) <= '0';
    outputs(2140) <= b and not a;
    outputs(2141) <= a;
    outputs(2142) <= a and not b;
    outputs(2143) <= not (a or b);
    outputs(2144) <= b;
    outputs(2145) <= not (a xor b);
    outputs(2146) <= b;
    outputs(2147) <= a;
    outputs(2148) <= b;
    outputs(2149) <= a and not b;
    outputs(2150) <= a and not b;
    outputs(2151) <= a and b;
    outputs(2152) <= not (a xor b);
    outputs(2153) <= b;
    outputs(2154) <= not (a xor b);
    outputs(2155) <= a and not b;
    outputs(2156) <= a;
    outputs(2157) <= not a or b;
    outputs(2158) <= a;
    outputs(2159) <= not (a and b);
    outputs(2160) <= not (a or b);
    outputs(2161) <= a and b;
    outputs(2162) <= b and not a;
    outputs(2163) <= a xor b;
    outputs(2164) <= not b;
    outputs(2165) <= b and not a;
    outputs(2166) <= b and not a;
    outputs(2167) <= not (a or b);
    outputs(2168) <= a and not b;
    outputs(2169) <= a or b;
    outputs(2170) <= not (a xor b);
    outputs(2171) <= not (a or b);
    outputs(2172) <= a and not b;
    outputs(2173) <= a and not b;
    outputs(2174) <= not (a xor b);
    outputs(2175) <= a and b;
    outputs(2176) <= b and not a;
    outputs(2177) <= not a;
    outputs(2178) <= not b;
    outputs(2179) <= b and not a;
    outputs(2180) <= not b;
    outputs(2181) <= a;
    outputs(2182) <= b;
    outputs(2183) <= a xor b;
    outputs(2184) <= b;
    outputs(2185) <= b;
    outputs(2186) <= a;
    outputs(2187) <= not a;
    outputs(2188) <= not a;
    outputs(2189) <= a xor b;
    outputs(2190) <= not (a xor b);
    outputs(2191) <= a;
    outputs(2192) <= a;
    outputs(2193) <= not (a or b);
    outputs(2194) <= not (a or b);
    outputs(2195) <= a xor b;
    outputs(2196) <= not b;
    outputs(2197) <= not (a or b);
    outputs(2198) <= not b;
    outputs(2199) <= a;
    outputs(2200) <= a and b;
    outputs(2201) <= a and not b;
    outputs(2202) <= a;
    outputs(2203) <= not b;
    outputs(2204) <= not (a or b);
    outputs(2205) <= not a;
    outputs(2206) <= a or b;
    outputs(2207) <= a;
    outputs(2208) <= b and not a;
    outputs(2209) <= not a;
    outputs(2210) <= not b;
    outputs(2211) <= not a;
    outputs(2212) <= not (a or b);
    outputs(2213) <= not b;
    outputs(2214) <= b;
    outputs(2215) <= a and not b;
    outputs(2216) <= not a;
    outputs(2217) <= not b;
    outputs(2218) <= not a;
    outputs(2219) <= a and b;
    outputs(2220) <= a xor b;
    outputs(2221) <= b;
    outputs(2222) <= not (a and b);
    outputs(2223) <= b and not a;
    outputs(2224) <= not a;
    outputs(2225) <= b and not a;
    outputs(2226) <= not (a xor b);
    outputs(2227) <= a and b;
    outputs(2228) <= not a;
    outputs(2229) <= a;
    outputs(2230) <= a and b;
    outputs(2231) <= b and not a;
    outputs(2232) <= not (a and b);
    outputs(2233) <= a xor b;
    outputs(2234) <= a and not b;
    outputs(2235) <= a and not b;
    outputs(2236) <= a and not b;
    outputs(2237) <= a xor b;
    outputs(2238) <= not a or b;
    outputs(2239) <= b and not a;
    outputs(2240) <= a xor b;
    outputs(2241) <= not (a or b);
    outputs(2242) <= b and not a;
    outputs(2243) <= not (a and b);
    outputs(2244) <= not b;
    outputs(2245) <= not (a or b);
    outputs(2246) <= not (a xor b);
    outputs(2247) <= b and not a;
    outputs(2248) <= a and b;
    outputs(2249) <= b;
    outputs(2250) <= a xor b;
    outputs(2251) <= a and not b;
    outputs(2252) <= a and not b;
    outputs(2253) <= not (a xor b);
    outputs(2254) <= not (a xor b);
    outputs(2255) <= a xor b;
    outputs(2256) <= not b;
    outputs(2257) <= not (a xor b);
    outputs(2258) <= a and not b;
    outputs(2259) <= b;
    outputs(2260) <= a and b;
    outputs(2261) <= not (a or b);
    outputs(2262) <= not (a or b);
    outputs(2263) <= not (a xor b);
    outputs(2264) <= not b or a;
    outputs(2265) <= not b;
    outputs(2266) <= b and not a;
    outputs(2267) <= a and not b;
    outputs(2268) <= a;
    outputs(2269) <= not (a xor b);
    outputs(2270) <= a xor b;
    outputs(2271) <= b and not a;
    outputs(2272) <= not b;
    outputs(2273) <= a and not b;
    outputs(2274) <= not b;
    outputs(2275) <= b;
    outputs(2276) <= a and not b;
    outputs(2277) <= b and not a;
    outputs(2278) <= not a;
    outputs(2279) <= a and b;
    outputs(2280) <= not a;
    outputs(2281) <= a xor b;
    outputs(2282) <= not (a or b);
    outputs(2283) <= a;
    outputs(2284) <= not a;
    outputs(2285) <= not a;
    outputs(2286) <= b;
    outputs(2287) <= b;
    outputs(2288) <= not (a or b);
    outputs(2289) <= not b;
    outputs(2290) <= not (a or b);
    outputs(2291) <= a xor b;
    outputs(2292) <= b;
    outputs(2293) <= b and not a;
    outputs(2294) <= a and b;
    outputs(2295) <= not (a and b);
    outputs(2296) <= a and b;
    outputs(2297) <= not (a or b);
    outputs(2298) <= b;
    outputs(2299) <= a and b;
    outputs(2300) <= a xor b;
    outputs(2301) <= not b;
    outputs(2302) <= a and not b;
    outputs(2303) <= b;
    outputs(2304) <= not a;
    outputs(2305) <= b and not a;
    outputs(2306) <= not b;
    outputs(2307) <= not (a xor b);
    outputs(2308) <= not a;
    outputs(2309) <= a xor b;
    outputs(2310) <= not (a xor b);
    outputs(2311) <= b;
    outputs(2312) <= a and not b;
    outputs(2313) <= not (a or b);
    outputs(2314) <= a xor b;
    outputs(2315) <= a and b;
    outputs(2316) <= not a;
    outputs(2317) <= a;
    outputs(2318) <= b and not a;
    outputs(2319) <= b and not a;
    outputs(2320) <= not b;
    outputs(2321) <= not a;
    outputs(2322) <= a and not b;
    outputs(2323) <= not (a or b);
    outputs(2324) <= a and not b;
    outputs(2325) <= a and b;
    outputs(2326) <= b and not a;
    outputs(2327) <= not (a xor b);
    outputs(2328) <= not b or a;
    outputs(2329) <= not a;
    outputs(2330) <= not a;
    outputs(2331) <= a or b;
    outputs(2332) <= not a;
    outputs(2333) <= b;
    outputs(2334) <= not b;
    outputs(2335) <= b and not a;
    outputs(2336) <= not b;
    outputs(2337) <= not b;
    outputs(2338) <= a and b;
    outputs(2339) <= a and not b;
    outputs(2340) <= not (a or b);
    outputs(2341) <= a and not b;
    outputs(2342) <= b;
    outputs(2343) <= a and not b;
    outputs(2344) <= a and b;
    outputs(2345) <= a;
    outputs(2346) <= not (a xor b);
    outputs(2347) <= not (a or b);
    outputs(2348) <= b and not a;
    outputs(2349) <= a and b;
    outputs(2350) <= a or b;
    outputs(2351) <= not a;
    outputs(2352) <= a and not b;
    outputs(2353) <= not a;
    outputs(2354) <= a or b;
    outputs(2355) <= b;
    outputs(2356) <= not b;
    outputs(2357) <= not (a or b);
    outputs(2358) <= not (a or b);
    outputs(2359) <= not (a xor b);
    outputs(2360) <= a;
    outputs(2361) <= a xor b;
    outputs(2362) <= a or b;
    outputs(2363) <= b and not a;
    outputs(2364) <= not a;
    outputs(2365) <= not (a or b);
    outputs(2366) <= not (a or b);
    outputs(2367) <= a xor b;
    outputs(2368) <= not b;
    outputs(2369) <= a and b;
    outputs(2370) <= not (a xor b);
    outputs(2371) <= a;
    outputs(2372) <= not (a and b);
    outputs(2373) <= not b;
    outputs(2374) <= a xor b;
    outputs(2375) <= not a;
    outputs(2376) <= b;
    outputs(2377) <= a xor b;
    outputs(2378) <= not (a xor b);
    outputs(2379) <= a and not b;
    outputs(2380) <= not (a or b);
    outputs(2381) <= b;
    outputs(2382) <= a;
    outputs(2383) <= not (a or b);
    outputs(2384) <= not (a or b);
    outputs(2385) <= b and not a;
    outputs(2386) <= a and b;
    outputs(2387) <= not (a or b);
    outputs(2388) <= a;
    outputs(2389) <= b and not a;
    outputs(2390) <= b;
    outputs(2391) <= a and not b;
    outputs(2392) <= b;
    outputs(2393) <= not b;
    outputs(2394) <= a;
    outputs(2395) <= not (a or b);
    outputs(2396) <= not (a xor b);
    outputs(2397) <= b;
    outputs(2398) <= b and not a;
    outputs(2399) <= b;
    outputs(2400) <= a or b;
    outputs(2401) <= a or b;
    outputs(2402) <= a;
    outputs(2403) <= b and not a;
    outputs(2404) <= b and not a;
    outputs(2405) <= b;
    outputs(2406) <= a xor b;
    outputs(2407) <= not (a or b);
    outputs(2408) <= a;
    outputs(2409) <= a and not b;
    outputs(2410) <= not (a or b);
    outputs(2411) <= not (a xor b);
    outputs(2412) <= not b;
    outputs(2413) <= not (a and b);
    outputs(2414) <= a xor b;
    outputs(2415) <= a and b;
    outputs(2416) <= b and not a;
    outputs(2417) <= a xor b;
    outputs(2418) <= not b;
    outputs(2419) <= a;
    outputs(2420) <= not (a or b);
    outputs(2421) <= a;
    outputs(2422) <= a and not b;
    outputs(2423) <= not (a or b);
    outputs(2424) <= a and not b;
    outputs(2425) <= a and b;
    outputs(2426) <= a;
    outputs(2427) <= not b;
    outputs(2428) <= a and b;
    outputs(2429) <= a and not b;
    outputs(2430) <= a and not b;
    outputs(2431) <= a and b;
    outputs(2432) <= not (a or b);
    outputs(2433) <= not (a or b);
    outputs(2434) <= not (a or b);
    outputs(2435) <= not (a xor b);
    outputs(2436) <= a and b;
    outputs(2437) <= a;
    outputs(2438) <= a and b;
    outputs(2439) <= b and not a;
    outputs(2440) <= not (a xor b);
    outputs(2441) <= a and b;
    outputs(2442) <= a and b;
    outputs(2443) <= a and b;
    outputs(2444) <= a xor b;
    outputs(2445) <= a and b;
    outputs(2446) <= not (a or b);
    outputs(2447) <= a;
    outputs(2448) <= b;
    outputs(2449) <= not b;
    outputs(2450) <= a and not b;
    outputs(2451) <= not b;
    outputs(2452) <= a xor b;
    outputs(2453) <= a xor b;
    outputs(2454) <= not (a xor b);
    outputs(2455) <= a xor b;
    outputs(2456) <= not b;
    outputs(2457) <= a;
    outputs(2458) <= b and not a;
    outputs(2459) <= a;
    outputs(2460) <= a and not b;
    outputs(2461) <= a;
    outputs(2462) <= not a;
    outputs(2463) <= not (a or b);
    outputs(2464) <= a xor b;
    outputs(2465) <= not (a or b);
    outputs(2466) <= not b;
    outputs(2467) <= a or b;
    outputs(2468) <= b and not a;
    outputs(2469) <= b;
    outputs(2470) <= not b;
    outputs(2471) <= not (a xor b);
    outputs(2472) <= a;
    outputs(2473) <= b and not a;
    outputs(2474) <= not b or a;
    outputs(2475) <= not (a xor b);
    outputs(2476) <= b and not a;
    outputs(2477) <= a xor b;
    outputs(2478) <= not a or b;
    outputs(2479) <= a and not b;
    outputs(2480) <= b;
    outputs(2481) <= a;
    outputs(2482) <= a;
    outputs(2483) <= not (a xor b);
    outputs(2484) <= not (a xor b);
    outputs(2485) <= b;
    outputs(2486) <= b;
    outputs(2487) <= not (a or b);
    outputs(2488) <= a and not b;
    outputs(2489) <= a and b;
    outputs(2490) <= not a;
    outputs(2491) <= not a;
    outputs(2492) <= not (a xor b);
    outputs(2493) <= a;
    outputs(2494) <= a;
    outputs(2495) <= a;
    outputs(2496) <= a;
    outputs(2497) <= a and b;
    outputs(2498) <= b;
    outputs(2499) <= not a;
    outputs(2500) <= not a;
    outputs(2501) <= not b;
    outputs(2502) <= b and not a;
    outputs(2503) <= a and not b;
    outputs(2504) <= not b;
    outputs(2505) <= a and b;
    outputs(2506) <= not b;
    outputs(2507) <= not b;
    outputs(2508) <= a xor b;
    outputs(2509) <= not (a or b);
    outputs(2510) <= not a;
    outputs(2511) <= b;
    outputs(2512) <= not (a or b);
    outputs(2513) <= not (a xor b);
    outputs(2514) <= a;
    outputs(2515) <= not b;
    outputs(2516) <= a or b;
    outputs(2517) <= not b;
    outputs(2518) <= b and not a;
    outputs(2519) <= not (a or b);
    outputs(2520) <= not (a or b);
    outputs(2521) <= a;
    outputs(2522) <= not a;
    outputs(2523) <= not a;
    outputs(2524) <= not b;
    outputs(2525) <= not a;
    outputs(2526) <= not (a or b);
    outputs(2527) <= not b;
    outputs(2528) <= b and not a;
    outputs(2529) <= a and not b;
    outputs(2530) <= a xor b;
    outputs(2531) <= a xor b;
    outputs(2532) <= a;
    outputs(2533) <= a and not b;
    outputs(2534) <= a or b;
    outputs(2535) <= a;
    outputs(2536) <= b;
    outputs(2537) <= b;
    outputs(2538) <= a xor b;
    outputs(2539) <= not (a or b);
    outputs(2540) <= '0';
    outputs(2541) <= a or b;
    outputs(2542) <= a and b;
    outputs(2543) <= not (a or b);
    outputs(2544) <= b;
    outputs(2545) <= a;
    outputs(2546) <= b;
    outputs(2547) <= not a;
    outputs(2548) <= a and b;
    outputs(2549) <= b;
    outputs(2550) <= not a;
    outputs(2551) <= a;
    outputs(2552) <= not b;
    outputs(2553) <= a and not b;
    outputs(2554) <= a and b;
    outputs(2555) <= not b or a;
    outputs(2556) <= a and not b;
    outputs(2557) <= b and not a;
    outputs(2558) <= not b;
    outputs(2559) <= not (a xor b);
    outputs(2560) <= not (a xor b);
    outputs(2561) <= a xor b;
    outputs(2562) <= a and not b;
    outputs(2563) <= not a;
    outputs(2564) <= not a;
    outputs(2565) <= a;
    outputs(2566) <= not b;
    outputs(2567) <= a and b;
    outputs(2568) <= a and b;
    outputs(2569) <= not a;
    outputs(2570) <= a and b;
    outputs(2571) <= a and b;
    outputs(2572) <= not (a xor b);
    outputs(2573) <= a xor b;
    outputs(2574) <= b;
    outputs(2575) <= not b;
    outputs(2576) <= a xor b;
    outputs(2577) <= a xor b;
    outputs(2578) <= a xor b;
    outputs(2579) <= not a;
    outputs(2580) <= not a;
    outputs(2581) <= not b or a;
    outputs(2582) <= not (a or b);
    outputs(2583) <= not (a and b);
    outputs(2584) <= b and not a;
    outputs(2585) <= not (a xor b);
    outputs(2586) <= not (a xor b);
    outputs(2587) <= a xor b;
    outputs(2588) <= not a;
    outputs(2589) <= not a;
    outputs(2590) <= a xor b;
    outputs(2591) <= not (a xor b);
    outputs(2592) <= b;
    outputs(2593) <= a;
    outputs(2594) <= a and not b;
    outputs(2595) <= a and not b;
    outputs(2596) <= a xor b;
    outputs(2597) <= not (a or b);
    outputs(2598) <= a;
    outputs(2599) <= a xor b;
    outputs(2600) <= a and b;
    outputs(2601) <= not (a xor b);
    outputs(2602) <= a;
    outputs(2603) <= a or b;
    outputs(2604) <= not a;
    outputs(2605) <= not (a xor b);
    outputs(2606) <= not a or b;
    outputs(2607) <= a and b;
    outputs(2608) <= not (a xor b);
    outputs(2609) <= not a;
    outputs(2610) <= b;
    outputs(2611) <= not a;
    outputs(2612) <= not b;
    outputs(2613) <= a or b;
    outputs(2614) <= a and b;
    outputs(2615) <= not (a or b);
    outputs(2616) <= b;
    outputs(2617) <= b;
    outputs(2618) <= not (a xor b);
    outputs(2619) <= b and not a;
    outputs(2620) <= not a;
    outputs(2621) <= a xor b;
    outputs(2622) <= a;
    outputs(2623) <= not b or a;
    outputs(2624) <= a xor b;
    outputs(2625) <= not (a xor b);
    outputs(2626) <= a and not b;
    outputs(2627) <= not (a or b);
    outputs(2628) <= a;
    outputs(2629) <= not (a xor b);
    outputs(2630) <= not a;
    outputs(2631) <= not b;
    outputs(2632) <= b;
    outputs(2633) <= a xor b;
    outputs(2634) <= a xor b;
    outputs(2635) <= not (a xor b);
    outputs(2636) <= a and not b;
    outputs(2637) <= a xor b;
    outputs(2638) <= not b;
    outputs(2639) <= not (a xor b);
    outputs(2640) <= not b;
    outputs(2641) <= not (a xor b);
    outputs(2642) <= not a;
    outputs(2643) <= not (a xor b);
    outputs(2644) <= b;
    outputs(2645) <= not a;
    outputs(2646) <= not a;
    outputs(2647) <= a and b;
    outputs(2648) <= a and b;
    outputs(2649) <= not b;
    outputs(2650) <= not b or a;
    outputs(2651) <= a or b;
    outputs(2652) <= not b;
    outputs(2653) <= not a;
    outputs(2654) <= b;
    outputs(2655) <= b;
    outputs(2656) <= a xor b;
    outputs(2657) <= b and not a;
    outputs(2658) <= not (a or b);
    outputs(2659) <= not (a xor b);
    outputs(2660) <= a and not b;
    outputs(2661) <= not (a and b);
    outputs(2662) <= not (a or b);
    outputs(2663) <= a and b;
    outputs(2664) <= not a;
    outputs(2665) <= a and b;
    outputs(2666) <= not (a xor b);
    outputs(2667) <= not a;
    outputs(2668) <= not a or b;
    outputs(2669) <= b;
    outputs(2670) <= not b or a;
    outputs(2671) <= not a;
    outputs(2672) <= not (a or b);
    outputs(2673) <= not (a xor b);
    outputs(2674) <= not (a xor b);
    outputs(2675) <= a xor b;
    outputs(2676) <= a and not b;
    outputs(2677) <= not (a or b);
    outputs(2678) <= not b or a;
    outputs(2679) <= not a or b;
    outputs(2680) <= b and not a;
    outputs(2681) <= not (a xor b);
    outputs(2682) <= a and not b;
    outputs(2683) <= not b or a;
    outputs(2684) <= a xor b;
    outputs(2685) <= a or b;
    outputs(2686) <= a and not b;
    outputs(2687) <= not (a xor b);
    outputs(2688) <= b and not a;
    outputs(2689) <= not b;
    outputs(2690) <= a xor b;
    outputs(2691) <= a;
    outputs(2692) <= not (a xor b);
    outputs(2693) <= b and not a;
    outputs(2694) <= a and b;
    outputs(2695) <= not b;
    outputs(2696) <= not (a xor b);
    outputs(2697) <= not (a xor b);
    outputs(2698) <= not (a or b);
    outputs(2699) <= not (a xor b);
    outputs(2700) <= not (a xor b);
    outputs(2701) <= a or b;
    outputs(2702) <= a and b;
    outputs(2703) <= not (a xor b);
    outputs(2704) <= not a;
    outputs(2705) <= a;
    outputs(2706) <= a xor b;
    outputs(2707) <= a and b;
    outputs(2708) <= a xor b;
    outputs(2709) <= a or b;
    outputs(2710) <= a;
    outputs(2711) <= a xor b;
    outputs(2712) <= a;
    outputs(2713) <= a and b;
    outputs(2714) <= b;
    outputs(2715) <= b;
    outputs(2716) <= not a or b;
    outputs(2717) <= a and b;
    outputs(2718) <= not a;
    outputs(2719) <= b;
    outputs(2720) <= a;
    outputs(2721) <= not (a or b);
    outputs(2722) <= not (a xor b);
    outputs(2723) <= not (a xor b);
    outputs(2724) <= a;
    outputs(2725) <= a and b;
    outputs(2726) <= not a;
    outputs(2727) <= not a;
    outputs(2728) <= a;
    outputs(2729) <= a and b;
    outputs(2730) <= not b;
    outputs(2731) <= b;
    outputs(2732) <= a xor b;
    outputs(2733) <= b;
    outputs(2734) <= not (a xor b);
    outputs(2735) <= a xor b;
    outputs(2736) <= a and not b;
    outputs(2737) <= not (a xor b);
    outputs(2738) <= not b or a;
    outputs(2739) <= not b;
    outputs(2740) <= b and not a;
    outputs(2741) <= a xor b;
    outputs(2742) <= not (a xor b);
    outputs(2743) <= not b or a;
    outputs(2744) <= a or b;
    outputs(2745) <= a or b;
    outputs(2746) <= not a;
    outputs(2747) <= not (a xor b);
    outputs(2748) <= a xor b;
    outputs(2749) <= not (a and b);
    outputs(2750) <= a;
    outputs(2751) <= b and not a;
    outputs(2752) <= a and b;
    outputs(2753) <= not (a and b);
    outputs(2754) <= not (a or b);
    outputs(2755) <= a and b;
    outputs(2756) <= a xor b;
    outputs(2757) <= b;
    outputs(2758) <= a;
    outputs(2759) <= a xor b;
    outputs(2760) <= a and not b;
    outputs(2761) <= a xor b;
    outputs(2762) <= b;
    outputs(2763) <= not a or b;
    outputs(2764) <= a;
    outputs(2765) <= not b;
    outputs(2766) <= not b;
    outputs(2767) <= not (a xor b);
    outputs(2768) <= a or b;
    outputs(2769) <= not (a xor b);
    outputs(2770) <= a and b;
    outputs(2771) <= b and not a;
    outputs(2772) <= a;
    outputs(2773) <= not (a xor b);
    outputs(2774) <= a and b;
    outputs(2775) <= a or b;
    outputs(2776) <= not b;
    outputs(2777) <= a xor b;
    outputs(2778) <= not (a xor b);
    outputs(2779) <= a and not b;
    outputs(2780) <= a;
    outputs(2781) <= a and b;
    outputs(2782) <= not b or a;
    outputs(2783) <= a;
    outputs(2784) <= not (a xor b);
    outputs(2785) <= not (a or b);
    outputs(2786) <= a and not b;
    outputs(2787) <= not (a or b);
    outputs(2788) <= a and b;
    outputs(2789) <= b;
    outputs(2790) <= not a;
    outputs(2791) <= not (a xor b);
    outputs(2792) <= b;
    outputs(2793) <= not a;
    outputs(2794) <= a;
    outputs(2795) <= a;
    outputs(2796) <= b;
    outputs(2797) <= not b or a;
    outputs(2798) <= not (a xor b);
    outputs(2799) <= a xor b;
    outputs(2800) <= a;
    outputs(2801) <= a xor b;
    outputs(2802) <= not b;
    outputs(2803) <= b;
    outputs(2804) <= not a;
    outputs(2805) <= b;
    outputs(2806) <= b;
    outputs(2807) <= not (a xor b);
    outputs(2808) <= a and not b;
    outputs(2809) <= a xor b;
    outputs(2810) <= a and not b;
    outputs(2811) <= a or b;
    outputs(2812) <= not a;
    outputs(2813) <= a xor b;
    outputs(2814) <= b;
    outputs(2815) <= not a;
    outputs(2816) <= not a;
    outputs(2817) <= not (a or b);
    outputs(2818) <= a and b;
    outputs(2819) <= not b or a;
    outputs(2820) <= not b;
    outputs(2821) <= not (a or b);
    outputs(2822) <= not (a or b);
    outputs(2823) <= not (a xor b);
    outputs(2824) <= b;
    outputs(2825) <= a xor b;
    outputs(2826) <= not (a and b);
    outputs(2827) <= not a;
    outputs(2828) <= not a;
    outputs(2829) <= a xor b;
    outputs(2830) <= not (a xor b);
    outputs(2831) <= a;
    outputs(2832) <= a;
    outputs(2833) <= b;
    outputs(2834) <= a xor b;
    outputs(2835) <= not (a or b);
    outputs(2836) <= not b;
    outputs(2837) <= a xor b;
    outputs(2838) <= a xor b;
    outputs(2839) <= not (a or b);
    outputs(2840) <= a and b;
    outputs(2841) <= not a;
    outputs(2842) <= a or b;
    outputs(2843) <= a and not b;
    outputs(2844) <= a and b;
    outputs(2845) <= not (a xor b);
    outputs(2846) <= not (a xor b);
    outputs(2847) <= not (a and b);
    outputs(2848) <= b and not a;
    outputs(2849) <= not (a or b);
    outputs(2850) <= not a;
    outputs(2851) <= a xor b;
    outputs(2852) <= a xor b;
    outputs(2853) <= not b;
    outputs(2854) <= a;
    outputs(2855) <= a and not b;
    outputs(2856) <= not (a xor b);
    outputs(2857) <= a xor b;
    outputs(2858) <= b;
    outputs(2859) <= not (a or b);
    outputs(2860) <= a and not b;
    outputs(2861) <= b and not a;
    outputs(2862) <= a and b;
    outputs(2863) <= not b;
    outputs(2864) <= a xor b;
    outputs(2865) <= a xor b;
    outputs(2866) <= not (a xor b);
    outputs(2867) <= not a;
    outputs(2868) <= not (a or b);
    outputs(2869) <= not (a or b);
    outputs(2870) <= not (a xor b);
    outputs(2871) <= not b or a;
    outputs(2872) <= a;
    outputs(2873) <= not b;
    outputs(2874) <= a xor b;
    outputs(2875) <= a xor b;
    outputs(2876) <= not a;
    outputs(2877) <= b;
    outputs(2878) <= b;
    outputs(2879) <= b;
    outputs(2880) <= b and not a;
    outputs(2881) <= not (a xor b);
    outputs(2882) <= not (a xor b);
    outputs(2883) <= not (a xor b);
    outputs(2884) <= b;
    outputs(2885) <= a xor b;
    outputs(2886) <= not (a xor b);
    outputs(2887) <= a or b;
    outputs(2888) <= not (a xor b);
    outputs(2889) <= not (a xor b);
    outputs(2890) <= a and b;
    outputs(2891) <= not a or b;
    outputs(2892) <= a xor b;
    outputs(2893) <= a xor b;
    outputs(2894) <= a and b;
    outputs(2895) <= not a or b;
    outputs(2896) <= a xor b;
    outputs(2897) <= a xor b;
    outputs(2898) <= a xor b;
    outputs(2899) <= b;
    outputs(2900) <= not b;
    outputs(2901) <= not (a xor b);
    outputs(2902) <= not (a or b);
    outputs(2903) <= not a;
    outputs(2904) <= b;
    outputs(2905) <= not a;
    outputs(2906) <= a;
    outputs(2907) <= not a;
    outputs(2908) <= a;
    outputs(2909) <= not (a xor b);
    outputs(2910) <= b and not a;
    outputs(2911) <= a;
    outputs(2912) <= b;
    outputs(2913) <= not a or b;
    outputs(2914) <= a xor b;
    outputs(2915) <= a or b;
    outputs(2916) <= not b or a;
    outputs(2917) <= b and not a;
    outputs(2918) <= a xor b;
    outputs(2919) <= not (a xor b);
    outputs(2920) <= not b or a;
    outputs(2921) <= a xor b;
    outputs(2922) <= a;
    outputs(2923) <= not a;
    outputs(2924) <= b;
    outputs(2925) <= a and b;
    outputs(2926) <= a and b;
    outputs(2927) <= not (a or b);
    outputs(2928) <= not (a xor b);
    outputs(2929) <= b;
    outputs(2930) <= not b;
    outputs(2931) <= not (a or b);
    outputs(2932) <= not b or a;
    outputs(2933) <= not (a xor b);
    outputs(2934) <= a;
    outputs(2935) <= b;
    outputs(2936) <= not (a xor b);
    outputs(2937) <= not b;
    outputs(2938) <= not (a xor b);
    outputs(2939) <= not (a xor b);
    outputs(2940) <= not (a xor b);
    outputs(2941) <= b;
    outputs(2942) <= a xor b;
    outputs(2943) <= b and not a;
    outputs(2944) <= not (a or b);
    outputs(2945) <= not (a or b);
    outputs(2946) <= not b;
    outputs(2947) <= not (a and b);
    outputs(2948) <= not b;
    outputs(2949) <= not b;
    outputs(2950) <= not (a xor b);
    outputs(2951) <= a and not b;
    outputs(2952) <= not (a xor b);
    outputs(2953) <= b and not a;
    outputs(2954) <= not (a xor b);
    outputs(2955) <= b;
    outputs(2956) <= not (a xor b);
    outputs(2957) <= a xor b;
    outputs(2958) <= not (a or b);
    outputs(2959) <= a and b;
    outputs(2960) <= not (a and b);
    outputs(2961) <= a and b;
    outputs(2962) <= a xor b;
    outputs(2963) <= a xor b;
    outputs(2964) <= a xor b;
    outputs(2965) <= a xor b;
    outputs(2966) <= b;
    outputs(2967) <= a;
    outputs(2968) <= a;
    outputs(2969) <= a xor b;
    outputs(2970) <= not b or a;
    outputs(2971) <= not a;
    outputs(2972) <= a xor b;
    outputs(2973) <= not a;
    outputs(2974) <= b and not a;
    outputs(2975) <= a;
    outputs(2976) <= not (a xor b);
    outputs(2977) <= not a or b;
    outputs(2978) <= not b;
    outputs(2979) <= not a;
    outputs(2980) <= a and b;
    outputs(2981) <= not (a xor b);
    outputs(2982) <= a;
    outputs(2983) <= not a or b;
    outputs(2984) <= b;
    outputs(2985) <= a and b;
    outputs(2986) <= not a;
    outputs(2987) <= not b;
    outputs(2988) <= not b;
    outputs(2989) <= not (a xor b);
    outputs(2990) <= not (a xor b);
    outputs(2991) <= a xor b;
    outputs(2992) <= a and not b;
    outputs(2993) <= a xor b;
    outputs(2994) <= a and not b;
    outputs(2995) <= not (a or b);
    outputs(2996) <= a and not b;
    outputs(2997) <= not (a xor b);
    outputs(2998) <= not (a and b);
    outputs(2999) <= b;
    outputs(3000) <= a;
    outputs(3001) <= a xor b;
    outputs(3002) <= a;
    outputs(3003) <= not a or b;
    outputs(3004) <= not (a or b);
    outputs(3005) <= b;
    outputs(3006) <= a and not b;
    outputs(3007) <= not (a xor b);
    outputs(3008) <= not a;
    outputs(3009) <= a or b;
    outputs(3010) <= a and b;
    outputs(3011) <= b;
    outputs(3012) <= not b;
    outputs(3013) <= a or b;
    outputs(3014) <= b;
    outputs(3015) <= a xor b;
    outputs(3016) <= not (a xor b);
    outputs(3017) <= not (a or b);
    outputs(3018) <= b;
    outputs(3019) <= not (a xor b);
    outputs(3020) <= not a;
    outputs(3021) <= a and b;
    outputs(3022) <= a xor b;
    outputs(3023) <= not (a or b);
    outputs(3024) <= b and not a;
    outputs(3025) <= not b;
    outputs(3026) <= a and not b;
    outputs(3027) <= a;
    outputs(3028) <= not (a and b);
    outputs(3029) <= not b or a;
    outputs(3030) <= b and not a;
    outputs(3031) <= not b;
    outputs(3032) <= a;
    outputs(3033) <= not a or b;
    outputs(3034) <= a;
    outputs(3035) <= not (a xor b);
    outputs(3036) <= not (a xor b);
    outputs(3037) <= a xor b;
    outputs(3038) <= b;
    outputs(3039) <= a or b;
    outputs(3040) <= b;
    outputs(3041) <= not a or b;
    outputs(3042) <= not a;
    outputs(3043) <= a;
    outputs(3044) <= not (a and b);
    outputs(3045) <= not a;
    outputs(3046) <= b;
    outputs(3047) <= not (a and b);
    outputs(3048) <= b;
    outputs(3049) <= not (a xor b);
    outputs(3050) <= b;
    outputs(3051) <= not b;
    outputs(3052) <= not b;
    outputs(3053) <= a xor b;
    outputs(3054) <= not (a and b);
    outputs(3055) <= a and b;
    outputs(3056) <= not (a and b);
    outputs(3057) <= not b;
    outputs(3058) <= a xor b;
    outputs(3059) <= a and not b;
    outputs(3060) <= a xor b;
    outputs(3061) <= a;
    outputs(3062) <= not b;
    outputs(3063) <= a and not b;
    outputs(3064) <= a xor b;
    outputs(3065) <= a;
    outputs(3066) <= not (a or b);
    outputs(3067) <= not a or b;
    outputs(3068) <= b and not a;
    outputs(3069) <= not b;
    outputs(3070) <= a xor b;
    outputs(3071) <= not a;
    outputs(3072) <= not (a and b);
    outputs(3073) <= a and not b;
    outputs(3074) <= b;
    outputs(3075) <= not (a and b);
    outputs(3076) <= not a;
    outputs(3077) <= b and not a;
    outputs(3078) <= not b;
    outputs(3079) <= a or b;
    outputs(3080) <= not (a xor b);
    outputs(3081) <= not (a xor b);
    outputs(3082) <= not (a xor b);
    outputs(3083) <= not (a xor b);
    outputs(3084) <= not a;
    outputs(3085) <= not (a or b);
    outputs(3086) <= not (a xor b);
    outputs(3087) <= a;
    outputs(3088) <= a and not b;
    outputs(3089) <= a and b;
    outputs(3090) <= not b;
    outputs(3091) <= not a or b;
    outputs(3092) <= b;
    outputs(3093) <= not (a or b);
    outputs(3094) <= a and not b;
    outputs(3095) <= not (a or b);
    outputs(3096) <= a;
    outputs(3097) <= not (a xor b);
    outputs(3098) <= not (a xor b);
    outputs(3099) <= a and b;
    outputs(3100) <= not (a xor b);
    outputs(3101) <= '1';
    outputs(3102) <= not (a xor b);
    outputs(3103) <= not a;
    outputs(3104) <= not a or b;
    outputs(3105) <= not (a xor b);
    outputs(3106) <= a xor b;
    outputs(3107) <= not b;
    outputs(3108) <= a and not b;
    outputs(3109) <= a;
    outputs(3110) <= not b;
    outputs(3111) <= not a;
    outputs(3112) <= not b;
    outputs(3113) <= not b;
    outputs(3114) <= not b;
    outputs(3115) <= not (a or b);
    outputs(3116) <= a;
    outputs(3117) <= a and not b;
    outputs(3118) <= a and b;
    outputs(3119) <= a xor b;
    outputs(3120) <= a;
    outputs(3121) <= b;
    outputs(3122) <= a and not b;
    outputs(3123) <= not b;
    outputs(3124) <= b;
    outputs(3125) <= not b;
    outputs(3126) <= a and b;
    outputs(3127) <= not b;
    outputs(3128) <= not a;
    outputs(3129) <= a and not b;
    outputs(3130) <= a;
    outputs(3131) <= b and not a;
    outputs(3132) <= a;
    outputs(3133) <= not b;
    outputs(3134) <= not (a and b);
    outputs(3135) <= not (a and b);
    outputs(3136) <= not (a or b);
    outputs(3137) <= not a;
    outputs(3138) <= not (a xor b);
    outputs(3139) <= b and not a;
    outputs(3140) <= not (a or b);
    outputs(3141) <= b and not a;
    outputs(3142) <= not a or b;
    outputs(3143) <= b;
    outputs(3144) <= not b;
    outputs(3145) <= b and not a;
    outputs(3146) <= a and b;
    outputs(3147) <= a or b;
    outputs(3148) <= a xor b;
    outputs(3149) <= not (a xor b);
    outputs(3150) <= a xor b;
    outputs(3151) <= not (a xor b);
    outputs(3152) <= not (a or b);
    outputs(3153) <= not (a or b);
    outputs(3154) <= not b;
    outputs(3155) <= not (a or b);
    outputs(3156) <= a and not b;
    outputs(3157) <= not (a xor b);
    outputs(3158) <= b and not a;
    outputs(3159) <= a and not b;
    outputs(3160) <= not (a or b);
    outputs(3161) <= a;
    outputs(3162) <= not (a or b);
    outputs(3163) <= not (a or b);
    outputs(3164) <= not (a or b);
    outputs(3165) <= not a or b;
    outputs(3166) <= not (a and b);
    outputs(3167) <= b;
    outputs(3168) <= b and not a;
    outputs(3169) <= b;
    outputs(3170) <= not a;
    outputs(3171) <= not (a xor b);
    outputs(3172) <= a and not b;
    outputs(3173) <= not a;
    outputs(3174) <= a xor b;
    outputs(3175) <= not (a or b);
    outputs(3176) <= not (a and b);
    outputs(3177) <= a and not b;
    outputs(3178) <= not (a xor b);
    outputs(3179) <= b;
    outputs(3180) <= a or b;
    outputs(3181) <= not (a or b);
    outputs(3182) <= not a;
    outputs(3183) <= not b or a;
    outputs(3184) <= a;
    outputs(3185) <= a xor b;
    outputs(3186) <= not a or b;
    outputs(3187) <= a xor b;
    outputs(3188) <= not a or b;
    outputs(3189) <= a and not b;
    outputs(3190) <= not (a xor b);
    outputs(3191) <= a xor b;
    outputs(3192) <= b;
    outputs(3193) <= not b;
    outputs(3194) <= a and not b;
    outputs(3195) <= a xor b;
    outputs(3196) <= b;
    outputs(3197) <= not a;
    outputs(3198) <= not a;
    outputs(3199) <= not a;
    outputs(3200) <= not (a xor b);
    outputs(3201) <= a and b;
    outputs(3202) <= not (a or b);
    outputs(3203) <= not (a xor b);
    outputs(3204) <= not b;
    outputs(3205) <= a and not b;
    outputs(3206) <= not a;
    outputs(3207) <= not b;
    outputs(3208) <= not (a xor b);
    outputs(3209) <= b;
    outputs(3210) <= a and b;
    outputs(3211) <= a and b;
    outputs(3212) <= not a;
    outputs(3213) <= not a;
    outputs(3214) <= b and not a;
    outputs(3215) <= not b;
    outputs(3216) <= a and b;
    outputs(3217) <= not (a xor b);
    outputs(3218) <= not a or b;
    outputs(3219) <= not b or a;
    outputs(3220) <= a xor b;
    outputs(3221) <= a and b;
    outputs(3222) <= a and not b;
    outputs(3223) <= a and not b;
    outputs(3224) <= a or b;
    outputs(3225) <= not (a xor b);
    outputs(3226) <= a xor b;
    outputs(3227) <= b and not a;
    outputs(3228) <= a and b;
    outputs(3229) <= not (a or b);
    outputs(3230) <= not (a xor b);
    outputs(3231) <= not a;
    outputs(3232) <= b;
    outputs(3233) <= not (a xor b);
    outputs(3234) <= a and b;
    outputs(3235) <= a and not b;
    outputs(3236) <= a xor b;
    outputs(3237) <= not (a xor b);
    outputs(3238) <= not (a xor b);
    outputs(3239) <= not (a or b);
    outputs(3240) <= a and not b;
    outputs(3241) <= b;
    outputs(3242) <= '0';
    outputs(3243) <= not (a xor b);
    outputs(3244) <= not b;
    outputs(3245) <= a;
    outputs(3246) <= not a;
    outputs(3247) <= a and b;
    outputs(3248) <= not (a xor b);
    outputs(3249) <= a;
    outputs(3250) <= not a or b;
    outputs(3251) <= a xor b;
    outputs(3252) <= not b;
    outputs(3253) <= b;
    outputs(3254) <= not (a xor b);
    outputs(3255) <= a and b;
    outputs(3256) <= a xor b;
    outputs(3257) <= b;
    outputs(3258) <= not a;
    outputs(3259) <= not a;
    outputs(3260) <= not a;
    outputs(3261) <= not a;
    outputs(3262) <= not b or a;
    outputs(3263) <= not (a or b);
    outputs(3264) <= not (a or b);
    outputs(3265) <= a xor b;
    outputs(3266) <= a xor b;
    outputs(3267) <= a and b;
    outputs(3268) <= not (a xor b);
    outputs(3269) <= a xor b;
    outputs(3270) <= not a;
    outputs(3271) <= not (a or b);
    outputs(3272) <= not a;
    outputs(3273) <= not (a xor b);
    outputs(3274) <= a;
    outputs(3275) <= a xor b;
    outputs(3276) <= a xor b;
    outputs(3277) <= a or b;
    outputs(3278) <= not (a or b);
    outputs(3279) <= b;
    outputs(3280) <= a and not b;
    outputs(3281) <= b;
    outputs(3282) <= not b;
    outputs(3283) <= a;
    outputs(3284) <= b;
    outputs(3285) <= not (a and b);
    outputs(3286) <= not (a xor b);
    outputs(3287) <= not b or a;
    outputs(3288) <= not b;
    outputs(3289) <= not (a and b);
    outputs(3290) <= not (a or b);
    outputs(3291) <= a;
    outputs(3292) <= not a;
    outputs(3293) <= not (a xor b);
    outputs(3294) <= a and not b;
    outputs(3295) <= a and not b;
    outputs(3296) <= not (a xor b);
    outputs(3297) <= a;
    outputs(3298) <= not a;
    outputs(3299) <= not a;
    outputs(3300) <= a and not b;
    outputs(3301) <= a xor b;
    outputs(3302) <= b and not a;
    outputs(3303) <= a and not b;
    outputs(3304) <= not b;
    outputs(3305) <= not (a xor b);
    outputs(3306) <= b;
    outputs(3307) <= a and b;
    outputs(3308) <= a;
    outputs(3309) <= a and b;
    outputs(3310) <= not (a and b);
    outputs(3311) <= a and b;
    outputs(3312) <= not (a or b);
    outputs(3313) <= not a;
    outputs(3314) <= not a;
    outputs(3315) <= not (a xor b);
    outputs(3316) <= not (a xor b);
    outputs(3317) <= a xor b;
    outputs(3318) <= not (a xor b);
    outputs(3319) <= not (a xor b);
    outputs(3320) <= a and not b;
    outputs(3321) <= not a;
    outputs(3322) <= a and not b;
    outputs(3323) <= not (a or b);
    outputs(3324) <= a;
    outputs(3325) <= a and b;
    outputs(3326) <= not a;
    outputs(3327) <= not a or b;
    outputs(3328) <= not a or b;
    outputs(3329) <= a and b;
    outputs(3330) <= not b;
    outputs(3331) <= a and not b;
    outputs(3332) <= not b;
    outputs(3333) <= not (a xor b);
    outputs(3334) <= not a or b;
    outputs(3335) <= not (a and b);
    outputs(3336) <= a xor b;
    outputs(3337) <= b and not a;
    outputs(3338) <= a and b;
    outputs(3339) <= not b;
    outputs(3340) <= not (a or b);
    outputs(3341) <= a or b;
    outputs(3342) <= not (a xor b);
    outputs(3343) <= not b;
    outputs(3344) <= not (a or b);
    outputs(3345) <= b and not a;
    outputs(3346) <= not (a xor b);
    outputs(3347) <= b and not a;
    outputs(3348) <= not b;
    outputs(3349) <= not (a or b);
    outputs(3350) <= a;
    outputs(3351) <= not b;
    outputs(3352) <= a and b;
    outputs(3353) <= a and not b;
    outputs(3354) <= not b;
    outputs(3355) <= b and not a;
    outputs(3356) <= a or b;
    outputs(3357) <= a xor b;
    outputs(3358) <= b and not a;
    outputs(3359) <= not b;
    outputs(3360) <= a;
    outputs(3361) <= a xor b;
    outputs(3362) <= not a;
    outputs(3363) <= not (a or b);
    outputs(3364) <= b and not a;
    outputs(3365) <= not b;
    outputs(3366) <= not b;
    outputs(3367) <= not (a xor b);
    outputs(3368) <= not a;
    outputs(3369) <= b and not a;
    outputs(3370) <= not a;
    outputs(3371) <= a xor b;
    outputs(3372) <= not (a xor b);
    outputs(3373) <= b;
    outputs(3374) <= not a;
    outputs(3375) <= b and not a;
    outputs(3376) <= not a;
    outputs(3377) <= a;
    outputs(3378) <= a and not b;
    outputs(3379) <= not b;
    outputs(3380) <= b;
    outputs(3381) <= not a or b;
    outputs(3382) <= not (a or b);
    outputs(3383) <= b and not a;
    outputs(3384) <= a and not b;
    outputs(3385) <= not b;
    outputs(3386) <= a xor b;
    outputs(3387) <= b and not a;
    outputs(3388) <= not b;
    outputs(3389) <= not b;
    outputs(3390) <= a xor b;
    outputs(3391) <= not b;
    outputs(3392) <= not b;
    outputs(3393) <= not a or b;
    outputs(3394) <= not (a xor b);
    outputs(3395) <= a and b;
    outputs(3396) <= a xor b;
    outputs(3397) <= not (a xor b);
    outputs(3398) <= a;
    outputs(3399) <= a;
    outputs(3400) <= b and not a;
    outputs(3401) <= b and not a;
    outputs(3402) <= a xor b;
    outputs(3403) <= a;
    outputs(3404) <= not (a or b);
    outputs(3405) <= a;
    outputs(3406) <= b;
    outputs(3407) <= b;
    outputs(3408) <= not b;
    outputs(3409) <= a and b;
    outputs(3410) <= b and not a;
    outputs(3411) <= not a;
    outputs(3412) <= not (a or b);
    outputs(3413) <= not a;
    outputs(3414) <= a xor b;
    outputs(3415) <= not a;
    outputs(3416) <= not b or a;
    outputs(3417) <= b;
    outputs(3418) <= a or b;
    outputs(3419) <= not (a xor b);
    outputs(3420) <= a and b;
    outputs(3421) <= a xor b;
    outputs(3422) <= not a or b;
    outputs(3423) <= not a or b;
    outputs(3424) <= a xor b;
    outputs(3425) <= b and not a;
    outputs(3426) <= a or b;
    outputs(3427) <= not (a xor b);
    outputs(3428) <= a and b;
    outputs(3429) <= b;
    outputs(3430) <= a xor b;
    outputs(3431) <= not b or a;
    outputs(3432) <= b;
    outputs(3433) <= not (a or b);
    outputs(3434) <= not a;
    outputs(3435) <= a xor b;
    outputs(3436) <= a and b;
    outputs(3437) <= a and b;
    outputs(3438) <= not b or a;
    outputs(3439) <= not b;
    outputs(3440) <= not b;
    outputs(3441) <= not b;
    outputs(3442) <= not a or b;
    outputs(3443) <= not a;
    outputs(3444) <= a xor b;
    outputs(3445) <= not a;
    outputs(3446) <= b and not a;
    outputs(3447) <= a;
    outputs(3448) <= a and not b;
    outputs(3449) <= a;
    outputs(3450) <= not b;
    outputs(3451) <= not (a or b);
    outputs(3452) <= b;
    outputs(3453) <= not b;
    outputs(3454) <= not b;
    outputs(3455) <= a;
    outputs(3456) <= not b;
    outputs(3457) <= not a;
    outputs(3458) <= not b;
    outputs(3459) <= not a;
    outputs(3460) <= not (a xor b);
    outputs(3461) <= b;
    outputs(3462) <= not (a xor b);
    outputs(3463) <= a xor b;
    outputs(3464) <= not b or a;
    outputs(3465) <= b and not a;
    outputs(3466) <= not a;
    outputs(3467) <= b;
    outputs(3468) <= a xor b;
    outputs(3469) <= not a;
    outputs(3470) <= a and not b;
    outputs(3471) <= b;
    outputs(3472) <= not a;
    outputs(3473) <= a and b;
    outputs(3474) <= a and not b;
    outputs(3475) <= not a or b;
    outputs(3476) <= b and not a;
    outputs(3477) <= a xor b;
    outputs(3478) <= not (a or b);
    outputs(3479) <= a xor b;
    outputs(3480) <= b;
    outputs(3481) <= not b;
    outputs(3482) <= a or b;
    outputs(3483) <= b and not a;
    outputs(3484) <= not b;
    outputs(3485) <= b and not a;
    outputs(3486) <= a;
    outputs(3487) <= not a or b;
    outputs(3488) <= a;
    outputs(3489) <= not b;
    outputs(3490) <= a xor b;
    outputs(3491) <= a or b;
    outputs(3492) <= b;
    outputs(3493) <= not (a xor b);
    outputs(3494) <= a xor b;
    outputs(3495) <= b and not a;
    outputs(3496) <= a and not b;
    outputs(3497) <= b;
    outputs(3498) <= a and b;
    outputs(3499) <= not (a and b);
    outputs(3500) <= not b;
    outputs(3501) <= not b or a;
    outputs(3502) <= b;
    outputs(3503) <= b;
    outputs(3504) <= not (a xor b);
    outputs(3505) <= a and b;
    outputs(3506) <= not (a xor b);
    outputs(3507) <= b;
    outputs(3508) <= not b or a;
    outputs(3509) <= a xor b;
    outputs(3510) <= b;
    outputs(3511) <= b;
    outputs(3512) <= a xor b;
    outputs(3513) <= a and b;
    outputs(3514) <= not b;
    outputs(3515) <= a;
    outputs(3516) <= not b;
    outputs(3517) <= not b or a;
    outputs(3518) <= a xor b;
    outputs(3519) <= not b;
    outputs(3520) <= a xor b;
    outputs(3521) <= b and not a;
    outputs(3522) <= b;
    outputs(3523) <= a or b;
    outputs(3524) <= b;
    outputs(3525) <= a and b;
    outputs(3526) <= b and not a;
    outputs(3527) <= b and not a;
    outputs(3528) <= a xor b;
    outputs(3529) <= b and not a;
    outputs(3530) <= not (a xor b);
    outputs(3531) <= not a;
    outputs(3532) <= a and b;
    outputs(3533) <= not (a and b);
    outputs(3534) <= b;
    outputs(3535) <= b;
    outputs(3536) <= not b;
    outputs(3537) <= a;
    outputs(3538) <= not a;
    outputs(3539) <= not a;
    outputs(3540) <= a xor b;
    outputs(3541) <= a and not b;
    outputs(3542) <= b;
    outputs(3543) <= a;
    outputs(3544) <= not (a xor b);
    outputs(3545) <= not (a xor b);
    outputs(3546) <= not a;
    outputs(3547) <= b;
    outputs(3548) <= b and not a;
    outputs(3549) <= not b or a;
    outputs(3550) <= b;
    outputs(3551) <= not b;
    outputs(3552) <= a xor b;
    outputs(3553) <= not a;
    outputs(3554) <= not a;
    outputs(3555) <= not a;
    outputs(3556) <= a;
    outputs(3557) <= not (a or b);
    outputs(3558) <= not (a or b);
    outputs(3559) <= a and not b;
    outputs(3560) <= a xor b;
    outputs(3561) <= not b;
    outputs(3562) <= not (a or b);
    outputs(3563) <= a;
    outputs(3564) <= not a or b;
    outputs(3565) <= a;
    outputs(3566) <= a xor b;
    outputs(3567) <= not b;
    outputs(3568) <= a and not b;
    outputs(3569) <= a or b;
    outputs(3570) <= a and not b;
    outputs(3571) <= not b;
    outputs(3572) <= a;
    outputs(3573) <= a xor b;
    outputs(3574) <= b;
    outputs(3575) <= a;
    outputs(3576) <= b and not a;
    outputs(3577) <= not (a xor b);
    outputs(3578) <= not (a xor b);
    outputs(3579) <= a;
    outputs(3580) <= not (a or b);
    outputs(3581) <= a xor b;
    outputs(3582) <= not b;
    outputs(3583) <= not (a or b);
    outputs(3584) <= a and b;
    outputs(3585) <= b;
    outputs(3586) <= not a;
    outputs(3587) <= b;
    outputs(3588) <= not a;
    outputs(3589) <= a;
    outputs(3590) <= b and not a;
    outputs(3591) <= a and b;
    outputs(3592) <= a;
    outputs(3593) <= not (a xor b);
    outputs(3594) <= a and b;
    outputs(3595) <= not (a xor b);
    outputs(3596) <= a xor b;
    outputs(3597) <= b;
    outputs(3598) <= not (a xor b);
    outputs(3599) <= not (a or b);
    outputs(3600) <= a;
    outputs(3601) <= a or b;
    outputs(3602) <= a and b;
    outputs(3603) <= not (a or b);
    outputs(3604) <= not (a xor b);
    outputs(3605) <= a and b;
    outputs(3606) <= a and not b;
    outputs(3607) <= not a or b;
    outputs(3608) <= not b or a;
    outputs(3609) <= not b or a;
    outputs(3610) <= not (a and b);
    outputs(3611) <= not (a or b);
    outputs(3612) <= b;
    outputs(3613) <= b and not a;
    outputs(3614) <= not (a or b);
    outputs(3615) <= a xor b;
    outputs(3616) <= not a;
    outputs(3617) <= a;
    outputs(3618) <= a;
    outputs(3619) <= a;
    outputs(3620) <= not (a or b);
    outputs(3621) <= not (a and b);
    outputs(3622) <= not b;
    outputs(3623) <= b and not a;
    outputs(3624) <= not a;
    outputs(3625) <= not (a or b);
    outputs(3626) <= b;
    outputs(3627) <= a and b;
    outputs(3628) <= b and not a;
    outputs(3629) <= b and not a;
    outputs(3630) <= a and b;
    outputs(3631) <= a and b;
    outputs(3632) <= not a;
    outputs(3633) <= not b or a;
    outputs(3634) <= b and not a;
    outputs(3635) <= not (a and b);
    outputs(3636) <= not a or b;
    outputs(3637) <= not (a or b);
    outputs(3638) <= not b;
    outputs(3639) <= a;
    outputs(3640) <= a and b;
    outputs(3641) <= not a;
    outputs(3642) <= not (a or b);
    outputs(3643) <= a or b;
    outputs(3644) <= a and not b;
    outputs(3645) <= a;
    outputs(3646) <= not a or b;
    outputs(3647) <= b and not a;
    outputs(3648) <= b;
    outputs(3649) <= not a;
    outputs(3650) <= b;
    outputs(3651) <= b;
    outputs(3652) <= not (a or b);
    outputs(3653) <= b and not a;
    outputs(3654) <= a and not b;
    outputs(3655) <= b;
    outputs(3656) <= not b;
    outputs(3657) <= not a;
    outputs(3658) <= a and not b;
    outputs(3659) <= b;
    outputs(3660) <= a and not b;
    outputs(3661) <= not a or b;
    outputs(3662) <= not a;
    outputs(3663) <= not (a or b);
    outputs(3664) <= a xor b;
    outputs(3665) <= b;
    outputs(3666) <= a and b;
    outputs(3667) <= not b;
    outputs(3668) <= a and b;
    outputs(3669) <= a xor b;
    outputs(3670) <= not (a xor b);
    outputs(3671) <= not b or a;
    outputs(3672) <= not a or b;
    outputs(3673) <= not (a or b);
    outputs(3674) <= a and not b;
    outputs(3675) <= a and b;
    outputs(3676) <= not b;
    outputs(3677) <= not a;
    outputs(3678) <= a xor b;
    outputs(3679) <= b and not a;
    outputs(3680) <= a or b;
    outputs(3681) <= a and not b;
    outputs(3682) <= a and not b;
    outputs(3683) <= a;
    outputs(3684) <= not b;
    outputs(3685) <= a;
    outputs(3686) <= a and b;
    outputs(3687) <= not (a or b);
    outputs(3688) <= b;
    outputs(3689) <= a;
    outputs(3690) <= not (a and b);
    outputs(3691) <= not a;
    outputs(3692) <= a and not b;
    outputs(3693) <= not b or a;
    outputs(3694) <= b;
    outputs(3695) <= not (a xor b);
    outputs(3696) <= a and not b;
    outputs(3697) <= not a;
    outputs(3698) <= a;
    outputs(3699) <= a and b;
    outputs(3700) <= not a;
    outputs(3701) <= a and b;
    outputs(3702) <= a;
    outputs(3703) <= not (a or b);
    outputs(3704) <= a xor b;
    outputs(3705) <= a and b;
    outputs(3706) <= a and b;
    outputs(3707) <= not (a or b);
    outputs(3708) <= not (a xor b);
    outputs(3709) <= not a;
    outputs(3710) <= a and b;
    outputs(3711) <= a;
    outputs(3712) <= not a;
    outputs(3713) <= not (a or b);
    outputs(3714) <= a and b;
    outputs(3715) <= b;
    outputs(3716) <= not b or a;
    outputs(3717) <= b;
    outputs(3718) <= not (a xor b);
    outputs(3719) <= a;
    outputs(3720) <= a or b;
    outputs(3721) <= not b;
    outputs(3722) <= not (a and b);
    outputs(3723) <= a xor b;
    outputs(3724) <= a or b;
    outputs(3725) <= not (a xor b);
    outputs(3726) <= a;
    outputs(3727) <= not (a xor b);
    outputs(3728) <= b and not a;
    outputs(3729) <= a;
    outputs(3730) <= b and not a;
    outputs(3731) <= a;
    outputs(3732) <= b;
    outputs(3733) <= a xor b;
    outputs(3734) <= b and not a;
    outputs(3735) <= a;
    outputs(3736) <= a;
    outputs(3737) <= b and not a;
    outputs(3738) <= a and b;
    outputs(3739) <= a xor b;
    outputs(3740) <= a and not b;
    outputs(3741) <= not (a or b);
    outputs(3742) <= b;
    outputs(3743) <= not (a and b);
    outputs(3744) <= not a;
    outputs(3745) <= b;
    outputs(3746) <= b;
    outputs(3747) <= not (a xor b);
    outputs(3748) <= not b or a;
    outputs(3749) <= a and b;
    outputs(3750) <= a and not b;
    outputs(3751) <= not (a or b);
    outputs(3752) <= not (a or b);
    outputs(3753) <= b and not a;
    outputs(3754) <= not a or b;
    outputs(3755) <= not a;
    outputs(3756) <= not a;
    outputs(3757) <= not b;
    outputs(3758) <= a xor b;
    outputs(3759) <= not a;
    outputs(3760) <= b;
    outputs(3761) <= a and b;
    outputs(3762) <= b and not a;
    outputs(3763) <= a or b;
    outputs(3764) <= a;
    outputs(3765) <= a xor b;
    outputs(3766) <= b;
    outputs(3767) <= a;
    outputs(3768) <= b and not a;
    outputs(3769) <= a;
    outputs(3770) <= b and not a;
    outputs(3771) <= a and not b;
    outputs(3772) <= b and not a;
    outputs(3773) <= not (a and b);
    outputs(3774) <= not a;
    outputs(3775) <= not b or a;
    outputs(3776) <= not b;
    outputs(3777) <= b and not a;
    outputs(3778) <= a;
    outputs(3779) <= a and b;
    outputs(3780) <= not b;
    outputs(3781) <= not b;
    outputs(3782) <= a xor b;
    outputs(3783) <= a and not b;
    outputs(3784) <= not (a or b);
    outputs(3785) <= a and not b;
    outputs(3786) <= not a;
    outputs(3787) <= b and not a;
    outputs(3788) <= a xor b;
    outputs(3789) <= not a;
    outputs(3790) <= not (a xor b);
    outputs(3791) <= not (a or b);
    outputs(3792) <= not (a or b);
    outputs(3793) <= not b;
    outputs(3794) <= b;
    outputs(3795) <= not a;
    outputs(3796) <= not a;
    outputs(3797) <= not (a xor b);
    outputs(3798) <= not (a and b);
    outputs(3799) <= not a;
    outputs(3800) <= not a;
    outputs(3801) <= a and not b;
    outputs(3802) <= a and b;
    outputs(3803) <= not a;
    outputs(3804) <= not a;
    outputs(3805) <= not a;
    outputs(3806) <= a and b;
    outputs(3807) <= not (a xor b);
    outputs(3808) <= b and not a;
    outputs(3809) <= not (a or b);
    outputs(3810) <= a;
    outputs(3811) <= a and b;
    outputs(3812) <= not b;
    outputs(3813) <= a and not b;
    outputs(3814) <= not b;
    outputs(3815) <= a;
    outputs(3816) <= a and b;
    outputs(3817) <= a and b;
    outputs(3818) <= b;
    outputs(3819) <= not b;
    outputs(3820) <= a xor b;
    outputs(3821) <= b;
    outputs(3822) <= a;
    outputs(3823) <= not b;
    outputs(3824) <= not (a or b);
    outputs(3825) <= not b;
    outputs(3826) <= not a;
    outputs(3827) <= not a;
    outputs(3828) <= not a;
    outputs(3829) <= not a or b;
    outputs(3830) <= not b;
    outputs(3831) <= a and b;
    outputs(3832) <= not a;
    outputs(3833) <= b and not a;
    outputs(3834) <= not (a xor b);
    outputs(3835) <= not a;
    outputs(3836) <= a and not b;
    outputs(3837) <= a and b;
    outputs(3838) <= not (a xor b);
    outputs(3839) <= b;
    outputs(3840) <= not a;
    outputs(3841) <= a and b;
    outputs(3842) <= not (a xor b);
    outputs(3843) <= not (a xor b);
    outputs(3844) <= b;
    outputs(3845) <= not (a xor b);
    outputs(3846) <= not (a xor b);
    outputs(3847) <= not (a xor b);
    outputs(3848) <= a;
    outputs(3849) <= not a;
    outputs(3850) <= a and not b;
    outputs(3851) <= not (a or b);
    outputs(3852) <= a xor b;
    outputs(3853) <= b and not a;
    outputs(3854) <= not a;
    outputs(3855) <= not (a or b);
    outputs(3856) <= a and not b;
    outputs(3857) <= not b or a;
    outputs(3858) <= b;
    outputs(3859) <= not (a or b);
    outputs(3860) <= a and b;
    outputs(3861) <= a;
    outputs(3862) <= not (a xor b);
    outputs(3863) <= b;
    outputs(3864) <= b and not a;
    outputs(3865) <= not a;
    outputs(3866) <= a;
    outputs(3867) <= a and b;
    outputs(3868) <= a;
    outputs(3869) <= a and not b;
    outputs(3870) <= a;
    outputs(3871) <= b;
    outputs(3872) <= not (a and b);
    outputs(3873) <= a xor b;
    outputs(3874) <= not b;
    outputs(3875) <= a and b;
    outputs(3876) <= a;
    outputs(3877) <= not a;
    outputs(3878) <= not a;
    outputs(3879) <= b;
    outputs(3880) <= b;
    outputs(3881) <= a xor b;
    outputs(3882) <= a xor b;
    outputs(3883) <= b;
    outputs(3884) <= a and b;
    outputs(3885) <= b and not a;
    outputs(3886) <= a and not b;
    outputs(3887) <= b;
    outputs(3888) <= not a;
    outputs(3889) <= a and b;
    outputs(3890) <= a and not b;
    outputs(3891) <= not b or a;
    outputs(3892) <= not a;
    outputs(3893) <= a;
    outputs(3894) <= not (a or b);
    outputs(3895) <= a;
    outputs(3896) <= a and b;
    outputs(3897) <= a xor b;
    outputs(3898) <= a or b;
    outputs(3899) <= not b or a;
    outputs(3900) <= not (a xor b);
    outputs(3901) <= not a or b;
    outputs(3902) <= a;
    outputs(3903) <= not b or a;
    outputs(3904) <= a and not b;
    outputs(3905) <= a and not b;
    outputs(3906) <= b and not a;
    outputs(3907) <= not b or a;
    outputs(3908) <= a;
    outputs(3909) <= not a;
    outputs(3910) <= a and b;
    outputs(3911) <= b;
    outputs(3912) <= not (a xor b);
    outputs(3913) <= not (a xor b);
    outputs(3914) <= b;
    outputs(3915) <= a or b;
    outputs(3916) <= b;
    outputs(3917) <= not (a and b);
    outputs(3918) <= not (a or b);
    outputs(3919) <= a and b;
    outputs(3920) <= a and b;
    outputs(3921) <= not a;
    outputs(3922) <= b;
    outputs(3923) <= a and not b;
    outputs(3924) <= a;
    outputs(3925) <= a xor b;
    outputs(3926) <= a;
    outputs(3927) <= a and b;
    outputs(3928) <= a and not b;
    outputs(3929) <= a and not b;
    outputs(3930) <= a xor b;
    outputs(3931) <= b;
    outputs(3932) <= not (a xor b);
    outputs(3933) <= a xor b;
    outputs(3934) <= a;
    outputs(3935) <= b and not a;
    outputs(3936) <= a and not b;
    outputs(3937) <= b and not a;
    outputs(3938) <= not b;
    outputs(3939) <= not b;
    outputs(3940) <= a xor b;
    outputs(3941) <= not (a and b);
    outputs(3942) <= not b or a;
    outputs(3943) <= not b;
    outputs(3944) <= b and not a;
    outputs(3945) <= b;
    outputs(3946) <= a;
    outputs(3947) <= not (a xor b);
    outputs(3948) <= b;
    outputs(3949) <= a and b;
    outputs(3950) <= a xor b;
    outputs(3951) <= a and not b;
    outputs(3952) <= not a;
    outputs(3953) <= not a;
    outputs(3954) <= not b;
    outputs(3955) <= b and not a;
    outputs(3956) <= a xor b;
    outputs(3957) <= not (a xor b);
    outputs(3958) <= not a;
    outputs(3959) <= not a;
    outputs(3960) <= not b;
    outputs(3961) <= not (a or b);
    outputs(3962) <= a or b;
    outputs(3963) <= a;
    outputs(3964) <= not (a xor b);
    outputs(3965) <= not (a xor b);
    outputs(3966) <= a and b;
    outputs(3967) <= not (a xor b);
    outputs(3968) <= not (a xor b);
    outputs(3969) <= a xor b;
    outputs(3970) <= a xor b;
    outputs(3971) <= not (a or b);
    outputs(3972) <= b and not a;
    outputs(3973) <= b;
    outputs(3974) <= b and not a;
    outputs(3975) <= a and not b;
    outputs(3976) <= not (a and b);
    outputs(3977) <= a;
    outputs(3978) <= not a;
    outputs(3979) <= not a;
    outputs(3980) <= not (a xor b);
    outputs(3981) <= not a;
    outputs(3982) <= not a;
    outputs(3983) <= b;
    outputs(3984) <= not a;
    outputs(3985) <= not b or a;
    outputs(3986) <= not b;
    outputs(3987) <= a xor b;
    outputs(3988) <= a;
    outputs(3989) <= a;
    outputs(3990) <= a and not b;
    outputs(3991) <= a and b;
    outputs(3992) <= not (a xor b);
    outputs(3993) <= not (a or b);
    outputs(3994) <= a;
    outputs(3995) <= b;
    outputs(3996) <= a and b;
    outputs(3997) <= b and not a;
    outputs(3998) <= not a or b;
    outputs(3999) <= a;
    outputs(4000) <= not a;
    outputs(4001) <= b;
    outputs(4002) <= not b;
    outputs(4003) <= b;
    outputs(4004) <= a or b;
    outputs(4005) <= a;
    outputs(4006) <= a xor b;
    outputs(4007) <= not (a or b);
    outputs(4008) <= not (a or b);
    outputs(4009) <= b;
    outputs(4010) <= not (a or b);
    outputs(4011) <= a;
    outputs(4012) <= a and b;
    outputs(4013) <= not (a xor b);
    outputs(4014) <= not (a xor b);
    outputs(4015) <= a xor b;
    outputs(4016) <= a and b;
    outputs(4017) <= a or b;
    outputs(4018) <= a;
    outputs(4019) <= not b;
    outputs(4020) <= not b or a;
    outputs(4021) <= a or b;
    outputs(4022) <= not a;
    outputs(4023) <= a xor b;
    outputs(4024) <= a xor b;
    outputs(4025) <= not a;
    outputs(4026) <= a xor b;
    outputs(4027) <= a xor b;
    outputs(4028) <= not (a and b);
    outputs(4029) <= not (a or b);
    outputs(4030) <= a xor b;
    outputs(4031) <= not (a xor b);
    outputs(4032) <= b and not a;
    outputs(4033) <= b;
    outputs(4034) <= not (a or b);
    outputs(4035) <= a xor b;
    outputs(4036) <= a and not b;
    outputs(4037) <= a;
    outputs(4038) <= b;
    outputs(4039) <= a and not b;
    outputs(4040) <= a and b;
    outputs(4041) <= a and b;
    outputs(4042) <= not (a or b);
    outputs(4043) <= a;
    outputs(4044) <= not (a and b);
    outputs(4045) <= not a or b;
    outputs(4046) <= a xor b;
    outputs(4047) <= b;
    outputs(4048) <= a;
    outputs(4049) <= b and not a;
    outputs(4050) <= not a or b;
    outputs(4051) <= not (a or b);
    outputs(4052) <= a and not b;
    outputs(4053) <= not b;
    outputs(4054) <= a and not b;
    outputs(4055) <= a and b;
    outputs(4056) <= a;
    outputs(4057) <= a and not b;
    outputs(4058) <= b and not a;
    outputs(4059) <= not a or b;
    outputs(4060) <= b;
    outputs(4061) <= a;
    outputs(4062) <= not a;
    outputs(4063) <= a and not b;
    outputs(4064) <= a;
    outputs(4065) <= b and not a;
    outputs(4066) <= a;
    outputs(4067) <= not (a xor b);
    outputs(4068) <= not a or b;
    outputs(4069) <= not (a and b);
    outputs(4070) <= not b or a;
    outputs(4071) <= b;
    outputs(4072) <= not b;
    outputs(4073) <= b;
    outputs(4074) <= a and not b;
    outputs(4075) <= b and not a;
    outputs(4076) <= a xor b;
    outputs(4077) <= b;
    outputs(4078) <= a and b;
    outputs(4079) <= b;
    outputs(4080) <= not (a or b);
    outputs(4081) <= not a or b;
    outputs(4082) <= a xor b;
    outputs(4083) <= a;
    outputs(4084) <= b;
    outputs(4085) <= not a or b;
    outputs(4086) <= b;
    outputs(4087) <= a;
    outputs(4088) <= b and not a;
    outputs(4089) <= a xor b;
    outputs(4090) <= a;
    outputs(4091) <= a xor b;
    outputs(4092) <= not b or a;
    outputs(4093) <= a and b;
    outputs(4094) <= not a;
    outputs(4095) <= not (a or b);
    outputs(4096) <= a xor b;
    outputs(4097) <= a;
    outputs(4098) <= b and not a;
    outputs(4099) <= not (a or b);
    outputs(4100) <= a and b;
    outputs(4101) <= not a;
    outputs(4102) <= a and not b;
    outputs(4103) <= a xor b;
    outputs(4104) <= not b;
    outputs(4105) <= not (a xor b);
    outputs(4106) <= not b or a;
    outputs(4107) <= not b;
    outputs(4108) <= a xor b;
    outputs(4109) <= b;
    outputs(4110) <= not a;
    outputs(4111) <= a;
    outputs(4112) <= b;
    outputs(4113) <= a;
    outputs(4114) <= b and not a;
    outputs(4115) <= b;
    outputs(4116) <= a or b;
    outputs(4117) <= a or b;
    outputs(4118) <= not b;
    outputs(4119) <= not a;
    outputs(4120) <= b;
    outputs(4121) <= a xor b;
    outputs(4122) <= b;
    outputs(4123) <= b;
    outputs(4124) <= not b or a;
    outputs(4125) <= a;
    outputs(4126) <= a and b;
    outputs(4127) <= a;
    outputs(4128) <= not (a xor b);
    outputs(4129) <= not b;
    outputs(4130) <= not b;
    outputs(4131) <= a and b;
    outputs(4132) <= a xor b;
    outputs(4133) <= a or b;
    outputs(4134) <= a and b;
    outputs(4135) <= not a or b;
    outputs(4136) <= not b;
    outputs(4137) <= a and b;
    outputs(4138) <= a;
    outputs(4139) <= a and b;
    outputs(4140) <= not b;
    outputs(4141) <= not a or b;
    outputs(4142) <= b;
    outputs(4143) <= not (a or b);
    outputs(4144) <= b;
    outputs(4145) <= b and not a;
    outputs(4146) <= not a;
    outputs(4147) <= b;
    outputs(4148) <= not a;
    outputs(4149) <= b;
    outputs(4150) <= not a;
    outputs(4151) <= b;
    outputs(4152) <= a and not b;
    outputs(4153) <= a and not b;
    outputs(4154) <= not (a and b);
    outputs(4155) <= a and not b;
    outputs(4156) <= not a;
    outputs(4157) <= a xor b;
    outputs(4158) <= a and not b;
    outputs(4159) <= b;
    outputs(4160) <= not b;
    outputs(4161) <= not a;
    outputs(4162) <= a and not b;
    outputs(4163) <= not a;
    outputs(4164) <= a xor b;
    outputs(4165) <= b;
    outputs(4166) <= a xor b;
    outputs(4167) <= not a;
    outputs(4168) <= not a;
    outputs(4169) <= a or b;
    outputs(4170) <= a;
    outputs(4171) <= b;
    outputs(4172) <= a xor b;
    outputs(4173) <= a and b;
    outputs(4174) <= a xor b;
    outputs(4175) <= not b;
    outputs(4176) <= not a;
    outputs(4177) <= b and not a;
    outputs(4178) <= not a;
    outputs(4179) <= b;
    outputs(4180) <= a;
    outputs(4181) <= a;
    outputs(4182) <= not b or a;
    outputs(4183) <= not a or b;
    outputs(4184) <= a;
    outputs(4185) <= not (a and b);
    outputs(4186) <= b;
    outputs(4187) <= not b or a;
    outputs(4188) <= a and b;
    outputs(4189) <= a;
    outputs(4190) <= a;
    outputs(4191) <= b;
    outputs(4192) <= not a or b;
    outputs(4193) <= a and not b;
    outputs(4194) <= not b;
    outputs(4195) <= not b;
    outputs(4196) <= not (a or b);
    outputs(4197) <= a and b;
    outputs(4198) <= not b or a;
    outputs(4199) <= a xor b;
    outputs(4200) <= not a or b;
    outputs(4201) <= not b;
    outputs(4202) <= a;
    outputs(4203) <= not (a or b);
    outputs(4204) <= a;
    outputs(4205) <= not (a xor b);
    outputs(4206) <= not (a xor b);
    outputs(4207) <= not b;
    outputs(4208) <= a and b;
    outputs(4209) <= not (a xor b);
    outputs(4210) <= a;
    outputs(4211) <= not (a xor b);
    outputs(4212) <= not a;
    outputs(4213) <= a;
    outputs(4214) <= not b;
    outputs(4215) <= b;
    outputs(4216) <= a and b;
    outputs(4217) <= a and b;
    outputs(4218) <= not (a or b);
    outputs(4219) <= b;
    outputs(4220) <= b and not a;
    outputs(4221) <= b;
    outputs(4222) <= not b or a;
    outputs(4223) <= b;
    outputs(4224) <= not (a xor b);
    outputs(4225) <= not a;
    outputs(4226) <= b;
    outputs(4227) <= b;
    outputs(4228) <= not (a and b);
    outputs(4229) <= not a;
    outputs(4230) <= b;
    outputs(4231) <= not a;
    outputs(4232) <= a or b;
    outputs(4233) <= not b;
    outputs(4234) <= a;
    outputs(4235) <= a or b;
    outputs(4236) <= not b;
    outputs(4237) <= not a;
    outputs(4238) <= a xor b;
    outputs(4239) <= a xor b;
    outputs(4240) <= b and not a;
    outputs(4241) <= a and b;
    outputs(4242) <= a and b;
    outputs(4243) <= not (a or b);
    outputs(4244) <= not (a xor b);
    outputs(4245) <= a and b;
    outputs(4246) <= a;
    outputs(4247) <= not b;
    outputs(4248) <= not (a xor b);
    outputs(4249) <= a and b;
    outputs(4250) <= b;
    outputs(4251) <= a and b;
    outputs(4252) <= not (a or b);
    outputs(4253) <= not (a or b);
    outputs(4254) <= not (a xor b);
    outputs(4255) <= not b;
    outputs(4256) <= not (a or b);
    outputs(4257) <= not (a or b);
    outputs(4258) <= a and not b;
    outputs(4259) <= not b or a;
    outputs(4260) <= not b;
    outputs(4261) <= a and not b;
    outputs(4262) <= not b;
    outputs(4263) <= not (a and b);
    outputs(4264) <= not b;
    outputs(4265) <= a and b;
    outputs(4266) <= a;
    outputs(4267) <= not b;
    outputs(4268) <= not (a or b);
    outputs(4269) <= b and not a;
    outputs(4270) <= a and not b;
    outputs(4271) <= not a;
    outputs(4272) <= not (a xor b);
    outputs(4273) <= not a or b;
    outputs(4274) <= not b;
    outputs(4275) <= not a;
    outputs(4276) <= a xor b;
    outputs(4277) <= a;
    outputs(4278) <= a and not b;
    outputs(4279) <= not (a or b);
    outputs(4280) <= not (a and b);
    outputs(4281) <= b;
    outputs(4282) <= not a or b;
    outputs(4283) <= not a or b;
    outputs(4284) <= not a;
    outputs(4285) <= a and b;
    outputs(4286) <= a;
    outputs(4287) <= not (a xor b);
    outputs(4288) <= a;
    outputs(4289) <= b;
    outputs(4290) <= b;
    outputs(4291) <= not b;
    outputs(4292) <= a;
    outputs(4293) <= not b;
    outputs(4294) <= a xor b;
    outputs(4295) <= a or b;
    outputs(4296) <= a;
    outputs(4297) <= a and b;
    outputs(4298) <= b;
    outputs(4299) <= not b or a;
    outputs(4300) <= a and not b;
    outputs(4301) <= a xor b;
    outputs(4302) <= not a or b;
    outputs(4303) <= not (a xor b);
    outputs(4304) <= a;
    outputs(4305) <= not a;
    outputs(4306) <= b;
    outputs(4307) <= not b or a;
    outputs(4308) <= a;
    outputs(4309) <= a;
    outputs(4310) <= b;
    outputs(4311) <= a and b;
    outputs(4312) <= not (a xor b);
    outputs(4313) <= a or b;
    outputs(4314) <= a and not b;
    outputs(4315) <= not b;
    outputs(4316) <= a and not b;
    outputs(4317) <= a xor b;
    outputs(4318) <= a;
    outputs(4319) <= not a or b;
    outputs(4320) <= b and not a;
    outputs(4321) <= not a;
    outputs(4322) <= not a;
    outputs(4323) <= a xor b;
    outputs(4324) <= not b;
    outputs(4325) <= b and not a;
    outputs(4326) <= not a;
    outputs(4327) <= a;
    outputs(4328) <= b;
    outputs(4329) <= b;
    outputs(4330) <= not a;
    outputs(4331) <= not b;
    outputs(4332) <= not (a or b);
    outputs(4333) <= not a;
    outputs(4334) <= a or b;
    outputs(4335) <= not a;
    outputs(4336) <= a xor b;
    outputs(4337) <= a;
    outputs(4338) <= not b;
    outputs(4339) <= not a;
    outputs(4340) <= not b;
    outputs(4341) <= b;
    outputs(4342) <= a or b;
    outputs(4343) <= a or b;
    outputs(4344) <= a and not b;
    outputs(4345) <= b;
    outputs(4346) <= b;
    outputs(4347) <= not a or b;
    outputs(4348) <= b;
    outputs(4349) <= not (a xor b);
    outputs(4350) <= a or b;
    outputs(4351) <= not b;
    outputs(4352) <= not (a and b);
    outputs(4353) <= not a;
    outputs(4354) <= not (a or b);
    outputs(4355) <= a xor b;
    outputs(4356) <= b and not a;
    outputs(4357) <= b;
    outputs(4358) <= not a;
    outputs(4359) <= a and b;
    outputs(4360) <= not a;
    outputs(4361) <= not (a and b);
    outputs(4362) <= not (a xor b);
    outputs(4363) <= a;
    outputs(4364) <= b;
    outputs(4365) <= not a;
    outputs(4366) <= b;
    outputs(4367) <= not b;
    outputs(4368) <= a xor b;
    outputs(4369) <= not (a xor b);
    outputs(4370) <= b and not a;
    outputs(4371) <= a;
    outputs(4372) <= a xor b;
    outputs(4373) <= a xor b;
    outputs(4374) <= a and b;
    outputs(4375) <= a;
    outputs(4376) <= not b;
    outputs(4377) <= not (a xor b);
    outputs(4378) <= not b;
    outputs(4379) <= a;
    outputs(4380) <= not a or b;
    outputs(4381) <= b and not a;
    outputs(4382) <= not (a xor b);
    outputs(4383) <= not a or b;
    outputs(4384) <= b and not a;
    outputs(4385) <= a and b;
    outputs(4386) <= a and b;
    outputs(4387) <= b and not a;
    outputs(4388) <= a;
    outputs(4389) <= a;
    outputs(4390) <= not (a xor b);
    outputs(4391) <= b;
    outputs(4392) <= not (a or b);
    outputs(4393) <= a xor b;
    outputs(4394) <= not (a xor b);
    outputs(4395) <= not b;
    outputs(4396) <= not a or b;
    outputs(4397) <= not (a xor b);
    outputs(4398) <= a and b;
    outputs(4399) <= a and b;
    outputs(4400) <= a or b;
    outputs(4401) <= not (a or b);
    outputs(4402) <= not (a or b);
    outputs(4403) <= not b;
    outputs(4404) <= a and not b;
    outputs(4405) <= not b;
    outputs(4406) <= b;
    outputs(4407) <= b and not a;
    outputs(4408) <= not (a and b);
    outputs(4409) <= not b;
    outputs(4410) <= not b or a;
    outputs(4411) <= not b;
    outputs(4412) <= b;
    outputs(4413) <= not a;
    outputs(4414) <= not a;
    outputs(4415) <= not (a and b);
    outputs(4416) <= a;
    outputs(4417) <= not b or a;
    outputs(4418) <= a and not b;
    outputs(4419) <= a and not b;
    outputs(4420) <= not (a xor b);
    outputs(4421) <= not (a or b);
    outputs(4422) <= a;
    outputs(4423) <= a xor b;
    outputs(4424) <= not a or b;
    outputs(4425) <= not (a or b);
    outputs(4426) <= b;
    outputs(4427) <= not (a xor b);
    outputs(4428) <= not (a and b);
    outputs(4429) <= a or b;
    outputs(4430) <= a and not b;
    outputs(4431) <= not a;
    outputs(4432) <= not (a or b);
    outputs(4433) <= b and not a;
    outputs(4434) <= b;
    outputs(4435) <= a xor b;
    outputs(4436) <= not (a xor b);
    outputs(4437) <= not (a and b);
    outputs(4438) <= not a;
    outputs(4439) <= a;
    outputs(4440) <= not b;
    outputs(4441) <= not (a or b);
    outputs(4442) <= not (a xor b);
    outputs(4443) <= a xor b;
    outputs(4444) <= a xor b;
    outputs(4445) <= b;
    outputs(4446) <= b and not a;
    outputs(4447) <= not a;
    outputs(4448) <= b;
    outputs(4449) <= a xor b;
    outputs(4450) <= not (a or b);
    outputs(4451) <= a and b;
    outputs(4452) <= not b;
    outputs(4453) <= b and not a;
    outputs(4454) <= b;
    outputs(4455) <= not b;
    outputs(4456) <= a;
    outputs(4457) <= a and b;
    outputs(4458) <= not (a or b);
    outputs(4459) <= a;
    outputs(4460) <= not a;
    outputs(4461) <= a and not b;
    outputs(4462) <= a and b;
    outputs(4463) <= not (a xor b);
    outputs(4464) <= not (a xor b);
    outputs(4465) <= not b;
    outputs(4466) <= not (a xor b);
    outputs(4467) <= not a;
    outputs(4468) <= not (a xor b);
    outputs(4469) <= a and b;
    outputs(4470) <= not (a xor b);
    outputs(4471) <= b and not a;
    outputs(4472) <= a;
    outputs(4473) <= not (a xor b);
    outputs(4474) <= b and not a;
    outputs(4475) <= not (a and b);
    outputs(4476) <= a and not b;
    outputs(4477) <= not b;
    outputs(4478) <= a;
    outputs(4479) <= a or b;
    outputs(4480) <= not b or a;
    outputs(4481) <= b;
    outputs(4482) <= a xor b;
    outputs(4483) <= b and not a;
    outputs(4484) <= a and b;
    outputs(4485) <= not (a or b);
    outputs(4486) <= not a;
    outputs(4487) <= not (a xor b);
    outputs(4488) <= a and b;
    outputs(4489) <= b;
    outputs(4490) <= not a;
    outputs(4491) <= not (a xor b);
    outputs(4492) <= a xor b;
    outputs(4493) <= a and not b;
    outputs(4494) <= not a;
    outputs(4495) <= not a;
    outputs(4496) <= b and not a;
    outputs(4497) <= not a or b;
    outputs(4498) <= a xor b;
    outputs(4499) <= b and not a;
    outputs(4500) <= b;
    outputs(4501) <= not (a or b);
    outputs(4502) <= a and b;
    outputs(4503) <= b;
    outputs(4504) <= a or b;
    outputs(4505) <= not a or b;
    outputs(4506) <= a xor b;
    outputs(4507) <= a xor b;
    outputs(4508) <= not (a xor b);
    outputs(4509) <= a;
    outputs(4510) <= a xor b;
    outputs(4511) <= a and not b;
    outputs(4512) <= not b;
    outputs(4513) <= a and b;
    outputs(4514) <= b;
    outputs(4515) <= not (a or b);
    outputs(4516) <= a and not b;
    outputs(4517) <= b and not a;
    outputs(4518) <= a;
    outputs(4519) <= a xor b;
    outputs(4520) <= a and not b;
    outputs(4521) <= a;
    outputs(4522) <= not (a and b);
    outputs(4523) <= not (a and b);
    outputs(4524) <= not (a or b);
    outputs(4525) <= not b;
    outputs(4526) <= not a;
    outputs(4527) <= a xor b;
    outputs(4528) <= a;
    outputs(4529) <= a and not b;
    outputs(4530) <= not (a or b);
    outputs(4531) <= not (a xor b);
    outputs(4532) <= not (a xor b);
    outputs(4533) <= a;
    outputs(4534) <= not a;
    outputs(4535) <= not b;
    outputs(4536) <= a and not b;
    outputs(4537) <= not b;
    outputs(4538) <= not (a xor b);
    outputs(4539) <= a or b;
    outputs(4540) <= not (a or b);
    outputs(4541) <= not b;
    outputs(4542) <= not (a or b);
    outputs(4543) <= a and b;
    outputs(4544) <= b and not a;
    outputs(4545) <= a and b;
    outputs(4546) <= a;
    outputs(4547) <= a and not b;
    outputs(4548) <= not (a and b);
    outputs(4549) <= a;
    outputs(4550) <= a xor b;
    outputs(4551) <= not (a xor b);
    outputs(4552) <= a;
    outputs(4553) <= not b;
    outputs(4554) <= not b or a;
    outputs(4555) <= not (a and b);
    outputs(4556) <= a xor b;
    outputs(4557) <= not (a xor b);
    outputs(4558) <= b and not a;
    outputs(4559) <= not a or b;
    outputs(4560) <= a xor b;
    outputs(4561) <= a;
    outputs(4562) <= a xor b;
    outputs(4563) <= not a;
    outputs(4564) <= a or b;
    outputs(4565) <= b;
    outputs(4566) <= b and not a;
    outputs(4567) <= a xor b;
    outputs(4568) <= not (a xor b);
    outputs(4569) <= a xor b;
    outputs(4570) <= not a;
    outputs(4571) <= a and b;
    outputs(4572) <= a and b;
    outputs(4573) <= a xor b;
    outputs(4574) <= not b;
    outputs(4575) <= not a or b;
    outputs(4576) <= b and not a;
    outputs(4577) <= not (a or b);
    outputs(4578) <= a;
    outputs(4579) <= not a or b;
    outputs(4580) <= not b;
    outputs(4581) <= a;
    outputs(4582) <= b and not a;
    outputs(4583) <= b and not a;
    outputs(4584) <= a xor b;
    outputs(4585) <= a and b;
    outputs(4586) <= a xor b;
    outputs(4587) <= not b or a;
    outputs(4588) <= a;
    outputs(4589) <= a xor b;
    outputs(4590) <= b and not a;
    outputs(4591) <= not b;
    outputs(4592) <= not (a xor b);
    outputs(4593) <= b and not a;
    outputs(4594) <= a or b;
    outputs(4595) <= b;
    outputs(4596) <= not a;
    outputs(4597) <= a and not b;
    outputs(4598) <= not a or b;
    outputs(4599) <= b and not a;
    outputs(4600) <= a xor b;
    outputs(4601) <= a xor b;
    outputs(4602) <= not b or a;
    outputs(4603) <= not a;
    outputs(4604) <= a;
    outputs(4605) <= not a or b;
    outputs(4606) <= not a;
    outputs(4607) <= a or b;
    outputs(4608) <= not (a or b);
    outputs(4609) <= not (a xor b);
    outputs(4610) <= a and b;
    outputs(4611) <= a and b;
    outputs(4612) <= a and b;
    outputs(4613) <= b;
    outputs(4614) <= not (a or b);
    outputs(4615) <= a or b;
    outputs(4616) <= a and b;
    outputs(4617) <= b and not a;
    outputs(4618) <= a and not b;
    outputs(4619) <= b;
    outputs(4620) <= a and b;
    outputs(4621) <= b and not a;
    outputs(4622) <= not (a or b);
    outputs(4623) <= not (a or b);
    outputs(4624) <= b and not a;
    outputs(4625) <= a and b;
    outputs(4626) <= a and b;
    outputs(4627) <= not a;
    outputs(4628) <= not a;
    outputs(4629) <= not a;
    outputs(4630) <= a xor b;
    outputs(4631) <= a and not b;
    outputs(4632) <= a;
    outputs(4633) <= a and b;
    outputs(4634) <= a;
    outputs(4635) <= a and b;
    outputs(4636) <= a;
    outputs(4637) <= not (a xor b);
    outputs(4638) <= b;
    outputs(4639) <= not (a or b);
    outputs(4640) <= not (a xor b);
    outputs(4641) <= a and not b;
    outputs(4642) <= a or b;
    outputs(4643) <= not a;
    outputs(4644) <= a and b;
    outputs(4645) <= a xor b;
    outputs(4646) <= a;
    outputs(4647) <= a and b;
    outputs(4648) <= a xor b;
    outputs(4649) <= not b;
    outputs(4650) <= a and b;
    outputs(4651) <= a xor b;
    outputs(4652) <= a xor b;
    outputs(4653) <= b and not a;
    outputs(4654) <= not (a xor b);
    outputs(4655) <= b and not a;
    outputs(4656) <= a and b;
    outputs(4657) <= a and not b;
    outputs(4658) <= not (a xor b);
    outputs(4659) <= a and b;
    outputs(4660) <= b and not a;
    outputs(4661) <= a and b;
    outputs(4662) <= not (a xor b);
    outputs(4663) <= a xor b;
    outputs(4664) <= b and not a;
    outputs(4665) <= not b;
    outputs(4666) <= a and not b;
    outputs(4667) <= a;
    outputs(4668) <= a and b;
    outputs(4669) <= a xor b;
    outputs(4670) <= a and not b;
    outputs(4671) <= not b;
    outputs(4672) <= a and not b;
    outputs(4673) <= a and not b;
    outputs(4674) <= a and b;
    outputs(4675) <= a;
    outputs(4676) <= b and not a;
    outputs(4677) <= a;
    outputs(4678) <= a or b;
    outputs(4679) <= not a;
    outputs(4680) <= a;
    outputs(4681) <= b and not a;
    outputs(4682) <= a xor b;
    outputs(4683) <= a xor b;
    outputs(4684) <= a;
    outputs(4685) <= not a;
    outputs(4686) <= a and not b;
    outputs(4687) <= not a;
    outputs(4688) <= a and not b;
    outputs(4689) <= not (a or b);
    outputs(4690) <= b and not a;
    outputs(4691) <= not a;
    outputs(4692) <= not (a xor b);
    outputs(4693) <= not b;
    outputs(4694) <= a xor b;
    outputs(4695) <= b;
    outputs(4696) <= a and b;
    outputs(4697) <= not (a xor b);
    outputs(4698) <= b and not a;
    outputs(4699) <= not b or a;
    outputs(4700) <= a and not b;
    outputs(4701) <= a and not b;
    outputs(4702) <= not (a or b);
    outputs(4703) <= a and b;
    outputs(4704) <= b;
    outputs(4705) <= a;
    outputs(4706) <= a and not b;
    outputs(4707) <= b and not a;
    outputs(4708) <= a and not b;
    outputs(4709) <= a xor b;
    outputs(4710) <= not a;
    outputs(4711) <= b and not a;
    outputs(4712) <= b;
    outputs(4713) <= b and not a;
    outputs(4714) <= not a;
    outputs(4715) <= a;
    outputs(4716) <= b and not a;
    outputs(4717) <= not (a xor b);
    outputs(4718) <= not b;
    outputs(4719) <= not (a or b);
    outputs(4720) <= a or b;
    outputs(4721) <= not (a and b);
    outputs(4722) <= not b;
    outputs(4723) <= a and b;
    outputs(4724) <= b and not a;
    outputs(4725) <= a and b;
    outputs(4726) <= b;
    outputs(4727) <= not (a xor b);
    outputs(4728) <= not b;
    outputs(4729) <= a and b;
    outputs(4730) <= not (a xor b);
    outputs(4731) <= not b;
    outputs(4732) <= a and not b;
    outputs(4733) <= not (a xor b);
    outputs(4734) <= a xor b;
    outputs(4735) <= a and not b;
    outputs(4736) <= a xor b;
    outputs(4737) <= not a;
    outputs(4738) <= not (a and b);
    outputs(4739) <= a and not b;
    outputs(4740) <= a and b;
    outputs(4741) <= a xor b;
    outputs(4742) <= a and not b;
    outputs(4743) <= a xor b;
    outputs(4744) <= a xor b;
    outputs(4745) <= b and not a;
    outputs(4746) <= not b or a;
    outputs(4747) <= b and not a;
    outputs(4748) <= a and not b;
    outputs(4749) <= a and b;
    outputs(4750) <= a;
    outputs(4751) <= not (a or b);
    outputs(4752) <= a and b;
    outputs(4753) <= not a or b;
    outputs(4754) <= a and not b;
    outputs(4755) <= not b;
    outputs(4756) <= not b;
    outputs(4757) <= a;
    outputs(4758) <= not (a or b);
    outputs(4759) <= not (a or b);
    outputs(4760) <= a and b;
    outputs(4761) <= b and not a;
    outputs(4762) <= b and not a;
    outputs(4763) <= a;
    outputs(4764) <= a and b;
    outputs(4765) <= a and b;
    outputs(4766) <= b;
    outputs(4767) <= a and not b;
    outputs(4768) <= not (a or b);
    outputs(4769) <= b;
    outputs(4770) <= not (a xor b);
    outputs(4771) <= not (a or b);
    outputs(4772) <= not b;
    outputs(4773) <= b and not a;
    outputs(4774) <= a xor b;
    outputs(4775) <= a and not b;
    outputs(4776) <= a and not b;
    outputs(4777) <= a;
    outputs(4778) <= not (a or b);
    outputs(4779) <= not b;
    outputs(4780) <= not (a xor b);
    outputs(4781) <= not (a or b);
    outputs(4782) <= a xor b;
    outputs(4783) <= not a or b;
    outputs(4784) <= a and b;
    outputs(4785) <= not a;
    outputs(4786) <= a and not b;
    outputs(4787) <= a and not b;
    outputs(4788) <= b;
    outputs(4789) <= a;
    outputs(4790) <= not (a and b);
    outputs(4791) <= not (a or b);
    outputs(4792) <= not (a xor b);
    outputs(4793) <= b and not a;
    outputs(4794) <= a and b;
    outputs(4795) <= not (a and b);
    outputs(4796) <= not a or b;
    outputs(4797) <= a and not b;
    outputs(4798) <= not a;
    outputs(4799) <= a and b;
    outputs(4800) <= not a;
    outputs(4801) <= a;
    outputs(4802) <= a and not b;
    outputs(4803) <= not a;
    outputs(4804) <= not (a or b);
    outputs(4805) <= not a;
    outputs(4806) <= a and not b;
    outputs(4807) <= not (a or b);
    outputs(4808) <= not b;
    outputs(4809) <= not (a or b);
    outputs(4810) <= not a;
    outputs(4811) <= not (a or b);
    outputs(4812) <= not a;
    outputs(4813) <= not b;
    outputs(4814) <= not (a xor b);
    outputs(4815) <= a and not b;
    outputs(4816) <= not (a or b);
    outputs(4817) <= b and not a;
    outputs(4818) <= b;
    outputs(4819) <= not a;
    outputs(4820) <= b and not a;
    outputs(4821) <= a and b;
    outputs(4822) <= b;
    outputs(4823) <= not (a xor b);
    outputs(4824) <= not a;
    outputs(4825) <= a or b;
    outputs(4826) <= a xor b;
    outputs(4827) <= a and not b;
    outputs(4828) <= a and not b;
    outputs(4829) <= not (a xor b);
    outputs(4830) <= not a;
    outputs(4831) <= a and b;
    outputs(4832) <= a or b;
    outputs(4833) <= not (a or b);
    outputs(4834) <= not a;
    outputs(4835) <= a;
    outputs(4836) <= a;
    outputs(4837) <= not b;
    outputs(4838) <= a and b;
    outputs(4839) <= '0';
    outputs(4840) <= a and not b;
    outputs(4841) <= not (a or b);
    outputs(4842) <= not b;
    outputs(4843) <= not (a xor b);
    outputs(4844) <= not (a or b);
    outputs(4845) <= a and not b;
    outputs(4846) <= b;
    outputs(4847) <= b;
    outputs(4848) <= not b;
    outputs(4849) <= a xor b;
    outputs(4850) <= a and not b;
    outputs(4851) <= a and not b;
    outputs(4852) <= a;
    outputs(4853) <= b;
    outputs(4854) <= a and not b;
    outputs(4855) <= not a;
    outputs(4856) <= b and not a;
    outputs(4857) <= b and not a;
    outputs(4858) <= a and b;
    outputs(4859) <= a and not b;
    outputs(4860) <= not b;
    outputs(4861) <= not b;
    outputs(4862) <= a;
    outputs(4863) <= b;
    outputs(4864) <= a and b;
    outputs(4865) <= not b or a;
    outputs(4866) <= not b or a;
    outputs(4867) <= not (a xor b);
    outputs(4868) <= not b;
    outputs(4869) <= not a or b;
    outputs(4870) <= b and not a;
    outputs(4871) <= a xor b;
    outputs(4872) <= not (a or b);
    outputs(4873) <= a xor b;
    outputs(4874) <= a and b;
    outputs(4875) <= a and b;
    outputs(4876) <= not a or b;
    outputs(4877) <= a xor b;
    outputs(4878) <= not a;
    outputs(4879) <= a;
    outputs(4880) <= b;
    outputs(4881) <= a xor b;
    outputs(4882) <= b and not a;
    outputs(4883) <= not a or b;
    outputs(4884) <= not (a xor b);
    outputs(4885) <= not a or b;
    outputs(4886) <= b;
    outputs(4887) <= not (a xor b);
    outputs(4888) <= a and not b;
    outputs(4889) <= not b;
    outputs(4890) <= a and not b;
    outputs(4891) <= a and b;
    outputs(4892) <= b;
    outputs(4893) <= not a or b;
    outputs(4894) <= a;
    outputs(4895) <= not (a and b);
    outputs(4896) <= a;
    outputs(4897) <= a and b;
    outputs(4898) <= b;
    outputs(4899) <= not (a or b);
    outputs(4900) <= b;
    outputs(4901) <= a;
    outputs(4902) <= not b;
    outputs(4903) <= a and not b;
    outputs(4904) <= b and not a;
    outputs(4905) <= not a;
    outputs(4906) <= not (a and b);
    outputs(4907) <= not a;
    outputs(4908) <= not (a xor b);
    outputs(4909) <= a xor b;
    outputs(4910) <= a xor b;
    outputs(4911) <= a and not b;
    outputs(4912) <= not b;
    outputs(4913) <= b and not a;
    outputs(4914) <= not (a or b);
    outputs(4915) <= not (a xor b);
    outputs(4916) <= not a;
    outputs(4917) <= not b or a;
    outputs(4918) <= a and not b;
    outputs(4919) <= not (a or b);
    outputs(4920) <= a xor b;
    outputs(4921) <= not a;
    outputs(4922) <= b;
    outputs(4923) <= a and not b;
    outputs(4924) <= a xor b;
    outputs(4925) <= a or b;
    outputs(4926) <= not (a xor b);
    outputs(4927) <= not (a or b);
    outputs(4928) <= b and not a;
    outputs(4929) <= b;
    outputs(4930) <= not b or a;
    outputs(4931) <= a and not b;
    outputs(4932) <= a and not b;
    outputs(4933) <= a;
    outputs(4934) <= not a;
    outputs(4935) <= a and b;
    outputs(4936) <= a xor b;
    outputs(4937) <= not b;
    outputs(4938) <= a and not b;
    outputs(4939) <= a xor b;
    outputs(4940) <= not b;
    outputs(4941) <= a;
    outputs(4942) <= a and not b;
    outputs(4943) <= not a or b;
    outputs(4944) <= not a;
    outputs(4945) <= b and not a;
    outputs(4946) <= a;
    outputs(4947) <= a and not b;
    outputs(4948) <= not a;
    outputs(4949) <= a and b;
    outputs(4950) <= a;
    outputs(4951) <= a;
    outputs(4952) <= b and not a;
    outputs(4953) <= a and b;
    outputs(4954) <= not b;
    outputs(4955) <= a or b;
    outputs(4956) <= a and b;
    outputs(4957) <= a and not b;
    outputs(4958) <= a and not b;
    outputs(4959) <= not b;
    outputs(4960) <= not (a xor b);
    outputs(4961) <= not a or b;
    outputs(4962) <= a xor b;
    outputs(4963) <= a and b;
    outputs(4964) <= a xor b;
    outputs(4965) <= not (a xor b);
    outputs(4966) <= b and not a;
    outputs(4967) <= not b or a;
    outputs(4968) <= a and not b;
    outputs(4969) <= not b or a;
    outputs(4970) <= not a;
    outputs(4971) <= not (a xor b);
    outputs(4972) <= a;
    outputs(4973) <= a xor b;
    outputs(4974) <= a and not b;
    outputs(4975) <= not b;
    outputs(4976) <= not a;
    outputs(4977) <= not b or a;
    outputs(4978) <= not a;
    outputs(4979) <= not b;
    outputs(4980) <= not b;
    outputs(4981) <= a and not b;
    outputs(4982) <= a or b;
    outputs(4983) <= not (a or b);
    outputs(4984) <= a;
    outputs(4985) <= b and not a;
    outputs(4986) <= not (a or b);
    outputs(4987) <= a;
    outputs(4988) <= not b;
    outputs(4989) <= a xor b;
    outputs(4990) <= a;
    outputs(4991) <= a and b;
    outputs(4992) <= a and b;
    outputs(4993) <= b;
    outputs(4994) <= b and not a;
    outputs(4995) <= not (a and b);
    outputs(4996) <= a and b;
    outputs(4997) <= a and not b;
    outputs(4998) <= a and not b;
    outputs(4999) <= not (a or b);
    outputs(5000) <= b;
    outputs(5001) <= b and not a;
    outputs(5002) <= a and b;
    outputs(5003) <= not (a or b);
    outputs(5004) <= b and not a;
    outputs(5005) <= not (a xor b);
    outputs(5006) <= b and not a;
    outputs(5007) <= b;
    outputs(5008) <= a or b;
    outputs(5009) <= not (a xor b);
    outputs(5010) <= not (a xor b);
    outputs(5011) <= b;
    outputs(5012) <= a and not b;
    outputs(5013) <= not (a and b);
    outputs(5014) <= not (a xor b);
    outputs(5015) <= not (a or b);
    outputs(5016) <= not b;
    outputs(5017) <= not a;
    outputs(5018) <= b;
    outputs(5019) <= not (a xor b);
    outputs(5020) <= not b;
    outputs(5021) <= not (a or b);
    outputs(5022) <= a or b;
    outputs(5023) <= a xor b;
    outputs(5024) <= a;
    outputs(5025) <= b and not a;
    outputs(5026) <= not b;
    outputs(5027) <= b;
    outputs(5028) <= not b or a;
    outputs(5029) <= not b;
    outputs(5030) <= a xor b;
    outputs(5031) <= a or b;
    outputs(5032) <= not a or b;
    outputs(5033) <= a;
    outputs(5034) <= not a;
    outputs(5035) <= b;
    outputs(5036) <= a or b;
    outputs(5037) <= b;
    outputs(5038) <= b and not a;
    outputs(5039) <= not (a xor b);
    outputs(5040) <= not a;
    outputs(5041) <= a and b;
    outputs(5042) <= not (a and b);
    outputs(5043) <= a and not b;
    outputs(5044) <= a;
    outputs(5045) <= a and not b;
    outputs(5046) <= a and not b;
    outputs(5047) <= b and not a;
    outputs(5048) <= not b;
    outputs(5049) <= not a or b;
    outputs(5050) <= a and b;
    outputs(5051) <= not (a xor b);
    outputs(5052) <= a;
    outputs(5053) <= not a or b;
    outputs(5054) <= not a;
    outputs(5055) <= a and b;
    outputs(5056) <= a;
    outputs(5057) <= b and not a;
    outputs(5058) <= a and not b;
    outputs(5059) <= a;
    outputs(5060) <= a and b;
    outputs(5061) <= b and not a;
    outputs(5062) <= a;
    outputs(5063) <= not (a or b);
    outputs(5064) <= not (a or b);
    outputs(5065) <= a;
    outputs(5066) <= a and not b;
    outputs(5067) <= not b or a;
    outputs(5068) <= not b;
    outputs(5069) <= a and not b;
    outputs(5070) <= a and b;
    outputs(5071) <= a xor b;
    outputs(5072) <= b and not a;
    outputs(5073) <= a xor b;
    outputs(5074) <= a xor b;
    outputs(5075) <= a and not b;
    outputs(5076) <= not (a or b);
    outputs(5077) <= a and b;
    outputs(5078) <= a and b;
    outputs(5079) <= not (a or b);
    outputs(5080) <= not a;
    outputs(5081) <= not (a and b);
    outputs(5082) <= not (a or b);
    outputs(5083) <= not b;
    outputs(5084) <= a xor b;
    outputs(5085) <= a and b;
    outputs(5086) <= not (a xor b);
    outputs(5087) <= b;
    outputs(5088) <= a;
    outputs(5089) <= a xor b;
    outputs(5090) <= a xor b;
    outputs(5091) <= not (a or b);
    outputs(5092) <= not a or b;
    outputs(5093) <= not b;
    outputs(5094) <= a xor b;
    outputs(5095) <= not (a or b);
    outputs(5096) <= b and not a;
    outputs(5097) <= b;
    outputs(5098) <= a and b;
    outputs(5099) <= not (a xor b);
    outputs(5100) <= not a;
    outputs(5101) <= b and not a;
    outputs(5102) <= b and not a;
    outputs(5103) <= a;
    outputs(5104) <= not b;
    outputs(5105) <= a and not b;
    outputs(5106) <= not a;
    outputs(5107) <= b;
    outputs(5108) <= b and not a;
    outputs(5109) <= a and not b;
    outputs(5110) <= not (a or b);
    outputs(5111) <= a xor b;
    outputs(5112) <= b and not a;
    outputs(5113) <= not (a and b);
    outputs(5114) <= not a or b;
    outputs(5115) <= not a;
    outputs(5116) <= not (a xor b);
    outputs(5117) <= not (a or b);
    outputs(5118) <= not (a xor b);
    outputs(5119) <= not a;
end Behavioral;
